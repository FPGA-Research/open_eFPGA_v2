magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect -170 4189 1721 5697
<< nwell >>
rect -250 22825 52 27807
rect 452 24950 958 25116
rect 452 23441 618 24950
rect 1692 23441 1858 24311
rect 452 23275 1858 23441
rect -250 22523 2297 22825
<< pwell >>
rect 170 27545 2976 27767
rect 170 23209 392 27545
rect 170 22987 2976 23209
rect 146 5057 1448 5279
rect 146 4163 368 5057
rect 1226 4163 1448 5057
<< mvpsubdiff >>
rect 196 27707 230 27741
rect 264 27707 299 27741
rect 333 27707 368 27741
rect 402 27707 437 27741
rect 471 27707 506 27741
rect 540 27707 575 27741
rect 609 27707 644 27741
rect 678 27707 713 27741
rect 747 27707 782 27741
rect 816 27707 851 27741
rect 885 27707 920 27741
rect 954 27707 988 27741
rect 1022 27707 1056 27741
rect 1090 27707 1124 27741
rect 1158 27707 1192 27741
rect 1226 27707 1260 27741
rect 1294 27707 1328 27741
rect 1362 27707 1396 27741
rect 1430 27707 1464 27741
rect 1498 27707 1532 27741
rect 1566 27707 1600 27741
rect 1634 27707 1668 27741
rect 1702 27707 1736 27741
rect 1770 27707 1804 27741
rect 1838 27707 1872 27741
rect 1906 27707 1940 27741
rect 1974 27707 2008 27741
rect 2042 27707 2076 27741
rect 2110 27707 2144 27741
rect 2178 27707 2212 27741
rect 2246 27707 2280 27741
rect 2314 27707 2348 27741
rect 2382 27707 2416 27741
rect 2450 27707 2484 27741
rect 2518 27707 2552 27741
rect 2586 27707 2620 27741
rect 2654 27707 2688 27741
rect 2722 27707 2756 27741
rect 2790 27707 2824 27741
rect 2858 27707 2892 27741
rect 2926 27707 2950 27741
rect 196 27673 2950 27707
rect 196 27639 264 27673
rect 298 27639 334 27673
rect 368 27639 404 27673
rect 438 27639 474 27673
rect 508 27639 544 27673
rect 578 27639 614 27673
rect 648 27639 684 27673
rect 718 27639 753 27673
rect 787 27639 822 27673
rect 856 27639 891 27673
rect 925 27639 960 27673
rect 994 27639 1029 27673
rect 1063 27639 1098 27673
rect 1132 27639 1167 27673
rect 1201 27639 1236 27673
rect 1270 27639 1305 27673
rect 1339 27639 1374 27673
rect 1408 27639 1443 27673
rect 1477 27639 1512 27673
rect 1546 27639 1581 27673
rect 1615 27639 1650 27673
rect 1684 27639 1719 27673
rect 1753 27639 1788 27673
rect 1822 27639 1857 27673
rect 1891 27639 1926 27673
rect 1960 27639 1995 27673
rect 2029 27639 2064 27673
rect 2098 27639 2133 27673
rect 2167 27639 2202 27673
rect 2236 27639 2271 27673
rect 2305 27639 2340 27673
rect 2374 27639 2409 27673
rect 2443 27639 2478 27673
rect 2512 27639 2547 27673
rect 2581 27639 2616 27673
rect 2650 27639 2685 27673
rect 2719 27639 2754 27673
rect 2788 27639 2823 27673
rect 2857 27639 2892 27673
rect 2926 27639 2950 27673
rect 196 27631 2950 27639
rect 230 27605 2950 27631
rect 230 27597 332 27605
rect 196 27586 332 27597
rect 196 27558 264 27586
rect 230 27552 264 27558
rect 298 27571 332 27586
rect 366 27571 402 27605
rect 436 27571 472 27605
rect 506 27571 542 27605
rect 576 27571 612 27605
rect 646 27571 682 27605
rect 716 27571 752 27605
rect 786 27571 822 27605
rect 856 27571 891 27605
rect 925 27571 960 27605
rect 994 27571 1029 27605
rect 1063 27571 1098 27605
rect 1132 27571 1167 27605
rect 1201 27571 1236 27605
rect 1270 27571 1305 27605
rect 1339 27571 1374 27605
rect 1408 27571 1443 27605
rect 1477 27571 1512 27605
rect 1546 27571 1581 27605
rect 1615 27571 1650 27605
rect 1684 27571 1719 27605
rect 1753 27571 1788 27605
rect 1822 27571 1857 27605
rect 1891 27571 1926 27605
rect 1960 27571 1995 27605
rect 2029 27571 2064 27605
rect 2098 27571 2133 27605
rect 2167 27571 2202 27605
rect 2236 27571 2271 27605
rect 2305 27571 2340 27605
rect 2374 27571 2409 27605
rect 2443 27571 2478 27605
rect 2512 27571 2547 27605
rect 2581 27571 2616 27605
rect 2650 27571 2685 27605
rect 2719 27571 2754 27605
rect 2788 27571 2823 27605
rect 2857 27571 2892 27605
rect 2926 27571 2950 27605
rect 298 27552 366 27571
rect 230 27524 366 27552
rect 196 27509 366 27524
rect 196 27499 332 27509
rect 196 27485 264 27499
rect 230 27465 264 27485
rect 298 27475 332 27499
rect 298 27465 366 27475
rect 230 27451 366 27465
rect 196 27412 366 27451
rect 230 27378 264 27412
rect 298 27378 332 27412
rect 196 27330 366 27378
rect 230 27296 264 27330
rect 298 27296 332 27330
rect 196 27261 366 27296
rect 230 27260 366 27261
rect 230 27227 264 27260
rect 196 27226 264 27227
rect 298 27226 332 27260
rect 196 27192 366 27226
rect 230 27190 366 27192
rect 230 27158 264 27190
rect 196 27156 264 27158
rect 298 27156 332 27190
rect 196 27123 366 27156
rect 230 27120 366 27123
rect 230 27089 264 27120
rect 196 27086 264 27089
rect 298 27086 332 27120
rect 196 27054 366 27086
rect 230 27050 366 27054
rect 230 27020 264 27050
rect 196 27016 264 27020
rect 298 27016 332 27050
rect 196 26985 366 27016
rect 230 26980 366 26985
rect 230 26951 264 26980
rect 196 26946 264 26951
rect 298 26946 332 26980
rect 196 26916 366 26946
rect 230 26910 366 26916
rect 230 26882 264 26910
rect 196 26876 264 26882
rect 298 26876 332 26910
rect 196 26847 366 26876
rect 230 26841 366 26847
rect 230 26813 264 26841
rect 196 26807 264 26813
rect 298 26840 366 26841
rect 298 26807 332 26840
rect 196 26806 332 26807
rect 196 26778 366 26806
rect 230 26772 366 26778
rect 230 26744 264 26772
rect 196 26738 264 26744
rect 298 26771 366 26772
rect 298 26738 332 26771
rect 196 26737 332 26738
rect 196 26709 366 26737
rect 230 26703 366 26709
rect 230 26675 264 26703
rect 196 26669 264 26675
rect 298 26702 366 26703
rect 298 26669 332 26702
rect 196 26668 332 26669
rect 196 26640 366 26668
rect 230 26634 366 26640
rect 230 26606 264 26634
rect 196 26600 264 26606
rect 298 26633 366 26634
rect 298 26600 332 26633
rect 196 26599 332 26600
rect 196 26571 366 26599
rect 230 26565 366 26571
rect 230 26537 264 26565
rect 196 26531 264 26537
rect 298 26564 366 26565
rect 298 26531 332 26564
rect 196 26530 332 26531
rect 196 26502 366 26530
rect 230 26496 366 26502
rect 230 26468 264 26496
rect 196 26462 264 26468
rect 298 26495 366 26496
rect 298 26462 332 26495
rect 196 26461 332 26462
rect 196 26433 366 26461
rect 230 26427 366 26433
rect 230 26399 264 26427
rect 196 26393 264 26399
rect 298 26426 366 26427
rect 298 26393 332 26426
rect 196 26392 332 26393
rect 196 26364 366 26392
rect 230 26358 366 26364
rect 230 26330 264 26358
rect 196 26324 264 26330
rect 298 26357 366 26358
rect 298 26324 332 26357
rect 196 26323 332 26324
rect 196 26295 366 26323
rect 230 26289 366 26295
rect 230 26261 264 26289
rect 196 26255 264 26261
rect 298 26288 366 26289
rect 298 26255 332 26288
rect 196 26254 332 26255
rect 196 26226 366 26254
rect 230 26220 366 26226
rect 230 26192 264 26220
rect 196 26186 264 26192
rect 298 26219 366 26220
rect 298 26186 332 26219
rect 196 26185 332 26186
rect 196 26157 366 26185
rect 230 26151 366 26157
rect 230 26123 264 26151
rect 196 26117 264 26123
rect 298 26150 366 26151
rect 298 26117 332 26150
rect 196 26116 332 26117
rect 196 26088 366 26116
rect 230 26082 366 26088
rect 230 26054 264 26082
rect 196 26048 264 26054
rect 298 26081 366 26082
rect 298 26048 332 26081
rect 196 26047 332 26048
rect 196 26019 366 26047
rect 230 26013 366 26019
rect 230 25985 264 26013
rect 196 25979 264 25985
rect 298 26012 366 26013
rect 298 25979 332 26012
rect 196 25978 332 25979
rect 196 25950 366 25978
rect 230 25944 366 25950
rect 230 25916 264 25944
rect 196 25910 264 25916
rect 298 25943 366 25944
rect 298 25910 332 25943
rect 196 25909 332 25910
rect 196 25881 366 25909
rect 230 25875 366 25881
rect 230 25847 264 25875
rect 196 25841 264 25847
rect 298 25874 366 25875
rect 298 25841 332 25874
rect 196 25840 332 25841
rect 196 25812 366 25840
rect 230 25806 366 25812
rect 230 25778 264 25806
rect 196 25772 264 25778
rect 298 25805 366 25806
rect 298 25772 332 25805
rect 196 25771 332 25772
rect 196 25743 366 25771
rect 230 25737 366 25743
rect 230 25709 264 25737
rect 196 25703 264 25709
rect 298 25736 366 25737
rect 298 25703 332 25736
rect 196 25702 332 25703
rect 196 25674 366 25702
rect 230 25668 366 25674
rect 230 25640 264 25668
rect 196 25634 264 25640
rect 298 25667 366 25668
rect 298 25634 332 25667
rect 196 25633 332 25634
rect 196 25605 366 25633
rect 230 25599 366 25605
rect 230 25571 264 25599
rect 196 25565 264 25571
rect 298 25598 366 25599
rect 298 25565 332 25598
rect 196 25564 332 25565
rect 196 25536 366 25564
rect 230 25530 366 25536
rect 230 25502 264 25530
rect 196 25496 264 25502
rect 298 25529 366 25530
rect 298 25496 332 25529
rect 196 25495 332 25496
rect 196 25467 366 25495
rect 230 25461 366 25467
rect 230 25433 264 25461
rect 196 25427 264 25433
rect 298 25460 366 25461
rect 298 25427 332 25460
rect 196 25426 332 25427
rect 196 25398 366 25426
rect 230 25392 366 25398
rect 230 25364 264 25392
rect 196 25358 264 25364
rect 298 25391 366 25392
rect 298 25358 332 25391
rect 196 25357 332 25358
rect 196 25329 366 25357
rect 230 25323 366 25329
rect 230 25295 264 25323
rect 196 25289 264 25295
rect 298 25322 366 25323
rect 298 25289 332 25322
rect 196 25288 332 25289
rect 196 25260 366 25288
rect 230 25254 366 25260
rect 230 25226 264 25254
rect 196 25220 264 25226
rect 298 25253 366 25254
rect 298 25220 332 25253
rect 196 25219 332 25220
rect 196 25191 366 25219
rect 230 25185 366 25191
rect 230 25157 264 25185
rect 196 25151 264 25157
rect 298 25184 366 25185
rect 298 25151 332 25184
rect 196 25150 332 25151
rect 196 25122 366 25150
rect 230 25116 366 25122
rect 230 25088 264 25116
rect 196 25082 264 25088
rect 298 25115 366 25116
rect 298 25082 332 25115
rect 196 25081 332 25082
rect 196 25053 366 25081
rect 230 25047 366 25053
rect 230 25019 264 25047
rect 196 25013 264 25019
rect 298 25046 366 25047
rect 298 25013 332 25046
rect 196 25012 332 25013
rect 196 24985 366 25012
rect 230 24978 366 24985
rect 230 24951 264 24978
rect 196 24944 264 24951
rect 298 24977 366 24978
rect 298 24944 332 24977
rect 196 24943 332 24944
rect 196 24917 366 24943
rect 230 24909 366 24917
rect 230 24883 264 24909
rect 196 24875 264 24883
rect 298 24908 366 24909
rect 298 24875 332 24908
rect 196 24874 332 24875
rect 196 24849 366 24874
rect 230 24840 366 24849
rect 230 24815 264 24840
rect 196 24806 264 24815
rect 298 24839 366 24840
rect 298 24806 332 24839
rect 196 24805 332 24806
rect 196 24781 366 24805
rect 230 24771 366 24781
rect 230 24747 264 24771
rect 196 24737 264 24747
rect 298 24770 366 24771
rect 298 24737 332 24770
rect 196 24736 332 24737
rect 196 24713 366 24736
rect 230 24702 366 24713
rect 230 24679 264 24702
rect 196 24668 264 24679
rect 298 24701 366 24702
rect 298 24668 332 24701
rect 196 24667 332 24668
rect 196 24645 366 24667
rect 230 24633 366 24645
rect 230 24611 264 24633
rect 196 24599 264 24611
rect 298 24632 366 24633
rect 298 24599 332 24632
rect 196 24598 332 24599
rect 196 24577 366 24598
rect 230 24564 366 24577
rect 230 24543 264 24564
rect 196 24530 264 24543
rect 298 24563 366 24564
rect 298 24530 332 24563
rect 196 24529 332 24530
rect 196 24509 366 24529
rect 230 24495 366 24509
rect 230 24475 264 24495
rect 196 24461 264 24475
rect 298 24494 366 24495
rect 298 24461 332 24494
rect 196 24460 332 24461
rect 196 24441 366 24460
rect 230 24426 366 24441
rect 230 24407 264 24426
rect 196 24392 264 24407
rect 298 24425 366 24426
rect 298 24392 332 24425
rect 196 24391 332 24392
rect 196 24373 366 24391
rect 230 24357 366 24373
rect 230 24339 264 24357
rect 196 24323 264 24339
rect 298 24356 366 24357
rect 298 24323 332 24356
rect 196 24322 332 24323
rect 196 24305 366 24322
rect 230 24288 366 24305
rect 230 24271 264 24288
rect 196 24254 264 24271
rect 298 24287 366 24288
rect 298 24254 332 24287
rect 196 24253 332 24254
rect 196 24237 366 24253
rect 230 24219 366 24237
rect 230 24203 264 24219
rect 196 24185 264 24203
rect 298 24218 366 24219
rect 298 24185 332 24218
rect 196 24184 332 24185
rect 196 24169 366 24184
rect 230 24150 366 24169
rect 230 24135 264 24150
rect 196 24116 264 24135
rect 298 24149 366 24150
rect 298 24116 332 24149
rect 196 24115 332 24116
rect 196 24101 366 24115
rect 230 24081 366 24101
rect 230 24067 264 24081
rect 196 24047 264 24067
rect 298 24080 366 24081
rect 298 24047 332 24080
rect 196 24046 332 24047
rect 196 24033 366 24046
rect 230 24012 366 24033
rect 230 23999 264 24012
rect 196 23978 264 23999
rect 298 24011 366 24012
rect 298 23978 332 24011
rect 196 23977 332 23978
rect 196 23965 366 23977
rect 230 23943 366 23965
rect 230 23931 264 23943
rect 196 23909 264 23931
rect 298 23942 366 23943
rect 298 23909 332 23942
rect 196 23908 332 23909
rect 196 23897 366 23908
rect 230 23874 366 23897
rect 230 23863 264 23874
rect 196 23840 264 23863
rect 298 23873 366 23874
rect 298 23840 332 23873
rect 196 23839 332 23840
rect 196 23829 366 23839
rect 230 23805 366 23829
rect 230 23795 264 23805
rect 196 23771 264 23795
rect 298 23804 366 23805
rect 298 23771 332 23804
rect 196 23770 332 23771
rect 196 23761 366 23770
rect 230 23736 366 23761
rect 230 23727 264 23736
rect 196 23702 264 23727
rect 298 23735 366 23736
rect 298 23702 332 23735
rect 196 23701 332 23702
rect 196 23693 366 23701
rect 230 23667 366 23693
rect 230 23659 264 23667
rect 196 23633 264 23659
rect 298 23666 366 23667
rect 298 23633 332 23666
rect 196 23632 332 23633
rect 196 23625 366 23632
rect 230 23598 366 23625
rect 230 23591 264 23598
rect 196 23564 264 23591
rect 298 23597 366 23598
rect 298 23564 332 23597
rect 196 23563 332 23564
rect 196 23557 366 23563
rect 230 23529 366 23557
rect 230 23523 264 23529
rect 196 23495 264 23523
rect 298 23528 366 23529
rect 298 23495 332 23528
rect 196 23494 332 23495
rect 196 23489 366 23494
rect 230 23460 366 23489
rect 230 23455 264 23460
rect 196 23426 264 23455
rect 298 23459 366 23460
rect 298 23426 332 23459
rect 196 23425 332 23426
rect 196 23421 366 23425
rect 230 23391 366 23421
rect 230 23387 264 23391
rect 196 23357 264 23387
rect 298 23390 366 23391
rect 298 23357 332 23390
rect 196 23356 332 23357
rect 196 23353 366 23356
rect 230 23322 366 23353
rect 230 23319 264 23322
rect 196 23288 264 23319
rect 298 23321 366 23322
rect 298 23288 332 23321
rect 196 23287 332 23288
rect 196 23285 366 23287
rect 230 23253 366 23285
rect 230 23251 264 23253
rect 196 23219 264 23251
rect 298 23252 366 23253
rect 298 23219 332 23252
rect 196 23218 332 23219
rect 196 23217 366 23218
rect 230 23184 366 23217
rect 230 23183 264 23184
rect 196 23150 264 23183
rect 298 23183 366 23184
rect 298 23150 332 23183
rect 196 23149 332 23150
rect 366 23149 402 23183
rect 436 23149 472 23183
rect 506 23149 542 23183
rect 576 23149 612 23183
rect 646 23149 682 23183
rect 716 23149 752 23183
rect 786 23149 822 23183
rect 856 23149 891 23183
rect 925 23149 960 23183
rect 994 23149 1029 23183
rect 1063 23149 1098 23183
rect 1132 23149 1167 23183
rect 1201 23149 1236 23183
rect 1270 23149 1305 23183
rect 1339 23149 1374 23183
rect 1408 23149 1443 23183
rect 1477 23149 1512 23183
rect 1546 23149 1581 23183
rect 1615 23149 1650 23183
rect 1684 23149 1719 23183
rect 1753 23149 1788 23183
rect 1822 23149 1857 23183
rect 1891 23149 1926 23183
rect 1960 23149 1995 23183
rect 2029 23149 2064 23183
rect 2098 23149 2133 23183
rect 2167 23149 2202 23183
rect 2236 23149 2271 23183
rect 2305 23149 2340 23183
rect 2374 23149 2409 23183
rect 2443 23149 2478 23183
rect 2512 23149 2547 23183
rect 2581 23149 2616 23183
rect 2650 23149 2685 23183
rect 2719 23149 2754 23183
rect 2788 23149 2823 23183
rect 2857 23149 2892 23183
rect 2926 23149 2950 23183
rect 230 23115 2950 23149
rect 196 23081 264 23115
rect 298 23081 334 23115
rect 368 23081 404 23115
rect 438 23081 474 23115
rect 508 23081 544 23115
rect 578 23081 614 23115
rect 648 23081 684 23115
rect 718 23081 753 23115
rect 787 23081 822 23115
rect 856 23081 891 23115
rect 925 23081 960 23115
rect 994 23081 1029 23115
rect 1063 23081 1098 23115
rect 1132 23081 1167 23115
rect 1201 23081 1236 23115
rect 1270 23081 1305 23115
rect 1339 23081 1374 23115
rect 1408 23081 1443 23115
rect 1477 23081 1512 23115
rect 1546 23081 1581 23115
rect 1615 23081 1650 23115
rect 1684 23081 1719 23115
rect 1753 23081 1788 23115
rect 1822 23081 1857 23115
rect 1891 23081 1926 23115
rect 1960 23081 1995 23115
rect 2029 23081 2064 23115
rect 2098 23081 2133 23115
rect 2167 23081 2202 23115
rect 2236 23081 2271 23115
rect 2305 23081 2340 23115
rect 2374 23081 2409 23115
rect 2443 23081 2478 23115
rect 2512 23081 2547 23115
rect 2581 23081 2616 23115
rect 2650 23081 2685 23115
rect 2719 23081 2754 23115
rect 2788 23081 2823 23115
rect 2857 23081 2892 23115
rect 2926 23081 2950 23115
rect 196 23047 2950 23081
rect 196 23013 230 23047
rect 264 23013 299 23047
rect 333 23013 368 23047
rect 402 23013 437 23047
rect 471 23013 506 23047
rect 540 23013 575 23047
rect 609 23013 644 23047
rect 678 23013 713 23047
rect 747 23013 782 23047
rect 816 23013 851 23047
rect 885 23013 920 23047
rect 954 23013 988 23047
rect 1022 23013 1056 23047
rect 1090 23013 1124 23047
rect 1158 23013 1192 23047
rect 1226 23013 1260 23047
rect 1294 23013 1328 23047
rect 1362 23013 1396 23047
rect 1430 23013 1464 23047
rect 1498 23013 1532 23047
rect 1566 23013 1600 23047
rect 1634 23013 1668 23047
rect 1702 23013 1736 23047
rect 1770 23013 1804 23047
rect 1838 23013 1872 23047
rect 1906 23013 1940 23047
rect 1974 23013 2008 23047
rect 2042 23013 2076 23047
rect 2110 23013 2144 23047
rect 2178 23013 2212 23047
rect 2246 23013 2280 23047
rect 2314 23013 2348 23047
rect 2382 23013 2416 23047
rect 2450 23013 2484 23047
rect 2518 23013 2552 23047
rect 2586 23013 2620 23047
rect 2654 23013 2688 23047
rect 2722 23013 2756 23047
rect 2790 23013 2824 23047
rect 2858 23013 2892 23047
rect 2926 23013 2950 23047
rect 172 5219 206 5253
rect 240 5219 278 5253
rect 312 5219 350 5253
rect 384 5219 422 5253
rect 456 5219 494 5253
rect 528 5219 566 5253
rect 600 5219 638 5253
rect 672 5219 710 5253
rect 744 5219 782 5253
rect 816 5219 854 5253
rect 888 5219 925 5253
rect 959 5219 996 5253
rect 1030 5219 1067 5253
rect 1101 5219 1138 5253
rect 1172 5219 1209 5253
rect 1243 5219 1280 5253
rect 1314 5219 1422 5253
rect 172 5185 1388 5219
rect 172 5151 240 5185
rect 274 5151 312 5185
rect 346 5151 384 5185
rect 418 5151 456 5185
rect 490 5151 528 5185
rect 562 5151 600 5185
rect 634 5151 672 5185
rect 706 5151 744 5185
rect 778 5151 816 5185
rect 850 5151 888 5185
rect 922 5151 960 5185
rect 994 5151 1032 5185
rect 1066 5151 1104 5185
rect 1138 5151 1176 5185
rect 1210 5151 1248 5185
rect 1282 5151 1320 5185
rect 1354 5151 1422 5185
rect 172 5149 1422 5151
rect 206 5117 1388 5149
rect 206 5115 308 5117
rect 172 5113 308 5115
rect 172 5080 240 5113
rect 206 5079 240 5080
rect 274 5083 308 5113
rect 342 5083 381 5117
rect 415 5083 454 5117
rect 488 5083 527 5117
rect 561 5083 600 5117
rect 634 5083 673 5117
rect 707 5083 746 5117
rect 780 5083 819 5117
rect 853 5083 892 5117
rect 926 5083 964 5117
rect 998 5083 1036 5117
rect 1070 5083 1108 5117
rect 1142 5083 1180 5117
rect 1214 5083 1252 5117
rect 1286 5115 1388 5117
rect 1286 5112 1422 5115
rect 1286 5083 1320 5112
rect 274 5079 342 5083
rect 206 5046 342 5079
rect 172 5045 342 5046
rect 172 5041 308 5045
rect 172 5011 240 5041
rect 206 5007 240 5011
rect 274 5011 308 5041
rect 274 5007 342 5011
rect 206 4977 342 5007
rect 172 4973 342 4977
rect 172 4969 308 4973
rect 172 4942 240 4969
rect 206 4935 240 4942
rect 274 4939 308 4969
rect 1252 5078 1320 5083
rect 1354 5079 1422 5112
rect 1354 5078 1388 5079
rect 1252 5045 1388 5078
rect 1252 5044 1422 5045
rect 1286 5039 1422 5044
rect 1286 5010 1320 5039
rect 1252 5005 1320 5010
rect 1354 5009 1422 5039
rect 1354 5005 1388 5009
rect 1252 4975 1388 5005
rect 1252 4971 1422 4975
rect 274 4935 342 4939
rect 206 4908 342 4935
rect 172 4901 342 4908
rect 172 4897 308 4901
rect 172 4873 240 4897
rect 206 4863 240 4873
rect 274 4867 308 4897
rect 274 4863 342 4867
rect 206 4839 342 4863
rect 172 4829 342 4839
rect 172 4825 308 4829
rect 172 4804 240 4825
rect 206 4791 240 4804
rect 274 4795 308 4825
rect 274 4791 342 4795
rect 206 4770 342 4791
rect 172 4757 342 4770
rect 172 4753 308 4757
rect 172 4735 240 4753
rect 206 4719 240 4735
rect 274 4723 308 4753
rect 274 4719 342 4723
rect 206 4701 342 4719
rect 172 4685 342 4701
rect 1286 4967 1422 4971
rect 1286 4937 1320 4967
rect 1252 4933 1320 4937
rect 1354 4939 1422 4967
rect 1354 4933 1388 4939
rect 1252 4905 1388 4933
rect 1252 4898 1422 4905
rect 1286 4895 1422 4898
rect 1286 4864 1320 4895
rect 1252 4861 1320 4864
rect 1354 4869 1422 4895
rect 1354 4861 1388 4869
rect 1252 4835 1388 4861
rect 1252 4825 1422 4835
rect 1286 4823 1422 4825
rect 1286 4791 1320 4823
rect 1252 4789 1320 4791
rect 1354 4799 1422 4823
rect 1354 4789 1388 4799
rect 1252 4765 1388 4789
rect 1252 4752 1422 4765
rect 1286 4751 1422 4752
rect 1286 4718 1320 4751
rect 1252 4717 1320 4718
rect 1354 4730 1422 4751
rect 1354 4717 1388 4730
rect 1252 4696 1388 4717
rect 172 4681 308 4685
rect 172 4666 240 4681
rect 206 4647 240 4666
rect 274 4651 308 4681
rect 274 4647 342 4651
rect 206 4632 342 4647
rect 172 4612 342 4632
rect 172 4609 308 4612
rect 172 4597 240 4609
rect 206 4575 240 4597
rect 274 4578 308 4609
rect 274 4575 342 4578
rect 206 4563 342 4575
rect 172 4539 342 4563
rect 1252 4679 1422 4696
rect 1286 4645 1320 4679
rect 1354 4661 1422 4679
rect 1354 4645 1388 4661
rect 1252 4627 1388 4645
rect 1252 4607 1422 4627
rect 1286 4573 1320 4607
rect 1354 4592 1422 4607
rect 1354 4573 1388 4592
rect 1252 4558 1388 4573
rect 172 4537 308 4539
rect 172 4527 240 4537
rect 206 4503 240 4527
rect 274 4505 308 4537
rect 274 4503 342 4505
rect 206 4493 342 4503
rect 172 4466 342 4493
rect 172 4465 308 4466
rect 172 4457 240 4465
rect 206 4431 240 4457
rect 274 4432 308 4465
rect 274 4431 342 4432
rect 206 4423 342 4431
rect 172 4393 342 4423
rect 172 4387 240 4393
rect 206 4359 240 4387
rect 274 4359 308 4393
rect 206 4353 342 4359
rect 172 4320 342 4353
rect 172 4317 240 4320
rect 206 4286 240 4317
rect 274 4286 308 4320
rect 206 4283 342 4286
rect 172 4247 342 4283
rect 1252 4535 1422 4558
rect 1286 4501 1320 4535
rect 1354 4523 1422 4535
rect 1354 4501 1388 4523
rect 1252 4489 1388 4501
rect 1252 4463 1422 4489
rect 1286 4429 1320 4463
rect 1354 4454 1422 4463
rect 1354 4429 1388 4454
rect 1252 4420 1388 4429
rect 1252 4391 1422 4420
rect 1286 4357 1320 4391
rect 1354 4385 1422 4391
rect 1354 4357 1388 4385
rect 1252 4351 1388 4357
rect 1252 4319 1422 4351
rect 1286 4285 1320 4319
rect 1354 4316 1422 4319
rect 1354 4285 1388 4316
rect 1252 4282 1388 4285
rect 206 4213 240 4247
rect 274 4213 308 4247
rect 172 4189 342 4213
rect 1252 4247 1422 4282
rect 1286 4213 1320 4247
rect 1354 4213 1388 4247
rect 1252 4189 1422 4213
<< mvnsubdiff >>
rect -184 27717 -14 27741
rect -150 27683 -116 27717
rect -82 27683 -48 27717
rect -184 27648 -14 27683
rect -150 27614 -116 27648
rect -82 27614 -48 27648
rect -184 27579 -14 27614
rect -150 27545 -116 27579
rect -82 27545 -48 27579
rect -184 27510 -14 27545
rect -150 27476 -116 27510
rect -82 27476 -48 27510
rect -184 27441 -14 27476
rect -150 27407 -116 27441
rect -82 27407 -48 27441
rect -184 27372 -14 27407
rect -150 27338 -116 27372
rect -82 27338 -48 27372
rect -184 27303 -14 27338
rect -150 27269 -116 27303
rect -82 27269 -48 27303
rect -184 27234 -14 27269
rect -150 27200 -116 27234
rect -82 27200 -48 27234
rect -184 27165 -14 27200
rect -150 27131 -116 27165
rect -82 27131 -48 27165
rect -184 27096 -14 27131
rect -150 27062 -116 27096
rect -82 27062 -48 27096
rect -184 27027 -14 27062
rect -150 26993 -116 27027
rect -82 26993 -48 27027
rect -184 26958 -14 26993
rect -150 26924 -116 26958
rect -82 26924 -48 26958
rect -184 26889 -14 26924
rect -150 26855 -116 26889
rect -82 26855 -48 26889
rect -184 26820 -14 26855
rect -150 26786 -116 26820
rect -82 26786 -48 26820
rect -184 26751 -14 26786
rect -150 26717 -116 26751
rect -82 26717 -48 26751
rect -184 26682 -14 26717
rect -150 26648 -116 26682
rect -82 26648 -48 26682
rect -184 26613 -14 26648
rect -150 26579 -116 26613
rect -82 26579 -48 26613
rect -184 26544 -14 26579
rect -150 26510 -116 26544
rect -82 26510 -48 26544
rect -184 26475 -14 26510
rect -150 26441 -116 26475
rect -82 26441 -48 26475
rect -184 26406 -14 26441
rect -150 26372 -116 26406
rect -82 26372 -48 26406
rect -184 26337 -14 26372
rect -150 26303 -116 26337
rect -82 26303 -48 26337
rect -184 26268 -14 26303
rect -150 26234 -116 26268
rect -82 26234 -48 26268
rect -184 26199 -14 26234
rect -150 26165 -116 26199
rect -82 26165 -48 26199
rect -184 26130 -14 26165
rect -150 26096 -116 26130
rect -82 26096 -48 26130
rect -184 26061 -14 26096
rect -150 26027 -116 26061
rect -82 26027 -48 26061
rect -184 25992 -14 26027
rect -150 25958 -116 25992
rect -82 25958 -48 25992
rect -184 25923 -14 25958
rect -150 25889 -116 25923
rect -82 25889 -48 25923
rect -184 25854 -14 25889
rect -150 25820 -116 25854
rect -82 25820 -48 25854
rect -184 25785 -14 25820
rect -150 25751 -116 25785
rect -82 25751 -48 25785
rect -184 25717 -14 25751
rect -150 25716 -14 25717
rect -150 25683 -116 25716
rect -184 25682 -116 25683
rect -82 25682 -48 25716
rect -184 25649 -14 25682
rect -150 25647 -14 25649
rect -150 25615 -116 25647
rect -184 25613 -116 25615
rect -82 25613 -48 25647
rect -184 25581 -14 25613
rect -150 25578 -14 25581
rect -150 25547 -116 25578
rect -184 25544 -116 25547
rect -82 25544 -48 25578
rect -184 25513 -14 25544
rect -150 25509 -14 25513
rect -150 25479 -116 25509
rect -184 25475 -116 25479
rect -82 25475 -48 25509
rect -184 25445 -14 25475
rect -150 25440 -14 25445
rect -150 25411 -116 25440
rect -184 25406 -116 25411
rect -82 25406 -48 25440
rect -184 25377 -14 25406
rect -150 25371 -14 25377
rect -150 25343 -116 25371
rect -184 25337 -116 25343
rect -82 25337 -48 25371
rect -184 25309 -14 25337
rect -150 25302 -14 25309
rect -150 25275 -116 25302
rect -184 25268 -116 25275
rect -82 25268 -48 25302
rect -184 25241 -14 25268
rect -150 25233 -14 25241
rect -150 25207 -116 25233
rect -184 25199 -116 25207
rect -82 25199 -48 25233
rect -184 25173 -14 25199
rect -150 25164 -14 25173
rect -150 25139 -116 25164
rect -184 25130 -116 25139
rect -82 25130 -48 25164
rect -184 25105 -14 25130
rect -150 25095 -14 25105
rect -150 25071 -116 25095
rect -184 25061 -116 25071
rect -82 25061 -48 25095
rect -184 25037 -14 25061
rect -150 25026 -14 25037
rect -150 25003 -116 25026
rect -184 24992 -116 25003
rect -82 24992 -48 25026
rect -184 24969 -14 24992
rect -150 24957 -14 24969
rect -150 24935 -116 24957
rect -184 24923 -116 24935
rect -82 24923 -48 24957
rect -184 24901 -14 24923
rect -150 24888 -14 24901
rect -150 24867 -116 24888
rect -184 24854 -116 24867
rect -82 24854 -48 24888
rect -184 24833 -14 24854
rect -150 24819 -14 24833
rect -150 24799 -116 24819
rect -184 24785 -116 24799
rect -82 24785 -48 24819
rect -184 24765 -14 24785
rect -150 24750 -14 24765
rect -150 24731 -116 24750
rect -184 24716 -116 24731
rect -82 24716 -48 24750
rect -184 24697 -14 24716
rect -150 24681 -14 24697
rect -150 24663 -116 24681
rect -184 24647 -116 24663
rect -82 24647 -48 24681
rect -184 24629 -14 24647
rect -150 24612 -14 24629
rect -150 24595 -116 24612
rect -184 24578 -116 24595
rect -82 24578 -48 24612
rect -184 24561 -14 24578
rect -150 24543 -14 24561
rect -150 24527 -116 24543
rect -184 24509 -116 24527
rect -82 24509 -48 24543
rect -184 24493 -14 24509
rect -150 24474 -14 24493
rect -150 24459 -116 24474
rect -184 24440 -116 24459
rect -82 24440 -48 24474
rect -184 24425 -14 24440
rect -150 24405 -14 24425
rect -150 24391 -116 24405
rect -184 24371 -116 24391
rect -82 24371 -48 24405
rect -184 24357 -14 24371
rect -150 24336 -14 24357
rect -150 24323 -116 24336
rect -184 24302 -116 24323
rect -82 24302 -48 24336
rect -184 24289 -14 24302
rect -150 24267 -14 24289
rect -150 24255 -116 24267
rect -184 24233 -116 24255
rect -82 24233 -48 24267
rect -184 24221 -14 24233
rect -150 24198 -14 24221
rect -150 24187 -116 24198
rect -184 24164 -116 24187
rect -82 24164 -48 24198
rect -184 24153 -14 24164
rect -150 24129 -14 24153
rect -150 24119 -116 24129
rect -184 24095 -116 24119
rect -82 24095 -48 24129
rect -184 24085 -14 24095
rect -150 24060 -14 24085
rect -150 24051 -116 24060
rect -184 24026 -116 24051
rect -82 24026 -48 24060
rect -184 24017 -14 24026
rect -150 23991 -14 24017
rect -150 23983 -116 23991
rect -184 23957 -116 23983
rect -82 23957 -48 23991
rect -184 23949 -14 23957
rect -150 23922 -14 23949
rect -150 23915 -116 23922
rect -184 23888 -116 23915
rect -82 23888 -48 23922
rect -184 23881 -14 23888
rect -150 23853 -14 23881
rect -150 23847 -116 23853
rect -184 23819 -116 23847
rect -82 23819 -48 23853
rect -184 23813 -14 23819
rect -150 23784 -14 23813
rect -150 23779 -116 23784
rect -184 23750 -116 23779
rect -82 23750 -48 23784
rect -184 23745 -14 23750
rect -150 23715 -14 23745
rect -150 23711 -116 23715
rect -184 23681 -116 23711
rect -82 23681 -48 23715
rect -184 23677 -14 23681
rect -150 23646 -14 23677
rect -150 23643 -116 23646
rect -184 23612 -116 23643
rect -82 23612 -48 23646
rect -184 23609 -14 23612
rect -150 23577 -14 23609
rect -150 23575 -116 23577
rect -184 23543 -116 23575
rect -82 23543 -48 23577
rect -184 23541 -14 23543
rect -150 23508 -14 23541
rect -150 23507 -116 23508
rect -184 23474 -116 23507
rect -82 23474 -48 23508
rect -184 23473 -14 23474
rect -150 23439 -14 23473
rect 518 24942 552 25050
rect 586 25016 623 25050
rect 657 25016 694 25050
rect 728 25016 764 25050
rect 798 25016 834 25050
rect 868 25016 892 25050
rect 518 24871 552 24908
rect 518 24800 552 24837
rect 518 24729 552 24766
rect 518 24658 552 24695
rect 518 24587 552 24624
rect 518 24516 552 24553
rect 518 24445 552 24482
rect 518 24374 552 24411
rect 518 24303 552 24340
rect 518 24221 552 24269
rect 1758 24221 1792 24245
rect 518 24148 552 24187
rect 518 24075 552 24114
rect 518 24001 552 24041
rect 518 23927 552 23967
rect 1758 24147 1792 24187
rect 1758 24073 1792 24113
rect 1758 23999 1792 24039
rect 1758 23925 1792 23965
rect 518 23853 552 23893
rect 518 23779 552 23819
rect 1758 23852 1792 23891
rect 518 23705 552 23745
rect 518 23631 552 23671
rect 518 23557 552 23597
rect 518 23483 552 23523
rect 1758 23779 1792 23818
rect 1758 23706 1792 23745
rect 1758 23633 1792 23672
rect 1758 23560 1792 23599
rect 518 23409 552 23449
rect 1758 23487 1792 23526
rect 518 23341 620 23375
rect 654 23341 689 23375
rect 723 23341 758 23375
rect 792 23341 827 23375
rect 861 23341 896 23375
rect 930 23341 965 23375
rect 999 23341 1034 23375
rect 1068 23341 1103 23375
rect 1137 23341 1172 23375
rect 1206 23341 1241 23375
rect 1275 23341 1310 23375
rect 1344 23341 1379 23375
rect 1413 23341 1448 23375
rect 1482 23341 1517 23375
rect 1551 23341 1586 23375
rect 1620 23341 1655 23375
rect 1689 23341 1724 23375
rect 1758 23341 1792 23453
rect -14 22725 21 22759
rect 55 22725 90 22759
rect 124 22725 159 22759
rect 193 22725 228 22759
rect 262 22725 297 22759
rect 331 22725 366 22759
rect 400 22725 435 22759
rect 469 22725 504 22759
rect 538 22725 573 22759
rect 607 22725 642 22759
rect 676 22725 711 22759
rect 745 22725 780 22759
rect -82 22691 780 22725
rect -184 22657 -116 22691
rect -82 22657 -47 22691
rect -13 22657 22 22691
rect 56 22657 91 22691
rect 125 22657 160 22691
rect 194 22657 229 22691
rect 263 22657 298 22691
rect 332 22657 367 22691
rect 401 22657 436 22691
rect 470 22657 505 22691
rect 539 22657 574 22691
rect 608 22657 643 22691
rect 677 22657 712 22691
rect 746 22657 780 22691
rect 2174 22657 2231 22759
rect -184 22623 2231 22657
rect -184 22589 -150 22623
rect -116 22589 -80 22623
rect -46 22589 -10 22623
rect 24 22589 60 22623
rect 94 22589 130 22623
rect 164 22589 200 22623
rect 234 22589 270 22623
rect 304 22589 340 22623
rect 374 22589 410 22623
rect 444 22589 480 22623
rect 514 22589 550 22623
rect 584 22589 620 22623
rect 654 22589 690 22623
rect 724 22589 760 22623
rect 794 22589 829 22623
rect 863 22589 898 22623
rect 932 22589 967 22623
rect 1001 22589 1036 22623
rect 1070 22589 1105 22623
rect 1139 22589 1174 22623
rect 1208 22589 1243 22623
rect 1277 22589 1312 22623
rect 1346 22589 1381 22623
rect 1415 22589 1450 22623
rect 1484 22589 1519 22623
rect 1553 22589 1588 22623
rect 1622 22589 1657 22623
rect 1691 22589 1726 22623
rect 1760 22589 1795 22623
rect 1829 22589 1864 22623
rect 1898 22589 1933 22623
rect 1967 22589 2002 22623
rect 2036 22589 2071 22623
rect 2105 22589 2140 22623
rect 2174 22589 2231 22623
<< mvpsubdiffcont >>
rect 230 27707 264 27741
rect 299 27707 333 27741
rect 368 27707 402 27741
rect 437 27707 471 27741
rect 506 27707 540 27741
rect 575 27707 609 27741
rect 644 27707 678 27741
rect 713 27707 747 27741
rect 782 27707 816 27741
rect 851 27707 885 27741
rect 920 27707 954 27741
rect 988 27707 1022 27741
rect 1056 27707 1090 27741
rect 1124 27707 1158 27741
rect 1192 27707 1226 27741
rect 1260 27707 1294 27741
rect 1328 27707 1362 27741
rect 1396 27707 1430 27741
rect 1464 27707 1498 27741
rect 1532 27707 1566 27741
rect 1600 27707 1634 27741
rect 1668 27707 1702 27741
rect 1736 27707 1770 27741
rect 1804 27707 1838 27741
rect 1872 27707 1906 27741
rect 1940 27707 1974 27741
rect 2008 27707 2042 27741
rect 2076 27707 2110 27741
rect 2144 27707 2178 27741
rect 2212 27707 2246 27741
rect 2280 27707 2314 27741
rect 2348 27707 2382 27741
rect 2416 27707 2450 27741
rect 2484 27707 2518 27741
rect 2552 27707 2586 27741
rect 2620 27707 2654 27741
rect 2688 27707 2722 27741
rect 2756 27707 2790 27741
rect 2824 27707 2858 27741
rect 2892 27707 2926 27741
rect 264 27639 298 27673
rect 334 27639 368 27673
rect 404 27639 438 27673
rect 474 27639 508 27673
rect 544 27639 578 27673
rect 614 27639 648 27673
rect 684 27639 718 27673
rect 753 27639 787 27673
rect 822 27639 856 27673
rect 891 27639 925 27673
rect 960 27639 994 27673
rect 1029 27639 1063 27673
rect 1098 27639 1132 27673
rect 1167 27639 1201 27673
rect 1236 27639 1270 27673
rect 1305 27639 1339 27673
rect 1374 27639 1408 27673
rect 1443 27639 1477 27673
rect 1512 27639 1546 27673
rect 1581 27639 1615 27673
rect 1650 27639 1684 27673
rect 1719 27639 1753 27673
rect 1788 27639 1822 27673
rect 1857 27639 1891 27673
rect 1926 27639 1960 27673
rect 1995 27639 2029 27673
rect 2064 27639 2098 27673
rect 2133 27639 2167 27673
rect 2202 27639 2236 27673
rect 2271 27639 2305 27673
rect 2340 27639 2374 27673
rect 2409 27639 2443 27673
rect 2478 27639 2512 27673
rect 2547 27639 2581 27673
rect 2616 27639 2650 27673
rect 2685 27639 2719 27673
rect 2754 27639 2788 27673
rect 2823 27639 2857 27673
rect 2892 27639 2926 27673
rect 196 27597 230 27631
rect 196 27524 230 27558
rect 264 27552 298 27586
rect 332 27571 366 27605
rect 402 27571 436 27605
rect 472 27571 506 27605
rect 542 27571 576 27605
rect 612 27571 646 27605
rect 682 27571 716 27605
rect 752 27571 786 27605
rect 822 27571 856 27605
rect 891 27571 925 27605
rect 960 27571 994 27605
rect 1029 27571 1063 27605
rect 1098 27571 1132 27605
rect 1167 27571 1201 27605
rect 1236 27571 1270 27605
rect 1305 27571 1339 27605
rect 1374 27571 1408 27605
rect 1443 27571 1477 27605
rect 1512 27571 1546 27605
rect 1581 27571 1615 27605
rect 1650 27571 1684 27605
rect 1719 27571 1753 27605
rect 1788 27571 1822 27605
rect 1857 27571 1891 27605
rect 1926 27571 1960 27605
rect 1995 27571 2029 27605
rect 2064 27571 2098 27605
rect 2133 27571 2167 27605
rect 2202 27571 2236 27605
rect 2271 27571 2305 27605
rect 2340 27571 2374 27605
rect 2409 27571 2443 27605
rect 2478 27571 2512 27605
rect 2547 27571 2581 27605
rect 2616 27571 2650 27605
rect 2685 27571 2719 27605
rect 2754 27571 2788 27605
rect 2823 27571 2857 27605
rect 2892 27571 2926 27605
rect 196 27451 230 27485
rect 264 27465 298 27499
rect 332 27475 366 27509
rect 196 27378 230 27412
rect 264 27378 298 27412
rect 332 27378 366 27412
rect 196 27296 230 27330
rect 264 27296 298 27330
rect 332 27296 366 27330
rect 196 27227 230 27261
rect 264 27226 298 27260
rect 332 27226 366 27260
rect 196 27158 230 27192
rect 264 27156 298 27190
rect 332 27156 366 27190
rect 196 27089 230 27123
rect 264 27086 298 27120
rect 332 27086 366 27120
rect 196 27020 230 27054
rect 264 27016 298 27050
rect 332 27016 366 27050
rect 196 26951 230 26985
rect 264 26946 298 26980
rect 332 26946 366 26980
rect 196 26882 230 26916
rect 264 26876 298 26910
rect 332 26876 366 26910
rect 196 26813 230 26847
rect 264 26807 298 26841
rect 332 26806 366 26840
rect 196 26744 230 26778
rect 264 26738 298 26772
rect 332 26737 366 26771
rect 196 26675 230 26709
rect 264 26669 298 26703
rect 332 26668 366 26702
rect 196 26606 230 26640
rect 264 26600 298 26634
rect 332 26599 366 26633
rect 196 26537 230 26571
rect 264 26531 298 26565
rect 332 26530 366 26564
rect 196 26468 230 26502
rect 264 26462 298 26496
rect 332 26461 366 26495
rect 196 26399 230 26433
rect 264 26393 298 26427
rect 332 26392 366 26426
rect 196 26330 230 26364
rect 264 26324 298 26358
rect 332 26323 366 26357
rect 196 26261 230 26295
rect 264 26255 298 26289
rect 332 26254 366 26288
rect 196 26192 230 26226
rect 264 26186 298 26220
rect 332 26185 366 26219
rect 196 26123 230 26157
rect 264 26117 298 26151
rect 332 26116 366 26150
rect 196 26054 230 26088
rect 264 26048 298 26082
rect 332 26047 366 26081
rect 196 25985 230 26019
rect 264 25979 298 26013
rect 332 25978 366 26012
rect 196 25916 230 25950
rect 264 25910 298 25944
rect 332 25909 366 25943
rect 196 25847 230 25881
rect 264 25841 298 25875
rect 332 25840 366 25874
rect 196 25778 230 25812
rect 264 25772 298 25806
rect 332 25771 366 25805
rect 196 25709 230 25743
rect 264 25703 298 25737
rect 332 25702 366 25736
rect 196 25640 230 25674
rect 264 25634 298 25668
rect 332 25633 366 25667
rect 196 25571 230 25605
rect 264 25565 298 25599
rect 332 25564 366 25598
rect 196 25502 230 25536
rect 264 25496 298 25530
rect 332 25495 366 25529
rect 196 25433 230 25467
rect 264 25427 298 25461
rect 332 25426 366 25460
rect 196 25364 230 25398
rect 264 25358 298 25392
rect 332 25357 366 25391
rect 196 25295 230 25329
rect 264 25289 298 25323
rect 332 25288 366 25322
rect 196 25226 230 25260
rect 264 25220 298 25254
rect 332 25219 366 25253
rect 196 25157 230 25191
rect 264 25151 298 25185
rect 332 25150 366 25184
rect 196 25088 230 25122
rect 264 25082 298 25116
rect 332 25081 366 25115
rect 196 25019 230 25053
rect 264 25013 298 25047
rect 332 25012 366 25046
rect 196 24951 230 24985
rect 264 24944 298 24978
rect 332 24943 366 24977
rect 196 24883 230 24917
rect 264 24875 298 24909
rect 332 24874 366 24908
rect 196 24815 230 24849
rect 264 24806 298 24840
rect 332 24805 366 24839
rect 196 24747 230 24781
rect 264 24737 298 24771
rect 332 24736 366 24770
rect 196 24679 230 24713
rect 264 24668 298 24702
rect 332 24667 366 24701
rect 196 24611 230 24645
rect 264 24599 298 24633
rect 332 24598 366 24632
rect 196 24543 230 24577
rect 264 24530 298 24564
rect 332 24529 366 24563
rect 196 24475 230 24509
rect 264 24461 298 24495
rect 332 24460 366 24494
rect 196 24407 230 24441
rect 264 24392 298 24426
rect 332 24391 366 24425
rect 196 24339 230 24373
rect 264 24323 298 24357
rect 332 24322 366 24356
rect 196 24271 230 24305
rect 264 24254 298 24288
rect 332 24253 366 24287
rect 196 24203 230 24237
rect 264 24185 298 24219
rect 332 24184 366 24218
rect 196 24135 230 24169
rect 264 24116 298 24150
rect 332 24115 366 24149
rect 196 24067 230 24101
rect 264 24047 298 24081
rect 332 24046 366 24080
rect 196 23999 230 24033
rect 264 23978 298 24012
rect 332 23977 366 24011
rect 196 23931 230 23965
rect 264 23909 298 23943
rect 332 23908 366 23942
rect 196 23863 230 23897
rect 264 23840 298 23874
rect 332 23839 366 23873
rect 196 23795 230 23829
rect 264 23771 298 23805
rect 332 23770 366 23804
rect 196 23727 230 23761
rect 264 23702 298 23736
rect 332 23701 366 23735
rect 196 23659 230 23693
rect 264 23633 298 23667
rect 332 23632 366 23666
rect 196 23591 230 23625
rect 264 23564 298 23598
rect 332 23563 366 23597
rect 196 23523 230 23557
rect 264 23495 298 23529
rect 332 23494 366 23528
rect 196 23455 230 23489
rect 264 23426 298 23460
rect 332 23425 366 23459
rect 196 23387 230 23421
rect 264 23357 298 23391
rect 332 23356 366 23390
rect 196 23319 230 23353
rect 264 23288 298 23322
rect 332 23287 366 23321
rect 196 23251 230 23285
rect 264 23219 298 23253
rect 332 23218 366 23252
rect 196 23183 230 23217
rect 264 23150 298 23184
rect 332 23149 366 23183
rect 402 23149 436 23183
rect 472 23149 506 23183
rect 542 23149 576 23183
rect 612 23149 646 23183
rect 682 23149 716 23183
rect 752 23149 786 23183
rect 822 23149 856 23183
rect 891 23149 925 23183
rect 960 23149 994 23183
rect 1029 23149 1063 23183
rect 1098 23149 1132 23183
rect 1167 23149 1201 23183
rect 1236 23149 1270 23183
rect 1305 23149 1339 23183
rect 1374 23149 1408 23183
rect 1443 23149 1477 23183
rect 1512 23149 1546 23183
rect 1581 23149 1615 23183
rect 1650 23149 1684 23183
rect 1719 23149 1753 23183
rect 1788 23149 1822 23183
rect 1857 23149 1891 23183
rect 1926 23149 1960 23183
rect 1995 23149 2029 23183
rect 2064 23149 2098 23183
rect 2133 23149 2167 23183
rect 2202 23149 2236 23183
rect 2271 23149 2305 23183
rect 2340 23149 2374 23183
rect 2409 23149 2443 23183
rect 2478 23149 2512 23183
rect 2547 23149 2581 23183
rect 2616 23149 2650 23183
rect 2685 23149 2719 23183
rect 2754 23149 2788 23183
rect 2823 23149 2857 23183
rect 2892 23149 2926 23183
rect 196 23115 230 23149
rect 264 23081 298 23115
rect 334 23081 368 23115
rect 404 23081 438 23115
rect 474 23081 508 23115
rect 544 23081 578 23115
rect 614 23081 648 23115
rect 684 23081 718 23115
rect 753 23081 787 23115
rect 822 23081 856 23115
rect 891 23081 925 23115
rect 960 23081 994 23115
rect 1029 23081 1063 23115
rect 1098 23081 1132 23115
rect 1167 23081 1201 23115
rect 1236 23081 1270 23115
rect 1305 23081 1339 23115
rect 1374 23081 1408 23115
rect 1443 23081 1477 23115
rect 1512 23081 1546 23115
rect 1581 23081 1615 23115
rect 1650 23081 1684 23115
rect 1719 23081 1753 23115
rect 1788 23081 1822 23115
rect 1857 23081 1891 23115
rect 1926 23081 1960 23115
rect 1995 23081 2029 23115
rect 2064 23081 2098 23115
rect 2133 23081 2167 23115
rect 2202 23081 2236 23115
rect 2271 23081 2305 23115
rect 2340 23081 2374 23115
rect 2409 23081 2443 23115
rect 2478 23081 2512 23115
rect 2547 23081 2581 23115
rect 2616 23081 2650 23115
rect 2685 23081 2719 23115
rect 2754 23081 2788 23115
rect 2823 23081 2857 23115
rect 2892 23081 2926 23115
rect 230 23013 264 23047
rect 299 23013 333 23047
rect 368 23013 402 23047
rect 437 23013 471 23047
rect 506 23013 540 23047
rect 575 23013 609 23047
rect 644 23013 678 23047
rect 713 23013 747 23047
rect 782 23013 816 23047
rect 851 23013 885 23047
rect 920 23013 954 23047
rect 988 23013 1022 23047
rect 1056 23013 1090 23047
rect 1124 23013 1158 23047
rect 1192 23013 1226 23047
rect 1260 23013 1294 23047
rect 1328 23013 1362 23047
rect 1396 23013 1430 23047
rect 1464 23013 1498 23047
rect 1532 23013 1566 23047
rect 1600 23013 1634 23047
rect 1668 23013 1702 23047
rect 1736 23013 1770 23047
rect 1804 23013 1838 23047
rect 1872 23013 1906 23047
rect 1940 23013 1974 23047
rect 2008 23013 2042 23047
rect 2076 23013 2110 23047
rect 2144 23013 2178 23047
rect 2212 23013 2246 23047
rect 2280 23013 2314 23047
rect 2348 23013 2382 23047
rect 2416 23013 2450 23047
rect 2484 23013 2518 23047
rect 2552 23013 2586 23047
rect 2620 23013 2654 23047
rect 2688 23013 2722 23047
rect 2756 23013 2790 23047
rect 2824 23013 2858 23047
rect 2892 23013 2926 23047
rect 206 5219 240 5253
rect 278 5219 312 5253
rect 350 5219 384 5253
rect 422 5219 456 5253
rect 494 5219 528 5253
rect 566 5219 600 5253
rect 638 5219 672 5253
rect 710 5219 744 5253
rect 782 5219 816 5253
rect 854 5219 888 5253
rect 925 5219 959 5253
rect 996 5219 1030 5253
rect 1067 5219 1101 5253
rect 1138 5219 1172 5253
rect 1209 5219 1243 5253
rect 1280 5219 1314 5253
rect 1388 5185 1422 5219
rect 240 5151 274 5185
rect 312 5151 346 5185
rect 384 5151 418 5185
rect 456 5151 490 5185
rect 528 5151 562 5185
rect 600 5151 634 5185
rect 672 5151 706 5185
rect 744 5151 778 5185
rect 816 5151 850 5185
rect 888 5151 922 5185
rect 960 5151 994 5185
rect 1032 5151 1066 5185
rect 1104 5151 1138 5185
rect 1176 5151 1210 5185
rect 1248 5151 1282 5185
rect 1320 5151 1354 5185
rect 172 5115 206 5149
rect 172 5046 206 5080
rect 240 5079 274 5113
rect 308 5083 342 5117
rect 381 5083 415 5117
rect 454 5083 488 5117
rect 527 5083 561 5117
rect 600 5083 634 5117
rect 673 5083 707 5117
rect 746 5083 780 5117
rect 819 5083 853 5117
rect 892 5083 926 5117
rect 964 5083 998 5117
rect 1036 5083 1070 5117
rect 1108 5083 1142 5117
rect 1180 5083 1214 5117
rect 1252 5083 1286 5117
rect 1388 5115 1422 5149
rect 172 4977 206 5011
rect 240 5007 274 5041
rect 308 5011 342 5045
rect 172 4908 206 4942
rect 240 4935 274 4969
rect 308 4939 342 4973
rect 1320 5078 1354 5112
rect 1388 5045 1422 5079
rect 1252 5010 1286 5044
rect 1320 5005 1354 5039
rect 1388 4975 1422 5009
rect 172 4839 206 4873
rect 240 4863 274 4897
rect 308 4867 342 4901
rect 172 4770 206 4804
rect 240 4791 274 4825
rect 308 4795 342 4829
rect 172 4701 206 4735
rect 240 4719 274 4753
rect 308 4723 342 4757
rect 1252 4937 1286 4971
rect 1320 4933 1354 4967
rect 1388 4905 1422 4939
rect 1252 4864 1286 4898
rect 1320 4861 1354 4895
rect 1388 4835 1422 4869
rect 1252 4791 1286 4825
rect 1320 4789 1354 4823
rect 1388 4765 1422 4799
rect 1252 4718 1286 4752
rect 1320 4717 1354 4751
rect 1388 4696 1422 4730
rect 172 4632 206 4666
rect 240 4647 274 4681
rect 308 4651 342 4685
rect 172 4563 206 4597
rect 240 4575 274 4609
rect 308 4578 342 4612
rect 1252 4645 1286 4679
rect 1320 4645 1354 4679
rect 1388 4627 1422 4661
rect 1252 4573 1286 4607
rect 1320 4573 1354 4607
rect 1388 4558 1422 4592
rect 172 4493 206 4527
rect 240 4503 274 4537
rect 308 4505 342 4539
rect 172 4423 206 4457
rect 240 4431 274 4465
rect 308 4432 342 4466
rect 172 4353 206 4387
rect 240 4359 274 4393
rect 308 4359 342 4393
rect 172 4283 206 4317
rect 240 4286 274 4320
rect 308 4286 342 4320
rect 1252 4501 1286 4535
rect 1320 4501 1354 4535
rect 1388 4489 1422 4523
rect 1252 4429 1286 4463
rect 1320 4429 1354 4463
rect 1388 4420 1422 4454
rect 1252 4357 1286 4391
rect 1320 4357 1354 4391
rect 1388 4351 1422 4385
rect 1252 4285 1286 4319
rect 1320 4285 1354 4319
rect 1388 4282 1422 4316
rect 172 4213 206 4247
rect 240 4213 274 4247
rect 308 4213 342 4247
rect 1252 4213 1286 4247
rect 1320 4213 1354 4247
rect 1388 4213 1422 4247
<< mvnsubdiffcont >>
rect -184 27683 -150 27717
rect -116 27683 -82 27717
rect -48 27683 -14 27717
rect -184 27614 -150 27648
rect -116 27614 -82 27648
rect -48 27614 -14 27648
rect -184 27545 -150 27579
rect -116 27545 -82 27579
rect -48 27545 -14 27579
rect -184 27476 -150 27510
rect -116 27476 -82 27510
rect -48 27476 -14 27510
rect -184 27407 -150 27441
rect -116 27407 -82 27441
rect -48 27407 -14 27441
rect -184 27338 -150 27372
rect -116 27338 -82 27372
rect -48 27338 -14 27372
rect -184 27269 -150 27303
rect -116 27269 -82 27303
rect -48 27269 -14 27303
rect -184 27200 -150 27234
rect -116 27200 -82 27234
rect -48 27200 -14 27234
rect -184 27131 -150 27165
rect -116 27131 -82 27165
rect -48 27131 -14 27165
rect -184 27062 -150 27096
rect -116 27062 -82 27096
rect -48 27062 -14 27096
rect -184 26993 -150 27027
rect -116 26993 -82 27027
rect -48 26993 -14 27027
rect -184 26924 -150 26958
rect -116 26924 -82 26958
rect -48 26924 -14 26958
rect -184 26855 -150 26889
rect -116 26855 -82 26889
rect -48 26855 -14 26889
rect -184 26786 -150 26820
rect -116 26786 -82 26820
rect -48 26786 -14 26820
rect -184 26717 -150 26751
rect -116 26717 -82 26751
rect -48 26717 -14 26751
rect -184 26648 -150 26682
rect -116 26648 -82 26682
rect -48 26648 -14 26682
rect -184 26579 -150 26613
rect -116 26579 -82 26613
rect -48 26579 -14 26613
rect -184 26510 -150 26544
rect -116 26510 -82 26544
rect -48 26510 -14 26544
rect -184 26441 -150 26475
rect -116 26441 -82 26475
rect -48 26441 -14 26475
rect -184 26372 -150 26406
rect -116 26372 -82 26406
rect -48 26372 -14 26406
rect -184 26303 -150 26337
rect -116 26303 -82 26337
rect -48 26303 -14 26337
rect -184 26234 -150 26268
rect -116 26234 -82 26268
rect -48 26234 -14 26268
rect -184 26165 -150 26199
rect -116 26165 -82 26199
rect -48 26165 -14 26199
rect -184 26096 -150 26130
rect -116 26096 -82 26130
rect -48 26096 -14 26130
rect -184 26027 -150 26061
rect -116 26027 -82 26061
rect -48 26027 -14 26061
rect -184 25958 -150 25992
rect -116 25958 -82 25992
rect -48 25958 -14 25992
rect -184 25889 -150 25923
rect -116 25889 -82 25923
rect -48 25889 -14 25923
rect -184 25820 -150 25854
rect -116 25820 -82 25854
rect -48 25820 -14 25854
rect -184 25751 -150 25785
rect -116 25751 -82 25785
rect -48 25751 -14 25785
rect -184 25683 -150 25717
rect -116 25682 -82 25716
rect -48 25682 -14 25716
rect -184 25615 -150 25649
rect -116 25613 -82 25647
rect -48 25613 -14 25647
rect -184 25547 -150 25581
rect -116 25544 -82 25578
rect -48 25544 -14 25578
rect -184 25479 -150 25513
rect -116 25475 -82 25509
rect -48 25475 -14 25509
rect -184 25411 -150 25445
rect -116 25406 -82 25440
rect -48 25406 -14 25440
rect -184 25343 -150 25377
rect -116 25337 -82 25371
rect -48 25337 -14 25371
rect -184 25275 -150 25309
rect -116 25268 -82 25302
rect -48 25268 -14 25302
rect -184 25207 -150 25241
rect -116 25199 -82 25233
rect -48 25199 -14 25233
rect -184 25139 -150 25173
rect -116 25130 -82 25164
rect -48 25130 -14 25164
rect -184 25071 -150 25105
rect -116 25061 -82 25095
rect -48 25061 -14 25095
rect -184 25003 -150 25037
rect -116 24992 -82 25026
rect -48 24992 -14 25026
rect -184 24935 -150 24969
rect -116 24923 -82 24957
rect -48 24923 -14 24957
rect -184 24867 -150 24901
rect -116 24854 -82 24888
rect -48 24854 -14 24888
rect -184 24799 -150 24833
rect -116 24785 -82 24819
rect -48 24785 -14 24819
rect -184 24731 -150 24765
rect -116 24716 -82 24750
rect -48 24716 -14 24750
rect -184 24663 -150 24697
rect -116 24647 -82 24681
rect -48 24647 -14 24681
rect -184 24595 -150 24629
rect -116 24578 -82 24612
rect -48 24578 -14 24612
rect -184 24527 -150 24561
rect -116 24509 -82 24543
rect -48 24509 -14 24543
rect -184 24459 -150 24493
rect -116 24440 -82 24474
rect -48 24440 -14 24474
rect -184 24391 -150 24425
rect -116 24371 -82 24405
rect -48 24371 -14 24405
rect -184 24323 -150 24357
rect -116 24302 -82 24336
rect -48 24302 -14 24336
rect -184 24255 -150 24289
rect -116 24233 -82 24267
rect -48 24233 -14 24267
rect -184 24187 -150 24221
rect -116 24164 -82 24198
rect -48 24164 -14 24198
rect -184 24119 -150 24153
rect -116 24095 -82 24129
rect -48 24095 -14 24129
rect -184 24051 -150 24085
rect -116 24026 -82 24060
rect -48 24026 -14 24060
rect -184 23983 -150 24017
rect -116 23957 -82 23991
rect -48 23957 -14 23991
rect -184 23915 -150 23949
rect -116 23888 -82 23922
rect -48 23888 -14 23922
rect -184 23847 -150 23881
rect -116 23819 -82 23853
rect -48 23819 -14 23853
rect -184 23779 -150 23813
rect -116 23750 -82 23784
rect -48 23750 -14 23784
rect -184 23711 -150 23745
rect -116 23681 -82 23715
rect -48 23681 -14 23715
rect -184 23643 -150 23677
rect -116 23612 -82 23646
rect -48 23612 -14 23646
rect -184 23575 -150 23609
rect -116 23543 -82 23577
rect -48 23543 -14 23577
rect -184 23507 -150 23541
rect -116 23474 -82 23508
rect -48 23474 -14 23508
rect -184 23439 -150 23473
rect -184 22725 -14 23439
rect 552 25016 586 25050
rect 623 25016 657 25050
rect 694 25016 728 25050
rect 764 25016 798 25050
rect 834 25016 868 25050
rect 518 24908 552 24942
rect 518 24837 552 24871
rect 518 24766 552 24800
rect 518 24695 552 24729
rect 518 24624 552 24658
rect 518 24553 552 24587
rect 518 24482 552 24516
rect 518 24411 552 24445
rect 518 24340 552 24374
rect 518 24269 552 24303
rect 518 24187 552 24221
rect 518 24114 552 24148
rect 518 24041 552 24075
rect 518 23967 552 24001
rect 518 23893 552 23927
rect 1758 24187 1792 24221
rect 1758 24113 1792 24147
rect 1758 24039 1792 24073
rect 1758 23965 1792 23999
rect 518 23819 552 23853
rect 1758 23891 1792 23925
rect 1758 23818 1792 23852
rect 518 23745 552 23779
rect 518 23671 552 23705
rect 518 23597 552 23631
rect 518 23523 552 23557
rect 1758 23745 1792 23779
rect 1758 23672 1792 23706
rect 1758 23599 1792 23633
rect 1758 23526 1792 23560
rect 518 23449 552 23483
rect 518 23375 552 23409
rect 1758 23453 1792 23487
rect 620 23341 654 23375
rect 689 23341 723 23375
rect 758 23341 792 23375
rect 827 23341 861 23375
rect 896 23341 930 23375
rect 965 23341 999 23375
rect 1034 23341 1068 23375
rect 1103 23341 1137 23375
rect 1172 23341 1206 23375
rect 1241 23341 1275 23375
rect 1310 23341 1344 23375
rect 1379 23341 1413 23375
rect 1448 23341 1482 23375
rect 1517 23341 1551 23375
rect 1586 23341 1620 23375
rect 1655 23341 1689 23375
rect 1724 23341 1758 23375
rect 21 22725 55 22759
rect 90 22725 124 22759
rect 159 22725 193 22759
rect 228 22725 262 22759
rect 297 22725 331 22759
rect 366 22725 400 22759
rect 435 22725 469 22759
rect 504 22725 538 22759
rect 573 22725 607 22759
rect 642 22725 676 22759
rect 711 22725 745 22759
rect -184 22691 -82 22725
rect -116 22657 -82 22691
rect -47 22657 -13 22691
rect 22 22657 56 22691
rect 91 22657 125 22691
rect 160 22657 194 22691
rect 229 22657 263 22691
rect 298 22657 332 22691
rect 367 22657 401 22691
rect 436 22657 470 22691
rect 505 22657 539 22691
rect 574 22657 608 22691
rect 643 22657 677 22691
rect 712 22657 746 22691
rect 780 22657 2174 22759
rect -150 22589 -116 22623
rect -80 22589 -46 22623
rect -10 22589 24 22623
rect 60 22589 94 22623
rect 130 22589 164 22623
rect 200 22589 234 22623
rect 270 22589 304 22623
rect 340 22589 374 22623
rect 410 22589 444 22623
rect 480 22589 514 22623
rect 550 22589 584 22623
rect 620 22589 654 22623
rect 690 22589 724 22623
rect 760 22589 794 22623
rect 829 22589 863 22623
rect 898 22589 932 22623
rect 967 22589 1001 22623
rect 1036 22589 1070 22623
rect 1105 22589 1139 22623
rect 1174 22589 1208 22623
rect 1243 22589 1277 22623
rect 1312 22589 1346 22623
rect 1381 22589 1415 22623
rect 1450 22589 1484 22623
rect 1519 22589 1553 22623
rect 1588 22589 1622 22623
rect 1657 22589 1691 22623
rect 1726 22589 1760 22623
rect 1795 22589 1829 22623
rect 1864 22589 1898 22623
rect 1933 22589 1967 22623
rect 2002 22589 2036 22623
rect 2071 22589 2105 22623
rect 2140 22589 2174 22623
<< poly >>
rect 4396 27009 4530 27025
rect 4396 26975 4412 27009
rect 4446 26975 4480 27009
rect 4514 26975 4530 27009
rect 4396 26959 4530 26975
rect 4808 27009 4942 27025
rect 4808 26975 4824 27009
rect 4858 26975 4892 27009
rect 4926 26975 4942 27009
rect 4808 26959 4942 26975
rect 5220 27009 5354 27025
rect 5220 26975 5236 27009
rect 5270 26975 5304 27009
rect 5338 26975 5354 27009
rect 5220 26959 5354 26975
rect 5632 27009 5766 27025
rect 5632 26975 5648 27009
rect 5682 26975 5716 27009
rect 5750 26975 5766 27009
rect 5632 26959 5766 26975
rect 6044 27009 6178 27025
rect 6044 26975 6060 27009
rect 6094 26975 6128 27009
rect 6162 26975 6178 27009
rect 6044 26959 6178 26975
rect 6456 27009 6590 27025
rect 6456 26975 6472 27009
rect 6506 26975 6540 27009
rect 6574 26975 6590 27009
rect 6456 26959 6590 26975
rect 6868 27009 7002 27025
rect 6868 26975 6884 27009
rect 6918 26975 6952 27009
rect 6986 26975 7002 27009
rect 6868 26959 7002 26975
rect 7280 27009 7414 27025
rect 7280 26975 7296 27009
rect 7330 26975 7364 27009
rect 7398 26975 7414 27009
rect 7280 26959 7414 26975
rect 7692 27009 7826 27025
rect 7692 26975 7708 27009
rect 7742 26975 7776 27009
rect 7810 26975 7826 27009
rect 7692 26959 7826 26975
rect 8104 27009 8238 27025
rect 8104 26975 8120 27009
rect 8154 26975 8188 27009
rect 8222 26975 8238 27009
rect 8104 26959 8238 26975
rect 8516 27009 8650 27025
rect 8516 26975 8532 27009
rect 8566 26975 8600 27009
rect 8634 26975 8650 27009
rect 8516 26959 8650 26975
rect 8928 27009 9062 27025
rect 8928 26975 8944 27009
rect 8978 26975 9012 27009
rect 9046 26975 9062 27009
rect 8928 26959 9062 26975
rect 9340 27009 9474 27025
rect 9340 26975 9356 27009
rect 9390 26975 9424 27009
rect 9458 26975 9474 27009
rect 9340 26959 9474 26975
rect 9752 27009 9886 27025
rect 9752 26975 9768 27009
rect 9802 26975 9836 27009
rect 9870 26975 9886 27009
rect 9752 26959 9886 26975
rect 10164 27009 10298 27025
rect 10164 26975 10180 27009
rect 10214 26975 10248 27009
rect 10282 26975 10298 27009
rect 10164 26959 10298 26975
rect 10576 27009 10710 27025
rect 10576 26975 10592 27009
rect 10626 26975 10660 27009
rect 10694 26975 10710 27009
rect 10576 26959 10710 26975
rect 10988 27009 11122 27025
rect 10988 26975 11004 27009
rect 11038 26975 11072 27009
rect 11106 26975 11122 27009
rect 10988 26959 11122 26975
rect 11400 27009 11534 27025
rect 11400 26975 11416 27009
rect 11450 26975 11484 27009
rect 11518 26975 11534 27009
rect 11400 26959 11534 26975
rect 11812 27009 11946 27025
rect 11812 26975 11828 27009
rect 11862 26975 11896 27009
rect 11930 26975 11946 27009
rect 11812 26959 11946 26975
rect 12224 27009 12358 27025
rect 12224 26975 12240 27009
rect 12274 26975 12308 27009
rect 12342 26975 12358 27009
rect 12224 26959 12358 26975
rect 12636 27009 12770 27025
rect 12636 26975 12652 27009
rect 12686 26975 12720 27009
rect 12754 26975 12770 27009
rect 12636 26959 12770 26975
rect 13048 27009 13182 27025
rect 13048 26975 13064 27009
rect 13098 26975 13132 27009
rect 13166 26975 13182 27009
rect 13048 26959 13182 26975
rect 13460 27009 13594 27025
rect 13460 26975 13476 27009
rect 13510 26975 13544 27009
rect 13578 26975 13594 27009
rect 13460 26959 13594 26975
rect 13872 27009 14006 27025
rect 13872 26975 13888 27009
rect 13922 26975 13956 27009
rect 13990 26975 14006 27009
rect 13872 26959 14006 26975
rect 14284 27009 14418 27025
rect 14284 26975 14300 27009
rect 14334 26975 14368 27009
rect 14402 26975 14418 27009
rect 14284 26959 14418 26975
rect 14696 27009 14830 27025
rect 14696 26975 14712 27009
rect 14746 26975 14780 27009
rect 14814 26975 14830 27009
rect 14696 26959 14830 26975
rect 2754 25475 2854 25491
rect 2754 25441 2787 25475
rect 2821 25441 2854 25475
rect 2754 25423 2854 25441
rect 574 24176 646 24192
rect 574 24142 590 24176
rect 624 24142 646 24176
rect 574 24108 646 24142
rect 574 24074 590 24108
rect 624 24092 646 24108
rect 624 24074 640 24092
rect 574 24040 640 24074
rect 574 24006 590 24040
rect 624 24036 640 24040
rect 624 24006 646 24036
rect 574 23972 646 24006
rect 574 23938 590 23972
rect 624 23938 646 23972
rect 574 23936 646 23938
rect 574 23922 640 23936
rect 574 23770 640 23784
rect 574 23768 646 23770
rect 574 23734 590 23768
rect 624 23734 646 23768
rect 574 23700 646 23734
rect 574 23666 590 23700
rect 624 23670 646 23700
rect 4396 23779 4530 23795
rect 4396 23745 4412 23779
rect 4446 23745 4480 23779
rect 4514 23745 4530 23779
rect 4396 23729 4530 23745
rect 4808 23779 4942 23795
rect 4808 23745 4824 23779
rect 4858 23745 4892 23779
rect 4926 23745 4942 23779
rect 4808 23729 4942 23745
rect 5220 23779 5354 23795
rect 5220 23745 5236 23779
rect 5270 23745 5304 23779
rect 5338 23745 5354 23779
rect 5220 23729 5354 23745
rect 5632 23779 5766 23795
rect 5632 23745 5648 23779
rect 5682 23745 5716 23779
rect 5750 23745 5766 23779
rect 5632 23729 5766 23745
rect 6044 23779 6178 23795
rect 6044 23745 6060 23779
rect 6094 23745 6128 23779
rect 6162 23745 6178 23779
rect 6044 23729 6178 23745
rect 6456 23779 6590 23795
rect 6456 23745 6472 23779
rect 6506 23745 6540 23779
rect 6574 23745 6590 23779
rect 6456 23729 6590 23745
rect 6868 23779 7002 23795
rect 6868 23745 6884 23779
rect 6918 23745 6952 23779
rect 6986 23745 7002 23779
rect 6868 23729 7002 23745
rect 7280 23779 7414 23795
rect 7280 23745 7296 23779
rect 7330 23745 7364 23779
rect 7398 23745 7414 23779
rect 7280 23729 7414 23745
rect 7692 23779 7826 23795
rect 7692 23745 7708 23779
rect 7742 23745 7776 23779
rect 7810 23745 7826 23779
rect 7692 23729 7826 23745
rect 8104 23779 8238 23795
rect 8104 23745 8120 23779
rect 8154 23745 8188 23779
rect 8222 23745 8238 23779
rect 8104 23729 8238 23745
rect 8516 23779 8650 23795
rect 8516 23745 8532 23779
rect 8566 23745 8600 23779
rect 8634 23745 8650 23779
rect 8516 23729 8650 23745
rect 8928 23779 9062 23795
rect 8928 23745 8944 23779
rect 8978 23745 9012 23779
rect 9046 23745 9062 23779
rect 8928 23729 9062 23745
rect 9340 23779 9474 23795
rect 9340 23745 9356 23779
rect 9390 23745 9424 23779
rect 9458 23745 9474 23779
rect 9340 23729 9474 23745
rect 9752 23779 9886 23795
rect 9752 23745 9768 23779
rect 9802 23745 9836 23779
rect 9870 23745 9886 23779
rect 9752 23729 9886 23745
rect 10164 23779 10298 23795
rect 10164 23745 10180 23779
rect 10214 23745 10248 23779
rect 10282 23745 10298 23779
rect 10164 23729 10298 23745
rect 10576 23779 10710 23795
rect 10576 23745 10592 23779
rect 10626 23745 10660 23779
rect 10694 23745 10710 23779
rect 10576 23729 10710 23745
rect 10988 23779 11122 23795
rect 10988 23745 11004 23779
rect 11038 23745 11072 23779
rect 11106 23745 11122 23779
rect 10988 23729 11122 23745
rect 11400 23779 11534 23795
rect 11400 23745 11416 23779
rect 11450 23745 11484 23779
rect 11518 23745 11534 23779
rect 11400 23729 11534 23745
rect 11812 23779 11946 23795
rect 11812 23745 11828 23779
rect 11862 23745 11896 23779
rect 11930 23745 11946 23779
rect 11812 23729 11946 23745
rect 12224 23779 12358 23795
rect 12224 23745 12240 23779
rect 12274 23745 12308 23779
rect 12342 23745 12358 23779
rect 12224 23729 12358 23745
rect 12636 23779 12770 23795
rect 12636 23745 12652 23779
rect 12686 23745 12720 23779
rect 12754 23745 12770 23779
rect 12636 23729 12770 23745
rect 13048 23779 13182 23795
rect 13048 23745 13064 23779
rect 13098 23745 13132 23779
rect 13166 23745 13182 23779
rect 13048 23729 13182 23745
rect 13460 23779 13594 23795
rect 13460 23745 13476 23779
rect 13510 23745 13544 23779
rect 13578 23745 13594 23779
rect 13460 23729 13594 23745
rect 13872 23779 14006 23795
rect 13872 23745 13888 23779
rect 13922 23745 13956 23779
rect 13990 23745 14006 23779
rect 13872 23729 14006 23745
rect 14284 23779 14418 23795
rect 14284 23745 14300 23779
rect 14334 23745 14368 23779
rect 14402 23745 14418 23779
rect 14284 23729 14418 23745
rect 14696 23779 14830 23795
rect 14696 23745 14712 23779
rect 14746 23745 14780 23779
rect 14814 23745 14830 23779
rect 14696 23729 14830 23745
rect 15108 23779 15242 23795
rect 15108 23745 15124 23779
rect 15158 23745 15192 23779
rect 15226 23745 15242 23779
rect 15108 23729 15242 23745
rect 15520 23779 15654 23795
rect 15520 23745 15536 23779
rect 15570 23745 15604 23779
rect 15638 23745 15654 23779
rect 15520 23729 15654 23745
rect 15932 23779 16066 23795
rect 15932 23745 15948 23779
rect 15982 23745 16016 23779
rect 16050 23745 16066 23779
rect 15932 23729 16066 23745
rect 16344 23779 16478 23795
rect 16344 23745 16360 23779
rect 16394 23745 16428 23779
rect 16462 23745 16478 23779
rect 16344 23729 16478 23745
rect 16756 23779 16890 23795
rect 16756 23745 16772 23779
rect 16806 23745 16840 23779
rect 16874 23745 16890 23779
rect 16756 23729 16890 23745
rect 17168 23779 17302 23795
rect 17168 23745 17184 23779
rect 17218 23745 17252 23779
rect 17286 23745 17302 23779
rect 17168 23729 17302 23745
rect 624 23666 640 23670
rect 574 23632 640 23666
rect 574 23598 590 23632
rect 624 23614 640 23632
rect 624 23598 646 23614
rect 574 23564 646 23598
rect 574 23530 590 23564
rect 624 23530 646 23564
rect 574 23514 646 23530
rect 2754 23265 2854 23283
rect 2754 23231 2787 23265
rect 2821 23231 2854 23265
rect 2754 23215 2854 23231
rect 374 4940 440 4956
rect 374 4906 390 4940
rect 424 4906 440 4940
rect 374 4872 440 4906
rect 374 4838 390 4872
rect 424 4838 440 4872
rect 374 4804 440 4838
rect 374 4770 390 4804
rect 424 4770 440 4804
rect 374 4736 440 4770
rect 374 4702 390 4736
rect 424 4702 440 4736
rect 374 4686 440 4702
rect 374 4532 440 4548
rect 374 4498 390 4532
rect 424 4498 440 4532
rect 374 4464 440 4498
rect 374 4430 390 4464
rect 424 4430 440 4464
rect 374 4396 440 4430
rect 374 4362 390 4396
rect 424 4362 440 4396
rect 374 4328 440 4362
rect 374 4294 390 4328
rect 424 4294 440 4328
rect 374 4278 440 4294
<< polycont >>
rect 4412 26975 4446 27009
rect 4480 26975 4514 27009
rect 4824 26975 4858 27009
rect 4892 26975 4926 27009
rect 5236 26975 5270 27009
rect 5304 26975 5338 27009
rect 5648 26975 5682 27009
rect 5716 26975 5750 27009
rect 6060 26975 6094 27009
rect 6128 26975 6162 27009
rect 6472 26975 6506 27009
rect 6540 26975 6574 27009
rect 6884 26975 6918 27009
rect 6952 26975 6986 27009
rect 7296 26975 7330 27009
rect 7364 26975 7398 27009
rect 7708 26975 7742 27009
rect 7776 26975 7810 27009
rect 8120 26975 8154 27009
rect 8188 26975 8222 27009
rect 8532 26975 8566 27009
rect 8600 26975 8634 27009
rect 8944 26975 8978 27009
rect 9012 26975 9046 27009
rect 9356 26975 9390 27009
rect 9424 26975 9458 27009
rect 9768 26975 9802 27009
rect 9836 26975 9870 27009
rect 10180 26975 10214 27009
rect 10248 26975 10282 27009
rect 10592 26975 10626 27009
rect 10660 26975 10694 27009
rect 11004 26975 11038 27009
rect 11072 26975 11106 27009
rect 11416 26975 11450 27009
rect 11484 26975 11518 27009
rect 11828 26975 11862 27009
rect 11896 26975 11930 27009
rect 12240 26975 12274 27009
rect 12308 26975 12342 27009
rect 12652 26975 12686 27009
rect 12720 26975 12754 27009
rect 13064 26975 13098 27009
rect 13132 26975 13166 27009
rect 13476 26975 13510 27009
rect 13544 26975 13578 27009
rect 13888 26975 13922 27009
rect 13956 26975 13990 27009
rect 14300 26975 14334 27009
rect 14368 26975 14402 27009
rect 14712 26975 14746 27009
rect 14780 26975 14814 27009
rect 2787 25441 2821 25475
rect 590 24142 624 24176
rect 590 24074 624 24108
rect 590 24006 624 24040
rect 590 23938 624 23972
rect 590 23734 624 23768
rect 590 23666 624 23700
rect 4412 23745 4446 23779
rect 4480 23745 4514 23779
rect 4824 23745 4858 23779
rect 4892 23745 4926 23779
rect 5236 23745 5270 23779
rect 5304 23745 5338 23779
rect 5648 23745 5682 23779
rect 5716 23745 5750 23779
rect 6060 23745 6094 23779
rect 6128 23745 6162 23779
rect 6472 23745 6506 23779
rect 6540 23745 6574 23779
rect 6884 23745 6918 23779
rect 6952 23745 6986 23779
rect 7296 23745 7330 23779
rect 7364 23745 7398 23779
rect 7708 23745 7742 23779
rect 7776 23745 7810 23779
rect 8120 23745 8154 23779
rect 8188 23745 8222 23779
rect 8532 23745 8566 23779
rect 8600 23745 8634 23779
rect 8944 23745 8978 23779
rect 9012 23745 9046 23779
rect 9356 23745 9390 23779
rect 9424 23745 9458 23779
rect 9768 23745 9802 23779
rect 9836 23745 9870 23779
rect 10180 23745 10214 23779
rect 10248 23745 10282 23779
rect 10592 23745 10626 23779
rect 10660 23745 10694 23779
rect 11004 23745 11038 23779
rect 11072 23745 11106 23779
rect 11416 23745 11450 23779
rect 11484 23745 11518 23779
rect 11828 23745 11862 23779
rect 11896 23745 11930 23779
rect 12240 23745 12274 23779
rect 12308 23745 12342 23779
rect 12652 23745 12686 23779
rect 12720 23745 12754 23779
rect 13064 23745 13098 23779
rect 13132 23745 13166 23779
rect 13476 23745 13510 23779
rect 13544 23745 13578 23779
rect 13888 23745 13922 23779
rect 13956 23745 13990 23779
rect 14300 23745 14334 23779
rect 14368 23745 14402 23779
rect 14712 23745 14746 23779
rect 14780 23745 14814 23779
rect 15124 23745 15158 23779
rect 15192 23745 15226 23779
rect 15536 23745 15570 23779
rect 15604 23745 15638 23779
rect 15948 23745 15982 23779
rect 16016 23745 16050 23779
rect 16360 23745 16394 23779
rect 16428 23745 16462 23779
rect 16772 23745 16806 23779
rect 16840 23745 16874 23779
rect 17184 23745 17218 23779
rect 17252 23745 17286 23779
rect 590 23598 624 23632
rect 590 23530 624 23564
rect 2787 23231 2821 23265
rect 390 4906 424 4940
rect 390 4838 424 4872
rect 390 4770 424 4804
rect 390 4702 424 4736
rect 390 4498 424 4532
rect 390 4430 424 4464
rect 390 4362 424 4396
rect 390 4294 424 4328
<< locali >>
rect -184 27729 -14 27741
rect -184 27717 -152 27729
rect -118 27717 -80 27729
rect -46 27717 -14 27729
rect -118 27695 -116 27717
rect -150 27683 -116 27695
rect -82 27695 -80 27717
rect -82 27683 -48 27695
rect -184 27656 -14 27683
rect -184 27648 -152 27656
rect -118 27648 -80 27656
rect -46 27648 -14 27656
rect -118 27622 -116 27648
rect -150 27614 -116 27622
rect -82 27622 -80 27648
rect -82 27614 -48 27622
rect -184 27583 -14 27614
rect -184 27579 -152 27583
rect -118 27579 -80 27583
rect -46 27579 -14 27583
rect -118 27549 -116 27579
rect -150 27545 -116 27549
rect -82 27549 -80 27579
rect -82 27545 -48 27549
rect -184 27510 -14 27545
rect -118 27476 -116 27510
rect -82 27476 -80 27510
rect -184 27441 -14 27476
rect -150 27437 -116 27441
rect -118 27407 -116 27437
rect -82 27437 -48 27441
rect -82 27407 -80 27437
rect -184 27403 -152 27407
rect -118 27403 -80 27407
rect -46 27403 -14 27407
rect -184 27372 -14 27403
rect -150 27364 -116 27372
rect -118 27338 -116 27364
rect -82 27364 -48 27372
rect -82 27338 -80 27364
rect -184 27330 -152 27338
rect -118 27330 -80 27338
rect -46 27330 -14 27338
rect -184 27303 -14 27330
rect -150 27291 -116 27303
rect -118 27269 -116 27291
rect -82 27291 -48 27303
rect -82 27269 -80 27291
rect -184 27257 -152 27269
rect -118 27257 -80 27269
rect -46 27257 -14 27269
rect -184 27234 -14 27257
rect -150 27218 -116 27234
rect -118 27200 -116 27218
rect -82 27218 -48 27234
rect -82 27200 -80 27218
rect -184 27184 -152 27200
rect -118 27184 -80 27200
rect -46 27184 -14 27200
rect -184 27165 -14 27184
rect -150 27145 -116 27165
rect -118 27131 -116 27145
rect -82 27145 -48 27165
rect -82 27131 -80 27145
rect -184 27111 -152 27131
rect -118 27111 -80 27131
rect -46 27111 -14 27131
rect -184 27096 -14 27111
rect -150 27072 -116 27096
rect -118 27062 -116 27072
rect -82 27072 -48 27096
rect -82 27062 -80 27072
rect -184 27038 -152 27062
rect -118 27038 -80 27062
rect -46 27038 -14 27062
rect -184 27027 -14 27038
rect -150 26999 -116 27027
rect -118 26993 -116 26999
rect -82 26999 -48 27027
rect -82 26993 -80 26999
rect -184 26965 -152 26993
rect -118 26965 -80 26993
rect -46 26965 -14 26993
rect -184 26958 -14 26965
rect -150 26926 -116 26958
rect -118 26924 -116 26926
rect -82 26926 -48 26958
rect -82 26924 -80 26926
rect -184 26892 -152 26924
rect -118 26892 -80 26924
rect -46 26892 -14 26924
rect -184 26889 -14 26892
rect -150 26855 -116 26889
rect -82 26855 -48 26889
rect -184 26853 -14 26855
rect -184 26820 -152 26853
rect -118 26820 -80 26853
rect -46 26820 -14 26853
rect -118 26819 -116 26820
rect -150 26786 -116 26819
rect -82 26819 -80 26820
rect -82 26786 -48 26819
rect -184 26780 -14 26786
rect -184 26751 -152 26780
rect -118 26751 -80 26780
rect -46 26751 -14 26780
rect -118 26746 -116 26751
rect -150 26717 -116 26746
rect -82 26746 -80 26751
rect -82 26717 -48 26746
rect -184 26707 -14 26717
rect -184 26682 -152 26707
rect -118 26682 -80 26707
rect -46 26682 -14 26707
rect -118 26673 -116 26682
rect -150 26648 -116 26673
rect -82 26673 -80 26682
rect -82 26648 -48 26673
rect -184 26634 -14 26648
rect -184 26613 -152 26634
rect -118 26613 -80 26634
rect -46 26613 -14 26634
rect -118 26600 -116 26613
rect -150 26579 -116 26600
rect -82 26600 -80 26613
rect -82 26579 -48 26600
rect -184 26561 -14 26579
rect -184 26544 -152 26561
rect -118 26544 -80 26561
rect -46 26544 -14 26561
rect -118 26527 -116 26544
rect -150 26510 -116 26527
rect -82 26527 -80 26544
rect -82 26510 -48 26527
rect -184 26488 -14 26510
rect -184 26475 -152 26488
rect -118 26475 -80 26488
rect -46 26475 -14 26488
rect -118 26454 -116 26475
rect -150 26441 -116 26454
rect -82 26454 -80 26475
rect -82 26441 -48 26454
rect -184 26415 -14 26441
rect -184 26406 -152 26415
rect -118 26406 -80 26415
rect -46 26406 -14 26415
rect -118 26381 -116 26406
rect -150 26372 -116 26381
rect -82 26381 -80 26406
rect -82 26372 -48 26381
rect -184 26342 -14 26372
rect -184 26337 -152 26342
rect -118 26337 -80 26342
rect -46 26337 -14 26342
rect -118 26308 -116 26337
rect -150 26303 -116 26308
rect -82 26308 -80 26337
rect -82 26303 -48 26308
rect -184 26269 -14 26303
rect -184 26268 -152 26269
rect -118 26268 -80 26269
rect -46 26268 -14 26269
rect -118 26235 -116 26268
rect -150 26234 -116 26235
rect -82 26235 -80 26268
rect -82 26234 -48 26235
rect -184 26199 -14 26234
rect -150 26196 -116 26199
rect -118 26165 -116 26196
rect -82 26196 -48 26199
rect -82 26165 -80 26196
rect -184 26162 -152 26165
rect -118 26162 -80 26165
rect -46 26162 -14 26165
rect -184 26130 -14 26162
rect -150 26123 -116 26130
rect -118 26096 -116 26123
rect -82 26123 -48 26130
rect -82 26096 -80 26123
rect -184 26089 -152 26096
rect -118 26089 -80 26096
rect -46 26089 -14 26096
rect -184 26061 -14 26089
rect -150 26050 -116 26061
rect -118 26027 -116 26050
rect -82 26050 -48 26061
rect -82 26027 -80 26050
rect -184 26016 -152 26027
rect -118 26016 -80 26027
rect -46 26016 -14 26027
rect -184 25992 -14 26016
rect -150 25977 -116 25992
rect -118 25958 -116 25977
rect -82 25977 -48 25992
rect -82 25958 -80 25977
rect -184 25943 -152 25958
rect -118 25943 -80 25958
rect -46 25943 -14 25958
rect -184 25923 -14 25943
rect -150 25904 -116 25923
rect -118 25889 -116 25904
rect -82 25904 -48 25923
rect -82 25889 -80 25904
rect -184 25870 -152 25889
rect -118 25870 -80 25889
rect -46 25870 -14 25889
rect -184 25854 -14 25870
rect -150 25831 -116 25854
rect -118 25820 -116 25831
rect -82 25831 -48 25854
rect -82 25820 -80 25831
rect -184 25797 -152 25820
rect -118 25797 -80 25820
rect -46 25797 -14 25820
rect -184 25785 -14 25797
rect -150 25758 -116 25785
rect -118 25751 -116 25758
rect -82 25758 -48 25785
rect -82 25751 -80 25758
rect -184 25724 -152 25751
rect -118 25724 -80 25751
rect -46 25724 -14 25751
rect -184 25717 -14 25724
rect -150 25716 -14 25717
rect -150 25685 -116 25716
rect -184 25651 -152 25683
rect -118 25682 -116 25685
rect -82 25685 -48 25716
rect -82 25682 -80 25685
rect -118 25651 -80 25682
rect -46 25651 -14 25682
rect -184 25649 -14 25651
rect -150 25647 -14 25649
rect -150 25615 -116 25647
rect -184 25613 -116 25615
rect -82 25613 -48 25647
rect -184 25612 -14 25613
rect -184 25581 -152 25612
rect -118 25578 -80 25612
rect -46 25578 -14 25612
rect -150 25547 -116 25578
rect -184 25544 -116 25547
rect -82 25544 -48 25578
rect -184 25539 -14 25544
rect -184 25513 -152 25539
rect -118 25509 -80 25539
rect -46 25509 -14 25539
rect -118 25505 -116 25509
rect -150 25479 -116 25505
rect -184 25475 -116 25479
rect -82 25505 -80 25509
rect -82 25475 -48 25505
rect -184 25466 -14 25475
rect -184 25445 -152 25466
rect -118 25440 -80 25466
rect -46 25440 -14 25466
rect -118 25432 -116 25440
rect -150 25411 -116 25432
rect -184 25406 -116 25411
rect -82 25432 -80 25440
rect -82 25406 -48 25432
rect -184 25393 -14 25406
rect -184 25377 -152 25393
rect -118 25371 -80 25393
rect -46 25371 -14 25393
rect -118 25359 -116 25371
rect -150 25343 -116 25359
rect -184 25337 -116 25343
rect -82 25359 -80 25371
rect -82 25337 -48 25359
rect -184 25320 -14 25337
rect -184 25309 -152 25320
rect -118 25302 -80 25320
rect -46 25302 -14 25320
rect -118 25286 -116 25302
rect -150 25275 -116 25286
rect -184 25268 -116 25275
rect -82 25286 -80 25302
rect -82 25268 -48 25286
rect -184 25247 -14 25268
rect -184 25241 -152 25247
rect -118 25233 -80 25247
rect -46 25233 -14 25247
rect -118 25213 -116 25233
rect -150 25207 -116 25213
rect -184 25199 -116 25207
rect -82 25213 -80 25233
rect -82 25199 -48 25213
rect -184 25175 -14 25199
rect -184 25174 -80 25175
rect -184 25173 -152 25174
rect -118 25164 -80 25174
rect -46 25164 -14 25175
rect -118 25140 -116 25164
rect -150 25139 -116 25140
rect -184 25130 -116 25139
rect -82 25141 -80 25164
rect -82 25130 -48 25141
rect -184 25105 -14 25130
rect -150 25103 -14 25105
rect -150 25101 -80 25103
rect -118 25095 -80 25101
rect -46 25095 -14 25103
rect -184 25067 -152 25071
rect -118 25067 -116 25095
rect -184 25061 -116 25067
rect -82 25069 -80 25095
rect -82 25061 -48 25069
rect -184 25037 -14 25061
rect -150 25031 -14 25037
rect -150 25028 -80 25031
rect -118 25026 -80 25028
rect -46 25026 -14 25031
rect -184 24994 -152 25003
rect -118 24994 -116 25026
rect -184 24992 -116 24994
rect -82 24997 -80 25026
rect -82 24992 -48 24997
rect -184 24969 -14 24992
rect -150 24959 -14 24969
rect -150 24957 -80 24959
rect -46 24957 -14 24959
rect -150 24955 -116 24957
rect -184 24921 -152 24935
rect -118 24923 -116 24955
rect -82 24925 -80 24957
rect -82 24923 -48 24925
rect -118 24921 -14 24923
rect -184 24901 -14 24921
rect -150 24888 -14 24901
rect -150 24882 -116 24888
rect -184 24848 -152 24867
rect -118 24854 -116 24882
rect -82 24887 -48 24888
rect -82 24854 -80 24887
rect -118 24853 -80 24854
rect -46 24853 -14 24854
rect -118 24848 -14 24853
rect -184 24833 -14 24848
rect -150 24819 -14 24833
rect -150 24809 -116 24819
rect -184 24775 -152 24799
rect -118 24785 -116 24809
rect -82 24815 -48 24819
rect -82 24785 -80 24815
rect -118 24781 -80 24785
rect -46 24781 -14 24785
rect -118 24775 -14 24781
rect -184 24765 -14 24775
rect -150 24750 -14 24765
rect -150 24736 -116 24750
rect -184 24702 -152 24731
rect -118 24716 -116 24736
rect -82 24743 -48 24750
rect -82 24716 -80 24743
rect -118 24709 -80 24716
rect -46 24709 -14 24716
rect -118 24702 -14 24709
rect -184 24697 -14 24702
rect -150 24681 -14 24697
rect -150 24663 -116 24681
rect -184 24629 -152 24663
rect -118 24647 -116 24663
rect -82 24671 -48 24681
rect -82 24647 -80 24671
rect -118 24637 -80 24647
rect -46 24637 -14 24647
rect -118 24629 -14 24637
rect -150 24612 -14 24629
rect -150 24595 -116 24612
rect -184 24590 -116 24595
rect -184 24561 -152 24590
rect -118 24578 -116 24590
rect -82 24599 -48 24612
rect -82 24578 -80 24599
rect -118 24565 -80 24578
rect -46 24565 -14 24578
rect -118 24556 -14 24565
rect -150 24543 -14 24556
rect -150 24527 -116 24543
rect -184 24517 -116 24527
rect -184 24493 -152 24517
rect -118 24509 -116 24517
rect -82 24527 -48 24543
rect -82 24509 -80 24527
rect -118 24493 -80 24509
rect -46 24493 -14 24509
rect -118 24483 -14 24493
rect -150 24474 -14 24483
rect -150 24459 -116 24474
rect -184 24444 -116 24459
rect -184 24425 -152 24444
rect -118 24440 -116 24444
rect -82 24455 -48 24474
rect -82 24440 -80 24455
rect -118 24421 -80 24440
rect -46 24421 -14 24440
rect -118 24410 -14 24421
rect -150 24405 -14 24410
rect -150 24391 -116 24405
rect -184 24371 -116 24391
rect -82 24383 -48 24405
rect -82 24371 -80 24383
rect -184 24357 -152 24371
rect -118 24349 -80 24371
rect -46 24349 -14 24371
rect -118 24337 -14 24349
rect -150 24336 -14 24337
rect -150 24323 -116 24336
rect -184 24302 -116 24323
rect -82 24311 -48 24336
rect -82 24302 -80 24311
rect -184 24298 -80 24302
rect -184 24289 -152 24298
rect -118 24277 -80 24298
rect -46 24277 -14 24302
rect -118 24267 -14 24277
rect -118 24264 -116 24267
rect -150 24255 -116 24264
rect -184 24233 -116 24255
rect -82 24239 -48 24267
rect -82 24233 -80 24239
rect -184 24225 -80 24233
rect -184 24221 -152 24225
rect -118 24205 -80 24225
rect -46 24205 -14 24233
rect -118 24198 -14 24205
rect -118 24191 -116 24198
rect -150 24187 -116 24191
rect -184 24164 -116 24187
rect -82 24167 -48 24198
rect -82 24164 -80 24167
rect -184 24153 -80 24164
rect -150 24152 -80 24153
rect -118 24133 -80 24152
rect -46 24133 -14 24164
rect -118 24129 -14 24133
rect -184 24118 -152 24119
rect -118 24118 -116 24129
rect -184 24095 -116 24118
rect -82 24095 -48 24129
rect -184 24085 -80 24095
rect -150 24079 -80 24085
rect -118 24061 -80 24079
rect -46 24061 -14 24095
rect -118 24060 -14 24061
rect -184 24045 -152 24051
rect -118 24045 -116 24060
rect -184 24026 -116 24045
rect -82 24026 -48 24060
rect -184 24023 -14 24026
rect -184 24017 -80 24023
rect -150 24006 -80 24017
rect -118 23991 -80 24006
rect -46 23991 -14 24023
rect -184 23972 -152 23983
rect -118 23972 -116 23991
rect -184 23957 -116 23972
rect -82 23989 -80 23991
rect -82 23957 -48 23989
rect -184 23951 -14 23957
rect -184 23949 -80 23951
rect -150 23933 -80 23949
rect -118 23922 -80 23933
rect -46 23922 -14 23951
rect -184 23899 -152 23915
rect -118 23899 -116 23922
rect -184 23888 -116 23899
rect -82 23917 -80 23922
rect -82 23888 -48 23917
rect -184 23881 -14 23888
rect -150 23879 -14 23881
rect -150 23860 -80 23879
rect -118 23853 -80 23860
rect -46 23853 -14 23879
rect -184 23826 -152 23847
rect -118 23826 -116 23853
rect -184 23819 -116 23826
rect -82 23845 -80 23853
rect -82 23819 -48 23845
rect -184 23813 -14 23819
rect -150 23807 -14 23813
rect -150 23787 -80 23807
rect -118 23784 -80 23787
rect -46 23784 -14 23807
rect -184 23753 -152 23779
rect -118 23753 -116 23784
rect -184 23750 -116 23753
rect -82 23773 -80 23784
rect -82 23750 -48 23773
rect -184 23745 -14 23750
rect -150 23735 -14 23745
rect -150 23715 -80 23735
rect -46 23715 -14 23735
rect -150 23714 -116 23715
rect -184 23680 -152 23711
rect -118 23681 -116 23714
rect -82 23701 -80 23715
rect -82 23681 -48 23701
rect -118 23680 -14 23681
rect -184 23677 -14 23680
rect -150 23663 -14 23677
rect -150 23646 -80 23663
rect -46 23646 -14 23663
rect -150 23643 -116 23646
rect -184 23641 -116 23643
rect -184 23609 -152 23641
rect -118 23612 -116 23641
rect -82 23629 -80 23646
rect -82 23612 -48 23629
rect -118 23607 -14 23612
rect -150 23591 -14 23607
rect -150 23577 -80 23591
rect -46 23577 -14 23591
rect -150 23575 -116 23577
rect -184 23568 -116 23575
rect -184 23541 -152 23568
rect -118 23543 -116 23568
rect -82 23557 -80 23577
rect -82 23543 -48 23557
rect -118 23534 -14 23543
rect -150 23519 -14 23534
rect -150 23508 -80 23519
rect -46 23508 -14 23519
rect -150 23507 -116 23508
rect -184 23495 -116 23507
rect -184 23473 -152 23495
rect -118 23474 -116 23495
rect -82 23485 -80 23508
rect -82 23474 -48 23485
rect -118 23461 -14 23474
rect -150 23447 -14 23461
rect -150 23439 -80 23447
rect -46 23439 -14 23447
rect 196 27707 230 27741
rect 264 27709 299 27741
rect 333 27709 368 27741
rect 402 27709 437 27741
rect 471 27709 506 27741
rect 540 27709 575 27741
rect 609 27709 644 27741
rect 264 27707 266 27709
rect 333 27707 341 27709
rect 402 27707 416 27709
rect 471 27707 491 27709
rect 540 27707 566 27709
rect 609 27707 640 27709
rect 678 27707 713 27741
rect 747 27707 782 27741
rect 816 27707 851 27741
rect 885 27709 920 27741
rect 954 27709 988 27741
rect 885 27707 908 27709
rect 954 27707 983 27709
rect 1022 27707 1056 27741
rect 1090 27709 1124 27741
rect 1158 27709 1192 27741
rect 1226 27709 1260 27741
rect 1294 27709 1328 27741
rect 1362 27709 1396 27741
rect 1092 27707 1124 27709
rect 1167 27707 1192 27709
rect 1242 27707 1260 27709
rect 1317 27707 1328 27709
rect 1392 27707 1396 27709
rect 1430 27709 1464 27741
rect 1498 27709 1532 27741
rect 1566 27709 1600 27741
rect 1634 27709 1668 27741
rect 1702 27709 1736 27741
rect 1430 27707 1433 27709
rect 1498 27707 1508 27709
rect 1566 27707 1583 27709
rect 1634 27707 1658 27709
rect 1702 27707 1732 27709
rect 1770 27707 1804 27741
rect 1838 27709 1872 27741
rect 1906 27709 1940 27741
rect 1974 27709 2008 27741
rect 2042 27709 2076 27741
rect 2110 27709 2144 27741
rect 2178 27709 2212 27741
rect 1840 27707 1872 27709
rect 1914 27707 1940 27709
rect 1988 27707 2008 27709
rect 2062 27707 2076 27709
rect 2136 27707 2144 27709
rect 2210 27707 2212 27709
rect 2246 27709 2280 27741
rect 2314 27709 2348 27741
rect 2382 27709 2416 27741
rect 2450 27709 2484 27741
rect 2518 27709 2552 27741
rect 2246 27707 2250 27709
rect 2314 27707 2324 27709
rect 2382 27707 2398 27709
rect 2450 27707 2472 27709
rect 2518 27707 2546 27709
rect 2586 27707 2620 27741
rect 2654 27707 2688 27741
rect 2722 27709 2756 27741
rect 2790 27709 2824 27741
rect 2858 27709 2892 27741
rect 2926 27709 2950 27741
rect 2728 27707 2756 27709
rect 2802 27707 2824 27709
rect 2876 27707 2892 27709
rect 196 27675 266 27707
rect 300 27675 341 27707
rect 375 27675 416 27707
rect 450 27675 491 27707
rect 525 27675 566 27707
rect 600 27675 640 27707
rect 674 27675 908 27707
rect 942 27675 983 27707
rect 1017 27675 1058 27707
rect 1092 27675 1133 27707
rect 1167 27675 1208 27707
rect 1242 27675 1283 27707
rect 1317 27675 1358 27707
rect 1392 27675 1433 27707
rect 1467 27675 1508 27707
rect 1542 27675 1583 27707
rect 1617 27675 1658 27707
rect 1692 27675 1732 27707
rect 1766 27675 1806 27707
rect 1840 27675 1880 27707
rect 1914 27675 1954 27707
rect 1988 27675 2028 27707
rect 2062 27675 2102 27707
rect 2136 27675 2176 27707
rect 2210 27675 2250 27707
rect 2284 27675 2324 27707
rect 2358 27675 2398 27707
rect 2432 27675 2472 27707
rect 2506 27675 2546 27707
rect 2580 27675 2620 27707
rect 2654 27675 2694 27707
rect 2728 27675 2768 27707
rect 2802 27675 2842 27707
rect 2876 27675 2916 27707
rect 196 27673 2950 27675
rect 196 27639 264 27673
rect 298 27639 334 27673
rect 368 27639 404 27673
rect 438 27639 474 27673
rect 508 27639 544 27673
rect 578 27639 614 27673
rect 648 27639 684 27673
rect 718 27639 753 27673
rect 787 27639 822 27673
rect 856 27639 891 27673
rect 925 27639 960 27673
rect 994 27639 1029 27673
rect 1063 27639 1098 27673
rect 1132 27639 1167 27673
rect 1201 27639 1236 27673
rect 1270 27639 1305 27673
rect 1339 27639 1374 27673
rect 1408 27639 1443 27673
rect 1477 27639 1512 27673
rect 1546 27639 1581 27673
rect 1615 27639 1650 27673
rect 1684 27639 1719 27673
rect 1753 27639 1788 27673
rect 1822 27639 1857 27673
rect 1891 27639 1926 27673
rect 1960 27639 1995 27673
rect 2029 27639 2064 27673
rect 2098 27639 2133 27673
rect 2167 27639 2202 27673
rect 2236 27639 2271 27673
rect 2305 27639 2340 27673
rect 2374 27639 2409 27673
rect 2443 27639 2478 27673
rect 2512 27639 2547 27673
rect 2581 27639 2616 27673
rect 2650 27639 2685 27673
rect 2719 27639 2754 27673
rect 2788 27639 2823 27673
rect 2857 27639 2892 27673
rect 2926 27639 2950 27673
rect 196 27637 2950 27639
rect 196 27631 300 27637
rect 230 27603 300 27631
rect 334 27605 385 27637
rect 419 27605 470 27637
rect 504 27605 555 27637
rect 589 27605 640 27637
rect 674 27605 908 27637
rect 942 27605 983 27637
rect 1017 27605 1058 27637
rect 1092 27605 1133 27637
rect 366 27603 385 27605
rect 436 27603 470 27605
rect 230 27597 332 27603
rect 196 27586 332 27597
rect 196 27558 228 27586
rect 262 27552 264 27586
rect 298 27571 332 27586
rect 366 27571 402 27603
rect 436 27571 472 27603
rect 506 27571 542 27605
rect 589 27603 612 27605
rect 674 27603 682 27605
rect 576 27571 612 27603
rect 646 27571 682 27603
rect 716 27571 752 27605
rect 786 27571 822 27605
rect 856 27571 891 27605
rect 942 27603 960 27605
rect 1017 27603 1029 27605
rect 1092 27603 1098 27605
rect 925 27571 960 27603
rect 994 27571 1029 27603
rect 1063 27571 1098 27603
rect 1132 27603 1133 27605
rect 1167 27605 1208 27637
rect 1242 27605 1283 27637
rect 1317 27605 1358 27637
rect 1392 27605 1433 27637
rect 1467 27605 1508 27637
rect 1542 27605 1583 27637
rect 1617 27605 1658 27637
rect 1692 27605 1732 27637
rect 1766 27605 1806 27637
rect 1840 27605 1880 27637
rect 1914 27605 1954 27637
rect 1988 27605 2028 27637
rect 2062 27605 2102 27637
rect 2136 27605 2176 27637
rect 2210 27605 2250 27637
rect 2284 27605 2324 27637
rect 2358 27605 2398 27637
rect 2432 27605 2472 27637
rect 2506 27605 2546 27637
rect 2580 27605 2620 27637
rect 2654 27605 2694 27637
rect 2728 27605 2768 27637
rect 2802 27605 2842 27637
rect 2876 27605 2916 27637
rect 1132 27571 1167 27603
rect 1201 27603 1208 27605
rect 1270 27603 1283 27605
rect 1339 27603 1358 27605
rect 1408 27603 1433 27605
rect 1477 27603 1508 27605
rect 1201 27571 1236 27603
rect 1270 27571 1305 27603
rect 1339 27571 1374 27603
rect 1408 27571 1443 27603
rect 1477 27571 1512 27603
rect 1546 27571 1581 27605
rect 1617 27603 1650 27605
rect 1692 27603 1719 27605
rect 1766 27603 1788 27605
rect 1840 27603 1857 27605
rect 1914 27603 1926 27605
rect 1988 27603 1995 27605
rect 2062 27603 2064 27605
rect 1615 27571 1650 27603
rect 1684 27571 1719 27603
rect 1753 27571 1788 27603
rect 1822 27571 1857 27603
rect 1891 27571 1926 27603
rect 1960 27571 1995 27603
rect 2029 27571 2064 27603
rect 2098 27603 2102 27605
rect 2167 27603 2176 27605
rect 2236 27603 2250 27605
rect 2305 27603 2324 27605
rect 2374 27603 2398 27605
rect 2443 27603 2472 27605
rect 2512 27603 2546 27605
rect 2098 27571 2133 27603
rect 2167 27571 2202 27603
rect 2236 27571 2271 27603
rect 2305 27571 2340 27603
rect 2374 27571 2409 27603
rect 2443 27571 2478 27603
rect 2512 27571 2547 27603
rect 2581 27571 2616 27605
rect 2654 27603 2685 27605
rect 2728 27603 2754 27605
rect 2802 27603 2823 27605
rect 2876 27603 2892 27605
rect 2650 27571 2685 27603
rect 2719 27571 2754 27603
rect 2788 27571 2823 27603
rect 2857 27571 2892 27603
rect 2926 27571 2950 27603
rect 298 27552 366 27571
rect 230 27533 366 27552
rect 230 27524 300 27533
rect 196 27507 300 27524
rect 334 27509 366 27533
rect 196 27485 228 27507
rect 262 27499 300 27507
rect 262 27473 264 27499
rect 230 27465 264 27473
rect 298 27475 332 27499
rect 298 27465 366 27475
rect 230 27451 366 27465
rect 196 27428 366 27451
rect 196 27412 228 27428
rect 262 27412 300 27428
rect 334 27412 366 27428
rect 262 27394 264 27412
rect 230 27378 264 27394
rect 298 27394 300 27412
rect 298 27378 332 27394
rect 196 27354 366 27378
rect 196 27330 228 27354
rect 262 27330 300 27354
rect 334 27330 366 27354
rect 262 27320 264 27330
rect 230 27296 264 27320
rect 298 27320 300 27330
rect 298 27296 332 27320
rect 196 27281 366 27296
rect 196 27280 300 27281
rect 196 27261 228 27280
rect 262 27260 300 27280
rect 334 27260 366 27281
rect 262 27246 264 27260
rect 230 27227 264 27246
rect 196 27226 264 27227
rect 298 27247 300 27260
rect 298 27226 332 27247
rect 196 27208 366 27226
rect 196 27206 300 27208
rect 196 27192 228 27206
rect 262 27190 300 27206
rect 334 27190 366 27208
rect 262 27172 264 27190
rect 230 27158 264 27172
rect 196 27156 264 27158
rect 298 27174 300 27190
rect 298 27156 332 27174
rect 196 27135 366 27156
rect 196 27133 300 27135
rect 196 27123 228 27133
rect 262 27120 300 27133
rect 334 27120 366 27135
rect 262 27099 264 27120
rect 230 27089 264 27099
rect 196 27086 264 27089
rect 298 27101 300 27120
rect 298 27086 332 27101
rect 196 27062 366 27086
rect 196 27060 300 27062
rect 196 27054 228 27060
rect 262 27050 300 27060
rect 334 27050 366 27062
rect 262 27026 264 27050
rect 230 27020 264 27026
rect 196 27016 264 27020
rect 298 27028 300 27050
rect 298 27016 332 27028
rect 196 26989 366 27016
rect 196 26987 300 26989
rect 196 26985 228 26987
rect 262 26980 300 26987
rect 334 26980 366 26989
rect 262 26953 264 26980
rect 230 26951 264 26953
rect 196 26946 264 26951
rect 298 26955 300 26980
rect 4396 26975 4412 27009
rect 4446 26975 4480 27009
rect 4514 26975 4530 27009
rect 4808 26975 4824 27009
rect 4858 26975 4892 27009
rect 4926 26975 4942 27009
rect 5220 26975 5236 27009
rect 5270 26975 5304 27009
rect 5338 26975 5354 27009
rect 5632 26975 5648 27009
rect 5682 26975 5716 27009
rect 5750 26975 5766 27009
rect 6044 26975 6060 27009
rect 6094 26975 6128 27009
rect 6162 26975 6178 27009
rect 6456 26975 6472 27009
rect 6506 26975 6540 27009
rect 6574 26975 6590 27009
rect 6868 26975 6884 27009
rect 6918 26975 6952 27009
rect 6986 26975 7002 27009
rect 7280 26975 7296 27009
rect 7330 26975 7364 27009
rect 7398 26975 7414 27009
rect 7692 26975 7708 27009
rect 7742 26975 7776 27009
rect 7810 26975 7826 27009
rect 8104 26975 8120 27009
rect 8154 26975 8188 27009
rect 8222 26975 8238 27009
rect 8516 26975 8532 27009
rect 8566 26975 8600 27009
rect 8634 26975 8650 27009
rect 8928 26975 8944 27009
rect 8978 26975 9012 27009
rect 9046 26975 9062 27009
rect 9340 26975 9356 27009
rect 9390 26975 9424 27009
rect 9458 26975 9474 27009
rect 9752 26975 9768 27009
rect 9802 26975 9836 27009
rect 9870 26975 9886 27009
rect 10164 26975 10180 27009
rect 10214 26975 10248 27009
rect 10282 26975 10298 27009
rect 10576 26975 10592 27009
rect 10626 26975 10660 27009
rect 10694 26975 10710 27009
rect 10988 26975 11004 27009
rect 11038 26975 11072 27009
rect 11106 26975 11122 27009
rect 11400 26975 11416 27009
rect 11450 26975 11484 27009
rect 11518 26975 11534 27009
rect 11812 26975 11828 27009
rect 11862 26975 11896 27009
rect 11930 26975 11946 27009
rect 12224 26975 12240 27009
rect 12274 26975 12308 27009
rect 12342 26975 12358 27009
rect 12636 26975 12652 27009
rect 12686 26975 12720 27009
rect 12754 26975 12770 27009
rect 13048 26975 13064 27009
rect 13098 26975 13132 27009
rect 13166 26975 13182 27009
rect 13460 26975 13476 27009
rect 13510 26975 13544 27009
rect 13578 26975 13594 27009
rect 13872 26975 13888 27009
rect 13922 26975 13956 27009
rect 13990 26975 14006 27009
rect 14284 26975 14300 27009
rect 14334 26975 14368 27009
rect 14402 26975 14418 27009
rect 14592 26998 14712 27009
rect 14626 26964 14664 26998
rect 14698 26975 14712 26998
rect 14746 26975 14780 27009
rect 14814 26975 14830 27009
rect 14698 26964 14830 26975
rect 298 26946 332 26955
rect 196 26916 366 26946
rect 230 26914 300 26916
rect 262 26910 300 26914
rect 334 26910 366 26916
rect 196 26880 228 26882
rect 262 26880 264 26910
rect 196 26876 264 26880
rect 298 26882 300 26910
rect 298 26876 332 26882
rect 196 26847 366 26876
rect 230 26843 366 26847
rect 230 26841 300 26843
rect 196 26807 228 26813
rect 262 26807 264 26841
rect 298 26809 300 26841
rect 334 26840 366 26843
rect 298 26807 332 26809
rect 196 26806 332 26807
rect 196 26778 366 26806
rect 230 26772 366 26778
rect 230 26768 264 26772
rect 196 26734 228 26744
rect 262 26738 264 26768
rect 298 26771 366 26772
rect 298 26770 332 26771
rect 298 26738 300 26770
rect 262 26736 300 26738
rect 334 26736 366 26737
rect 262 26734 366 26736
rect 196 26709 366 26734
rect 230 26703 366 26709
rect 230 26695 264 26703
rect 196 26661 228 26675
rect 262 26669 264 26695
rect 298 26702 366 26703
rect 298 26697 332 26702
rect 298 26669 300 26697
rect 262 26663 300 26669
rect 334 26663 366 26668
rect 262 26661 366 26663
rect 196 26640 366 26661
rect 230 26634 366 26640
rect 230 26622 264 26634
rect 196 26588 228 26606
rect 262 26600 264 26622
rect 298 26633 366 26634
rect 298 26624 332 26633
rect 298 26600 300 26624
rect 262 26590 300 26600
rect 334 26590 366 26599
rect 262 26588 366 26590
rect 196 26571 366 26588
rect 230 26565 366 26571
rect 230 26549 264 26565
rect 196 26515 228 26537
rect 262 26531 264 26549
rect 298 26564 366 26565
rect 298 26551 332 26564
rect 298 26531 300 26551
rect 262 26517 300 26531
rect 334 26517 366 26530
rect 262 26515 366 26517
rect 196 26502 366 26515
rect 230 26496 366 26502
rect 230 26476 264 26496
rect 196 26442 228 26468
rect 262 26462 264 26476
rect 298 26495 366 26496
rect 298 26478 332 26495
rect 298 26462 300 26478
rect 262 26444 300 26462
rect 334 26444 366 26461
rect 262 26442 366 26444
rect 196 26433 366 26442
rect 230 26427 366 26433
rect 230 26403 264 26427
rect 196 26369 228 26399
rect 262 26393 264 26403
rect 298 26426 366 26427
rect 298 26405 332 26426
rect 298 26393 300 26405
rect 262 26371 300 26393
rect 334 26371 366 26392
rect 262 26369 366 26371
rect 196 26364 366 26369
rect 230 26358 366 26364
rect 230 26330 264 26358
rect 196 26296 228 26330
rect 262 26324 264 26330
rect 298 26357 366 26358
rect 298 26332 332 26357
rect 298 26324 300 26332
rect 262 26298 300 26324
rect 334 26298 366 26323
rect 262 26296 366 26298
rect 196 26295 366 26296
rect 230 26289 366 26295
rect 230 26261 264 26289
rect 196 26257 264 26261
rect 196 26226 228 26257
rect 262 26255 264 26257
rect 298 26288 366 26289
rect 298 26259 332 26288
rect 298 26255 300 26259
rect 262 26225 300 26255
rect 334 26225 366 26254
rect 262 26223 366 26225
rect 230 26220 366 26223
rect 230 26192 264 26220
rect 196 26186 264 26192
rect 298 26219 366 26220
rect 298 26186 332 26219
rect 196 26184 300 26186
rect 196 26157 228 26184
rect 262 26152 300 26184
rect 334 26152 366 26185
rect 262 26151 366 26152
rect 262 26150 264 26151
rect 230 26123 264 26150
rect 196 26117 264 26123
rect 298 26150 366 26151
rect 298 26117 332 26150
rect 196 26116 332 26117
rect 196 26113 366 26116
rect 196 26111 300 26113
rect 196 26088 228 26111
rect 262 26082 300 26111
rect 262 26077 264 26082
rect 230 26054 264 26077
rect 196 26048 264 26054
rect 298 26079 300 26082
rect 334 26081 366 26113
rect 298 26048 332 26079
rect 196 26047 332 26048
rect 196 26040 366 26047
rect 196 26038 300 26040
rect 196 26019 228 26038
rect 262 26013 300 26038
rect 262 26004 264 26013
rect 230 25985 264 26004
rect 196 25979 264 25985
rect 298 26006 300 26013
rect 334 26012 366 26040
rect 298 25979 332 26006
rect 196 25978 332 25979
rect 196 25967 366 25978
rect 196 25965 300 25967
rect 196 25950 228 25965
rect 262 25944 300 25965
rect 262 25931 264 25944
rect 230 25916 264 25931
rect 196 25910 264 25916
rect 298 25933 300 25944
rect 334 25943 366 25967
rect 298 25910 332 25933
rect 196 25909 332 25910
rect 196 25894 366 25909
rect 196 25892 300 25894
rect 196 25881 228 25892
rect 262 25875 300 25892
rect 262 25858 264 25875
rect 230 25847 264 25858
rect 196 25841 264 25847
rect 298 25860 300 25875
rect 334 25874 366 25894
rect 298 25841 332 25860
rect 196 25840 332 25841
rect 196 25821 366 25840
rect 196 25819 300 25821
rect 196 25812 228 25819
rect 262 25806 300 25819
rect 262 25785 264 25806
rect 230 25778 264 25785
rect 196 25772 264 25778
rect 298 25787 300 25806
rect 334 25805 366 25821
rect 298 25772 332 25787
rect 196 25771 332 25772
rect 196 25748 366 25771
rect 196 25746 300 25748
rect 196 25743 228 25746
rect 262 25737 300 25746
rect 262 25712 264 25737
rect 230 25709 264 25712
rect 196 25703 264 25709
rect 298 25714 300 25737
rect 334 25736 366 25748
rect 298 25703 332 25714
rect 196 25702 332 25703
rect 196 25675 366 25702
rect 196 25674 300 25675
rect 230 25673 300 25674
rect 262 25668 300 25673
rect 196 25639 228 25640
rect 262 25639 264 25668
rect 196 25634 264 25639
rect 298 25641 300 25668
rect 334 25667 366 25675
rect 298 25634 332 25641
rect 196 25633 332 25634
rect 196 25605 366 25633
rect 230 25602 366 25605
rect 230 25600 300 25602
rect 262 25599 300 25600
rect 196 25566 228 25571
rect 262 25566 264 25599
rect 196 25565 264 25566
rect 298 25568 300 25599
rect 334 25598 366 25602
rect 298 25565 332 25568
rect 196 25564 332 25565
rect 196 25536 366 25564
rect 230 25530 366 25536
rect 230 25527 264 25530
rect 196 25493 228 25502
rect 262 25496 264 25527
rect 298 25529 366 25530
rect 298 25496 300 25529
rect 262 25495 300 25496
rect 262 25493 366 25495
rect 196 25467 366 25493
rect 230 25461 366 25467
rect 230 25454 264 25461
rect 196 25420 228 25433
rect 262 25427 264 25454
rect 298 25460 366 25461
rect 298 25456 332 25460
rect 298 25427 300 25456
rect 262 25422 300 25427
rect 334 25422 366 25426
rect 262 25420 366 25422
rect 196 25398 366 25420
rect 230 25392 366 25398
rect 230 25381 264 25392
rect 196 25347 228 25364
rect 262 25358 264 25381
rect 298 25391 366 25392
rect 298 25383 332 25391
rect 298 25358 300 25383
rect 262 25349 300 25358
rect 2771 25441 2787 25475
rect 2821 25441 2882 25475
rect 2771 25403 2916 25441
rect 2771 25369 2882 25403
rect 334 25349 366 25357
rect 262 25347 366 25349
rect 196 25329 366 25347
rect 230 25323 366 25329
rect 230 25308 264 25323
rect 196 25274 228 25295
rect 262 25289 264 25308
rect 298 25322 366 25323
rect 298 25311 332 25322
rect 298 25289 300 25311
rect 262 25277 300 25289
rect 334 25277 366 25288
rect 262 25274 366 25277
rect 196 25260 366 25274
rect 230 25254 366 25260
rect 230 25235 264 25254
rect 196 25201 228 25226
rect 262 25220 264 25235
rect 298 25253 366 25254
rect 298 25239 332 25253
rect 298 25220 300 25239
rect 262 25205 300 25220
rect 334 25205 366 25219
rect 262 25201 366 25205
rect 196 25191 366 25201
rect 230 25185 366 25191
rect 230 25162 264 25185
rect 196 25128 228 25157
rect 262 25151 264 25162
rect 298 25184 366 25185
rect 298 25167 332 25184
rect 298 25151 300 25167
rect 262 25133 300 25151
rect 334 25133 366 25150
rect 262 25128 366 25133
rect 196 25122 366 25128
rect 230 25116 366 25122
rect 230 25089 264 25116
rect 196 25055 228 25088
rect 262 25082 264 25089
rect 298 25115 366 25116
rect 298 25095 332 25115
rect 298 25082 300 25095
rect 262 25061 300 25082
rect 334 25061 366 25081
rect 262 25055 366 25061
rect 196 25053 366 25055
rect 230 25047 366 25053
rect 230 25019 264 25047
rect 196 25016 264 25019
rect 196 24985 228 25016
rect 262 25013 264 25016
rect 298 25046 366 25047
rect 298 25023 332 25046
rect 298 25013 300 25023
rect 262 24989 300 25013
rect 334 24989 366 25012
rect 262 24982 366 24989
rect 230 24978 366 24982
rect 230 24951 264 24978
rect 196 24944 264 24951
rect 298 24977 366 24978
rect 298 24951 332 24977
rect 298 24944 300 24951
rect 196 24943 300 24944
rect 196 24917 228 24943
rect 262 24917 300 24943
rect 334 24917 366 24943
rect 262 24909 366 24917
rect 230 24883 264 24909
rect 196 24875 264 24883
rect 298 24908 366 24909
rect 298 24879 332 24908
rect 298 24875 300 24879
rect 196 24870 300 24875
rect 196 24849 228 24870
rect 262 24845 300 24870
rect 334 24845 366 24874
rect 262 24840 366 24845
rect 262 24836 264 24840
rect 230 24815 264 24836
rect 196 24806 264 24815
rect 298 24839 366 24840
rect 298 24807 332 24839
rect 298 24806 300 24807
rect 196 24797 300 24806
rect 196 24781 228 24797
rect 262 24773 300 24797
rect 334 24773 366 24805
rect 262 24771 366 24773
rect 262 24763 264 24771
rect 230 24747 264 24763
rect 196 24737 264 24747
rect 298 24770 366 24771
rect 298 24737 332 24770
rect 196 24736 332 24737
rect 196 24735 366 24736
rect 196 24724 300 24735
rect 196 24713 228 24724
rect 262 24702 300 24724
rect 262 24690 264 24702
rect 230 24679 264 24690
rect 196 24668 264 24679
rect 298 24701 300 24702
rect 334 24701 366 24735
rect 298 24668 332 24701
rect 196 24667 332 24668
rect 196 24663 366 24667
rect 196 24651 300 24663
rect 196 24645 228 24651
rect 262 24633 300 24651
rect 262 24617 264 24633
rect 230 24611 264 24617
rect 196 24599 264 24611
rect 298 24629 300 24633
rect 334 24632 366 24663
rect 298 24599 332 24629
rect 196 24598 332 24599
rect 196 24591 366 24598
rect 196 24578 300 24591
rect 196 24577 228 24578
rect 262 24564 300 24578
rect 262 24544 264 24564
rect 230 24543 264 24544
rect 196 24530 264 24543
rect 298 24557 300 24564
rect 334 24563 366 24591
rect 298 24530 332 24557
rect 196 24529 332 24530
rect 196 24519 366 24529
rect 196 24509 300 24519
rect 230 24505 300 24509
rect 262 24495 300 24505
rect 196 24471 228 24475
rect 262 24471 264 24495
rect 196 24461 264 24471
rect 298 24485 300 24495
rect 334 24494 366 24519
rect 298 24461 332 24485
rect 196 24460 332 24461
rect 196 24447 366 24460
rect 196 24441 300 24447
rect 230 24432 300 24441
rect 262 24426 300 24432
rect 196 24398 228 24407
rect 262 24398 264 24426
rect 196 24392 264 24398
rect 298 24413 300 24426
rect 334 24425 366 24447
rect 298 24392 332 24413
rect 196 24391 332 24392
rect 196 24375 366 24391
rect 196 24373 300 24375
rect 230 24359 300 24373
rect 262 24357 300 24359
rect 196 24325 228 24339
rect 262 24325 264 24357
rect 196 24323 264 24325
rect 298 24341 300 24357
rect 334 24356 366 24375
rect 298 24323 332 24341
rect 196 24322 332 24323
rect 196 24305 366 24322
rect 230 24303 366 24305
rect 230 24288 300 24303
rect 230 24286 264 24288
rect 196 24252 228 24271
rect 262 24254 264 24286
rect 298 24269 300 24288
rect 334 24287 366 24303
rect 298 24254 332 24269
rect 262 24253 332 24254
rect 262 24252 366 24253
rect 196 24237 366 24252
rect 230 24231 366 24237
rect 230 24219 300 24231
rect 230 24213 264 24219
rect 196 24179 228 24203
rect 262 24185 264 24213
rect 298 24197 300 24219
rect 334 24218 366 24231
rect 298 24185 332 24197
rect 262 24184 332 24185
rect 262 24179 366 24184
rect 196 24169 366 24179
rect 230 24159 366 24169
rect 230 24150 300 24159
rect 230 24140 264 24150
rect 196 24106 228 24135
rect 262 24116 264 24140
rect 298 24125 300 24150
rect 334 24149 366 24159
rect 298 24116 332 24125
rect 262 24115 332 24116
rect 262 24106 366 24115
rect 196 24101 366 24106
rect 230 24087 366 24101
rect 230 24081 300 24087
rect 230 24067 264 24081
rect 196 24033 228 24067
rect 262 24047 264 24067
rect 298 24053 300 24081
rect 334 24080 366 24087
rect 298 24047 332 24053
rect 262 24046 332 24047
rect 262 24033 366 24046
rect 230 24015 366 24033
rect 230 24012 300 24015
rect 230 23999 264 24012
rect 196 23994 264 23999
rect 196 23965 228 23994
rect 262 23978 264 23994
rect 298 23981 300 24012
rect 334 24011 366 24015
rect 298 23978 332 23981
rect 262 23977 332 23978
rect 262 23960 366 23977
rect 230 23943 366 23960
rect 230 23931 264 23943
rect 196 23921 264 23931
rect 196 23897 228 23921
rect 262 23909 264 23921
rect 298 23909 300 23943
rect 334 23942 366 23943
rect 262 23908 332 23909
rect 262 23887 366 23908
rect 230 23874 366 23887
rect 230 23863 264 23874
rect 196 23848 264 23863
rect 196 23829 228 23848
rect 262 23840 264 23848
rect 298 23873 366 23874
rect 298 23871 332 23873
rect 298 23840 300 23871
rect 262 23837 300 23840
rect 334 23837 366 23839
rect 262 23814 366 23837
rect 230 23805 366 23814
rect 230 23795 264 23805
rect 196 23775 264 23795
rect 196 23761 228 23775
rect 262 23771 264 23775
rect 298 23804 366 23805
rect 298 23799 332 23804
rect 298 23771 300 23799
rect 262 23765 300 23771
rect 334 23765 366 23770
rect 262 23741 366 23765
rect 230 23736 366 23741
rect 230 23727 264 23736
rect 196 23702 264 23727
rect 298 23735 366 23736
rect 298 23727 332 23735
rect 298 23702 300 23727
rect 196 23693 228 23702
rect 262 23693 300 23702
rect 334 23693 366 23701
rect 262 23668 366 23693
rect 230 23667 366 23668
rect 230 23659 264 23667
rect 196 23633 264 23659
rect 298 23666 366 23667
rect 298 23655 332 23666
rect 298 23633 300 23655
rect 196 23629 300 23633
rect 196 23625 228 23629
rect 262 23621 300 23629
rect 334 23621 366 23632
rect 262 23598 366 23621
rect 262 23595 264 23598
rect 230 23591 264 23595
rect 196 23564 264 23591
rect 298 23597 366 23598
rect 298 23583 332 23597
rect 298 23564 300 23583
rect 196 23557 300 23564
rect 230 23556 300 23557
rect 262 23549 300 23556
rect 334 23549 366 23563
rect 262 23529 366 23549
rect 196 23522 228 23523
rect 262 23522 264 23529
rect 196 23495 264 23522
rect 298 23528 366 23529
rect 298 23511 332 23528
rect 298 23495 300 23511
rect 196 23489 300 23495
rect 230 23483 300 23489
rect 262 23477 300 23483
rect 334 23477 366 23494
rect 262 23460 366 23477
rect 196 23449 228 23455
rect 262 23449 264 23460
rect 196 23426 264 23449
rect 298 23459 366 23460
rect 298 23439 332 23459
rect 298 23426 300 23439
rect 196 23421 300 23426
rect 230 23410 300 23421
rect 262 23405 300 23410
rect 334 23405 366 23425
rect 262 23391 366 23405
rect 196 23376 228 23387
rect 262 23376 264 23391
rect 196 23357 264 23376
rect 298 23390 366 23391
rect 298 23367 332 23390
rect 298 23357 300 23367
rect 196 23353 300 23357
rect 230 23337 300 23353
rect 262 23333 300 23337
rect 334 23333 366 23356
rect 518 24942 552 25050
rect 586 25016 623 25050
rect 657 25016 694 25050
rect 728 25016 764 25050
rect 798 25016 834 25050
rect 868 25016 892 25050
rect 518 24871 552 24908
rect 518 24800 552 24837
rect 518 24729 552 24766
rect 518 24658 552 24695
rect 518 24587 552 24624
rect 518 24516 552 24553
rect 518 24445 552 24482
rect 518 24374 552 24411
rect 518 24303 552 24340
rect 518 24221 552 24269
rect 735 24203 778 24237
rect 812 24203 855 24237
rect 889 24203 932 24237
rect 966 24203 1009 24237
rect 1043 24203 1086 24237
rect 1120 24203 1162 24237
rect 1196 24203 1238 24237
rect 1272 24203 1314 24237
rect 1348 24203 1390 24237
rect 1424 24203 1466 24237
rect 1500 24203 1542 24237
rect 1576 24203 1618 24237
rect 1758 24221 1792 24245
rect 518 24148 552 24187
rect 518 24075 552 24114
rect 518 24001 552 24041
rect 518 23927 552 23967
rect 590 24182 624 24192
rect 590 24176 615 24182
rect 624 24142 649 24148
rect 590 24110 649 24142
rect 590 24108 615 24110
rect 1758 24147 1792 24187
rect 624 24074 649 24076
rect 590 24040 649 24074
rect 735 24047 778 24081
rect 812 24047 855 24081
rect 889 24047 932 24081
rect 966 24047 1009 24081
rect 1043 24047 1086 24081
rect 1120 24047 1162 24081
rect 1196 24047 1238 24081
rect 1272 24047 1314 24081
rect 1348 24047 1390 24081
rect 1424 24047 1466 24081
rect 1500 24047 1542 24081
rect 1576 24047 1618 24081
rect 1758 24073 1792 24113
rect 624 24038 649 24040
rect 590 24004 615 24006
rect 590 23972 649 24004
rect 624 23966 649 23972
rect 590 23932 615 23938
rect 1758 23999 1792 24039
rect 590 23922 624 23932
rect 1758 23925 1792 23965
rect 518 23853 552 23893
rect 735 23891 778 23925
rect 812 23891 855 23925
rect 889 23891 932 23925
rect 966 23891 1009 23925
rect 1043 23891 1086 23925
rect 1120 23891 1162 23925
rect 1196 23891 1238 23925
rect 1272 23891 1314 23925
rect 1348 23891 1390 23925
rect 1424 23891 1466 23925
rect 1500 23891 1542 23925
rect 1576 23891 1618 23925
rect 518 23779 552 23819
rect 1758 23852 1792 23891
rect 518 23705 552 23745
rect 518 23631 552 23671
rect 518 23557 552 23597
rect 518 23483 552 23523
rect 590 23779 624 23784
rect 735 23781 778 23815
rect 812 23781 855 23815
rect 889 23781 932 23815
rect 966 23781 1009 23815
rect 1043 23781 1086 23815
rect 1120 23781 1162 23815
rect 1196 23781 1238 23815
rect 1272 23781 1314 23815
rect 1348 23781 1390 23815
rect 1424 23781 1466 23815
rect 1500 23781 1542 23815
rect 1576 23781 1618 23815
rect 1758 23779 1792 23818
rect 14696 23779 14830 26964
rect 590 23768 615 23779
rect 624 23734 649 23745
rect 590 23707 649 23734
rect 590 23700 615 23707
rect 624 23666 649 23673
rect 590 23635 649 23666
rect 1758 23706 1792 23745
rect 590 23632 615 23635
rect 735 23625 778 23659
rect 812 23625 855 23659
rect 889 23625 932 23659
rect 966 23625 1009 23659
rect 1043 23625 1086 23659
rect 1120 23625 1162 23659
rect 1196 23625 1238 23659
rect 1272 23625 1314 23659
rect 1348 23625 1390 23659
rect 1424 23625 1466 23659
rect 1500 23625 1542 23659
rect 1576 23625 1618 23659
rect 1758 23633 1792 23672
rect 4396 23745 4410 23779
rect 4446 23745 4480 23779
rect 4516 23745 4530 23779
rect 4808 23745 4822 23779
rect 4858 23745 4892 23779
rect 4928 23745 4942 23779
rect 5220 23745 5234 23779
rect 5270 23745 5304 23779
rect 5340 23745 5354 23779
rect 5632 23745 5646 23779
rect 5682 23745 5716 23779
rect 5752 23745 5766 23779
rect 6044 23745 6058 23779
rect 6094 23745 6128 23779
rect 6164 23745 6178 23779
rect 6456 23745 6470 23779
rect 6506 23745 6540 23779
rect 6576 23745 6590 23779
rect 6868 23745 6882 23779
rect 6918 23745 6952 23779
rect 6988 23745 7002 23779
rect 7280 23745 7294 23779
rect 7330 23745 7364 23779
rect 7400 23745 7414 23779
rect 7692 23745 7706 23779
rect 7742 23745 7776 23779
rect 7812 23745 7826 23779
rect 8104 23745 8118 23779
rect 8154 23745 8188 23779
rect 8224 23745 8238 23779
rect 8516 23745 8530 23779
rect 8566 23745 8600 23779
rect 8636 23745 8650 23779
rect 8928 23745 8942 23779
rect 8978 23745 9012 23779
rect 9048 23745 9062 23779
rect 9340 23745 9354 23779
rect 9390 23745 9424 23779
rect 9460 23745 9474 23779
rect 9752 23745 9766 23779
rect 9802 23745 9836 23779
rect 9872 23745 9886 23779
rect 10164 23745 10178 23779
rect 10214 23745 10248 23779
rect 10284 23745 10298 23779
rect 10576 23745 10590 23779
rect 10626 23745 10660 23779
rect 10696 23745 10710 23779
rect 10988 23745 11002 23779
rect 11038 23745 11072 23779
rect 11108 23745 11122 23779
rect 11278 23745 11316 23779
rect 11400 23745 11414 23779
rect 11450 23745 11484 23779
rect 11520 23745 11534 23779
rect 11654 23745 11692 23779
rect 11812 23745 11826 23779
rect 11862 23745 11896 23779
rect 11932 23745 11946 23779
rect 12066 23745 12104 23779
rect 12224 23745 12238 23779
rect 12274 23745 12308 23779
rect 12344 23745 12358 23779
rect 12478 23745 12516 23779
rect 12636 23745 12650 23779
rect 12686 23745 12720 23779
rect 12756 23745 12770 23779
rect 12890 23745 12928 23779
rect 13048 23745 13062 23779
rect 13098 23745 13132 23779
rect 13168 23745 13182 23779
rect 13302 23745 13340 23779
rect 13460 23745 13474 23779
rect 13510 23745 13544 23779
rect 13580 23745 13594 23779
rect 13714 23745 13752 23779
rect 13872 23745 13886 23779
rect 13922 23745 13956 23779
rect 13992 23745 14006 23779
rect 14126 23745 14164 23779
rect 14284 23745 14298 23779
rect 14334 23745 14368 23779
rect 14404 23745 14418 23779
rect 14502 23745 14540 23779
rect 14690 23745 14712 23779
rect 14762 23745 14780 23779
rect 14814 23745 14830 23779
rect 15108 23745 15124 23779
rect 15158 23745 15192 23779
rect 15230 23745 15242 23779
rect 15520 23745 15536 23779
rect 15570 23745 15604 23779
rect 15642 23745 15654 23779
rect 15932 23745 15948 23779
rect 15982 23745 16016 23779
rect 16054 23745 16066 23779
rect 16344 23745 16360 23779
rect 16394 23745 16428 23779
rect 16466 23745 16478 23779
rect 16756 23745 16772 23779
rect 16806 23745 16840 23779
rect 16878 23745 16890 23779
rect 17149 23745 17184 23779
rect 17221 23745 17252 23779
rect 17286 23745 17302 23779
rect 4396 23699 4528 23745
rect 4396 23665 4410 23699
rect 4444 23665 4482 23699
rect 4516 23665 4528 23699
rect 624 23598 649 23601
rect 590 23564 649 23598
rect 624 23563 649 23564
rect 590 23529 615 23530
rect 1758 23560 1792 23599
rect 11002 23622 11108 23745
rect 11244 23699 11350 23745
rect 11278 23665 11316 23699
rect 11036 23588 11074 23622
rect 11620 23622 11726 23745
rect 12032 23699 12138 23745
rect 12066 23665 12104 23699
rect 11654 23588 11692 23622
rect 12444 23622 12550 23745
rect 12856 23699 12962 23745
rect 12890 23665 12928 23699
rect 12478 23588 12516 23622
rect 13268 23622 13374 23745
rect 13680 23699 13786 23745
rect 13714 23665 13752 23699
rect 13302 23588 13340 23622
rect 14092 23622 14198 23745
rect 14468 23699 14574 23745
rect 14502 23665 14540 23699
rect 14126 23588 14164 23622
rect 590 23514 624 23529
rect 735 23469 778 23503
rect 812 23469 855 23503
rect 889 23469 932 23503
rect 966 23469 1009 23503
rect 1043 23469 1086 23503
rect 1120 23469 1162 23503
rect 1196 23469 1238 23503
rect 1272 23469 1314 23503
rect 1348 23469 1390 23503
rect 1424 23469 1466 23503
rect 1500 23469 1542 23503
rect 1576 23469 1618 23503
rect 1758 23487 1792 23526
rect 518 23409 552 23449
rect 518 23341 620 23375
rect 654 23341 689 23375
rect 723 23341 758 23375
rect 792 23341 827 23375
rect 861 23341 896 23375
rect 930 23341 965 23375
rect 999 23341 1034 23375
rect 1068 23341 1103 23375
rect 1137 23341 1172 23375
rect 1206 23341 1241 23375
rect 1275 23341 1310 23375
rect 1344 23341 1379 23375
rect 1413 23341 1448 23375
rect 1482 23341 1517 23375
rect 1551 23341 1586 23375
rect 1620 23341 1655 23375
rect 1689 23341 1724 23375
rect 1758 23341 1792 23453
rect 2651 23425 2689 23459
rect 2723 23425 2837 23459
rect 262 23322 366 23333
rect 196 23303 228 23319
rect 262 23303 264 23322
rect 196 23288 264 23303
rect 298 23321 366 23322
rect 298 23295 332 23321
rect 298 23288 300 23295
rect 196 23285 300 23288
rect 230 23264 300 23285
rect 262 23261 300 23264
rect 334 23261 366 23287
rect 262 23253 366 23261
rect 196 23230 228 23251
rect 262 23230 264 23253
rect 196 23219 264 23230
rect 298 23252 366 23253
rect 298 23223 332 23252
rect 2771 23265 2837 23425
rect 2771 23231 2787 23265
rect 2821 23231 2837 23265
rect 298 23219 300 23223
rect 196 23217 300 23219
rect 230 23191 300 23217
rect 262 23189 300 23191
rect 334 23189 366 23218
rect 262 23184 366 23189
rect 196 23157 228 23183
rect 262 23157 264 23184
rect 196 23150 264 23157
rect 298 23183 366 23184
rect 298 23151 332 23183
rect 366 23151 402 23183
rect 436 23151 472 23183
rect 506 23151 542 23183
rect 576 23151 612 23183
rect 646 23151 682 23183
rect 716 23151 752 23183
rect 786 23151 822 23183
rect 856 23151 891 23183
rect 925 23151 960 23183
rect 298 23150 300 23151
rect 196 23149 300 23150
rect 366 23149 373 23151
rect 436 23149 446 23151
rect 506 23149 519 23151
rect 576 23149 592 23151
rect 646 23149 665 23151
rect 716 23149 738 23151
rect 786 23149 811 23151
rect 856 23149 884 23151
rect 925 23149 957 23151
rect 994 23149 1029 23183
rect 1063 23151 1098 23183
rect 1132 23151 1167 23183
rect 1201 23151 1236 23183
rect 1270 23151 1305 23183
rect 1339 23151 1374 23183
rect 1408 23151 1443 23183
rect 1477 23151 1512 23183
rect 1546 23151 1581 23183
rect 1615 23151 1650 23183
rect 1064 23149 1098 23151
rect 1137 23149 1167 23151
rect 1210 23149 1236 23151
rect 1283 23149 1305 23151
rect 1356 23149 1374 23151
rect 1429 23149 1443 23151
rect 1502 23149 1512 23151
rect 1575 23149 1581 23151
rect 1648 23149 1650 23151
rect 1684 23151 1719 23183
rect 1753 23151 1788 23183
rect 1822 23151 1857 23183
rect 1891 23151 1926 23183
rect 1960 23151 1995 23183
rect 2029 23151 2064 23183
rect 2098 23151 2133 23183
rect 2167 23151 2202 23183
rect 2236 23151 2271 23183
rect 1684 23149 1687 23151
rect 1753 23149 1760 23151
rect 1822 23149 1833 23151
rect 1891 23149 1906 23151
rect 1960 23149 1979 23151
rect 2029 23149 2052 23151
rect 2098 23149 2124 23151
rect 2167 23149 2196 23151
rect 2236 23149 2268 23151
rect 2305 23149 2340 23183
rect 2374 23149 2409 23183
rect 2443 23151 2478 23183
rect 2512 23151 2547 23183
rect 2581 23151 2616 23183
rect 2650 23151 2685 23183
rect 2719 23151 2754 23183
rect 2788 23151 2823 23183
rect 2857 23151 2892 23183
rect 2926 23151 2950 23183
rect 2446 23149 2478 23151
rect 2518 23149 2547 23151
rect 2590 23149 2616 23151
rect 2662 23149 2685 23151
rect 2734 23149 2754 23151
rect 2806 23149 2823 23151
rect 2878 23149 2892 23151
rect 230 23117 300 23149
rect 334 23117 373 23149
rect 407 23117 446 23149
rect 480 23117 519 23149
rect 553 23117 592 23149
rect 626 23117 665 23149
rect 699 23117 738 23149
rect 772 23117 811 23149
rect 845 23117 884 23149
rect 918 23117 957 23149
rect 991 23117 1030 23149
rect 1064 23117 1103 23149
rect 1137 23117 1176 23149
rect 1210 23117 1249 23149
rect 1283 23117 1322 23149
rect 1356 23117 1395 23149
rect 1429 23117 1468 23149
rect 1502 23117 1541 23149
rect 1575 23117 1614 23149
rect 1648 23117 1687 23149
rect 1721 23117 1760 23149
rect 1794 23117 1833 23149
rect 1867 23117 1906 23149
rect 1940 23117 1979 23149
rect 2013 23117 2052 23149
rect 2086 23117 2124 23149
rect 2158 23117 2196 23149
rect 2230 23117 2268 23149
rect 2302 23117 2340 23149
rect 2374 23117 2412 23149
rect 2446 23117 2484 23149
rect 2518 23117 2556 23149
rect 2590 23117 2628 23149
rect 2662 23117 2700 23149
rect 2734 23117 2772 23149
rect 2806 23117 2844 23149
rect 2878 23117 2916 23149
rect 230 23115 2950 23117
rect 196 23081 264 23115
rect 298 23081 334 23115
rect 368 23081 404 23115
rect 438 23081 474 23115
rect 508 23081 544 23115
rect 578 23081 614 23115
rect 648 23081 684 23115
rect 718 23081 753 23115
rect 787 23081 822 23115
rect 856 23081 891 23115
rect 925 23081 960 23115
rect 994 23081 1029 23115
rect 1063 23081 1098 23115
rect 1132 23081 1167 23115
rect 1201 23081 1236 23115
rect 1270 23081 1305 23115
rect 1339 23081 1374 23115
rect 1408 23081 1443 23115
rect 1477 23081 1512 23115
rect 1546 23081 1581 23115
rect 1615 23081 1650 23115
rect 1684 23081 1719 23115
rect 1753 23081 1788 23115
rect 1822 23081 1857 23115
rect 1891 23081 1926 23115
rect 1960 23081 1995 23115
rect 2029 23081 2064 23115
rect 2098 23081 2133 23115
rect 2167 23081 2202 23115
rect 2236 23081 2271 23115
rect 2305 23081 2340 23115
rect 2374 23081 2409 23115
rect 2443 23081 2478 23115
rect 2512 23081 2547 23115
rect 2581 23081 2616 23115
rect 2650 23081 2685 23115
rect 2719 23081 2754 23115
rect 2788 23081 2823 23115
rect 2857 23081 2892 23115
rect 2926 23081 2950 23115
rect 196 23079 2950 23081
rect 196 23047 266 23079
rect 300 23047 340 23079
rect 374 23047 414 23079
rect 448 23047 488 23079
rect 522 23047 562 23079
rect 596 23047 636 23079
rect 670 23047 710 23079
rect 744 23047 784 23079
rect 818 23047 858 23079
rect 892 23047 932 23079
rect 966 23047 1006 23079
rect 1040 23047 1080 23079
rect 1114 23047 1154 23079
rect 1188 23047 1228 23079
rect 1262 23047 1302 23079
rect 1336 23047 1376 23079
rect 1410 23047 1450 23079
rect 1484 23047 1524 23079
rect 1558 23047 1598 23079
rect 1632 23047 1672 23079
rect 1706 23047 1746 23079
rect 1780 23047 1820 23079
rect 1854 23047 1894 23079
rect 1928 23047 1967 23079
rect 2001 23047 2040 23079
rect 2074 23047 2113 23079
rect 2147 23047 2186 23079
rect 2220 23047 2259 23079
rect 2293 23047 2332 23079
rect 2366 23047 2405 23079
rect 2439 23047 2478 23079
rect 2512 23047 2551 23079
rect 2585 23047 2624 23079
rect 2658 23047 2697 23079
rect 2731 23047 2770 23079
rect 2804 23047 2843 23079
rect 2877 23047 2916 23079
rect 196 23013 230 23047
rect 264 23045 266 23047
rect 333 23045 340 23047
rect 402 23045 414 23047
rect 471 23045 488 23047
rect 540 23045 562 23047
rect 609 23045 636 23047
rect 678 23045 710 23047
rect 264 23013 299 23045
rect 333 23013 368 23045
rect 402 23013 437 23045
rect 471 23013 506 23045
rect 540 23013 575 23045
rect 609 23013 644 23045
rect 678 23013 713 23045
rect 747 23013 782 23047
rect 818 23045 851 23047
rect 892 23045 920 23047
rect 966 23045 988 23047
rect 1040 23045 1056 23047
rect 1114 23045 1124 23047
rect 1188 23045 1192 23047
rect 816 23013 851 23045
rect 885 23013 920 23045
rect 954 23013 988 23045
rect 1022 23013 1056 23045
rect 1090 23013 1124 23045
rect 1158 23013 1192 23045
rect 1226 23045 1228 23047
rect 1294 23045 1302 23047
rect 1362 23045 1376 23047
rect 1430 23045 1450 23047
rect 1498 23045 1524 23047
rect 1566 23045 1598 23047
rect 1226 23013 1260 23045
rect 1294 23013 1328 23045
rect 1362 23013 1396 23045
rect 1430 23013 1464 23045
rect 1498 23013 1532 23045
rect 1566 23013 1600 23045
rect 1634 23013 1668 23047
rect 1706 23045 1736 23047
rect 1780 23045 1804 23047
rect 1854 23045 1872 23047
rect 1928 23045 1940 23047
rect 2001 23045 2008 23047
rect 2074 23045 2076 23047
rect 1702 23013 1736 23045
rect 1770 23013 1804 23045
rect 1838 23013 1872 23045
rect 1906 23013 1940 23045
rect 1974 23013 2008 23045
rect 2042 23013 2076 23045
rect 2110 23045 2113 23047
rect 2178 23045 2186 23047
rect 2246 23045 2259 23047
rect 2314 23045 2332 23047
rect 2382 23045 2405 23047
rect 2450 23045 2478 23047
rect 2518 23045 2551 23047
rect 2110 23013 2144 23045
rect 2178 23013 2212 23045
rect 2246 23013 2280 23045
rect 2314 23013 2348 23045
rect 2382 23013 2416 23045
rect 2450 23013 2484 23045
rect 2518 23013 2552 23045
rect 2586 23013 2620 23047
rect 2658 23045 2688 23047
rect 2731 23045 2756 23047
rect 2804 23045 2824 23047
rect 2877 23045 2892 23047
rect 2654 23013 2688 23045
rect 2722 23013 2756 23045
rect 2790 23013 2824 23045
rect 2858 23013 2892 23045
rect 2926 23013 2950 23045
rect -14 22727 21 22759
rect 55 22727 90 22759
rect 124 22727 159 22759
rect 193 22727 228 22759
rect 262 22727 297 22759
rect -14 22725 -5 22727
rect 55 22725 70 22727
rect 124 22725 144 22727
rect 193 22725 218 22727
rect 262 22725 292 22727
rect 331 22725 366 22759
rect 400 22725 435 22759
rect 469 22727 504 22759
rect 538 22727 573 22759
rect 607 22727 642 22759
rect 676 22727 711 22759
rect 745 22727 780 22759
rect 2174 22727 2208 22759
rect 474 22725 504 22727
rect 548 22725 573 22727
rect 622 22725 642 22727
rect 696 22725 711 22727
rect -82 22693 -80 22725
rect -46 22693 -5 22725
rect 29 22693 70 22725
rect 104 22693 144 22725
rect 178 22693 218 22725
rect 252 22693 292 22725
rect 326 22693 366 22725
rect 400 22693 440 22725
rect 474 22693 514 22725
rect 548 22693 588 22725
rect 622 22693 662 22725
rect 696 22693 736 22725
rect 770 22693 780 22727
rect 2176 22693 2208 22727
rect -82 22691 780 22693
rect -184 22657 -116 22691
rect -82 22657 -47 22691
rect -13 22657 22 22691
rect 56 22657 91 22691
rect 125 22657 160 22691
rect 194 22657 229 22691
rect 263 22657 298 22691
rect 332 22657 367 22691
rect 401 22657 436 22691
rect 470 22657 505 22691
rect 539 22657 574 22691
rect 608 22657 643 22691
rect 677 22657 712 22691
rect 746 22657 780 22691
rect 2174 22657 2208 22693
rect -184 22655 2208 22657
rect -184 22623 -114 22655
rect -184 22589 -150 22623
rect -116 22621 -114 22623
rect -80 22623 -41 22655
rect -7 22623 32 22655
rect 66 22623 105 22655
rect 139 22623 178 22655
rect 212 22623 251 22655
rect 285 22623 324 22655
rect 358 22623 397 22655
rect 431 22623 470 22655
rect 504 22623 543 22655
rect 577 22623 616 22655
rect 650 22623 689 22655
rect 723 22623 762 22655
rect 796 22623 835 22655
rect 869 22623 908 22655
rect 942 22623 981 22655
rect 1015 22623 1054 22655
rect 1088 22623 1127 22655
rect 1161 22623 1200 22655
rect 1234 22623 1273 22655
rect 1307 22623 1346 22655
rect -116 22589 -80 22621
rect -46 22621 -41 22623
rect 24 22621 32 22623
rect 94 22621 105 22623
rect 164 22621 178 22623
rect 234 22621 251 22623
rect 304 22621 324 22623
rect 374 22621 397 22623
rect 444 22621 470 22623
rect 514 22621 543 22623
rect 584 22621 616 22623
rect 654 22621 689 22623
rect -46 22589 -10 22621
rect 24 22589 60 22621
rect 94 22589 130 22621
rect 164 22589 200 22621
rect 234 22589 270 22621
rect 304 22589 340 22621
rect 374 22589 410 22621
rect 444 22589 480 22621
rect 514 22589 550 22621
rect 584 22589 620 22621
rect 654 22589 690 22621
rect 724 22589 760 22623
rect 796 22621 829 22623
rect 869 22621 898 22623
rect 942 22621 967 22623
rect 1015 22621 1036 22623
rect 1088 22621 1105 22623
rect 1161 22621 1174 22623
rect 1234 22621 1243 22623
rect 1307 22621 1312 22623
rect 794 22589 829 22621
rect 863 22589 898 22621
rect 932 22589 967 22621
rect 1001 22589 1036 22621
rect 1070 22589 1105 22621
rect 1139 22589 1174 22621
rect 1208 22589 1243 22621
rect 1277 22589 1312 22621
rect 1380 22623 1419 22655
rect 1453 22623 1492 22655
rect 1526 22623 1565 22655
rect 1599 22623 1638 22655
rect 1672 22623 1710 22655
rect 1744 22623 1782 22655
rect 1816 22623 1854 22655
rect 1888 22623 1926 22655
rect 1960 22623 1998 22655
rect 2032 22623 2070 22655
rect 2104 22623 2142 22655
rect 1380 22621 1381 22623
rect 1346 22589 1381 22621
rect 1415 22621 1419 22623
rect 1484 22621 1492 22623
rect 1553 22621 1565 22623
rect 1622 22621 1638 22623
rect 1691 22621 1710 22623
rect 1760 22621 1782 22623
rect 1829 22621 1854 22623
rect 1898 22621 1926 22623
rect 1967 22621 1998 22623
rect 2036 22621 2070 22623
rect 1415 22589 1450 22621
rect 1484 22589 1519 22621
rect 1553 22589 1588 22621
rect 1622 22589 1657 22621
rect 1691 22589 1726 22621
rect 1760 22589 1795 22621
rect 1829 22589 1864 22621
rect 1898 22589 1933 22621
rect 1967 22589 2002 22621
rect 2036 22589 2071 22621
rect 2105 22589 2140 22623
rect 2176 22621 2208 22655
rect 2174 22589 2208 22621
rect -2199 18309 -2089 18343
rect -2055 18309 -2016 18343
rect -1982 18309 -1943 18343
rect -1909 18309 -1870 18343
rect -1836 18309 -1797 18343
rect -1763 18309 -1724 18343
rect -1690 18309 -1651 18343
rect -1617 18309 -1578 18343
rect -1544 18309 -1505 18343
rect -1471 18309 -1432 18343
rect -1398 18309 -1359 18343
rect -1325 18309 -1286 18343
rect -1252 18309 -1213 18343
rect -1179 18309 -1140 18343
rect -1106 18309 -1067 18343
rect -1033 18309 -994 18343
rect -960 18309 -921 18343
rect -887 18309 -848 18343
rect -814 18309 -775 18343
rect -741 18309 -702 18343
rect -668 18309 -629 18343
rect -595 18309 -556 18343
rect -522 18309 -483 18343
rect -449 18309 -410 18343
rect -376 18309 -337 18343
rect -303 18309 -264 18343
rect -230 18309 -191 18343
rect -157 18309 -118 18343
rect -84 18309 -45 18343
rect -11 18309 28 18343
rect 62 18309 101 18343
rect 135 18309 174 18343
rect 208 18309 247 18343
rect 281 18309 320 18343
rect 354 18309 393 18343
rect 427 18309 466 18343
rect 500 18309 539 18343
rect 573 18309 612 18343
rect 646 18309 685 18343
rect 719 18309 758 18343
rect 792 18309 831 18343
rect 865 18309 904 18343
rect 938 18309 977 18343
rect 1011 18309 1050 18343
rect 1084 18309 1123 18343
rect 1157 18309 1196 18343
rect 1230 18309 1269 18343
rect 1303 18309 1342 18343
rect 1376 18309 1415 18343
rect 1449 18309 1488 18343
rect 1522 18309 1561 18343
rect 1595 18309 1634 18343
rect 1668 18309 1707 18343
rect -2199 18305 1741 18309
rect -2165 18271 1741 18305
rect -2199 18237 -2127 18271
rect -2093 18237 -2055 18271
rect -2021 18237 -1983 18271
rect -1949 18237 -1911 18271
rect -1877 18237 -1839 18271
rect -1805 18237 -1767 18271
rect -1733 18237 -1695 18271
rect -1661 18237 -1623 18271
rect -1589 18237 -1551 18271
rect -1517 18237 -1479 18271
rect -1445 18237 -1407 18271
rect -1373 18237 -1335 18271
rect -1301 18237 -1263 18271
rect -1229 18237 -1191 18271
rect -1157 18237 -1119 18271
rect -1085 18237 -1047 18271
rect -1013 18237 -975 18271
rect -941 18237 -903 18271
rect -869 18237 -831 18271
rect -797 18237 -759 18271
rect -725 18237 -687 18271
rect -653 18237 -615 18271
rect -581 18237 -543 18271
rect -509 18237 -471 18271
rect -437 18237 -399 18271
rect -365 18237 -327 18271
rect -293 18237 -255 18271
rect -221 18237 -183 18271
rect -149 18237 -111 18271
rect -77 18237 -39 18271
rect -5 18237 33 18271
rect 67 18237 105 18271
rect 139 18237 177 18271
rect 211 18237 249 18271
rect 283 18237 321 18271
rect 355 18237 393 18271
rect 427 18237 466 18271
rect 500 18237 539 18271
rect 573 18237 612 18271
rect 646 18237 685 18271
rect 719 18237 758 18271
rect 792 18237 831 18271
rect 865 18237 904 18271
rect 938 18237 977 18271
rect 1011 18237 1050 18271
rect 1084 18237 1123 18271
rect 1157 18237 1196 18271
rect 1230 18237 1269 18271
rect 1303 18237 1342 18271
rect 1376 18237 1415 18271
rect 1449 18237 1488 18271
rect 1522 18237 1561 18271
rect 1595 18237 1634 18271
rect 1668 18237 1707 18271
rect -2199 18233 -2093 18237
rect -2165 18199 -2093 18233
rect -2199 18180 -2093 18199
rect -2199 18161 -2127 18180
rect -2165 18146 -2127 18161
rect -2165 18127 -2093 18146
rect -2199 18089 -2093 18127
rect -2165 18055 -2127 18089
rect 172 5219 206 5253
rect 240 5219 278 5253
rect 312 5219 350 5253
rect 384 5219 422 5253
rect 456 5219 494 5253
rect 528 5219 566 5253
rect 600 5219 638 5253
rect 672 5219 710 5253
rect 744 5219 782 5253
rect 816 5219 854 5253
rect 888 5219 925 5253
rect 959 5219 996 5253
rect 1030 5219 1067 5253
rect 1101 5219 1138 5253
rect 1172 5219 1209 5253
rect 1243 5219 1280 5253
rect 1314 5219 1422 5253
rect 172 5185 1388 5219
rect 172 5151 240 5185
rect 274 5151 312 5185
rect 346 5151 384 5185
rect 418 5151 456 5185
rect 490 5151 528 5185
rect 562 5151 600 5185
rect 634 5151 672 5185
rect 706 5151 744 5185
rect 778 5151 816 5185
rect 850 5151 888 5185
rect 922 5151 960 5185
rect 994 5151 1032 5185
rect 1066 5151 1104 5185
rect 1138 5151 1176 5185
rect 1210 5151 1248 5185
rect 1282 5151 1320 5185
rect 1354 5151 1422 5185
rect 172 5149 1422 5151
rect 206 5117 1388 5149
rect 206 5115 308 5117
rect 172 5113 308 5115
rect 172 5080 240 5113
rect 206 5079 240 5080
rect 274 5083 308 5113
rect 342 5083 381 5117
rect 415 5083 454 5117
rect 488 5083 527 5117
rect 561 5083 600 5117
rect 634 5083 673 5117
rect 707 5083 746 5117
rect 780 5083 819 5117
rect 853 5083 892 5117
rect 926 5083 964 5117
rect 998 5083 1036 5117
rect 1070 5083 1108 5117
rect 1142 5083 1180 5117
rect 1214 5083 1252 5117
rect 1286 5115 1388 5117
rect 1286 5112 1422 5115
rect 1286 5083 1320 5112
rect 274 5079 342 5083
rect 206 5046 342 5079
rect 172 5045 342 5046
rect 172 5041 308 5045
rect 172 5011 240 5041
rect 206 5007 240 5011
rect 274 5011 308 5041
rect 274 5007 342 5011
rect 206 4977 342 5007
rect 1252 5078 1320 5083
rect 1354 5079 1422 5112
rect 1354 5078 1388 5079
rect 1252 5045 1388 5078
rect 1252 5044 1422 5045
rect 1286 5039 1422 5044
rect 1286 5010 1320 5039
rect 1252 5005 1320 5010
rect 1354 5009 1422 5039
rect 1354 5005 1388 5009
rect 172 4973 342 4977
rect 172 4969 308 4973
rect 172 4942 240 4969
rect 206 4935 240 4942
rect 274 4939 308 4969
rect 527 4967 569 5001
rect 603 4967 645 5001
rect 679 4967 721 5001
rect 755 4967 797 5001
rect 831 4967 873 5001
rect 907 4967 948 5001
rect 982 4967 1023 5001
rect 1252 4975 1388 5005
rect 1252 4971 1422 4975
rect 274 4935 342 4939
rect 206 4908 342 4935
rect 172 4901 342 4908
rect 172 4897 308 4901
rect 172 4873 240 4897
rect 206 4863 240 4873
rect 274 4867 308 4897
rect 274 4863 342 4867
rect 206 4839 342 4863
rect 172 4829 342 4839
rect 172 4825 308 4829
rect 172 4804 240 4825
rect 206 4791 240 4804
rect 274 4795 308 4825
rect 274 4791 342 4795
rect 206 4770 342 4791
rect 172 4757 342 4770
rect 172 4753 308 4757
rect 172 4735 240 4753
rect 206 4719 240 4735
rect 274 4723 308 4753
rect 274 4719 342 4723
rect 206 4701 342 4719
rect 172 4685 342 4701
rect 378 4940 436 4956
rect 378 4906 390 4940
rect 424 4906 436 4940
rect 378 4872 436 4906
rect 378 4838 390 4872
rect 424 4838 436 4872
rect 1286 4967 1422 4971
rect 1286 4937 1320 4967
rect 1252 4933 1320 4937
rect 1354 4939 1422 4967
rect 1354 4933 1388 4939
rect 1252 4905 1388 4933
rect 1252 4898 1422 4905
rect 1286 4895 1422 4898
rect 1286 4864 1320 4895
rect 1252 4861 1320 4864
rect 1354 4869 1422 4895
rect 1354 4861 1388 4869
rect 378 4804 436 4838
rect 527 4811 569 4845
rect 603 4811 645 4845
rect 679 4811 721 4845
rect 755 4811 797 4845
rect 831 4811 873 4845
rect 907 4811 948 4845
rect 982 4811 1023 4845
rect 1252 4835 1388 4861
rect 1252 4825 1422 4835
rect 378 4770 390 4804
rect 424 4770 436 4804
rect 378 4736 436 4770
rect 378 4702 390 4736
rect 424 4702 436 4736
rect 378 4686 436 4702
rect 1286 4823 1422 4825
rect 1286 4791 1320 4823
rect 1252 4789 1320 4791
rect 1354 4799 1422 4823
rect 1354 4789 1388 4799
rect 1252 4765 1388 4789
rect 1252 4752 1422 4765
rect 1286 4751 1422 4752
rect 1286 4718 1320 4751
rect 1252 4717 1320 4718
rect 1354 4730 1422 4751
rect 1354 4717 1388 4730
rect 1252 4696 1388 4717
rect 172 4681 308 4685
rect 172 4666 240 4681
rect 206 4647 240 4666
rect 274 4651 308 4681
rect 527 4655 569 4689
rect 603 4655 645 4689
rect 679 4655 721 4689
rect 755 4655 797 4689
rect 831 4655 873 4689
rect 907 4655 948 4689
rect 982 4655 1023 4689
rect 1252 4679 1422 4696
rect 274 4647 342 4651
rect 206 4632 342 4647
rect 172 4612 342 4632
rect 172 4609 308 4612
rect 172 4597 240 4609
rect 206 4575 240 4597
rect 274 4578 308 4609
rect 1286 4645 1320 4679
rect 1354 4661 1422 4679
rect 1354 4645 1388 4661
rect 1252 4627 1388 4645
rect 1252 4607 1422 4627
rect 274 4575 342 4578
rect 206 4563 342 4575
rect 172 4539 342 4563
rect 172 4537 308 4539
rect 172 4527 240 4537
rect 206 4503 240 4527
rect 274 4505 308 4537
rect 274 4503 342 4505
rect 206 4493 342 4503
rect 172 4466 342 4493
rect 390 4532 424 4548
rect 527 4545 569 4579
rect 603 4545 645 4579
rect 679 4545 721 4579
rect 755 4545 797 4579
rect 831 4545 873 4579
rect 907 4545 948 4579
rect 982 4545 1023 4579
rect 1286 4573 1320 4607
rect 1354 4592 1422 4607
rect 1354 4573 1388 4592
rect 1252 4558 1388 4573
rect 390 4476 424 4498
rect 1252 4535 1422 4558
rect 1286 4501 1320 4535
rect 1354 4523 1422 4535
rect 1354 4501 1388 4523
rect 1252 4489 1388 4501
rect 172 4465 308 4466
rect 172 4457 240 4465
rect 206 4431 240 4457
rect 274 4432 308 4465
rect 382 4464 429 4476
rect 382 4449 390 4464
rect 274 4431 342 4432
rect 206 4423 342 4431
rect 172 4393 342 4423
rect 172 4387 240 4393
rect 206 4359 240 4387
rect 274 4359 308 4393
rect 206 4353 342 4359
rect 172 4320 342 4353
rect 172 4317 240 4320
rect 206 4286 240 4317
rect 274 4286 308 4320
rect 206 4283 342 4286
rect 172 4247 342 4283
rect 424 4449 429 4464
rect 1252 4463 1422 4489
rect 390 4396 424 4430
rect 1286 4429 1320 4463
rect 1354 4454 1422 4463
rect 1354 4429 1388 4454
rect 527 4389 569 4423
rect 603 4389 645 4423
rect 679 4389 721 4423
rect 755 4389 797 4423
rect 831 4389 873 4423
rect 907 4389 948 4423
rect 982 4389 1023 4423
rect 1252 4420 1388 4429
rect 1252 4391 1422 4420
rect 390 4328 424 4362
rect 390 4278 424 4294
rect 1286 4357 1320 4391
rect 1354 4385 1422 4391
rect 1354 4357 1388 4385
rect 1252 4351 1388 4357
rect 1252 4319 1422 4351
rect 1286 4285 1320 4319
rect 1354 4316 1422 4319
rect 1354 4285 1388 4316
rect 1252 4282 1388 4285
rect 206 4213 240 4247
rect 274 4213 308 4247
rect 527 4233 569 4267
rect 603 4233 645 4267
rect 679 4233 721 4267
rect 755 4233 797 4267
rect 831 4233 873 4267
rect 907 4233 948 4267
rect 982 4233 1023 4267
rect 1252 4247 1422 4282
rect 172 4189 342 4213
rect 1286 4213 1320 4247
rect 1354 4213 1388 4247
rect 1252 4189 1422 4213
<< viali >>
rect -152 27717 -118 27729
rect -80 27717 -46 27729
rect -152 27695 -150 27717
rect -150 27695 -118 27717
rect -80 27695 -48 27717
rect -48 27695 -46 27717
rect -152 27648 -118 27656
rect -80 27648 -46 27656
rect -152 27622 -150 27648
rect -150 27622 -118 27648
rect -80 27622 -48 27648
rect -48 27622 -46 27648
rect -152 27579 -118 27583
rect -80 27579 -46 27583
rect -152 27549 -150 27579
rect -150 27549 -118 27579
rect -80 27549 -48 27579
rect -48 27549 -46 27579
rect -152 27476 -150 27510
rect -150 27476 -118 27510
rect -80 27476 -48 27510
rect -48 27476 -46 27510
rect -152 27407 -150 27437
rect -150 27407 -118 27437
rect -80 27407 -48 27437
rect -48 27407 -46 27437
rect -152 27403 -118 27407
rect -80 27403 -46 27407
rect -152 27338 -150 27364
rect -150 27338 -118 27364
rect -80 27338 -48 27364
rect -48 27338 -46 27364
rect -152 27330 -118 27338
rect -80 27330 -46 27338
rect -152 27269 -150 27291
rect -150 27269 -118 27291
rect -80 27269 -48 27291
rect -48 27269 -46 27291
rect -152 27257 -118 27269
rect -80 27257 -46 27269
rect -152 27200 -150 27218
rect -150 27200 -118 27218
rect -80 27200 -48 27218
rect -48 27200 -46 27218
rect -152 27184 -118 27200
rect -80 27184 -46 27200
rect -152 27131 -150 27145
rect -150 27131 -118 27145
rect -80 27131 -48 27145
rect -48 27131 -46 27145
rect -152 27111 -118 27131
rect -80 27111 -46 27131
rect -152 27062 -150 27072
rect -150 27062 -118 27072
rect -80 27062 -48 27072
rect -48 27062 -46 27072
rect -152 27038 -118 27062
rect -80 27038 -46 27062
rect -152 26993 -150 26999
rect -150 26993 -118 26999
rect -80 26993 -48 26999
rect -48 26993 -46 26999
rect -152 26965 -118 26993
rect -80 26965 -46 26993
rect -152 26924 -150 26926
rect -150 26924 -118 26926
rect -80 26924 -48 26926
rect -48 26924 -46 26926
rect -152 26892 -118 26924
rect -80 26892 -46 26924
rect -152 26820 -118 26853
rect -80 26820 -46 26853
rect -152 26819 -150 26820
rect -150 26819 -118 26820
rect -80 26819 -48 26820
rect -48 26819 -46 26820
rect -152 26751 -118 26780
rect -80 26751 -46 26780
rect -152 26746 -150 26751
rect -150 26746 -118 26751
rect -80 26746 -48 26751
rect -48 26746 -46 26751
rect -152 26682 -118 26707
rect -80 26682 -46 26707
rect -152 26673 -150 26682
rect -150 26673 -118 26682
rect -80 26673 -48 26682
rect -48 26673 -46 26682
rect -152 26613 -118 26634
rect -80 26613 -46 26634
rect -152 26600 -150 26613
rect -150 26600 -118 26613
rect -80 26600 -48 26613
rect -48 26600 -46 26613
rect -152 26544 -118 26561
rect -80 26544 -46 26561
rect -152 26527 -150 26544
rect -150 26527 -118 26544
rect -80 26527 -48 26544
rect -48 26527 -46 26544
rect -152 26475 -118 26488
rect -80 26475 -46 26488
rect -152 26454 -150 26475
rect -150 26454 -118 26475
rect -80 26454 -48 26475
rect -48 26454 -46 26475
rect -152 26406 -118 26415
rect -80 26406 -46 26415
rect -152 26381 -150 26406
rect -150 26381 -118 26406
rect -80 26381 -48 26406
rect -48 26381 -46 26406
rect -152 26337 -118 26342
rect -80 26337 -46 26342
rect -152 26308 -150 26337
rect -150 26308 -118 26337
rect -80 26308 -48 26337
rect -48 26308 -46 26337
rect -152 26268 -118 26269
rect -80 26268 -46 26269
rect -152 26235 -150 26268
rect -150 26235 -118 26268
rect -80 26235 -48 26268
rect -48 26235 -46 26268
rect -152 26165 -150 26196
rect -150 26165 -118 26196
rect -80 26165 -48 26196
rect -48 26165 -46 26196
rect -152 26162 -118 26165
rect -80 26162 -46 26165
rect -152 26096 -150 26123
rect -150 26096 -118 26123
rect -80 26096 -48 26123
rect -48 26096 -46 26123
rect -152 26089 -118 26096
rect -80 26089 -46 26096
rect -152 26027 -150 26050
rect -150 26027 -118 26050
rect -80 26027 -48 26050
rect -48 26027 -46 26050
rect -152 26016 -118 26027
rect -80 26016 -46 26027
rect -152 25958 -150 25977
rect -150 25958 -118 25977
rect -80 25958 -48 25977
rect -48 25958 -46 25977
rect -152 25943 -118 25958
rect -80 25943 -46 25958
rect -152 25889 -150 25904
rect -150 25889 -118 25904
rect -80 25889 -48 25904
rect -48 25889 -46 25904
rect -152 25870 -118 25889
rect -80 25870 -46 25889
rect -152 25820 -150 25831
rect -150 25820 -118 25831
rect -80 25820 -48 25831
rect -48 25820 -46 25831
rect -152 25797 -118 25820
rect -80 25797 -46 25820
rect -152 25751 -150 25758
rect -150 25751 -118 25758
rect -80 25751 -48 25758
rect -48 25751 -46 25758
rect -152 25724 -118 25751
rect -80 25724 -46 25751
rect -152 25683 -150 25685
rect -150 25683 -118 25685
rect -152 25651 -118 25683
rect -80 25682 -48 25685
rect -48 25682 -46 25685
rect -80 25651 -46 25682
rect -152 25581 -118 25612
rect -152 25578 -150 25581
rect -150 25578 -118 25581
rect -80 25578 -46 25612
rect -152 25513 -118 25539
rect -152 25505 -150 25513
rect -150 25505 -118 25513
rect -80 25509 -46 25539
rect -80 25505 -48 25509
rect -48 25505 -46 25509
rect -152 25445 -118 25466
rect -152 25432 -150 25445
rect -150 25432 -118 25445
rect -80 25440 -46 25466
rect -80 25432 -48 25440
rect -48 25432 -46 25440
rect -152 25377 -118 25393
rect -152 25359 -150 25377
rect -150 25359 -118 25377
rect -80 25371 -46 25393
rect -80 25359 -48 25371
rect -48 25359 -46 25371
rect -152 25309 -118 25320
rect -152 25286 -150 25309
rect -150 25286 -118 25309
rect -80 25302 -46 25320
rect -80 25286 -48 25302
rect -48 25286 -46 25302
rect -152 25241 -118 25247
rect -152 25213 -150 25241
rect -150 25213 -118 25241
rect -80 25233 -46 25247
rect -80 25213 -48 25233
rect -48 25213 -46 25233
rect -152 25173 -118 25174
rect -152 25140 -150 25173
rect -150 25140 -118 25173
rect -80 25164 -46 25175
rect -80 25141 -48 25164
rect -48 25141 -46 25164
rect -152 25071 -150 25101
rect -150 25071 -118 25101
rect -80 25095 -46 25103
rect -152 25067 -118 25071
rect -80 25069 -48 25095
rect -48 25069 -46 25095
rect -152 25003 -150 25028
rect -150 25003 -118 25028
rect -80 25026 -46 25031
rect -152 24994 -118 25003
rect -80 24997 -48 25026
rect -48 24997 -46 25026
rect -80 24957 -46 24959
rect -152 24935 -150 24955
rect -150 24935 -118 24955
rect -152 24921 -118 24935
rect -80 24925 -48 24957
rect -48 24925 -46 24957
rect -152 24867 -150 24882
rect -150 24867 -118 24882
rect -152 24848 -118 24867
rect -80 24854 -48 24887
rect -48 24854 -46 24887
rect -80 24853 -46 24854
rect -152 24799 -150 24809
rect -150 24799 -118 24809
rect -152 24775 -118 24799
rect -80 24785 -48 24815
rect -48 24785 -46 24815
rect -80 24781 -46 24785
rect -152 24731 -150 24736
rect -150 24731 -118 24736
rect -152 24702 -118 24731
rect -80 24716 -48 24743
rect -48 24716 -46 24743
rect -80 24709 -46 24716
rect -152 24629 -118 24663
rect -80 24647 -48 24671
rect -48 24647 -46 24671
rect -80 24637 -46 24647
rect -152 24561 -118 24590
rect -80 24578 -48 24599
rect -48 24578 -46 24599
rect -80 24565 -46 24578
rect -152 24556 -150 24561
rect -150 24556 -118 24561
rect -152 24493 -118 24517
rect -80 24509 -48 24527
rect -48 24509 -46 24527
rect -80 24493 -46 24509
rect -152 24483 -150 24493
rect -150 24483 -118 24493
rect -152 24425 -118 24444
rect -80 24440 -48 24455
rect -48 24440 -46 24455
rect -152 24410 -150 24425
rect -150 24410 -118 24425
rect -80 24421 -46 24440
rect -80 24371 -48 24383
rect -48 24371 -46 24383
rect -152 24357 -118 24371
rect -152 24337 -150 24357
rect -150 24337 -118 24357
rect -80 24349 -46 24371
rect -80 24302 -48 24311
rect -48 24302 -46 24311
rect -152 24289 -118 24298
rect -152 24264 -150 24289
rect -150 24264 -118 24289
rect -80 24277 -46 24302
rect -80 24233 -48 24239
rect -48 24233 -46 24239
rect -152 24221 -118 24225
rect -152 24191 -150 24221
rect -150 24191 -118 24221
rect -80 24205 -46 24233
rect -80 24164 -48 24167
rect -48 24164 -46 24167
rect -152 24119 -150 24152
rect -150 24119 -118 24152
rect -80 24133 -46 24164
rect -152 24118 -118 24119
rect -152 24051 -150 24079
rect -150 24051 -118 24079
rect -80 24061 -46 24095
rect -152 24045 -118 24051
rect -152 23983 -150 24006
rect -150 23983 -118 24006
rect -80 23991 -46 24023
rect -152 23972 -118 23983
rect -80 23989 -48 23991
rect -48 23989 -46 23991
rect -152 23915 -150 23933
rect -150 23915 -118 23933
rect -80 23922 -46 23951
rect -152 23899 -118 23915
rect -80 23917 -48 23922
rect -48 23917 -46 23922
rect -152 23847 -150 23860
rect -150 23847 -118 23860
rect -80 23853 -46 23879
rect -152 23826 -118 23847
rect -80 23845 -48 23853
rect -48 23845 -46 23853
rect -152 23779 -150 23787
rect -150 23779 -118 23787
rect -80 23784 -46 23807
rect -152 23753 -118 23779
rect -80 23773 -48 23784
rect -48 23773 -46 23784
rect -80 23715 -46 23735
rect -152 23711 -150 23714
rect -150 23711 -118 23714
rect -152 23680 -118 23711
rect -80 23701 -48 23715
rect -48 23701 -46 23715
rect -80 23646 -46 23663
rect -152 23609 -118 23641
rect -80 23629 -48 23646
rect -48 23629 -46 23646
rect -152 23607 -150 23609
rect -150 23607 -118 23609
rect -80 23577 -46 23591
rect -152 23541 -118 23568
rect -80 23557 -48 23577
rect -48 23557 -46 23577
rect -152 23534 -150 23541
rect -150 23534 -118 23541
rect -80 23508 -46 23519
rect -152 23473 -118 23495
rect -80 23485 -48 23508
rect -48 23485 -46 23508
rect -152 23461 -150 23473
rect -150 23461 -118 23473
rect -80 23439 -46 23447
rect -152 23388 -118 23422
rect -80 23413 -46 23439
rect -152 23315 -118 23349
rect -80 23341 -46 23375
rect -152 23242 -118 23276
rect -80 23269 -46 23303
rect -152 23169 -118 23203
rect -80 23197 -46 23231
rect -152 23096 -118 23130
rect -80 23125 -46 23159
rect -152 23023 -118 23057
rect -80 23053 -46 23087
rect -152 22950 -118 22984
rect -80 22981 -46 23015
rect 266 27707 299 27709
rect 299 27707 300 27709
rect 341 27707 368 27709
rect 368 27707 375 27709
rect 416 27707 437 27709
rect 437 27707 450 27709
rect 491 27707 506 27709
rect 506 27707 525 27709
rect 566 27707 575 27709
rect 575 27707 600 27709
rect 640 27707 644 27709
rect 644 27707 674 27709
rect 908 27707 920 27709
rect 920 27707 942 27709
rect 983 27707 988 27709
rect 988 27707 1017 27709
rect 1058 27707 1090 27709
rect 1090 27707 1092 27709
rect 1133 27707 1158 27709
rect 1158 27707 1167 27709
rect 1208 27707 1226 27709
rect 1226 27707 1242 27709
rect 1283 27707 1294 27709
rect 1294 27707 1317 27709
rect 1358 27707 1362 27709
rect 1362 27707 1392 27709
rect 1433 27707 1464 27709
rect 1464 27707 1467 27709
rect 1508 27707 1532 27709
rect 1532 27707 1542 27709
rect 1583 27707 1600 27709
rect 1600 27707 1617 27709
rect 1658 27707 1668 27709
rect 1668 27707 1692 27709
rect 1732 27707 1736 27709
rect 1736 27707 1766 27709
rect 1806 27707 1838 27709
rect 1838 27707 1840 27709
rect 1880 27707 1906 27709
rect 1906 27707 1914 27709
rect 1954 27707 1974 27709
rect 1974 27707 1988 27709
rect 2028 27707 2042 27709
rect 2042 27707 2062 27709
rect 2102 27707 2110 27709
rect 2110 27707 2136 27709
rect 2176 27707 2178 27709
rect 2178 27707 2210 27709
rect 2250 27707 2280 27709
rect 2280 27707 2284 27709
rect 2324 27707 2348 27709
rect 2348 27707 2358 27709
rect 2398 27707 2416 27709
rect 2416 27707 2432 27709
rect 2472 27707 2484 27709
rect 2484 27707 2506 27709
rect 2546 27707 2552 27709
rect 2552 27707 2580 27709
rect 2620 27707 2654 27709
rect 2694 27707 2722 27709
rect 2722 27707 2728 27709
rect 2768 27707 2790 27709
rect 2790 27707 2802 27709
rect 2842 27707 2858 27709
rect 2858 27707 2876 27709
rect 2916 27707 2926 27709
rect 2926 27707 2950 27709
rect 266 27675 300 27707
rect 341 27675 375 27707
rect 416 27675 450 27707
rect 491 27675 525 27707
rect 566 27675 600 27707
rect 640 27675 674 27707
rect 908 27675 942 27707
rect 983 27675 1017 27707
rect 1058 27675 1092 27707
rect 1133 27675 1167 27707
rect 1208 27675 1242 27707
rect 1283 27675 1317 27707
rect 1358 27675 1392 27707
rect 1433 27675 1467 27707
rect 1508 27675 1542 27707
rect 1583 27675 1617 27707
rect 1658 27675 1692 27707
rect 1732 27675 1766 27707
rect 1806 27675 1840 27707
rect 1880 27675 1914 27707
rect 1954 27675 1988 27707
rect 2028 27675 2062 27707
rect 2102 27675 2136 27707
rect 2176 27675 2210 27707
rect 2250 27675 2284 27707
rect 2324 27675 2358 27707
rect 2398 27675 2432 27707
rect 2472 27675 2506 27707
rect 2546 27675 2580 27707
rect 2620 27675 2654 27707
rect 2694 27675 2728 27707
rect 2768 27675 2802 27707
rect 2842 27675 2876 27707
rect 2916 27675 2950 27707
rect 300 27605 334 27637
rect 385 27605 419 27637
rect 470 27605 504 27637
rect 555 27605 589 27637
rect 640 27605 674 27637
rect 908 27605 942 27637
rect 983 27605 1017 27637
rect 1058 27605 1092 27637
rect 300 27603 332 27605
rect 332 27603 334 27605
rect 385 27603 402 27605
rect 402 27603 419 27605
rect 470 27603 472 27605
rect 472 27603 504 27605
rect 228 27558 262 27586
rect 228 27552 230 27558
rect 230 27552 262 27558
rect 555 27603 576 27605
rect 576 27603 589 27605
rect 640 27603 646 27605
rect 646 27603 674 27605
rect 908 27603 925 27605
rect 925 27603 942 27605
rect 983 27603 994 27605
rect 994 27603 1017 27605
rect 1058 27603 1063 27605
rect 1063 27603 1092 27605
rect 1133 27603 1167 27637
rect 1208 27605 1242 27637
rect 1283 27605 1317 27637
rect 1358 27605 1392 27637
rect 1433 27605 1467 27637
rect 1508 27605 1542 27637
rect 1583 27605 1617 27637
rect 1658 27605 1692 27637
rect 1732 27605 1766 27637
rect 1806 27605 1840 27637
rect 1880 27605 1914 27637
rect 1954 27605 1988 27637
rect 2028 27605 2062 27637
rect 2102 27605 2136 27637
rect 2176 27605 2210 27637
rect 2250 27605 2284 27637
rect 2324 27605 2358 27637
rect 2398 27605 2432 27637
rect 2472 27605 2506 27637
rect 2546 27605 2580 27637
rect 2620 27605 2654 27637
rect 2694 27605 2728 27637
rect 2768 27605 2802 27637
rect 2842 27605 2876 27637
rect 2916 27605 2950 27637
rect 1208 27603 1236 27605
rect 1236 27603 1242 27605
rect 1283 27603 1305 27605
rect 1305 27603 1317 27605
rect 1358 27603 1374 27605
rect 1374 27603 1392 27605
rect 1433 27603 1443 27605
rect 1443 27603 1467 27605
rect 1508 27603 1512 27605
rect 1512 27603 1542 27605
rect 1583 27603 1615 27605
rect 1615 27603 1617 27605
rect 1658 27603 1684 27605
rect 1684 27603 1692 27605
rect 1732 27603 1753 27605
rect 1753 27603 1766 27605
rect 1806 27603 1822 27605
rect 1822 27603 1840 27605
rect 1880 27603 1891 27605
rect 1891 27603 1914 27605
rect 1954 27603 1960 27605
rect 1960 27603 1988 27605
rect 2028 27603 2029 27605
rect 2029 27603 2062 27605
rect 2102 27603 2133 27605
rect 2133 27603 2136 27605
rect 2176 27603 2202 27605
rect 2202 27603 2210 27605
rect 2250 27603 2271 27605
rect 2271 27603 2284 27605
rect 2324 27603 2340 27605
rect 2340 27603 2358 27605
rect 2398 27603 2409 27605
rect 2409 27603 2432 27605
rect 2472 27603 2478 27605
rect 2478 27603 2506 27605
rect 2546 27603 2547 27605
rect 2547 27603 2580 27605
rect 2620 27603 2650 27605
rect 2650 27603 2654 27605
rect 2694 27603 2719 27605
rect 2719 27603 2728 27605
rect 2768 27603 2788 27605
rect 2788 27603 2802 27605
rect 2842 27603 2857 27605
rect 2857 27603 2876 27605
rect 2916 27603 2926 27605
rect 2926 27603 2950 27605
rect 300 27509 334 27533
rect 228 27485 262 27507
rect 300 27499 332 27509
rect 332 27499 334 27509
rect 228 27473 230 27485
rect 230 27473 262 27485
rect 228 27412 262 27428
rect 300 27412 334 27428
rect 228 27394 230 27412
rect 230 27394 262 27412
rect 300 27394 332 27412
rect 332 27394 334 27412
rect 228 27330 262 27354
rect 300 27330 334 27354
rect 228 27320 230 27330
rect 230 27320 262 27330
rect 300 27320 332 27330
rect 332 27320 334 27330
rect 228 27261 262 27280
rect 228 27246 230 27261
rect 230 27246 262 27261
rect 300 27260 334 27281
rect 300 27247 332 27260
rect 332 27247 334 27260
rect 228 27192 262 27206
rect 228 27172 230 27192
rect 230 27172 262 27192
rect 300 27190 334 27208
rect 300 27174 332 27190
rect 332 27174 334 27190
rect 228 27123 262 27133
rect 228 27099 230 27123
rect 230 27099 262 27123
rect 300 27120 334 27135
rect 300 27101 332 27120
rect 332 27101 334 27120
rect 228 27054 262 27060
rect 228 27026 230 27054
rect 230 27026 262 27054
rect 300 27050 334 27062
rect 300 27028 332 27050
rect 332 27028 334 27050
rect 228 26985 262 26987
rect 228 26953 230 26985
rect 230 26953 262 26985
rect 300 26980 334 26989
rect 300 26955 332 26980
rect 332 26955 334 26980
rect 14592 26964 14626 26998
rect 14664 26964 14698 26998
rect 228 26882 230 26914
rect 230 26882 262 26914
rect 300 26910 334 26916
rect 228 26880 262 26882
rect 300 26882 332 26910
rect 332 26882 334 26910
rect 228 26813 230 26841
rect 230 26813 262 26841
rect 228 26807 262 26813
rect 300 26840 334 26843
rect 300 26809 332 26840
rect 332 26809 334 26840
rect 228 26744 230 26768
rect 230 26744 262 26768
rect 228 26734 262 26744
rect 300 26737 332 26770
rect 332 26737 334 26770
rect 300 26736 334 26737
rect 228 26675 230 26695
rect 230 26675 262 26695
rect 228 26661 262 26675
rect 300 26668 332 26697
rect 332 26668 334 26697
rect 300 26663 334 26668
rect 228 26606 230 26622
rect 230 26606 262 26622
rect 228 26588 262 26606
rect 300 26599 332 26624
rect 332 26599 334 26624
rect 300 26590 334 26599
rect 228 26537 230 26549
rect 230 26537 262 26549
rect 228 26515 262 26537
rect 300 26530 332 26551
rect 332 26530 334 26551
rect 300 26517 334 26530
rect 228 26468 230 26476
rect 230 26468 262 26476
rect 228 26442 262 26468
rect 300 26461 332 26478
rect 332 26461 334 26478
rect 300 26444 334 26461
rect 228 26399 230 26403
rect 230 26399 262 26403
rect 228 26369 262 26399
rect 300 26392 332 26405
rect 332 26392 334 26405
rect 300 26371 334 26392
rect 228 26296 262 26330
rect 300 26323 332 26332
rect 332 26323 334 26332
rect 300 26298 334 26323
rect 228 26226 262 26257
rect 228 26223 230 26226
rect 230 26223 262 26226
rect 300 26254 332 26259
rect 332 26254 334 26259
rect 300 26225 334 26254
rect 300 26185 332 26186
rect 332 26185 334 26186
rect 228 26157 262 26184
rect 228 26150 230 26157
rect 230 26150 262 26157
rect 300 26152 334 26185
rect 228 26088 262 26111
rect 228 26077 230 26088
rect 230 26077 262 26088
rect 300 26081 334 26113
rect 300 26079 332 26081
rect 332 26079 334 26081
rect 228 26019 262 26038
rect 228 26004 230 26019
rect 230 26004 262 26019
rect 300 26012 334 26040
rect 300 26006 332 26012
rect 332 26006 334 26012
rect 228 25950 262 25965
rect 228 25931 230 25950
rect 230 25931 262 25950
rect 300 25943 334 25967
rect 300 25933 332 25943
rect 332 25933 334 25943
rect 228 25881 262 25892
rect 228 25858 230 25881
rect 230 25858 262 25881
rect 300 25874 334 25894
rect 300 25860 332 25874
rect 332 25860 334 25874
rect 228 25812 262 25819
rect 228 25785 230 25812
rect 230 25785 262 25812
rect 300 25805 334 25821
rect 300 25787 332 25805
rect 332 25787 334 25805
rect 228 25743 262 25746
rect 228 25712 230 25743
rect 230 25712 262 25743
rect 300 25736 334 25748
rect 300 25714 332 25736
rect 332 25714 334 25736
rect 228 25640 230 25673
rect 230 25640 262 25673
rect 228 25639 262 25640
rect 300 25667 334 25675
rect 300 25641 332 25667
rect 332 25641 334 25667
rect 228 25571 230 25600
rect 230 25571 262 25600
rect 228 25566 262 25571
rect 300 25598 334 25602
rect 300 25568 332 25598
rect 332 25568 334 25598
rect 228 25502 230 25527
rect 230 25502 262 25527
rect 228 25493 262 25502
rect 300 25495 332 25529
rect 332 25495 334 25529
rect 228 25433 230 25454
rect 230 25433 262 25454
rect 228 25420 262 25433
rect 300 25426 332 25456
rect 332 25426 334 25456
rect 300 25422 334 25426
rect 228 25364 230 25381
rect 230 25364 262 25381
rect 228 25347 262 25364
rect 300 25357 332 25383
rect 332 25357 334 25383
rect 2882 25441 2916 25475
rect 2882 25369 2916 25403
rect 300 25349 334 25357
rect 228 25295 230 25308
rect 230 25295 262 25308
rect 228 25274 262 25295
rect 300 25288 332 25311
rect 332 25288 334 25311
rect 300 25277 334 25288
rect 228 25226 230 25235
rect 230 25226 262 25235
rect 228 25201 262 25226
rect 300 25219 332 25239
rect 332 25219 334 25239
rect 300 25205 334 25219
rect 228 25157 230 25162
rect 230 25157 262 25162
rect 228 25128 262 25157
rect 300 25150 332 25167
rect 332 25150 334 25167
rect 300 25133 334 25150
rect 228 25088 230 25089
rect 230 25088 262 25089
rect 228 25055 262 25088
rect 300 25081 332 25095
rect 332 25081 334 25095
rect 300 25061 334 25081
rect 228 24985 262 25016
rect 300 25012 332 25023
rect 332 25012 334 25023
rect 300 24989 334 25012
rect 228 24982 230 24985
rect 230 24982 262 24985
rect 300 24943 332 24951
rect 332 24943 334 24951
rect 228 24917 262 24943
rect 300 24917 334 24943
rect 228 24909 230 24917
rect 230 24909 262 24917
rect 300 24874 332 24879
rect 332 24874 334 24879
rect 228 24849 262 24870
rect 228 24836 230 24849
rect 230 24836 262 24849
rect 300 24845 334 24874
rect 300 24805 332 24807
rect 332 24805 334 24807
rect 228 24781 262 24797
rect 228 24763 230 24781
rect 230 24763 262 24781
rect 300 24773 334 24805
rect 228 24713 262 24724
rect 228 24690 230 24713
rect 230 24690 262 24713
rect 300 24701 334 24735
rect 228 24645 262 24651
rect 228 24617 230 24645
rect 230 24617 262 24645
rect 300 24632 334 24663
rect 300 24629 332 24632
rect 332 24629 334 24632
rect 228 24577 262 24578
rect 228 24544 230 24577
rect 230 24544 262 24577
rect 300 24563 334 24591
rect 300 24557 332 24563
rect 332 24557 334 24563
rect 228 24475 230 24505
rect 230 24475 262 24505
rect 228 24471 262 24475
rect 300 24494 334 24519
rect 300 24485 332 24494
rect 332 24485 334 24494
rect 228 24407 230 24432
rect 230 24407 262 24432
rect 228 24398 262 24407
rect 300 24425 334 24447
rect 300 24413 332 24425
rect 332 24413 334 24425
rect 228 24339 230 24359
rect 230 24339 262 24359
rect 228 24325 262 24339
rect 300 24356 334 24375
rect 300 24341 332 24356
rect 332 24341 334 24356
rect 228 24271 230 24286
rect 230 24271 262 24286
rect 228 24252 262 24271
rect 300 24287 334 24303
rect 300 24269 332 24287
rect 332 24269 334 24287
rect 228 24203 230 24213
rect 230 24203 262 24213
rect 228 24179 262 24203
rect 300 24218 334 24231
rect 300 24197 332 24218
rect 332 24197 334 24218
rect 228 24135 230 24140
rect 230 24135 262 24140
rect 228 24106 262 24135
rect 300 24149 334 24159
rect 300 24125 332 24149
rect 332 24125 334 24149
rect 228 24033 262 24067
rect 300 24080 334 24087
rect 300 24053 332 24080
rect 332 24053 334 24080
rect 228 23965 262 23994
rect 300 24011 334 24015
rect 300 23981 332 24011
rect 332 23981 334 24011
rect 228 23960 230 23965
rect 230 23960 262 23965
rect 228 23897 262 23921
rect 300 23942 334 23943
rect 300 23909 332 23942
rect 332 23909 334 23942
rect 228 23887 230 23897
rect 230 23887 262 23897
rect 228 23829 262 23848
rect 300 23839 332 23871
rect 332 23839 334 23871
rect 300 23837 334 23839
rect 228 23814 230 23829
rect 230 23814 262 23829
rect 228 23761 262 23775
rect 300 23770 332 23799
rect 332 23770 334 23799
rect 300 23765 334 23770
rect 228 23741 230 23761
rect 230 23741 262 23761
rect 228 23693 262 23702
rect 300 23701 332 23727
rect 332 23701 334 23727
rect 300 23693 334 23701
rect 228 23668 230 23693
rect 230 23668 262 23693
rect 300 23632 332 23655
rect 332 23632 334 23655
rect 228 23625 262 23629
rect 228 23595 230 23625
rect 230 23595 262 23625
rect 300 23621 334 23632
rect 300 23563 332 23583
rect 332 23563 334 23583
rect 228 23523 230 23556
rect 230 23523 262 23556
rect 300 23549 334 23563
rect 228 23522 262 23523
rect 300 23494 332 23511
rect 332 23494 334 23511
rect 228 23455 230 23483
rect 230 23455 262 23483
rect 300 23477 334 23494
rect 228 23449 262 23455
rect 300 23425 332 23439
rect 332 23425 334 23439
rect 228 23387 230 23410
rect 230 23387 262 23410
rect 300 23405 334 23425
rect 228 23376 262 23387
rect 300 23356 332 23367
rect 332 23356 334 23367
rect 228 23319 230 23337
rect 230 23319 262 23337
rect 300 23333 334 23356
rect 701 24203 735 24237
rect 778 24203 812 24237
rect 855 24203 889 24237
rect 932 24203 966 24237
rect 1009 24203 1043 24237
rect 1086 24203 1120 24237
rect 1162 24203 1196 24237
rect 1238 24203 1272 24237
rect 1314 24203 1348 24237
rect 1390 24203 1424 24237
rect 1466 24203 1500 24237
rect 1542 24203 1576 24237
rect 1618 24203 1652 24237
rect 615 24176 649 24182
rect 615 24148 624 24176
rect 624 24148 649 24176
rect 615 24108 649 24110
rect 615 24076 624 24108
rect 624 24076 649 24108
rect 701 24047 735 24081
rect 778 24047 812 24081
rect 855 24047 889 24081
rect 932 24047 966 24081
rect 1009 24047 1043 24081
rect 1086 24047 1120 24081
rect 1162 24047 1196 24081
rect 1238 24047 1272 24081
rect 1314 24047 1348 24081
rect 1390 24047 1424 24081
rect 1466 24047 1500 24081
rect 1542 24047 1576 24081
rect 1618 24047 1652 24081
rect 615 24006 624 24038
rect 624 24006 649 24038
rect 615 24004 649 24006
rect 615 23938 624 23966
rect 624 23938 649 23966
rect 615 23932 649 23938
rect 701 23891 735 23925
rect 778 23891 812 23925
rect 855 23891 889 23925
rect 932 23891 966 23925
rect 1009 23891 1043 23925
rect 1086 23891 1120 23925
rect 1162 23891 1196 23925
rect 1238 23891 1272 23925
rect 1314 23891 1348 23925
rect 1390 23891 1424 23925
rect 1466 23891 1500 23925
rect 1542 23891 1576 23925
rect 1618 23891 1652 23925
rect 701 23781 735 23815
rect 778 23781 812 23815
rect 855 23781 889 23815
rect 932 23781 966 23815
rect 1009 23781 1043 23815
rect 1086 23781 1120 23815
rect 1162 23781 1196 23815
rect 1238 23781 1272 23815
rect 1314 23781 1348 23815
rect 1390 23781 1424 23815
rect 1466 23781 1500 23815
rect 1542 23781 1576 23815
rect 1618 23781 1652 23815
rect 615 23768 649 23779
rect 615 23745 624 23768
rect 624 23745 649 23768
rect 615 23700 649 23707
rect 615 23673 624 23700
rect 624 23673 649 23700
rect 615 23632 649 23635
rect 615 23601 624 23632
rect 624 23601 649 23632
rect 701 23625 735 23659
rect 778 23625 812 23659
rect 855 23625 889 23659
rect 932 23625 966 23659
rect 1009 23625 1043 23659
rect 1086 23625 1120 23659
rect 1162 23625 1196 23659
rect 1238 23625 1272 23659
rect 1314 23625 1348 23659
rect 1390 23625 1424 23659
rect 1466 23625 1500 23659
rect 1542 23625 1576 23659
rect 1618 23625 1652 23659
rect 4410 23745 4412 23779
rect 4412 23745 4444 23779
rect 4482 23745 4514 23779
rect 4514 23745 4516 23779
rect 4822 23745 4824 23779
rect 4824 23745 4856 23779
rect 4894 23745 4926 23779
rect 4926 23745 4928 23779
rect 5234 23745 5236 23779
rect 5236 23745 5268 23779
rect 5306 23745 5338 23779
rect 5338 23745 5340 23779
rect 5646 23745 5648 23779
rect 5648 23745 5680 23779
rect 5718 23745 5750 23779
rect 5750 23745 5752 23779
rect 6058 23745 6060 23779
rect 6060 23745 6092 23779
rect 6130 23745 6162 23779
rect 6162 23745 6164 23779
rect 6470 23745 6472 23779
rect 6472 23745 6504 23779
rect 6542 23745 6574 23779
rect 6574 23745 6576 23779
rect 6882 23745 6884 23779
rect 6884 23745 6916 23779
rect 6954 23745 6986 23779
rect 6986 23745 6988 23779
rect 7294 23745 7296 23779
rect 7296 23745 7328 23779
rect 7366 23745 7398 23779
rect 7398 23745 7400 23779
rect 7706 23745 7708 23779
rect 7708 23745 7740 23779
rect 7778 23745 7810 23779
rect 7810 23745 7812 23779
rect 8118 23745 8120 23779
rect 8120 23745 8152 23779
rect 8190 23745 8222 23779
rect 8222 23745 8224 23779
rect 8530 23745 8532 23779
rect 8532 23745 8564 23779
rect 8602 23745 8634 23779
rect 8634 23745 8636 23779
rect 8942 23745 8944 23779
rect 8944 23745 8976 23779
rect 9014 23745 9046 23779
rect 9046 23745 9048 23779
rect 9354 23745 9356 23779
rect 9356 23745 9388 23779
rect 9426 23745 9458 23779
rect 9458 23745 9460 23779
rect 9766 23745 9768 23779
rect 9768 23745 9800 23779
rect 9838 23745 9870 23779
rect 9870 23745 9872 23779
rect 10178 23745 10180 23779
rect 10180 23745 10212 23779
rect 10250 23745 10282 23779
rect 10282 23745 10284 23779
rect 10590 23745 10592 23779
rect 10592 23745 10624 23779
rect 10662 23745 10694 23779
rect 10694 23745 10696 23779
rect 11002 23745 11004 23779
rect 11004 23745 11036 23779
rect 11074 23745 11106 23779
rect 11106 23745 11108 23779
rect 11244 23745 11278 23779
rect 11316 23745 11350 23779
rect 11414 23745 11416 23779
rect 11416 23745 11448 23779
rect 11486 23745 11518 23779
rect 11518 23745 11520 23779
rect 11620 23745 11654 23779
rect 11692 23745 11726 23779
rect 11826 23745 11828 23779
rect 11828 23745 11860 23779
rect 11898 23745 11930 23779
rect 11930 23745 11932 23779
rect 12032 23745 12066 23779
rect 12104 23745 12138 23779
rect 12238 23745 12240 23779
rect 12240 23745 12272 23779
rect 12310 23745 12342 23779
rect 12342 23745 12344 23779
rect 12444 23745 12478 23779
rect 12516 23745 12550 23779
rect 12650 23745 12652 23779
rect 12652 23745 12684 23779
rect 12722 23745 12754 23779
rect 12754 23745 12756 23779
rect 12856 23745 12890 23779
rect 12928 23745 12962 23779
rect 13062 23745 13064 23779
rect 13064 23745 13096 23779
rect 13134 23745 13166 23779
rect 13166 23745 13168 23779
rect 13268 23745 13302 23779
rect 13340 23745 13374 23779
rect 13474 23745 13476 23779
rect 13476 23745 13508 23779
rect 13546 23745 13578 23779
rect 13578 23745 13580 23779
rect 13680 23745 13714 23779
rect 13752 23745 13786 23779
rect 13886 23745 13888 23779
rect 13888 23745 13920 23779
rect 13958 23745 13990 23779
rect 13990 23745 13992 23779
rect 14092 23745 14126 23779
rect 14164 23745 14198 23779
rect 14298 23745 14300 23779
rect 14300 23745 14332 23779
rect 14370 23745 14402 23779
rect 14402 23745 14404 23779
rect 14468 23745 14502 23779
rect 14540 23745 14574 23779
rect 14656 23745 14690 23779
rect 14728 23745 14746 23779
rect 14746 23745 14762 23779
rect 15124 23745 15158 23779
rect 15196 23745 15226 23779
rect 15226 23745 15230 23779
rect 15536 23745 15570 23779
rect 15608 23745 15638 23779
rect 15638 23745 15642 23779
rect 15948 23745 15982 23779
rect 16020 23745 16050 23779
rect 16050 23745 16054 23779
rect 16360 23745 16394 23779
rect 16432 23745 16462 23779
rect 16462 23745 16466 23779
rect 16772 23745 16806 23779
rect 16844 23745 16874 23779
rect 16874 23745 16878 23779
rect 17115 23745 17149 23779
rect 17187 23745 17218 23779
rect 17218 23745 17221 23779
rect 4410 23665 4444 23699
rect 4482 23665 4516 23699
rect 615 23530 624 23563
rect 624 23530 649 23563
rect 615 23529 649 23530
rect 11244 23665 11278 23699
rect 11316 23665 11350 23699
rect 11002 23588 11036 23622
rect 11074 23588 11108 23622
rect 12032 23665 12066 23699
rect 12104 23665 12138 23699
rect 11620 23588 11654 23622
rect 11692 23588 11726 23622
rect 12856 23665 12890 23699
rect 12928 23665 12962 23699
rect 12444 23588 12478 23622
rect 12516 23588 12550 23622
rect 13680 23665 13714 23699
rect 13752 23665 13786 23699
rect 13268 23588 13302 23622
rect 13340 23588 13374 23622
rect 14468 23665 14502 23699
rect 14540 23665 14574 23699
rect 14092 23588 14126 23622
rect 14164 23588 14198 23622
rect 701 23469 735 23503
rect 778 23469 812 23503
rect 855 23469 889 23503
rect 932 23469 966 23503
rect 1009 23469 1043 23503
rect 1086 23469 1120 23503
rect 1162 23469 1196 23503
rect 1238 23469 1272 23503
rect 1314 23469 1348 23503
rect 1390 23469 1424 23503
rect 1466 23469 1500 23503
rect 1542 23469 1576 23503
rect 1618 23469 1652 23503
rect 2617 23425 2651 23459
rect 2689 23425 2723 23459
rect 228 23303 262 23319
rect 300 23287 332 23295
rect 332 23287 334 23295
rect 228 23251 230 23264
rect 230 23251 262 23264
rect 300 23261 334 23287
rect 228 23230 262 23251
rect 300 23218 332 23223
rect 332 23218 334 23223
rect 228 23183 230 23191
rect 230 23183 262 23191
rect 300 23189 334 23218
rect 228 23157 262 23183
rect 300 23149 332 23151
rect 332 23149 334 23151
rect 373 23149 402 23151
rect 402 23149 407 23151
rect 446 23149 472 23151
rect 472 23149 480 23151
rect 519 23149 542 23151
rect 542 23149 553 23151
rect 592 23149 612 23151
rect 612 23149 626 23151
rect 665 23149 682 23151
rect 682 23149 699 23151
rect 738 23149 752 23151
rect 752 23149 772 23151
rect 811 23149 822 23151
rect 822 23149 845 23151
rect 884 23149 891 23151
rect 891 23149 918 23151
rect 957 23149 960 23151
rect 960 23149 991 23151
rect 1030 23149 1063 23151
rect 1063 23149 1064 23151
rect 1103 23149 1132 23151
rect 1132 23149 1137 23151
rect 1176 23149 1201 23151
rect 1201 23149 1210 23151
rect 1249 23149 1270 23151
rect 1270 23149 1283 23151
rect 1322 23149 1339 23151
rect 1339 23149 1356 23151
rect 1395 23149 1408 23151
rect 1408 23149 1429 23151
rect 1468 23149 1477 23151
rect 1477 23149 1502 23151
rect 1541 23149 1546 23151
rect 1546 23149 1575 23151
rect 1614 23149 1615 23151
rect 1615 23149 1648 23151
rect 1687 23149 1719 23151
rect 1719 23149 1721 23151
rect 1760 23149 1788 23151
rect 1788 23149 1794 23151
rect 1833 23149 1857 23151
rect 1857 23149 1867 23151
rect 1906 23149 1926 23151
rect 1926 23149 1940 23151
rect 1979 23149 1995 23151
rect 1995 23149 2013 23151
rect 2052 23149 2064 23151
rect 2064 23149 2086 23151
rect 2124 23149 2133 23151
rect 2133 23149 2158 23151
rect 2196 23149 2202 23151
rect 2202 23149 2230 23151
rect 2268 23149 2271 23151
rect 2271 23149 2302 23151
rect 2340 23149 2374 23151
rect 2412 23149 2443 23151
rect 2443 23149 2446 23151
rect 2484 23149 2512 23151
rect 2512 23149 2518 23151
rect 2556 23149 2581 23151
rect 2581 23149 2590 23151
rect 2628 23149 2650 23151
rect 2650 23149 2662 23151
rect 2700 23149 2719 23151
rect 2719 23149 2734 23151
rect 2772 23149 2788 23151
rect 2788 23149 2806 23151
rect 2844 23149 2857 23151
rect 2857 23149 2878 23151
rect 2916 23149 2926 23151
rect 2926 23149 2950 23151
rect 300 23117 334 23149
rect 373 23117 407 23149
rect 446 23117 480 23149
rect 519 23117 553 23149
rect 592 23117 626 23149
rect 665 23117 699 23149
rect 738 23117 772 23149
rect 811 23117 845 23149
rect 884 23117 918 23149
rect 957 23117 991 23149
rect 1030 23117 1064 23149
rect 1103 23117 1137 23149
rect 1176 23117 1210 23149
rect 1249 23117 1283 23149
rect 1322 23117 1356 23149
rect 1395 23117 1429 23149
rect 1468 23117 1502 23149
rect 1541 23117 1575 23149
rect 1614 23117 1648 23149
rect 1687 23117 1721 23149
rect 1760 23117 1794 23149
rect 1833 23117 1867 23149
rect 1906 23117 1940 23149
rect 1979 23117 2013 23149
rect 2052 23117 2086 23149
rect 2124 23117 2158 23149
rect 2196 23117 2230 23149
rect 2268 23117 2302 23149
rect 2340 23117 2374 23149
rect 2412 23117 2446 23149
rect 2484 23117 2518 23149
rect 2556 23117 2590 23149
rect 2628 23117 2662 23149
rect 2700 23117 2734 23149
rect 2772 23117 2806 23149
rect 2844 23117 2878 23149
rect 2916 23117 2950 23149
rect 266 23047 300 23079
rect 340 23047 374 23079
rect 414 23047 448 23079
rect 488 23047 522 23079
rect 562 23047 596 23079
rect 636 23047 670 23079
rect 710 23047 744 23079
rect 784 23047 818 23079
rect 858 23047 892 23079
rect 932 23047 966 23079
rect 1006 23047 1040 23079
rect 1080 23047 1114 23079
rect 1154 23047 1188 23079
rect 1228 23047 1262 23079
rect 1302 23047 1336 23079
rect 1376 23047 1410 23079
rect 1450 23047 1484 23079
rect 1524 23047 1558 23079
rect 1598 23047 1632 23079
rect 1672 23047 1706 23079
rect 1746 23047 1780 23079
rect 1820 23047 1854 23079
rect 1894 23047 1928 23079
rect 1967 23047 2001 23079
rect 2040 23047 2074 23079
rect 2113 23047 2147 23079
rect 2186 23047 2220 23079
rect 2259 23047 2293 23079
rect 2332 23047 2366 23079
rect 2405 23047 2439 23079
rect 2478 23047 2512 23079
rect 2551 23047 2585 23079
rect 2624 23047 2658 23079
rect 2697 23047 2731 23079
rect 2770 23047 2804 23079
rect 2843 23047 2877 23079
rect 2916 23047 2950 23079
rect 266 23045 299 23047
rect 299 23045 300 23047
rect 340 23045 368 23047
rect 368 23045 374 23047
rect 414 23045 437 23047
rect 437 23045 448 23047
rect 488 23045 506 23047
rect 506 23045 522 23047
rect 562 23045 575 23047
rect 575 23045 596 23047
rect 636 23045 644 23047
rect 644 23045 670 23047
rect 710 23045 713 23047
rect 713 23045 744 23047
rect 784 23045 816 23047
rect 816 23045 818 23047
rect 858 23045 885 23047
rect 885 23045 892 23047
rect 932 23045 954 23047
rect 954 23045 966 23047
rect 1006 23045 1022 23047
rect 1022 23045 1040 23047
rect 1080 23045 1090 23047
rect 1090 23045 1114 23047
rect 1154 23045 1158 23047
rect 1158 23045 1188 23047
rect 1228 23045 1260 23047
rect 1260 23045 1262 23047
rect 1302 23045 1328 23047
rect 1328 23045 1336 23047
rect 1376 23045 1396 23047
rect 1396 23045 1410 23047
rect 1450 23045 1464 23047
rect 1464 23045 1484 23047
rect 1524 23045 1532 23047
rect 1532 23045 1558 23047
rect 1598 23045 1600 23047
rect 1600 23045 1632 23047
rect 1672 23045 1702 23047
rect 1702 23045 1706 23047
rect 1746 23045 1770 23047
rect 1770 23045 1780 23047
rect 1820 23045 1838 23047
rect 1838 23045 1854 23047
rect 1894 23045 1906 23047
rect 1906 23045 1928 23047
rect 1967 23045 1974 23047
rect 1974 23045 2001 23047
rect 2040 23045 2042 23047
rect 2042 23045 2074 23047
rect 2113 23045 2144 23047
rect 2144 23045 2147 23047
rect 2186 23045 2212 23047
rect 2212 23045 2220 23047
rect 2259 23045 2280 23047
rect 2280 23045 2293 23047
rect 2332 23045 2348 23047
rect 2348 23045 2366 23047
rect 2405 23045 2416 23047
rect 2416 23045 2439 23047
rect 2478 23045 2484 23047
rect 2484 23045 2512 23047
rect 2551 23045 2552 23047
rect 2552 23045 2585 23047
rect 2624 23045 2654 23047
rect 2654 23045 2658 23047
rect 2697 23045 2722 23047
rect 2722 23045 2731 23047
rect 2770 23045 2790 23047
rect 2790 23045 2804 23047
rect 2843 23045 2858 23047
rect 2858 23045 2877 23047
rect 2916 23045 2926 23047
rect 2926 23045 2950 23047
rect -152 22877 -118 22911
rect -80 22909 -46 22943
rect -152 22804 -118 22838
rect -80 22837 -46 22871
rect -80 22765 -46 22799
rect -152 22731 -118 22765
rect -80 22725 -46 22727
rect -5 22725 21 22727
rect 21 22725 29 22727
rect 70 22725 90 22727
rect 90 22725 104 22727
rect 144 22725 159 22727
rect 159 22725 178 22727
rect 218 22725 228 22727
rect 228 22725 252 22727
rect 292 22725 297 22727
rect 297 22725 326 22727
rect 366 22725 400 22727
rect 440 22725 469 22727
rect 469 22725 474 22727
rect 514 22725 538 22727
rect 538 22725 548 22727
rect 588 22725 607 22727
rect 607 22725 622 22727
rect 662 22725 676 22727
rect 676 22725 696 22727
rect 736 22725 745 22727
rect 745 22725 770 22727
rect -80 22693 -46 22725
rect -5 22693 29 22725
rect 70 22693 104 22725
rect 144 22693 178 22725
rect 218 22693 252 22725
rect 292 22693 326 22725
rect 366 22693 400 22725
rect 440 22693 474 22725
rect 514 22693 548 22725
rect 588 22693 622 22725
rect 662 22693 696 22725
rect 736 22693 770 22725
rect 810 22693 844 22727
rect 884 22693 918 22727
rect 958 22693 992 22727
rect 1032 22693 1066 22727
rect 1106 22693 1140 22727
rect 1180 22693 1214 22727
rect 1254 22693 1288 22727
rect 1328 22693 1362 22727
rect 1402 22693 1436 22727
rect 1476 22693 1510 22727
rect 1550 22693 1584 22727
rect 1624 22693 1658 22727
rect 1698 22693 1732 22727
rect 1772 22693 1806 22727
rect 1846 22693 1880 22727
rect 1920 22693 1954 22727
rect 1994 22693 2028 22727
rect 2068 22693 2102 22727
rect 2142 22693 2174 22727
rect 2174 22693 2176 22727
rect -114 22621 -80 22655
rect -41 22623 -7 22655
rect 32 22623 66 22655
rect 105 22623 139 22655
rect 178 22623 212 22655
rect 251 22623 285 22655
rect 324 22623 358 22655
rect 397 22623 431 22655
rect 470 22623 504 22655
rect 543 22623 577 22655
rect 616 22623 650 22655
rect 689 22623 723 22655
rect 762 22623 796 22655
rect 835 22623 869 22655
rect 908 22623 942 22655
rect 981 22623 1015 22655
rect 1054 22623 1088 22655
rect 1127 22623 1161 22655
rect 1200 22623 1234 22655
rect 1273 22623 1307 22655
rect -41 22621 -10 22623
rect -10 22621 -7 22623
rect 32 22621 60 22623
rect 60 22621 66 22623
rect 105 22621 130 22623
rect 130 22621 139 22623
rect 178 22621 200 22623
rect 200 22621 212 22623
rect 251 22621 270 22623
rect 270 22621 285 22623
rect 324 22621 340 22623
rect 340 22621 358 22623
rect 397 22621 410 22623
rect 410 22621 431 22623
rect 470 22621 480 22623
rect 480 22621 504 22623
rect 543 22621 550 22623
rect 550 22621 577 22623
rect 616 22621 620 22623
rect 620 22621 650 22623
rect 689 22621 690 22623
rect 690 22621 723 22623
rect 762 22621 794 22623
rect 794 22621 796 22623
rect 835 22621 863 22623
rect 863 22621 869 22623
rect 908 22621 932 22623
rect 932 22621 942 22623
rect 981 22621 1001 22623
rect 1001 22621 1015 22623
rect 1054 22621 1070 22623
rect 1070 22621 1088 22623
rect 1127 22621 1139 22623
rect 1139 22621 1161 22623
rect 1200 22621 1208 22623
rect 1208 22621 1234 22623
rect 1273 22621 1277 22623
rect 1277 22621 1307 22623
rect 1346 22621 1380 22655
rect 1419 22623 1453 22655
rect 1492 22623 1526 22655
rect 1565 22623 1599 22655
rect 1638 22623 1672 22655
rect 1710 22623 1744 22655
rect 1782 22623 1816 22655
rect 1854 22623 1888 22655
rect 1926 22623 1960 22655
rect 1998 22623 2032 22655
rect 2070 22623 2104 22655
rect 2142 22623 2176 22655
rect 1419 22621 1450 22623
rect 1450 22621 1453 22623
rect 1492 22621 1519 22623
rect 1519 22621 1526 22623
rect 1565 22621 1588 22623
rect 1588 22621 1599 22623
rect 1638 22621 1657 22623
rect 1657 22621 1672 22623
rect 1710 22621 1726 22623
rect 1726 22621 1744 22623
rect 1782 22621 1795 22623
rect 1795 22621 1816 22623
rect 1854 22621 1864 22623
rect 1864 22621 1888 22623
rect 1926 22621 1933 22623
rect 1933 22621 1960 22623
rect 1998 22621 2002 22623
rect 2002 22621 2032 22623
rect 2070 22621 2071 22623
rect 2071 22621 2104 22623
rect 2142 22621 2174 22623
rect 2174 22621 2176 22623
rect -2089 18309 -2055 18343
rect -2016 18309 -1982 18343
rect -1943 18309 -1909 18343
rect -1870 18309 -1836 18343
rect -1797 18309 -1763 18343
rect -1724 18309 -1690 18343
rect -1651 18309 -1617 18343
rect -1578 18309 -1544 18343
rect -1505 18309 -1471 18343
rect -1432 18309 -1398 18343
rect -1359 18309 -1325 18343
rect -1286 18309 -1252 18343
rect -1213 18309 -1179 18343
rect -1140 18309 -1106 18343
rect -1067 18309 -1033 18343
rect -994 18309 -960 18343
rect -921 18309 -887 18343
rect -848 18309 -814 18343
rect -775 18309 -741 18343
rect -702 18309 -668 18343
rect -629 18309 -595 18343
rect -556 18309 -522 18343
rect -483 18309 -449 18343
rect -410 18309 -376 18343
rect -337 18309 -303 18343
rect -264 18309 -230 18343
rect -191 18309 -157 18343
rect -118 18309 -84 18343
rect -45 18309 -11 18343
rect 28 18309 62 18343
rect 101 18309 135 18343
rect 174 18309 208 18343
rect 247 18309 281 18343
rect 320 18309 354 18343
rect 393 18309 427 18343
rect 466 18309 500 18343
rect 539 18309 573 18343
rect 612 18309 646 18343
rect 685 18309 719 18343
rect 758 18309 792 18343
rect 831 18309 865 18343
rect 904 18309 938 18343
rect 977 18309 1011 18343
rect 1050 18309 1084 18343
rect 1123 18309 1157 18343
rect 1196 18309 1230 18343
rect 1269 18309 1303 18343
rect 1342 18309 1376 18343
rect 1415 18309 1449 18343
rect 1488 18309 1522 18343
rect 1561 18309 1595 18343
rect 1634 18309 1668 18343
rect 1707 18309 1741 18343
rect -2199 18271 -2165 18305
rect -2127 18237 -2093 18271
rect -2055 18237 -2021 18271
rect -1983 18237 -1949 18271
rect -1911 18237 -1877 18271
rect -1839 18237 -1805 18271
rect -1767 18237 -1733 18271
rect -1695 18237 -1661 18271
rect -1623 18237 -1589 18271
rect -1551 18237 -1517 18271
rect -1479 18237 -1445 18271
rect -1407 18237 -1373 18271
rect -1335 18237 -1301 18271
rect -1263 18237 -1229 18271
rect -1191 18237 -1157 18271
rect -1119 18237 -1085 18271
rect -1047 18237 -1013 18271
rect -975 18237 -941 18271
rect -903 18237 -869 18271
rect -831 18237 -797 18271
rect -759 18237 -725 18271
rect -687 18237 -653 18271
rect -615 18237 -581 18271
rect -543 18237 -509 18271
rect -471 18237 -437 18271
rect -399 18237 -365 18271
rect -327 18237 -293 18271
rect -255 18237 -221 18271
rect -183 18237 -149 18271
rect -111 18237 -77 18271
rect -39 18237 -5 18271
rect 33 18237 67 18271
rect 105 18237 139 18271
rect 177 18237 211 18271
rect 249 18237 283 18271
rect 321 18237 355 18271
rect 393 18237 427 18271
rect 466 18237 500 18271
rect 539 18237 573 18271
rect 612 18237 646 18271
rect 685 18237 719 18271
rect 758 18237 792 18271
rect 831 18237 865 18271
rect 904 18237 938 18271
rect 977 18237 1011 18271
rect 1050 18237 1084 18271
rect 1123 18237 1157 18271
rect 1196 18237 1230 18271
rect 1269 18237 1303 18271
rect 1342 18237 1376 18271
rect 1415 18237 1449 18271
rect 1488 18237 1522 18271
rect 1561 18237 1595 18271
rect 1634 18237 1668 18271
rect 1707 18237 1741 18271
rect -2199 18199 -2165 18233
rect -2199 18127 -2165 18161
rect -2127 18146 -2093 18180
rect -2199 18055 -2165 18089
rect -2127 18055 -2093 18089
rect 493 4967 527 5001
rect 569 4967 603 5001
rect 645 4967 679 5001
rect 721 4967 755 5001
rect 797 4967 831 5001
rect 873 4967 907 5001
rect 948 4967 982 5001
rect 1023 4967 1057 5001
rect 493 4811 527 4845
rect 569 4811 603 4845
rect 645 4811 679 4845
rect 721 4811 755 4845
rect 797 4811 831 4845
rect 873 4811 907 4845
rect 948 4811 982 4845
rect 1023 4811 1057 4845
rect 493 4655 527 4689
rect 569 4655 603 4689
rect 645 4655 679 4689
rect 721 4655 755 4689
rect 797 4655 831 4689
rect 873 4655 907 4689
rect 948 4655 982 4689
rect 1023 4655 1057 4689
rect 493 4545 527 4579
rect 569 4545 603 4579
rect 645 4545 679 4579
rect 721 4545 755 4579
rect 797 4545 831 4579
rect 873 4545 907 4579
rect 948 4545 982 4579
rect 1023 4545 1057 4579
rect 493 4389 527 4423
rect 569 4389 603 4423
rect 645 4389 679 4423
rect 721 4389 755 4423
rect 797 4389 831 4423
rect 873 4389 907 4423
rect 948 4389 982 4423
rect 1023 4389 1057 4423
rect 493 4233 527 4267
rect 569 4233 603 4267
rect 645 4233 679 4267
rect 721 4233 755 4267
rect 797 4233 831 4267
rect 873 4233 907 4267
rect 948 4233 982 4267
rect 1023 4233 1057 4267
<< metal1 >>
rect -158 27729 -40 27741
rect -158 27695 -152 27729
rect -118 27695 -80 27729
rect -46 27695 -40 27729
rect -158 27656 -40 27695
rect -158 27622 -152 27656
rect -118 27622 -80 27656
rect -46 27622 -40 27656
rect -158 27583 -40 27622
rect -158 27549 -152 27583
rect -118 27549 -80 27583
rect -46 27549 -40 27583
rect -158 27510 -40 27549
rect -158 27476 -152 27510
rect -118 27476 -80 27510
rect -46 27476 -40 27510
rect -158 27437 -40 27476
rect -158 27403 -152 27437
rect -118 27403 -80 27437
rect -46 27403 -40 27437
rect -158 27364 -40 27403
rect -158 27330 -152 27364
rect -118 27330 -80 27364
rect -46 27330 -40 27364
rect -158 27291 -40 27330
rect -158 27257 -152 27291
rect -118 27257 -80 27291
rect -46 27257 -40 27291
rect -158 27218 -40 27257
rect -158 27184 -152 27218
rect -118 27184 -80 27218
rect -46 27184 -40 27218
rect -158 27145 -40 27184
rect -158 27111 -152 27145
rect -118 27111 -80 27145
rect -46 27111 -40 27145
rect -158 27072 -40 27111
rect -158 27038 -152 27072
rect -118 27038 -80 27072
rect -46 27038 -40 27072
rect -158 26999 -40 27038
rect -158 26965 -152 26999
rect -118 26965 -80 26999
rect -46 26965 -40 26999
rect -158 26926 -40 26965
rect -158 26892 -152 26926
rect -118 26892 -80 26926
rect -46 26892 -40 26926
rect -158 26853 -40 26892
rect -158 26819 -152 26853
rect -118 26819 -80 26853
rect -46 26819 -40 26853
rect -158 26780 -40 26819
rect -158 26746 -152 26780
rect -118 26746 -80 26780
rect -46 26746 -40 26780
rect -158 26707 -40 26746
rect -158 26673 -152 26707
rect -118 26673 -80 26707
rect -46 26673 -40 26707
rect -158 26634 -40 26673
rect -158 26600 -152 26634
rect -118 26600 -80 26634
rect -46 26600 -40 26634
rect -158 26561 -40 26600
rect -158 26527 -152 26561
rect -118 26527 -80 26561
rect -46 26527 -40 26561
rect -158 26488 -40 26527
rect -158 26454 -152 26488
rect -118 26454 -80 26488
rect -46 26454 -40 26488
rect -158 26415 -40 26454
rect -158 26381 -152 26415
rect -118 26381 -80 26415
rect -46 26381 -40 26415
rect -158 26342 -40 26381
rect -158 26308 -152 26342
rect -118 26308 -80 26342
rect -46 26308 -40 26342
rect -158 26269 -40 26308
rect -158 26235 -152 26269
rect -118 26235 -80 26269
rect -46 26235 -40 26269
rect -158 26196 -40 26235
rect -158 26162 -152 26196
rect -118 26162 -80 26196
rect -46 26162 -40 26196
rect -158 26123 -40 26162
rect -158 26089 -152 26123
rect -118 26089 -80 26123
rect -46 26089 -40 26123
rect -158 26050 -40 26089
rect -158 26016 -152 26050
rect -118 26016 -80 26050
rect -46 26016 -40 26050
rect -158 25977 -40 26016
rect -158 25943 -152 25977
rect -118 25943 -80 25977
rect -46 25943 -40 25977
rect -158 25904 -40 25943
rect -158 25870 -152 25904
rect -118 25870 -80 25904
rect -46 25870 -40 25904
rect -158 25831 -40 25870
rect -158 25797 -152 25831
rect -118 25797 -80 25831
rect -46 25797 -40 25831
rect -158 25758 -40 25797
rect -158 25724 -152 25758
rect -118 25724 -80 25758
rect -46 25724 -40 25758
rect -158 25685 -40 25724
rect -158 25651 -152 25685
rect -118 25651 -80 25685
rect -46 25651 -40 25685
rect -158 25612 -40 25651
rect -158 25578 -152 25612
rect -118 25578 -80 25612
rect -46 25578 -40 25612
rect -158 25539 -40 25578
rect -158 25505 -152 25539
rect -118 25505 -80 25539
rect -46 25505 -40 25539
rect -158 25466 -40 25505
rect -158 25432 -152 25466
rect -118 25432 -80 25466
rect -46 25432 -40 25466
rect -158 25393 -40 25432
rect -158 25359 -152 25393
rect -118 25359 -80 25393
rect -46 25359 -40 25393
rect -158 25320 -40 25359
rect -158 25286 -152 25320
rect -118 25286 -80 25320
rect -46 25286 -40 25320
rect -158 25247 -40 25286
rect -158 25213 -152 25247
rect -118 25213 -80 25247
rect -46 25213 -40 25247
rect -158 25175 -40 25213
rect -158 25174 -80 25175
rect -158 25140 -152 25174
rect -118 25141 -80 25174
rect -46 25141 -40 25175
rect -118 25140 -40 25141
rect -158 25103 -40 25140
rect -158 25101 -80 25103
rect -158 25067 -152 25101
rect -118 25069 -80 25101
rect -46 25069 -40 25103
rect -118 25067 -40 25069
rect -158 25031 -40 25067
rect -158 25028 -80 25031
rect -158 24994 -152 25028
rect -118 24997 -80 25028
rect -46 24997 -40 25031
rect -118 24994 -40 24997
rect -158 24959 -40 24994
rect -158 24955 -80 24959
rect -158 24921 -152 24955
rect -118 24925 -80 24955
rect -46 24925 -40 24959
rect -118 24921 -40 24925
rect -158 24887 -40 24921
rect -158 24882 -80 24887
rect -158 24848 -152 24882
rect -118 24853 -80 24882
rect -46 24853 -40 24887
rect -118 24848 -40 24853
rect -158 24815 -40 24848
rect -158 24809 -80 24815
rect -158 24775 -152 24809
rect -118 24781 -80 24809
rect -46 24781 -40 24815
rect -118 24775 -40 24781
rect -158 24743 -40 24775
rect -158 24736 -80 24743
rect -158 24702 -152 24736
rect -118 24709 -80 24736
rect -46 24709 -40 24743
rect -118 24702 -40 24709
rect -158 24671 -40 24702
rect -158 24663 -80 24671
rect -158 24629 -152 24663
rect -118 24637 -80 24663
rect -46 24637 -40 24671
rect -118 24629 -40 24637
rect -158 24599 -40 24629
rect -158 24590 -80 24599
rect -158 24556 -152 24590
rect -118 24565 -80 24590
rect -46 24565 -40 24599
rect -118 24556 -40 24565
rect -158 24527 -40 24556
rect -158 24517 -80 24527
rect -158 24483 -152 24517
rect -118 24493 -80 24517
rect -46 24493 -40 24527
rect -118 24483 -40 24493
rect -158 24455 -40 24483
rect -158 24444 -80 24455
rect -158 24410 -152 24444
rect -118 24421 -80 24444
rect -46 24421 -40 24455
rect -118 24410 -40 24421
rect -158 24383 -40 24410
rect -158 24371 -80 24383
rect -158 24337 -152 24371
rect -118 24349 -80 24371
rect -46 24349 -40 24383
rect -118 24337 -40 24349
rect -158 24311 -40 24337
rect -158 24298 -80 24311
rect -158 24264 -152 24298
rect -118 24277 -80 24298
rect -46 24277 -40 24311
rect -118 24264 -40 24277
rect -158 24239 -40 24264
rect -158 24225 -80 24239
rect -158 24191 -152 24225
rect -118 24205 -80 24225
rect -46 24205 -40 24239
rect -118 24191 -40 24205
rect -158 24167 -40 24191
rect -158 24152 -80 24167
rect -158 24118 -152 24152
rect -118 24133 -80 24152
rect -46 24133 -40 24167
rect -118 24118 -40 24133
rect -158 24095 -40 24118
rect -158 24079 -80 24095
rect -158 24045 -152 24079
rect -118 24061 -80 24079
rect -46 24061 -40 24095
rect -118 24045 -40 24061
rect -158 24023 -40 24045
rect -158 24006 -80 24023
rect -158 23972 -152 24006
rect -118 23989 -80 24006
rect -46 23989 -40 24023
rect -118 23972 -40 23989
rect -158 23951 -40 23972
rect -158 23933 -80 23951
rect -158 23899 -152 23933
rect -118 23917 -80 23933
rect -46 23917 -40 23951
rect -118 23899 -40 23917
rect -158 23879 -40 23899
rect -158 23860 -80 23879
rect -158 23826 -152 23860
rect -118 23845 -80 23860
rect -46 23845 -40 23879
rect -118 23826 -40 23845
rect -158 23807 -40 23826
rect -158 23787 -80 23807
rect -158 23753 -152 23787
rect -118 23773 -80 23787
rect -46 23773 -40 23807
rect -118 23753 -40 23773
rect -158 23735 -40 23753
rect -158 23714 -80 23735
rect -158 23680 -152 23714
rect -118 23701 -80 23714
rect -46 23701 -40 23735
rect -118 23680 -40 23701
rect -158 23663 -40 23680
rect -158 23641 -80 23663
rect -158 23607 -152 23641
rect -118 23629 -80 23641
rect -46 23629 -40 23663
rect -118 23607 -40 23629
rect -158 23591 -40 23607
rect -158 23568 -80 23591
rect -158 23534 -152 23568
rect -118 23557 -80 23568
rect -46 23557 -40 23591
rect -118 23534 -40 23557
rect -158 23519 -40 23534
rect -158 23495 -80 23519
rect -158 23461 -152 23495
rect -118 23485 -80 23495
rect -46 23485 -40 23519
rect -118 23461 -40 23485
rect -158 23447 -40 23461
rect -158 23422 -80 23447
rect -158 23388 -152 23422
rect -118 23413 -80 23422
rect -46 23413 -40 23447
rect -118 23388 -40 23413
rect -158 23375 -40 23388
rect -158 23349 -80 23375
rect -158 23315 -152 23349
rect -118 23341 -80 23349
rect -46 23341 -40 23375
rect -118 23315 -40 23341
rect -158 23303 -40 23315
rect -158 23276 -80 23303
rect -158 23242 -152 23276
rect -118 23269 -80 23276
rect -46 23269 -40 23303
rect -118 23242 -40 23269
rect -158 23231 -40 23242
rect -158 23203 -80 23231
rect -158 23169 -152 23203
rect -118 23197 -80 23203
rect -46 23197 -40 23231
rect -118 23169 -40 23197
rect -158 23159 -40 23169
rect -158 23130 -80 23159
rect -158 23096 -152 23130
rect -118 23125 -80 23130
rect -46 23125 -40 23159
rect -118 23096 -40 23125
rect -158 23087 -40 23096
rect -158 23057 -80 23087
tri -178 23023 -158 23043 se
rect -158 23023 -152 23057
rect -118 23053 -80 23057
rect -46 23053 -40 23087
rect -118 23023 -40 23053
rect 222 27709 686 27721
rect 222 27675 266 27709
rect 300 27675 341 27709
rect 375 27675 416 27709
rect 450 27675 491 27709
rect 525 27675 566 27709
rect 600 27675 640 27709
rect 674 27675 686 27709
rect 222 27637 686 27675
rect 222 27603 300 27637
rect 334 27603 385 27637
rect 419 27603 470 27637
rect 504 27603 555 27637
rect 589 27603 640 27637
rect 674 27603 686 27637
rect 222 27597 686 27603
rect 896 27709 3100 27721
rect 896 27675 908 27709
rect 942 27675 983 27709
rect 1017 27675 1058 27709
rect 1092 27675 1133 27709
rect 1167 27675 1208 27709
rect 1242 27675 1283 27709
rect 1317 27675 1358 27709
rect 1392 27675 1433 27709
rect 1467 27675 1508 27709
rect 1542 27675 1583 27709
rect 1617 27675 1658 27709
rect 1692 27675 1732 27709
rect 1766 27675 1806 27709
rect 1840 27675 1880 27709
rect 1914 27675 1954 27709
rect 1988 27675 2028 27709
rect 2062 27675 2102 27709
rect 2136 27675 2176 27709
rect 2210 27675 2250 27709
rect 2284 27675 2324 27709
rect 2358 27675 2398 27709
rect 2432 27675 2472 27709
rect 2506 27675 2546 27709
rect 2580 27675 2620 27709
rect 2654 27675 2694 27709
rect 2728 27675 2768 27709
rect 2802 27675 2842 27709
rect 2876 27675 2916 27709
rect 2950 27675 3100 27709
rect 896 27637 3100 27675
rect 896 27603 908 27637
rect 942 27603 983 27637
rect 1017 27603 1058 27637
rect 1092 27603 1133 27637
rect 1167 27603 1208 27637
rect 1242 27603 1283 27637
rect 1317 27603 1358 27637
rect 1392 27603 1433 27637
rect 1467 27603 1508 27637
rect 1542 27603 1583 27637
rect 1617 27603 1658 27637
rect 1692 27603 1732 27637
rect 1766 27603 1806 27637
rect 1840 27603 1880 27637
rect 1914 27603 1954 27637
rect 1988 27603 2028 27637
rect 2062 27603 2102 27637
rect 2136 27603 2176 27637
rect 2210 27603 2250 27637
rect 2284 27603 2324 27637
rect 2358 27603 2398 27637
rect 2432 27603 2472 27637
rect 2506 27603 2546 27637
rect 2580 27603 2620 27637
rect 2654 27603 2694 27637
rect 2728 27603 2768 27637
rect 2802 27603 2842 27637
rect 2876 27603 2916 27637
rect 2950 27603 3100 27637
rect 896 27597 3100 27603
rect 222 27586 340 27597
rect 222 27552 228 27586
rect 262 27552 340 27586
tri 2845 27563 2879 27597 ne
rect 2879 27563 3100 27597
rect 222 27533 340 27552
rect 222 27507 300 27533
rect 222 27473 228 27507
rect 262 27499 300 27507
rect 334 27499 340 27533
tri 2879 27511 2931 27563 ne
rect 2931 27511 3100 27563
rect 10777 27511 10783 27563
rect 10835 27511 10847 27563
rect 10899 27511 18478 27563
rect 262 27473 340 27499
tri 2931 27483 2959 27511 ne
rect 2959 27483 3100 27511
rect 222 27428 340 27473
tri 2959 27472 2970 27483 ne
rect 2970 27472 3100 27483
rect 10820 27431 10826 27483
rect 10878 27431 10890 27483
rect 10942 27473 18397 27483
tri 18397 27473 18407 27483 sw
rect 10942 27431 18407 27473
tri 18407 27431 18449 27473 sw
rect 222 27394 228 27428
rect 262 27394 300 27428
rect 334 27394 340 27428
tri 18375 27399 18407 27431 ne
rect 18407 27399 18449 27431
tri 18449 27399 18481 27431 sw
rect 222 27354 340 27394
tri 18407 27382 18424 27399 ne
rect 18424 27382 18481 27399
tri 18424 27377 18429 27382 ne
rect 222 27320 228 27354
rect 262 27320 300 27354
rect 334 27320 340 27354
rect 18429 27351 18481 27382
rect 222 27281 340 27320
rect 222 27280 300 27281
rect 222 27246 228 27280
rect 262 27247 300 27280
rect 334 27247 340 27281
rect 262 27246 340 27247
rect 222 27208 340 27246
rect 6633 27229 6639 27345
rect 6819 27229 6825 27345
rect 222 27206 300 27208
rect 222 27172 228 27206
rect 262 27174 300 27206
rect 334 27174 340 27208
rect 262 27172 340 27174
rect 222 27135 340 27172
rect 222 27133 300 27135
rect 222 27099 228 27133
rect 262 27101 300 27133
rect 334 27101 340 27135
rect 262 27099 340 27101
rect 222 27062 340 27099
rect 222 27060 300 27062
rect 222 27026 228 27060
rect 262 27028 300 27060
rect 334 27028 340 27062
rect 262 27026 340 27028
rect 222 26989 340 27026
tri 14672 27024 14869 27221 ne
rect 222 26987 300 26989
rect 222 26953 228 26987
rect 262 26955 300 26987
rect 334 26955 340 26989
rect 4191 26955 4197 27007
rect 4249 26955 4261 27007
rect 4313 26998 14722 27007
rect 4313 26964 14592 26998
rect 14626 26964 14664 26998
rect 14698 26964 14722 26998
rect 4313 26955 14722 26964
rect 262 26953 340 26955
rect 222 26916 340 26953
rect 222 26914 300 26916
rect 222 26880 228 26914
rect 262 26882 300 26914
rect 334 26882 340 26916
rect 262 26880 340 26882
rect 14869 26880 15069 27221
tri 15069 27024 15266 27221 nw
tri 15496 27024 15693 27221 ne
rect 15693 26972 15893 27221
tri 15893 27024 16090 27221 nw
tri 16320 27024 16517 27221 ne
rect 15694 26970 15892 26971
rect 15693 26934 15893 26970
rect 15694 26933 15892 26934
rect 15693 26880 15893 26932
rect 16517 26972 16717 27221
tri 16717 27024 16914 27221 nw
tri 17144 27024 17341 27221 ne
rect 16518 26970 16716 26971
rect 16517 26934 16717 26970
rect 16518 26933 16716 26934
rect 16517 26880 16717 26932
rect 17341 26994 17634 27221
tri 17550 26992 17552 26994 ne
rect 17552 26992 17634 26994
rect 17341 26990 17550 26992
tri 17550 26990 17552 26992 sw
tri 17552 26990 17554 26992 ne
rect 17554 26990 17634 26992
rect 17341 26988 17552 26990
tri 17552 26988 17554 26990 sw
tri 17554 26988 17556 26990 ne
rect 17556 26988 17634 26990
rect 17341 26986 17554 26988
tri 17554 26986 17556 26988 sw
tri 17556 26986 17558 26988 ne
rect 17558 26986 17634 26988
rect 17341 26984 17556 26986
tri 17556 26984 17558 26986 sw
tri 17558 26984 17560 26986 ne
rect 17560 26984 17634 26986
rect 17341 26982 17558 26984
tri 17558 26982 17560 26984 sw
tri 17560 26982 17562 26984 ne
rect 17562 26982 17634 26984
rect 17341 26980 17560 26982
tri 17560 26980 17562 26982 sw
tri 17562 26980 17564 26982 ne
rect 17564 26980 17634 26982
rect 17341 26978 17562 26980
tri 17562 26978 17564 26980 sw
tri 17564 26978 17566 26980 ne
rect 17566 26978 17634 26980
rect 17341 26976 17564 26978
tri 17564 26976 17566 26978 sw
tri 17566 26976 17568 26978 ne
rect 17568 26976 17634 26978
rect 17341 26974 17566 26976
tri 17566 26974 17568 26976 sw
tri 17568 26974 17570 26976 ne
rect 17570 26974 17634 26976
rect 17341 26972 17568 26974
tri 17568 26972 17570 26974 sw
tri 17570 26972 17572 26974 ne
rect 17572 26972 17634 26974
rect 17341 26970 17570 26972
tri 17570 26970 17572 26972 sw
tri 17572 26970 17574 26972 ne
rect 17574 26970 17634 26972
rect 17341 26968 17572 26970
tri 17572 26968 17574 26970 sw
tri 17574 26968 17576 26970 ne
rect 17576 26968 17634 26970
rect 17341 26966 17574 26968
tri 17574 26966 17576 26968 sw
tri 17576 26966 17578 26968 ne
rect 17578 26966 17634 26968
rect 17341 26964 17576 26966
tri 17576 26964 17578 26966 sw
tri 17578 26964 17580 26966 ne
rect 17580 26964 17634 26966
tri 17512 26962 17514 26964 ne
rect 17514 26962 17578 26964
tri 17578 26962 17580 26964 sw
tri 17580 26962 17582 26964 ne
rect 17341 26960 17512 26962
tri 17512 26960 17514 26962 sw
tri 17514 26960 17516 26962 ne
rect 17516 26960 17580 26962
rect 17341 26958 17514 26960
tri 17514 26958 17516 26960 sw
tri 17516 26958 17518 26960 ne
rect 17518 26958 17580 26960
rect 17341 26956 17516 26958
tri 17516 26956 17518 26958 sw
tri 17518 26956 17520 26958 ne
rect 17520 26956 17580 26958
rect 17341 26954 17518 26956
tri 17518 26954 17520 26956 sw
tri 17520 26954 17522 26956 ne
rect 17522 26954 17580 26956
rect 17341 26952 17520 26954
tri 17520 26952 17522 26954 sw
tri 17522 26952 17524 26954 ne
rect 17524 26952 17580 26954
rect 17341 26950 17522 26952
tri 17522 26950 17524 26952 sw
tri 17524 26950 17526 26952 ne
rect 17526 26950 17580 26952
rect 17341 26948 17524 26950
tri 17524 26948 17526 26950 sw
tri 17526 26948 17528 26950 ne
rect 17528 26948 17580 26950
rect 17341 26946 17526 26948
tri 17526 26946 17528 26948 sw
tri 17528 26946 17530 26948 ne
rect 17530 26946 17580 26948
rect 17341 26944 17528 26946
tri 17528 26944 17530 26946 sw
tri 17530 26944 17532 26946 ne
rect 17532 26944 17580 26946
rect 17341 26942 17530 26944
tri 17530 26942 17532 26944 sw
tri 17532 26942 17534 26944 ne
rect 17534 26942 17580 26944
rect 17341 26940 17532 26942
tri 17532 26940 17534 26942 sw
tri 17534 26940 17536 26942 ne
rect 17536 26940 17580 26942
rect 17341 26938 17534 26940
tri 17534 26938 17536 26940 sw
tri 17536 26938 17538 26940 ne
rect 17538 26938 17580 26940
rect 17341 26936 17536 26938
tri 17536 26936 17538 26938 sw
tri 17538 26936 17540 26938 ne
rect 17540 26936 17580 26938
rect 17341 26934 17538 26936
tri 17538 26934 17540 26936 sw
tri 17540 26934 17542 26936 ne
rect 17542 26934 17580 26936
rect 17341 26932 17540 26934
tri 17540 26932 17542 26934 sw
tri 17542 26932 17544 26934 ne
rect 17341 26880 17542 26932
rect 222 26843 340 26880
rect 222 26841 300 26843
rect 222 26807 228 26841
rect 262 26809 300 26841
rect 334 26809 340 26843
rect 262 26807 340 26809
rect 222 26770 340 26807
rect 222 26768 300 26770
rect 222 26734 228 26768
rect 262 26736 300 26768
rect 334 26736 340 26770
rect 262 26734 340 26736
rect 222 26697 340 26734
rect 222 26695 300 26697
rect 222 26661 228 26695
rect 262 26663 300 26695
rect 334 26663 340 26697
rect 262 26661 340 26663
rect 222 26624 340 26661
rect 222 26622 300 26624
rect 222 26588 228 26622
rect 262 26590 300 26622
rect 334 26590 340 26624
rect 262 26588 340 26590
rect 222 26551 340 26588
rect 10665 26836 10721 26843
rect 10665 26784 10667 26836
rect 10719 26784 10721 26836
rect 10665 26772 10721 26784
rect 10665 26720 10667 26772
rect 10719 26720 10721 26772
rect 222 26549 300 26551
rect 222 26515 228 26549
rect 262 26517 300 26549
rect 334 26517 340 26551
rect 262 26515 340 26517
rect 222 26478 340 26515
rect 222 26476 300 26478
rect 222 26442 228 26476
rect 262 26444 300 26476
rect 334 26444 340 26478
rect 262 26442 340 26444
rect 222 26405 340 26442
rect 222 26403 300 26405
rect 222 26369 228 26403
rect 262 26371 300 26403
rect 334 26371 340 26405
rect 262 26369 340 26371
rect 222 26332 340 26369
rect 222 26330 300 26332
rect 222 26296 228 26330
rect 262 26298 300 26330
rect 334 26298 340 26332
rect 262 26296 340 26298
rect 222 26259 340 26296
rect 222 26257 300 26259
rect 222 26223 228 26257
rect 262 26225 300 26257
rect 334 26225 340 26259
rect 262 26223 340 26225
rect 222 26186 340 26223
rect 222 26184 300 26186
rect 222 26150 228 26184
rect 262 26152 300 26184
rect 334 26152 340 26186
rect 262 26150 340 26152
rect 222 26113 340 26150
rect 222 26111 300 26113
rect 222 26077 228 26111
rect 262 26079 300 26111
rect 334 26079 340 26113
rect 262 26077 340 26079
rect 222 26040 340 26077
rect 222 26038 300 26040
rect 222 26004 228 26038
rect 262 26006 300 26038
rect 334 26006 340 26040
rect 262 26004 340 26006
rect 222 25967 340 26004
rect 222 25965 300 25967
rect 222 25931 228 25965
rect 262 25933 300 25965
rect 334 25933 340 25967
rect 262 25931 340 25933
rect 222 25894 340 25931
rect 222 25892 300 25894
rect 222 25858 228 25892
rect 262 25860 300 25892
rect 334 25860 340 25894
rect 262 25858 340 25860
rect 222 25821 340 25858
rect 222 25819 300 25821
rect 222 25785 228 25819
rect 262 25787 300 25819
rect 334 25787 340 25821
rect 262 25785 340 25787
rect 222 25748 340 25785
rect 222 25746 300 25748
rect 222 25712 228 25746
rect 262 25714 300 25746
rect 334 25714 340 25748
rect 262 25712 340 25714
rect 222 25675 340 25712
rect 222 25673 300 25675
rect 222 25639 228 25673
rect 262 25641 300 25673
rect 334 25641 340 25675
rect 262 25639 340 25641
rect 222 25602 340 25639
rect 222 25600 300 25602
rect 222 25566 228 25600
rect 262 25568 300 25600
rect 334 25568 340 25602
rect 262 25566 340 25568
rect 222 25529 340 25566
rect 222 25527 300 25529
rect 222 25493 228 25527
rect 262 25495 300 25527
rect 334 25495 340 25529
rect 262 25493 340 25495
rect 222 25456 340 25493
rect 222 25454 300 25456
rect 222 25420 228 25454
rect 262 25422 300 25454
rect 334 25422 340 25456
rect 262 25420 340 25422
rect 222 25383 340 25420
rect 222 25381 300 25383
rect 222 25347 228 25381
rect 262 25349 300 25381
rect 334 25349 340 25383
rect 262 25347 340 25349
rect 222 25311 340 25347
rect 222 25308 300 25311
rect 222 25274 228 25308
rect 262 25277 300 25308
rect 334 25277 340 25311
rect 262 25274 340 25277
rect 222 25239 340 25274
rect 222 25235 300 25239
rect 222 25201 228 25235
rect 262 25205 300 25235
rect 334 25205 340 25239
rect 262 25201 340 25205
rect 222 25167 340 25201
rect 222 25162 300 25167
rect 222 25128 228 25162
rect 262 25133 300 25162
rect 334 25133 340 25167
rect 2876 26580 2928 26586
rect 2876 26516 2928 26528
rect 7009 26510 7015 26562
rect 7067 26510 7079 26562
rect 7131 26510 7143 26562
rect 7195 26510 7207 26562
rect 7259 26510 7271 26562
rect 7323 26510 7329 26562
rect 8593 26510 8599 26562
rect 8651 26510 8663 26562
rect 8715 26510 8727 26562
rect 8779 26510 8791 26562
rect 8843 26510 8855 26562
rect 8907 26510 8913 26562
rect 2876 25475 2928 26464
rect 5049 26458 5055 26510
rect 5107 26458 5119 26510
rect 5171 26458 5177 26510
rect 2876 25441 2882 25475
rect 2916 25441 2928 25475
rect 2876 25403 2928 25441
rect 2876 25369 2882 25403
rect 2916 25369 2928 25403
rect 262 25128 340 25133
rect 222 25095 340 25128
rect 660 25097 666 25149
rect 718 25097 730 25149
rect 782 25097 788 25149
rect 222 25089 300 25095
rect 222 25055 228 25089
rect 262 25061 300 25089
rect 334 25061 340 25095
rect 262 25055 340 25061
rect 222 25023 340 25055
rect 222 25016 300 25023
rect 222 24982 228 25016
rect 262 24989 300 25016
rect 334 24989 340 25023
rect 262 24982 340 24989
rect 222 24951 340 24982
rect 222 24943 300 24951
rect 222 24909 228 24943
rect 262 24917 300 24943
rect 334 24917 340 24951
rect 262 24909 340 24917
rect 222 24879 340 24909
rect 222 24870 300 24879
rect 222 24836 228 24870
rect 262 24845 300 24870
rect 334 24845 340 24879
rect 262 24836 340 24845
rect 222 24807 340 24836
rect 222 24797 300 24807
rect 222 24763 228 24797
rect 262 24773 300 24797
rect 334 24773 340 24807
rect 262 24763 340 24773
rect 222 24735 340 24763
rect 222 24724 300 24735
rect 222 24690 228 24724
rect 262 24701 300 24724
rect 334 24701 340 24735
rect 262 24690 340 24701
rect 222 24663 340 24690
rect 222 24651 300 24663
rect 222 24617 228 24651
rect 262 24629 300 24651
rect 334 24629 340 24663
rect 262 24617 340 24629
rect 222 24591 340 24617
rect 222 24578 300 24591
rect 222 24544 228 24578
rect 262 24557 300 24578
rect 334 24557 340 24591
rect 262 24544 340 24557
rect 222 24519 340 24544
rect 222 24505 300 24519
rect 222 24471 228 24505
rect 262 24485 300 24505
rect 334 24485 340 24519
rect 262 24471 340 24485
rect 222 24447 340 24471
rect 222 24432 300 24447
rect 222 24398 228 24432
rect 262 24413 300 24432
rect 334 24413 340 24447
rect 262 24398 340 24413
rect 222 24375 340 24398
rect 222 24359 300 24375
rect 222 24325 228 24359
rect 262 24341 300 24359
rect 334 24341 340 24375
rect 262 24325 340 24341
rect 222 24303 340 24325
rect 222 24286 300 24303
rect 222 24252 228 24286
rect 262 24269 300 24286
rect 334 24269 340 24303
rect 262 24252 340 24269
tri 1074 24252 1090 24268 se
rect 1090 24252 1142 24268
tri 1142 24252 1158 24268 sw
rect 222 24231 340 24252
tri 1065 24243 1074 24252 se
rect 1074 24246 1158 24252
rect 1074 24243 1090 24246
rect 222 24213 300 24231
rect 222 24179 228 24213
rect 262 24197 300 24213
rect 334 24197 340 24231
rect 689 24237 1090 24243
rect 1142 24243 1158 24246
tri 1158 24243 1167 24252 sw
rect 1142 24237 1664 24243
rect 689 24203 701 24237
rect 735 24203 778 24237
rect 812 24203 855 24237
rect 889 24203 932 24237
rect 966 24203 1009 24237
rect 1043 24203 1086 24237
rect 1142 24203 1162 24237
rect 1196 24203 1238 24237
rect 1272 24203 1314 24237
rect 1348 24203 1390 24237
rect 1424 24203 1466 24237
rect 1500 24203 1542 24237
rect 1576 24203 1618 24237
rect 1652 24203 1664 24237
rect 689 24197 1090 24203
rect 262 24179 340 24197
rect 1142 24197 1664 24203
rect 222 24159 340 24179
rect 222 24140 300 24159
rect 222 24106 228 24140
rect 262 24125 300 24140
rect 334 24125 340 24159
rect 262 24106 340 24125
rect 222 24087 340 24106
rect 222 24067 300 24087
rect 222 24033 228 24067
rect 262 24053 300 24067
rect 334 24053 340 24087
rect 262 24033 340 24053
rect 222 24015 340 24033
rect 222 23994 300 24015
rect 222 23960 228 23994
rect 262 23981 300 23994
rect 334 23981 340 24015
rect 262 23960 340 23981
rect 222 23943 340 23960
rect 222 23921 300 23943
rect 222 23887 228 23921
rect 262 23909 300 23921
rect 334 23909 340 23943
rect 603 24182 661 24188
rect 603 24148 615 24182
rect 649 24148 661 24182
rect 603 24110 661 24148
rect 1090 24182 1142 24194
rect 1090 24124 1142 24130
rect 603 24076 615 24110
rect 649 24076 661 24110
rect 1170 24122 1222 24128
rect 603 24038 661 24076
rect 689 24081 1170 24087
rect 1222 24081 1664 24087
rect 689 24047 701 24081
rect 735 24047 778 24081
rect 812 24047 855 24081
rect 889 24047 932 24081
rect 966 24047 1009 24081
rect 1043 24047 1086 24081
rect 1120 24047 1162 24081
rect 1222 24070 1238 24081
rect 1196 24058 1238 24070
rect 1222 24047 1238 24058
rect 1272 24047 1314 24081
rect 1348 24047 1390 24081
rect 1424 24047 1466 24081
rect 1500 24047 1542 24081
rect 1576 24047 1618 24081
rect 1652 24047 1664 24081
rect 689 24041 1170 24047
rect 603 24004 615 24038
rect 649 24004 661 24038
rect 1222 24041 1664 24047
rect 603 23966 661 24004
rect 603 23932 615 23966
rect 649 23932 661 23966
rect 603 23926 661 23932
rect 1090 23998 1142 24004
rect 1170 24000 1222 24006
rect 1090 23934 1142 23946
rect 262 23887 340 23909
rect 222 23871 340 23887
rect 689 23925 1090 23931
rect 1142 23925 1664 23931
rect 689 23891 701 23925
rect 735 23891 778 23925
rect 812 23891 855 23925
rect 889 23891 932 23925
rect 966 23891 1009 23925
rect 1043 23891 1086 23925
rect 1142 23891 1162 23925
rect 1196 23891 1238 23925
rect 1272 23891 1314 23925
rect 1348 23891 1390 23925
rect 1424 23891 1466 23925
rect 1500 23891 1542 23925
rect 1576 23891 1618 23925
rect 1652 23891 1664 23925
rect 689 23885 1090 23891
tri 1065 23876 1074 23885 ne
rect 1074 23882 1090 23885
rect 1142 23885 1664 23891
tri 2575 23885 2605 23915 se
rect 2605 23885 2657 23915
rect 1142 23882 1158 23885
rect 1074 23876 1158 23882
tri 1158 23876 1167 23885 nw
tri 2569 23879 2575 23885 se
rect 2575 23879 2657 23885
rect 222 23848 300 23871
rect 222 23814 228 23848
rect 262 23837 300 23848
rect 334 23837 340 23871
tri 1074 23860 1090 23876 ne
rect 1090 23860 1142 23876
tri 1142 23860 1158 23876 nw
rect 262 23814 340 23837
tri 1234 23830 1250 23846 se
rect 1250 23830 1302 23846
tri 1302 23830 1318 23846 sw
tri 1225 23821 1234 23830 se
rect 1234 23824 1318 23830
rect 1234 23821 1250 23824
rect 222 23799 340 23814
rect 222 23775 300 23799
rect 222 23741 228 23775
rect 262 23765 300 23775
rect 334 23765 340 23799
rect 689 23815 1250 23821
rect 1302 23821 1318 23824
tri 1318 23821 1327 23830 sw
rect 1302 23815 1664 23821
rect 262 23741 340 23765
rect 222 23727 340 23741
rect 222 23702 300 23727
rect 222 23668 228 23702
rect 262 23693 300 23702
rect 334 23693 340 23727
rect 262 23668 340 23693
rect 222 23655 340 23668
rect 222 23629 300 23655
rect 222 23595 228 23629
rect 262 23621 300 23629
rect 334 23621 340 23655
rect 262 23595 340 23621
rect 222 23583 340 23595
rect 222 23556 300 23583
rect 222 23522 228 23556
rect 262 23549 300 23556
rect 334 23549 340 23583
rect 262 23522 340 23549
rect 603 23779 661 23785
rect 603 23745 615 23779
rect 649 23745 661 23779
rect 689 23781 701 23815
rect 735 23781 778 23815
rect 812 23781 855 23815
rect 889 23781 932 23815
rect 966 23781 1009 23815
rect 1043 23781 1086 23815
rect 1120 23781 1162 23815
rect 1196 23781 1238 23815
rect 1302 23781 1314 23815
rect 1348 23781 1390 23815
rect 1424 23781 1466 23815
rect 1500 23781 1542 23815
rect 1576 23781 1618 23815
rect 1652 23781 1664 23815
rect 689 23775 1250 23781
rect 603 23707 661 23745
rect 603 23673 615 23707
rect 649 23673 661 23707
rect 1302 23775 1664 23781
rect 2569 23816 2657 23879
rect 2569 23813 2642 23816
tri 2642 23813 2645 23816 nw
rect 1250 23760 1302 23772
rect 1250 23702 1302 23708
rect 2569 23717 2620 23813
tri 2620 23791 2642 23813 nw
tri 2854 23791 2876 23813 se
rect 2876 23791 2928 25369
rect 4502 24216 4508 24268
rect 4560 24216 4572 24268
rect 4624 24216 4636 24268
rect 4688 24216 4700 24268
rect 4752 24216 4764 24268
rect 4816 24216 4822 24268
rect 5326 24216 5332 24268
rect 5384 24216 5396 24268
rect 5448 24216 5460 24268
rect 5512 24216 5524 24268
rect 5576 24216 5588 24268
rect 5640 24216 5646 24268
rect 6150 24216 6156 24268
rect 6208 24216 6220 24268
rect 6272 24216 6284 24268
rect 6336 24216 6348 24268
rect 6400 24216 6412 24268
rect 6464 24216 6470 24268
rect 6974 24216 6980 24268
rect 7032 24216 7044 24268
rect 7096 24216 7108 24268
rect 7160 24216 7172 24268
rect 7224 24216 7236 24268
rect 7288 24216 7294 24268
rect 7798 24216 7804 24268
rect 7856 24216 7868 24268
rect 7920 24216 7932 24268
rect 7984 24216 7996 24268
rect 8048 24216 8060 24268
rect 8112 24216 8118 24268
rect 8622 24216 8628 24268
rect 8680 24216 8692 24268
rect 8744 24216 8756 24268
rect 8808 24216 8820 24268
rect 8872 24216 8884 24268
rect 8936 24216 8942 24268
rect 9460 24216 9466 24268
rect 9518 24216 9530 24268
rect 9582 24216 9594 24268
rect 9646 24216 9658 24268
rect 9710 24216 9722 24268
rect 9774 24216 9780 24268
rect 10270 24216 10276 24268
rect 10328 24216 10340 24268
rect 10392 24216 10404 24268
rect 10456 24216 10468 24268
rect 10520 24216 10532 24268
rect 10584 24216 10590 24268
rect 10665 24149 10721 26720
rect 10665 24097 10667 24149
rect 10719 24097 10721 24149
rect 10665 24085 10721 24097
rect 10665 24033 10667 24085
rect 10719 24033 10721 24085
rect 10665 24027 10721 24033
rect 10977 26552 11033 26559
rect 10977 26500 10979 26552
rect 11031 26500 11033 26552
rect 11196 26510 11202 26562
rect 11254 26510 11266 26562
rect 11318 26510 11330 26562
rect 11382 26510 11394 26562
rect 11446 26510 11452 26562
rect 12716 26510 12722 26562
rect 12774 26510 12786 26562
rect 12838 26510 12850 26562
rect 12902 26510 12914 26562
rect 12966 26510 12978 26562
rect 13030 26510 13036 26562
rect 15254 26510 15260 26562
rect 15312 26510 15324 26562
rect 15376 26510 15388 26562
rect 15440 26510 15452 26562
rect 15504 26510 15516 26562
rect 15568 26510 15574 26562
rect 16838 26510 16844 26562
rect 16896 26510 16908 26562
rect 16960 26510 16972 26562
rect 17024 26510 17036 26562
rect 17088 26510 17100 26562
rect 17152 26510 17158 26562
rect 10977 26488 11033 26500
rect 10977 26436 10979 26488
rect 11031 26436 11033 26488
rect 10977 24149 11033 26436
rect 11080 24216 11086 24268
rect 11138 24216 11150 24268
rect 11202 24216 11214 24268
rect 11266 24216 11278 24268
rect 11330 24216 11342 24268
rect 11394 24216 11400 24268
rect 11918 24216 11924 24268
rect 11976 24216 11988 24268
rect 12040 24216 12052 24268
rect 12104 24216 12116 24268
rect 12168 24216 12180 24268
rect 12232 24216 12238 24268
rect 12742 24216 12748 24268
rect 12800 24216 12812 24268
rect 12864 24216 12876 24268
rect 12928 24216 12940 24268
rect 12992 24216 13004 24268
rect 13056 24216 13062 24268
rect 13566 24216 13572 24268
rect 13624 24216 13636 24268
rect 13688 24216 13700 24268
rect 13752 24216 13764 24268
rect 13816 24216 13828 24268
rect 13880 24216 13886 24268
rect 14390 24216 14396 24268
rect 14448 24216 14460 24268
rect 14512 24216 14524 24268
rect 14576 24216 14588 24268
rect 14640 24216 14652 24268
rect 14704 24216 14710 24268
rect 15214 24216 15220 24268
rect 15272 24216 15284 24268
rect 15336 24216 15348 24268
rect 15400 24216 15412 24268
rect 15464 24216 15476 24268
rect 15528 24216 15534 24268
rect 16038 24216 16044 24268
rect 16096 24216 16108 24268
rect 16160 24216 16172 24268
rect 16224 24216 16236 24268
rect 16288 24216 16300 24268
rect 16352 24216 16358 24268
rect 16862 24216 16868 24268
rect 16920 24216 16932 24268
rect 16984 24216 16996 24268
rect 17048 24216 17060 24268
rect 17112 24216 17124 24268
rect 17176 24216 17182 24268
rect 10977 24097 10979 24149
rect 11031 24097 11033 24149
rect 10977 24085 11033 24097
rect 10977 24033 10979 24085
rect 11031 24033 11033 24085
rect 10977 24027 11033 24033
rect 4477 23877 4861 23973
rect 4983 23892 5178 23976
rect 5299 23877 5683 23973
rect 5807 23892 6002 23976
rect 6123 23877 6507 23973
rect 6631 23892 6826 23976
rect 6947 23877 7331 23973
rect 7455 23892 7650 23976
rect 7771 23877 8155 23973
rect 8279 23892 8474 23976
rect 8595 23877 8979 23973
rect 9103 23892 9298 23976
rect 9419 23877 9803 23973
rect 9927 23892 10122 23976
rect 10243 23877 10627 23973
rect 10751 23892 10946 23976
rect 11067 23877 11451 23973
rect 11575 23892 11770 23976
rect 11891 23877 12275 23973
rect 12399 23892 12594 23976
rect 12715 23877 13099 23973
rect 13223 23892 13418 23976
rect 13539 23877 13923 23973
rect 14047 23892 14242 23976
rect 14363 23877 14747 23973
rect 15187 23877 15571 23973
rect 16011 23877 16395 23973
rect 16835 23877 17219 23973
rect 17490 23874 17542 26880
rect 17544 26879 17580 26934
rect 17543 23875 17581 26879
tri 2851 23788 2854 23791 se
rect 2854 23788 2928 23791
rect 17341 23822 17542 23874
rect 17341 23820 17540 23822
tri 17540 23820 17542 23822 nw
tri 17542 23820 17544 23822 se
rect 17544 23820 17580 23875
rect 17341 23818 17538 23820
tri 17538 23818 17540 23820 nw
tri 17540 23818 17542 23820 se
rect 17542 23818 17580 23820
rect 17341 23816 17536 23818
tri 17536 23816 17538 23818 nw
tri 17538 23816 17540 23818 se
rect 17540 23816 17580 23818
rect 17341 23814 17534 23816
tri 17534 23814 17536 23816 nw
tri 17536 23814 17538 23816 se
rect 17538 23814 17580 23816
rect 17341 23812 17532 23814
tri 17532 23812 17534 23814 nw
tri 17534 23812 17536 23814 se
rect 17536 23812 17580 23814
rect 17341 23810 17530 23812
tri 17530 23810 17532 23812 nw
tri 17532 23810 17534 23812 se
rect 17534 23810 17580 23812
rect 17341 23808 17528 23810
tri 17528 23808 17530 23810 nw
tri 17530 23808 17532 23810 se
rect 17532 23808 17580 23810
rect 17341 23806 17526 23808
tri 17526 23806 17528 23808 nw
tri 17528 23806 17530 23808 se
rect 17530 23806 17580 23808
rect 17341 23804 17524 23806
tri 17524 23804 17526 23806 nw
tri 17526 23804 17528 23806 se
rect 17528 23804 17580 23806
rect 17341 23802 17522 23804
tri 17522 23802 17524 23804 nw
tri 17524 23802 17526 23804 se
rect 17526 23802 17580 23804
rect 17341 23800 17520 23802
tri 17520 23800 17522 23802 nw
tri 17522 23800 17524 23802 se
rect 17524 23800 17580 23802
rect 17341 23798 17518 23800
tri 17518 23798 17520 23800 nw
tri 17520 23798 17522 23800 se
rect 17522 23798 17580 23800
rect 17341 23796 17516 23798
tri 17516 23796 17518 23798 nw
tri 17518 23796 17520 23798 se
rect 17520 23796 17580 23798
rect 17341 23794 17514 23796
tri 17514 23794 17516 23796 nw
tri 17516 23794 17518 23796 se
rect 17518 23794 17580 23796
rect 17341 23792 17512 23794
tri 17512 23792 17514 23794 nw
tri 17514 23792 17516 23794 se
rect 17516 23792 17580 23794
tri 17512 23790 17514 23792 se
rect 17514 23790 17578 23792
tri 17578 23790 17580 23792 nw
tri 17580 23790 17582 23792 se
rect 17582 23790 17634 26964
rect 17341 23788 17576 23790
tri 17576 23788 17578 23790 nw
tri 17578 23788 17580 23790 se
rect 17580 23788 17634 23790
rect 2657 23736 2663 23788
rect 2715 23736 2727 23788
rect 2779 23736 2785 23788
rect 2787 23787 2823 23788
rect 2786 23737 2824 23787
rect 2787 23736 2823 23737
rect 2825 23736 2928 23788
rect 4398 23779 4649 23788
rect 4651 23787 4687 23788
rect 4398 23745 4410 23779
rect 4444 23745 4482 23779
rect 4516 23745 4649 23779
rect 4398 23736 4649 23745
rect 4650 23737 4688 23787
rect 4689 23779 5061 23788
rect 5063 23787 5099 23788
rect 4689 23745 4822 23779
rect 4856 23745 4894 23779
rect 4928 23745 5061 23779
rect 4651 23736 4687 23737
rect 4689 23736 5061 23745
rect 5062 23737 5100 23787
rect 5101 23779 5473 23788
rect 5475 23787 5511 23788
rect 5101 23745 5234 23779
rect 5268 23745 5306 23779
rect 5340 23745 5473 23779
rect 5063 23736 5099 23737
rect 5101 23736 5473 23745
rect 5474 23737 5512 23787
rect 5513 23779 5885 23788
rect 5887 23787 5923 23788
rect 5513 23745 5646 23779
rect 5680 23745 5718 23779
rect 5752 23745 5885 23779
rect 5475 23736 5511 23737
rect 5513 23736 5885 23745
rect 5886 23737 5924 23787
rect 5925 23779 6297 23788
rect 6299 23787 6335 23788
rect 5925 23745 6058 23779
rect 6092 23745 6130 23779
rect 6164 23745 6297 23779
rect 5887 23736 5923 23737
rect 5925 23736 6297 23745
rect 6298 23737 6336 23787
rect 6337 23779 6709 23788
rect 6337 23745 6470 23779
rect 6504 23745 6542 23779
rect 6576 23745 6709 23779
rect 6299 23736 6335 23737
rect 6337 23736 6709 23745
rect 6710 23737 6711 23787
rect 6747 23737 6748 23787
rect 6749 23779 6998 23788
rect 6749 23745 6882 23779
rect 6916 23745 6954 23779
rect 6988 23745 6998 23779
rect 6749 23736 6998 23745
rect 7050 23736 7062 23788
rect 7114 23736 7121 23788
rect 7123 23787 7159 23788
rect 7122 23737 7160 23787
rect 7161 23779 7533 23788
rect 7535 23787 7571 23788
rect 7161 23745 7294 23779
rect 7328 23745 7366 23779
rect 7400 23745 7533 23779
rect 7123 23736 7159 23737
rect 7161 23736 7533 23745
rect 7534 23737 7572 23787
rect 7573 23779 7850 23788
rect 7852 23787 7888 23788
rect 7573 23745 7706 23779
rect 7740 23745 7778 23779
rect 7812 23745 7850 23779
rect 7535 23736 7571 23737
rect 7573 23736 7850 23745
rect 7851 23737 7889 23787
rect 7852 23736 7888 23737
rect 7890 23736 7904 23788
rect 7956 23736 7968 23788
rect 8020 23736 8039 23788
rect 8041 23787 8077 23788
rect 8040 23737 8078 23787
rect 8079 23779 8357 23788
rect 8359 23787 8395 23788
rect 8079 23745 8118 23779
rect 8152 23745 8190 23779
rect 8224 23745 8357 23779
rect 8041 23736 8077 23737
rect 8079 23736 8357 23745
rect 8358 23737 8396 23787
rect 8397 23779 8769 23788
rect 8397 23745 8530 23779
rect 8564 23745 8602 23779
rect 8636 23745 8769 23779
rect 8359 23736 8395 23737
rect 8397 23736 8769 23745
rect 8770 23737 8771 23787
rect 8807 23737 8808 23787
rect 8809 23779 9181 23788
rect 9183 23787 9219 23788
rect 8809 23745 8942 23779
rect 8976 23745 9014 23779
rect 9048 23745 9181 23779
rect 8809 23736 9181 23745
rect 9182 23737 9220 23787
rect 9221 23779 9593 23788
rect 9595 23787 9631 23788
rect 9221 23745 9354 23779
rect 9388 23745 9426 23779
rect 9460 23745 9593 23779
rect 9183 23736 9219 23737
rect 9221 23736 9593 23745
rect 9594 23737 9632 23787
rect 9633 23779 10005 23788
rect 10007 23787 10043 23788
rect 9633 23745 9766 23779
rect 9800 23745 9838 23779
rect 9872 23745 10005 23779
rect 9595 23736 9631 23737
rect 9633 23736 10005 23745
rect 10006 23737 10044 23787
rect 10045 23779 10417 23788
rect 10419 23787 10455 23788
rect 10045 23745 10178 23779
rect 10212 23745 10250 23779
rect 10284 23745 10417 23779
rect 10007 23736 10043 23737
rect 10045 23736 10417 23745
rect 10418 23737 10456 23787
rect 10457 23779 10829 23788
rect 10831 23787 10867 23788
rect 10457 23745 10590 23779
rect 10624 23745 10662 23779
rect 10696 23745 10829 23779
rect 10419 23736 10455 23737
rect 10457 23736 10829 23745
rect 10830 23737 10868 23787
rect 10869 23779 11120 23788
rect 10869 23745 11002 23779
rect 11036 23745 11074 23779
rect 11108 23745 11120 23779
rect 10831 23736 10867 23737
rect 10869 23736 11120 23745
rect 11232 23779 11362 23788
rect 11364 23787 11400 23788
rect 11232 23745 11244 23779
rect 11278 23745 11316 23779
rect 11350 23745 11362 23779
rect 11232 23736 11362 23745
rect 11363 23737 11401 23787
rect 11402 23779 11532 23788
rect 11402 23745 11414 23779
rect 11448 23745 11486 23779
rect 11520 23745 11532 23779
rect 11364 23736 11400 23737
rect 11402 23736 11532 23745
rect 11533 23737 11534 23787
rect 11570 23737 11571 23787
rect 11572 23779 11774 23788
rect 11572 23745 11620 23779
rect 11654 23745 11692 23779
rect 11726 23745 11774 23779
rect 11572 23736 11774 23745
rect 11775 23737 11776 23787
rect 11812 23737 11813 23787
rect 11814 23779 11944 23788
rect 11946 23787 11982 23788
rect 11814 23745 11826 23779
rect 11860 23745 11898 23779
rect 11932 23745 11944 23779
rect 11814 23736 11944 23745
rect 11945 23737 11983 23787
rect 11984 23779 12186 23788
rect 12188 23787 12224 23788
rect 11984 23745 12032 23779
rect 12066 23745 12104 23779
rect 12138 23745 12186 23779
rect 11946 23736 11982 23737
rect 11984 23736 12186 23745
rect 12187 23737 12225 23787
rect 12226 23779 12356 23788
rect 12226 23745 12238 23779
rect 12272 23745 12310 23779
rect 12344 23745 12356 23779
rect 12188 23736 12224 23737
rect 12226 23736 12356 23745
rect 12357 23737 12358 23787
rect 12394 23737 12395 23787
rect 12396 23779 12598 23788
rect 12396 23745 12444 23779
rect 12478 23745 12516 23779
rect 12550 23745 12598 23779
rect 12396 23736 12598 23745
rect 12599 23737 12600 23787
rect 12636 23737 12637 23787
rect 12638 23779 12768 23788
rect 12770 23787 12806 23788
rect 12638 23745 12650 23779
rect 12684 23745 12722 23779
rect 12756 23745 12768 23779
rect 12638 23736 12768 23745
rect 12769 23737 12807 23787
rect 12808 23779 13010 23788
rect 13012 23787 13048 23788
rect 12808 23745 12856 23779
rect 12890 23745 12928 23779
rect 12962 23745 13010 23779
rect 12770 23736 12806 23737
rect 12808 23736 13010 23745
rect 13011 23737 13049 23787
rect 13050 23779 13180 23788
rect 13050 23745 13062 23779
rect 13096 23745 13134 23779
rect 13168 23745 13180 23779
rect 13012 23736 13048 23737
rect 13050 23736 13180 23745
rect 13181 23737 13182 23787
rect 13218 23737 13219 23787
rect 13220 23779 13422 23788
rect 13220 23745 13268 23779
rect 13302 23745 13340 23779
rect 13374 23745 13422 23779
rect 13220 23736 13422 23745
rect 13423 23737 13424 23787
rect 13460 23737 13461 23787
rect 13462 23779 13592 23788
rect 13594 23787 13630 23788
rect 13462 23745 13474 23779
rect 13508 23745 13546 23779
rect 13580 23745 13592 23779
rect 13462 23736 13592 23745
rect 13593 23737 13631 23787
rect 13632 23779 13834 23788
rect 13632 23745 13680 23779
rect 13714 23745 13752 23779
rect 13786 23745 13834 23779
rect 13594 23736 13630 23737
rect 13632 23736 13834 23745
rect 13835 23737 13836 23787
rect 13872 23737 13873 23787
rect 13874 23779 14004 23788
rect 14006 23787 14042 23788
rect 13874 23745 13886 23779
rect 13920 23745 13958 23779
rect 13992 23745 14004 23779
rect 13874 23736 14004 23745
rect 14005 23737 14043 23787
rect 14044 23779 14246 23788
rect 14248 23787 14284 23788
rect 14044 23745 14092 23779
rect 14126 23745 14164 23779
rect 14198 23745 14246 23779
rect 14006 23736 14042 23737
rect 14044 23736 14246 23745
rect 14247 23737 14285 23787
rect 14286 23779 14416 23788
rect 14286 23745 14298 23779
rect 14332 23745 14370 23779
rect 14404 23745 14416 23779
rect 14248 23736 14284 23737
rect 14286 23736 14416 23745
rect 14417 23737 14418 23787
rect 14454 23737 14455 23787
rect 14456 23779 14586 23788
rect 17341 23786 17574 23788
tri 17574 23786 17576 23788 nw
tri 17576 23786 17578 23788 se
rect 17578 23786 17634 23788
rect 17341 23785 17573 23786
tri 17573 23785 17574 23786 nw
tri 17575 23785 17576 23786 se
rect 17576 23785 17634 23786
rect 14456 23745 14468 23779
rect 14502 23745 14540 23779
rect 14574 23745 14586 23779
rect 14456 23736 14586 23745
rect 14644 23779 14947 23785
rect 14644 23745 14656 23779
rect 14690 23745 14728 23779
rect 14762 23745 14947 23779
rect 14644 23739 14947 23745
rect 14948 23740 14949 23784
rect 14985 23740 14986 23784
rect 14987 23779 15173 23785
rect 15225 23779 15238 23785
rect 14987 23745 15124 23779
rect 15158 23745 15173 23779
rect 15230 23745 15238 23779
rect 14987 23739 15173 23745
tri 15161 23736 15164 23739 ne
rect 15164 23736 15173 23739
tri 2851 23733 2854 23736 ne
rect 2854 23733 2928 23736
tri 15164 23733 15167 23736 ne
rect 15167 23733 15173 23736
rect 15225 23733 15238 23745
rect 15290 23733 15296 23785
rect 15336 23733 15342 23785
rect 15394 23733 15407 23785
rect 15459 23779 15895 23785
rect 15897 23784 15933 23785
rect 15459 23745 15536 23779
rect 15570 23745 15608 23779
rect 15642 23745 15895 23779
rect 15459 23739 15895 23745
rect 15896 23740 15934 23784
rect 15935 23779 16296 23785
rect 16298 23784 16334 23785
rect 15935 23745 15948 23779
rect 15982 23745 16020 23779
rect 16054 23745 16296 23779
rect 15897 23739 15933 23740
rect 15935 23739 16296 23745
rect 16297 23740 16335 23784
rect 16336 23779 16719 23785
rect 16721 23784 16757 23785
rect 16336 23745 16360 23779
rect 16394 23745 16432 23779
rect 16466 23745 16719 23779
rect 16298 23739 16334 23740
rect 16336 23739 16719 23745
rect 16720 23740 16758 23784
rect 16759 23779 16890 23785
rect 16892 23784 16928 23785
rect 16759 23745 16772 23779
rect 16806 23745 16844 23779
rect 16878 23745 16890 23779
rect 16721 23739 16757 23740
rect 16759 23739 16890 23745
rect 16891 23740 16929 23784
rect 16930 23779 17233 23785
rect 16930 23745 17115 23779
rect 17149 23745 17187 23779
rect 17221 23745 17233 23779
rect 16892 23739 16928 23740
rect 16930 23739 17233 23745
rect 17341 23784 17572 23785
tri 17572 23784 17573 23785 nw
tri 17574 23784 17575 23785 se
rect 17575 23784 17634 23785
rect 17341 23782 17570 23784
tri 17570 23782 17572 23784 nw
tri 17572 23782 17574 23784 se
rect 17574 23782 17634 23784
rect 17341 23780 17568 23782
tri 17568 23780 17570 23782 nw
tri 17570 23780 17572 23782 se
rect 17572 23780 17634 23782
rect 17341 23778 17566 23780
tri 17566 23778 17568 23780 nw
tri 17568 23778 17570 23780 se
rect 17570 23778 17634 23780
rect 17341 23776 17564 23778
tri 17564 23776 17566 23778 nw
tri 17566 23776 17568 23778 se
rect 17568 23776 17634 23778
rect 17341 23774 17562 23776
tri 17562 23774 17564 23776 nw
tri 17564 23774 17566 23776 se
rect 17566 23774 17634 23776
rect 17341 23772 17560 23774
tri 17560 23772 17562 23774 nw
tri 17562 23772 17564 23774 se
rect 17564 23772 17634 23774
rect 17341 23770 17558 23772
tri 17558 23770 17560 23772 nw
tri 17560 23770 17562 23772 se
rect 17562 23770 17634 23772
rect 17341 23768 17556 23770
tri 17556 23768 17558 23770 nw
tri 17558 23768 17560 23770 se
rect 17560 23768 17634 23770
rect 17341 23766 17554 23768
tri 17554 23766 17556 23768 nw
tri 17556 23766 17558 23768 se
rect 17558 23766 17634 23768
rect 17341 23764 17552 23766
tri 17552 23764 17554 23766 nw
tri 17554 23764 17556 23766 se
rect 17556 23764 17634 23766
rect 17341 23762 17550 23764
tri 17550 23762 17552 23764 nw
tri 17552 23762 17554 23764 se
rect 17554 23762 17634 23764
tri 17550 23760 17552 23762 se
rect 17552 23760 17634 23762
rect 15459 23736 15468 23739
tri 15468 23736 15471 23739 nw
tri 16934 23736 16937 23739 ne
rect 16937 23736 17084 23739
rect 15459 23733 15465 23736
tri 15465 23733 15468 23736 nw
tri 16937 23733 16940 23736 ne
rect 16940 23733 17084 23736
tri 2620 23717 2636 23733 sw
tri 2854 23717 2870 23733 ne
rect 2870 23717 2928 23733
tri 16940 23717 16956 23733 ne
rect 2569 23711 2636 23717
tri 2636 23711 2642 23717 sw
tri 2870 23711 2876 23717 ne
rect 2569 23706 2642 23711
tri 2642 23706 2647 23711 sw
rect 603 23635 661 23673
rect 1330 23700 1382 23706
rect 603 23601 615 23635
rect 649 23601 661 23635
rect 689 23659 1330 23665
rect 2569 23699 2647 23706
tri 2647 23699 2654 23706 sw
rect 1382 23659 1664 23665
rect 689 23625 701 23659
rect 735 23625 778 23659
rect 812 23625 855 23659
rect 889 23625 932 23659
rect 966 23625 1009 23659
rect 1043 23625 1086 23659
rect 1120 23625 1162 23659
rect 1196 23625 1238 23659
rect 1272 23625 1314 23659
rect 1382 23648 1390 23659
rect 1348 23636 1390 23648
rect 1382 23625 1390 23636
rect 1424 23625 1466 23659
rect 1500 23625 1542 23659
rect 1576 23625 1618 23659
rect 1652 23625 1664 23659
rect 689 23619 1330 23625
rect 603 23563 661 23601
rect 1382 23619 1664 23625
rect 603 23529 615 23563
rect 649 23529 661 23563
rect 603 23523 661 23529
rect 1250 23576 1302 23582
rect 1330 23578 1382 23584
rect 2569 23585 2654 23699
rect 2569 23578 2647 23585
tri 2647 23578 2654 23585 nw
rect 222 23511 340 23522
rect 222 23483 300 23511
rect 222 23449 228 23483
rect 262 23477 300 23483
rect 334 23477 340 23511
rect 1250 23512 1302 23524
rect 262 23449 340 23477
rect 689 23503 1250 23509
rect 2569 23573 2642 23578
tri 2642 23573 2647 23578 nw
rect 2569 23572 2641 23573
tri 2641 23572 2642 23573 nw
tri 2875 23572 2876 23573 se
rect 2876 23572 2928 23717
rect 4217 23656 4223 23708
rect 4275 23656 4287 23708
rect 4339 23699 15107 23708
rect 4339 23665 4410 23699
rect 4444 23665 4482 23699
rect 4516 23665 11244 23699
rect 11278 23665 11316 23699
rect 11350 23665 12032 23699
rect 12066 23665 12104 23699
rect 12138 23665 12856 23699
rect 12890 23665 12928 23699
rect 12962 23665 13680 23699
rect 13714 23665 13752 23699
rect 13786 23665 14468 23699
rect 14502 23665 14540 23699
rect 14574 23665 15107 23699
rect 16828 23695 16880 23701
rect 4339 23656 15107 23665
tri 16794 23661 16828 23695 se
rect 4217 23576 4223 23628
rect 4275 23576 4287 23628
rect 4339 23622 14998 23628
rect 4339 23588 11002 23622
rect 11036 23588 11074 23622
rect 11108 23588 11620 23622
rect 11654 23588 11692 23622
rect 11726 23588 12444 23622
rect 12478 23588 12516 23622
rect 12550 23588 13268 23622
rect 13302 23588 13340 23622
rect 13374 23588 14092 23622
rect 14126 23588 14164 23622
rect 14198 23588 14998 23622
rect 15210 23609 15216 23661
rect 15268 23609 15285 23661
rect 15337 23609 15353 23661
rect 15405 23643 16828 23661
rect 15405 23630 16880 23643
rect 15405 23609 16828 23630
rect 4339 23576 14998 23588
tri 16794 23576 16827 23609 ne
rect 16827 23578 16828 23609
rect 16827 23576 16880 23578
tri 16827 23575 16828 23576 ne
rect 16828 23572 16880 23576
rect 16956 23665 17084 23733
tri 17084 23717 17106 23739 nw
rect 16957 23663 17083 23664
rect 16956 23627 17084 23663
tri 17328 23627 17341 23640 se
rect 17341 23627 17634 23760
rect 16957 23626 17083 23627
tri 17327 23626 17328 23627 se
rect 17328 23626 17634 23627
tri 17326 23625 17327 23626 se
rect 17327 23625 17634 23626
rect 16956 23613 17084 23625
rect 2569 23561 2630 23572
tri 2630 23561 2641 23572 nw
tri 2864 23561 2875 23572 se
rect 2875 23561 2928 23572
rect 16956 23561 16962 23613
rect 17014 23561 17026 23613
rect 17078 23561 17084 23613
tri 17262 23561 17326 23625 se
rect 17326 23561 17634 23625
rect 17647 26035 18349 26041
rect 17647 24767 17652 26035
rect 18344 24767 18349 26035
rect 17647 24754 18349 24767
rect 17647 24702 17652 24754
rect 17704 24702 17716 24754
rect 17768 24702 17780 24754
rect 17832 24702 17844 24754
rect 17896 24702 17908 24754
rect 17960 24702 17972 24754
rect 18024 24702 18036 24754
rect 18088 24702 18100 24754
rect 18152 24702 18164 24754
rect 18216 24702 18228 24754
rect 18280 24702 18292 24754
rect 18344 24702 18349 24754
rect 17647 24689 18349 24702
rect 17647 24637 17652 24689
rect 17704 24637 17716 24689
rect 17768 24637 17780 24689
rect 17832 24637 17844 24689
rect 17896 24637 17908 24689
rect 17960 24637 17972 24689
rect 18024 24637 18036 24689
rect 18088 24637 18100 24689
rect 18152 24637 18164 24689
rect 18216 24637 18228 24689
rect 18280 24637 18292 24689
rect 18344 24637 18349 24689
rect 17647 24624 18349 24637
rect 17647 24572 17652 24624
rect 17704 24572 17716 24624
rect 17768 24572 17780 24624
rect 17832 24572 17844 24624
rect 17896 24572 17908 24624
rect 17960 24572 17972 24624
rect 18024 24572 18036 24624
rect 18088 24572 18100 24624
rect 18152 24572 18164 24624
rect 18216 24572 18228 24624
rect 18280 24572 18292 24624
rect 18344 24572 18349 24624
rect 17647 24559 18349 24572
rect 17647 24507 17652 24559
rect 17704 24507 17716 24559
rect 17768 24507 17780 24559
rect 17832 24507 17844 24559
rect 17896 24507 17908 24559
rect 17960 24507 17972 24559
rect 18024 24507 18036 24559
rect 18088 24507 18100 24559
rect 18152 24507 18164 24559
rect 18216 24507 18228 24559
rect 18280 24507 18292 24559
rect 18344 24507 18349 24559
rect 17647 24494 18349 24507
rect 17647 24442 17652 24494
rect 17704 24442 17716 24494
rect 17768 24442 17780 24494
rect 17832 24442 17844 24494
rect 17896 24442 17908 24494
rect 17960 24442 17972 24494
rect 18024 24442 18036 24494
rect 18088 24442 18100 24494
rect 18152 24442 18164 24494
rect 18216 24442 18228 24494
rect 18280 24442 18292 24494
rect 18344 24442 18349 24494
rect 17647 24429 18349 24442
rect 17647 24377 17652 24429
rect 17704 24377 17716 24429
rect 17768 24377 17780 24429
rect 17832 24377 17844 24429
rect 17896 24377 17908 24429
rect 17960 24377 17972 24429
rect 18024 24377 18036 24429
rect 18088 24377 18100 24429
rect 18152 24377 18164 24429
rect 18216 24377 18228 24429
rect 18280 24377 18292 24429
rect 18344 24377 18349 24429
rect 17647 24364 18349 24377
rect 17647 24312 17652 24364
rect 17704 24312 17716 24364
rect 17768 24312 17780 24364
rect 17832 24312 17844 24364
rect 17896 24312 17908 24364
rect 17960 24312 17972 24364
rect 18024 24312 18036 24364
rect 18088 24312 18100 24364
rect 18152 24312 18164 24364
rect 18216 24312 18228 24364
rect 18280 24312 18292 24364
rect 18344 24312 18349 24364
rect 17647 24299 18349 24312
rect 17647 24247 17652 24299
rect 17704 24247 17716 24299
rect 17768 24247 17780 24299
rect 17832 24247 17844 24299
rect 17896 24247 17908 24299
rect 17960 24247 17972 24299
rect 18024 24247 18036 24299
rect 18088 24247 18100 24299
rect 18152 24247 18164 24299
rect 18216 24247 18228 24299
rect 18280 24247 18292 24299
rect 18344 24247 18349 24299
rect 17647 24234 18349 24247
rect 17647 24182 17652 24234
rect 17704 24182 17716 24234
rect 17768 24182 17780 24234
rect 17832 24182 17844 24234
rect 17896 24182 17908 24234
rect 17960 24182 17972 24234
rect 18024 24182 18036 24234
rect 18088 24182 18100 24234
rect 18152 24182 18164 24234
rect 18216 24182 18228 24234
rect 18280 24182 18292 24234
rect 18344 24182 18349 24234
rect 17647 24169 18349 24182
rect 17647 24117 17652 24169
rect 17704 24117 17716 24169
rect 17768 24117 17780 24169
rect 17832 24117 17844 24169
rect 17896 24117 17908 24169
rect 17960 24117 17972 24169
rect 18024 24117 18036 24169
rect 18088 24117 18100 24169
rect 18152 24117 18164 24169
rect 18216 24117 18228 24169
rect 18280 24117 18292 24169
rect 18344 24117 18349 24169
rect 17647 24104 18349 24117
rect 17647 24052 17652 24104
rect 17704 24052 17716 24104
rect 17768 24052 17780 24104
rect 17832 24052 17844 24104
rect 17896 24052 17908 24104
rect 17960 24052 17972 24104
rect 18024 24052 18036 24104
rect 18088 24052 18100 24104
rect 18152 24052 18164 24104
rect 18216 24052 18228 24104
rect 18280 24052 18292 24104
rect 18344 24052 18349 24104
rect 17647 24039 18349 24052
rect 17647 23987 17652 24039
rect 17704 23987 17716 24039
rect 17768 23987 17780 24039
rect 17832 23987 17844 24039
rect 17896 23987 17908 24039
rect 17960 23987 17972 24039
rect 18024 23987 18036 24039
rect 18088 23987 18100 24039
rect 18152 23987 18164 24039
rect 18216 23987 18228 24039
rect 18280 23987 18292 24039
rect 18344 23987 18349 24039
rect 17647 23974 18349 23987
rect 17647 23922 17652 23974
rect 17704 23922 17716 23974
rect 17768 23922 17780 23974
rect 17832 23922 17844 23974
rect 17896 23922 17908 23974
rect 17960 23922 17972 23974
rect 18024 23922 18036 23974
rect 18088 23922 18100 23974
rect 18152 23922 18164 23974
rect 18216 23922 18228 23974
rect 18280 23922 18292 23974
rect 18344 23922 18349 23974
rect 17647 23909 18349 23922
rect 17647 23857 17652 23909
rect 17704 23857 17716 23909
rect 17768 23857 17780 23909
rect 17832 23857 17844 23909
rect 17896 23857 17908 23909
rect 17960 23857 17972 23909
rect 18024 23857 18036 23909
rect 18088 23857 18100 23909
rect 18152 23857 18164 23909
rect 18216 23857 18228 23909
rect 18280 23857 18292 23909
rect 18344 23857 18349 23909
rect 17647 23844 18349 23857
rect 17647 23792 17652 23844
rect 17704 23792 17716 23844
rect 17768 23792 17780 23844
rect 17832 23792 17844 23844
rect 17896 23792 17908 23844
rect 17960 23792 17972 23844
rect 18024 23792 18036 23844
rect 18088 23792 18100 23844
rect 18152 23792 18164 23844
rect 18216 23792 18228 23844
rect 18280 23792 18292 23844
rect 18344 23792 18349 23844
rect 17647 23779 18349 23792
rect 17647 23727 17652 23779
rect 17704 23727 17716 23779
rect 17768 23727 17780 23779
rect 17832 23727 17844 23779
rect 17896 23727 17908 23779
rect 17960 23727 17972 23779
rect 18024 23727 18036 23779
rect 18088 23727 18100 23779
rect 18152 23727 18164 23779
rect 18216 23727 18228 23779
rect 18280 23727 18292 23779
rect 18344 23727 18349 23779
rect 17647 23714 18349 23727
rect 17647 23662 17652 23714
rect 17704 23662 17716 23714
rect 17768 23662 17780 23714
rect 17832 23662 17844 23714
rect 17896 23662 17908 23714
rect 17960 23662 17972 23714
rect 18024 23662 18036 23714
rect 18088 23662 18100 23714
rect 18152 23662 18164 23714
rect 18216 23662 18228 23714
rect 18280 23662 18292 23714
rect 18344 23662 18349 23714
rect 17647 23649 18349 23662
rect 17647 23597 17652 23649
rect 17704 23597 17716 23649
rect 17768 23597 17780 23649
rect 17832 23597 17844 23649
rect 17896 23597 17908 23649
rect 17960 23597 17972 23649
rect 18024 23597 18036 23649
rect 18088 23597 18100 23649
rect 18152 23597 18164 23649
rect 18216 23597 18228 23649
rect 18280 23597 18292 23649
rect 18344 23597 18349 23649
rect 17647 23591 18349 23597
rect 1302 23503 1664 23509
rect 689 23469 701 23503
rect 735 23469 778 23503
rect 812 23469 855 23503
rect 889 23469 932 23503
rect 966 23469 1009 23503
rect 1043 23469 1086 23503
rect 1120 23469 1162 23503
rect 1196 23469 1238 23503
rect 1302 23469 1314 23503
rect 1348 23469 1390 23503
rect 1424 23469 1466 23503
rect 1500 23469 1542 23503
rect 1576 23469 1618 23503
rect 1652 23469 1664 23503
rect 689 23463 1250 23469
tri 1225 23459 1229 23463 ne
rect 1229 23460 1250 23463
rect 1302 23463 1664 23469
rect 2569 23468 2620 23561
tri 2620 23551 2630 23561 nw
tri 2854 23551 2864 23561 se
rect 2864 23551 2928 23561
tri 2851 23548 2854 23551 se
rect 2854 23548 2928 23551
tri 17249 23548 17262 23561 se
rect 17262 23548 17634 23561
rect 17855 23553 18076 23591
rect 2657 23496 2663 23548
rect 2715 23496 2727 23548
rect 2779 23496 2785 23548
rect 2787 23547 2823 23548
rect 2786 23497 2824 23547
rect 2787 23496 2823 23497
rect 2825 23496 2928 23548
tri 17234 23533 17249 23548 se
rect 17249 23533 17634 23548
tri 2620 23468 2645 23493 sw
rect 1302 23460 1323 23463
rect 1229 23459 1323 23460
tri 1323 23459 1327 23463 nw
tri 1229 23454 1234 23459 ne
rect 1234 23454 1318 23459
tri 1318 23454 1323 23459 nw
rect 222 23439 340 23449
rect 222 23410 300 23439
rect 222 23376 228 23410
rect 262 23405 300 23410
rect 334 23405 340 23439
tri 1234 23438 1250 23454 ne
rect 1250 23438 1302 23454
tri 1302 23438 1318 23454 nw
rect 2569 23416 2611 23468
rect 2663 23416 2675 23468
rect 2727 23416 2735 23468
rect 3485 23416 3491 23468
rect 3543 23416 3555 23468
rect 3607 23416 3619 23468
rect 3671 23416 3677 23468
rect 262 23376 340 23405
rect 222 23367 340 23376
rect 222 23337 300 23367
rect 222 23303 228 23337
rect 262 23333 300 23337
rect 334 23333 340 23367
rect 262 23303 340 23333
rect 222 23295 340 23303
rect 222 23264 300 23295
rect 222 23230 228 23264
rect 262 23261 300 23264
rect 334 23261 340 23295
rect 262 23230 340 23261
rect 222 23223 340 23230
rect 222 23191 300 23223
rect 222 23157 228 23191
rect 262 23189 300 23191
rect 334 23189 340 23223
rect 262 23157 340 23189
tri 2870 23182 2970 23282 se
rect 2970 23182 3100 23282
tri 340 23157 365 23182 sw
tri 2845 23157 2870 23182 se
rect 2870 23157 3100 23182
rect 222 23151 3100 23157
rect 222 23117 300 23151
rect 334 23117 373 23151
rect 407 23117 446 23151
rect 480 23117 519 23151
rect 553 23117 592 23151
rect 626 23117 665 23151
rect 699 23117 738 23151
rect 772 23117 811 23151
rect 845 23117 884 23151
rect 918 23117 957 23151
rect 991 23117 1030 23151
rect 1064 23117 1103 23151
rect 1137 23117 1176 23151
rect 1210 23117 1249 23151
rect 1283 23117 1322 23151
rect 1356 23117 1395 23151
rect 1429 23117 1468 23151
rect 1502 23117 1541 23151
rect 1575 23117 1614 23151
rect 1648 23117 1687 23151
rect 1721 23117 1760 23151
rect 1794 23117 1833 23151
rect 1867 23117 1906 23151
rect 1940 23117 1979 23151
rect 2013 23117 2052 23151
rect 2086 23117 2124 23151
rect 2158 23117 2196 23151
rect 2230 23117 2268 23151
rect 2302 23117 2340 23151
rect 2374 23117 2412 23151
rect 2446 23117 2484 23151
rect 2518 23117 2556 23151
rect 2590 23117 2628 23151
rect 2662 23117 2700 23151
rect 2734 23117 2772 23151
rect 2806 23117 2844 23151
rect 2878 23117 2916 23151
rect 2950 23117 3100 23151
rect 222 23079 3100 23117
rect 222 23045 266 23079
rect 300 23045 340 23079
rect 374 23045 414 23079
rect 448 23045 488 23079
rect 522 23045 562 23079
rect 596 23045 636 23079
rect 670 23045 710 23079
rect 744 23045 784 23079
rect 818 23045 858 23079
rect 892 23045 932 23079
rect 966 23045 1006 23079
rect 1040 23045 1080 23079
rect 1114 23045 1154 23079
rect 1188 23045 1228 23079
rect 1262 23045 1302 23079
rect 1336 23045 1376 23079
rect 1410 23045 1450 23079
rect 1484 23045 1524 23079
rect 1558 23045 1598 23079
rect 1632 23045 1672 23079
rect 1706 23045 1746 23079
rect 1780 23045 1820 23079
rect 1854 23045 1894 23079
rect 1928 23045 1967 23079
rect 2001 23045 2040 23079
rect 2074 23045 2113 23079
rect 2147 23045 2186 23079
rect 2220 23045 2259 23079
rect 2293 23045 2332 23079
rect 2366 23045 2405 23079
rect 2439 23045 2478 23079
rect 2512 23045 2551 23079
rect 2585 23045 2624 23079
rect 2658 23045 2697 23079
rect 2731 23045 2770 23079
rect 2804 23045 2843 23079
rect 2877 23045 2916 23079
rect 2950 23045 3100 23079
rect 222 23033 3100 23045
tri -186 23015 -178 23023 se
rect -178 23015 -40 23023
tri -214 22987 -186 23015 se
rect -186 22987 -80 23015
rect -158 22984 -80 22987
rect -158 22950 -152 22984
rect -118 22981 -80 22984
rect -46 22981 -40 23015
rect -118 22950 -40 22981
rect -158 22943 -40 22950
rect -158 22911 -80 22943
rect -158 22877 -152 22911
rect -118 22909 -80 22911
rect -46 22909 -40 22943
rect -118 22877 -40 22909
rect -158 22871 -40 22877
rect -158 22838 -80 22871
rect -158 22804 -152 22838
rect -118 22837 -80 22838
rect -46 22837 -40 22871
rect -118 22804 -40 22837
rect -158 22799 -40 22804
rect -158 22765 -80 22799
rect -46 22765 -40 22799
rect -158 22731 -152 22765
rect -118 22733 -40 22765
tri -40 22733 -15 22758 sw
rect -118 22731 2188 22733
rect -158 22727 2188 22731
rect -158 22693 -80 22727
rect -46 22693 -5 22727
rect 29 22693 70 22727
rect 104 22693 144 22727
rect 178 22693 218 22727
rect 252 22693 292 22727
rect 326 22693 366 22727
rect 400 22693 440 22727
rect 474 22693 514 22727
rect 548 22693 588 22727
rect 622 22693 662 22727
rect 696 22693 736 22727
rect 770 22693 810 22727
rect 844 22693 884 22727
rect 918 22693 958 22727
rect 992 22693 1032 22727
rect 1066 22693 1106 22727
rect 1140 22693 1180 22727
rect 1214 22693 1254 22727
rect 1288 22693 1328 22727
rect 1362 22693 1402 22727
rect 1436 22693 1476 22727
rect 1510 22693 1550 22727
rect 1584 22693 1624 22727
rect 1658 22693 1698 22727
rect 1732 22693 1772 22727
rect 1806 22693 1846 22727
rect 1880 22693 1920 22727
rect 1954 22693 1994 22727
rect 2028 22693 2068 22727
rect 2102 22693 2142 22727
rect 2176 22693 2188 22727
rect -158 22655 2188 22693
rect -158 22621 -114 22655
rect -80 22621 -41 22655
rect -7 22621 32 22655
rect 66 22621 105 22655
rect 139 22621 178 22655
rect 212 22621 251 22655
rect 285 22621 324 22655
rect 358 22621 397 22655
rect 431 22621 470 22655
rect 504 22621 543 22655
rect 577 22621 616 22655
rect 650 22621 689 22655
rect 723 22621 762 22655
rect 796 22621 835 22655
rect 869 22621 908 22655
rect 942 22621 981 22655
rect 1015 22621 1054 22655
rect 1088 22621 1127 22655
rect 1161 22621 1200 22655
rect 1234 22621 1273 22655
rect 1307 22621 1346 22655
rect 1380 22621 1419 22655
rect 1453 22621 1492 22655
rect 1526 22621 1565 22655
rect 1599 22621 1638 22655
rect 1672 22621 1710 22655
rect 1744 22621 1782 22655
rect 1816 22621 1854 22655
rect 1888 22621 1926 22655
rect 1960 22621 1998 22655
rect 2032 22621 2070 22655
rect 2104 22621 2142 22655
rect 2176 22621 2188 22655
rect -158 22615 2188 22621
rect 236 22581 448 22587
rect 288 22529 396 22581
rect 236 22517 448 22529
rect 288 22465 396 22517
rect 236 22459 448 22465
rect -25 20619 27 20625
rect -25 20555 27 20567
rect -25 20445 27 20503
tri -25 20418 2 20445 ne
rect 2 20418 27 20445
tri 27 20418 76 20467 sw
tri 2 20393 27 20418 ne
rect 27 20393 396 20418
tri 27 20366 54 20393 ne
rect 54 20366 396 20393
tri 396 20366 448 20418 sw
tri 368 20357 377 20366 ne
rect 377 20357 448 20366
tri 377 20338 396 20357 ne
rect 396 20351 448 20357
rect 396 20287 448 20299
rect 396 20229 448 20235
rect -2205 18343 1753 18349
rect -2205 18309 -2089 18343
rect -2055 18309 -2016 18343
rect -1982 18309 -1943 18343
rect -1909 18309 -1870 18343
rect -1836 18309 -1797 18343
rect -1763 18309 -1724 18343
rect -1690 18309 -1651 18343
rect -1617 18309 -1578 18343
rect -1544 18309 -1505 18343
rect -1471 18309 -1432 18343
rect -1398 18309 -1359 18343
rect -1325 18309 -1286 18343
rect -1252 18309 -1213 18343
rect -1179 18309 -1140 18343
rect -1106 18309 -1067 18343
rect -1033 18309 -994 18343
rect -960 18309 -921 18343
rect -887 18309 -848 18343
rect -814 18309 -775 18343
rect -741 18309 -702 18343
rect -668 18309 -629 18343
rect -595 18309 -556 18343
rect -522 18309 -483 18343
rect -449 18309 -410 18343
rect -376 18309 -337 18343
rect -303 18309 -264 18343
rect -230 18309 -191 18343
rect -157 18309 -118 18343
rect -84 18309 -45 18343
rect -11 18309 28 18343
rect 62 18309 101 18343
rect 135 18309 174 18343
rect 208 18309 247 18343
rect 281 18309 320 18343
rect 354 18309 393 18343
rect 427 18309 466 18343
rect 500 18309 539 18343
rect 573 18309 612 18343
rect 646 18309 685 18343
rect 719 18309 758 18343
rect 792 18309 831 18343
rect 865 18309 904 18343
rect 938 18309 977 18343
rect 1011 18309 1050 18343
rect 1084 18309 1123 18343
rect 1157 18309 1196 18343
rect 1230 18309 1269 18343
rect 1303 18309 1342 18343
rect 1376 18309 1415 18343
rect 1449 18309 1488 18343
rect 1522 18309 1561 18343
rect 1595 18309 1634 18343
rect 1668 18309 1707 18343
rect 1741 18309 1753 18343
rect -2205 18305 1753 18309
rect -2205 18271 -2199 18305
rect -2165 18271 1753 18305
rect -2205 18237 -2127 18271
rect -2093 18237 -2055 18271
rect -2021 18237 -1983 18271
rect -1949 18237 -1911 18271
rect -1877 18237 -1839 18271
rect -1805 18237 -1767 18271
rect -1733 18237 -1695 18271
rect -1661 18237 -1623 18271
rect -1589 18237 -1551 18271
rect -1517 18237 -1479 18271
rect -1445 18237 -1407 18271
rect -1373 18237 -1335 18271
rect -1301 18237 -1263 18271
rect -1229 18237 -1191 18271
rect -1157 18237 -1119 18271
rect -1085 18237 -1047 18271
rect -1013 18237 -975 18271
rect -941 18237 -903 18271
rect -869 18237 -831 18271
rect -797 18237 -759 18271
rect -725 18237 -687 18271
rect -653 18237 -615 18271
rect -581 18237 -543 18271
rect -509 18237 -471 18271
rect -437 18237 -399 18271
rect -365 18237 -327 18271
rect -293 18237 -255 18271
rect -221 18237 -183 18271
rect -149 18237 -111 18271
rect -77 18237 -39 18271
rect -5 18237 33 18271
rect 67 18237 105 18271
rect 139 18237 177 18271
rect 211 18237 249 18271
rect 283 18237 321 18271
rect 355 18237 393 18271
rect 427 18237 466 18271
rect 500 18237 539 18271
rect 573 18237 612 18271
rect 646 18237 685 18271
rect 719 18237 758 18271
rect 792 18237 831 18271
rect 865 18237 904 18271
rect 938 18237 977 18271
rect 1011 18237 1050 18271
rect 1084 18237 1123 18271
rect 1157 18237 1196 18271
rect 1230 18237 1269 18271
rect 1303 18237 1342 18271
rect 1376 18237 1415 18271
rect 1449 18237 1488 18271
rect 1522 18237 1561 18271
rect 1595 18237 1634 18271
rect 1668 18237 1707 18271
rect 1741 18237 1753 18271
rect -2205 18233 1753 18237
rect -2205 18199 -2199 18233
rect -2165 18231 1753 18233
rect -2165 18199 -2087 18231
rect -2205 18180 -2087 18199
rect -2205 18161 -2127 18180
rect -2205 18127 -2199 18161
rect -2165 18146 -2127 18161
rect -2093 18146 -2087 18180
rect -2165 18127 -2087 18146
rect -2205 18089 -2087 18127
rect -2205 18055 -2199 18089
rect -2165 18055 -2127 18089
rect -2093 18055 -2087 18089
rect -2205 18043 -2087 18055
rect 481 5001 927 5007
rect 979 5001 991 5007
rect 1043 5001 1069 5007
rect 481 4967 493 5001
rect 527 4967 569 5001
rect 603 4967 645 5001
rect 679 4967 721 5001
rect 755 4967 797 5001
rect 831 4967 873 5001
rect 907 4967 927 5001
rect 982 4967 991 5001
rect 1057 4967 1069 5001
rect 481 4961 927 4967
tri 915 4955 921 4961 ne
rect 921 4955 927 4961
rect 979 4955 991 4967
rect 1043 4961 1069 4967
rect 1043 4955 1049 4961
tri 1049 4955 1055 4961 nw
rect -3494 4902 -405 4954
rect 1036 4886 1088 4892
tri 1014 4854 1036 4876 se
rect -2848 4802 -2842 4854
rect -2790 4802 -2778 4854
rect -2726 4851 -2720 4854
tri 1011 4851 1014 4854 se
rect 1014 4851 1036 4854
rect -2726 4845 1036 4851
rect -2726 4811 493 4845
rect 527 4811 569 4845
rect 603 4811 645 4845
rect 679 4811 721 4845
rect 755 4811 797 4845
rect 831 4811 873 4845
rect 907 4811 948 4845
rect 982 4811 1023 4845
rect 1057 4822 1088 4834
rect -2726 4805 1036 4811
rect -2726 4802 -2720 4805
tri 1011 4802 1014 4805 ne
rect 1014 4802 1036 4805
tri 1014 4780 1036 4802 ne
rect 956 4762 1008 4768
rect 1036 4764 1088 4770
rect 956 4698 1008 4710
rect -3088 4641 -3036 4647
rect -2928 4643 -2922 4695
rect -2870 4643 -2858 4695
rect -2806 4689 956 4695
tri 1008 4695 1033 4720 sw
rect 1008 4689 1069 4695
rect -2806 4655 493 4689
rect 527 4655 569 4689
rect 603 4655 645 4689
rect 679 4655 721 4689
rect 755 4655 797 4689
rect 831 4655 873 4689
rect 907 4655 948 4689
rect 1008 4655 1023 4689
rect 1057 4655 1069 4689
rect -2806 4649 956 4655
rect -2806 4643 -2800 4649
tri 931 4643 937 4649 ne
rect 937 4646 956 4649
rect 1008 4649 1069 4655
rect 1008 4646 1024 4649
rect 937 4643 1024 4646
tri 937 4640 940 4643 ne
rect 940 4640 1024 4643
tri 1024 4640 1033 4649 nw
tri 940 4624 956 4640 ne
rect 956 4624 1008 4640
tri 1008 4624 1024 4640 nw
tri 780 4594 796 4610 se
rect 796 4594 848 4610
tri 848 4594 864 4610 sw
rect -3088 4585 -3036 4589
tri 771 4585 780 4594 se
rect 780 4588 864 4594
rect 780 4585 796 4588
rect -3088 4579 796 4585
rect 848 4585 864 4588
tri 864 4585 873 4594 sw
rect 848 4579 1069 4585
rect -3088 4577 493 4579
rect -3036 4545 493 4577
rect 527 4545 569 4579
rect 603 4545 645 4579
rect 679 4545 721 4579
rect 755 4545 796 4579
rect 848 4545 873 4579
rect 907 4545 948 4579
rect 982 4545 1023 4579
rect 1057 4545 1069 4579
rect -3036 4539 796 4545
rect -3088 4519 -3036 4525
tri 771 4519 791 4539 ne
rect 791 4536 796 4539
rect 848 4539 1069 4545
rect 791 4524 848 4536
rect 791 4519 796 4524
tri 791 4514 796 4519 ne
tri 848 4514 873 4539 nw
rect 796 4466 848 4472
rect 876 4464 928 4470
tri 855 4433 876 4454 se
rect -3008 4381 -3002 4433
rect -2950 4381 -2938 4433
rect -2886 4430 -2880 4433
tri 852 4430 855 4433 se
rect 855 4430 876 4433
rect -2886 4429 481 4430
tri 851 4429 852 4430 se
rect 852 4429 876 4430
rect -2886 4423 876 4429
rect 928 4423 1069 4429
rect -2886 4389 493 4423
rect 527 4389 569 4423
rect 603 4389 645 4423
rect 679 4389 721 4423
rect 755 4389 797 4423
rect 831 4389 873 4423
rect 928 4412 948 4423
rect 907 4400 948 4412
rect 928 4389 948 4400
rect 982 4389 1023 4423
rect 1057 4389 1069 4423
rect -2886 4384 876 4389
rect -2886 4381 -2880 4384
rect 481 4383 876 4384
tri 851 4381 853 4383 ne
rect 853 4381 876 4383
tri 853 4358 876 4381 ne
rect 928 4383 1069 4389
rect 796 4340 848 4346
rect 876 4342 928 4348
tri 771 4273 796 4298 se
rect 796 4276 848 4288
rect 481 4267 796 4273
tri 848 4273 873 4298 sw
rect 848 4267 1069 4273
rect 481 4233 493 4267
rect 527 4233 569 4267
rect 603 4233 645 4267
rect 679 4233 721 4267
rect 755 4233 796 4267
rect 848 4233 873 4267
rect 907 4233 948 4267
rect 982 4233 1023 4267
rect 1057 4233 1069 4267
rect 481 4227 796 4233
tri 771 4218 780 4227 ne
rect 780 4224 796 4227
rect 848 4227 1069 4233
rect 848 4224 864 4227
rect 780 4218 864 4224
tri 864 4218 873 4227 nw
tri 780 4202 796 4218 ne
rect 796 4202 848 4218
tri 848 4202 864 4218 nw
<< rmetal1 >>
rect 15693 26971 15893 26972
rect 15693 26970 15694 26971
rect 15892 26970 15893 26971
rect 15693 26933 15694 26934
rect 15892 26933 15893 26934
rect 15693 26932 15893 26933
rect 16517 26971 16717 26972
rect 16517 26970 16518 26971
rect 16716 26970 16717 26971
rect 16517 26933 16518 26934
rect 16716 26933 16717 26934
rect 16517 26932 16717 26933
rect 17341 26992 17550 26994
tri 17550 26992 17552 26994 sw
tri 17550 26990 17552 26992 ne
tri 17552 26990 17554 26992 sw
tri 17552 26988 17554 26990 ne
tri 17554 26988 17556 26990 sw
tri 17554 26986 17556 26988 ne
tri 17556 26986 17558 26988 sw
tri 17556 26984 17558 26986 ne
tri 17558 26984 17560 26986 sw
tri 17558 26982 17560 26984 ne
tri 17560 26982 17562 26984 sw
tri 17560 26980 17562 26982 ne
tri 17562 26980 17564 26982 sw
tri 17562 26978 17564 26980 ne
tri 17564 26978 17566 26980 sw
tri 17564 26976 17566 26978 ne
tri 17566 26976 17568 26978 sw
tri 17566 26974 17568 26976 ne
tri 17568 26974 17570 26976 sw
tri 17568 26972 17570 26974 ne
tri 17570 26972 17572 26974 sw
tri 17570 26970 17572 26972 ne
tri 17572 26970 17574 26972 sw
tri 17572 26968 17574 26970 ne
tri 17574 26968 17576 26970 sw
tri 17574 26966 17576 26968 ne
tri 17576 26966 17578 26968 sw
tri 17576 26964 17578 26966 ne
tri 17578 26964 17580 26966 sw
rect 17341 26962 17512 26964
tri 17512 26962 17514 26964 sw
tri 17578 26962 17580 26964 ne
tri 17580 26962 17582 26964 sw
tri 17512 26960 17514 26962 ne
tri 17514 26960 17516 26962 sw
tri 17514 26958 17516 26960 ne
tri 17516 26958 17518 26960 sw
tri 17516 26956 17518 26958 ne
tri 17518 26956 17520 26958 sw
tri 17518 26954 17520 26956 ne
tri 17520 26954 17522 26956 sw
tri 17520 26952 17522 26954 ne
tri 17522 26952 17524 26954 sw
tri 17522 26950 17524 26952 ne
tri 17524 26950 17526 26952 sw
tri 17524 26948 17526 26950 ne
tri 17526 26948 17528 26950 sw
tri 17526 26946 17528 26948 ne
tri 17528 26946 17530 26948 sw
tri 17528 26944 17530 26946 ne
tri 17530 26944 17532 26946 sw
tri 17530 26942 17532 26944 ne
tri 17532 26942 17534 26944 sw
tri 17532 26940 17534 26942 ne
tri 17534 26940 17536 26942 sw
tri 17534 26938 17536 26940 ne
tri 17536 26938 17538 26940 sw
tri 17536 26936 17538 26938 ne
tri 17538 26936 17540 26938 sw
tri 17538 26934 17540 26936 ne
tri 17540 26934 17542 26936 sw
tri 17540 26932 17542 26934 ne
tri 17542 26932 17544 26934 sw
rect 17542 26879 17544 26932
rect 17580 26879 17582 26962
rect 17542 23875 17543 26879
rect 17581 23875 17582 26879
rect 17542 23822 17544 23875
tri 17540 23820 17542 23822 se
tri 17542 23820 17544 23822 nw
tri 17538 23818 17540 23820 se
tri 17540 23818 17542 23820 nw
tri 17536 23816 17538 23818 se
tri 17538 23816 17540 23818 nw
tri 17534 23814 17536 23816 se
tri 17536 23814 17538 23816 nw
tri 17532 23812 17534 23814 se
tri 17534 23812 17536 23814 nw
tri 17530 23810 17532 23812 se
tri 17532 23810 17534 23812 nw
tri 17528 23808 17530 23810 se
tri 17530 23808 17532 23810 nw
tri 17526 23806 17528 23808 se
tri 17528 23806 17530 23808 nw
tri 17524 23804 17526 23806 se
tri 17526 23804 17528 23806 nw
tri 17522 23802 17524 23804 se
tri 17524 23802 17526 23804 nw
tri 17520 23800 17522 23802 se
tri 17522 23800 17524 23802 nw
tri 17518 23798 17520 23800 se
tri 17520 23798 17522 23800 nw
tri 17516 23796 17518 23798 se
tri 17518 23796 17520 23798 nw
tri 17514 23794 17516 23796 se
tri 17516 23794 17518 23796 nw
tri 17512 23792 17514 23794 se
tri 17514 23792 17516 23794 nw
rect 17580 23792 17582 23875
rect 17341 23790 17512 23792
tri 17512 23790 17514 23792 nw
tri 17578 23790 17580 23792 se
tri 17580 23790 17582 23792 nw
tri 17576 23788 17578 23790 se
tri 17578 23788 17580 23790 nw
rect 2785 23787 2787 23788
rect 2823 23787 2825 23788
rect 2785 23737 2786 23787
rect 2824 23737 2825 23787
rect 2785 23736 2787 23737
rect 2823 23736 2825 23737
rect 4649 23787 4651 23788
rect 4687 23787 4689 23788
rect 4649 23737 4650 23787
rect 4688 23737 4689 23787
rect 5061 23787 5063 23788
rect 5099 23787 5101 23788
rect 4649 23736 4651 23737
rect 4687 23736 4689 23737
rect 5061 23737 5062 23787
rect 5100 23737 5101 23787
rect 5473 23787 5475 23788
rect 5511 23787 5513 23788
rect 5061 23736 5063 23737
rect 5099 23736 5101 23737
rect 5473 23737 5474 23787
rect 5512 23737 5513 23787
rect 5885 23787 5887 23788
rect 5923 23787 5925 23788
rect 5473 23736 5475 23737
rect 5511 23736 5513 23737
rect 5885 23737 5886 23787
rect 5924 23737 5925 23787
rect 6297 23787 6299 23788
rect 6335 23787 6337 23788
rect 5885 23736 5887 23737
rect 5923 23736 5925 23737
rect 6297 23737 6298 23787
rect 6336 23737 6337 23787
rect 6709 23787 6711 23788
rect 6297 23736 6299 23737
rect 6335 23736 6337 23737
rect 6709 23737 6710 23787
rect 6709 23736 6711 23737
rect 6747 23787 6749 23788
rect 6748 23737 6749 23787
rect 6747 23736 6749 23737
rect 7121 23787 7123 23788
rect 7159 23787 7161 23788
rect 7121 23737 7122 23787
rect 7160 23737 7161 23787
rect 7533 23787 7535 23788
rect 7571 23787 7573 23788
rect 7121 23736 7123 23737
rect 7159 23736 7161 23737
rect 7533 23737 7534 23787
rect 7572 23737 7573 23787
rect 7850 23787 7852 23788
rect 7888 23787 7890 23788
rect 7533 23736 7535 23737
rect 7571 23736 7573 23737
rect 7850 23737 7851 23787
rect 7889 23737 7890 23787
rect 7850 23736 7852 23737
rect 7888 23736 7890 23737
rect 8039 23787 8041 23788
rect 8077 23787 8079 23788
rect 8039 23737 8040 23787
rect 8078 23737 8079 23787
rect 8357 23787 8359 23788
rect 8395 23787 8397 23788
rect 8039 23736 8041 23737
rect 8077 23736 8079 23737
rect 8357 23737 8358 23787
rect 8396 23737 8397 23787
rect 8769 23787 8771 23788
rect 8357 23736 8359 23737
rect 8395 23736 8397 23737
rect 8769 23737 8770 23787
rect 8769 23736 8771 23737
rect 8807 23787 8809 23788
rect 8808 23737 8809 23787
rect 9181 23787 9183 23788
rect 9219 23787 9221 23788
rect 8807 23736 8809 23737
rect 9181 23737 9182 23787
rect 9220 23737 9221 23787
rect 9593 23787 9595 23788
rect 9631 23787 9633 23788
rect 9181 23736 9183 23737
rect 9219 23736 9221 23737
rect 9593 23737 9594 23787
rect 9632 23737 9633 23787
rect 10005 23787 10007 23788
rect 10043 23787 10045 23788
rect 9593 23736 9595 23737
rect 9631 23736 9633 23737
rect 10005 23737 10006 23787
rect 10044 23737 10045 23787
rect 10417 23787 10419 23788
rect 10455 23787 10457 23788
rect 10005 23736 10007 23737
rect 10043 23736 10045 23737
rect 10417 23737 10418 23787
rect 10456 23737 10457 23787
rect 10829 23787 10831 23788
rect 10867 23787 10869 23788
rect 10417 23736 10419 23737
rect 10455 23736 10457 23737
rect 10829 23737 10830 23787
rect 10868 23737 10869 23787
rect 10829 23736 10831 23737
rect 10867 23736 10869 23737
rect 11362 23787 11364 23788
rect 11400 23787 11402 23788
rect 11362 23737 11363 23787
rect 11401 23737 11402 23787
rect 11532 23787 11534 23788
rect 11362 23736 11364 23737
rect 11400 23736 11402 23737
rect 11532 23737 11533 23787
rect 11532 23736 11534 23737
rect 11570 23787 11572 23788
rect 11571 23737 11572 23787
rect 11774 23787 11776 23788
rect 11570 23736 11572 23737
rect 11774 23737 11775 23787
rect 11774 23736 11776 23737
rect 11812 23787 11814 23788
rect 11813 23737 11814 23787
rect 11944 23787 11946 23788
rect 11982 23787 11984 23788
rect 11812 23736 11814 23737
rect 11944 23737 11945 23787
rect 11983 23737 11984 23787
rect 12186 23787 12188 23788
rect 12224 23787 12226 23788
rect 11944 23736 11946 23737
rect 11982 23736 11984 23737
rect 12186 23737 12187 23787
rect 12225 23737 12226 23787
rect 12356 23787 12358 23788
rect 12186 23736 12188 23737
rect 12224 23736 12226 23737
rect 12356 23737 12357 23787
rect 12356 23736 12358 23737
rect 12394 23787 12396 23788
rect 12395 23737 12396 23787
rect 12598 23787 12600 23788
rect 12394 23736 12396 23737
rect 12598 23737 12599 23787
rect 12598 23736 12600 23737
rect 12636 23787 12638 23788
rect 12637 23737 12638 23787
rect 12768 23787 12770 23788
rect 12806 23787 12808 23788
rect 12636 23736 12638 23737
rect 12768 23737 12769 23787
rect 12807 23737 12808 23787
rect 13010 23787 13012 23788
rect 13048 23787 13050 23788
rect 12768 23736 12770 23737
rect 12806 23736 12808 23737
rect 13010 23737 13011 23787
rect 13049 23737 13050 23787
rect 13180 23787 13182 23788
rect 13010 23736 13012 23737
rect 13048 23736 13050 23737
rect 13180 23737 13181 23787
rect 13180 23736 13182 23737
rect 13218 23787 13220 23788
rect 13219 23737 13220 23787
rect 13422 23787 13424 23788
rect 13218 23736 13220 23737
rect 13422 23737 13423 23787
rect 13422 23736 13424 23737
rect 13460 23787 13462 23788
rect 13461 23737 13462 23787
rect 13592 23787 13594 23788
rect 13630 23787 13632 23788
rect 13460 23736 13462 23737
rect 13592 23737 13593 23787
rect 13631 23737 13632 23787
rect 13834 23787 13836 23788
rect 13592 23736 13594 23737
rect 13630 23736 13632 23737
rect 13834 23737 13835 23787
rect 13834 23736 13836 23737
rect 13872 23787 13874 23788
rect 13873 23737 13874 23787
rect 14004 23787 14006 23788
rect 14042 23787 14044 23788
rect 13872 23736 13874 23737
rect 14004 23737 14005 23787
rect 14043 23737 14044 23787
rect 14246 23787 14248 23788
rect 14284 23787 14286 23788
rect 14004 23736 14006 23737
rect 14042 23736 14044 23737
rect 14246 23737 14247 23787
rect 14285 23737 14286 23787
rect 14416 23787 14418 23788
rect 14246 23736 14248 23737
rect 14284 23736 14286 23737
rect 14416 23737 14417 23787
rect 14416 23736 14418 23737
rect 14454 23787 14456 23788
rect 14455 23737 14456 23787
tri 17574 23786 17576 23788 se
tri 17576 23786 17578 23788 nw
tri 17573 23785 17574 23786 se
rect 17574 23785 17575 23786
tri 17575 23785 17576 23786 nw
rect 14454 23736 14456 23737
rect 14947 23784 14949 23785
rect 14947 23740 14948 23784
rect 14947 23739 14949 23740
rect 14985 23784 14987 23785
rect 14986 23740 14987 23784
rect 14985 23739 14987 23740
rect 15895 23784 15897 23785
rect 15933 23784 15935 23785
rect 15895 23740 15896 23784
rect 15934 23740 15935 23784
rect 16296 23784 16298 23785
rect 16334 23784 16336 23785
rect 15895 23739 15897 23740
rect 15933 23739 15935 23740
rect 16296 23740 16297 23784
rect 16335 23740 16336 23784
rect 16719 23784 16721 23785
rect 16757 23784 16759 23785
rect 16296 23739 16298 23740
rect 16334 23739 16336 23740
rect 16719 23740 16720 23784
rect 16758 23740 16759 23784
rect 16890 23784 16892 23785
rect 16928 23784 16930 23785
rect 16719 23739 16721 23740
rect 16757 23739 16759 23740
rect 16890 23740 16891 23784
rect 16929 23740 16930 23784
rect 16890 23739 16892 23740
rect 16928 23739 16930 23740
tri 17572 23784 17573 23785 se
rect 17573 23784 17574 23785
tri 17574 23784 17575 23785 nw
tri 17570 23782 17572 23784 se
tri 17572 23782 17574 23784 nw
tri 17568 23780 17570 23782 se
tri 17570 23780 17572 23782 nw
tri 17566 23778 17568 23780 se
tri 17568 23778 17570 23780 nw
tri 17564 23776 17566 23778 se
tri 17566 23776 17568 23778 nw
tri 17562 23774 17564 23776 se
tri 17564 23774 17566 23776 nw
tri 17560 23772 17562 23774 se
tri 17562 23772 17564 23774 nw
tri 17558 23770 17560 23772 se
tri 17560 23770 17562 23772 nw
tri 17556 23768 17558 23770 se
tri 17558 23768 17560 23770 nw
tri 17554 23766 17556 23768 se
tri 17556 23766 17558 23768 nw
tri 17552 23764 17554 23766 se
tri 17554 23764 17556 23766 nw
tri 17550 23762 17552 23764 se
tri 17552 23762 17554 23764 nw
rect 17341 23760 17550 23762
tri 17550 23760 17552 23762 nw
rect 16956 23664 17084 23665
rect 16956 23663 16957 23664
rect 17083 23663 17084 23664
rect 16956 23626 16957 23627
rect 17083 23626 17084 23627
rect 16956 23625 17084 23626
rect 2785 23547 2787 23548
rect 2823 23547 2825 23548
rect 2785 23497 2786 23547
rect 2824 23497 2825 23547
rect 2785 23496 2787 23497
rect 2823 23496 2825 23497
<< via1 >>
rect 10783 27511 10835 27563
rect 10847 27511 10899 27563
rect 10826 27431 10878 27483
rect 10890 27431 10942 27483
rect 6639 27229 6819 27345
rect 4197 26955 4249 27007
rect 4261 26955 4313 27007
rect 10667 26784 10719 26836
rect 10667 26720 10719 26772
rect 2876 26528 2928 26580
rect 2876 26464 2928 26516
rect 7015 26510 7067 26562
rect 7079 26510 7131 26562
rect 7143 26510 7195 26562
rect 7207 26510 7259 26562
rect 7271 26510 7323 26562
rect 8599 26510 8651 26562
rect 8663 26510 8715 26562
rect 8727 26510 8779 26562
rect 8791 26510 8843 26562
rect 8855 26510 8907 26562
rect 5055 26458 5107 26510
rect 5119 26458 5171 26510
rect 666 25097 718 25149
rect 730 25097 782 25149
rect 1090 24237 1142 24246
rect 1090 24203 1120 24237
rect 1120 24203 1142 24237
rect 1090 24194 1142 24203
rect 1090 24130 1142 24182
rect 1170 24081 1222 24122
rect 1170 24070 1196 24081
rect 1196 24070 1222 24081
rect 1170 24047 1196 24058
rect 1196 24047 1222 24058
rect 1170 24006 1222 24047
rect 1090 23946 1142 23998
rect 1090 23925 1142 23934
rect 1090 23891 1120 23925
rect 1120 23891 1142 23925
rect 1090 23882 1142 23891
rect 1250 23815 1302 23824
rect 1250 23781 1272 23815
rect 1272 23781 1302 23815
rect 1250 23772 1302 23781
rect 1250 23708 1302 23760
rect 4508 24216 4560 24268
rect 4572 24216 4624 24268
rect 4636 24216 4688 24268
rect 4700 24216 4752 24268
rect 4764 24216 4816 24268
rect 5332 24216 5384 24268
rect 5396 24216 5448 24268
rect 5460 24216 5512 24268
rect 5524 24216 5576 24268
rect 5588 24216 5640 24268
rect 6156 24216 6208 24268
rect 6220 24216 6272 24268
rect 6284 24216 6336 24268
rect 6348 24216 6400 24268
rect 6412 24216 6464 24268
rect 6980 24216 7032 24268
rect 7044 24216 7096 24268
rect 7108 24216 7160 24268
rect 7172 24216 7224 24268
rect 7236 24216 7288 24268
rect 7804 24216 7856 24268
rect 7868 24216 7920 24268
rect 7932 24216 7984 24268
rect 7996 24216 8048 24268
rect 8060 24216 8112 24268
rect 8628 24216 8680 24268
rect 8692 24216 8744 24268
rect 8756 24216 8808 24268
rect 8820 24216 8872 24268
rect 8884 24216 8936 24268
rect 9466 24216 9518 24268
rect 9530 24216 9582 24268
rect 9594 24216 9646 24268
rect 9658 24216 9710 24268
rect 9722 24216 9774 24268
rect 10276 24216 10328 24268
rect 10340 24216 10392 24268
rect 10404 24216 10456 24268
rect 10468 24216 10520 24268
rect 10532 24216 10584 24268
rect 10667 24097 10719 24149
rect 10667 24033 10719 24085
rect 10979 26500 11031 26552
rect 11202 26510 11254 26562
rect 11266 26510 11318 26562
rect 11330 26510 11382 26562
rect 11394 26510 11446 26562
rect 12722 26510 12774 26562
rect 12786 26510 12838 26562
rect 12850 26510 12902 26562
rect 12914 26510 12966 26562
rect 12978 26510 13030 26562
rect 15260 26510 15312 26562
rect 15324 26510 15376 26562
rect 15388 26510 15440 26562
rect 15452 26510 15504 26562
rect 15516 26510 15568 26562
rect 16844 26510 16896 26562
rect 16908 26510 16960 26562
rect 16972 26510 17024 26562
rect 17036 26510 17088 26562
rect 17100 26510 17152 26562
rect 10979 26436 11031 26488
rect 11086 24216 11138 24268
rect 11150 24216 11202 24268
rect 11214 24216 11266 24268
rect 11278 24216 11330 24268
rect 11342 24216 11394 24268
rect 11924 24216 11976 24268
rect 11988 24216 12040 24268
rect 12052 24216 12104 24268
rect 12116 24216 12168 24268
rect 12180 24216 12232 24268
rect 12748 24216 12800 24268
rect 12812 24216 12864 24268
rect 12876 24216 12928 24268
rect 12940 24216 12992 24268
rect 13004 24216 13056 24268
rect 13572 24216 13624 24268
rect 13636 24216 13688 24268
rect 13700 24216 13752 24268
rect 13764 24216 13816 24268
rect 13828 24216 13880 24268
rect 14396 24216 14448 24268
rect 14460 24216 14512 24268
rect 14524 24216 14576 24268
rect 14588 24216 14640 24268
rect 14652 24216 14704 24268
rect 15220 24216 15272 24268
rect 15284 24216 15336 24268
rect 15348 24216 15400 24268
rect 15412 24216 15464 24268
rect 15476 24216 15528 24268
rect 16044 24216 16096 24268
rect 16108 24216 16160 24268
rect 16172 24216 16224 24268
rect 16236 24216 16288 24268
rect 16300 24216 16352 24268
rect 16868 24216 16920 24268
rect 16932 24216 16984 24268
rect 16996 24216 17048 24268
rect 17060 24216 17112 24268
rect 17124 24216 17176 24268
rect 10979 24097 11031 24149
rect 10979 24033 11031 24085
rect 2663 23736 2715 23788
rect 2727 23736 2779 23788
rect 6998 23736 7050 23788
rect 7062 23736 7114 23788
rect 7904 23736 7956 23788
rect 7968 23736 8020 23788
rect 15173 23779 15225 23785
rect 15173 23745 15196 23779
rect 15196 23745 15225 23779
rect 15173 23733 15225 23745
rect 15238 23733 15290 23785
rect 15342 23733 15394 23785
rect 15407 23733 15459 23785
rect 1330 23659 1382 23700
rect 1330 23648 1348 23659
rect 1348 23648 1382 23659
rect 1330 23625 1348 23636
rect 1348 23625 1382 23636
rect 1330 23584 1382 23625
rect 1250 23524 1302 23576
rect 1250 23503 1302 23512
rect 4223 23656 4275 23708
rect 4287 23656 4339 23708
rect 4223 23576 4275 23628
rect 4287 23576 4339 23628
rect 15216 23609 15268 23661
rect 15285 23609 15337 23661
rect 15353 23609 15405 23661
rect 16828 23643 16880 23695
rect 16828 23578 16880 23630
rect 16962 23561 17014 23613
rect 17026 23561 17078 23613
rect 17652 24767 18344 26035
rect 17652 24702 17704 24754
rect 17716 24702 17768 24754
rect 17780 24702 17832 24754
rect 17844 24702 17896 24754
rect 17908 24702 17960 24754
rect 17972 24702 18024 24754
rect 18036 24702 18088 24754
rect 18100 24702 18152 24754
rect 18164 24702 18216 24754
rect 18228 24702 18280 24754
rect 18292 24702 18344 24754
rect 17652 24637 17704 24689
rect 17716 24637 17768 24689
rect 17780 24637 17832 24689
rect 17844 24637 17896 24689
rect 17908 24637 17960 24689
rect 17972 24637 18024 24689
rect 18036 24637 18088 24689
rect 18100 24637 18152 24689
rect 18164 24637 18216 24689
rect 18228 24637 18280 24689
rect 18292 24637 18344 24689
rect 17652 24572 17704 24624
rect 17716 24572 17768 24624
rect 17780 24572 17832 24624
rect 17844 24572 17896 24624
rect 17908 24572 17960 24624
rect 17972 24572 18024 24624
rect 18036 24572 18088 24624
rect 18100 24572 18152 24624
rect 18164 24572 18216 24624
rect 18228 24572 18280 24624
rect 18292 24572 18344 24624
rect 17652 24507 17704 24559
rect 17716 24507 17768 24559
rect 17780 24507 17832 24559
rect 17844 24507 17896 24559
rect 17908 24507 17960 24559
rect 17972 24507 18024 24559
rect 18036 24507 18088 24559
rect 18100 24507 18152 24559
rect 18164 24507 18216 24559
rect 18228 24507 18280 24559
rect 18292 24507 18344 24559
rect 17652 24442 17704 24494
rect 17716 24442 17768 24494
rect 17780 24442 17832 24494
rect 17844 24442 17896 24494
rect 17908 24442 17960 24494
rect 17972 24442 18024 24494
rect 18036 24442 18088 24494
rect 18100 24442 18152 24494
rect 18164 24442 18216 24494
rect 18228 24442 18280 24494
rect 18292 24442 18344 24494
rect 17652 24377 17704 24429
rect 17716 24377 17768 24429
rect 17780 24377 17832 24429
rect 17844 24377 17896 24429
rect 17908 24377 17960 24429
rect 17972 24377 18024 24429
rect 18036 24377 18088 24429
rect 18100 24377 18152 24429
rect 18164 24377 18216 24429
rect 18228 24377 18280 24429
rect 18292 24377 18344 24429
rect 17652 24312 17704 24364
rect 17716 24312 17768 24364
rect 17780 24312 17832 24364
rect 17844 24312 17896 24364
rect 17908 24312 17960 24364
rect 17972 24312 18024 24364
rect 18036 24312 18088 24364
rect 18100 24312 18152 24364
rect 18164 24312 18216 24364
rect 18228 24312 18280 24364
rect 18292 24312 18344 24364
rect 17652 24247 17704 24299
rect 17716 24247 17768 24299
rect 17780 24247 17832 24299
rect 17844 24247 17896 24299
rect 17908 24247 17960 24299
rect 17972 24247 18024 24299
rect 18036 24247 18088 24299
rect 18100 24247 18152 24299
rect 18164 24247 18216 24299
rect 18228 24247 18280 24299
rect 18292 24247 18344 24299
rect 17652 24182 17704 24234
rect 17716 24182 17768 24234
rect 17780 24182 17832 24234
rect 17844 24182 17896 24234
rect 17908 24182 17960 24234
rect 17972 24182 18024 24234
rect 18036 24182 18088 24234
rect 18100 24182 18152 24234
rect 18164 24182 18216 24234
rect 18228 24182 18280 24234
rect 18292 24182 18344 24234
rect 17652 24117 17704 24169
rect 17716 24117 17768 24169
rect 17780 24117 17832 24169
rect 17844 24117 17896 24169
rect 17908 24117 17960 24169
rect 17972 24117 18024 24169
rect 18036 24117 18088 24169
rect 18100 24117 18152 24169
rect 18164 24117 18216 24169
rect 18228 24117 18280 24169
rect 18292 24117 18344 24169
rect 17652 24052 17704 24104
rect 17716 24052 17768 24104
rect 17780 24052 17832 24104
rect 17844 24052 17896 24104
rect 17908 24052 17960 24104
rect 17972 24052 18024 24104
rect 18036 24052 18088 24104
rect 18100 24052 18152 24104
rect 18164 24052 18216 24104
rect 18228 24052 18280 24104
rect 18292 24052 18344 24104
rect 17652 23987 17704 24039
rect 17716 23987 17768 24039
rect 17780 23987 17832 24039
rect 17844 23987 17896 24039
rect 17908 23987 17960 24039
rect 17972 23987 18024 24039
rect 18036 23987 18088 24039
rect 18100 23987 18152 24039
rect 18164 23987 18216 24039
rect 18228 23987 18280 24039
rect 18292 23987 18344 24039
rect 17652 23922 17704 23974
rect 17716 23922 17768 23974
rect 17780 23922 17832 23974
rect 17844 23922 17896 23974
rect 17908 23922 17960 23974
rect 17972 23922 18024 23974
rect 18036 23922 18088 23974
rect 18100 23922 18152 23974
rect 18164 23922 18216 23974
rect 18228 23922 18280 23974
rect 18292 23922 18344 23974
rect 17652 23857 17704 23909
rect 17716 23857 17768 23909
rect 17780 23857 17832 23909
rect 17844 23857 17896 23909
rect 17908 23857 17960 23909
rect 17972 23857 18024 23909
rect 18036 23857 18088 23909
rect 18100 23857 18152 23909
rect 18164 23857 18216 23909
rect 18228 23857 18280 23909
rect 18292 23857 18344 23909
rect 17652 23792 17704 23844
rect 17716 23792 17768 23844
rect 17780 23792 17832 23844
rect 17844 23792 17896 23844
rect 17908 23792 17960 23844
rect 17972 23792 18024 23844
rect 18036 23792 18088 23844
rect 18100 23792 18152 23844
rect 18164 23792 18216 23844
rect 18228 23792 18280 23844
rect 18292 23792 18344 23844
rect 17652 23727 17704 23779
rect 17716 23727 17768 23779
rect 17780 23727 17832 23779
rect 17844 23727 17896 23779
rect 17908 23727 17960 23779
rect 17972 23727 18024 23779
rect 18036 23727 18088 23779
rect 18100 23727 18152 23779
rect 18164 23727 18216 23779
rect 18228 23727 18280 23779
rect 18292 23727 18344 23779
rect 17652 23662 17704 23714
rect 17716 23662 17768 23714
rect 17780 23662 17832 23714
rect 17844 23662 17896 23714
rect 17908 23662 17960 23714
rect 17972 23662 18024 23714
rect 18036 23662 18088 23714
rect 18100 23662 18152 23714
rect 18164 23662 18216 23714
rect 18228 23662 18280 23714
rect 18292 23662 18344 23714
rect 17652 23597 17704 23649
rect 17716 23597 17768 23649
rect 17780 23597 17832 23649
rect 17844 23597 17896 23649
rect 17908 23597 17960 23649
rect 17972 23597 18024 23649
rect 18036 23597 18088 23649
rect 18100 23597 18152 23649
rect 18164 23597 18216 23649
rect 18228 23597 18280 23649
rect 18292 23597 18344 23649
rect 1250 23469 1272 23503
rect 1272 23469 1302 23503
rect 1250 23460 1302 23469
rect 2663 23496 2715 23548
rect 2727 23496 2779 23548
rect 2611 23459 2663 23468
rect 2611 23425 2617 23459
rect 2617 23425 2651 23459
rect 2651 23425 2663 23459
rect 2611 23416 2663 23425
rect 2675 23459 2727 23468
rect 2675 23425 2689 23459
rect 2689 23425 2723 23459
rect 2723 23425 2727 23459
rect 2675 23416 2727 23425
rect 3491 23416 3543 23468
rect 3555 23416 3607 23468
rect 3619 23416 3671 23468
rect 236 22529 288 22581
rect 396 22529 448 22581
rect 236 22465 288 22517
rect 396 22465 448 22517
rect -25 20567 27 20619
rect -25 20503 27 20555
rect 396 20299 448 20351
rect 396 20235 448 20287
rect 927 5001 979 5007
rect 991 5001 1043 5007
rect 927 4967 948 5001
rect 948 4967 979 5001
rect 991 4967 1023 5001
rect 1023 4967 1043 5001
rect 927 4955 979 4967
rect 991 4955 1043 4967
rect -2842 4802 -2790 4854
rect -2778 4802 -2726 4854
rect 1036 4845 1088 4886
rect 1036 4834 1057 4845
rect 1057 4834 1088 4845
rect 1036 4811 1057 4822
rect 1057 4811 1088 4822
rect 1036 4770 1088 4811
rect 956 4710 1008 4762
rect -2922 4643 -2870 4695
rect -2858 4643 -2806 4695
rect 956 4689 1008 4698
rect 956 4655 982 4689
rect 982 4655 1008 4689
rect 956 4646 1008 4655
rect -3088 4589 -3036 4641
rect 796 4579 848 4588
rect -3088 4525 -3036 4577
rect 796 4545 797 4579
rect 797 4545 831 4579
rect 831 4545 848 4579
rect 796 4536 848 4545
rect 796 4472 848 4524
rect -3002 4381 -2950 4433
rect -2938 4381 -2886 4433
rect 876 4423 928 4464
rect 876 4412 907 4423
rect 907 4412 928 4423
rect 876 4389 907 4400
rect 907 4389 928 4400
rect 876 4348 928 4389
rect 796 4288 848 4340
rect 796 4267 848 4276
rect 796 4233 797 4267
rect 797 4233 831 4267
rect 831 4233 848 4267
rect 796 4224 848 4233
<< metal2 >>
tri 3115 26955 3167 27007 se
rect 3167 26955 4197 27007
rect 4249 26955 4261 27007
rect 4313 26955 4319 27007
tri 3093 26933 3115 26955 se
rect 3115 26933 3167 26955
tri 3167 26933 3189 26955 nw
tri 3019 26859 3093 26933 se
tri 3093 26859 3167 26933 nw
tri 2996 26836 3019 26859 se
rect 3019 26836 3070 26859
tri 3070 26836 3093 26859 nw
tri 2945 26785 2996 26836 se
rect 2996 26785 3019 26836
tri 3019 26785 3070 26836 nw
tri 2944 26784 2945 26785 se
rect 2945 26784 3018 26785
tri 3018 26784 3019 26785 nw
tri 2932 26772 2944 26784 se
rect 2944 26772 3006 26784
tri 3006 26772 3018 26784 nw
tri 2880 26720 2932 26772 se
rect 2932 26720 2954 26772
tri 2954 26720 3006 26772 nw
tri 2876 26716 2880 26720 se
rect 2880 26716 2950 26720
tri 2950 26716 2954 26720 nw
rect 2876 26580 2928 26716
tri 2928 26694 2950 26716 nw
tri 4477 26544 4478 26545 se
rect 4478 26544 4862 27929
rect 2876 26516 2928 26528
tri 4443 26510 4477 26544 se
rect 4477 26510 4862 26544
tri 4862 26510 4896 26544 sw
rect 4985 26522 5177 27929
tri 4985 26510 4997 26522 ne
rect 4997 26510 5177 26522
rect 2876 26458 2928 26464
tri 4391 26458 4443 26510 se
rect 4443 26458 4896 26510
tri 4896 26458 4948 26510 sw
tri 4997 26458 5049 26510 ne
rect 5049 26458 5055 26510
rect 5107 26458 5119 26510
rect 5171 26458 5177 26510
rect 5302 26458 5686 27929
rect 5809 26458 6001 27929
rect 6126 26458 6510 27929
rect 6633 27345 6825 27929
rect 6633 27229 6639 27345
rect 6819 27229 6825 27345
tri 4369 26436 4391 26458 se
rect 4391 26455 4948 26458
tri 4948 26455 4951 26458 sw
rect 4391 26436 4951 26455
tri 4951 26436 4970 26455 sw
tri 6614 26436 6633 26455 se
rect 6633 26436 6825 27229
rect 6945 26574 8977 27929
tri 6945 26562 6957 26574 ne
rect 6957 26562 8965 26574
tri 8965 26562 8977 26574 nw
rect 9102 27749 10855 27929
rect 9102 27563 10494 27749
tri 10494 27563 10680 27749 nw
rect 9102 27511 10442 27563
tri 10442 27511 10494 27563 nw
tri 10702 27511 10754 27563 se
rect 10754 27511 10783 27563
rect 10835 27511 10847 27563
rect 10899 27511 10905 27563
tri 6957 26510 7009 26562 ne
rect 7009 26510 7015 26562
rect 7067 26510 7079 26562
rect 7131 26510 7143 26562
rect 7195 26510 7207 26562
rect 7259 26510 7271 26562
rect 7323 26510 8599 26562
rect 8651 26510 8663 26562
rect 8715 26510 8727 26562
rect 8779 26510 8791 26562
rect 8843 26510 8855 26562
rect 8907 26552 8955 26562
tri 8955 26552 8965 26562 nw
rect 8907 26544 8947 26552
tri 8947 26544 8955 26552 nw
rect 8907 26510 8913 26544
tri 8913 26510 8947 26544 nw
tri 9068 26510 9102 26544 se
rect 9102 26510 10431 27511
tri 10431 27500 10442 27511 nw
tri 10691 27500 10702 27511 se
rect 10702 27500 10748 27511
tri 10674 27483 10691 27500 se
rect 10691 27483 10748 27500
tri 10748 27483 10776 27511 nw
tri 10667 27476 10674 27483 se
rect 10674 27476 10719 27483
rect 10667 26836 10719 27476
tri 10719 27454 10748 27483 nw
rect 10820 27431 10826 27483
rect 10878 27431 10890 27483
rect 10942 27432 10980 27483
tri 10980 27432 11031 27483 sw
rect 10942 27431 11031 27432
tri 10954 27406 10979 27431 ne
rect 10667 26772 10719 26784
rect 10667 26714 10719 26720
rect 10979 26552 11031 27431
rect 11131 26575 13100 27929
tri 11131 26562 11144 26575 ne
rect 11144 26574 13100 26575
rect 11144 26562 13088 26574
tri 13088 26562 13100 26574 nw
tri 10431 26510 10467 26546 sw
tri 9058 26500 9068 26510 se
rect 9068 26500 10467 26510
tri 10467 26500 10477 26510 sw
tri 11144 26510 11196 26562 ne
rect 11196 26510 11202 26562
rect 11254 26510 11266 26562
rect 11318 26510 11330 26562
rect 11382 26510 11394 26562
rect 11446 26510 12722 26562
rect 12774 26510 12786 26562
rect 12838 26510 12850 26562
rect 12902 26510 12914 26562
rect 12966 26510 12978 26562
rect 13030 26544 13070 26562
tri 13070 26544 13088 26562 nw
rect 13030 26510 13036 26544
tri 13036 26510 13070 26544 nw
tri 13191 26510 13225 26544 se
rect 13225 26510 15073 27929
rect 15190 26574 17222 27929
tri 15190 26562 15202 26574 ne
rect 15202 26562 17210 26574
tri 17210 26562 17222 26574 nw
tri 15202 26544 15220 26562 ne
rect 15220 26544 15260 26562
tri 15073 26510 15107 26544 sw
tri 15220 26510 15254 26544 ne
rect 15254 26510 15260 26544
rect 15312 26510 15324 26562
rect 15376 26510 15388 26562
rect 15440 26510 15452 26562
rect 15504 26510 15516 26562
rect 15568 26510 16844 26562
rect 16896 26510 16908 26562
rect 16960 26510 16972 26562
rect 17024 26510 17036 26562
rect 17088 26510 17100 26562
rect 17152 26544 17192 26562
tri 17192 26544 17210 26562 nw
rect 17152 26510 17158 26544
tri 17158 26510 17192 26544 nw
tri 17339 26510 17373 26544 se
rect 17373 26510 18369 27929
tri 9046 26488 9058 26500 se
rect 9058 26488 10477 26500
tri 10477 26488 10489 26500 sw
rect 10979 26488 11031 26500
tri 9016 26458 9046 26488 se
rect 9046 26458 10489 26488
tri 10489 26458 10519 26488 sw
tri 9013 26455 9016 26458 se
rect 9016 26455 10519 26458
tri 6825 26436 6844 26455 sw
tri 8994 26436 9013 26455 se
rect 9013 26436 10519 26455
tri 10519 26436 10541 26458 sw
tri 4363 26430 4369 26436 se
rect 4369 26430 4970 26436
rect 3313 26402 4020 26430
tri 4020 26402 4048 26430 sw
tri 4335 26402 4363 26430 se
rect 4363 26402 4970 26430
tri 4970 26402 5004 26436 sw
tri 6580 26402 6614 26436 se
rect 6614 26402 6844 26436
tri 6844 26402 6878 26436 sw
tri 8960 26402 8994 26436 se
rect 8994 26430 10541 26436
tri 10541 26430 10547 26436 sw
rect 10979 26430 11031 26436
tri 13111 26430 13191 26510 se
rect 13191 26430 15107 26510
tri 15107 26430 15187 26510 sw
tri 17259 26430 17339 26510 se
rect 17339 26430 18369 26510
rect 8994 26402 10547 26430
tri 10547 26402 10575 26430 sw
tri 13083 26402 13111 26430 se
rect 13111 26402 15187 26430
tri 15187 26402 15215 26430 sw
tri 17231 26402 17259 26430 se
rect 17259 26402 18369 26430
rect 3313 26090 18369 26402
tri 17485 26035 17540 26090 ne
rect 17540 26035 18369 26090
tri 17540 25982 17593 26035 ne
rect 17593 25982 17652 26035
rect 4160 25946 17440 25982
tri 17440 25946 17476 25982 sw
tri 17593 25946 17629 25982 ne
rect 4160 25849 17476 25946
tri 17476 25849 17573 25946 sw
tri 620 25097 650 25127 se
rect 650 25097 666 25149
rect 718 25097 730 25149
rect 782 25097 788 25149
tri 576 25053 620 25097 se
rect 620 25053 650 25097
tri 650 25053 694 25097 nw
tri 502 24979 576 25053 se
tri 576 24979 650 25053 nw
tri 428 24905 502 24979 se
tri 502 24905 576 24979 nw
tri 410 24887 428 24905 se
rect 428 24887 484 24905
tri 484 24887 502 24905 nw
tri 346 23284 410 23348 se
rect 410 23326 462 24887
tri 462 24865 484 24887 nw
rect 4160 24435 17573 25849
tri 8064 24429 8070 24435 ne
rect 8070 24429 8673 24435
tri 8673 24429 8679 24435 nw
tri 8879 24429 8885 24435 ne
rect 8885 24429 11969 24435
tri 11969 24429 11975 24435 nw
tri 12175 24429 12181 24435 ne
rect 12181 24429 12793 24435
tri 12793 24429 12799 24435 nw
tri 12999 24429 13005 24435 ne
rect 13005 24429 13617 24435
tri 13617 24429 13623 24435 nw
tri 13823 24429 13829 24435 ne
rect 13829 24429 14441 24435
tri 14441 24429 14447 24435 nw
tri 14647 24429 14653 24435 ne
rect 14653 24429 15265 24435
tri 15265 24429 15271 24435 nw
tri 15471 24429 15477 24435 ne
rect 15477 24429 16089 24435
tri 16089 24429 16095 24435 nw
tri 16295 24429 16301 24435 ne
rect 16301 24429 16913 24435
tri 16913 24429 16919 24435 nw
tri 17119 24429 17125 24435 ne
rect 17125 24429 17573 24435
tri 8070 24377 8122 24429 ne
rect 8122 24377 8621 24429
tri 8621 24377 8673 24429 nw
tri 8885 24377 8937 24429 ne
rect 8937 24399 11939 24429
tri 11939 24399 11969 24429 nw
tri 12181 24399 12211 24429 ne
rect 12211 24399 12741 24429
rect 8937 24377 9483 24399
tri 9483 24377 9505 24399 nw
tri 11351 24377 11373 24399 ne
rect 11373 24377 11917 24399
tri 11917 24377 11939 24399 nw
tri 12211 24377 12233 24399 ne
rect 12233 24377 12741 24399
tri 12741 24377 12793 24429 nw
tri 13005 24377 13057 24429 ne
rect 13057 24377 13565 24429
tri 13565 24377 13617 24429 nw
tri 13829 24377 13881 24429 ne
rect 13881 24377 14389 24429
tri 14389 24377 14441 24429 nw
tri 14653 24377 14705 24429 ne
rect 14705 24377 15213 24429
tri 15213 24377 15265 24429 nw
tri 15477 24377 15529 24429 ne
rect 15529 24377 16037 24429
tri 16037 24377 16089 24429 nw
tri 16301 24377 16353 24429 ne
rect 16353 24377 16861 24429
tri 16861 24377 16913 24429 nw
tri 17125 24377 17177 24429 ne
rect 17177 24377 17573 24429
tri 8122 24364 8135 24377 ne
rect 8135 24364 8608 24377
tri 8608 24364 8621 24377 nw
tri 8937 24364 8950 24377 ne
rect 8950 24364 9470 24377
tri 9470 24364 9483 24377 nw
tri 11373 24364 11386 24377 ne
rect 11386 24364 11904 24377
tri 11904 24364 11917 24377 nw
tri 12233 24364 12246 24377 ne
rect 12246 24364 12728 24377
tri 12728 24364 12741 24377 nw
tri 13057 24364 13070 24377 ne
rect 13070 24364 13552 24377
tri 13552 24364 13565 24377 nw
tri 13881 24364 13894 24377 ne
rect 13894 24364 14376 24377
tri 14376 24364 14389 24377 nw
tri 14705 24364 14718 24377 ne
rect 14718 24364 15200 24377
tri 15200 24364 15213 24377 nw
tri 15529 24364 15542 24377 ne
rect 15542 24364 16024 24377
tri 16024 24364 16037 24377 nw
tri 16353 24364 16366 24377 ne
rect 16366 24364 16848 24377
tri 16848 24364 16861 24377 nw
tri 17177 24364 17190 24377 ne
rect 17190 24364 17573 24377
tri 8135 24312 8187 24364 ne
rect 8187 24312 8556 24364
tri 8556 24312 8608 24364 nw
tri 8950 24312 9002 24364 ne
rect 9002 24312 9418 24364
tri 9418 24312 9470 24364 nw
tri 11386 24312 11438 24364 ne
rect 11438 24312 11852 24364
tri 11852 24312 11904 24364 nw
tri 12246 24312 12298 24364 ne
rect 12298 24312 12676 24364
tri 12676 24312 12728 24364 nw
tri 13070 24312 13122 24364 ne
rect 13122 24312 13500 24364
tri 13500 24312 13552 24364 nw
tri 13894 24312 13946 24364 ne
rect 13946 24312 14324 24364
tri 14324 24312 14376 24364 nw
tri 14718 24312 14770 24364 ne
rect 14770 24312 15148 24364
tri 15148 24312 15200 24364 nw
tri 15542 24312 15594 24364 ne
rect 15594 24312 15972 24364
tri 15972 24312 16024 24364 nw
tri 16366 24312 16418 24364 ne
rect 16418 24312 16796 24364
tri 16796 24312 16848 24364 nw
tri 17190 24312 17242 24364 ne
rect 17242 24312 17573 24364
tri 8187 24301 8198 24312 ne
rect 8198 24301 8543 24312
tri 502 23326 529 23353 se
rect 529 23331 581 24301
rect 529 23326 534 23331
rect 410 23286 422 23326
tri 422 23286 462 23326 nw
tri 462 23286 502 23326 se
rect 502 23286 534 23326
rect 410 23284 420 23286
tri 420 23284 422 23286 nw
tri 460 23284 462 23286 se
rect 462 23284 534 23286
tri 534 23284 581 23331 nw
tri 341 23279 346 23284 se
rect 346 23279 415 23284
tri 415 23279 420 23284 nw
tri 455 23279 460 23284 se
rect 460 23279 529 23284
tri 529 23279 534 23284 nw
tri 604 23279 609 23284 se
rect 609 23279 661 24301
tri 336 23274 341 23279 se
rect 341 23274 410 23279
tri 410 23274 415 23279 nw
tri 450 23274 455 23279 se
rect 455 23274 498 23279
tri 310 23248 336 23274 se
rect 336 23248 384 23274
tri 384 23248 410 23274 nw
tri 424 23248 450 23274 se
rect 450 23248 498 23274
tri 498 23248 529 23279 nw
tri 573 23248 604 23279 se
rect 604 23262 661 23279
rect 604 23251 650 23262
tri 650 23251 661 23262 nw
rect 604 23248 647 23251
tri 647 23248 650 23251 nw
tri 687 23248 690 23251 se
rect 690 23248 742 24301
tri 267 23205 310 23248 se
rect 310 23234 370 23248
tri 370 23234 384 23248 nw
tri 410 23234 424 23248 se
rect 424 23234 460 23248
rect 310 23205 341 23234
tri 341 23205 370 23234 nw
tri 381 23205 410 23234 se
rect 410 23210 460 23234
tri 460 23210 498 23248 nw
tri 535 23210 573 23248 se
rect 573 23217 616 23248
tri 616 23217 647 23248 nw
tri 656 23217 687 23248 se
rect 687 23229 742 23248
rect 687 23217 730 23229
tri 730 23217 742 23229 nw
rect 573 23210 609 23217
tri 609 23210 616 23217 nw
tri 649 23210 656 23217 se
rect 656 23210 690 23217
rect 410 23205 455 23210
tri 455 23205 460 23210 nw
tri 530 23205 535 23210 se
rect 535 23205 576 23210
tri 262 23200 267 23205 se
rect 267 23200 336 23205
tri 336 23200 341 23205 nw
tri 376 23200 381 23205 se
rect 381 23200 450 23205
tri 450 23200 455 23205 nw
tri 525 23200 530 23205 se
rect 530 23200 576 23205
tri 193 23131 262 23200 se
rect 262 23160 296 23200
tri 296 23160 336 23200 nw
tri 336 23160 376 23200 se
rect 376 23160 386 23200
rect 262 23131 267 23160
tri 267 23131 296 23160 nw
tri 307 23131 336 23160 se
rect 336 23136 386 23160
tri 386 23136 450 23200 nw
tri 461 23136 525 23200 se
rect 525 23177 576 23200
tri 576 23177 609 23210 nw
tri 616 23177 649 23210 se
rect 649 23177 690 23210
tri 690 23177 730 23217 nw
tri 730 23177 770 23217 se
rect 770 23189 822 24301
rect 770 23177 810 23189
tri 810 23177 822 23189 nw
rect 525 23143 542 23177
tri 542 23143 576 23177 nw
tri 582 23143 616 23177 se
rect 616 23143 650 23177
rect 525 23136 535 23143
tri 535 23136 542 23143 nw
tri 575 23136 582 23143 se
rect 582 23137 650 23143
tri 650 23137 690 23177 nw
tri 690 23137 730 23177 se
rect 730 23143 776 23177
tri 776 23143 810 23177 nw
tri 816 23143 850 23177 se
rect 850 23155 902 24301
rect 850 23143 884 23155
rect 730 23137 770 23143
tri 770 23137 776 23143 nw
tri 810 23137 816 23143 se
rect 816 23137 884 23143
tri 884 23137 902 23155 nw
rect 582 23136 616 23137
rect 336 23131 381 23136
tri 381 23131 386 23136 nw
tri 456 23131 461 23136 se
rect 461 23131 502 23136
tri 188 23126 193 23131 se
rect 193 23126 262 23131
tri 262 23126 267 23131 nw
tri 302 23126 307 23131 se
rect 307 23126 376 23131
tri 376 23126 381 23131 nw
tri 451 23126 456 23131 se
rect 456 23126 502 23131
tri 114 23052 188 23126 se
rect 188 23086 222 23126
tri 222 23086 262 23126 nw
tri 262 23086 302 23126 se
rect 302 23086 312 23126
tri 188 23052 222 23086 nw
tri 235 23059 262 23086 se
rect 262 23062 312 23086
tri 312 23062 376 23126 nw
tri 387 23062 451 23126 se
rect 451 23103 502 23126
tri 502 23103 535 23136 nw
tri 542 23103 575 23136 se
rect 575 23103 616 23136
tri 616 23103 650 23137 nw
tri 656 23103 690 23137 se
rect 690 23103 736 23137
tri 736 23103 770 23137 nw
tri 776 23103 810 23137 se
rect 810 23109 856 23137
tri 856 23109 884 23137 nw
tri 902 23109 930 23137 se
rect 930 23115 982 24301
rect 930 23109 970 23115
rect 810 23103 850 23109
tri 850 23103 856 23109 nw
tri 896 23103 902 23109 se
rect 902 23103 970 23109
tri 970 23103 982 23115 nw
rect 451 23069 468 23103
tri 468 23069 502 23103 nw
tri 508 23069 542 23103 se
rect 542 23097 610 23103
tri 610 23097 616 23103 nw
tri 650 23097 656 23103 se
rect 656 23097 702 23103
rect 542 23069 570 23097
rect 451 23062 461 23069
tri 461 23062 468 23069 nw
tri 501 23062 508 23069 se
rect 508 23062 570 23069
rect 262 23059 309 23062
tri 309 23059 312 23062 nw
tri 384 23059 387 23062 se
rect 387 23059 428 23062
tri 76 23014 114 23052 se
rect 114 23014 150 23052
tri 150 23014 188 23052 nw
rect -166 22599 -38 22753
tri 42 21090 76 21124 se
rect 76 21102 128 23014
tri 128 22992 150 23014 nw
tri 161 22660 235 22734 se
rect 235 22712 287 23059
tri 287 23037 309 23059 nw
tri 362 23037 384 23059 se
rect 384 23037 428 23059
tri 235 22660 287 22712 nw
tri 316 22991 362 23037 se
rect 362 23029 428 23037
tri 428 23029 461 23062 nw
tri 468 23029 501 23062 se
rect 501 23057 570 23062
tri 570 23057 610 23097 nw
tri 610 23057 650 23097 se
rect 650 23069 702 23097
tri 702 23069 736 23103 nw
tri 742 23069 776 23103 se
rect 776 23069 810 23103
rect 650 23057 690 23069
tri 690 23057 702 23069 nw
tri 730 23057 742 23069 se
rect 742 23063 810 23069
tri 810 23063 850 23103 nw
tri 856 23063 896 23103 se
rect 896 23079 946 23103
tri 946 23079 970 23103 nw
tri 986 23079 1010 23103 se
rect 1010 23091 1062 24301
tri 8198 24299 8200 24301 ne
rect 8200 24299 8543 24301
tri 8543 24299 8556 24312 nw
tri 9002 24299 9015 24312 ne
rect 9015 24299 9405 24312
tri 9405 24299 9418 24312 nw
tri 11438 24299 11451 24312 ne
rect 11451 24299 11839 24312
tri 11839 24299 11852 24312 nw
tri 12298 24299 12311 24312 ne
rect 12311 24299 12663 24312
tri 12663 24299 12676 24312 nw
tri 13122 24299 13135 24312 ne
rect 13135 24299 13487 24312
tri 13487 24299 13500 24312 nw
tri 13946 24299 13959 24312 ne
rect 13959 24299 14311 24312
tri 14311 24299 14324 24312 nw
tri 14770 24299 14783 24312 ne
rect 14783 24299 15135 24312
tri 15135 24299 15148 24312 nw
tri 15594 24299 15607 24312 ne
rect 15607 24299 15959 24312
tri 15959 24299 15972 24312 nw
tri 16418 24299 16431 24312 ne
rect 16431 24299 16783 24312
tri 16783 24299 16796 24312 nw
tri 17242 24299 17255 24312 ne
rect 17255 24299 17573 24312
tri 4373 24268 4404 24299 se
rect 4404 24268 4815 24299
tri 4815 24268 4846 24299 sw
tri 5296 24268 5327 24299 se
rect 5327 24268 5639 24299
tri 5639 24268 5670 24299 sw
tri 6120 24268 6151 24299 se
rect 6151 24268 6463 24299
tri 6463 24268 6494 24299 sw
tri 6944 24268 6975 24299 se
rect 6975 24268 7287 24299
tri 7287 24268 7318 24299 sw
tri 7768 24268 7799 24299 se
rect 7799 24291 8111 24299
tri 8111 24291 8119 24299 sw
tri 8200 24291 8208 24299 ne
rect 7799 24268 8119 24291
tri 8119 24268 8142 24291 sw
rect 1010 23079 1050 23091
tri 1050 23079 1062 23091 nw
rect 1090 24246 1142 24252
rect 1090 24182 1142 24194
rect 1090 23998 1142 24130
rect 4373 24216 4508 24268
rect 4560 24216 4572 24268
rect 4624 24216 4636 24268
rect 4688 24216 4700 24268
rect 4752 24216 4764 24268
rect 4816 24261 4846 24268
tri 4846 24261 4853 24268 sw
rect 4816 24216 4853 24261
rect 1090 23934 1142 23946
rect 896 23063 930 23079
tri 930 23063 946 23079 nw
tri 970 23063 986 23079 se
rect 986 23063 1016 23079
rect 742 23057 782 23063
rect 501 23029 542 23057
tri 542 23029 570 23057 nw
tri 582 23029 610 23057 se
rect 610 23029 662 23057
tri 662 23029 690 23057 nw
tri 702 23029 730 23057 se
rect 730 23035 782 23057
tri 782 23035 810 23063 nw
tri 828 23035 856 23063 se
rect 856 23039 906 23063
tri 906 23039 930 23063 nw
tri 946 23039 970 23063 se
rect 970 23045 1016 23063
tri 1016 23045 1050 23079 nw
tri 1056 23045 1090 23079 se
rect 1090 23057 1142 23882
rect 1090 23045 1130 23057
tri 1130 23045 1142 23057 nw
rect 1170 24122 1222 24128
rect 1170 24058 1222 24070
rect 1170 23927 1222 24006
tri 1222 23927 1247 23952 sw
rect 1170 23922 1319 23927
tri 1319 23922 1324 23927 sw
rect 1170 23909 1324 23922
tri 1324 23909 1337 23922 sw
rect 1170 23890 1337 23909
tri 1337 23890 1356 23909 sw
rect 4373 23890 4853 24216
rect 5296 24216 5332 24268
rect 5384 24216 5396 24268
rect 5448 24216 5460 24268
rect 5512 24216 5524 24268
rect 5576 24216 5588 24268
rect 5640 24261 5670 24268
tri 5670 24261 5677 24268 sw
rect 5640 24216 5677 24261
rect 5296 23890 5677 24216
rect 6120 24216 6156 24268
rect 6208 24216 6220 24268
rect 6272 24216 6284 24268
rect 6336 24216 6348 24268
rect 6400 24216 6412 24268
rect 6464 24261 6494 24268
tri 6494 24261 6501 24268 sw
rect 6464 24216 6501 24261
rect 6120 23890 6501 24216
rect 6944 24216 6980 24268
rect 7032 24216 7044 24268
rect 7096 24216 7108 24268
rect 7160 24216 7172 24268
rect 7224 24216 7236 24268
rect 7288 24261 7318 24268
tri 7318 24261 7325 24268 sw
rect 7288 24216 7325 24261
rect 6944 23890 7325 24216
rect 7768 24216 7804 24268
rect 7856 24216 7868 24268
rect 7920 24216 7932 24268
rect 7984 24216 7996 24268
rect 8048 24216 8060 24268
rect 8112 24261 8142 24268
tri 8142 24261 8149 24268 sw
rect 8112 24216 8149 24261
rect 7768 23890 8149 24216
rect 1170 23875 1356 23890
rect 1170 23857 1229 23875
tri 1229 23857 1247 23875 nw
tri 1297 23857 1315 23875 ne
rect 1315 23857 1356 23875
tri 1356 23857 1389 23890 sw
rect 1170 23856 1228 23857
tri 1228 23856 1229 23857 nw
tri 1315 23856 1316 23857 ne
rect 1316 23856 1389 23857
tri 1389 23856 1390 23857 sw
rect 970 23039 1010 23045
tri 1010 23039 1016 23045 nw
tri 1050 23039 1056 23045 se
rect 1056 23039 1096 23045
rect 856 23035 882 23039
rect 730 23029 776 23035
tri 776 23029 782 23035 nw
tri 822 23029 828 23035 se
rect 828 23029 882 23035
rect 362 22997 396 23029
tri 396 22997 428 23029 nw
tri 436 22997 468 23029 se
rect 468 23017 530 23029
tri 530 23017 542 23029 nw
tri 570 23017 582 23029 se
rect 582 23017 628 23029
rect 468 22997 490 23017
rect 362 22991 390 22997
tri 390 22991 396 22997 nw
tri 430 22991 436 22997 se
rect 436 22991 490 22997
rect 76 21090 116 21102
tri 116 21090 128 21102 nw
tri 156 22655 161 22660 se
rect 161 22655 230 22660
tri 230 22655 235 22660 nw
tri 2 21050 42 21090 se
rect 42 21062 88 21090
tri 88 21062 116 21090 nw
tri 128 21062 156 21090 se
rect 156 21068 208 22655
tri 208 22633 230 22655 nw
rect 156 21062 196 21068
rect 42 21050 76 21062
tri 76 21050 88 21062 nw
tri 116 21050 128 21062 se
rect 128 21056 196 21062
tri 196 21056 208 21068 nw
rect 236 22581 288 22587
rect 236 22517 288 22529
rect 128 21050 187 21056
tri -25 21023 2 21050 se
rect 2 21023 49 21050
tri 49 21023 76 21050 nw
tri 89 21023 116 21050 se
rect 116 21047 187 21050
tri 187 21047 196 21056 nw
tri 227 21047 236 21056 se
rect 236 21047 288 22465
rect 116 21023 156 21047
rect -25 21016 42 21023
tri 42 21016 49 21023 nw
tri 82 21016 89 21023 se
rect 89 21016 156 21023
tri 156 21016 187 21047 nw
tri 214 21034 227 21047 se
rect 227 21034 288 21047
tri 196 21016 214 21034 se
rect 214 21022 276 21034
tri 276 21022 288 21034 nw
rect 214 21016 270 21022
tri 270 21016 276 21022 nw
tri 310 21016 316 21022 se
rect 316 21016 368 22991
tri 368 22969 390 22991 nw
tri 408 22969 430 22991 se
rect 430 22977 490 22991
tri 490 22977 530 23017 nw
tri 530 22977 570 23017 se
rect 570 22995 628 23017
tri 628 22995 662 23029 nw
tri 668 22995 702 23029 se
rect 702 22995 736 23029
rect 570 22977 610 22995
tri 610 22977 628 22995 nw
tri 650 22977 668 22995 se
rect 668 22989 736 22995
tri 736 22989 776 23029 nw
tri 782 22989 822 23029 se
rect 822 23015 882 23029
tri 882 23015 906 23039 nw
tri 922 23015 946 23039 se
rect 946 23015 976 23039
rect 822 22989 856 23015
tri 856 22989 882 23015 nw
tri 896 22989 922 23015 se
rect 922 23005 976 23015
tri 976 23005 1010 23039 nw
tri 1016 23005 1050 23039 se
rect 1050 23011 1096 23039
tri 1096 23011 1130 23045 nw
tri 1136 23011 1170 23045 se
rect 1170 23023 1222 23856
tri 1222 23850 1228 23856 nw
tri 1316 23853 1319 23856 ne
rect 1319 23853 1390 23856
tri 1319 23850 1322 23853 ne
rect 1322 23850 1390 23853
tri 1322 23844 1328 23850 ne
rect 1328 23844 1390 23850
tri 1390 23844 1402 23856 sw
tri 1328 23830 1342 23844 ne
rect 1342 23830 1402 23844
tri 1402 23830 1416 23844 sw
rect 1170 23011 1210 23023
tri 1210 23011 1222 23023 nw
rect 1250 23824 1302 23830
tri 1342 23792 1380 23830 ne
rect 1380 23792 1416 23830
tri 1416 23792 1454 23830 sw
tri 1380 23788 1384 23792 ne
rect 1384 23788 1454 23792
tri 1454 23788 1458 23792 sw
tri 1384 23782 1390 23788 ne
rect 1390 23782 1458 23788
tri 1458 23782 1464 23788 sw
rect 1250 23760 1302 23772
tri 1390 23736 1436 23782 ne
rect 1436 23736 1464 23782
tri 1464 23736 1510 23782 sw
rect 2657 23736 2663 23788
rect 2715 23736 2727 23788
rect 2779 23736 6998 23788
rect 7050 23736 7062 23788
rect 7114 23736 7120 23788
tri 7782 23736 7834 23788 se
rect 7834 23736 7904 23788
rect 7956 23736 7968 23788
rect 8020 23736 8026 23788
tri 1436 23733 1439 23736 ne
rect 1439 23733 1510 23736
tri 1510 23733 1513 23736 sw
tri 7779 23733 7782 23736 se
rect 7782 23733 7853 23736
tri 7853 23733 7856 23736 nw
tri 1439 23727 1445 23733 ne
rect 1445 23727 1513 23733
tri 1513 23727 1519 23733 sw
tri 7773 23727 7779 23733 se
rect 7779 23727 7847 23733
tri 7847 23727 7853 23733 nw
tri 1445 23714 1458 23727 ne
rect 1458 23714 1519 23727
tri 1519 23714 1532 23727 sw
tri 7760 23714 7773 23727 se
rect 7773 23714 7834 23727
tri 7834 23714 7847 23727 nw
tri 1458 23708 1464 23714 ne
rect 1464 23710 1532 23714
tri 1532 23710 1536 23714 sw
tri 7756 23710 7760 23714 se
rect 7760 23710 7830 23714
tri 7830 23710 7834 23714 nw
rect 1464 23708 1536 23710
tri 1536 23708 1538 23710 sw
tri 7754 23708 7756 23710 se
rect 7756 23708 7828 23710
tri 7828 23708 7830 23710 nw
rect 1250 23576 1302 23708
tri 1464 23706 1466 23708 ne
rect 1466 23706 4223 23708
rect 1250 23512 1302 23524
rect 1050 23005 1090 23011
tri 1090 23005 1096 23011 nw
tri 1130 23005 1136 23011 se
rect 1136 23005 1204 23011
tri 1204 23005 1210 23011 nw
tri 1244 23005 1250 23011 se
rect 1250 23005 1302 23460
rect 922 22989 946 23005
rect 668 22977 708 22989
rect 430 22969 476 22977
tri 396 22957 408 22969 se
rect 408 22963 476 22969
tri 476 22963 490 22977 nw
tri 516 22963 530 22977 se
rect 530 22963 588 22977
rect 408 22957 470 22963
tri 470 22957 476 22963 nw
tri 510 22957 516 22963 se
rect 516 22957 588 22963
rect 396 22581 448 22957
tri 448 22935 470 22957 nw
tri 488 22935 510 22957 se
rect 510 22955 588 22957
tri 588 22955 610 22977 nw
tri 628 22955 650 22977 se
rect 650 22961 708 22977
tri 708 22961 736 22989 nw
tri 754 22961 782 22989 se
rect 782 22975 842 22989
tri 842 22975 856 22989 nw
tri 882 22975 896 22989 se
rect 896 22975 946 22989
tri 946 22975 976 23005 nw
tri 986 22975 1016 23005 se
rect 1016 22975 1056 23005
rect 782 22961 818 22975
rect 650 22955 702 22961
tri 702 22955 708 22961 nw
tri 748 22955 754 22961 se
rect 754 22955 818 22961
rect 510 22935 556 22955
rect 396 22517 448 22529
rect 396 22459 448 22465
tri 476 22923 488 22935 se
rect 488 22923 556 22935
tri 556 22923 588 22955 nw
tri 596 22923 628 22955 se
rect 628 22923 662 22955
rect 476 22902 535 22923
tri 535 22902 556 22923 nw
tri 575 22902 596 22923 se
rect 596 22915 662 22923
tri 662 22915 702 22955 nw
tri 708 22915 748 22955 se
rect 748 22951 818 22955
tri 818 22951 842 22975 nw
tri 858 22951 882 22975 se
rect 882 22971 942 22975
tri 942 22971 946 22975 nw
tri 982 22971 986 22975 se
rect 986 22971 1056 22975
tri 1056 22971 1090 23005 nw
tri 1096 22971 1130 23005 se
rect 1130 22983 1182 23005
tri 1182 22983 1204 23005 nw
tri 1222 22983 1244 23005 se
rect 1244 22989 1302 23005
rect 1244 22983 1290 22989
rect 1130 22971 1170 22983
tri 1170 22971 1182 22983 nw
tri 1210 22971 1222 22983 se
rect 1222 22977 1290 22983
tri 1290 22977 1302 22989 nw
rect 1330 23700 1382 23706
tri 1466 23665 1507 23706 ne
rect 1507 23665 4223 23706
tri 1382 23656 1391 23665 sw
tri 1507 23656 1516 23665 ne
rect 1516 23656 4223 23665
rect 4275 23656 4287 23708
rect 4339 23656 4345 23708
tri 7741 23695 7754 23708 se
rect 7754 23695 7815 23708
tri 7815 23695 7828 23708 nw
tri 7707 23661 7741 23695 se
rect 7741 23661 7781 23695
tri 7781 23661 7815 23695 nw
tri 7702 23656 7707 23661 se
rect 7707 23656 7776 23661
tri 7776 23656 7781 23661 nw
rect 1382 23648 1391 23656
rect 1330 23636 1391 23648
tri 1391 23636 1411 23656 sw
tri 7686 23640 7702 23656 se
rect 7702 23640 7760 23656
tri 7760 23640 7776 23656 nw
tri 7682 23636 7686 23640 se
rect 7686 23636 7756 23640
tri 7756 23636 7760 23640 nw
rect 1382 23628 1411 23636
tri 1411 23628 1419 23636 sw
tri 7674 23628 7682 23636 se
rect 7682 23628 7748 23636
tri 7748 23628 7756 23636 nw
rect 1382 23584 4223 23628
rect 1330 23576 4223 23584
rect 4275 23576 4287 23628
rect 4339 23576 4345 23628
tri 4419 23609 4438 23628 se
rect 4438 23609 7729 23628
tri 7729 23609 7748 23628 nw
tri 4410 23600 4419 23609 se
rect 4419 23600 7720 23609
tri 7720 23600 7729 23609 nw
tri 4388 23578 4410 23600 se
rect 4410 23578 7698 23600
tri 7698 23578 7720 23600 nw
tri 4386 23576 4388 23578 se
rect 4388 23576 7696 23578
tri 7696 23576 7698 23578 nw
rect 1222 22971 1256 22977
rect 882 22951 902 22971
rect 748 22915 782 22951
tri 782 22915 818 22951 nw
tri 822 22915 858 22951 se
rect 858 22931 902 22951
tri 902 22931 942 22971 nw
tri 942 22931 982 22971 se
rect 982 22937 1022 22971
tri 1022 22937 1056 22971 nw
tri 1062 22937 1096 22971 se
rect 1096 22937 1136 22971
tri 1136 22937 1170 22971 nw
tri 1176 22937 1210 22971 se
rect 1210 22943 1256 22971
tri 1256 22943 1290 22977 nw
tri 1296 22943 1330 22977 se
rect 1330 22955 1382 23576
tri 1382 23563 1395 23576 nw
tri 4373 23563 4386 23576 se
rect 4386 23563 4445 23576
tri 4371 23561 4373 23563 se
rect 4373 23561 4445 23563
tri 4445 23561 4460 23576 nw
tri 4364 23554 4371 23561 se
rect 4371 23554 4438 23561
tri 4438 23554 4445 23561 nw
tri 4358 23548 4364 23554 se
rect 4364 23548 4432 23554
tri 4432 23548 4438 23554 nw
rect 2657 23496 2663 23548
rect 2715 23496 2727 23548
rect 2779 23496 4380 23548
tri 4380 23496 4432 23548 nw
rect 2605 23416 2611 23468
rect 2663 23416 2675 23468
rect 2727 23416 3491 23468
rect 3543 23416 3555 23468
rect 3607 23416 3619 23468
rect 3671 23416 3677 23468
rect 1210 22937 1250 22943
tri 1250 22937 1256 22943 nw
tri 1290 22937 1296 22943 se
rect 1296 22937 1330 22943
rect 982 22931 1016 22937
tri 1016 22931 1022 22937 nw
tri 1056 22931 1062 22937 se
rect 1062 22931 1130 22937
tri 1130 22931 1136 22937 nw
tri 1170 22931 1176 22937 se
rect 1176 22931 1216 22937
rect 858 22915 882 22931
rect 596 22902 649 22915
tri 649 22902 662 22915 nw
tri 695 22902 708 22915 se
rect 708 22911 778 22915
tri 778 22911 782 22915 nw
tri 818 22911 822 22915 se
rect 822 22911 882 22915
tri 882 22911 902 22931 nw
tri 922 22911 942 22931 se
rect 942 22911 987 22931
rect 708 22902 769 22911
tri 769 22902 778 22911 nw
tri 809 22902 818 22911 se
rect 818 22902 873 22911
tri 873 22902 882 22911 nw
tri 913 22902 922 22911 se
rect 922 22902 987 22911
tri 987 22902 1016 22931 nw
tri 1027 22902 1056 22931 se
rect 1056 22902 1101 22931
tri 1101 22902 1130 22931 nw
tri 1141 22902 1170 22931 se
rect 1170 22903 1216 22931
tri 1216 22903 1250 22937 nw
tri 1256 22903 1290 22937 se
rect 1290 22903 1330 22937
tri 1330 22903 1382 22955 nw
rect 1170 22902 1215 22903
tri 1215 22902 1216 22903 nw
tri 1255 22902 1256 22903 se
rect 1256 22902 1329 22903
tri 1329 22902 1330 22903 nw
rect -25 21010 36 21016
tri 36 21010 42 21016 nw
tri 76 21010 82 21016 se
rect 82 21010 147 21016
rect -25 20619 27 21010
tri 27 21001 36 21010 nw
tri 67 21001 76 21010 se
rect 76 21007 147 21010
tri 147 21007 156 21016 nw
tri 187 21007 196 21016 se
rect 196 21007 261 21016
tri 261 21007 270 21016 nw
tri 301 21007 310 21016 se
rect 310 21007 368 21016
rect 76 21001 135 21007
rect -25 20555 27 20567
rect -25 20497 27 20503
tri 55 20989 67 21001 se
rect 67 20995 135 21001
tri 135 20995 147 21007 nw
tri 175 20995 187 21007 se
rect 187 20995 243 21007
rect 67 20989 129 20995
tri 129 20989 135 20995 nw
tri 169 20989 175 20995 se
rect 175 20989 243 20995
tri 243 20989 261 21007 nw
tri 283 20989 301 21007 se
rect 301 21000 368 21007
rect 301 20989 316 21000
rect 55 20374 107 20989
tri 107 20967 129 20989 nw
tri 147 20967 169 20989 se
rect 169 20967 221 20989
tri 221 20967 243 20989 nw
tri 261 20967 283 20989 se
rect 283 20967 316 20989
tri 135 20955 147 20967 se
rect 147 20955 202 20967
rect 135 20948 202 20955
tri 202 20948 221 20967 nw
tri 242 20948 261 20967 se
rect 261 20948 316 20967
tri 316 20948 368 21000 nw
rect 135 20409 187 20948
tri 187 20933 202 20948 nw
tri 227 20933 242 20948 se
rect 242 20933 289 20948
tri 215 20921 227 20933 se
rect 227 20921 289 20933
tri 289 20921 316 20948 nw
rect 215 20443 267 20921
tri 267 20899 289 20921 nw
tri 267 20443 289 20465 sw
tri 215 20431 227 20443 ne
rect 227 20431 289 20443
tri 135 20404 140 20409 ne
rect 140 20404 187 20409
tri 187 20404 214 20431 sw
tri 227 20404 254 20431 ne
rect 254 20416 289 20431
tri 289 20416 316 20443 sw
rect 254 20404 316 20416
tri 140 20396 148 20404 ne
rect 148 20396 214 20404
tri 214 20396 222 20404 sw
tri 254 20396 262 20404 ne
rect 262 20396 316 20404
tri 107 20374 129 20396 sw
tri 148 20374 170 20396 ne
rect 170 20374 222 20396
tri 222 20374 244 20396 sw
tri 262 20374 284 20396 ne
rect 284 20374 316 20396
tri 55 20357 72 20374 ne
rect 72 20368 129 20374
tri 129 20368 135 20374 sw
tri 170 20368 176 20374 ne
rect 176 20370 244 20374
tri 244 20370 248 20374 sw
tri 284 20370 288 20374 ne
rect 288 20370 316 20374
rect 176 20369 248 20370
tri 248 20369 249 20370 sw
tri 288 20369 289 20370 ne
rect 289 20369 316 20370
tri 316 20369 363 20416 sw
rect 176 20368 249 20369
rect 72 20357 135 20368
tri 135 20357 146 20368 sw
tri 176 20357 187 20368 ne
rect 187 20357 249 20368
tri 249 20357 261 20369 sw
tri 289 20357 301 20369 ne
rect 301 20364 363 20369
tri 363 20364 368 20369 sw
rect 301 20357 368 20364
tri 72 20351 78 20357 ne
rect 78 20351 146 20357
tri 146 20351 152 20357 sw
tri 187 20351 193 20357 ne
rect 193 20351 261 20357
tri 261 20351 267 20357 sw
tri 301 20351 307 20357 ne
rect 307 20351 368 20357
tri 78 20300 129 20351 ne
rect 129 20347 152 20351
tri 152 20347 156 20351 sw
tri 193 20347 197 20351 ne
rect 197 20347 267 20351
tri 267 20347 271 20351 sw
tri 307 20347 311 20351 ne
rect 311 20347 368 20351
rect 129 20330 156 20347
tri 156 20330 173 20347 sw
tri 197 20330 214 20347 ne
rect 214 20342 271 20347
tri 271 20342 276 20347 sw
tri 311 20342 316 20347 ne
rect 214 20330 276 20342
tri 276 20330 288 20342 sw
rect 129 20300 173 20330
tri 173 20300 203 20330 sw
tri 214 20308 236 20330 ne
tri 129 20299 130 20300 ne
rect 130 20299 203 20300
tri 203 20299 204 20300 sw
tri 130 20287 142 20299 ne
rect 142 20295 204 20299
tri 204 20295 208 20299 sw
rect 142 20287 208 20295
tri 142 20273 156 20287 ne
rect 156 19152 208 20287
rect 236 19152 288 20330
rect 316 19152 368 20347
rect 396 20351 448 20357
rect 396 20287 448 20299
rect 396 19152 448 20235
rect 476 19152 528 22902
tri 528 22895 535 22902 nw
tri 568 22895 575 22902 se
rect 575 22895 636 22902
tri 556 22883 568 22895 se
rect 568 22889 636 22895
tri 636 22889 649 22902 nw
tri 682 22889 695 22902 se
rect 695 22889 754 22902
rect 568 22883 630 22889
tri 630 22883 636 22889 nw
tri 676 22883 682 22889 se
rect 682 22887 754 22889
tri 754 22887 769 22902 nw
tri 794 22887 809 22902 se
rect 809 22897 868 22902
tri 868 22897 873 22902 nw
tri 908 22897 913 22902 se
rect 913 22897 982 22902
tri 982 22897 987 22902 nw
tri 1022 22897 1027 22902 se
rect 1027 22897 1096 22902
tri 1096 22897 1101 22902 nw
tri 1136 22897 1141 22902 se
rect 1141 22897 1185 22902
rect 809 22887 843 22897
rect 682 22883 739 22887
rect 556 22872 619 22883
tri 619 22872 630 22883 nw
tri 665 22872 676 22883 se
rect 676 22872 739 22883
tri 739 22872 754 22887 nw
tri 779 22872 794 22887 se
rect 794 22872 843 22887
tri 843 22872 868 22897 nw
tri 883 22872 908 22897 se
rect 908 22872 957 22897
tri 957 22872 982 22897 nw
tri 997 22872 1022 22897 se
rect 1022 22872 1071 22897
tri 1071 22872 1096 22897 nw
tri 1111 22872 1136 22897 se
rect 1136 22872 1185 22897
tri 1185 22872 1215 22902 nw
tri 1225 22872 1255 22902 se
rect 1255 22872 1299 22902
tri 1299 22872 1329 22902 nw
rect 556 19152 608 22872
tri 608 22861 619 22872 nw
tri 654 22861 665 22872 se
rect 665 22861 714 22872
tri 636 22843 654 22861 se
rect 654 22847 714 22861
tri 714 22847 739 22872 nw
tri 754 22847 779 22872 se
rect 779 22857 828 22872
tri 828 22857 843 22872 nw
tri 868 22857 883 22872 se
rect 883 22863 948 22872
tri 948 22863 957 22872 nw
tri 988 22863 997 22872 se
rect 997 22863 1062 22872
tri 1062 22863 1071 22872 nw
tri 1102 22863 1111 22872 se
rect 1111 22869 1182 22872
tri 1182 22869 1185 22872 nw
tri 1222 22869 1225 22872 se
rect 1225 22869 1256 22872
rect 1111 22863 1176 22869
tri 1176 22863 1182 22869 nw
tri 1216 22863 1222 22869 se
rect 1222 22863 1256 22869
rect 883 22857 942 22863
tri 942 22857 948 22863 nw
tri 982 22857 988 22863 se
rect 988 22857 1056 22863
tri 1056 22857 1062 22863 nw
tri 1096 22857 1102 22863 se
rect 1102 22857 1142 22863
rect 779 22847 818 22857
tri 818 22847 828 22857 nw
tri 858 22847 868 22857 se
rect 868 22847 908 22857
rect 654 22843 710 22847
tri 710 22843 714 22847 nw
tri 750 22843 754 22847 se
rect 754 22843 796 22847
rect 636 19152 688 22843
tri 688 22821 710 22843 nw
tri 728 22821 750 22843 se
rect 750 22825 796 22843
tri 796 22825 818 22847 nw
tri 836 22825 858 22847 se
rect 858 22825 908 22847
rect 750 22821 780 22825
tri 716 22809 728 22821 se
rect 728 22809 780 22821
tri 780 22809 796 22825 nw
tri 820 22809 836 22825 se
rect 836 22823 908 22825
tri 908 22823 942 22857 nw
tri 948 22823 982 22857 se
rect 982 22823 1022 22857
tri 1022 22823 1056 22857 nw
tri 1062 22823 1096 22857 se
rect 1096 22829 1142 22857
tri 1142 22829 1176 22863 nw
tri 1182 22829 1216 22863 se
rect 1216 22829 1256 22863
tri 1256 22829 1299 22872 nw
rect 1096 22823 1108 22829
rect 836 22809 876 22823
rect 716 19152 768 22809
tri 768 22797 780 22809 nw
tri 808 22797 820 22809 se
rect 820 22797 876 22809
tri 796 22785 808 22797 se
rect 808 22791 876 22797
tri 876 22791 908 22823 nw
tri 916 22791 948 22823 se
rect 948 22791 988 22823
rect 808 22785 870 22791
tri 870 22785 876 22791 nw
tri 914 22789 916 22791 se
rect 916 22789 988 22791
tri 988 22789 1022 22823 nw
tri 1028 22789 1062 22823 se
rect 1062 22795 1108 22823
tri 1108 22795 1142 22829 nw
tri 1148 22795 1182 22829 se
rect 1062 22789 1102 22795
tri 1102 22789 1108 22795 nw
tri 1142 22789 1148 22795 se
rect 1148 22789 1182 22795
tri 910 22785 914 22789 se
rect 914 22785 984 22789
tri 984 22785 988 22789 nw
tri 1024 22785 1028 22789 se
rect 1028 22785 1068 22789
tri 774 18411 796 18433 se
rect 796 18411 848 22785
tri 848 22763 870 22785 nw
tri 888 22763 910 22785 se
rect 910 22783 982 22785
tri 982 22783 984 22785 nw
tri 1022 22783 1024 22785 se
rect 1024 22783 1068 22785
rect 910 22763 962 22783
tri 962 22763 982 22783 nw
tri 1002 22763 1022 22783 se
rect 1022 22763 1068 22783
tri 721 18358 774 18411 se
rect 774 18399 836 18411
tri 836 18399 848 18411 nw
tri 876 22751 888 22763 se
rect 888 22751 950 22763
tri 950 22751 962 22763 nw
tri 990 22751 1002 22763 se
rect 1002 22755 1068 22763
tri 1068 22755 1102 22789 nw
tri 1108 22755 1142 22789 se
rect 1142 22755 1182 22789
tri 1182 22755 1256 22829 nw
rect 1002 22751 1036 22755
rect 774 18392 829 18399
tri 829 18392 836 18399 nw
tri 869 18392 876 18399 se
rect 876 18392 928 22751
tri 928 22729 950 22751 nw
tri 968 22729 990 22751 se
rect 990 22729 1036 22751
rect 774 18358 795 18392
tri 795 18358 829 18392 nw
tri 854 18377 869 18392 se
rect 869 18377 928 18392
tri 835 18358 854 18377 se
rect 854 18358 909 18377
tri 909 18358 928 18377 nw
tri 956 22717 968 22729 se
rect 968 22723 1036 22729
tri 1036 22723 1068 22755 nw
tri 1076 22723 1108 22755 se
rect 1108 22723 1110 22755
rect 968 22717 1030 22723
tri 1030 22717 1036 22723 nw
tri 1070 22717 1076 22723 se
rect 1076 22717 1110 22723
tri 949 18358 956 18365 se
rect 956 18358 1008 22717
tri 1008 22695 1030 22717 nw
tri 1048 22695 1070 22717 se
rect 1070 22695 1110 22717
tri 647 18284 721 18358 se
rect 721 18352 789 18358
tri 789 18352 795 18358 nw
tri 829 18352 835 18358 se
rect 835 18352 903 18358
tri 903 18352 909 18358 nw
tri 943 18352 949 18358 se
rect 949 18352 1008 18358
rect 721 18318 755 18352
tri 755 18318 789 18352 nw
tri 795 18318 829 18352 se
rect 829 18343 894 18352
tri 894 18343 903 18352 nw
tri 934 18343 943 18352 se
rect 943 18343 1008 18352
rect 829 18318 863 18343
tri 721 18284 755 18318 nw
tri 761 18284 795 18318 se
rect 795 18312 863 18318
tri 863 18312 894 18343 nw
tri 903 18312 934 18343 se
rect 934 18331 996 18343
tri 996 18331 1008 18343 nw
tri 1036 22683 1048 22695 se
rect 1048 22683 1110 22695
tri 1110 22683 1182 22755 nw
rect 934 18312 971 18331
rect 795 18284 835 18312
tri 835 18284 863 18312 nw
tri 875 18284 903 18312 se
rect 903 18306 971 18312
tri 971 18306 996 18331 nw
tri 1014 18309 1036 18331 se
rect 1036 18309 1088 22683
tri 1088 22661 1110 22683 nw
rect 8208 22523 8536 24299
tri 8536 24292 8543 24299 nw
tri 8616 24292 8623 24299 se
rect 8623 24292 8935 24299
tri 8592 24268 8616 24292 se
rect 8616 24282 8935 24292
tri 8935 24282 8952 24299 sw
tri 9015 24291 9023 24299 ne
rect 9023 24291 9397 24299
tri 9397 24291 9405 24299 nw
tri 11451 24291 11459 24299 ne
rect 11459 24291 11832 24299
tri 11832 24292 11839 24299 nw
tri 11912 24292 11919 24299 se
rect 11919 24292 12231 24299
tri 9023 24282 9032 24291 ne
rect 9032 24282 9388 24291
tri 9388 24282 9397 24291 nw
tri 9468 24282 9477 24291 se
rect 9477 24282 9759 24291
rect 8616 24268 8952 24282
tri 8952 24268 8966 24282 sw
rect 9032 24268 9374 24282
tri 9374 24268 9388 24282 nw
tri 9454 24268 9468 24282 se
rect 9468 24268 9759 24282
tri 9759 24268 9782 24291 sw
tri 10248 24268 10271 24291 se
rect 10271 24268 10583 24291
tri 10583 24268 10606 24291 sw
tri 11072 24268 11095 24291 se
rect 11095 24268 11379 24291
tri 11379 24268 11402 24291 sw
tri 11459 24268 11482 24291 ne
rect 11482 24268 11832 24291
rect 8592 24216 8628 24268
rect 8680 24216 8692 24268
rect 8744 24216 8756 24268
rect 8808 24216 8820 24268
rect 8872 24216 8884 24268
rect 8936 24261 8966 24268
tri 8966 24261 8973 24268 sw
rect 8936 24216 8973 24261
rect 8592 23890 8973 24216
rect 9032 22523 9360 24268
tri 9360 24254 9374 24268 nw
tri 9440 24254 9454 24268 se
rect 9454 24254 9466 24268
tri 9416 24230 9440 24254 se
rect 9440 24230 9466 24254
rect 9416 24216 9466 24230
rect 9518 24216 9530 24268
rect 9582 24216 9594 24268
rect 9646 24216 9658 24268
rect 9710 24216 9722 24268
rect 9774 24253 9782 24268
tri 9782 24253 9797 24268 sw
rect 9774 24216 9797 24253
rect 9416 23890 9797 24216
tri 10240 24260 10248 24268 se
rect 10248 24260 10276 24268
rect 10240 24216 10276 24260
rect 10328 24216 10340 24268
rect 10392 24216 10404 24268
rect 10456 24216 10468 24268
rect 10520 24216 10532 24268
rect 10584 24253 10606 24268
tri 10606 24253 10621 24268 sw
rect 10584 24216 10621 24253
rect 10240 23890 10621 24216
tri 11064 24260 11072 24268 se
rect 11072 24260 11086 24268
rect 11064 24216 11086 24260
rect 11138 24216 11150 24268
rect 11202 24216 11214 24268
rect 11266 24216 11278 24268
rect 11330 24216 11342 24268
rect 11394 24246 11402 24268
tri 11402 24246 11424 24268 sw
tri 11482 24246 11504 24268 ne
rect 11394 24225 11424 24246
tri 11424 24225 11445 24246 sw
rect 11394 24216 11445 24225
rect 10667 24149 10719 24155
rect 10667 24085 10719 24097
tri 10665 23708 10667 23710 se
rect 10667 23708 10719 24033
tri 10652 23695 10665 23708 se
rect 10665 23695 10719 23708
tri 10618 23661 10652 23695 se
rect 10652 23688 10719 23695
rect 10652 23661 10692 23688
tri 10692 23661 10719 23688 nw
rect 10979 24149 11031 24155
rect 10979 24085 11031 24097
tri 10613 23656 10618 23661 se
rect 10618 23656 10667 23661
tri 10593 23636 10613 23656 se
rect 10613 23636 10667 23656
tri 10667 23636 10692 23661 nw
tri 10585 23628 10593 23636 se
rect 10593 23628 10640 23636
tri 10566 23609 10585 23628 se
rect 10585 23609 10640 23628
tri 10640 23609 10667 23636 nw
tri 10557 23600 10566 23609 se
rect 10566 23600 10631 23609
tri 10631 23600 10640 23609 nw
tri 9997 23578 10019 23600 se
rect 10019 23578 10609 23600
tri 10609 23578 10631 23600 nw
tri 9995 23576 9997 23578 se
rect 9997 23576 10592 23578
tri 9980 23561 9995 23576 se
rect 9995 23561 10592 23576
tri 10592 23561 10609 23578 nw
tri 9967 23548 9980 23561 se
rect 9980 23548 10579 23561
tri 10579 23548 10592 23561 nw
tri 9915 23496 9967 23548 se
rect 9967 23496 10019 23548
tri 9899 23480 9915 23496 se
rect 9915 23480 10019 23496
tri 10019 23480 10087 23548 nw
tri 9887 23468 9899 23480 se
tri 9835 23416 9887 23468 se
rect 9887 23416 9899 23468
tri 9779 23360 9835 23416 se
rect 9835 23360 9899 23416
tri 9899 23360 10019 23480 nw
tri 9777 23358 9779 23360 se
rect 9779 23358 9897 23360
tri 9897 23358 9899 23360 nw
tri 9703 23284 9777 23358 se
rect 9777 23284 9823 23358
tri 9823 23284 9897 23358 nw
tri 10905 23284 10979 23358 se
rect 10979 23336 11031 24033
rect 11064 23890 11445 24216
tri 10979 23284 11031 23336 nw
tri 9667 23248 9703 23284 se
rect 9703 23248 9787 23284
tri 9787 23248 9823 23284 nw
tri 10869 23248 10905 23284 se
rect 10905 23248 10943 23284
tri 10943 23248 10979 23284 nw
tri 9660 23241 9667 23248 se
rect 9667 23241 9780 23248
tri 9780 23241 9787 23248 nw
tri 10205 23241 10212 23248 se
rect 10212 23241 10891 23248
rect 9660 22902 9776 23241
tri 9776 23237 9780 23241 nw
tri 10201 23237 10205 23241 se
rect 10205 23237 10891 23241
tri 10092 23128 10201 23237 se
rect 10201 23196 10891 23237
tri 10891 23196 10943 23248 nw
rect 10201 23128 10212 23196
tri 10212 23128 10280 23196 nw
tri 10076 23112 10092 23128 se
rect 10092 23112 10196 23128
tri 10196 23112 10212 23128 nw
rect 10076 22902 10192 23112
tri 10192 23108 10196 23112 nw
rect 11504 22523 11832 24268
tri 11888 24268 11912 24292 se
rect 11912 24282 12231 24292
tri 12231 24282 12248 24299 sw
tri 12311 24282 12328 24299 ne
rect 11912 24268 12248 24282
tri 12248 24268 12262 24282 sw
rect 11888 24216 11924 24268
rect 11976 24216 11988 24268
rect 12040 24216 12052 24268
rect 12104 24216 12116 24268
rect 12168 24216 12180 24268
rect 12232 24261 12262 24268
tri 12262 24261 12269 24268 sw
rect 12232 24216 12269 24261
rect 11888 23890 12269 24216
rect 12328 22523 12656 24299
tri 12656 24292 12663 24299 nw
tri 12736 24292 12743 24299 se
rect 12743 24292 13055 24299
tri 12712 24268 12736 24292 se
rect 12736 24282 13055 24292
tri 13055 24282 13072 24299 sw
tri 13135 24282 13152 24299 ne
rect 12736 24268 13072 24282
tri 13072 24268 13086 24282 sw
rect 12712 24216 12748 24268
rect 12800 24216 12812 24268
rect 12864 24216 12876 24268
rect 12928 24216 12940 24268
rect 12992 24216 13004 24268
rect 13056 24261 13086 24268
tri 13086 24261 13093 24268 sw
rect 13056 24216 13093 24261
rect 12712 23890 13093 24216
rect 13152 22523 13480 24299
tri 13480 24292 13487 24299 nw
tri 13560 24292 13567 24299 se
rect 13567 24292 13879 24299
tri 13536 24268 13560 24292 se
rect 13560 24282 13879 24292
tri 13879 24282 13896 24299 sw
tri 13959 24282 13976 24299 ne
rect 13560 24268 13896 24282
tri 13896 24268 13910 24282 sw
rect 13536 24216 13572 24268
rect 13624 24216 13636 24268
rect 13688 24216 13700 24268
rect 13752 24216 13764 24268
rect 13816 24216 13828 24268
rect 13880 24261 13910 24268
tri 13910 24261 13917 24268 sw
rect 13880 24216 13917 24261
rect 13536 23890 13917 24216
rect 13976 22523 14304 24299
tri 14304 24292 14311 24299 nw
tri 14384 24292 14391 24299 se
rect 14391 24292 14703 24299
tri 14360 24268 14384 24292 se
rect 14384 24282 14703 24292
tri 14703 24282 14720 24299 sw
tri 14783 24282 14800 24299 ne
rect 14384 24268 14720 24282
tri 14720 24268 14734 24282 sw
rect 14360 24216 14396 24268
rect 14448 24216 14460 24268
rect 14512 24216 14524 24268
rect 14576 24216 14588 24268
rect 14640 24216 14652 24268
rect 14704 24261 14734 24268
tri 14734 24261 14741 24268 sw
rect 14704 24216 14741 24261
rect 14360 23890 14741 24216
rect 14800 22523 15128 24299
tri 15128 24292 15135 24299 nw
tri 15208 24292 15215 24299 se
rect 15215 24292 15527 24299
tri 15184 24268 15208 24292 se
rect 15208 24282 15527 24292
tri 15527 24282 15544 24299 sw
tri 15607 24282 15624 24299 ne
rect 15208 24268 15544 24282
tri 15544 24268 15558 24282 sw
rect 15184 24216 15220 24268
rect 15272 24216 15284 24268
rect 15336 24216 15348 24268
rect 15400 24216 15412 24268
rect 15464 24216 15476 24268
rect 15528 24261 15558 24268
tri 15558 24261 15565 24268 sw
rect 15528 24216 15565 24261
rect 15184 23890 15565 24216
rect 15167 23733 15173 23785
rect 15225 23733 15238 23785
rect 15290 23733 15296 23785
rect 15336 23733 15342 23785
rect 15394 23733 15407 23785
rect 15459 23733 15465 23785
tri 15176 23727 15182 23733 ne
rect 15182 23727 15296 23733
tri 15182 23714 15195 23727 ne
rect 15195 23714 15296 23727
tri 15195 23699 15210 23714 ne
rect 15210 23661 15296 23714
tri 15296 23661 15330 23695 sw
rect 15210 23609 15216 23661
rect 15268 23609 15285 23661
rect 15337 23609 15353 23661
rect 15405 23609 15411 23661
rect 15624 22523 15952 24299
tri 15952 24292 15959 24299 nw
tri 16032 24292 16039 24299 se
rect 16039 24292 16351 24299
tri 16008 24268 16032 24292 se
rect 16032 24282 16351 24292
tri 16351 24282 16368 24299 sw
tri 16431 24282 16448 24299 ne
rect 16032 24268 16368 24282
tri 16368 24268 16382 24282 sw
rect 16008 24216 16044 24268
rect 16096 24216 16108 24268
rect 16160 24216 16172 24268
rect 16224 24216 16236 24268
rect 16288 24216 16300 24268
rect 16352 24261 16382 24268
tri 16382 24261 16389 24268 sw
rect 16352 24216 16389 24261
rect 16008 23890 16389 24216
rect 16448 22523 16776 24299
tri 16776 24292 16783 24299 nw
tri 16856 24292 16863 24299 se
rect 16863 24292 17175 24299
tri 16832 24268 16856 24292 se
rect 16856 24291 17175 24292
tri 17175 24291 17183 24299 sw
tri 17255 24291 17263 24299 ne
rect 16856 24268 17183 24291
tri 17183 24268 17206 24291 sw
rect 16832 24216 16868 24268
rect 16920 24216 16932 24268
rect 16984 24216 16996 24268
rect 17048 24216 17060 24268
rect 17112 24216 17124 24268
rect 17176 24261 17206 24268
tri 17206 24261 17213 24268 sw
rect 17176 24216 17213 24261
rect 16832 23890 17213 24216
rect 16828 23695 17130 23701
rect 16880 23664 17130 23695
tri 17130 23664 17167 23701 sw
rect 16880 23651 17167 23664
rect 16880 23649 16912 23651
tri 16912 23649 16914 23651 nw
tri 17090 23649 17092 23651 ne
rect 17092 23649 17167 23651
rect 16828 23630 16880 23643
tri 16880 23617 16912 23649 nw
tri 17092 23624 17117 23649 ne
rect 16828 23572 16880 23578
rect 16956 23561 16962 23613
rect 17014 23561 17026 23613
rect 17078 23561 17084 23613
rect 16956 22872 17084 23561
rect 17117 22994 17167 23649
tri 17167 22994 17233 23060 sw
rect 17263 22523 17573 24299
rect 17629 24767 17652 25982
rect 18344 24767 18369 26035
rect 17629 24754 18369 24767
rect 17629 24702 17652 24754
rect 17704 24702 17716 24754
rect 17768 24702 17780 24754
rect 17832 24702 17844 24754
rect 17896 24702 17908 24754
rect 17960 24702 17972 24754
rect 18024 24702 18036 24754
rect 18088 24702 18100 24754
rect 18152 24702 18164 24754
rect 18216 24702 18228 24754
rect 18280 24702 18292 24754
rect 18344 24702 18369 24754
rect 17629 24689 18369 24702
rect 17629 24637 17652 24689
rect 17704 24637 17716 24689
rect 17768 24637 17780 24689
rect 17832 24637 17844 24689
rect 17896 24637 17908 24689
rect 17960 24637 17972 24689
rect 18024 24637 18036 24689
rect 18088 24637 18100 24689
rect 18152 24637 18164 24689
rect 18216 24637 18228 24689
rect 18280 24637 18292 24689
rect 18344 24637 18369 24689
rect 17629 24624 18369 24637
rect 17629 24572 17652 24624
rect 17704 24572 17716 24624
rect 17768 24572 17780 24624
rect 17832 24572 17844 24624
rect 17896 24572 17908 24624
rect 17960 24572 17972 24624
rect 18024 24572 18036 24624
rect 18088 24572 18100 24624
rect 18152 24572 18164 24624
rect 18216 24572 18228 24624
rect 18280 24572 18292 24624
rect 18344 24572 18369 24624
rect 17629 24559 18369 24572
rect 17629 24507 17652 24559
rect 17704 24507 17716 24559
rect 17768 24507 17780 24559
rect 17832 24507 17844 24559
rect 17896 24507 17908 24559
rect 17960 24507 17972 24559
rect 18024 24507 18036 24559
rect 18088 24507 18100 24559
rect 18152 24507 18164 24559
rect 18216 24507 18228 24559
rect 18280 24507 18292 24559
rect 18344 24507 18369 24559
rect 17629 24494 18369 24507
rect 17629 24442 17652 24494
rect 17704 24442 17716 24494
rect 17768 24442 17780 24494
rect 17832 24442 17844 24494
rect 17896 24442 17908 24494
rect 17960 24442 17972 24494
rect 18024 24442 18036 24494
rect 18088 24442 18100 24494
rect 18152 24442 18164 24494
rect 18216 24442 18228 24494
rect 18280 24442 18292 24494
rect 18344 24442 18369 24494
rect 17629 24429 18369 24442
rect 17629 24377 17652 24429
rect 17704 24377 17716 24429
rect 17768 24377 17780 24429
rect 17832 24377 17844 24429
rect 17896 24377 17908 24429
rect 17960 24377 17972 24429
rect 18024 24377 18036 24429
rect 18088 24377 18100 24429
rect 18152 24377 18164 24429
rect 18216 24377 18228 24429
rect 18280 24377 18292 24429
rect 18344 24377 18369 24429
rect 17629 24364 18369 24377
rect 17629 24312 17652 24364
rect 17704 24312 17716 24364
rect 17768 24312 17780 24364
rect 17832 24312 17844 24364
rect 17896 24312 17908 24364
rect 17960 24312 17972 24364
rect 18024 24312 18036 24364
rect 18088 24312 18100 24364
rect 18152 24312 18164 24364
rect 18216 24312 18228 24364
rect 18280 24312 18292 24364
rect 18344 24312 18369 24364
rect 17629 24299 18369 24312
rect 17629 24247 17652 24299
rect 17704 24247 17716 24299
rect 17768 24247 17780 24299
rect 17832 24247 17844 24299
rect 17896 24247 17908 24299
rect 17960 24247 17972 24299
rect 18024 24247 18036 24299
rect 18088 24247 18100 24299
rect 18152 24247 18164 24299
rect 18216 24247 18228 24299
rect 18280 24247 18292 24299
rect 18344 24247 18369 24299
rect 17629 24234 18369 24247
rect 17629 24182 17652 24234
rect 17704 24182 17716 24234
rect 17768 24182 17780 24234
rect 17832 24182 17844 24234
rect 17896 24182 17908 24234
rect 17960 24182 17972 24234
rect 18024 24182 18036 24234
rect 18088 24182 18100 24234
rect 18152 24182 18164 24234
rect 18216 24182 18228 24234
rect 18280 24182 18292 24234
rect 18344 24182 18369 24234
rect 17629 24169 18369 24182
rect 17629 24117 17652 24169
rect 17704 24117 17716 24169
rect 17768 24117 17780 24169
rect 17832 24117 17844 24169
rect 17896 24117 17908 24169
rect 17960 24117 17972 24169
rect 18024 24117 18036 24169
rect 18088 24117 18100 24169
rect 18152 24117 18164 24169
rect 18216 24117 18228 24169
rect 18280 24117 18292 24169
rect 18344 24117 18369 24169
rect 17629 24104 18369 24117
rect 17629 24052 17652 24104
rect 17704 24052 17716 24104
rect 17768 24052 17780 24104
rect 17832 24052 17844 24104
rect 17896 24052 17908 24104
rect 17960 24052 17972 24104
rect 18024 24052 18036 24104
rect 18088 24052 18100 24104
rect 18152 24052 18164 24104
rect 18216 24052 18228 24104
rect 18280 24052 18292 24104
rect 18344 24052 18369 24104
rect 17629 24039 18369 24052
rect 17629 23987 17652 24039
rect 17704 23987 17716 24039
rect 17768 23987 17780 24039
rect 17832 23987 17844 24039
rect 17896 23987 17908 24039
rect 17960 23987 17972 24039
rect 18024 23987 18036 24039
rect 18088 23987 18100 24039
rect 18152 23987 18164 24039
rect 18216 23987 18228 24039
rect 18280 23987 18292 24039
rect 18344 23987 18369 24039
rect 17629 23974 18369 23987
rect 17629 23922 17652 23974
rect 17704 23922 17716 23974
rect 17768 23922 17780 23974
rect 17832 23922 17844 23974
rect 17896 23922 17908 23974
rect 17960 23922 17972 23974
rect 18024 23922 18036 23974
rect 18088 23922 18100 23974
rect 18152 23922 18164 23974
rect 18216 23922 18228 23974
rect 18280 23922 18292 23974
rect 18344 23922 18369 23974
rect 17629 23909 18369 23922
rect 17629 23857 17652 23909
rect 17704 23857 17716 23909
rect 17768 23857 17780 23909
rect 17832 23857 17844 23909
rect 17896 23857 17908 23909
rect 17960 23857 17972 23909
rect 18024 23857 18036 23909
rect 18088 23857 18100 23909
rect 18152 23857 18164 23909
rect 18216 23857 18228 23909
rect 18280 23857 18292 23909
rect 18344 23857 18369 23909
rect 17629 23844 18369 23857
rect 17629 23792 17652 23844
rect 17704 23792 17716 23844
rect 17768 23792 17780 23844
rect 17832 23792 17844 23844
rect 17896 23792 17908 23844
rect 17960 23792 17972 23844
rect 18024 23792 18036 23844
rect 18088 23792 18100 23844
rect 18152 23792 18164 23844
rect 18216 23792 18228 23844
rect 18280 23792 18292 23844
rect 18344 23792 18369 23844
rect 17629 23779 18369 23792
rect 17629 23727 17652 23779
rect 17704 23727 17716 23779
rect 17768 23727 17780 23779
rect 17832 23727 17844 23779
rect 17896 23727 17908 23779
rect 17960 23727 17972 23779
rect 18024 23727 18036 23779
rect 18088 23727 18100 23779
rect 18152 23727 18164 23779
rect 18216 23727 18228 23779
rect 18280 23727 18292 23779
rect 18344 23727 18369 23779
rect 17629 23714 18369 23727
rect 17629 23662 17652 23714
rect 17704 23662 17716 23714
rect 17768 23662 17780 23714
rect 17832 23662 17844 23714
rect 17896 23662 17908 23714
rect 17960 23662 17972 23714
rect 18024 23662 18036 23714
rect 18088 23662 18100 23714
rect 18152 23662 18164 23714
rect 18216 23662 18228 23714
rect 18280 23662 18292 23714
rect 18344 23662 18369 23714
rect 17629 23649 18369 23662
rect 17629 23597 17652 23649
rect 17704 23597 17716 23649
rect 17768 23597 17780 23649
rect 17832 23597 17844 23649
rect 17896 23597 17908 23649
rect 17960 23597 17972 23649
rect 18024 23597 18036 23649
rect 18088 23597 18100 23649
rect 18152 23597 18164 23649
rect 18216 23597 18228 23649
rect 18280 23597 18292 23649
rect 18344 23597 18369 23649
rect 17629 22523 18369 23597
tri 1011 18306 1014 18309 se
rect 1014 18306 1063 18309
rect 903 18284 949 18306
tri 949 18284 971 18306 nw
tri 989 18284 1011 18306 se
rect 1011 18284 1063 18306
tri 1063 18284 1088 18309 nw
tri 573 18210 647 18284 se
rect 647 18278 715 18284
tri 715 18278 721 18284 nw
tri 755 18278 761 18284 se
rect 761 18278 829 18284
tri 829 18278 835 18284 nw
tri 869 18278 875 18284 se
rect 875 18278 943 18284
tri 943 18278 949 18284 nw
tri 983 18278 989 18284 se
rect 989 18278 1057 18284
tri 1057 18278 1063 18284 nw
rect 647 18244 681 18278
tri 681 18244 715 18278 nw
tri 721 18244 755 18278 se
rect 755 18272 823 18278
tri 823 18272 829 18278 nw
tri 863 18272 869 18278 se
rect 869 18272 937 18278
tri 937 18272 943 18278 nw
tri 977 18272 983 18278 se
rect 983 18272 1051 18278
tri 1051 18272 1057 18278 nw
rect 755 18244 789 18272
tri 647 18210 681 18244 nw
tri 687 18210 721 18244 se
rect 721 18238 789 18244
tri 789 18238 823 18272 nw
tri 829 18238 863 18272 se
rect 863 18266 931 18272
tri 931 18266 937 18272 nw
tri 971 18266 977 18272 se
rect 977 18266 1045 18272
tri 1045 18266 1051 18272 nw
rect 863 18238 897 18266
rect 721 18210 761 18238
tri 761 18210 789 18238 nw
tri 801 18210 829 18238 se
rect 829 18232 897 18238
tri 897 18232 931 18266 nw
tri 937 18232 971 18266 se
rect 971 18232 989 18266
rect 829 18210 875 18232
tri 875 18210 897 18232 nw
tri 915 18210 937 18232 se
rect 937 18210 989 18232
tri 989 18210 1045 18266 nw
tri 499 18136 573 18210 se
rect 573 18204 641 18210
tri 641 18204 647 18210 nw
tri 681 18204 687 18210 se
rect 687 18204 755 18210
tri 755 18204 761 18210 nw
tri 795 18204 801 18210 se
rect 801 18204 869 18210
tri 869 18204 875 18210 nw
tri 909 18204 915 18210 se
rect 915 18204 983 18210
tri 983 18204 989 18210 nw
rect 573 18170 607 18204
tri 607 18170 641 18204 nw
tri 647 18170 681 18204 se
rect 681 18198 749 18204
tri 749 18198 755 18204 nw
tri 789 18198 795 18204 se
rect 795 18198 863 18204
tri 863 18198 869 18204 nw
tri 903 18198 909 18204 se
rect 909 18198 977 18204
tri 977 18198 983 18204 nw
rect 681 18170 715 18198
tri 573 18136 607 18170 nw
tri 613 18136 647 18170 se
rect 647 18164 715 18170
tri 715 18164 749 18198 nw
tri 755 18164 789 18198 se
rect 789 18192 857 18198
tri 857 18192 863 18198 nw
tri 897 18192 903 18198 se
rect 903 18192 971 18198
tri 971 18192 977 18198 nw
rect 789 18164 823 18192
rect 647 18136 687 18164
tri 687 18136 715 18164 nw
tri 727 18136 755 18164 se
rect 755 18158 823 18164
tri 823 18158 857 18192 nw
tri 863 18158 897 18192 se
rect 897 18158 915 18192
rect 755 18136 801 18158
tri 801 18136 823 18158 nw
tri 841 18136 863 18158 se
rect 863 18136 915 18158
tri 915 18136 971 18192 nw
tri 425 18062 499 18136 se
rect 499 18130 567 18136
tri 567 18130 573 18136 nw
tri 607 18130 613 18136 se
rect 613 18130 681 18136
tri 681 18130 687 18136 nw
tri 721 18130 727 18136 se
rect 727 18130 795 18136
tri 795 18130 801 18136 nw
tri 835 18130 841 18136 se
rect 841 18130 909 18136
tri 909 18130 915 18136 nw
rect 499 18096 533 18130
tri 533 18096 567 18130 nw
tri 573 18096 607 18130 se
rect 607 18124 675 18130
tri 675 18124 681 18130 nw
tri 715 18124 721 18130 se
rect 721 18124 789 18130
tri 789 18124 795 18130 nw
tri 829 18124 835 18130 se
rect 835 18124 903 18130
tri 903 18124 909 18130 nw
rect 607 18096 641 18124
tri 499 18062 533 18096 nw
tri 539 18062 573 18096 se
rect 573 18090 641 18096
tri 641 18090 675 18124 nw
tri 681 18090 715 18124 se
rect 715 18118 783 18124
tri 783 18118 789 18124 nw
tri 823 18118 829 18124 se
rect 829 18118 897 18124
tri 897 18118 903 18124 nw
rect 715 18090 749 18118
rect 573 18062 613 18090
tri 613 18062 641 18090 nw
tri 653 18062 681 18090 se
rect 681 18084 749 18090
tri 749 18084 783 18118 nw
tri 789 18084 823 18118 se
rect 823 18084 841 18118
rect 681 18062 727 18084
tri 727 18062 749 18084 nw
tri 767 18062 789 18084 se
rect 789 18062 841 18084
tri 841 18062 897 18118 nw
tri 351 17988 425 18062 se
rect 425 18056 493 18062
tri 493 18056 499 18062 nw
tri 533 18056 539 18062 se
rect 539 18056 607 18062
tri 607 18056 613 18062 nw
tri 647 18056 653 18062 se
rect 653 18056 721 18062
tri 721 18056 727 18062 nw
tri 761 18056 767 18062 se
rect 767 18056 835 18062
tri 835 18056 841 18062 nw
rect 425 18022 459 18056
tri 459 18022 493 18056 nw
tri 499 18022 533 18056 se
rect 533 18050 601 18056
tri 601 18050 607 18056 nw
tri 641 18050 647 18056 se
rect 647 18050 715 18056
tri 715 18050 721 18056 nw
tri 755 18050 761 18056 se
rect 761 18050 829 18056
tri 829 18050 835 18056 nw
rect 533 18022 567 18050
tri 425 17988 459 18022 nw
tri 465 17988 499 18022 se
rect 499 18016 567 18022
tri 567 18016 601 18050 nw
tri 607 18016 641 18050 se
rect 641 18044 709 18050
tri 709 18044 715 18050 nw
tri 749 18044 755 18050 se
rect 755 18044 823 18050
tri 823 18044 829 18050 nw
rect 641 18016 675 18044
rect 499 17988 539 18016
tri 539 17988 567 18016 nw
tri 579 17988 607 18016 se
rect 607 18010 675 18016
tri 675 18010 709 18044 nw
tri 715 18010 749 18044 se
rect 749 18010 767 18044
rect 607 17988 653 18010
tri 653 17988 675 18010 nw
tri 693 17988 715 18010 se
rect 715 17988 767 18010
tri 767 17988 823 18044 nw
tri 329 17966 351 17988 se
rect 351 17982 419 17988
tri 419 17982 425 17988 nw
tri 459 17982 465 17988 se
rect 465 17982 533 17988
tri 533 17982 539 17988 nw
tri 573 17982 579 17988 se
rect 579 17982 647 17988
tri 647 17982 653 17988 nw
tri 687 17982 693 17988 se
rect 693 17982 761 17988
tri 761 17982 767 17988 nw
rect 351 17966 403 17982
tri 403 17966 419 17982 nw
tri 443 17966 459 17982 se
rect 459 17976 527 17982
tri 527 17976 533 17982 nw
tri 567 17976 573 17982 se
rect 573 17976 641 17982
tri 641 17976 647 17982 nw
tri 681 17976 687 17982 se
rect 687 17976 755 17982
tri 755 17976 761 17982 nw
rect 459 17966 517 17976
tri 517 17966 527 17976 nw
tri 557 17966 567 17976 se
rect 567 17970 635 17976
tri 635 17970 641 17976 nw
tri 675 17970 681 17976 se
rect 681 17970 749 17976
tri 749 17970 755 17976 nw
rect 567 17966 631 17970
tri 631 17966 635 17970 nw
tri 671 17966 675 17970 se
rect 675 17966 745 17970
tri 745 17966 749 17970 nw
tri -2873 17914 -2821 17966 se
rect -2821 17948 385 17966
tri 385 17948 403 17966 nw
tri 425 17948 443 17966 se
rect 443 17948 493 17966
rect -2821 17914 351 17948
tri 351 17914 385 17948 nw
tri 391 17914 425 17948 se
rect 425 17942 493 17948
tri 493 17942 517 17966 nw
tri 533 17942 557 17966 se
rect 557 17942 601 17966
rect 425 17914 465 17942
tri 465 17914 493 17942 nw
tri 505 17914 533 17942 se
rect 533 17936 601 17942
tri 601 17936 631 17966 nw
tri 641 17936 671 17966 se
rect 671 17936 693 17966
rect 533 17914 579 17936
tri 579 17914 601 17936 nw
tri 619 17914 641 17936 se
rect 641 17914 693 17936
tri 693 17914 745 17966 nw
tri -2895 17892 -2873 17914 se
rect -2873 17892 -2821 17914
tri -2821 17892 -2799 17914 nw
tri 385 17908 391 17914 se
rect 391 17908 459 17914
tri 459 17908 465 17914 nw
tri 499 17908 505 17914 se
rect 505 17908 573 17914
tri 573 17908 579 17914 nw
tri 613 17908 619 17914 se
rect 619 17908 687 17914
tri 687 17908 693 17914 nw
tri 369 17892 385 17908 se
rect 385 17902 453 17908
tri 453 17902 459 17908 nw
tri 493 17902 499 17908 se
rect 499 17902 567 17908
tri 567 17902 573 17908 nw
tri 607 17902 613 17908 se
rect 613 17902 681 17908
tri 681 17902 687 17908 nw
rect 385 17892 443 17902
tri 443 17892 453 17902 nw
tri 483 17892 493 17902 se
rect 493 17896 561 17902
tri 561 17896 567 17902 nw
tri 601 17896 607 17902 se
rect 607 17896 675 17902
tri 675 17896 681 17902 nw
rect 493 17892 557 17896
tri 557 17892 561 17896 nw
tri 597 17892 601 17896 se
rect 601 17892 671 17896
tri 671 17892 675 17896 nw
tri -2901 17886 -2895 17892 se
rect -2895 17886 -2827 17892
tri -2827 17886 -2821 17892 nw
tri 363 17886 369 17892 se
rect 369 17886 437 17892
tri 437 17886 443 17892 nw
tri 477 17886 483 17892 se
rect 483 17886 551 17892
tri 551 17886 557 17892 nw
tri 591 17886 597 17892 se
rect 597 17886 665 17892
tri 665 17886 671 17892 nw
tri -2969 17818 -2901 17886 se
rect -2901 17852 -2861 17886
tri -2861 17852 -2827 17886 nw
tri -2821 17852 -2787 17886 se
rect -2787 17868 419 17886
tri 419 17868 437 17886 nw
tri 459 17868 477 17886 se
rect 477 17868 527 17886
rect -2787 17852 385 17868
rect -2901 17818 -2895 17852
tri -2895 17818 -2861 17852 nw
tri -2855 17818 -2821 17852 se
rect -2821 17834 385 17852
tri 385 17834 419 17868 nw
tri 425 17834 459 17868 se
rect 459 17862 527 17868
tri 527 17862 551 17886 nw
tri 567 17862 591 17886 se
rect 591 17862 613 17886
rect 459 17834 499 17862
tri 499 17834 527 17862 nw
tri 539 17834 567 17862 se
rect 567 17834 613 17862
tri 613 17834 665 17886 nw
rect -2821 17818 -2787 17834
tri -2975 17812 -2969 17818 se
rect -2969 17812 -2901 17818
tri -2901 17812 -2895 17818 nw
tri -2861 17812 -2855 17818 se
rect -2855 17812 -2787 17818
tri -2787 17812 -2765 17834 nw
tri 419 17828 425 17834 se
rect 425 17828 493 17834
tri 493 17828 499 17834 nw
tri 533 17828 539 17834 se
rect 539 17828 607 17834
tri 607 17828 613 17834 nw
tri 403 17812 419 17828 se
rect 419 17822 487 17828
tri 487 17822 493 17828 nw
tri 527 17822 533 17828 se
rect 533 17822 601 17828
tri 601 17822 607 17828 nw
rect 419 17812 477 17822
tri 477 17812 487 17822 nw
tri 517 17812 527 17822 se
rect 527 17812 591 17822
tri 591 17812 601 17822 nw
tri -3043 17744 -2975 17812 se
rect -2975 17778 -2935 17812
tri -2935 17778 -2901 17812 nw
tri -2895 17778 -2861 17812 se
rect -2861 17806 -2793 17812
tri -2793 17806 -2787 17812 nw
tri 397 17806 403 17812 se
rect 403 17806 471 17812
tri 471 17806 477 17812 nw
tri 511 17806 517 17812 se
rect 517 17806 585 17812
tri 585 17806 591 17812 nw
rect -2861 17778 -2827 17806
rect -2975 17744 -2969 17778
tri -2969 17744 -2935 17778 nw
tri -2929 17744 -2895 17778 se
rect -2895 17772 -2827 17778
tri -2827 17772 -2793 17806 nw
tri -2787 17772 -2753 17806 se
rect -2753 17788 453 17806
tri 453 17788 471 17806 nw
tri 493 17788 511 17806 se
rect 511 17788 533 17806
rect -2753 17772 419 17788
rect -2895 17744 -2861 17772
tri -3049 17738 -3043 17744 se
rect -3043 17738 -2975 17744
tri -2975 17738 -2969 17744 nw
tri -2935 17738 -2929 17744 se
rect -2929 17738 -2861 17744
tri -2861 17738 -2827 17772 nw
tri -2821 17738 -2787 17772 se
rect -2787 17754 419 17772
tri 419 17754 453 17788 nw
tri 459 17754 493 17788 se
rect 493 17754 533 17788
tri 533 17754 585 17806 nw
rect -2787 17738 -2753 17754
tri -3088 17699 -3049 17738 se
rect -3049 17704 -3009 17738
tri -3009 17704 -2975 17738 nw
tri -2969 17704 -2935 17738 se
rect -2935 17732 -2867 17738
tri -2867 17732 -2861 17738 nw
tri -2827 17732 -2821 17738 se
rect -2821 17732 -2753 17738
tri -2753 17732 -2731 17754 nw
tri 453 17748 459 17754 se
rect 459 17748 527 17754
tri 527 17748 533 17754 nw
tri 437 17732 453 17748 se
rect 453 17732 511 17748
tri 511 17732 527 17748 nw
rect -2935 17704 -2901 17732
rect -3049 17699 -3014 17704
tri -3014 17699 -3009 17704 nw
tri -2974 17699 -2969 17704 se
rect -2969 17699 -2901 17704
tri -3356 5051 -3328 5079 se
rect -3088 4641 -3036 17699
tri -3036 17677 -3014 17699 nw
tri -2996 17677 -2974 17699 se
rect -2974 17698 -2901 17699
tri -2901 17698 -2867 17732 nw
tri -2861 17698 -2827 17732 se
rect -2827 17726 -2759 17732
tri -2759 17726 -2753 17732 nw
tri 431 17726 437 17732 se
rect 437 17726 505 17732
tri 505 17726 511 17732 nw
rect -2827 17698 -2793 17726
rect -2974 17677 -2934 17698
rect -3088 4577 -3036 4589
rect -3088 4218 -3036 4525
tri -3008 17665 -2996 17677 se
rect -2996 17665 -2934 17677
tri -2934 17665 -2901 17698 nw
tri -2894 17665 -2861 17698 se
rect -2861 17692 -2793 17698
tri -2793 17692 -2759 17726 nw
tri -2753 17692 -2719 17726 se
rect -2719 17692 453 17726
rect -2861 17665 -2827 17692
rect -3008 4472 -2956 17665
tri -2956 17643 -2934 17665 nw
tri -2901 17658 -2894 17665 se
rect -2894 17658 -2827 17665
tri -2827 17658 -2793 17692 nw
tri -2787 17658 -2753 17692 se
rect -2753 17674 453 17692
tri 453 17674 505 17726 nw
rect -2753 17658 -2719 17674
tri -2916 17643 -2901 17658 se
rect -2901 17652 -2833 17658
tri -2833 17652 -2827 17658 nw
tri -2793 17652 -2787 17658 se
rect -2787 17652 -2719 17658
tri -2719 17652 -2697 17674 nw
rect -2901 17643 -2848 17652
tri -2928 17631 -2916 17643 se
rect -2916 17637 -2848 17643
tri -2848 17637 -2833 17652 nw
tri -2808 17637 -2793 17652 se
rect -2793 17637 -2774 17652
rect -2916 17631 -2854 17637
tri -2854 17631 -2848 17637 nw
tri -2814 17631 -2808 17637 se
rect -2808 17631 -2774 17637
rect -2928 4710 -2876 17631
tri -2876 17609 -2854 17631 nw
tri -2836 17609 -2814 17631 se
rect -2814 17609 -2774 17631
tri -2848 17597 -2836 17609 se
rect -2836 17597 -2774 17609
tri -2774 17597 -2719 17652 nw
rect -2848 4892 -2796 17597
tri -2796 17575 -2774 17597 nw
rect 921 4955 927 5007
rect 979 4955 991 5007
rect 1043 4955 1049 5007
tri 931 4930 956 4955 ne
tri -2796 4892 -2792 4896 sw
rect -2848 4886 -2792 4892
tri -2792 4886 -2786 4892 sw
rect -2848 4854 -2786 4886
tri -2786 4854 -2754 4886 sw
rect -2848 4802 -2842 4854
rect -2790 4802 -2778 4854
rect -2726 4802 -2720 4854
rect 956 4762 1008 4955
tri 1008 4930 1033 4955 nw
rect 1036 4886 1088 4892
rect 1036 4822 1088 4834
rect 1036 4764 1088 4770
tri -2876 4710 -2849 4737 sw
rect -2928 4698 -2849 4710
tri -2849 4698 -2837 4710 sw
rect 956 4698 1008 4710
rect -2928 4695 -2837 4698
tri -2837 4695 -2834 4698 sw
rect -2928 4643 -2922 4695
rect -2870 4643 -2858 4695
rect -2806 4643 -2800 4695
rect 956 4640 1008 4646
rect 796 4588 848 4594
rect 796 4524 848 4536
tri -2956 4472 -2953 4475 sw
rect -3008 4466 -2953 4472
tri -2953 4466 -2947 4472 sw
rect -3008 4464 -2947 4466
tri -2947 4464 -2945 4466 sw
rect -3008 4433 -2945 4464
tri -2945 4433 -2914 4464 sw
rect -3008 4381 -3002 4433
rect -2950 4381 -2938 4433
rect -2886 4381 -2880 4433
rect 796 4340 848 4472
rect 876 4464 928 4470
rect 876 4400 928 4412
rect 876 4342 928 4348
rect 796 4276 848 4288
rect 796 4218 848 4224
<< metal3 >>
rect 7768 23899 8154 24135
rect 8592 23904 8980 24140
rect 9416 23904 9804 24140
rect 10240 23904 10628 24140
rect 11064 23904 11452 24140
rect 11888 23904 12276 24140
rect 12712 23904 13100 24140
rect 13536 23904 13924 24140
rect 14360 23904 14748 24140
rect 15184 23904 15572 24140
rect 16008 23904 16396 24140
rect 16832 23904 17220 24140
tri 13922 23902 13924 23904 nw
tri -244 22966 -170 23040 se
rect -170 22966 72 23040
tri 72 22966 146 23040 sw
rect -244 17883 146 22966
<< metal4 >>
tri 4177 23939 4472 24234 se
rect 4472 23939 17218 24376
rect 4177 23909 17218 23939
rect 4177 23404 15403 23909
tri 15403 23622 15690 23909 nw
tri 12098 22414 13088 23404 ne
rect 13088 22516 15403 23404
rect 13088 22414 15301 22516
tri 15301 22414 15403 22516 nw
rect 13088 20701 13588 22414
tri 13588 20701 15301 22414 nw
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 11350 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 11726 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 12138 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 12550 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 12962 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 13374 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 13786 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 14198 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 14574 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 11726 0 1 23588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 11350 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 12138 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 12550 0 1 23588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 12962 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform -1 0 13374 0 1 23588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform -1 0 13786 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform -1 0 14198 0 1 23588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform -1 0 14574 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 0 -1 2916 1 0 25369
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 4410 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 4822 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 5234 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 5646 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 6058 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 6470 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 6882 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 7294 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 1 0 7706 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 1 0 14656 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1707688321
transform 1 0 8118 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1707688321
transform 1 0 8530 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1707688321
transform 1 0 8942 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1707688321
transform 1 0 9354 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1707688321
transform 1 0 9766 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1707688321
transform 1 0 10178 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1707688321
transform 1 0 10590 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1707688321
transform 1 0 4410 0 1 23665
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1707688321
transform 1 0 11414 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1707688321
transform 1 0 13062 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1707688321
transform 1 0 13886 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1707688321
transform 1 0 13474 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1707688321
transform 1 0 11826 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1707688321
transform 1 0 12238 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1707688321
transform 1 0 14298 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1707688321
transform 1 0 12650 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1707688321
transform 1 0 11002 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1707688321
transform 1 0 11002 0 1 23588
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_47
timestamp 1707688321
transform 1 0 15536 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_48
timestamp 1707688321
transform 1 0 15124 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_49
timestamp 1707688321
transform 1 0 16360 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_50
timestamp 1707688321
transform 1 0 15948 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_51
timestamp 1707688321
transform 1 0 16772 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_52
timestamp 1707688321
transform 1 0 17115 0 1 23745
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_53
timestamp 1707688321
transform 1 0 2617 0 1 23425
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_54
timestamp 1707688321
transform 1 0 14592 0 1 26964
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1707688321
transform 1 0 615 0 1 23932
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_1
timestamp 1707688321
transform 1 0 615 0 1 23529
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 1008 -1 0 4768
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 848 -1 0 4346
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 848 -1 0 4594
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 -1 928 -1 0 4470
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 -1 1088 -1 0 4892
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform -1 0 10948 0 -1 27483
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform -1 0 10905 0 -1 27563
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 0 -1 448 1 0 22459
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 0 -1 27 1 0 20497
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform 0 -1 448 1 0 20229
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform 0 -1 1142 1 0 23876
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform 0 -1 1302 1 0 23454
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform 0 -1 1302 1 0 23702
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform 0 -1 1382 1 0 23578
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform 0 -1 1222 1 0 24000
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 0 -1 1142 1 0 24124
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 0 -1 2928 1 0 26458
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 0 -1 10719 1 0 26714
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 0 -1 11031 1 0 26430
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 0 -1 11031 1 0 24027
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 0 -1 10719 1 0 24027
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 0 -1 288 1 0 22459
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 1 0 921 0 -1 5007
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 1 0 2657 0 1 23496
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 1 0 16956 0 1 23561
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1707688321
transform 1 0 4217 0 1 23656
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1707688321
transform 1 0 4217 0 1 23576
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1707688321
transform 1 0 7898 0 1 23736
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1707688321
transform 1 0 2605 0 1 23416
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1707688321
transform 1 0 6992 0 1 23736
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1707688321
transform 1 0 2657 0 1 23736
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1707688321
transform 1 0 4191 0 1 26955
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1707688321
transform 1 0 5049 0 1 26458
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1707688321
transform 1 0 660 0 1 25097
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 1 0 6633 0 1 27229
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1707688321
transform -1 0 13036 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1707688321
transform -1 0 8913 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1707688321
transform -1 0 17158 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1707688321
transform 1 0 6974 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_4
timestamp 1707688321
transform 1 0 6150 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_5
timestamp 1707688321
transform 1 0 7009 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_6
timestamp 1707688321
transform 1 0 7798 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_7
timestamp 1707688321
transform 1 0 5326 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_8
timestamp 1707688321
transform 1 0 9460 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_9
timestamp 1707688321
transform 1 0 10270 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_10
timestamp 1707688321
transform 1 0 11080 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_11
timestamp 1707688321
transform 1 0 11918 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_12
timestamp 1707688321
transform 1 0 12742 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_13
timestamp 1707688321
transform 1 0 15254 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_14
timestamp 1707688321
transform 1 0 16862 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_15
timestamp 1707688321
transform 1 0 16038 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_16
timestamp 1707688321
transform 1 0 15214 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_17
timestamp 1707688321
transform 1 0 4502 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_18
timestamp 1707688321
transform 1 0 14390 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_19
timestamp 1707688321
transform 1 0 8622 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_20
timestamp 1707688321
transform 1 0 13566 0 1 24216
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 1 0 3485 0 1 23416
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform -1 0 11452 0 1 26510
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 1 0 4985 0 1 27749
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 1 0 5809 0 1 27749
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1707688321
transform 1 0 6633 0 1 27749
box 0 0 192 180
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_0
timestamp 1707688321
transform 1 0 -214 0 1 22615
box 0 0 128 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1707688321
transform 1 0 5809 0 1 26458
box 0 0 192 372
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1707688321
transform 1 0 4478 0 1 27749
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_1
timestamp 1707688321
transform 1 0 5302 0 1 27749
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_2
timestamp 1707688321
transform 1 0 6126 0 1 27749
box 0 0 384 180
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 4478 0 1 27229
box 0 0 384 116
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1707688321
transform 1 0 4985 0 -1 26830
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_1
timestamp 1707688321
transform 1 0 14873 0 1 26093
box 0 0 192 308
use M1M2_CDNS_524688791851193  M1M2_CDNS_524688791851193_0
timestamp 1707688321
transform 1 0 6966 0 1 27749
box 0 0 704 180
use M1M2_CDNS_524688791851246  M1M2_CDNS_524688791851246_0
timestamp 1707688321
transform -1 0 11452 0 -1 26882
box 0 0 320 308
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_0
timestamp 1707688321
transform 1 0 12369 0 1 27800
box 0 0 704 116
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_1
timestamp 1707688321
transform 1 0 11131 0 1 27800
box 0 0 704 116
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_2
timestamp 1707688321
transform 1 0 15211 0 1 27800
box 0 0 704 116
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_3
timestamp 1707688321
transform 1 0 8246 0 1 27800
box 0 0 704 116
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_4
timestamp 1707688321
transform 1 0 16491 0 1 27800
box 0 0 704 116
use M1M2_CDNS_524688791851540  M1M2_CDNS_524688791851540_0
timestamp 1707688321
transform 1 0 3328 0 1 26093
box 0 0 768 308
use M1M2_CDNS_524688791851541  M1M2_CDNS_524688791851541_0
timestamp 1707688321
transform 1 0 7769 0 -1 26882
box 0 0 384 372
use M1M2_CDNS_524688791851541  M1M2_CDNS_524688791851541_1
timestamp 1707688321
transform 1 0 11892 0 -1 26882
box 0 0 384 372
use M1M2_CDNS_524688791851541  M1M2_CDNS_524688791851541_2
timestamp 1707688321
transform 1 0 16014 0 -1 26882
box 0 0 384 372
use M1M2_CDNS_524688791851541  M1M2_CDNS_524688791851541_3
timestamp 1707688321
transform 1 0 5302 0 1 26458
box 0 0 384 372
use M1M2_CDNS_524688791851541  M1M2_CDNS_524688791851541_4
timestamp 1707688321
transform 1 0 6126 0 1 26458
box 0 0 384 372
use M1M2_CDNS_524688791851542  M1M2_CDNS_524688791851542_0
timestamp 1707688321
transform 1 0 17601 0 1 26093
box 0 0 768 1076
use M1M2_CDNS_524688791851543  M1M2_CDNS_524688791851543_0
timestamp 1707688321
transform 1 0 17385 0 1 27749
box 0 0 960 180
use M1M2_CDNS_524688791851544  M1M2_CDNS_524688791851544_0
timestamp 1707688321
transform 1 0 9127 0 1 27749
box 0 0 1728 180
use M1M2_CDNS_524688791851544  M1M2_CDNS_524688791851544_1
timestamp 1707688321
transform 1 0 13252 0 1 27749
box 0 0 1728 180
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_0
timestamp 1707688321
transform 1 0 4160 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_1
timestamp 1707688321
transform 1 0 14048 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_2
timestamp 1707688321
transform 1 0 13224 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_3
timestamp 1707688321
transform 1 0 12400 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_4
timestamp 1707688321
transform 1 0 4984 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_5
timestamp 1707688321
transform 1 0 5808 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_6
timestamp 1707688321
transform 1 0 6632 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_7
timestamp 1707688321
transform 1 0 7456 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_8
timestamp 1707688321
transform 1 0 8280 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_9
timestamp 1707688321
transform 1 0 9104 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_10
timestamp 1707688321
transform 1 0 9928 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_11
timestamp 1707688321
transform 1 0 10752 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851545  M1M2_CDNS_524688791851545_12
timestamp 1707688321
transform 1 0 11576 0 1 24435
box 0 0 192 1524
use M1M2_CDNS_524688791851546  M1M2_CDNS_524688791851546_0
timestamp 1707688321
transform 1 0 6945 0 -1 26882
box 0 0 384 308
use M1M2_CDNS_524688791851546  M1M2_CDNS_524688791851546_1
timestamp 1707688321
transform 1 0 8593 0 -1 26882
box 0 0 384 308
use M1M2_CDNS_524688791851546  M1M2_CDNS_524688791851546_2
timestamp 1707688321
transform 1 0 12716 0 -1 26882
box 0 0 384 308
use M1M2_CDNS_524688791851546  M1M2_CDNS_524688791851546_3
timestamp 1707688321
transform 1 0 15190 0 -1 26882
box 0 0 384 308
use M1M2_CDNS_524688791851546  M1M2_CDNS_524688791851546_4
timestamp 1707688321
transform 1 0 16838 0 -1 26882
box 0 0 384 308
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_0
timestamp 1707688321
transform 1 0 8592 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_1
timestamp 1707688321
transform 1 0 6944 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_2
timestamp 1707688321
transform 1 0 9416 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_3
timestamp 1707688321
transform 1 0 10240 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_4
timestamp 1707688321
transform 1 0 11064 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_5
timestamp 1707688321
transform 1 0 11888 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_6
timestamp 1707688321
transform 1 0 7768 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_7
timestamp 1707688321
transform 1 0 12712 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_8
timestamp 1707688321
transform 1 0 6120 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_9
timestamp 1707688321
transform 1 0 16832 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_10
timestamp 1707688321
transform 1 0 5296 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_11
timestamp 1707688321
transform 1 0 16008 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_12
timestamp 1707688321
transform 1 0 15184 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_13
timestamp 1707688321
transform 1 0 14360 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_14
timestamp 1707688321
transform 1 0 4472 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851547  M1M2_CDNS_524688791851547_15
timestamp 1707688321
transform 1 0 13536 0 1 23896
box 0 -6 384 314
use M1M2_CDNS_524688791851548  M1M2_CDNS_524688791851548_0
timestamp 1707688321
transform 1 0 9110 0 1 27229
box 0 0 1280 116
use M1M2_CDNS_524688791851549  M1M2_CDNS_524688791851549_0
timestamp 1707688321
transform 1 0 13233 0 1 27229
box 0 0 1792 116
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_0
timestamp 1707688321
transform 1 0 9421 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_1
timestamp 1707688321
transform 1 0 10245 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_2
timestamp 1707688321
transform 1 0 4373 0 1 23900
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_3
timestamp 1707688321
transform 1 0 5301 0 1 23900
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_4
timestamp 1707688321
transform 1 0 6125 0 1 23900
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_5
timestamp 1707688321
transform 1 0 6949 0 1 23900
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_6
timestamp 1707688321
transform 1 0 7773 0 1 23900
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_7
timestamp 1707688321
transform 1 0 8597 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_8
timestamp 1707688321
transform 1 0 11069 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_9
timestamp 1707688321
transform 1 0 11893 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_10
timestamp 1707688321
transform 1 0 12717 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_11
timestamp 1707688321
transform 1 0 13541 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_12
timestamp 1707688321
transform 1 0 16837 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_13
timestamp 1707688321
transform 1 0 16013 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_14
timestamp 1707688321
transform 1 0 15189 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851550  M2M3_CDNS_524688791851550_15
timestamp 1707688321
transform 1 0 14365 0 1 23905
box -5 0 381 234
use M2M3_CDNS_524688791851551  M2M3_CDNS_524688791851551_0
timestamp 1707688321
transform 1 0 -214 0 1 22599
box -5 0 221 394
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_0
timestamp 1707688321
transform 1 0 6945 0 1 23899
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_1
timestamp 1707688321
transform 1 0 6121 0 1 23899
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_2
timestamp 1707688321
transform 1 0 5297 0 1 23899
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_3
timestamp 1707688321
transform 1 0 4369 0 1 23899
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_4
timestamp 1707688321
transform 1 0 7769 0 1 23899
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_5
timestamp 1707688321
transform 1 0 8593 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_6
timestamp 1707688321
transform 1 0 9417 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_7
timestamp 1707688321
transform 1 0 10241 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_8
timestamp 1707688321
transform 1 0 11065 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_9
timestamp 1707688321
transform 1 0 11889 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_10
timestamp 1707688321
transform 1 0 12713 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_11
timestamp 1707688321
transform 1 0 13537 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_12
timestamp 1707688321
transform 1 0 14361 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_13
timestamp 1707688321
transform 1 0 15185 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_14
timestamp 1707688321
transform 1 0 16009 0 1 23904
box -1 0 385 236
use M3M4_CDNS_524688791851539  M3M4_CDNS_524688791851539_15
timestamp 1707688321
transform 1 0 16833 0 1 23904
box -1 0 385 236
use nfet_CDNS_52468879185391  nfet_CDNS_52468879185391_0
timestamp 1707688321
transform 0 -1 1062 -1 0 4534
box -79 -26 335 626
use nfet_CDNS_52468879185391  nfet_CDNS_52468879185391_1
timestamp 1707688321
transform 0 -1 1062 1 0 4700
box -79 -26 335 626
use pEsdFet_CDNS_524688791851555  pEsdFet_CDNS_524688791851555_0
timestamp 1707688321
transform 1 0 4408 0 1 23827
box -1484 -840 14366 3940
use pfet_CDNS_52468879185397  pfet_CDNS_52468879185397_0
timestamp 1707688321
transform 0 -1 1672 -1 0 23770
box -119 -66 375 1066
use pfet_CDNS_52468879185397  pfet_CDNS_52468879185397_1
timestamp 1707688321
transform 0 -1 1672 1 0 23936
box -119 -66 375 1066
use PYbentRes_CDNS_524688791851554  PYbentRes_CDNS_524688791851554_0
timestamp 1707688321
transform 0 -1 2854 1 0 23333
box -50 0 2090 100
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1707688321
transform 0 -1 2837 -1 0 25491
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1707688321
transform 0 -1 2837 1 0 23215
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 11812 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 11400 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 1 13048 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 13460 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 1 12636 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 1 12224 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 1 7692 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 1 8516 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 0 1 8104 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1707688321
transform 0 1 9752 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1707688321
transform 0 1 10164 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1707688321
transform 0 1 9340 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_12
timestamp 1707688321
transform 0 1 8928 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_13
timestamp 1707688321
transform 0 1 6044 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_14
timestamp 1707688321
transform 0 1 6456 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_15
timestamp 1707688321
transform 0 1 7280 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_16
timestamp 1707688321
transform 0 1 6868 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_17
timestamp 1707688321
transform 0 1 5220 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_18
timestamp 1707688321
transform 0 1 5632 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_19
timestamp 1707688321
transform 0 1 4808 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_20
timestamp 1707688321
transform 0 1 4396 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_21
timestamp 1707688321
transform 0 1 10988 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_22
timestamp 1707688321
transform 0 1 10576 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_23
timestamp 1707688321
transform 0 1 13872 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_24
timestamp 1707688321
transform 0 1 14284 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_25
timestamp 1707688321
transform 0 1 14696 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_26
timestamp 1707688321
transform 0 1 14284 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_27
timestamp 1707688321
transform 0 1 10988 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_28
timestamp 1707688321
transform 0 1 11400 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_29
timestamp 1707688321
transform 0 1 12224 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_30
timestamp 1707688321
transform 0 1 11812 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_31
timestamp 1707688321
transform 0 1 13460 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_32
timestamp 1707688321
transform 0 1 13872 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_33
timestamp 1707688321
transform 0 1 13048 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_34
timestamp 1707688321
transform 0 1 12636 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_35
timestamp 1707688321
transform 0 1 7692 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_36
timestamp 1707688321
transform 0 1 8104 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_37
timestamp 1707688321
transform 0 1 8928 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_38
timestamp 1707688321
transform 0 1 8516 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_39
timestamp 1707688321
transform 0 1 10164 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_40
timestamp 1707688321
transform 0 1 10576 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_41
timestamp 1707688321
transform 0 1 9752 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_42
timestamp 1707688321
transform 0 1 9340 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_43
timestamp 1707688321
transform 0 1 6044 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_44
timestamp 1707688321
transform 0 1 6456 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_45
timestamp 1707688321
transform 0 1 7280 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_46
timestamp 1707688321
transform 0 1 6868 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_47
timestamp 1707688321
transform 0 1 5220 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_48
timestamp 1707688321
transform 0 1 5632 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_49
timestamp 1707688321
transform 0 1 4808 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_50
timestamp 1707688321
transform 0 1 4396 1 0 26959
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_51
timestamp 1707688321
transform 0 1 14696 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_52
timestamp 1707688321
transform 0 1 16344 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_53
timestamp 1707688321
transform 0 1 16756 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_54
timestamp 1707688321
transform 0 1 17168 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_55
timestamp 1707688321
transform 0 1 15932 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_56
timestamp 1707688321
transform 0 1 15520 1 0 23729
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_57
timestamp 1707688321
transform 0 1 15108 1 0 23729
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 1 0 374 0 1 4686
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1707688321
transform 1 0 374 0 1 4278
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_2
timestamp 1707688321
transform 1 0 574 0 1 23922
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_3
timestamp 1707688321
transform 1 0 574 0 1 23514
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1707688321
transform -1 0 11624 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1707688321
transform -1 0 6801 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_2
timestamp 1707688321
transform -1 0 12690 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_3
timestamp 1707688321
transform -1 0 13514 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_4
timestamp 1707688321
transform -1 0 14508 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_5
timestamp 1707688321
transform 1 0 11722 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_6
timestamp 1707688321
transform 1 0 8717 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_7
timestamp 1707688321
transform 1 0 12304 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_8
timestamp 1707688321
transform 1 0 13128 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_9
timestamp 1707688321
transform 1 0 13782 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1707688321
transform 1 0 14895 0 1 23739
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1707688321
transform -1 0 11454 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1707688321
transform -1 0 4741 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_2
timestamp 1707688321
transform -1 0 5153 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_3
timestamp 1707688321
transform -1 0 5565 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_4
timestamp 1707688321
transform -1 0 5977 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_5
timestamp 1707688321
transform -1 0 6389 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_6
timestamp 1707688321
transform -1 0 7213 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_7
timestamp 1707688321
transform -1 0 7625 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_8
timestamp 1707688321
transform -1 0 7942 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_9
timestamp 1707688321
transform -1 0 12860 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_10
timestamp 1707688321
transform -1 0 13684 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_11
timestamp 1707688321
transform -1 0 14338 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_12
timestamp 1707688321
transform -1 0 2877 0 1 23496
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_13
timestamp 1707688321
transform -1 0 2877 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_14
timestamp 1707688321
transform 1 0 11892 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_15
timestamp 1707688321
transform 1 0 7987 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_16
timestamp 1707688321
transform 1 0 8305 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_17
timestamp 1707688321
transform 1 0 9129 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_18
timestamp 1707688321
transform 1 0 9541 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_19
timestamp 1707688321
transform 1 0 9953 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_20
timestamp 1707688321
transform 1 0 10365 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_21
timestamp 1707688321
transform 1 0 10777 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_22
timestamp 1707688321
transform 1 0 12134 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_23
timestamp 1707688321
transform 1 0 12958 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_24
timestamp 1707688321
transform 1 0 13952 0 1 23736
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1707688321
transform 1 0 15843 0 -1 23785
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_1
timestamp 1707688321
transform 1 0 16667 0 -1 23785
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_2
timestamp 1707688321
transform 1 0 16838 0 -1 23785
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_3
timestamp 1707688321
transform 1 0 16244 0 -1 23785
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_0
timestamp 1707688321
transform 0 1 16956 1 0 23573
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851552  sky130_fd_io__tk_em1s_CDNS_524688791851552_0
timestamp 1707688321
transform 0 1 15693 -1 0 27024
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851552  sky130_fd_io__tk_em1s_CDNS_524688791851552_1
timestamp 1707688321
transform 0 1 16517 -1 0 27024
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851553  sky130_fd_io__tk_em1s_CDNS_524688791851553_0
timestamp 1707688321
transform -1 0 17634 0 1 23874
box 0 0 1 1
<< labels >>
flabel comment s 9717 22945 9717 22945 0 FreeSans 300 0 0 0 pug<0>
flabel comment s 10138 22956 10138 22956 0 FreeSans 300 0 0 0 pug<1>
flabel comment s 842 25124 842 25124 0 FreeSans 300 90 0 0 nghs_h
flabel comment s 17028 23886 17028 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 16204 23886 16204 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 15380 23886 15380 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 14556 23886 14556 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 13732 23886 13732 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 12908 23886 12908 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 12084 23886 12084 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 11260 23886 11260 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 10436 23886 10436 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 9612 23886 9612 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 8788 23886 8788 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 7964 23886 7964 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 7140 23886 7140 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 6316 23886 6316 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 5492 23886 5492 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 4668 23886 4668 23886 0 FreeSans 200 0 0 0 pad
flabel comment s 17439 23886 17439 23886 0 FreeSans 200 0 0 0 vpb_drvr
flabel comment s 16630 23886 16630 23886 0 FreeSans 200 0 0 0 vpb_drvr
flabel comment s 15795 23886 15795 23886 0 FreeSans 200 0 0 0 vpb_drvr
flabel comment s 14969 23886 14969 23886 0 FreeSans 200 0 0 0 vpb_drvr
flabel comment s 14140 23886 14140 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 13317 23886 13317 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 12493 23886 12493 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 11678 23886 11678 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 10844 23886 10844 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 7566 23886 7566 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 8390 23886 8390 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 10040 23886 10040 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 9216 23886 9216 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 5908 23886 5908 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 6732 23886 6732 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 5082 23886 5082 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 4258 23886 4258 23886 0 FreeSans 200 0 0 0 vcc_io
flabel comment s 4280 23688 4280 23688 0 FreeSans 200 0 0 0 pug<2>
flabel comment s 663 16908 663 16908 0 FreeSans 100 0 0 0 pu_h_n<1>
flabel comment s 517 23300 517 23300 0 FreeSans 100 0 0 0 pu_h_n<0>
flabel comment s 952 23293 952 23293 0 FreeSans 100 0 0 0 pu_h_n<1>
flabel comment s 1115 23293 1115 23293 0 FreeSans 100 0 0 0 pu_h_n<2>
flabel comment s 1276 23292 1276 23292 0 FreeSans 100 0 0 0 pu_h_n<3>
flabel comment s 719 23298 719 23298 0 FreeSans 100 0 0 0 pug<0>
flabel comment s 1033 23294 1033 23294 0 FreeSans 100 0 0 0 pug<1>
flabel comment s 1193 23291 1193 23291 0 FreeSans 100 0 0 0 pug<2>
flabel comment s 189 16908 189 16908 0 FreeSans 100 0 0 0 pu_h_n<0>
flabel comment s 794 23285 794 23285 0 FreeSans 100 90 0 0 pad_weak
flabel comment s 786 4758 786 4758 0 FreeSans 200 0 0 0 I183
flabel comment s 779 4902 779 4902 0 FreeSans 200 0 0 0 I183
flabel comment s 576 17018 576 17018 0 FreeSans 200 90 0 0 pad_strong_slow
flabel comment s 497 16962 497 16962 0 FreeSans 200 90 0 0 pad_weak
flabel comment s 14525 23686 14525 23686 0 FreeSans 200 0 0 0 pug<2>
flabel comment s 4280 23604 4280 23604 0 FreeSans 200 0 0 0 pug<3>
flabel comment s 420 16903 420 16903 0 FreeSans 100 0 0 0 nghs
flabel comment s 340 16902 340 16902 0 FreeSans 100 0 0 0 pghs
flabel comment s 1063 16909 1063 16909 0 FreeSans 100 0 0 0 pug<3>
flabel comment s 901 16908 901 16908 0 FreeSans 100 0 0 0 pug<2>
flabel comment s 743 16907 743 16907 0 FreeSans 100 0 0 0 pug<1>
flabel comment s 267 16908 267 16908 0 FreeSans 100 0 0 0 pug<0>
flabel comment s 985 16908 985 16908 0 FreeSans 100 0 0 0 pu_h_n<3>
flabel comment s 822 16908 822 16908 0 FreeSans 100 0 0 0 pu_h_n<2>
flabel comment s 873 23263 873 23263 0 FreeSans 100 90 0 0 pad_strong_slow
flabel comment s 1062 24135 1062 24135 0 FreeSans 200 0 0 0 I48
flabel comment s 1059 23983 1059 23983 0 FreeSans 200 0 0 0 I48
flabel comment s 1059 23712 1059 23712 0 FreeSans 200 0 0 0 I184
flabel comment s 1052 23568 1052 23568 0 FreeSans 200 0 0 0 I184
flabel comment s 789 17033 789 17033 0 FreeSans 200 0 0 0 I49
flabel comment s 786 17185 786 17185 0 FreeSans 200 0 0 0 I49
flabel comment s 786 17456 786 17456 0 FreeSans 200 0 0 0 I183
flabel comment s 779 17600 779 17600 0 FreeSans 200 0 0 0 I183
flabel comment s 14353 23698 14353 23698 0 FreeSans 400 0 0 0 <19.8>
flabel comment s 13941 23698 13941 23698 0 FreeSans 400 0 0 0 <19.7>
flabel comment s 13534 23698 13534 23698 0 FreeSans 400 0 0 0 <19.6>
flabel comment s 13122 23698 13122 23698 0 FreeSans 400 0 0 0 <19.5>
flabel comment s 12706 23698 12706 23698 0 FreeSans 400 0 0 0 <19.4>
flabel comment s 12297 23698 12297 23698 0 FreeSans 400 0 0 0 <19.3>
flabel comment s 11882 23698 11882 23698 0 FreeSans 400 0 0 0 <19.2>
flabel comment s 11467 23698 11467 23698 0 FreeSans 400 0 0 0 <19.1>
flabel comment s 14767 23761 14767 23761 0 FreeSans 400 0 0 0 <18>
flabel comment s 7753 23698 7753 23698 0 FreeSans 400 0 0 0 <17>
flabel comment s 11053 23698 11053 23698 0 FreeSans 400 0 0 0 <16>
flabel comment s 10632 23698 10632 23698 0 FreeSans 400 0 0 0 <15>
flabel comment s 10222 23698 10222 23698 0 FreeSans 400 0 0 0 <14>
flabel comment s 9809 23698 9809 23698 0 FreeSans 400 0 0 0 <13>
flabel comment s 9405 23698 9405 23698 0 FreeSans 400 0 0 0 <12>
flabel comment s 8990 23698 8990 23698 0 FreeSans 400 0 0 0 <11>
flabel comment s 8576 23698 8576 23698 0 FreeSans 400 0 0 0 <10>
flabel comment s 8164 23698 8164 23698 0 FreeSans 400 0 0 0 <9>
flabel comment s 7344 23698 7344 23698 0 FreeSans 400 0 0 0 <8>
flabel comment s 6937 23698 6937 23698 0 FreeSans 400 0 0 0 <7>
flabel comment s 6530 23698 6530 23698 0 FreeSans 400 0 0 0 <6>
flabel comment s 6105 23698 6105 23698 0 FreeSans 400 0 0 0 <5>
flabel comment s 5697 23698 5697 23698 0 FreeSans 400 0 0 0 <4>
flabel comment s 5287 23698 5287 23698 0 FreeSans 400 0 0 0 <3>
flabel comment s 4875 23698 4875 23698 0 FreeSans 400 0 0 0 <2>
flabel comment s 4465 23698 4465 23698 0 FreeSans 400 0 0 0 <1>
flabel comment s 1357 23296 1357 23296 0 FreeSans 100 0 0 0 pug<3>
flabel comment s 636 23286 636 23286 0 FreeSans 100 0 0 0 pghs
flabel metal1 s 4477 23877 4861 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 2669 23524 2669 23524 0 FreeSans 200 0 0 0 tie_hi_opt
flabel metal1 s 2901 23983 2901 23983 0 FreeSans 200 0 0 0 tie_hi
flabel metal1 s 7756 23762 7756 23762 0 FreeSans 200 0 0 0 p17g
flabel metal1 s 10640 23765 10640 23765 0 FreeSans 200 0 0 0 p15g
flabel metal1 s 10232 23761 10232 23761 0 FreeSans 200 0 0 0 p14g
flabel metal1 s 9817 23760 9817 23760 0 FreeSans 200 0 0 0 p13g
flabel metal1 s 9404 23762 9404 23762 0 FreeSans 200 0 0 0 p12g
flabel metal1 s 8996 23761 8996 23761 0 FreeSans 200 0 0 0 p11g
flabel metal1 s 8584 23763 8584 23763 0 FreeSans 200 0 0 0 p10g
flabel metal1 s 8174 23763 8174 23763 0 FreeSans 200 0 0 0 p9g
flabel metal1 s 7346 23761 7346 23761 0 FreeSans 200 0 0 0 p8g
flabel metal1 s 6935 23759 6935 23759 0 FreeSans 200 0 0 0 p7g
flabel metal1 s 6520 23760 6520 23760 0 FreeSans 200 0 0 0 p6g
flabel metal1 s 6106 23765 6106 23765 0 FreeSans 200 0 0 0 p5g
flabel metal1 s 5698 23765 5698 23765 0 FreeSans 200 0 0 0 p4g
flabel metal1 s 5287 23762 5287 23762 0 FreeSans 200 0 0 0 p3g
flabel metal1 s 4875 23763 4875 23763 0 FreeSans 200 0 0 0 p2g
flabel metal1 s 14363 23877 14747 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 15187 23877 15571 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 16011 23877 16395 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 16835 23877 17219 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 4983 23892 5178 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 5807 23892 6002 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 6631 23892 6826 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 7455 23892 7650 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 8279 23892 8474 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 9103 23892 9298 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 9927 23892 10122 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 10751 23892 10946 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 11575 23892 11770 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 12399 23892 12594 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 13223 23892 13418 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 14047 23892 14242 23976 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 17855 23553 18076 23653 0 FreeSans 200 0 0 0 vpb_drvr
port 6 nsew
flabel metal1 s 5299 23877 5683 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 10243 23877 10627 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 11891 23877 12275 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 6123 23877 6507 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 7771 23877 8155 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 13539 23877 13923 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 11067 23877 11451 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 9419 23877 9803 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 6947 23877 7331 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 8595 23877 8979 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 12715 23877 13099 23973 0 FreeSans 200 0 0 0 pad
port 2 nsew
flabel metal1 s 610 23638 653 23662 0 FreeSans 200 0 0 0 pghs_h<3>
port 4 nsew
flabel metal1 s 612 24043 647 24069 0 FreeSans 200 0 0 0 pghs_h<2>
port 5 nsew
flabel locali s 1758 23958 1792 24179 0 FreeSans 200 90 0 0 vpb_drvr
port 6 nsew
flabel locali s 382 4449 429 4476 0 FreeSans 200 0 0 0 nghs_h<2>
port 7 nsew
flabel locali s 1277 4189 1395 4235 0 FreeSans 200 0 0 0 vgnd_io
port 8 nsew
flabel locali s 382 4760 429 4787 0 FreeSans 200 0 0 0 nghs_h<3>
port 9 nsew
flabel metal2 s 17629 22523 18369 22563 0 FreeSans 200 0 0 0 vpb_drvr
port 6 nsew
flabel metal2 s 16956 22872 17084 22912 0 FreeSans 200 0 0 0 p2gate
port 10 nsew
flabel metal2 s 13976 22523 14304 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 13152 22523 13480 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 12328 22523 12656 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 11504 22523 11832 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 9032 22523 9360 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 8208 22523 8536 22563 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal2 s 796 19152 848 19162 0 FreeSans 100 0 0 0 pu_h_n<2>
port 11 nsew
flabel metal2 s 956 19152 1008 19162 0 FreeSans 100 0 0 0 pu_h_n<3>
port 12 nsew
flabel metal2 s 876 19152 928 19162 0 FreeSans 100 0 0 0 pug<2>
port 13 nsew
flabel metal2 s 1036 19152 1088 19162 0 FreeSans 100 0 0 0 pug<3>
port 14 nsew
flabel metal2 s 17117 23218 17167 23258 0 FreeSans 200 0 0 0 vcc_io_soft
port 15 nsew
<< properties >>
string GDS_END 91954012
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91767150
string path 421.350 589.300 421.350 592.525 
<< end >>
