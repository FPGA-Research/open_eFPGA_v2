magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 1175 157 1357 201
rect 1660 157 2196 203
rect 1 145 825 157
rect 1029 145 2196 157
rect 1 21 2196 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 355 47 385 131
rect 457 47 487 131
rect 535 47 565 131
rect 631 47 661 131
rect 707 47 737 131
rect 911 47 941 119
rect 1007 47 1037 119
rect 1105 47 1135 131
rect 1251 47 1281 175
rect 1352 47 1382 119
rect 1455 47 1485 119
rect 1550 47 1580 131
rect 1738 47 1768 177
rect 1833 47 1863 177
rect 1917 47 1947 177
rect 2003 47 2033 177
rect 2087 47 2117 177
<< scpmoshvt >>
rect 80 363 110 491
rect 164 363 194 491
rect 352 369 382 497
rect 436 369 466 497
rect 530 369 560 497
rect 614 369 644 497
rect 707 369 737 497
rect 910 413 940 497
rect 1003 413 1033 497
rect 1099 413 1129 497
rect 1231 347 1261 497
rect 1326 413 1356 497
rect 1410 413 1440 497
rect 1527 413 1557 497
rect 1738 297 1768 497
rect 1833 297 1863 497
rect 1917 297 1947 497
rect 2003 297 2033 497
rect 2087 297 2117 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 89 355 131
rect 299 55 311 89
rect 345 55 355 89
rect 299 47 355 55
rect 385 89 457 131
rect 385 55 411 89
rect 445 55 457 89
rect 385 47 457 55
rect 487 47 535 131
rect 565 89 631 131
rect 565 55 586 89
rect 620 55 631 89
rect 565 47 631 55
rect 661 47 707 131
rect 737 89 799 131
rect 1201 131 1251 175
rect 1055 119 1105 131
rect 737 55 753 89
rect 787 55 799 89
rect 737 47 799 55
rect 855 107 911 119
rect 855 73 863 107
rect 897 73 911 107
rect 855 47 911 73
rect 941 107 1007 119
rect 941 73 963 107
rect 997 73 1007 107
rect 941 47 1007 73
rect 1037 47 1105 119
rect 1135 101 1251 131
rect 1135 67 1179 101
rect 1213 67 1251 101
rect 1135 47 1251 67
rect 1281 119 1331 175
rect 1686 162 1738 177
rect 1500 119 1550 131
rect 1281 107 1352 119
rect 1281 73 1297 107
rect 1331 73 1352 107
rect 1281 47 1352 73
rect 1382 107 1455 119
rect 1382 73 1409 107
rect 1443 73 1455 107
rect 1382 47 1455 73
rect 1485 47 1550 119
rect 1580 107 1632 131
rect 1580 73 1590 107
rect 1624 73 1632 107
rect 1580 47 1632 73
rect 1686 128 1694 162
rect 1728 128 1738 162
rect 1686 94 1738 128
rect 1686 60 1694 94
rect 1728 60 1738 94
rect 1686 47 1738 60
rect 1768 123 1833 177
rect 1768 89 1785 123
rect 1819 89 1833 123
rect 1768 47 1833 89
rect 1863 164 1917 177
rect 1863 130 1873 164
rect 1907 130 1917 164
rect 1863 96 1917 130
rect 1863 62 1873 96
rect 1907 62 1917 96
rect 1863 47 1917 62
rect 1947 96 2003 177
rect 1947 62 1959 96
rect 1993 62 2003 96
rect 1947 47 2003 62
rect 2033 164 2087 177
rect 2033 130 2043 164
rect 2077 130 2087 164
rect 2033 96 2087 130
rect 2033 62 2043 96
rect 2077 62 2087 96
rect 2033 47 2087 62
rect 2117 96 2170 177
rect 2117 62 2127 96
rect 2161 62 2170 96
rect 2117 47 2170 62
<< pdiff >>
rect 28 477 80 491
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 363 80 375
rect 110 461 164 491
rect 110 427 120 461
rect 154 427 164 461
rect 110 363 164 427
rect 194 477 246 491
rect 194 443 204 477
rect 238 443 246 477
rect 194 409 246 443
rect 194 375 204 409
rect 238 375 246 409
rect 194 363 246 375
rect 300 452 352 497
rect 300 418 308 452
rect 342 418 352 452
rect 300 369 352 418
rect 382 483 436 497
rect 382 449 392 483
rect 426 449 436 483
rect 382 369 436 449
rect 466 369 530 497
rect 560 483 614 497
rect 560 449 570 483
rect 604 449 614 483
rect 560 369 614 449
rect 644 369 707 497
rect 737 483 794 497
rect 737 449 752 483
rect 786 449 794 483
rect 737 369 794 449
rect 848 472 910 497
rect 848 438 856 472
rect 890 438 910 472
rect 848 413 910 438
rect 940 472 1003 497
rect 940 438 955 472
rect 989 438 1003 472
rect 940 413 1003 438
rect 1033 413 1099 497
rect 1129 485 1231 497
rect 1129 451 1187 485
rect 1221 451 1231 485
rect 1129 417 1231 451
rect 1129 413 1187 417
rect 1144 383 1187 413
rect 1221 383 1231 417
rect 1144 347 1231 383
rect 1261 477 1326 497
rect 1261 443 1271 477
rect 1305 443 1326 477
rect 1261 413 1326 443
rect 1356 467 1410 497
rect 1356 433 1366 467
rect 1400 433 1410 467
rect 1356 413 1410 433
rect 1440 413 1527 497
rect 1557 477 1632 497
rect 1557 443 1589 477
rect 1623 443 1632 477
rect 1557 413 1632 443
rect 1686 475 1738 497
rect 1686 441 1694 475
rect 1728 441 1738 475
rect 1261 347 1311 413
rect 1686 407 1738 441
rect 1686 373 1694 407
rect 1728 373 1738 407
rect 1686 297 1738 373
rect 1768 455 1833 497
rect 1768 421 1785 455
rect 1819 421 1833 455
rect 1768 375 1833 421
rect 1768 341 1785 375
rect 1819 341 1833 375
rect 1768 297 1833 341
rect 1863 479 1917 497
rect 1863 445 1873 479
rect 1907 445 1917 479
rect 1863 411 1917 445
rect 1863 377 1873 411
rect 1907 377 1917 411
rect 1863 343 1917 377
rect 1863 309 1873 343
rect 1907 309 1917 343
rect 1863 297 1917 309
rect 1947 487 2003 497
rect 1947 453 1959 487
rect 1993 453 2003 487
rect 1947 419 2003 453
rect 1947 385 1959 419
rect 1993 385 2003 419
rect 1947 297 2003 385
rect 2033 479 2087 497
rect 2033 445 2043 479
rect 2077 445 2087 479
rect 2033 411 2087 445
rect 2033 377 2043 411
rect 2077 377 2087 411
rect 2033 343 2087 377
rect 2033 309 2043 343
rect 2077 309 2087 343
rect 2033 297 2087 309
rect 2117 487 2175 497
rect 2117 453 2127 487
rect 2161 453 2175 487
rect 2117 419 2175 453
rect 2117 385 2127 419
rect 2161 385 2175 419
rect 2117 297 2175 385
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 311 55 345 89
rect 411 55 445 89
rect 586 55 620 89
rect 753 55 787 89
rect 863 73 897 107
rect 963 73 997 107
rect 1179 67 1213 101
rect 1297 73 1331 107
rect 1409 73 1443 107
rect 1590 73 1624 107
rect 1694 128 1728 162
rect 1694 60 1728 94
rect 1785 89 1819 123
rect 1873 130 1907 164
rect 1873 62 1907 96
rect 1959 62 1993 96
rect 2043 130 2077 164
rect 2043 62 2077 96
rect 2127 62 2161 96
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 120 427 154 461
rect 204 443 238 477
rect 204 375 238 409
rect 308 418 342 452
rect 392 449 426 483
rect 570 449 604 483
rect 752 449 786 483
rect 856 438 890 472
rect 955 438 989 472
rect 1187 451 1221 485
rect 1187 383 1221 417
rect 1271 443 1305 477
rect 1366 433 1400 467
rect 1589 443 1623 477
rect 1694 441 1728 475
rect 1694 373 1728 407
rect 1785 421 1819 455
rect 1785 341 1819 375
rect 1873 445 1907 479
rect 1873 377 1907 411
rect 1873 309 1907 343
rect 1959 453 1993 487
rect 1959 385 1993 419
rect 2043 445 2077 479
rect 2043 377 2077 411
rect 2043 309 2077 343
rect 2127 453 2161 487
rect 2127 385 2161 419
<< poly >>
rect 80 491 110 517
rect 164 491 194 517
rect 352 497 382 523
rect 436 497 466 523
rect 530 497 560 523
rect 614 497 644 523
rect 707 497 737 523
rect 910 497 940 523
rect 1003 497 1033 523
rect 1099 497 1129 523
rect 1231 497 1261 523
rect 1326 497 1356 523
rect 1410 497 1440 523
rect 1527 497 1557 523
rect 1738 497 1768 523
rect 1833 497 1863 523
rect 1917 497 1947 523
rect 2003 497 2033 523
rect 2087 497 2117 523
rect 910 375 940 413
rect 1003 381 1033 413
rect 80 348 110 363
rect 47 318 110 348
rect 47 265 77 318
rect 164 274 194 363
rect 352 331 382 369
rect 436 331 466 369
rect 530 337 560 369
rect 614 337 644 369
rect 340 321 466 331
rect 340 287 356 321
rect 390 301 466 321
rect 515 321 569 337
rect 390 287 406 301
rect 340 277 406 287
rect 515 287 525 321
rect 559 287 569 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 194 274
rect 119 230 135 264
rect 169 230 194 264
rect 119 220 194 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 355 131 385 277
rect 515 271 569 287
rect 611 321 665 337
rect 611 287 621 321
rect 655 287 665 321
rect 611 271 665 287
rect 707 304 737 369
rect 895 365 961 375
rect 895 331 911 365
rect 945 331 961 365
rect 895 321 961 331
rect 1003 365 1057 381
rect 1003 331 1013 365
rect 1047 331 1057 365
rect 1003 315 1057 331
rect 707 288 761 304
rect 427 225 493 235
rect 427 191 443 225
rect 477 191 493 225
rect 427 181 493 191
rect 457 131 487 181
rect 535 131 565 271
rect 707 254 717 288
rect 751 254 761 288
rect 1003 279 1033 315
rect 707 238 761 254
rect 911 249 1033 279
rect 607 207 661 223
rect 607 173 617 207
rect 651 173 661 207
rect 607 157 661 173
rect 631 131 661 157
rect 707 131 737 238
rect 911 119 941 249
rect 1099 213 1129 413
rect 1231 309 1261 347
rect 1326 315 1356 413
rect 1410 375 1440 413
rect 1527 381 1557 413
rect 1409 365 1475 375
rect 1409 331 1425 365
rect 1459 331 1475 365
rect 1409 321 1475 331
rect 1527 365 1605 381
rect 1527 331 1561 365
rect 1595 331 1605 365
rect 1527 315 1605 331
rect 1171 299 1261 309
rect 1171 265 1187 299
rect 1221 265 1261 299
rect 1171 255 1261 265
rect 1231 220 1261 255
rect 1313 299 1367 315
rect 1313 265 1323 299
rect 1357 279 1367 299
rect 1357 265 1485 279
rect 1313 249 1485 265
rect 983 191 1037 207
rect 983 157 993 191
rect 1027 157 1037 191
rect 1099 203 1179 213
rect 1099 183 1129 203
rect 983 141 1037 157
rect 1007 119 1037 141
rect 1105 169 1129 183
rect 1163 169 1179 203
rect 1231 190 1281 220
rect 1251 175 1281 190
rect 1352 191 1413 207
rect 1105 159 1179 169
rect 1105 131 1135 159
rect 1352 157 1369 191
rect 1403 157 1413 191
rect 1352 141 1413 157
rect 1352 119 1382 141
rect 1455 119 1485 249
rect 1550 131 1580 315
rect 1738 265 1768 297
rect 1636 249 1768 265
rect 1636 215 1646 249
rect 1680 215 1768 249
rect 1636 199 1768 215
rect 1738 177 1768 199
rect 1833 265 1863 297
rect 1917 265 1947 297
rect 2003 265 2033 297
rect 2087 265 2117 297
rect 1833 249 2117 265
rect 1833 215 1843 249
rect 1877 215 1911 249
rect 1945 215 1979 249
rect 2013 215 2047 249
rect 2081 215 2117 249
rect 1833 199 2117 215
rect 1833 177 1863 199
rect 1917 177 1947 199
rect 2003 177 2033 199
rect 2087 177 2117 199
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 457 21 487 47
rect 535 21 565 47
rect 631 21 661 47
rect 707 21 737 47
rect 911 21 941 47
rect 1007 21 1037 47
rect 1105 21 1135 47
rect 1251 21 1281 47
rect 1352 21 1382 47
rect 1455 21 1485 47
rect 1550 21 1580 47
rect 1738 21 1768 47
rect 1833 21 1863 47
rect 1917 21 1947 47
rect 2003 21 2033 47
rect 2087 21 2117 47
<< polycont >>
rect 356 287 390 321
rect 525 287 559 321
rect 33 215 67 249
rect 135 230 169 264
rect 621 287 655 321
rect 911 331 945 365
rect 1013 331 1047 365
rect 443 191 477 225
rect 717 254 751 288
rect 617 173 651 207
rect 1425 331 1459 365
rect 1561 331 1595 365
rect 1187 265 1221 299
rect 1323 265 1357 299
rect 993 157 1027 191
rect 1129 169 1163 203
rect 1369 157 1403 191
rect 1646 215 1680 249
rect 1843 215 1877 249
rect 1911 215 1945 249
rect 1979 215 2013 249
rect 2047 215 2081 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 170 527
rect 104 427 120 461
rect 154 427 170 461
rect 204 477 249 493
rect 238 443 249 477
rect 204 409 249 443
rect 70 391 169 393
rect 70 375 123 391
rect 36 359 123 375
rect 157 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 194 169 230
rect 238 375 249 409
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 249 375
rect 204 153 211 187
rect 245 153 249 187
rect 204 143 249 153
rect 35 119 69 127
rect 203 119 249 143
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 249 119
rect 203 69 249 85
rect 287 452 342 489
rect 287 418 308 452
rect 376 483 442 527
rect 752 483 786 527
rect 376 449 392 483
rect 426 449 442 483
rect 539 449 570 483
rect 604 449 718 483
rect 287 415 342 418
rect 287 372 650 415
rect 287 89 321 372
rect 356 321 390 337
rect 356 157 390 287
rect 424 225 458 372
rect 616 337 650 372
rect 684 399 718 449
rect 752 433 786 449
rect 843 472 890 488
rect 1187 485 1221 527
rect 843 438 856 472
rect 939 438 955 472
rect 989 438 1153 472
rect 843 413 890 438
rect 843 399 877 413
rect 684 365 877 399
rect 997 391 1085 402
rect 492 321 559 337
rect 492 287 525 321
rect 492 271 559 287
rect 616 321 655 337
rect 616 287 621 321
rect 616 271 655 287
rect 707 288 805 331
rect 707 254 717 288
rect 751 254 805 288
rect 424 191 443 225
rect 477 191 493 225
rect 617 207 651 223
rect 707 207 805 254
rect 843 173 877 365
rect 617 157 651 173
rect 356 123 651 157
rect 685 139 877 173
rect 911 365 959 381
rect 945 331 959 365
rect 997 365 1043 391
rect 997 331 1013 365
rect 1077 357 1085 391
rect 1047 331 1085 357
rect 911 207 959 331
rect 1119 315 1153 438
rect 1187 417 1221 451
rect 1187 367 1221 383
rect 1255 477 1305 493
rect 1255 443 1271 477
rect 1563 477 1624 527
rect 1255 427 1305 443
rect 1350 433 1366 467
rect 1400 433 1527 467
rect 1119 299 1221 315
rect 1119 297 1187 299
rect 1061 265 1187 297
rect 1061 263 1221 265
rect 911 191 1027 207
rect 911 187 993 191
rect 911 153 951 187
rect 985 157 993 187
rect 985 153 1027 157
rect 911 141 1027 153
rect 103 17 169 59
rect 287 55 311 89
rect 345 55 361 89
rect 395 55 411 89
rect 445 55 461 89
rect 495 61 530 123
rect 685 89 719 139
rect 843 107 877 139
rect 1061 107 1095 263
rect 1187 249 1221 263
rect 1129 213 1163 219
rect 1255 213 1289 427
rect 1323 391 1361 393
rect 1323 357 1325 391
rect 1359 357 1361 391
rect 1323 299 1361 357
rect 1357 265 1361 299
rect 1323 249 1361 265
rect 1395 365 1459 381
rect 1395 331 1425 365
rect 1395 315 1459 331
rect 1129 203 1289 213
rect 1395 207 1433 315
rect 1493 281 1527 433
rect 1563 443 1589 477
rect 1623 443 1624 477
rect 1563 427 1624 443
rect 1694 475 1751 491
rect 1728 441 1751 475
rect 1694 407 1751 441
rect 1561 373 1694 381
rect 1728 373 1751 407
rect 1561 365 1751 373
rect 1595 331 1751 365
rect 1561 315 1751 331
rect 1785 455 1821 527
rect 1959 487 1993 527
rect 1819 421 1821 455
rect 1785 375 1821 421
rect 1819 341 1821 375
rect 1785 325 1821 341
rect 1857 445 1873 479
rect 1907 445 1923 479
rect 1857 411 1923 445
rect 1857 377 1873 411
rect 1907 377 1923 411
rect 1857 343 1923 377
rect 2127 487 2161 527
rect 1959 419 1993 453
rect 1959 369 1993 385
rect 2027 445 2043 479
rect 2077 445 2093 479
rect 2027 411 2093 445
rect 2027 377 2043 411
rect 2077 377 2093 411
rect 1163 169 1289 203
rect 1129 153 1289 169
rect 564 55 586 89
rect 620 55 719 89
rect 753 89 793 105
rect 787 55 793 89
rect 843 73 863 107
rect 897 73 913 107
rect 947 73 963 107
rect 997 73 1095 107
rect 1145 101 1219 117
rect 395 17 461 55
rect 753 17 793 55
rect 1145 67 1179 101
rect 1213 67 1219 101
rect 1255 107 1289 153
rect 1323 191 1433 207
rect 1323 187 1369 191
rect 1323 153 1325 187
rect 1359 157 1369 187
rect 1403 157 1433 191
rect 1359 153 1433 157
rect 1323 141 1433 153
rect 1467 265 1527 281
rect 1714 265 1751 315
rect 1857 309 1873 343
rect 1907 335 1923 343
rect 2027 343 2093 377
rect 2127 419 2161 453
rect 2127 369 2161 385
rect 2027 335 2043 343
rect 1907 309 2043 335
rect 2077 335 2093 343
rect 2077 309 2191 335
rect 1857 301 2191 309
rect 1467 249 1680 265
rect 1467 215 1646 249
rect 1467 199 1680 215
rect 1714 249 2097 265
rect 1714 215 1843 249
rect 1877 215 1911 249
rect 1945 215 1979 249
rect 2013 215 2047 249
rect 2081 215 2097 249
rect 1467 107 1501 199
rect 1714 165 1750 215
rect 2131 181 2191 301
rect 1678 162 1750 165
rect 1678 128 1694 162
rect 1728 128 1750 162
rect 1857 164 2191 181
rect 1255 73 1297 107
rect 1331 73 1347 107
rect 1393 73 1409 107
rect 1443 73 1501 107
rect 1550 107 1624 123
rect 1550 73 1590 107
rect 1145 17 1219 67
rect 1550 17 1624 73
rect 1678 94 1750 128
rect 1678 60 1694 94
rect 1728 60 1750 94
rect 1785 123 1819 139
rect 1785 17 1819 89
rect 1857 130 1873 164
rect 1907 147 2043 164
rect 1907 130 1923 147
rect 1857 96 1923 130
rect 2027 130 2043 147
rect 2077 147 2191 164
rect 2077 130 2093 147
rect 1857 62 1873 96
rect 1907 62 1923 96
rect 1857 61 1923 62
rect 1959 96 1993 113
rect 1959 17 1993 62
rect 2027 96 2093 130
rect 2027 62 2043 96
rect 2077 62 2093 96
rect 2027 61 2093 62
rect 2127 96 2161 113
rect 2127 17 2161 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 123 357 157 391
rect 211 153 245 187
rect 1043 365 1077 391
rect 1043 357 1047 365
rect 1047 357 1077 365
rect 951 153 985 187
rect 1325 357 1359 391
rect 1325 153 1359 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
<< metal1 >>
rect 0 561 2208 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2208 561
rect 0 496 2208 527
rect 111 391 169 397
rect 111 357 123 391
rect 157 388 169 391
rect 1031 391 1089 397
rect 1031 388 1043 391
rect 157 360 1043 388
rect 157 357 169 360
rect 111 351 169 357
rect 1031 357 1043 360
rect 1077 388 1089 391
rect 1313 391 1371 397
rect 1313 388 1325 391
rect 1077 360 1325 388
rect 1077 357 1089 360
rect 1031 351 1089 357
rect 1313 357 1325 360
rect 1359 357 1371 391
rect 1313 351 1371 357
rect 199 187 257 193
rect 199 153 211 187
rect 245 184 257 187
rect 939 187 997 193
rect 939 184 951 187
rect 245 156 951 184
rect 245 153 257 156
rect 199 147 257 153
rect 939 153 951 156
rect 985 184 997 187
rect 1313 187 1371 193
rect 1313 184 1325 187
rect 985 156 1325 184
rect 985 153 997 156
rect 939 147 997 153
rect 1313 153 1325 156
rect 1359 153 1371 187
rect 1313 147 1371 153
rect 0 17 2208 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2208 17
rect 0 -48 2208 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 765 221 799 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel locali s 510 289 544 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 495 85 529 119 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 2145 221 2179 255 0 FreeSans 300 0 0 0 Q
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 sdfxtp_4
rlabel metal1 s 0 -48 2208 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2208 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2208 544
string GDS_END 408676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 392218
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.040 0.000 
<< end >>
