magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 349 0 352 90
<< via1 >>
rect 3 0 349 90
<< metal2 >>
rect 0 0 3 90
rect 349 0 352 90
<< properties >>
string GDS_END 85880402
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85878158
<< end >>
