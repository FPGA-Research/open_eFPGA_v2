magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1163 203
rect 30 -17 64 21
<< locali >>
rect 103 333 169 493
rect 375 333 441 425
rect 103 301 441 333
rect 122 289 441 301
rect 21 215 88 255
rect 122 177 169 289
rect 300 215 465 255
rect 519 215 716 255
rect 756 215 908 255
rect 944 215 1179 255
rect 103 127 169 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 299 69 527
rect 203 367 253 527
rect 291 459 509 493
rect 291 367 341 459
rect 475 323 509 459
rect 543 459 889 493
rect 543 367 609 459
rect 643 323 693 425
rect 475 289 693 323
rect 739 323 789 425
rect 823 367 889 459
rect 923 323 957 493
rect 991 357 1057 527
rect 1091 323 1141 493
rect 739 289 1141 323
rect 17 93 69 181
rect 203 147 1141 181
rect 203 93 253 147
rect 17 51 253 93
rect 291 17 341 109
rect 375 51 441 147
rect 475 17 509 109
rect 543 51 609 147
rect 643 17 690 109
rect 739 51 805 147
rect 839 17 873 109
rect 907 51 973 147
rect 1007 17 1041 109
rect 1075 51 1141 147
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 944 215 1179 255 6 A1
port 1 nsew signal input
rlabel locali s 756 215 908 255 6 A2
port 2 nsew signal input
rlabel locali s 519 215 716 255 6 A3
port 3 nsew signal input
rlabel locali s 300 215 465 255 6 A4
port 4 nsew signal input
rlabel locali s 21 215 88 255 6 B1
port 5 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1163 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 127 169 177 6 Y
port 10 nsew signal output
rlabel locali s 122 177 169 289 6 Y
port 10 nsew signal output
rlabel locali s 122 289 441 301 6 Y
port 10 nsew signal output
rlabel locali s 103 301 441 333 6 Y
port 10 nsew signal output
rlabel locali s 375 333 441 425 6 Y
port 10 nsew signal output
rlabel locali s 103 333 169 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 730510
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 719466
<< end >>
