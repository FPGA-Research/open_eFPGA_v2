magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 6060 4720 15316 4838
rect 3769 4650 15316 4720
rect 0 3991 15316 4650
rect 0 2500 15320 3991
rect 0 769 15000 2500
rect 0 766 12808 769
rect 0 90 8354 766
rect 11143 90 12808 766
<< nwell >>
rect -185 4561 15401 4921
rect -185 3937 11916 4561
rect -185 3907 10300 3937
rect -185 2240 290 3907
rect 897 3621 10300 3907
rect 3099 3589 10300 3621
rect 15114 2706 15401 4561
rect 14720 2420 15401 2706
rect -185 2024 1330 2240
rect 3110 2066 4530 2248
rect -185 970 660 2024
rect 8787 1705 9287 2020
rect 10118 1713 10556 2335
rect 10055 1705 10556 1713
rect 14720 1705 15084 2420
rect 8787 970 9089 1705
rect 11614 970 15084 1705
rect -185 823 15084 970
rect -185 370 11614 823
rect 14720 370 15084 823
rect -185 10 15084 370
<< pwell >>
rect 382 2308 1012 3144
rect 9145 2873 9307 3525
rect 8437 1038 8727 1980
<< mvpsubdiff >>
rect 9171 3475 9281 3499
rect 9171 3441 9175 3475
rect 9209 3441 9243 3475
rect 9277 3441 9281 3475
rect 9171 3401 9281 3441
rect 9171 3367 9175 3401
rect 9209 3367 9243 3401
rect 9277 3367 9281 3401
rect 9171 3327 9281 3367
rect 9171 3293 9175 3327
rect 9209 3293 9243 3327
rect 9277 3293 9281 3327
rect 9171 3253 9281 3293
rect 9171 3219 9175 3253
rect 9209 3219 9243 3253
rect 9277 3219 9281 3253
rect 9171 3179 9281 3219
rect 9171 3145 9175 3179
rect 9209 3145 9243 3179
rect 9277 3145 9281 3179
rect 408 3094 986 3118
rect 442 3060 476 3094
rect 510 3060 544 3094
rect 578 3060 612 3094
rect 646 3060 680 3094
rect 714 3060 748 3094
rect 782 3060 816 3094
rect 850 3060 884 3094
rect 918 3060 952 3094
rect 408 3023 986 3060
rect 442 2989 476 3023
rect 510 2989 544 3023
rect 578 2989 612 3023
rect 646 2989 680 3023
rect 714 2989 748 3023
rect 782 2989 816 3023
rect 850 2989 884 3023
rect 918 2989 952 3023
rect 408 2952 986 2989
rect 442 2918 476 2952
rect 510 2918 544 2952
rect 578 2918 612 2952
rect 646 2918 680 2952
rect 714 2918 748 2952
rect 782 2918 816 2952
rect 850 2918 884 2952
rect 918 2918 952 2952
rect 408 2882 986 2918
rect 9171 3105 9281 3145
rect 9171 3071 9175 3105
rect 9209 3071 9243 3105
rect 9277 3071 9281 3105
rect 9171 3031 9281 3071
rect 9171 2997 9175 3031
rect 9209 2997 9243 3031
rect 9277 2997 9281 3031
rect 9171 2957 9281 2997
rect 9171 2923 9175 2957
rect 9209 2923 9243 2957
rect 9277 2923 9281 2957
rect 9171 2899 9281 2923
rect 442 2848 476 2882
rect 510 2848 544 2882
rect 578 2848 612 2882
rect 646 2848 680 2882
rect 714 2848 748 2882
rect 782 2848 816 2882
rect 850 2848 884 2882
rect 918 2848 952 2882
rect 408 2812 986 2848
rect 442 2778 476 2812
rect 510 2778 544 2812
rect 578 2778 612 2812
rect 646 2778 680 2812
rect 714 2778 748 2812
rect 782 2778 816 2812
rect 850 2778 884 2812
rect 918 2778 952 2812
rect 408 2742 986 2778
rect 442 2708 476 2742
rect 510 2708 544 2742
rect 578 2708 612 2742
rect 646 2708 680 2742
rect 714 2708 748 2742
rect 782 2708 816 2742
rect 850 2708 884 2742
rect 918 2708 952 2742
rect 408 2672 986 2708
rect 442 2638 476 2672
rect 510 2638 544 2672
rect 578 2638 612 2672
rect 646 2638 680 2672
rect 714 2638 748 2672
rect 782 2638 816 2672
rect 850 2638 884 2672
rect 918 2638 952 2672
rect 408 2602 986 2638
rect 442 2568 476 2602
rect 510 2568 544 2602
rect 578 2568 612 2602
rect 646 2568 680 2602
rect 714 2568 748 2602
rect 782 2568 816 2602
rect 850 2568 884 2602
rect 918 2568 952 2602
rect 408 2532 986 2568
rect 442 2498 476 2532
rect 510 2498 544 2532
rect 578 2498 612 2532
rect 646 2498 680 2532
rect 714 2498 748 2532
rect 782 2498 816 2532
rect 850 2498 884 2532
rect 918 2498 952 2532
rect 408 2462 986 2498
rect 442 2428 476 2462
rect 510 2428 544 2462
rect 578 2428 612 2462
rect 646 2428 680 2462
rect 714 2428 748 2462
rect 782 2428 816 2462
rect 850 2428 884 2462
rect 918 2428 952 2462
rect 408 2392 986 2428
rect 442 2358 476 2392
rect 510 2358 544 2392
rect 578 2358 612 2392
rect 646 2358 680 2392
rect 714 2358 748 2392
rect 782 2358 816 2392
rect 850 2358 884 2392
rect 918 2358 952 2392
rect 408 2334 986 2358
rect 8463 1930 8701 1954
rect 8497 1896 8531 1930
rect 8565 1896 8599 1930
rect 8633 1896 8667 1930
rect 8463 1856 8701 1896
rect 8497 1822 8531 1856
rect 8565 1822 8599 1856
rect 8633 1822 8667 1856
rect 8463 1782 8701 1822
rect 8497 1748 8531 1782
rect 8565 1748 8599 1782
rect 8633 1748 8667 1782
rect 8463 1708 8701 1748
rect 8497 1674 8531 1708
rect 8565 1674 8599 1708
rect 8633 1674 8667 1708
rect 8463 1634 8701 1674
rect 8497 1600 8531 1634
rect 8565 1600 8599 1634
rect 8633 1600 8667 1634
rect 8463 1560 8701 1600
rect 8497 1526 8531 1560
rect 8565 1526 8599 1560
rect 8633 1526 8667 1560
rect 8463 1487 8701 1526
rect 8497 1453 8531 1487
rect 8565 1453 8599 1487
rect 8633 1453 8667 1487
rect 8463 1414 8701 1453
rect 8497 1380 8531 1414
rect 8565 1380 8599 1414
rect 8633 1380 8667 1414
rect 8463 1341 8701 1380
rect 8497 1307 8531 1341
rect 8565 1307 8599 1341
rect 8633 1307 8667 1341
rect 8463 1268 8701 1307
rect 8497 1234 8531 1268
rect 8565 1234 8599 1268
rect 8633 1234 8667 1268
rect 8463 1195 8701 1234
rect 8497 1161 8531 1195
rect 8565 1161 8599 1195
rect 8633 1161 8667 1195
rect 8463 1122 8701 1161
rect 8497 1088 8531 1122
rect 8565 1088 8599 1122
rect 8633 1088 8667 1122
rect 8463 1064 8701 1088
<< mvnsubdiff >>
rect -17 4821 43 4855
rect 77 4821 151 4855
rect 185 4821 220 4855
rect 254 4821 289 4855
rect 323 4821 358 4855
rect 392 4821 427 4855
rect 461 4821 496 4855
rect 530 4821 565 4855
rect 599 4821 634 4855
rect 668 4821 703 4855
rect 737 4821 772 4855
rect 806 4821 841 4855
rect 875 4821 910 4855
rect 944 4821 979 4855
rect 1013 4821 1048 4855
rect 1082 4821 1117 4855
rect 1151 4821 1186 4855
rect 1220 4821 1255 4855
rect 1289 4821 1324 4855
rect 1358 4821 1393 4855
rect 1427 4821 1462 4855
rect 1496 4821 1531 4855
rect 1565 4821 1600 4855
rect 1634 4821 1669 4855
rect 1703 4821 1738 4855
rect 1772 4821 1807 4855
rect 1841 4821 1875 4855
rect 1909 4821 1943 4855
rect 1977 4821 2011 4855
rect 2045 4821 2079 4855
rect 2113 4821 2147 4855
rect 2181 4821 2215 4855
rect 2249 4821 2283 4855
rect 2317 4821 2351 4855
rect 2385 4821 2419 4855
rect 2453 4821 2487 4855
rect 2521 4821 2555 4855
rect 3971 4821 3983 4855
rect 4017 4821 4051 4855
rect 4085 4821 4119 4855
rect 4153 4821 4187 4855
rect 4221 4821 4255 4855
rect 4289 4821 4323 4855
rect 4357 4821 4391 4855
rect 4425 4821 4459 4855
rect 4493 4821 4527 4855
rect 4561 4821 4595 4855
rect 4629 4821 4663 4855
rect 4697 4821 4731 4855
rect 4765 4821 4799 4855
rect 4833 4821 4867 4855
rect 4901 4821 4935 4855
rect 4969 4821 5003 4855
rect 5037 4821 5071 4855
rect 5105 4821 5139 4855
rect 5173 4821 5207 4855
rect 5241 4821 5275 4855
rect 5309 4821 5343 4855
rect 5377 4821 5411 4855
rect 5445 4821 5479 4855
rect 5513 4821 5547 4855
rect 5581 4821 5615 4855
rect 5649 4821 5683 4855
rect 5717 4821 5751 4855
rect 5785 4821 5819 4855
rect 5853 4821 5887 4855
rect 5921 4821 5955 4855
rect 5989 4821 6023 4855
rect 6057 4821 6091 4855
rect 6125 4821 6159 4855
rect 6193 4821 6227 4855
rect 6261 4821 6295 4855
rect 6329 4821 6363 4855
rect 6397 4821 6431 4855
rect 6465 4821 6499 4855
rect 6533 4821 6567 4855
rect 6601 4821 6635 4855
rect 6669 4821 6703 4855
rect 6737 4821 6771 4855
rect 6805 4821 6839 4855
rect 6873 4821 6907 4855
rect 6941 4821 6975 4855
rect 7009 4821 7043 4855
rect 7077 4821 7111 4855
rect 7145 4821 7179 4855
rect 7213 4821 7247 4855
rect 7281 4821 7315 4855
rect 7349 4821 7383 4855
rect 7417 4821 7451 4855
rect 7485 4821 7519 4855
rect 7553 4821 7587 4855
rect 7621 4821 7655 4855
rect 7689 4821 7723 4855
rect 7757 4821 7791 4855
rect 7825 4821 7859 4855
rect 7893 4821 7927 4855
rect 7961 4821 7995 4855
rect 8029 4821 8063 4855
rect 8097 4821 8131 4855
rect 8165 4821 8199 4855
rect 8233 4821 8267 4855
rect 8301 4821 8335 4855
rect 8369 4821 8403 4855
rect 8437 4821 8471 4855
rect 8505 4821 8539 4855
rect 8573 4821 8607 4855
rect 8641 4821 8675 4855
rect 8709 4821 8743 4855
rect 8777 4821 8811 4855
rect 8845 4821 8879 4855
rect 8913 4821 8947 4855
rect 8981 4821 9015 4855
rect 9049 4821 9083 4855
rect 9117 4821 9151 4855
rect 9185 4821 9219 4855
rect 9253 4821 9287 4855
rect 9321 4821 9355 4855
rect 9389 4821 9423 4855
rect 9457 4821 9491 4855
rect 9525 4821 9559 4855
rect 9593 4821 9627 4855
rect 9661 4821 9695 4855
rect 9729 4821 9763 4855
rect 9797 4821 9831 4855
rect 9865 4821 9899 4855
rect 9933 4821 9967 4855
rect 10001 4821 10035 4855
rect 10069 4821 10103 4855
rect 10137 4821 10171 4855
rect 10205 4821 10239 4855
rect 10273 4821 10307 4855
rect 10341 4821 10375 4855
rect 10409 4821 10443 4855
rect 10477 4821 10511 4855
rect 10545 4821 10579 4855
rect 10613 4821 10647 4855
rect 10681 4821 10715 4855
rect 10749 4821 10783 4855
rect 10817 4821 10851 4855
rect 10885 4821 10919 4855
rect 10953 4821 10987 4855
rect 11021 4821 11055 4855
rect 11089 4821 11123 4855
rect 11157 4821 11191 4855
rect 11225 4821 11259 4855
rect 11293 4821 11327 4855
rect 11361 4821 11395 4855
rect 11429 4821 11463 4855
rect 11497 4821 11531 4855
rect 11565 4821 11599 4855
rect 11633 4821 11667 4855
rect 11701 4821 11735 4855
rect 11769 4821 11803 4855
rect 11837 4821 11871 4855
rect 11905 4821 11939 4855
rect 11973 4821 12007 4855
rect 12041 4821 12075 4855
rect 12109 4821 12143 4855
rect 12177 4821 12201 4855
rect -17 4787 2577 4821
rect -17 4753 93 4787
rect 127 4753 162 4787
rect 196 4753 231 4787
rect 265 4753 300 4787
rect 334 4753 369 4787
rect 403 4753 438 4787
rect 472 4753 507 4787
rect 541 4753 576 4787
rect 610 4753 645 4787
rect 679 4753 714 4787
rect 748 4753 783 4787
rect 817 4753 852 4787
rect 886 4753 921 4787
rect 955 4753 990 4787
rect 1024 4753 1059 4787
rect 1093 4753 1128 4787
rect 1162 4753 1197 4787
rect 1231 4753 1266 4787
rect 1300 4753 1335 4787
rect 1369 4753 1404 4787
rect 1438 4753 1473 4787
rect 1507 4753 1542 4787
rect 1576 4753 1611 4787
rect 1645 4753 1680 4787
rect 1714 4753 1749 4787
rect 1783 4753 1818 4787
rect 1852 4753 1887 4787
rect 1921 4753 1956 4787
rect 1990 4753 2025 4787
rect 2059 4753 2094 4787
rect 2128 4753 2163 4787
rect 2197 4753 2232 4787
rect 2266 4753 2301 4787
rect 2335 4753 2370 4787
rect 2404 4753 2439 4787
rect 2473 4753 2508 4787
rect 2542 4753 2577 4787
rect 17 4719 2577 4753
rect -17 4685 93 4719
rect 127 4685 162 4719
rect 196 4685 231 4719
rect 265 4685 300 4719
rect 334 4685 369 4719
rect 403 4685 438 4719
rect 472 4685 507 4719
rect 541 4685 576 4719
rect 610 4685 645 4719
rect 679 4685 714 4719
rect 748 4685 783 4719
rect 817 4685 852 4719
rect 886 4685 921 4719
rect 955 4685 990 4719
rect 1024 4685 1059 4719
rect 1093 4685 1128 4719
rect 1162 4685 1197 4719
rect 1231 4685 1266 4719
rect 1300 4685 1335 4719
rect 1369 4685 1404 4719
rect 1438 4685 1473 4719
rect 1507 4685 1542 4719
rect 1576 4685 1611 4719
rect 1645 4685 1680 4719
rect 1714 4685 1749 4719
rect 1783 4685 1818 4719
rect 1852 4685 1887 4719
rect 1921 4685 1956 4719
rect 1990 4685 2025 4719
rect 2059 4685 2094 4719
rect 2128 4685 2163 4719
rect 2197 4685 2232 4719
rect 2266 4685 2301 4719
rect 2335 4685 2370 4719
rect 2404 4685 2439 4719
rect 2473 4685 2508 4719
rect 2542 4685 2577 4719
rect 17 4651 2577 4685
rect -17 4617 93 4651
rect 127 4617 162 4651
rect 196 4617 231 4651
rect 265 4617 300 4651
rect 334 4617 369 4651
rect 403 4617 438 4651
rect 472 4617 507 4651
rect 541 4617 576 4651
rect 610 4617 645 4651
rect 679 4617 714 4651
rect 748 4617 783 4651
rect 817 4617 852 4651
rect 886 4617 921 4651
rect 955 4617 990 4651
rect 1024 4617 1059 4651
rect 1093 4617 1128 4651
rect 1162 4617 1197 4651
rect 1231 4617 1266 4651
rect 1300 4617 1335 4651
rect 1369 4617 1404 4651
rect 1438 4617 1473 4651
rect 1507 4617 1542 4651
rect 1576 4617 1611 4651
rect 1645 4617 1680 4651
rect 1714 4617 1749 4651
rect 1783 4617 1818 4651
rect 1852 4617 1887 4651
rect 1921 4617 1956 4651
rect 1990 4617 2025 4651
rect 2059 4617 2094 4651
rect 2128 4617 2163 4651
rect 2197 4617 2232 4651
rect 2266 4617 2301 4651
rect 2335 4617 2370 4651
rect 2404 4617 2439 4651
rect 2473 4617 2508 4651
rect 2542 4617 2577 4651
rect 3971 4752 4674 4821
rect 3971 4718 4056 4752
rect 4090 4718 4126 4752
rect 4160 4718 4196 4752
rect 4230 4718 4266 4752
rect 4300 4718 4336 4752
rect 4370 4718 4406 4752
rect 4440 4718 4476 4752
rect 4510 4718 4546 4752
rect 4580 4718 4616 4752
rect 4650 4718 4674 4752
rect 3971 4695 4674 4718
rect 3971 4617 3995 4695
rect 4636 4663 4674 4695
rect 7833 4752 8428 4821
rect 7833 4718 7857 4752
rect 7891 4718 7931 4752
rect 7965 4718 8005 4752
rect 8039 4718 8078 4752
rect 8112 4718 8151 4752
rect 8185 4718 8224 4752
rect 8258 4718 8297 4752
rect 8331 4718 8370 4752
rect 8404 4718 8428 4752
rect 7833 4663 8428 4718
rect 17 4583 3995 4617
rect -17 4581 3995 4583
rect -17 4549 93 4581
rect 17 4547 93 4549
rect 127 4547 167 4581
rect 201 4547 241 4581
rect 275 4547 315 4581
rect 349 4547 388 4581
rect 422 4547 461 4581
rect 495 4547 534 4581
rect 568 4547 607 4581
rect 641 4547 680 4581
rect 714 4547 753 4581
rect 787 4571 3995 4581
rect 7833 4629 7857 4663
rect 7891 4629 7931 4663
rect 7965 4629 8005 4663
rect 8039 4629 8078 4663
rect 8112 4629 8151 4663
rect 8185 4629 8224 4663
rect 8258 4629 8297 4663
rect 8331 4629 8370 4663
rect 8404 4629 8428 4663
rect 7833 4595 8428 4629
rect 787 4547 811 4571
rect 17 4515 811 4547
rect -17 4513 811 4515
rect -17 4481 93 4513
rect 17 4479 93 4481
rect 127 4479 167 4513
rect 201 4479 241 4513
rect 275 4479 315 4513
rect 349 4479 388 4513
rect 422 4479 461 4513
rect 495 4479 534 4513
rect 568 4479 607 4513
rect 641 4479 680 4513
rect 714 4479 753 4513
rect 787 4479 811 4513
rect 17 4447 811 4479
rect -17 4445 811 4447
rect -17 4413 93 4445
rect 17 4411 93 4413
rect 127 4411 167 4445
rect 201 4411 241 4445
rect 275 4411 315 4445
rect 349 4411 388 4445
rect 422 4411 461 4445
rect 495 4411 534 4445
rect 568 4411 607 4445
rect 641 4411 680 4445
rect 714 4411 753 4445
rect 787 4411 811 4445
rect 7833 4561 7857 4595
rect 7891 4561 7931 4595
rect 7965 4561 8005 4595
rect 8039 4561 8078 4595
rect 8112 4561 8151 4595
rect 8185 4561 8224 4595
rect 8258 4561 8297 4595
rect 8331 4561 8370 4595
rect 8404 4561 8428 4595
rect 7833 4527 8428 4561
rect 7833 4493 7857 4527
rect 7891 4493 7931 4527
rect 7965 4493 8005 4527
rect 8039 4493 8078 4527
rect 8112 4493 8151 4527
rect 8185 4493 8224 4527
rect 8258 4493 8297 4527
rect 8331 4493 8370 4527
rect 8404 4493 8428 4527
rect 7833 4459 8428 4493
rect 7833 4425 7857 4459
rect 7891 4425 7931 4459
rect 7965 4425 8005 4459
rect 8039 4425 8078 4459
rect 8112 4425 8151 4459
rect 8185 4425 8224 4459
rect 8258 4425 8297 4459
rect 8331 4425 8370 4459
rect 8404 4425 8428 4459
rect 17 4379 197 4411
rect 7833 4392 8428 4425
rect -17 4377 197 4379
rect -17 4345 140 4377
rect 17 4343 140 4345
rect 174 4343 197 4377
rect 17 4311 197 4343
rect -17 4309 197 4311
rect -17 4277 140 4309
rect 17 4275 140 4277
rect 174 4275 197 4309
rect 17 4243 197 4275
rect -17 4241 197 4243
rect -17 4209 140 4241
rect 17 4207 140 4209
rect 174 4207 197 4241
rect 17 4175 197 4207
rect -17 4173 197 4175
rect -17 4141 140 4173
rect 17 4139 140 4141
rect 174 4139 197 4173
rect 17 4107 197 4139
rect -17 4105 197 4107
rect -17 4073 140 4105
rect 17 4071 140 4073
rect 174 4071 197 4105
rect 17 4039 197 4071
rect -17 4037 197 4039
rect -17 4005 140 4037
rect 17 4003 140 4005
rect 174 4003 197 4037
rect 17 3971 197 4003
rect -17 3969 197 3971
rect -17 3937 140 3969
rect 17 3935 140 3937
rect 174 3935 197 3969
rect 17 3903 197 3935
rect -17 3901 197 3903
rect -17 3869 140 3901
rect 17 3867 140 3869
rect 174 3867 197 3901
rect 17 3835 197 3867
rect -17 3833 197 3835
rect -17 3801 140 3833
rect 17 3799 140 3801
rect 174 3799 197 3833
rect 17 3767 197 3799
rect -17 3765 197 3767
rect -17 3733 140 3765
rect 17 3731 140 3733
rect 174 3731 197 3765
rect 17 3699 197 3731
rect -17 3697 197 3699
rect -17 3665 140 3697
rect 17 3663 140 3665
rect 174 3663 197 3697
rect 17 3631 197 3663
rect -17 3629 197 3631
rect -17 3597 140 3629
rect 17 3595 140 3597
rect 174 3595 197 3629
rect 17 3563 197 3595
rect -17 3561 197 3563
rect -17 3529 140 3561
rect 17 3527 140 3529
rect 174 3527 197 3561
rect 17 3495 197 3527
rect -17 3493 197 3495
rect -17 3461 140 3493
rect 17 3459 140 3461
rect 174 3459 197 3493
rect 17 3427 197 3459
rect -17 3425 197 3427
rect -17 3393 140 3425
rect 17 3391 140 3393
rect 174 3391 197 3425
rect 17 3359 197 3391
rect -17 3357 197 3359
rect -17 3325 140 3357
rect 17 3323 140 3325
rect 174 3323 197 3357
rect 17 3291 197 3323
rect -17 3289 197 3291
rect -17 3257 140 3289
rect 17 3255 140 3257
rect 174 3255 197 3289
rect 17 3223 197 3255
rect -17 3221 197 3223
rect -17 3189 140 3221
rect 17 3187 140 3189
rect 174 3187 197 3221
rect 17 3155 197 3187
rect -17 3152 197 3155
rect -17 3121 140 3152
rect 17 3118 140 3121
rect 174 3118 197 3152
rect 17 3087 197 3118
rect -17 3083 197 3087
rect -17 3053 140 3083
rect 17 3049 140 3053
rect 174 3049 197 3083
rect 17 3019 197 3049
rect -17 3014 197 3019
rect -17 2985 140 3014
rect 17 2980 140 2985
rect 174 2980 197 3014
rect 17 2951 197 2980
rect -17 2945 197 2951
rect -17 2917 140 2945
rect 17 2911 140 2917
rect 174 2911 197 2945
rect 17 2883 197 2911
rect -17 2876 197 2883
rect -17 2849 140 2876
rect 17 2842 140 2849
rect 174 2842 197 2876
rect 17 2815 197 2842
rect -17 2807 197 2815
rect -17 2781 140 2807
rect 17 2773 140 2781
rect 174 2773 197 2807
rect 17 2747 197 2773
rect -17 2738 197 2747
rect -17 2713 140 2738
rect 17 2704 140 2713
rect 174 2704 197 2738
rect 17 2679 197 2704
rect -17 2669 197 2679
rect -17 2645 140 2669
rect 17 2635 140 2645
rect 174 2635 197 2669
rect 17 2611 197 2635
rect -17 2600 197 2611
rect -17 2577 140 2600
rect 17 2566 140 2577
rect 174 2566 197 2600
rect 17 2543 197 2566
rect -17 2531 197 2543
rect -17 2509 140 2531
rect 17 2497 140 2509
rect 174 2497 197 2531
rect 17 2475 197 2497
rect -17 2462 197 2475
rect -17 2441 140 2462
rect 17 2428 140 2441
rect 174 2428 197 2462
rect 17 2407 197 2428
rect -17 2393 197 2407
rect -17 2372 140 2393
rect 17 2359 140 2372
rect 174 2359 197 2393
rect 17 2338 197 2359
rect -17 2324 197 2338
rect 14983 2486 15038 2520
rect 14983 2418 15017 2452
rect 14983 2350 15017 2384
rect -17 2303 140 2324
rect 17 2290 140 2303
rect 174 2290 197 2324
rect 17 2269 197 2290
rect 14983 2282 15017 2316
rect -17 2255 197 2269
rect -17 2234 140 2255
rect 17 2221 140 2234
rect 174 2221 197 2255
rect 17 2200 197 2221
rect -17 2186 197 2200
rect -17 2165 140 2186
rect 17 2152 140 2165
rect 174 2152 197 2186
rect 10184 2245 10490 2269
rect 17 2131 197 2152
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect -17 2117 197 2131
rect -17 2096 140 2117
rect 17 2083 140 2096
rect 174 2083 197 2117
rect 17 2062 197 2083
rect -17 2048 197 2062
rect -17 2027 140 2048
rect 17 2014 140 2027
rect 174 2014 197 2048
rect 17 2004 197 2014
rect 17 1993 587 2004
rect -17 1980 587 1993
rect -17 1958 145 1980
rect 17 1946 145 1958
rect 179 1946 213 1980
rect 247 1946 281 1980
rect 315 1946 349 1980
rect 383 1946 417 1980
rect 451 1946 485 1980
rect 519 1946 553 1980
rect 17 1924 587 1946
rect -17 1909 587 1924
rect -17 1889 145 1909
rect 17 1875 145 1889
rect 179 1875 213 1909
rect 247 1875 281 1909
rect 315 1875 349 1909
rect 383 1875 417 1909
rect 451 1875 485 1909
rect 519 1875 553 1909
rect 17 1855 587 1875
rect -17 1838 587 1855
rect -17 1820 145 1838
rect 17 1804 145 1820
rect 179 1804 213 1838
rect 247 1804 281 1838
rect 315 1804 349 1838
rect 383 1804 417 1838
rect 451 1804 485 1838
rect 519 1804 553 1838
rect 17 1786 587 1804
rect -17 1767 587 1786
rect -17 1751 145 1767
rect 17 1733 145 1751
rect 179 1733 213 1767
rect 247 1733 281 1767
rect 315 1733 349 1767
rect 383 1733 417 1767
rect 451 1733 485 1767
rect 519 1733 553 1767
rect 17 1717 587 1733
rect -17 1696 587 1717
rect -17 1682 145 1696
rect 17 1662 145 1682
rect 179 1662 213 1696
rect 247 1662 281 1696
rect 315 1662 349 1696
rect 383 1662 417 1696
rect 451 1662 485 1696
rect 519 1662 553 1696
rect 17 1648 587 1662
rect -17 1625 587 1648
rect -17 1613 145 1625
rect 17 1591 145 1613
rect 179 1591 213 1625
rect 247 1591 281 1625
rect 315 1591 349 1625
rect 383 1591 417 1625
rect 451 1591 485 1625
rect 519 1591 553 1625
rect 17 1579 587 1591
rect -17 1554 587 1579
rect -17 1544 145 1554
rect 17 1520 145 1544
rect 179 1520 213 1554
rect 247 1520 281 1554
rect 315 1520 349 1554
rect 383 1520 417 1554
rect 451 1520 485 1554
rect 519 1520 553 1554
rect 17 1510 587 1520
rect -17 1483 587 1510
rect -17 1475 145 1483
rect 17 1449 145 1475
rect 179 1449 213 1483
rect 247 1449 281 1483
rect 315 1449 349 1483
rect 383 1449 417 1483
rect 451 1449 485 1483
rect 519 1449 553 1483
rect 17 1441 587 1449
rect -17 1412 587 1441
rect -17 1406 145 1412
rect 17 1378 145 1406
rect 179 1378 213 1412
rect 247 1378 281 1412
rect 315 1378 349 1412
rect 383 1378 417 1412
rect 451 1378 485 1412
rect 519 1378 553 1412
rect 17 1372 587 1378
rect -17 1342 587 1372
rect -17 1337 145 1342
rect 17 1308 145 1337
rect 179 1308 213 1342
rect 247 1308 281 1342
rect 315 1308 349 1342
rect 383 1308 417 1342
rect 451 1308 485 1342
rect 519 1308 553 1342
rect 17 1303 587 1308
rect -17 1272 587 1303
rect -17 1268 145 1272
rect 17 1238 145 1268
rect 179 1238 213 1272
rect 247 1238 281 1272
rect 315 1238 349 1272
rect 383 1238 417 1272
rect 451 1238 485 1272
rect 519 1238 553 1272
rect 17 1234 587 1238
rect -17 1202 587 1234
rect -17 1199 145 1202
rect 17 1168 145 1199
rect 179 1168 213 1202
rect 247 1168 281 1202
rect 315 1168 349 1202
rect 383 1168 417 1202
rect 451 1168 485 1202
rect 519 1168 553 1202
rect 17 1165 587 1168
rect -17 1132 587 1165
rect -17 1130 145 1132
rect 17 1098 145 1130
rect 179 1098 213 1132
rect 247 1098 281 1132
rect 315 1098 349 1132
rect 383 1098 417 1132
rect 451 1098 485 1132
rect 519 1098 553 1132
rect 17 1096 587 1098
rect -17 1062 587 1096
rect 8853 1930 9023 1954
rect 8887 1896 8921 1930
rect 8955 1896 8989 1930
rect 8853 1860 9023 1896
rect 8887 1826 8921 1860
rect 8955 1826 8989 1860
rect 8853 1790 9023 1826
rect 8887 1756 8921 1790
rect 8955 1756 8989 1790
rect 9155 1930 9221 1954
rect 9155 1896 9171 1930
rect 9205 1896 9221 1930
rect 9155 1829 9221 1896
rect 9155 1795 9171 1829
rect 9205 1795 9221 1829
rect 9155 1771 9221 1795
rect 10184 1779 10490 1803
rect 14983 2214 15017 2248
rect 14983 2146 15017 2180
rect 14983 2078 15017 2112
rect 14983 2010 15017 2044
rect 14983 1942 15017 1976
rect 14983 1874 15017 1908
rect 14983 1806 15017 1840
rect 8853 1721 9023 1756
rect 8887 1687 8921 1721
rect 8955 1687 8989 1721
rect 8853 1652 9023 1687
rect 8887 1618 8921 1652
rect 8955 1618 8989 1652
rect 8853 1583 9023 1618
rect 8887 1549 8921 1583
rect 8955 1549 8989 1583
rect 8853 1514 9023 1549
rect 8887 1480 8921 1514
rect 8955 1480 8989 1514
rect 8853 1445 9023 1480
rect 8887 1411 8921 1445
rect 8955 1411 8989 1445
rect 8853 1376 9023 1411
rect 8887 1342 8921 1376
rect 8955 1342 8989 1376
rect 8853 1307 9023 1342
rect 8887 1273 8921 1307
rect 8955 1273 8989 1307
rect 8853 1238 9023 1273
rect 8887 1204 8921 1238
rect 8955 1204 8989 1238
rect 8853 1169 9023 1204
rect 8887 1135 8921 1169
rect 8955 1135 8989 1169
rect 8853 1100 9023 1135
rect 8887 1066 8921 1100
rect 8955 1066 8989 1100
rect -17 1061 145 1062
rect 17 1028 145 1061
rect 179 1028 213 1062
rect 247 1028 281 1062
rect 315 1028 349 1062
rect 383 1028 417 1062
rect 451 1028 485 1062
rect 519 1028 553 1062
rect 17 1027 587 1028
rect -17 1004 587 1027
rect 8853 1031 9023 1066
rect -17 992 17 1004
rect 8887 997 8921 1031
rect 8955 997 8989 1031
rect 8853 973 9023 997
rect 14983 1738 15017 1772
rect 14983 1670 15017 1704
rect 14983 1602 15017 1636
rect 14983 1534 15017 1568
rect 14983 1466 15017 1500
rect 14983 1398 15017 1432
rect 14983 1330 15017 1364
rect 14983 1262 15017 1296
rect 14983 1194 15017 1228
rect 14983 1126 15017 1160
rect 14983 1058 15017 1092
rect 14983 990 15017 1024
rect -17 923 17 958
rect -17 854 17 889
rect -17 785 17 820
rect 14983 922 15017 956
rect 14983 854 15017 888
rect 14983 786 15017 820
rect -17 727 17 751
rect 14893 752 14983 766
rect 14893 718 15017 752
rect 14893 684 14983 718
rect 14893 650 15017 684
rect 14893 616 14983 650
rect 14893 582 15017 616
rect 14893 548 14983 582
rect 14893 514 15017 548
rect 14893 480 14983 514
rect 14893 446 15017 480
rect 14893 412 14983 446
rect 14893 378 15017 412
rect 14893 344 14983 378
rect 14893 310 15017 344
rect 14893 276 14983 310
rect 14893 242 15017 276
rect 14893 208 14983 242
rect 14893 174 15017 208
rect 14893 140 14983 174
rect 14893 76 15017 140
<< mvpsubdiffcont >>
rect 9175 3441 9209 3475
rect 9243 3441 9277 3475
rect 9175 3367 9209 3401
rect 9243 3367 9277 3401
rect 9175 3293 9209 3327
rect 9243 3293 9277 3327
rect 9175 3219 9209 3253
rect 9243 3219 9277 3253
rect 9175 3145 9209 3179
rect 9243 3145 9277 3179
rect 408 3060 442 3094
rect 476 3060 510 3094
rect 544 3060 578 3094
rect 612 3060 646 3094
rect 680 3060 714 3094
rect 748 3060 782 3094
rect 816 3060 850 3094
rect 884 3060 918 3094
rect 952 3060 986 3094
rect 408 2989 442 3023
rect 476 2989 510 3023
rect 544 2989 578 3023
rect 612 2989 646 3023
rect 680 2989 714 3023
rect 748 2989 782 3023
rect 816 2989 850 3023
rect 884 2989 918 3023
rect 952 2989 986 3023
rect 408 2918 442 2952
rect 476 2918 510 2952
rect 544 2918 578 2952
rect 612 2918 646 2952
rect 680 2918 714 2952
rect 748 2918 782 2952
rect 816 2918 850 2952
rect 884 2918 918 2952
rect 952 2918 986 2952
rect 9175 3071 9209 3105
rect 9243 3071 9277 3105
rect 9175 2997 9209 3031
rect 9243 2997 9277 3031
rect 9175 2923 9209 2957
rect 9243 2923 9277 2957
rect 408 2848 442 2882
rect 476 2848 510 2882
rect 544 2848 578 2882
rect 612 2848 646 2882
rect 680 2848 714 2882
rect 748 2848 782 2882
rect 816 2848 850 2882
rect 884 2848 918 2882
rect 952 2848 986 2882
rect 408 2778 442 2812
rect 476 2778 510 2812
rect 544 2778 578 2812
rect 612 2778 646 2812
rect 680 2778 714 2812
rect 748 2778 782 2812
rect 816 2778 850 2812
rect 884 2778 918 2812
rect 952 2778 986 2812
rect 408 2708 442 2742
rect 476 2708 510 2742
rect 544 2708 578 2742
rect 612 2708 646 2742
rect 680 2708 714 2742
rect 748 2708 782 2742
rect 816 2708 850 2742
rect 884 2708 918 2742
rect 952 2708 986 2742
rect 408 2638 442 2672
rect 476 2638 510 2672
rect 544 2638 578 2672
rect 612 2638 646 2672
rect 680 2638 714 2672
rect 748 2638 782 2672
rect 816 2638 850 2672
rect 884 2638 918 2672
rect 952 2638 986 2672
rect 408 2568 442 2602
rect 476 2568 510 2602
rect 544 2568 578 2602
rect 612 2568 646 2602
rect 680 2568 714 2602
rect 748 2568 782 2602
rect 816 2568 850 2602
rect 884 2568 918 2602
rect 952 2568 986 2602
rect 408 2498 442 2532
rect 476 2498 510 2532
rect 544 2498 578 2532
rect 612 2498 646 2532
rect 680 2498 714 2532
rect 748 2498 782 2532
rect 816 2498 850 2532
rect 884 2498 918 2532
rect 952 2498 986 2532
rect 408 2428 442 2462
rect 476 2428 510 2462
rect 544 2428 578 2462
rect 612 2428 646 2462
rect 680 2428 714 2462
rect 748 2428 782 2462
rect 816 2428 850 2462
rect 884 2428 918 2462
rect 952 2428 986 2462
rect 408 2358 442 2392
rect 476 2358 510 2392
rect 544 2358 578 2392
rect 612 2358 646 2392
rect 680 2358 714 2392
rect 748 2358 782 2392
rect 816 2358 850 2392
rect 884 2358 918 2392
rect 952 2358 986 2392
rect 8463 1896 8497 1930
rect 8531 1896 8565 1930
rect 8599 1896 8633 1930
rect 8667 1896 8701 1930
rect 8463 1822 8497 1856
rect 8531 1822 8565 1856
rect 8599 1822 8633 1856
rect 8667 1822 8701 1856
rect 8463 1748 8497 1782
rect 8531 1748 8565 1782
rect 8599 1748 8633 1782
rect 8667 1748 8701 1782
rect 8463 1674 8497 1708
rect 8531 1674 8565 1708
rect 8599 1674 8633 1708
rect 8667 1674 8701 1708
rect 8463 1600 8497 1634
rect 8531 1600 8565 1634
rect 8599 1600 8633 1634
rect 8667 1600 8701 1634
rect 8463 1526 8497 1560
rect 8531 1526 8565 1560
rect 8599 1526 8633 1560
rect 8667 1526 8701 1560
rect 8463 1453 8497 1487
rect 8531 1453 8565 1487
rect 8599 1453 8633 1487
rect 8667 1453 8701 1487
rect 8463 1380 8497 1414
rect 8531 1380 8565 1414
rect 8599 1380 8633 1414
rect 8667 1380 8701 1414
rect 8463 1307 8497 1341
rect 8531 1307 8565 1341
rect 8599 1307 8633 1341
rect 8667 1307 8701 1341
rect 8463 1234 8497 1268
rect 8531 1234 8565 1268
rect 8599 1234 8633 1268
rect 8667 1234 8701 1268
rect 8463 1161 8497 1195
rect 8531 1161 8565 1195
rect 8599 1161 8633 1195
rect 8667 1161 8701 1195
rect 8463 1088 8497 1122
rect 8531 1088 8565 1122
rect 8599 1088 8633 1122
rect 8667 1088 8701 1122
<< mvnsubdiffcont >>
rect 43 4821 77 4855
rect 151 4821 185 4855
rect 220 4821 254 4855
rect 289 4821 323 4855
rect 358 4821 392 4855
rect 427 4821 461 4855
rect 496 4821 530 4855
rect 565 4821 599 4855
rect 634 4821 668 4855
rect 703 4821 737 4855
rect 772 4821 806 4855
rect 841 4821 875 4855
rect 910 4821 944 4855
rect 979 4821 1013 4855
rect 1048 4821 1082 4855
rect 1117 4821 1151 4855
rect 1186 4821 1220 4855
rect 1255 4821 1289 4855
rect 1324 4821 1358 4855
rect 1393 4821 1427 4855
rect 1462 4821 1496 4855
rect 1531 4821 1565 4855
rect 1600 4821 1634 4855
rect 1669 4821 1703 4855
rect 1738 4821 1772 4855
rect 1807 4821 1841 4855
rect 1875 4821 1909 4855
rect 1943 4821 1977 4855
rect 2011 4821 2045 4855
rect 2079 4821 2113 4855
rect 2147 4821 2181 4855
rect 2215 4821 2249 4855
rect 2283 4821 2317 4855
rect 2351 4821 2385 4855
rect 2419 4821 2453 4855
rect 2487 4821 2521 4855
rect 2555 4821 3971 4855
rect 3983 4821 4017 4855
rect 4051 4821 4085 4855
rect 4119 4821 4153 4855
rect 4187 4821 4221 4855
rect 4255 4821 4289 4855
rect 4323 4821 4357 4855
rect 4391 4821 4425 4855
rect 4459 4821 4493 4855
rect 4527 4821 4561 4855
rect 4595 4821 4629 4855
rect 4663 4821 4697 4855
rect 4731 4821 4765 4855
rect 4799 4821 4833 4855
rect 4867 4821 4901 4855
rect 4935 4821 4969 4855
rect 5003 4821 5037 4855
rect 5071 4821 5105 4855
rect 5139 4821 5173 4855
rect 5207 4821 5241 4855
rect 5275 4821 5309 4855
rect 5343 4821 5377 4855
rect 5411 4821 5445 4855
rect 5479 4821 5513 4855
rect 5547 4821 5581 4855
rect 5615 4821 5649 4855
rect 5683 4821 5717 4855
rect 5751 4821 5785 4855
rect 5819 4821 5853 4855
rect 5887 4821 5921 4855
rect 5955 4821 5989 4855
rect 6023 4821 6057 4855
rect 6091 4821 6125 4855
rect 6159 4821 6193 4855
rect 6227 4821 6261 4855
rect 6295 4821 6329 4855
rect 6363 4821 6397 4855
rect 6431 4821 6465 4855
rect 6499 4821 6533 4855
rect 6567 4821 6601 4855
rect 6635 4821 6669 4855
rect 6703 4821 6737 4855
rect 6771 4821 6805 4855
rect 6839 4821 6873 4855
rect 6907 4821 6941 4855
rect 6975 4821 7009 4855
rect 7043 4821 7077 4855
rect 7111 4821 7145 4855
rect 7179 4821 7213 4855
rect 7247 4821 7281 4855
rect 7315 4821 7349 4855
rect 7383 4821 7417 4855
rect 7451 4821 7485 4855
rect 7519 4821 7553 4855
rect 7587 4821 7621 4855
rect 7655 4821 7689 4855
rect 7723 4821 7757 4855
rect 7791 4821 7825 4855
rect 7859 4821 7893 4855
rect 7927 4821 7961 4855
rect 7995 4821 8029 4855
rect 8063 4821 8097 4855
rect 8131 4821 8165 4855
rect 8199 4821 8233 4855
rect 8267 4821 8301 4855
rect 8335 4821 8369 4855
rect 8403 4821 8437 4855
rect 8471 4821 8505 4855
rect 8539 4821 8573 4855
rect 8607 4821 8641 4855
rect 8675 4821 8709 4855
rect 8743 4821 8777 4855
rect 8811 4821 8845 4855
rect 8879 4821 8913 4855
rect 8947 4821 8981 4855
rect 9015 4821 9049 4855
rect 9083 4821 9117 4855
rect 9151 4821 9185 4855
rect 9219 4821 9253 4855
rect 9287 4821 9321 4855
rect 9355 4821 9389 4855
rect 9423 4821 9457 4855
rect 9491 4821 9525 4855
rect 9559 4821 9593 4855
rect 9627 4821 9661 4855
rect 9695 4821 9729 4855
rect 9763 4821 9797 4855
rect 9831 4821 9865 4855
rect 9899 4821 9933 4855
rect 9967 4821 10001 4855
rect 10035 4821 10069 4855
rect 10103 4821 10137 4855
rect 10171 4821 10205 4855
rect 10239 4821 10273 4855
rect 10307 4821 10341 4855
rect 10375 4821 10409 4855
rect 10443 4821 10477 4855
rect 10511 4821 10545 4855
rect 10579 4821 10613 4855
rect 10647 4821 10681 4855
rect 10715 4821 10749 4855
rect 10783 4821 10817 4855
rect 10851 4821 10885 4855
rect 10919 4821 10953 4855
rect 10987 4821 11021 4855
rect 11055 4821 11089 4855
rect 11123 4821 11157 4855
rect 11191 4821 11225 4855
rect 11259 4821 11293 4855
rect 11327 4821 11361 4855
rect 11395 4821 11429 4855
rect 11463 4821 11497 4855
rect 11531 4821 11565 4855
rect 11599 4821 11633 4855
rect 11667 4821 11701 4855
rect 11735 4821 11769 4855
rect 11803 4821 11837 4855
rect 11871 4821 11905 4855
rect 11939 4821 11973 4855
rect 12007 4821 12041 4855
rect 12075 4821 12109 4855
rect 12143 4821 12177 4855
rect 93 4753 127 4787
rect 162 4753 196 4787
rect 231 4753 265 4787
rect 300 4753 334 4787
rect 369 4753 403 4787
rect 438 4753 472 4787
rect 507 4753 541 4787
rect 576 4753 610 4787
rect 645 4753 679 4787
rect 714 4753 748 4787
rect 783 4753 817 4787
rect 852 4753 886 4787
rect 921 4753 955 4787
rect 990 4753 1024 4787
rect 1059 4753 1093 4787
rect 1128 4753 1162 4787
rect 1197 4753 1231 4787
rect 1266 4753 1300 4787
rect 1335 4753 1369 4787
rect 1404 4753 1438 4787
rect 1473 4753 1507 4787
rect 1542 4753 1576 4787
rect 1611 4753 1645 4787
rect 1680 4753 1714 4787
rect 1749 4753 1783 4787
rect 1818 4753 1852 4787
rect 1887 4753 1921 4787
rect 1956 4753 1990 4787
rect 2025 4753 2059 4787
rect 2094 4753 2128 4787
rect 2163 4753 2197 4787
rect 2232 4753 2266 4787
rect 2301 4753 2335 4787
rect 2370 4753 2404 4787
rect 2439 4753 2473 4787
rect 2508 4753 2542 4787
rect -17 4719 17 4753
rect 93 4685 127 4719
rect 162 4685 196 4719
rect 231 4685 265 4719
rect 300 4685 334 4719
rect 369 4685 403 4719
rect 438 4685 472 4719
rect 507 4685 541 4719
rect 576 4685 610 4719
rect 645 4685 679 4719
rect 714 4685 748 4719
rect 783 4685 817 4719
rect 852 4685 886 4719
rect 921 4685 955 4719
rect 990 4685 1024 4719
rect 1059 4685 1093 4719
rect 1128 4685 1162 4719
rect 1197 4685 1231 4719
rect 1266 4685 1300 4719
rect 1335 4685 1369 4719
rect 1404 4685 1438 4719
rect 1473 4685 1507 4719
rect 1542 4685 1576 4719
rect 1611 4685 1645 4719
rect 1680 4685 1714 4719
rect 1749 4685 1783 4719
rect 1818 4685 1852 4719
rect 1887 4685 1921 4719
rect 1956 4685 1990 4719
rect 2025 4685 2059 4719
rect 2094 4685 2128 4719
rect 2163 4685 2197 4719
rect 2232 4685 2266 4719
rect 2301 4685 2335 4719
rect 2370 4685 2404 4719
rect 2439 4685 2473 4719
rect 2508 4685 2542 4719
rect -17 4651 17 4685
rect 93 4617 127 4651
rect 162 4617 196 4651
rect 231 4617 265 4651
rect 300 4617 334 4651
rect 369 4617 403 4651
rect 438 4617 472 4651
rect 507 4617 541 4651
rect 576 4617 610 4651
rect 645 4617 679 4651
rect 714 4617 748 4651
rect 783 4617 817 4651
rect 852 4617 886 4651
rect 921 4617 955 4651
rect 990 4617 1024 4651
rect 1059 4617 1093 4651
rect 1128 4617 1162 4651
rect 1197 4617 1231 4651
rect 1266 4617 1300 4651
rect 1335 4617 1369 4651
rect 1404 4617 1438 4651
rect 1473 4617 1507 4651
rect 1542 4617 1576 4651
rect 1611 4617 1645 4651
rect 1680 4617 1714 4651
rect 1749 4617 1783 4651
rect 1818 4617 1852 4651
rect 1887 4617 1921 4651
rect 1956 4617 1990 4651
rect 2025 4617 2059 4651
rect 2094 4617 2128 4651
rect 2163 4617 2197 4651
rect 2232 4617 2266 4651
rect 2301 4617 2335 4651
rect 2370 4617 2404 4651
rect 2439 4617 2473 4651
rect 2508 4617 2542 4651
rect 2577 4617 3971 4821
rect 4056 4718 4090 4752
rect 4126 4718 4160 4752
rect 4196 4718 4230 4752
rect 4266 4718 4300 4752
rect 4336 4718 4370 4752
rect 4406 4718 4440 4752
rect 4476 4718 4510 4752
rect 4546 4718 4580 4752
rect 4616 4718 4650 4752
rect 7857 4718 7891 4752
rect 7931 4718 7965 4752
rect 8005 4718 8039 4752
rect 8078 4718 8112 4752
rect 8151 4718 8185 4752
rect 8224 4718 8258 4752
rect 8297 4718 8331 4752
rect 8370 4718 8404 4752
rect -17 4583 17 4617
rect -17 4515 17 4549
rect 93 4547 127 4581
rect 167 4547 201 4581
rect 241 4547 275 4581
rect 315 4547 349 4581
rect 388 4547 422 4581
rect 461 4547 495 4581
rect 534 4547 568 4581
rect 607 4547 641 4581
rect 680 4547 714 4581
rect 753 4547 787 4581
rect 7857 4629 7891 4663
rect 7931 4629 7965 4663
rect 8005 4629 8039 4663
rect 8078 4629 8112 4663
rect 8151 4629 8185 4663
rect 8224 4629 8258 4663
rect 8297 4629 8331 4663
rect 8370 4629 8404 4663
rect -17 4447 17 4481
rect 93 4479 127 4513
rect 167 4479 201 4513
rect 241 4479 275 4513
rect 315 4479 349 4513
rect 388 4479 422 4513
rect 461 4479 495 4513
rect 534 4479 568 4513
rect 607 4479 641 4513
rect 680 4479 714 4513
rect 753 4479 787 4513
rect -17 4379 17 4413
rect 93 4411 127 4445
rect 167 4411 201 4445
rect 241 4411 275 4445
rect 315 4411 349 4445
rect 388 4411 422 4445
rect 461 4411 495 4445
rect 534 4411 568 4445
rect 607 4411 641 4445
rect 680 4411 714 4445
rect 753 4411 787 4445
rect 7857 4561 7891 4595
rect 7931 4561 7965 4595
rect 8005 4561 8039 4595
rect 8078 4561 8112 4595
rect 8151 4561 8185 4595
rect 8224 4561 8258 4595
rect 8297 4561 8331 4595
rect 8370 4561 8404 4595
rect 7857 4493 7891 4527
rect 7931 4493 7965 4527
rect 8005 4493 8039 4527
rect 8078 4493 8112 4527
rect 8151 4493 8185 4527
rect 8224 4493 8258 4527
rect 8297 4493 8331 4527
rect 8370 4493 8404 4527
rect 7857 4425 7891 4459
rect 7931 4425 7965 4459
rect 8005 4425 8039 4459
rect 8078 4425 8112 4459
rect 8151 4425 8185 4459
rect 8224 4425 8258 4459
rect 8297 4425 8331 4459
rect 8370 4425 8404 4459
rect -17 4311 17 4345
rect 140 4343 174 4377
rect -17 4243 17 4277
rect 140 4275 174 4309
rect -17 4175 17 4209
rect 140 4207 174 4241
rect -17 4107 17 4141
rect 140 4139 174 4173
rect -17 4039 17 4073
rect 140 4071 174 4105
rect -17 3971 17 4005
rect 140 4003 174 4037
rect -17 3903 17 3937
rect 140 3935 174 3969
rect -17 3835 17 3869
rect 140 3867 174 3901
rect -17 3767 17 3801
rect 140 3799 174 3833
rect -17 3699 17 3733
rect 140 3731 174 3765
rect -17 3631 17 3665
rect 140 3663 174 3697
rect -17 3563 17 3597
rect 140 3595 174 3629
rect -17 3495 17 3529
rect 140 3527 174 3561
rect -17 3427 17 3461
rect 140 3459 174 3493
rect -17 3359 17 3393
rect 140 3391 174 3425
rect -17 3291 17 3325
rect 140 3323 174 3357
rect -17 3223 17 3257
rect 140 3255 174 3289
rect -17 3155 17 3189
rect 140 3187 174 3221
rect -17 3087 17 3121
rect 140 3118 174 3152
rect -17 3019 17 3053
rect 140 3049 174 3083
rect -17 2951 17 2985
rect 140 2980 174 3014
rect -17 2883 17 2917
rect 140 2911 174 2945
rect -17 2815 17 2849
rect 140 2842 174 2876
rect -17 2747 17 2781
rect 140 2773 174 2807
rect -17 2679 17 2713
rect 140 2704 174 2738
rect -17 2611 17 2645
rect 140 2635 174 2669
rect -17 2543 17 2577
rect 140 2566 174 2600
rect -17 2475 17 2509
rect 140 2497 174 2531
rect -17 2407 17 2441
rect 140 2428 174 2462
rect -17 2338 17 2372
rect 140 2359 174 2393
rect 14983 2452 15017 2486
rect 14983 2384 15017 2418
rect -17 2269 17 2303
rect 140 2290 174 2324
rect 14983 2316 15017 2350
rect -17 2200 17 2234
rect 140 2221 174 2255
rect -17 2131 17 2165
rect 140 2152 174 2186
rect 3200 2140 3234 2174
rect 3271 2140 3305 2174
rect 3342 2140 3376 2174
rect 3413 2140 3447 2174
rect 3484 2140 3518 2174
rect 3555 2140 3589 2174
rect 3626 2140 3660 2174
rect 3697 2140 3731 2174
rect 3768 2140 3802 2174
rect 3839 2140 3873 2174
rect 3910 2140 3944 2174
rect 3981 2140 4015 2174
rect 4052 2140 4086 2174
rect 4123 2140 4157 2174
rect 4194 2140 4228 2174
rect 4265 2140 4299 2174
rect 4336 2140 4370 2174
rect 4406 2140 4440 2174
rect -17 2062 17 2096
rect 140 2083 174 2117
rect -17 1993 17 2027
rect 140 2014 174 2048
rect -17 1924 17 1958
rect 145 1946 179 1980
rect 213 1946 247 1980
rect 281 1946 315 1980
rect 349 1946 383 1980
rect 417 1946 451 1980
rect 485 1946 519 1980
rect 553 1946 587 1980
rect -17 1855 17 1889
rect 145 1875 179 1909
rect 213 1875 247 1909
rect 281 1875 315 1909
rect 349 1875 383 1909
rect 417 1875 451 1909
rect 485 1875 519 1909
rect 553 1875 587 1909
rect -17 1786 17 1820
rect 145 1804 179 1838
rect 213 1804 247 1838
rect 281 1804 315 1838
rect 349 1804 383 1838
rect 417 1804 451 1838
rect 485 1804 519 1838
rect 553 1804 587 1838
rect -17 1717 17 1751
rect 145 1733 179 1767
rect 213 1733 247 1767
rect 281 1733 315 1767
rect 349 1733 383 1767
rect 417 1733 451 1767
rect 485 1733 519 1767
rect 553 1733 587 1767
rect -17 1648 17 1682
rect 145 1662 179 1696
rect 213 1662 247 1696
rect 281 1662 315 1696
rect 349 1662 383 1696
rect 417 1662 451 1696
rect 485 1662 519 1696
rect 553 1662 587 1696
rect -17 1579 17 1613
rect 145 1591 179 1625
rect 213 1591 247 1625
rect 281 1591 315 1625
rect 349 1591 383 1625
rect 417 1591 451 1625
rect 485 1591 519 1625
rect 553 1591 587 1625
rect -17 1510 17 1544
rect 145 1520 179 1554
rect 213 1520 247 1554
rect 281 1520 315 1554
rect 349 1520 383 1554
rect 417 1520 451 1554
rect 485 1520 519 1554
rect 553 1520 587 1554
rect -17 1441 17 1475
rect 145 1449 179 1483
rect 213 1449 247 1483
rect 281 1449 315 1483
rect 349 1449 383 1483
rect 417 1449 451 1483
rect 485 1449 519 1483
rect 553 1449 587 1483
rect -17 1372 17 1406
rect 145 1378 179 1412
rect 213 1378 247 1412
rect 281 1378 315 1412
rect 349 1378 383 1412
rect 417 1378 451 1412
rect 485 1378 519 1412
rect 553 1378 587 1412
rect -17 1303 17 1337
rect 145 1308 179 1342
rect 213 1308 247 1342
rect 281 1308 315 1342
rect 349 1308 383 1342
rect 417 1308 451 1342
rect 485 1308 519 1342
rect 553 1308 587 1342
rect -17 1234 17 1268
rect 145 1238 179 1272
rect 213 1238 247 1272
rect 281 1238 315 1272
rect 349 1238 383 1272
rect 417 1238 451 1272
rect 485 1238 519 1272
rect 553 1238 587 1272
rect -17 1165 17 1199
rect 145 1168 179 1202
rect 213 1168 247 1202
rect 281 1168 315 1202
rect 349 1168 383 1202
rect 417 1168 451 1202
rect 485 1168 519 1202
rect 553 1168 587 1202
rect -17 1096 17 1130
rect 145 1098 179 1132
rect 213 1098 247 1132
rect 281 1098 315 1132
rect 349 1098 383 1132
rect 417 1098 451 1132
rect 485 1098 519 1132
rect 553 1098 587 1132
rect 8853 1896 8887 1930
rect 8921 1896 8955 1930
rect 8989 1896 9023 1930
rect 8853 1826 8887 1860
rect 8921 1826 8955 1860
rect 8989 1826 9023 1860
rect 8853 1756 8887 1790
rect 8921 1756 8955 1790
rect 8989 1756 9023 1790
rect 9171 1896 9205 1930
rect 9171 1795 9205 1829
rect 10184 1803 10490 2245
rect 14983 2248 15017 2282
rect 14983 2180 15017 2214
rect 14983 2112 15017 2146
rect 14983 2044 15017 2078
rect 14983 1976 15017 2010
rect 14983 1908 15017 1942
rect 14983 1840 15017 1874
rect 14983 1772 15017 1806
rect 8853 1687 8887 1721
rect 8921 1687 8955 1721
rect 8989 1687 9023 1721
rect 8853 1618 8887 1652
rect 8921 1618 8955 1652
rect 8989 1618 9023 1652
rect 8853 1549 8887 1583
rect 8921 1549 8955 1583
rect 8989 1549 9023 1583
rect 8853 1480 8887 1514
rect 8921 1480 8955 1514
rect 8989 1480 9023 1514
rect 8853 1411 8887 1445
rect 8921 1411 8955 1445
rect 8989 1411 9023 1445
rect 8853 1342 8887 1376
rect 8921 1342 8955 1376
rect 8989 1342 9023 1376
rect 8853 1273 8887 1307
rect 8921 1273 8955 1307
rect 8989 1273 9023 1307
rect 8853 1204 8887 1238
rect 8921 1204 8955 1238
rect 8989 1204 9023 1238
rect 8853 1135 8887 1169
rect 8921 1135 8955 1169
rect 8989 1135 9023 1169
rect 8853 1066 8887 1100
rect 8921 1066 8955 1100
rect 8989 1066 9023 1100
rect -17 1027 17 1061
rect 145 1028 179 1062
rect 213 1028 247 1062
rect 281 1028 315 1062
rect 349 1028 383 1062
rect 417 1028 451 1062
rect 485 1028 519 1062
rect 553 1028 587 1062
rect -17 958 17 992
rect 8853 997 8887 1031
rect 8921 997 8955 1031
rect 8989 997 9023 1031
rect 14983 1704 15017 1738
rect 14983 1636 15017 1670
rect 14983 1568 15017 1602
rect 14983 1500 15017 1534
rect 14983 1432 15017 1466
rect 14983 1364 15017 1398
rect 14983 1296 15017 1330
rect 14983 1228 15017 1262
rect 14983 1160 15017 1194
rect 14983 1092 15017 1126
rect 14983 1024 15017 1058
rect -17 889 17 923
rect -17 820 17 854
rect -17 751 17 785
rect 14983 956 15017 990
rect 14983 888 15017 922
rect 14983 820 15017 854
rect 14983 752 15017 786
rect 14983 684 15017 718
rect 14983 616 15017 650
rect 14983 548 15017 582
rect 14983 480 15017 514
rect 14983 412 15017 446
rect 14983 344 15017 378
rect 14983 276 15017 310
rect 14983 208 15017 242
rect 14983 140 15017 174
<< locali >>
rect -17 4821 43 4855
rect 77 4821 151 4855
rect 185 4821 220 4855
rect 254 4821 289 4855
rect 323 4821 358 4855
rect 392 4821 427 4855
rect 461 4821 496 4855
rect 530 4821 565 4855
rect 599 4821 634 4855
rect 668 4821 703 4855
rect 737 4821 772 4855
rect 806 4821 841 4855
rect 875 4821 910 4855
rect 944 4821 979 4855
rect 1013 4821 1048 4855
rect 1082 4821 1117 4855
rect 1151 4821 1186 4855
rect 1220 4821 1255 4855
rect 1289 4821 1324 4855
rect 1358 4821 1393 4855
rect 1427 4821 1462 4855
rect 1496 4821 1531 4855
rect 1565 4821 1600 4855
rect 1634 4821 1669 4855
rect 1703 4821 1738 4855
rect 1772 4821 1807 4855
rect 1841 4821 1875 4855
rect 1909 4821 1943 4855
rect 1977 4821 2011 4855
rect 2045 4821 2079 4855
rect 2113 4821 2147 4855
rect 2181 4821 2215 4855
rect 2249 4821 2283 4855
rect 2317 4821 2351 4855
rect 2385 4821 2419 4855
rect 2453 4821 2487 4855
rect 2521 4821 2555 4855
rect 3971 4821 3983 4855
rect 4017 4821 4051 4855
rect 4085 4821 4119 4855
rect 4153 4821 4187 4855
rect 4221 4821 4255 4855
rect 4289 4821 4323 4855
rect 4357 4821 4391 4855
rect 4425 4821 4459 4855
rect 4493 4821 4527 4855
rect 4561 4821 4595 4855
rect 4629 4821 4663 4855
rect 4697 4821 4731 4855
rect 4765 4821 4799 4855
rect 4833 4821 4867 4855
rect 4901 4821 4935 4855
rect 4969 4821 5003 4855
rect 5037 4821 5071 4855
rect 5105 4821 5139 4855
rect 5173 4821 5207 4855
rect 5241 4821 5275 4855
rect 5309 4821 5343 4855
rect 5377 4821 5411 4855
rect 5445 4821 5479 4855
rect 5513 4821 5547 4855
rect 5581 4821 5615 4855
rect 5649 4821 5683 4855
rect 5717 4821 5751 4855
rect 5785 4821 5819 4855
rect 5853 4821 5887 4855
rect 5921 4821 5955 4855
rect 5989 4821 6023 4855
rect 6057 4821 6091 4855
rect 6125 4821 6159 4855
rect 6193 4821 6227 4855
rect 6261 4821 6295 4855
rect 6329 4821 6363 4855
rect 6397 4821 6431 4855
rect 6465 4821 6499 4855
rect 6533 4821 6567 4855
rect 6601 4821 6635 4855
rect 6669 4821 6703 4855
rect 6737 4821 6771 4855
rect 6805 4821 6839 4855
rect 6873 4821 6907 4855
rect 6941 4821 6975 4855
rect 7009 4821 7043 4855
rect 7077 4821 7111 4855
rect 7145 4821 7179 4855
rect 7213 4821 7247 4855
rect 7281 4821 7315 4855
rect 7349 4821 7383 4855
rect 7417 4821 7451 4855
rect 7485 4821 7519 4855
rect 7553 4821 7587 4855
rect 7621 4821 7655 4855
rect 7689 4821 7723 4855
rect 7757 4821 7791 4855
rect 7825 4821 7859 4855
rect 7893 4821 7927 4855
rect 7961 4821 7995 4855
rect 8029 4821 8063 4855
rect 8097 4821 8131 4855
rect 8165 4821 8199 4855
rect 8233 4821 8267 4855
rect 8301 4821 8335 4855
rect 8369 4821 8403 4855
rect 8437 4821 8471 4855
rect 8505 4821 8539 4855
rect 8573 4821 8607 4855
rect 8641 4821 8675 4855
rect 8709 4821 8743 4855
rect 8777 4821 8811 4855
rect 8845 4821 8879 4855
rect 8913 4821 8947 4855
rect 8981 4821 9015 4855
rect 9049 4821 9083 4855
rect 9117 4821 9151 4855
rect 9185 4821 9219 4855
rect 9253 4821 9287 4855
rect 9321 4821 9355 4855
rect 9389 4821 9423 4855
rect 9457 4821 9491 4855
rect 9525 4821 9559 4855
rect 9593 4821 9627 4855
rect 9661 4821 9695 4855
rect 9729 4821 9763 4855
rect 9797 4821 9831 4855
rect 9865 4821 9899 4855
rect 9933 4821 9967 4855
rect 10001 4821 10035 4855
rect 10069 4821 10103 4855
rect 10137 4821 10171 4855
rect 10205 4821 10239 4855
rect 10273 4821 10307 4855
rect 10341 4821 10375 4855
rect 10409 4821 10443 4855
rect 10477 4821 10511 4855
rect 10545 4821 10579 4855
rect 10613 4821 10647 4855
rect 10681 4821 10715 4855
rect 10749 4821 10783 4855
rect 10817 4821 10851 4855
rect 10885 4821 10919 4855
rect 10953 4821 10987 4855
rect 11021 4821 11055 4855
rect 11089 4821 11123 4855
rect 11157 4821 11191 4855
rect 11225 4821 11259 4855
rect 11293 4821 11327 4855
rect 11361 4821 11395 4855
rect 11429 4821 11463 4855
rect 11497 4821 11531 4855
rect 11565 4821 11599 4855
rect 11633 4821 11667 4855
rect 11701 4821 11735 4855
rect 11769 4821 11803 4855
rect 11837 4821 11871 4855
rect 11905 4821 11939 4855
rect 11973 4821 12007 4855
rect 12041 4821 12075 4855
rect 12109 4821 12143 4855
rect 12177 4821 12201 4855
rect -17 4787 2577 4821
rect -17 4753 93 4787
rect 127 4753 162 4787
rect 196 4753 231 4787
rect 265 4753 300 4787
rect 334 4753 369 4787
rect 403 4753 438 4787
rect 472 4753 507 4787
rect 541 4753 576 4787
rect 610 4753 645 4787
rect 679 4753 714 4787
rect 748 4753 783 4787
rect 817 4753 852 4787
rect 886 4753 921 4787
rect 955 4753 990 4787
rect 1024 4753 1059 4787
rect 1093 4753 1128 4787
rect 1162 4753 1197 4787
rect 1231 4753 1266 4787
rect 1300 4753 1335 4787
rect 1369 4753 1404 4787
rect 1438 4753 1473 4787
rect 1507 4753 1542 4787
rect 1576 4753 1611 4787
rect 1645 4753 1680 4787
rect 1714 4753 1749 4787
rect 1783 4753 1818 4787
rect 1852 4753 1887 4787
rect 1921 4753 1956 4787
rect 1990 4753 2025 4787
rect 2059 4753 2094 4787
rect 2128 4753 2163 4787
rect 2197 4753 2232 4787
rect 2266 4753 2301 4787
rect 2335 4753 2370 4787
rect 2404 4753 2439 4787
rect 2473 4753 2508 4787
rect 2542 4753 2577 4787
rect 17 4719 2577 4753
rect -17 4685 93 4719
rect 127 4685 162 4719
rect 196 4685 231 4719
rect 265 4685 300 4719
rect 334 4685 369 4719
rect 403 4685 438 4719
rect 472 4685 507 4719
rect 541 4685 576 4719
rect 610 4685 645 4719
rect 679 4685 714 4719
rect 748 4685 783 4719
rect 817 4685 852 4719
rect 886 4685 921 4719
rect 955 4685 990 4719
rect 1024 4685 1059 4719
rect 1093 4685 1128 4719
rect 1162 4685 1197 4719
rect 1231 4685 1266 4719
rect 1300 4685 1335 4719
rect 1369 4685 1404 4719
rect 1438 4685 1473 4719
rect 1507 4685 1542 4719
rect 1576 4685 1611 4719
rect 1645 4685 1680 4719
rect 1714 4685 1749 4719
rect 1783 4685 1818 4719
rect 1852 4685 1887 4719
rect 1921 4685 1956 4719
rect 1990 4685 2025 4719
rect 2059 4685 2094 4719
rect 2128 4685 2163 4719
rect 2197 4685 2232 4719
rect 2266 4685 2301 4719
rect 2335 4685 2370 4719
rect 2404 4685 2439 4719
rect 2473 4685 2508 4719
rect 2542 4685 2577 4719
rect 17 4651 2577 4685
rect -17 4617 93 4651
rect 127 4617 162 4651
rect 196 4617 231 4651
rect 265 4617 300 4651
rect 334 4617 369 4651
rect 403 4617 438 4651
rect 472 4617 507 4651
rect 541 4617 576 4651
rect 610 4617 645 4651
rect 679 4617 714 4651
rect 748 4617 783 4651
rect 817 4617 852 4651
rect 886 4617 921 4651
rect 955 4617 990 4651
rect 1024 4617 1059 4651
rect 1093 4617 1128 4651
rect 1162 4617 1197 4651
rect 1231 4617 1266 4651
rect 1300 4617 1335 4651
rect 1369 4617 1404 4651
rect 1438 4617 1473 4651
rect 1507 4617 1542 4651
rect 1576 4617 1611 4651
rect 1645 4617 1680 4651
rect 1714 4617 1749 4651
rect 1783 4617 1818 4651
rect 1852 4617 1887 4651
rect 1921 4617 1956 4651
rect 1990 4617 2025 4651
rect 2059 4617 2094 4651
rect 2128 4617 2163 4651
rect 2197 4617 2232 4651
rect 2266 4617 2301 4651
rect 2335 4617 2370 4651
rect 2404 4617 2439 4651
rect 2473 4617 2508 4651
rect 2542 4617 2577 4651
rect 3971 4752 4674 4821
rect 3971 4718 4056 4752
rect 4090 4718 4126 4752
rect 4160 4718 4196 4752
rect 4230 4718 4266 4752
rect 4300 4718 4336 4752
rect 4370 4718 4406 4752
rect 4440 4718 4476 4752
rect 4510 4718 4546 4752
rect 4580 4718 4616 4752
rect 4650 4718 4674 4752
rect 3971 4695 4674 4718
rect 7833 4752 8428 4821
rect 7833 4718 7857 4752
rect 7891 4718 7931 4752
rect 7965 4718 8005 4752
rect 8039 4718 8078 4752
rect 8112 4718 8151 4752
rect 8185 4718 8224 4752
rect 8258 4718 8297 4752
rect 8331 4718 8370 4752
rect 8404 4718 8428 4752
rect 11990 4736 12503 4776
rect 3971 4617 3995 4695
rect 4638 4634 4672 4695
rect 7833 4663 8428 4718
rect 17 4583 3995 4617
rect -17 4581 3995 4583
rect -17 4549 93 4581
rect 17 4547 93 4549
rect 127 4547 167 4581
rect 201 4547 241 4581
rect 275 4547 315 4581
rect 349 4547 388 4581
rect 422 4547 461 4581
rect 495 4547 534 4581
rect 568 4547 607 4581
rect 641 4547 680 4581
rect 714 4547 753 4581
rect 787 4556 3995 4581
rect 7833 4629 7857 4663
rect 7891 4629 7931 4663
rect 7965 4629 8005 4663
rect 8039 4629 8078 4663
rect 8112 4629 8151 4663
rect 8185 4629 8224 4663
rect 8258 4629 8297 4663
rect 8331 4629 8370 4663
rect 8404 4629 8428 4663
rect 7833 4595 8428 4629
rect 7833 4561 7857 4595
rect 7891 4561 7931 4595
rect 7965 4561 8005 4595
rect 8039 4561 8078 4595
rect 8112 4561 8151 4595
rect 8185 4561 8224 4595
rect 8258 4561 8297 4595
rect 8331 4561 8370 4595
rect 8404 4561 8428 4595
rect 787 4547 811 4556
rect 17 4513 811 4547
rect 17 4510 93 4513
rect -17 4481 93 4510
rect 17 4479 93 4481
rect 127 4479 167 4513
rect 201 4479 241 4513
rect 275 4479 315 4513
rect 349 4479 388 4513
rect 422 4479 461 4513
rect 495 4479 534 4513
rect 568 4479 607 4513
rect 641 4479 680 4513
rect 714 4479 753 4513
rect 787 4479 811 4513
rect 17 4445 811 4479
rect 4638 4479 4672 4517
rect 7038 4479 7072 4517
rect 7833 4527 8428 4561
rect 7833 4493 7857 4527
rect 7891 4493 7931 4527
rect 7965 4493 8005 4527
rect 8039 4493 8078 4527
rect 8112 4493 8151 4527
rect 8185 4493 8224 4527
rect 8258 4493 8297 4527
rect 8331 4493 8370 4527
rect 8404 4493 8428 4527
rect 7833 4459 8428 4493
rect 17 4438 93 4445
rect -17 4413 93 4438
rect 17 4411 93 4413
rect 127 4411 167 4445
rect 201 4411 241 4445
rect 275 4411 315 4445
rect 349 4411 388 4445
rect 422 4411 461 4445
rect 495 4411 534 4445
rect 568 4411 607 4445
rect 641 4411 680 4445
rect 714 4411 753 4445
rect 787 4411 811 4445
rect 7833 4425 7857 4459
rect 7891 4425 7931 4459
rect 7965 4425 8005 4459
rect 8039 4425 8078 4459
rect 8112 4425 8151 4459
rect 8185 4425 8224 4459
rect 8258 4425 8297 4459
rect 8331 4425 8370 4459
rect 8404 4425 8428 4459
rect 17 4379 197 4411
rect -17 4377 197 4379
rect -17 4345 140 4377
rect 17 4343 140 4345
rect 174 4343 197 4377
rect 17 4311 197 4343
rect -17 4309 197 4311
rect -17 4277 140 4309
rect 17 4275 140 4277
rect 174 4275 197 4309
rect 364 4299 398 4411
rect 716 4299 750 4411
rect 7833 4392 8428 4425
rect 17 4243 197 4275
rect -17 4241 197 4243
rect -17 4209 140 4241
rect 17 4207 140 4209
rect 174 4207 197 4241
rect 17 4175 197 4207
rect -17 4173 197 4175
rect -17 4141 140 4173
rect 17 4139 140 4141
rect 174 4139 197 4173
rect 17 4107 197 4139
rect -17 4105 197 4107
rect -17 4073 140 4105
rect 17 4071 140 4073
rect 174 4071 197 4105
rect 17 4039 197 4071
rect -17 4037 197 4039
rect -17 4005 140 4037
rect 17 4003 140 4005
rect 174 4003 197 4037
rect 17 3971 197 4003
rect -17 3969 197 3971
rect -17 3937 140 3969
rect 17 3935 140 3937
rect 174 3935 197 3969
rect 17 3903 197 3935
rect -17 3901 197 3903
rect -17 3893 140 3901
rect 17 3867 140 3893
rect 174 3867 197 3901
rect 17 3835 197 3867
rect -17 3833 197 3835
rect -17 3821 140 3833
rect 17 3799 140 3821
rect 174 3799 197 3833
rect 17 3767 197 3799
rect -17 3765 197 3767
rect -17 3749 140 3765
rect 17 3731 140 3749
rect 174 3731 197 3765
rect 17 3699 197 3731
rect -17 3697 197 3699
rect -17 3665 140 3697
rect 17 3663 140 3665
rect 174 3663 197 3697
rect 17 3631 197 3663
rect -17 3629 197 3631
rect -17 3597 140 3629
rect 17 3595 140 3597
rect 174 3595 197 3629
rect 7122 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 7256 3669
rect 9440 3642 9454 3669
rect 7122 3605 7256 3635
rect 9434 3635 9454 3642
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 17 3563 197 3595
rect 7603 3567 7653 3601
rect 7885 3580 7896 3595
rect -17 3561 197 3563
rect 7930 3561 7968 3595
rect 8002 3580 8019 3595
rect -17 3529 140 3561
rect 17 3527 140 3529
rect 174 3527 197 3561
rect 8183 3556 8233 3590
rect 9132 3580 9144 3595
rect 9178 3561 9216 3595
rect 9250 3580 9266 3595
rect 9434 3582 9704 3635
rect 10031 3549 10069 3583
rect 10103 3549 10141 3583
rect 17 3495 197 3527
rect 8648 3519 8765 3548
rect -17 3493 197 3495
rect -17 3461 140 3493
rect 17 3459 140 3461
rect 174 3459 197 3493
rect 8693 3485 8731 3519
rect 17 3427 197 3459
rect -17 3425 197 3427
rect -17 3393 140 3425
rect 17 3391 140 3393
rect 174 3391 197 3425
rect 17 3359 197 3391
rect -17 3357 197 3359
rect -17 3325 140 3357
rect 17 3323 140 3325
rect 174 3323 197 3357
rect 17 3291 197 3323
rect -17 3289 197 3291
rect -17 3257 140 3289
rect 17 3255 140 3257
rect 174 3255 197 3289
rect 17 3223 197 3255
rect -17 3221 197 3223
rect -17 3189 140 3221
rect 17 3187 140 3189
rect 174 3187 197 3221
rect 17 3155 197 3187
rect -17 3152 197 3155
rect -17 3121 140 3152
rect 17 3118 140 3121
rect 174 3118 197 3152
rect 9171 3475 9281 3499
rect 9171 3441 9175 3475
rect 9209 3441 9243 3475
rect 9277 3441 9281 3475
rect 9171 3401 9281 3441
rect 9171 3372 9175 3401
rect 9209 3372 9243 3401
rect 9277 3372 9281 3401
rect 9171 3194 9173 3372
rect 9279 3194 9281 3372
rect 9171 3179 9281 3194
rect 9171 3145 9175 3179
rect 9209 3145 9243 3179
rect 9277 3145 9281 3179
rect 17 3087 197 3118
rect -17 3083 197 3087
rect -17 3053 140 3083
rect 17 3049 140 3053
rect 174 3049 197 3083
rect 17 3019 197 3049
rect -17 3014 197 3019
rect -17 2985 140 3014
rect 17 2980 140 2985
rect 174 2980 197 3014
rect 17 2951 197 2980
rect -17 2945 197 2951
rect -17 2917 140 2945
rect 17 2911 140 2917
rect 174 2911 197 2945
rect 17 2883 197 2911
rect -17 2876 197 2883
rect -17 2849 140 2876
rect 17 2842 140 2849
rect 174 2842 197 2876
rect 17 2815 197 2842
rect -17 2807 197 2815
rect -17 2781 140 2807
rect 17 2773 140 2781
rect 174 2773 197 2807
rect 17 2747 197 2773
rect -17 2738 197 2747
rect -17 2713 140 2738
rect 17 2704 140 2713
rect 174 2704 197 2738
rect 17 2679 197 2704
rect -17 2669 197 2679
rect -17 2645 140 2669
rect 17 2635 140 2645
rect 174 2635 197 2669
rect 17 2611 197 2635
rect -17 2600 197 2611
rect -17 2577 140 2600
rect 17 2566 140 2577
rect 174 2566 197 2600
rect 17 2543 197 2566
rect -17 2531 197 2543
rect -17 2509 140 2531
rect 17 2497 140 2509
rect 174 2497 197 2531
rect 17 2475 197 2497
rect -17 2462 197 2475
rect -17 2441 140 2462
rect 17 2428 140 2441
rect 174 2428 197 2462
rect 17 2407 197 2428
rect -17 2393 197 2407
rect -17 2372 140 2393
rect 17 2359 140 2372
rect 174 2359 197 2393
rect 17 2338 197 2359
rect -17 2324 197 2338
rect 408 3094 986 3118
rect 442 3060 476 3094
rect 510 3060 544 3094
rect 578 3060 612 3094
rect 646 3060 680 3094
rect 714 3060 748 3094
rect 782 3060 816 3094
rect 850 3060 884 3094
rect 918 3060 952 3094
rect 408 3023 986 3060
rect 442 2989 476 3023
rect 510 2989 544 3023
rect 578 2989 612 3023
rect 646 2989 680 3023
rect 714 2989 748 3023
rect 782 2989 816 3023
rect 850 2989 884 3023
rect 918 2989 952 3023
rect 408 2952 986 2989
rect 442 2918 476 2952
rect 510 2918 544 2952
rect 578 2918 612 2952
rect 646 2918 680 2952
rect 714 2918 748 2952
rect 782 2918 816 2952
rect 850 2918 884 2952
rect 918 2918 952 2952
rect 408 2882 986 2918
rect 9171 3105 9281 3145
rect 9171 3071 9175 3105
rect 9209 3071 9243 3105
rect 9277 3071 9281 3105
rect 9171 3031 9281 3071
rect 9171 2997 9175 3031
rect 9209 2997 9243 3031
rect 9277 2997 9281 3031
rect 9171 2957 9281 2997
rect 9171 2923 9175 2957
rect 9209 2923 9243 2957
rect 9277 2923 9281 2957
rect 9171 2899 9281 2923
rect 442 2848 476 2882
rect 510 2848 544 2882
rect 578 2848 612 2882
rect 646 2848 680 2882
rect 714 2848 748 2882
rect 782 2848 816 2882
rect 850 2848 884 2882
rect 918 2848 952 2882
rect 408 2812 986 2848
rect 442 2778 476 2812
rect 510 2778 544 2812
rect 578 2778 612 2812
rect 646 2778 680 2812
rect 714 2778 748 2812
rect 782 2778 816 2812
rect 850 2778 884 2812
rect 918 2778 952 2812
rect 408 2742 986 2778
rect 442 2708 476 2742
rect 510 2708 544 2742
rect 578 2708 612 2742
rect 646 2708 680 2742
rect 714 2708 748 2742
rect 782 2708 816 2742
rect 850 2708 884 2742
rect 918 2708 952 2742
rect 408 2672 986 2708
rect 442 2638 476 2672
rect 510 2638 544 2672
rect 578 2638 612 2672
rect 646 2638 680 2672
rect 714 2638 748 2672
rect 782 2638 816 2672
rect 850 2638 884 2672
rect 918 2638 952 2672
rect 408 2602 986 2638
rect 442 2568 476 2602
rect 510 2568 544 2602
rect 578 2568 612 2602
rect 646 2568 680 2602
rect 714 2568 748 2602
rect 782 2568 816 2602
rect 850 2568 884 2602
rect 918 2568 952 2602
rect 408 2532 986 2568
rect 442 2498 476 2532
rect 510 2498 544 2532
rect 578 2498 612 2532
rect 646 2498 680 2532
rect 714 2498 748 2532
rect 782 2498 816 2532
rect 850 2498 884 2532
rect 918 2498 952 2532
rect 408 2462 986 2498
rect 442 2428 476 2462
rect 510 2428 544 2462
rect 578 2428 612 2462
rect 646 2428 680 2462
rect 714 2428 748 2462
rect 782 2428 816 2462
rect 850 2428 884 2462
rect 918 2428 952 2462
rect 408 2392 986 2428
rect 442 2358 476 2392
rect 510 2358 544 2392
rect 578 2358 612 2392
rect 646 2358 680 2392
rect 714 2358 748 2392
rect 782 2358 816 2392
rect 850 2358 884 2392
rect 918 2358 952 2392
rect 408 2334 986 2358
rect 14983 2486 15038 2520
rect 14983 2418 15017 2452
rect 14983 2350 15017 2384
rect -17 2303 140 2324
rect 17 2290 140 2303
rect 174 2290 197 2324
rect 17 2269 197 2290
rect 14983 2282 15017 2316
rect -17 2255 197 2269
rect -17 2234 140 2255
rect 17 2221 140 2234
rect 174 2221 197 2255
rect 17 2200 197 2221
rect -17 2186 197 2200
rect -17 2165 140 2186
rect 17 2152 140 2165
rect 174 2152 197 2186
rect 10184 2245 10563 2269
rect 17 2131 197 2152
rect 3176 2174 4464 2182
rect 3176 2140 3200 2174
rect 3234 2140 3271 2174
rect 3305 2140 3342 2174
rect 3376 2140 3413 2174
rect 3447 2140 3484 2174
rect 3518 2140 3555 2174
rect 3589 2140 3626 2174
rect 3660 2140 3697 2174
rect 3731 2140 3768 2174
rect 3802 2140 3839 2174
rect 3873 2140 3910 2174
rect 3944 2140 3981 2174
rect 4015 2140 4052 2174
rect 4086 2140 4123 2174
rect 4157 2140 4194 2174
rect 4228 2140 4265 2174
rect 4299 2140 4336 2174
rect 4370 2140 4406 2174
rect 4440 2140 4464 2174
rect 3176 2132 4464 2140
rect -17 2117 197 2131
rect -17 2096 140 2117
rect 17 2083 140 2096
rect 174 2083 197 2117
rect 17 2062 197 2083
rect -17 2048 197 2062
rect -17 2027 140 2048
rect 17 2014 140 2027
rect 174 2014 197 2048
rect 17 2004 197 2014
rect 3316 2008 3350 2132
rect 3628 2008 3662 2132
rect 17 1993 587 2004
rect -17 1980 587 1993
rect -17 1958 145 1980
rect 17 1946 145 1958
rect 179 1946 213 1980
rect 247 1946 281 1980
rect 315 1946 349 1980
rect 383 1946 417 1980
rect 451 1946 485 1980
rect 519 1946 553 1980
rect 17 1924 587 1946
rect -17 1909 587 1924
rect -17 1889 145 1909
rect 17 1875 145 1889
rect 179 1875 213 1909
rect 247 1875 281 1909
rect 315 1875 349 1909
rect 383 1875 417 1909
rect 451 1875 485 1909
rect 519 1875 553 1909
rect 17 1855 587 1875
rect -17 1838 587 1855
rect -17 1820 145 1838
rect 17 1804 145 1820
rect 179 1804 213 1838
rect 247 1804 281 1838
rect 315 1804 349 1838
rect 383 1804 417 1838
rect 451 1804 485 1838
rect 519 1804 553 1838
rect 17 1786 587 1804
rect -17 1767 587 1786
rect -17 1751 145 1767
rect 17 1733 145 1751
rect 179 1733 213 1767
rect 247 1733 281 1767
rect 315 1733 349 1767
rect 383 1733 417 1767
rect 451 1733 485 1767
rect 519 1733 553 1767
rect 17 1717 587 1733
rect -17 1696 587 1717
rect -17 1682 145 1696
rect 17 1662 145 1682
rect 179 1662 213 1696
rect 247 1662 281 1696
rect 315 1662 349 1696
rect 383 1662 417 1696
rect 451 1662 485 1696
rect 519 1662 553 1696
rect 17 1648 587 1662
rect -17 1625 587 1648
rect -17 1613 145 1625
rect 17 1591 145 1613
rect 179 1591 213 1625
rect 247 1591 281 1625
rect 315 1591 349 1625
rect 383 1591 417 1625
rect 451 1591 485 1625
rect 519 1591 553 1625
rect 17 1579 587 1591
rect -17 1554 587 1579
rect -17 1544 145 1554
rect 17 1520 145 1544
rect 179 1520 213 1554
rect 247 1520 281 1554
rect 315 1520 349 1554
rect 383 1520 417 1554
rect 451 1520 485 1554
rect 519 1520 553 1554
rect 17 1510 587 1520
rect -17 1483 587 1510
rect -17 1475 145 1483
rect 17 1449 145 1475
rect 179 1449 213 1483
rect 247 1449 281 1483
rect 315 1449 349 1483
rect 383 1449 417 1483
rect 451 1449 485 1483
rect 519 1449 553 1483
rect 17 1441 587 1449
rect -17 1412 587 1441
rect -17 1406 145 1412
rect 17 1378 145 1406
rect 179 1378 213 1412
rect 247 1378 281 1412
rect 315 1378 349 1412
rect 383 1378 417 1412
rect 451 1378 485 1412
rect 519 1378 553 1412
rect 17 1372 587 1378
rect -17 1342 587 1372
rect -17 1337 145 1342
rect 17 1308 145 1337
rect 179 1308 213 1342
rect 247 1308 281 1342
rect 315 1308 349 1342
rect 383 1308 417 1342
rect 451 1308 485 1342
rect 519 1308 553 1342
rect 17 1303 587 1308
rect -17 1272 587 1303
rect -17 1268 145 1272
rect 17 1238 145 1268
rect 179 1238 213 1272
rect 247 1238 281 1272
rect 315 1238 349 1272
rect 383 1238 417 1272
rect 451 1238 485 1272
rect 519 1238 553 1272
rect 17 1234 587 1238
rect -17 1202 587 1234
rect -17 1199 145 1202
rect 17 1168 145 1199
rect 179 1168 213 1202
rect 247 1168 281 1202
rect 315 1168 349 1202
rect 383 1168 417 1202
rect 451 1168 485 1202
rect 519 1168 553 1202
rect 17 1165 587 1168
rect -17 1132 587 1165
rect -17 1130 145 1132
rect 17 1098 145 1130
rect 179 1098 213 1132
rect 247 1098 281 1132
rect 315 1098 349 1132
rect 383 1098 417 1132
rect 451 1098 485 1132
rect 519 1098 553 1132
rect 17 1096 587 1098
rect -17 1062 587 1096
rect -17 1061 145 1062
rect 17 1028 145 1061
rect 179 1028 213 1062
rect 247 1028 281 1062
rect 315 1028 349 1062
rect 383 1028 417 1062
rect 451 1028 485 1062
rect 519 1028 553 1062
rect 17 1027 587 1028
rect -17 1004 587 1027
rect 3940 1008 4072 2132
rect 8463 1930 8701 1954
rect 8497 1896 8531 1930
rect 8565 1896 8599 1930
rect 8633 1896 8667 1930
rect 8463 1856 8701 1896
rect 8497 1822 8531 1856
rect 8565 1822 8599 1856
rect 8633 1822 8667 1856
rect 8463 1782 8701 1822
rect 8497 1748 8531 1782
rect 8565 1748 8599 1782
rect 8633 1748 8667 1782
rect 8463 1708 8701 1748
rect 8497 1674 8531 1708
rect 8565 1674 8599 1708
rect 8633 1674 8667 1708
rect 8463 1634 8701 1674
rect 8497 1600 8531 1634
rect 8565 1600 8599 1634
rect 8633 1600 8667 1634
rect 8463 1560 8701 1600
rect 8497 1526 8531 1560
rect 8565 1526 8599 1560
rect 8633 1526 8667 1560
rect 8463 1487 8701 1526
rect 8497 1453 8531 1487
rect 8565 1453 8599 1487
rect 8633 1453 8667 1487
rect 8463 1414 8701 1453
rect 8497 1380 8531 1414
rect 8565 1380 8599 1414
rect 8633 1380 8667 1414
rect 8463 1341 8701 1380
rect 8497 1307 8531 1341
rect 8565 1307 8599 1341
rect 8633 1307 8667 1341
rect 8463 1268 8701 1307
rect 8497 1234 8531 1268
rect 8565 1234 8599 1268
rect 8633 1234 8667 1268
rect 8463 1195 8701 1234
rect 8497 1161 8531 1195
rect 8565 1161 8599 1195
rect 8633 1161 8667 1195
rect 8463 1122 8701 1161
rect 8497 1088 8531 1122
rect 8565 1088 8599 1122
rect 8633 1088 8667 1122
rect 8463 1064 8701 1088
rect 8853 1930 9221 1954
rect 8887 1896 8921 1930
rect 8955 1896 8989 1930
rect 9023 1896 9171 1930
rect 9205 1896 9221 1930
rect 8853 1860 9221 1896
rect 8887 1826 8921 1860
rect 8955 1826 8989 1860
rect 9023 1829 9221 1860
rect 9023 1826 9171 1829
rect 8853 1795 9171 1826
rect 9205 1795 9221 1829
rect 8853 1790 9221 1795
rect 8887 1756 8921 1790
rect 8955 1756 8989 1790
rect 9023 1771 9221 1790
rect 10490 1803 10563 2245
rect 10184 1779 10563 1803
rect 8853 1721 9023 1756
rect 8887 1687 8921 1721
rect 8955 1687 8989 1721
rect 8853 1652 9023 1687
rect 8887 1618 8921 1652
rect 8955 1618 8989 1652
rect 8853 1583 9023 1618
rect 8887 1549 8921 1583
rect 8955 1549 8989 1583
rect 10195 1742 10563 1779
rect 10301 1564 10457 1742
rect 14983 2214 15017 2248
rect 14983 2146 15017 2180
rect 14983 2078 15017 2112
rect 14983 2010 15017 2044
rect 14983 1942 15017 1976
rect 14983 1874 15017 1908
rect 14983 1806 15017 1840
rect 14983 1742 15017 1772
rect 14983 1670 15017 1704
rect 14983 1602 15017 1636
rect 8853 1514 9023 1549
rect 8887 1480 8921 1514
rect 8955 1480 8989 1514
rect 8853 1445 9023 1480
rect 8887 1411 8921 1445
rect 8955 1411 8989 1445
rect 8853 1376 9023 1411
rect 8887 1342 8921 1376
rect 8955 1342 8989 1376
rect 8853 1307 9023 1342
rect 8887 1273 8921 1307
rect 8955 1273 8989 1307
rect 8853 1238 9023 1273
rect 8887 1204 8921 1238
rect 8955 1204 8989 1238
rect 8853 1169 9023 1204
rect 8887 1135 8921 1169
rect 8955 1135 8989 1169
rect 8853 1100 9023 1135
rect 8887 1066 8921 1100
rect 8955 1066 8989 1100
rect 8853 1031 9023 1066
rect -17 992 17 1004
rect 8887 997 8921 1031
rect 8955 997 8989 1031
rect 8853 973 9023 997
rect 14983 1534 15017 1564
rect 14983 1466 15017 1500
rect 14983 1398 15017 1432
rect 14983 1330 15017 1364
rect 14983 1262 15017 1296
rect 14983 1194 15017 1228
rect 14983 1126 15017 1160
rect 14983 1058 15017 1092
rect 14983 990 15017 1024
rect -17 923 17 958
rect -17 854 17 889
rect -17 785 17 820
rect 14983 922 15017 956
rect 14983 854 15017 888
rect 14983 786 15017 820
rect -17 727 17 751
rect 14893 752 14983 766
rect 14893 718 15017 752
rect 14893 684 14983 718
rect 14893 650 15017 684
rect 14893 616 14983 650
rect 14893 582 15017 616
rect 14893 548 14983 582
rect 14893 514 15017 548
rect 14893 480 14983 514
rect 14893 446 15017 480
rect 14893 412 14983 446
rect 14893 378 15017 412
rect 14893 344 14983 378
rect 14893 310 15017 344
rect 14893 276 14983 310
rect 14893 242 15017 276
rect 14893 208 14983 242
rect 14893 174 15017 208
rect 14893 140 14983 174
rect 14893 76 15017 140
<< viali >>
rect -17 4515 17 4544
rect -17 4510 17 4515
rect -17 4447 17 4472
rect -17 4438 17 4447
rect 4638 4517 4672 4551
rect 4638 4445 4672 4479
rect 7038 4517 7072 4551
rect 7038 4445 7072 4479
rect -17 3869 17 3893
rect -17 3859 17 3869
rect -17 3801 17 3821
rect -17 3787 17 3801
rect -17 3733 17 3749
rect -17 3715 17 3733
rect 7138 3635 7172 3669
rect 7210 3635 7244 3669
rect 9454 3635 9488 3669
rect 9526 3635 9560 3669
rect 9598 3635 9632 3669
rect 9670 3635 9704 3669
rect 7896 3561 7930 3595
rect 7968 3561 8002 3595
rect 9144 3561 9178 3595
rect 9216 3561 9250 3595
rect 9997 3549 10031 3583
rect 10069 3549 10103 3583
rect 10141 3549 10175 3583
rect 8659 3485 8693 3519
rect 8731 3485 8765 3519
rect 9173 3367 9175 3372
rect 9175 3367 9209 3372
rect 9209 3367 9243 3372
rect 9243 3367 9277 3372
rect 9277 3367 9279 3372
rect 9173 3327 9279 3367
rect 9173 3293 9175 3327
rect 9175 3293 9209 3327
rect 9209 3293 9243 3327
rect 9243 3293 9277 3327
rect 9277 3293 9279 3327
rect 9173 3253 9279 3293
rect 9173 3219 9175 3253
rect 9175 3219 9209 3253
rect 9209 3219 9243 3253
rect 9243 3219 9277 3253
rect 9277 3219 9279 3253
rect 9173 3194 9279 3219
rect 10195 1564 10301 1742
rect 10457 1564 10563 1742
rect 14983 1738 15017 1742
rect 14983 1708 15017 1738
rect 14983 1636 15017 1670
rect 14983 1568 15017 1598
rect 14983 1564 15017 1568
<< metal1 >>
rect 14655 4638 14695 4676
rect -23 4551 12576 4563
rect -23 4544 4638 4551
rect -23 4510 -17 4544
rect 17 4517 4638 4544
rect 4672 4517 7038 4551
rect 7072 4517 12576 4551
rect 17 4510 12576 4517
rect -23 4479 12576 4510
rect -23 4472 4638 4479
rect -23 4438 -17 4472
rect 17 4445 4638 4472
rect 4672 4445 7038 4479
rect 7072 4445 12576 4479
rect 17 4438 12576 4445
rect -23 4417 12576 4438
rect 10155 4327 10207 4333
rect 10155 4263 10207 4275
tri 10130 4233 10155 4258 se
rect 7138 4211 10155 4233
rect 13704 4223 13743 4244
rect 7138 4205 10207 4211
rect 7860 4131 7906 4177
rect 9102 4131 9148 4177
rect 10098 4089 10138 4135
rect 7668 4013 7708 4059
rect 5766 3933 5806 3979
rect 5902 3933 5943 3979
rect -23 3893 11740 3905
rect -23 3859 -17 3893
rect 17 3859 11740 3893
rect -23 3821 11740 3859
rect -23 3787 -17 3821
rect 17 3787 11740 3821
rect -23 3749 11740 3787
rect -23 3715 -17 3749
rect 17 3739 11740 3749
rect 17 3715 1511 3739
rect -23 3703 1511 3715
tri 1511 3703 1547 3739 nw
tri 1661 3703 1697 3739 ne
rect 1697 3703 11740 3739
rect 66 3629 103 3675
rect 6875 3669 9716 3675
rect 6927 3635 7138 3669
rect 7172 3635 7210 3669
rect 7244 3635 9454 3669
rect 9488 3635 9526 3669
rect 9560 3635 9598 3669
rect 9632 3635 9670 3669
rect 9704 3635 9716 3669
rect 6927 3629 9716 3635
rect 6875 3605 6927 3617
tri 6927 3604 6952 3629 nw
rect 7884 3595 9886 3601
tri 9886 3595 9892 3601 sw
rect 7884 3561 7896 3595
rect 7930 3561 7968 3595
rect 8002 3561 9144 3595
rect 9178 3561 9216 3595
rect 9250 3589 9892 3595
tri 9892 3589 9898 3595 sw
rect 9250 3583 9898 3589
tri 9898 3583 9904 3589 sw
rect 9985 3583 10085 3595
rect 10137 3583 10149 3595
rect 9250 3561 9904 3583
rect 7884 3555 9904 3561
tri 9904 3555 9932 3583 sw
rect 6875 3547 6927 3553
tri 9858 3549 9864 3555 ne
rect 9864 3549 9932 3555
tri 9932 3549 9938 3555 sw
rect 9985 3549 9997 3583
rect 10031 3549 10069 3583
rect 10137 3549 10141 3583
tri 9864 3547 9866 3549 ne
rect 9866 3547 9938 3549
tri 9938 3547 9940 3549 sw
tri 9866 3527 9886 3547 ne
rect 9886 3543 9940 3547
tri 9940 3543 9944 3547 sw
rect 9985 3543 10085 3549
rect 10137 3543 10149 3549
rect 10201 3543 10207 3595
rect 9886 3527 9944 3543
tri 9944 3527 9960 3543 sw
rect 8647 3519 9386 3527
rect 8647 3485 8659 3519
rect 8693 3485 8731 3519
rect 8765 3485 9386 3519
rect 8647 3475 9386 3485
rect 9438 3475 9450 3527
rect 9502 3475 9508 3527
tri 9886 3515 9898 3527 ne
rect 9898 3515 9960 3527
tri 9960 3515 9972 3527 sw
tri 9898 3475 9938 3515 ne
rect 9938 3475 12101 3515
tri 9938 3463 9950 3475 ne
rect 9950 3463 12101 3475
rect 12153 3463 12165 3515
rect 12217 3463 12223 3515
rect 0 3372 10260 3379
rect 0 3194 9173 3372
rect 9279 3334 10260 3372
tri 10260 3334 10305 3379 sw
tri 10471 3334 10516 3379 se
rect 10516 3334 12576 3379
rect 9279 3194 12576 3334
rect 0 3177 12576 3194
rect 0 2765 15001 2895
rect 9781 2307 9827 2353
rect 0 2149 15001 2279
rect 0 1742 15023 1754
rect 0 1564 10195 1742
rect 10301 1564 10457 1742
rect 10563 1708 14983 1742
rect 15017 1708 15023 1742
rect 10563 1670 15023 1708
rect 10563 1643 14983 1670
rect 10563 1564 11508 1643
rect 0 1552 11508 1564
rect 12095 1636 14983 1643
rect 15017 1636 15023 1670
rect 12095 1598 15023 1636
rect 12095 1564 14983 1598
rect 15017 1564 15023 1598
rect 12095 1552 15023 1564
rect 0 1100 14511 1228
rect 0 1026 10097 1100
<< via1 >>
rect 10155 4275 10207 4327
rect 10155 4211 10207 4263
rect 6875 3617 6927 3669
rect 6875 3553 6927 3605
rect 10085 3583 10137 3595
rect 10149 3583 10201 3595
rect 10085 3549 10103 3583
rect 10103 3549 10137 3583
rect 10149 3549 10175 3583
rect 10175 3549 10201 3583
rect 10085 3543 10137 3549
rect 10149 3543 10201 3549
rect 9386 3475 9438 3527
rect 9450 3475 9502 3527
rect 12101 3463 12153 3515
rect 12165 3463 12217 3515
<< metal2 >>
rect 10155 4327 10207 4333
rect 10155 4263 10207 4275
rect 6875 3669 6927 3675
rect 6875 3605 6927 3617
rect 6875 3535 6927 3553
tri 9451 3547 9456 3552 se
rect 9456 3547 9508 4061
tri 10130 3595 10155 3620 se
rect 10155 3595 10207 4211
rect 10324 3623 10382 3675
tri 9447 3543 9451 3547 se
rect 9451 3543 9508 3547
rect 10079 3543 10085 3595
rect 10137 3543 10149 3595
rect 10201 3543 10207 3595
tri 9439 3535 9447 3543 se
rect 9447 3535 9508 3543
tri 9431 3527 9439 3535 se
rect 9439 3527 9508 3535
rect 9380 3475 9386 3527
rect 9438 3475 9450 3527
rect 9502 3475 9508 3527
tri 9431 3463 9443 3475 ne
rect 9443 3463 9456 3475
rect 12095 3463 12101 3515
rect 12153 3463 12165 3515
rect 12217 3463 12223 3515
tri 9443 3450 9456 3463 ne
rect 9855 1940 9902 1992
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 17 -1 0 4544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 9250 0 1 3561
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 8002 0 1 3561
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 1 0 7138 0 1 3635
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 1 0 8659 0 1 3485
box 0 0 1 1
use L1M1_CDNS_5246887918558  L1M1_CDNS_5246887918558_0
timestamp 1707688321
transform 1 0 9173 0 -1 3372
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform -1 0 10175 0 1 3549
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 17 1 0 3715
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 15017 1 0 1564
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 1 0 9454 0 1 3635
box 0 0 1 1
use L1M1_CDNS_52468879185300  L1M1_CDNS_52468879185300_0
timestamp 1707688321
transform 0 -1 599 1 0 1564
box -12 -6 190 616
use L1M1_CDNS_52468879185301  L1M1_CDNS_52468879185301_0
timestamp 1707688321
transform 0 1 400 -1 0 2883
box -12 -6 118 616
use L1M1_CDNS_52468879185302  L1M1_CDNS_52468879185302_0
timestamp 1707688321
transform -1 0 8713 0 -1 1221
box -12 -6 262 184
use L1M1_CDNS_52468879185303  L1M1_CDNS_52468879185303_0
timestamp 1707688321
transform 0 -1 799 -1 0 4543
box -12 -6 118 472
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_0
timestamp 1707688321
transform 1 0 8845 0 -1 1747
box -12 -6 190 184
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1707688321
transform 0 1 10195 -1 0 1742
box 0 0 1 1
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_1
timestamp 1707688321
transform 0 1 10457 -1 0 1742
box 0 0 1 1
use L1M1_CDNS_524688791851402  L1M1_CDNS_524688791851402_0
timestamp 1707688321
transform -1 0 8455 0 -1 4544
box -12 -6 622 112
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 10207 -1 0 4333
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 9508 0 -1 3527
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 1 6875 1 0 3547
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 1 0 10079 0 -1 3595
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 1 0 12095 0 1 3463
box 0 0 1 1
use sky130_fd_io__sio_com_pdpredrvr_strong_slow  sky130_fd_io__sio_com_pdpredrvr_strong_slow_0
timestamp 1707688321
transform -1 0 9387 0 1 2797
box 0 0 872 1568
use sky130_fd_io__sio_com_pdpredrvr_weak  sky130_fd_io__sio_com_pdpredrvr_weak_0
timestamp 1707688321
transform -1 0 8515 0 1 2797
box -85 8 809 1568
use sky130_fd_io__sio_com_pupredrvr_strong_slow  sky130_fd_io__sio_com_pupredrvr_strong_slow_0
timestamp 1707688321
transform -1 0 10215 0 1 2797
box -85 0 913 1568
use sky130_fd_io__sio_com_pupredrvr_weak  sky130_fd_io__sio_com_pupredrvr_weak_0
timestamp 1707688321
transform -1 0 7791 0 1 2798
box 21 7 731 1967
use sky130_fd_io__sio_pdpredrvr_strong  sky130_fd_io__sio_pdpredrvr_strong_0
timestamp 1707688321
transform 1 0 509 0 1 691
box -6 38 14735 4493
use sky130_fd_io__sio_pupredrvr_strong  sky130_fd_io__sio_pupredrvr_strong_0
timestamp 1707688321
transform 1 0 66 0 1 2133
box -66 10 7230 2632
<< labels >>
flabel comment s 14689 2495 14689 2495 0 FreeSans 440 90 0 0 condiode
flabel comment s 560 2408 560 2408 0 FreeSans 300 0 0 0 condiode
flabel comment s 10707 3958 10707 3958 0 FreeSans 300 0 0 0 pden_h_n1
flabel comment s 9376 4044 9376 4044 0 FreeSans 300 0 0 0 pden_h_n1
flabel comment s 7497 3968 7497 3968 0 FreeSans 300 0 0 0 pden_h_n1
flabel comment s 7988 3576 7988 3576 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 9129 3579 9129 3579 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 10392 3490 10392 3490 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 8484 4228 8484 4228 0 FreeSans 300 0 0 0 puen_h1
flabel comment s 9328 4228 9328 4228 0 FreeSans 300 0 0 0 puen_h1
flabel metal1 s 5902 3933 5943 3979 3 FreeSans 300 0 0 0 pu_h_n<3>
port 4 nsew
flabel metal1 s 5766 3933 5806 3979 7 FreeSans 300 0 0 0 pu_h_n<2>
port 5 nsew
flabel metal1 s 10098 4089 10138 4135 3 FreeSans 300 0 0 0 pu_h_n<1>
port 6 nsew
flabel metal1 s 7668 4013 7708 4059 3 FreeSans 300 0 0 0 pu_h_n<0>
port 7 nsew
flabel metal1 s 9102 4131 9148 4177 3 FreeSans 300 0 0 0 pd_h<1>
port 8 nsew
flabel metal1 s 7860 4131 7906 4177 3 FreeSans 300 0 0 0 pd_h<0>
port 9 nsew
flabel metal1 s 9781 2307 9827 2353 3 FreeSans 300 0 0 0 slow_h
port 10 nsew
flabel metal1 s 12534 3177 12576 3379 7 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 11698 3703 11740 3905 7 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 12539 4417 12576 4563 7 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 14958 2765 15000 2895 7 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 14958 2149 15000 2279 7 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 14469 1100 14511 1228 7 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 14958 1552 15000 1754 7 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 0 1552 42 1754 3 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 0 1026 42 1228 3 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 0 2149 42 2279 3 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 0 2765 42 2895 3 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 0 4417 37 4563 3 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 0 3703 42 3905 3 FreeSans 300 0 0 0 vcc_io
port 12 nsew
flabel metal1 s 0 3177 42 3379 3 FreeSans 300 0 0 0 vgnd_io
port 11 nsew
flabel metal1 s 66 3629 103 3675 3 FreeSans 300 180 0 0 slow_h_n
port 13 nsew
flabel metal1 s 13704 4223 13743 4244 0 FreeSans 200 0 0 0 pd_h<4>
port 2 nsew
flabel metal1 s 14655 4638 14695 4676 0 FreeSans 200 0 0 0 i2c_mode_h_n
port 3 nsew
flabel locali s 7603 3567 7653 3601 3 FreeSans 300 0 0 0 puen_h<0>
port 14 nsew
flabel locali s 8183 3556 8233 3590 3 FreeSans 300 0 0 0 pden_h_n<0>
port 15 nsew
flabel metal2 s 10324 3623 10382 3675 3 FreeSans 300 0 0 0 pd_h<3>
port 16 nsew
flabel metal2 s 9855 1940 9902 1992 3 FreeSans 300 180 0 0 pd_h<2>
port 17 nsew
flabel metal2 s 12176 3463 12223 3515 3 FreeSans 300 180 0 0 drvlo_h_n
port 18 nsew
flabel metal2 s 6875 3535 6927 3587 3 FreeSans 300 0 0 0 drvhi_h
port 19 nsew
flabel metal2 s 10160 3543 10207 3595 3 FreeSans 300 180 0 0 puen_h<1>
port 20 nsew
flabel metal2 s 9456 4009 9508 4061 3 FreeSans 300 0 0 0 pden_h_n<1>
port 21 nsew
<< properties >>
string GDS_END 88078116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88002672
string path 229.700 49.500 229.700 43.625 
<< end >>
