magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 2566 1426
<< nmos >>
rect 0 0 36 1400
rect 238 0 274 1400
rect 554 0 590 1400
rect 792 0 828 1400
rect 1108 0 1144 1400
rect 1346 0 1382 1400
rect 1662 0 1698 1400
rect 1900 0 1936 1400
rect 2216 0 2252 1400
rect 2454 0 2490 1400
<< ndiff >>
rect -50 0 0 1400
rect 36 0 238 1400
rect 274 0 314 1400
rect 514 0 554 1400
rect 590 0 792 1400
rect 828 0 868 1400
rect 1068 0 1108 1400
rect 1144 0 1346 1400
rect 1382 0 1422 1400
rect 1622 0 1662 1400
rect 1698 0 1900 1400
rect 1936 0 1976 1400
rect 2176 0 2216 1400
rect 2252 0 2454 1400
rect 2490 0 2540 1400
<< poly >>
rect 0 1400 36 1432
rect 238 1400 274 1432
rect 554 1400 590 1432
rect 792 1400 828 1432
rect 1108 1400 1144 1432
rect 1346 1400 1382 1432
rect 1662 1400 1698 1432
rect 1900 1400 1936 1432
rect 2216 1400 2252 1432
rect 2454 1400 2490 1432
rect 0 -32 36 0
rect 238 -32 274 0
rect 554 -32 590 0
rect 792 -32 828 0
rect 1108 -32 1144 0
rect 1346 -32 1382 0
rect 1662 -32 1698 0
rect 1900 -32 1936 0
rect 2216 -32 2252 0
rect 2454 -32 2490 0
<< locali >>
rect -229 -4 -51 1354
rect 325 -4 503 1354
rect 879 -4 1057 1354
rect 1433 -4 1611 1354
rect 1987 -4 2165 1354
rect 2541 -4 2719 1354
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_0
timestamp 1707688321
transform -1 0 -40 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_1
timestamp 1707688321
transform 1 0 314 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_2
timestamp 1707688321
transform 1 0 868 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_3
timestamp 1707688321
transform 1 0 1422 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_4
timestamp 1707688321
transform 1 0 1976 0 1 0
box -26 -26 226 1426
use DFTPL1s2_CDNS_55959141808702  DFTPL1s2_CDNS_55959141808702_5
timestamp 1707688321
transform 1 0 2530 0 1 0
box -26 -26 226 1426
<< labels >>
flabel comment s 2630 675 2630 675 0 FreeSans 300 0 0 0 S
flabel comment s 2353 700 2353 700 0 FreeSans 300 0 0 0 D
flabel comment s 2076 675 2076 675 0 FreeSans 300 0 0 0 S
flabel comment s 1799 700 1799 700 0 FreeSans 300 0 0 0 D
flabel comment s 1522 675 1522 675 0 FreeSans 300 0 0 0 S
flabel comment s 1245 700 1245 700 0 FreeSans 300 0 0 0 D
flabel comment s 968 675 968 675 0 FreeSans 300 0 0 0 S
flabel comment s 691 700 691 700 0 FreeSans 300 0 0 0 D
flabel comment s 414 675 414 675 0 FreeSans 300 0 0 0 S
flabel comment s 137 700 137 700 0 FreeSans 300 0 0 0 D
flabel comment s -140 675 -140 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 2760200
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2754832
<< end >>
