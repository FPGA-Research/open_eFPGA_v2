magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -79 -26 483 226
<< nmos >>
rect 0 0 36 200
rect 92 0 128 200
rect 184 0 220 200
rect 276 0 312 200
rect 368 0 404 200
<< ndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 36 182 92 200
rect 36 148 47 182
rect 81 148 92 182
rect 36 114 92 148
rect 36 80 47 114
rect 81 80 92 114
rect 36 46 92 80
rect 36 12 47 46
rect 81 12 92 46
rect 36 0 92 12
rect 128 182 184 200
rect 128 148 139 182
rect 173 148 184 182
rect 128 114 184 148
rect 128 80 139 114
rect 173 80 184 114
rect 128 46 184 80
rect 128 12 139 46
rect 173 12 184 46
rect 128 0 184 12
rect 220 182 276 200
rect 220 148 231 182
rect 265 148 276 182
rect 220 114 276 148
rect 220 80 231 114
rect 265 80 276 114
rect 220 46 276 80
rect 220 12 231 46
rect 265 12 276 46
rect 220 0 276 12
rect 312 182 368 200
rect 312 148 323 182
rect 357 148 368 182
rect 312 114 368 148
rect 312 80 323 114
rect 357 80 368 114
rect 312 46 368 80
rect 312 12 323 46
rect 357 12 368 46
rect 312 0 368 12
rect 404 182 457 200
rect 404 148 415 182
rect 449 148 457 182
rect 404 114 457 148
rect 404 80 415 114
rect 449 80 457 114
rect 404 46 457 80
rect 404 12 415 46
rect 449 12 457 46
rect 404 0 457 12
<< ndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 47 148 81 182
rect 47 80 81 114
rect 47 12 81 46
rect 139 148 173 182
rect 139 80 173 114
rect 139 12 173 46
rect 231 148 265 182
rect 231 80 265 114
rect 231 12 265 46
rect 323 148 357 182
rect 323 80 357 114
rect 323 12 357 46
rect 415 148 449 182
rect 415 80 449 114
rect 415 12 449 46
<< poly >>
rect 0 200 36 226
rect 92 200 128 226
rect 184 200 220 226
rect 276 200 312 226
rect 368 200 404 226
rect 0 -26 36 0
rect 92 -26 128 0
rect 184 -26 220 0
rect 276 -26 312 0
rect 368 -26 404 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 47 182 81 198
rect 47 114 81 148
rect 47 46 81 80
rect 47 -4 81 12
rect 139 182 173 198
rect 139 114 173 148
rect 139 46 173 80
rect 139 -4 173 12
rect 231 182 265 198
rect 231 114 265 148
rect 231 46 265 80
rect 231 -4 265 12
rect 323 182 357 198
rect 323 114 357 148
rect 323 46 357 80
rect 323 -4 357 12
rect 415 182 449 198
rect 415 114 449 148
rect 415 46 449 80
rect 415 -4 449 12
use DFL1sd2_CDNS_5246887918539  DFL1sd2_CDNS_5246887918539_0
timestamp 1707688321
transform 1 0 312 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_5246887918539  DFL1sd2_CDNS_5246887918539_1
timestamp 1707688321
transform 1 0 220 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_5246887918539  DFL1sd2_CDNS_5246887918539_2
timestamp 1707688321
transform 1 0 128 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_5246887918539  DFL1sd2_CDNS_5246887918539_3
timestamp 1707688321
transform 1 0 36 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_1
timestamp 1707688321
transform 1 0 404 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 64 97 64 97 0 FreeSans 300 0 0 0 D
flabel comment s 156 97 156 97 0 FreeSans 300 0 0 0 S
flabel comment s 248 97 248 97 0 FreeSans 300 0 0 0 D
flabel comment s 340 97 340 97 0 FreeSans 300 0 0 0 S
flabel comment s 432 97 432 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85797274
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85794468
<< end >>
