magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 679 1592 1471
<< pwell >>
rect 1420 25 1522 159
<< psubdiff >>
rect 1446 109 1496 133
rect 1446 75 1454 109
rect 1488 75 1496 109
rect 1446 51 1496 75
<< nsubdiff >>
rect 1446 1339 1496 1363
rect 1446 1305 1454 1339
rect 1488 1305 1496 1339
rect 1446 1281 1496 1305
<< psubdiffcont >>
rect 1454 75 1488 109
<< nsubdiffcont >>
rect 1454 1305 1488 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1556 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1350 1130 1384 1397
rect 1454 1339 1488 1397
rect 1454 1289 1488 1305
rect 64 724 98 740
rect 64 674 98 690
rect 706 724 740 1096
rect 706 690 757 724
rect 706 318 740 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1350 17 1384 218
rect 1454 109 1488 125
rect 1454 17 1488 75
rect 0 -17 1556 17
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_16  sky130_sram_1kbyte_1rw1r_32x256_8_contact_16_0
timestamp 1707688321
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_28  sky130_sram_1kbyte_1rw1r_32x256_8_contact_28_0
timestamp 1707688321
transform 1 0 1446 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_29  sky130_sram_1kbyte_1rw1r_32x256_8_contact_29_0
timestamp 1707688321
transform 1 0 1446 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m12_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m12_w2_000_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 51
box -26 -26 1364 456
use sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m12_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m12_w2_000_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 963
box -59 -56 1397 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 740 707 740 707 4 Z
rlabel locali s 778 0 778 0 4 gnd
rlabel locali s 778 1414 778 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1556 1414
string GDS_END 352868
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 350230
<< end >>
