magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect -2289 -120 5161 1874
<< nwell >>
rect -2369 1595 5241 1954
rect -2369 160 -2009 1595
rect -2369 -200 5241 160
rect 7513 -200 8129 1209
<< pwell >>
rect -1949 1448 5169 1534
rect -1949 306 -1863 1448
rect -1949 220 5169 306
<< mvpsubdiff >>
rect -1923 1474 -1833 1508
rect -1799 1474 -1765 1508
rect -1731 1474 -1697 1508
rect -1663 1474 -1629 1508
rect -1595 1474 -1485 1508
rect -1451 1474 -1417 1508
rect -1383 1474 -1349 1508
rect -1315 1474 -1281 1508
rect -1247 1474 -1213 1508
rect -1179 1474 -1145 1508
rect -1111 1474 -1077 1508
rect -1043 1474 -1009 1508
rect -975 1474 -941 1508
rect -907 1474 -873 1508
rect -839 1474 -805 1508
rect -771 1474 -737 1508
rect -703 1474 -669 1508
rect -635 1474 -601 1508
rect -567 1474 -533 1508
rect -499 1474 -465 1508
rect -431 1474 -397 1508
rect -363 1474 -329 1508
rect -295 1474 -261 1508
rect -227 1474 -193 1508
rect -159 1474 -125 1508
rect -91 1474 -57 1508
rect -23 1474 11 1508
rect 45 1474 79 1508
rect 113 1474 147 1508
rect 181 1474 215 1508
rect 249 1474 283 1508
rect 317 1474 351 1508
rect 385 1474 419 1508
rect 453 1474 487 1508
rect 521 1474 555 1508
rect 589 1474 623 1508
rect 657 1474 691 1508
rect 725 1474 759 1508
rect 793 1474 827 1508
rect 861 1474 895 1508
rect 929 1474 963 1508
rect 997 1474 1031 1508
rect 1065 1474 1099 1508
rect 1133 1474 1167 1508
rect 1201 1474 1235 1508
rect 1269 1474 1303 1508
rect 1337 1474 1371 1508
rect 1405 1474 1439 1508
rect 1473 1474 1507 1508
rect 1541 1474 1575 1508
rect 1609 1474 1643 1508
rect 1677 1474 1711 1508
rect 1745 1474 1779 1508
rect 1813 1474 1847 1508
rect 1881 1474 1915 1508
rect 1949 1474 1983 1508
rect 2017 1474 2051 1508
rect 2085 1474 2119 1508
rect 2153 1474 2187 1508
rect 2221 1474 2255 1508
rect 2289 1474 2323 1508
rect 2357 1474 2391 1508
rect 2425 1474 2459 1508
rect 2493 1474 2527 1508
rect 2561 1474 2595 1508
rect 2629 1474 2663 1508
rect 2697 1474 2731 1508
rect 2765 1474 2799 1508
rect 2833 1474 2867 1508
rect 2901 1474 2935 1508
rect 2969 1474 3003 1508
rect 3037 1474 3071 1508
rect 3105 1474 3139 1508
rect 3173 1474 3239 1508
rect 3273 1474 3307 1508
rect 3341 1474 3375 1508
rect 3409 1474 3443 1508
rect 3477 1474 3511 1508
rect 3545 1474 3579 1508
rect 3613 1474 3647 1508
rect 3681 1474 3715 1508
rect 3749 1474 3783 1508
rect 3817 1474 3851 1508
rect 3885 1474 3919 1508
rect 3953 1474 3987 1508
rect 4021 1474 4055 1508
rect 4089 1474 4123 1508
rect 4157 1474 4191 1508
rect 4225 1474 4259 1508
rect 4293 1474 4327 1508
rect 4361 1474 4395 1508
rect 4429 1474 4463 1508
rect 4497 1474 4531 1508
rect 4565 1474 4599 1508
rect 4633 1474 4667 1508
rect 4701 1474 4735 1508
rect 4769 1474 4803 1508
rect 4837 1474 4871 1508
rect 4905 1474 4939 1508
rect 4973 1474 5007 1508
rect 5041 1474 5075 1508
rect 5109 1474 5143 1508
rect -1923 1406 -1889 1440
rect -1923 1338 -1889 1372
rect -1923 1270 -1889 1304
rect -1923 1202 -1889 1236
rect -1923 1134 -1889 1168
rect -1923 1066 -1889 1100
rect -1923 998 -1889 1032
rect -1923 930 -1889 964
rect -1923 862 -1889 896
rect -1923 794 -1889 828
rect -1923 726 -1889 760
rect -1923 658 -1889 692
rect -1923 590 -1889 624
rect -1923 522 -1889 556
rect -1923 454 -1889 488
rect -1923 386 -1889 420
rect -1923 246 -1889 352
rect -1855 246 -1821 280
rect -1787 246 -1753 280
rect -1719 246 -1685 280
rect -1651 246 -1617 280
rect -1583 246 -1549 280
rect -1515 246 -1481 280
rect -1447 246 -1413 280
rect -1379 246 -1345 280
rect -1311 246 -1277 280
rect -1243 246 -1209 280
rect -1175 246 -1141 280
rect -1107 246 -1073 280
rect -1039 246 -1005 280
rect -971 246 -937 280
rect -903 246 -869 280
rect -835 246 -801 280
rect -767 246 -733 280
rect -699 246 -665 280
rect -631 246 -597 280
rect -563 246 -529 280
rect -495 246 -461 280
rect -427 246 -393 280
rect -359 246 -325 280
rect -291 246 -257 280
rect -223 246 -189 280
rect -155 246 -121 280
rect -87 246 -53 280
rect -19 246 15 280
rect 49 246 83 280
rect 117 246 151 280
rect 185 246 219 280
rect 253 246 287 280
rect 321 246 355 280
rect 389 246 423 280
rect 457 246 491 280
rect 525 246 559 280
rect 593 246 627 280
rect 661 246 695 280
rect 729 246 763 280
rect 797 246 831 280
rect 865 246 899 280
rect 933 246 967 280
rect 1001 246 1035 280
rect 1069 246 1103 280
rect 1137 246 1171 280
rect 1205 246 1239 280
rect 1273 246 1307 280
rect 1341 246 1375 280
rect 1409 246 1443 280
rect 1477 246 1511 280
rect 1545 246 1579 280
rect 1613 246 1647 280
rect 1681 246 1715 280
rect 1749 246 1783 280
rect 1817 246 1851 280
rect 1885 246 1919 280
rect 1953 246 1987 280
rect 2021 246 2055 280
rect 2089 246 2123 280
rect 2157 246 2191 280
rect 2225 246 2259 280
rect 2293 246 2327 280
rect 2361 246 2395 280
rect 2429 246 2463 280
rect 2497 246 2531 280
rect 2565 246 2599 280
rect 2633 246 2667 280
rect 2701 246 2735 280
rect 2769 246 2803 280
rect 2837 246 2871 280
rect 2905 246 2939 280
rect 2973 246 3007 280
rect 3041 246 3075 280
rect 3109 246 3143 280
rect 3177 246 3211 280
rect 3245 246 3279 280
rect 3313 246 3347 280
rect 3381 246 3415 280
rect 3449 246 3483 280
rect 3517 246 3551 280
rect 3585 246 3619 280
rect 3653 246 3687 280
rect 3721 246 3755 280
rect 3789 246 3823 280
rect 3857 246 3891 280
rect 3925 246 3959 280
rect 3993 246 4027 280
rect 4061 246 4095 280
rect 4129 246 4163 280
rect 4197 246 4231 280
rect 4265 246 4299 280
rect 4333 246 4367 280
rect 4401 246 4435 280
rect 4469 246 4503 280
rect 4537 246 4571 280
rect 4605 246 4639 280
rect 4673 246 4707 280
rect 4741 246 4775 280
rect 4809 246 4843 280
rect 4877 246 4911 280
rect 4945 246 4979 280
rect 5013 246 5047 280
rect 5081 246 5143 280
<< mvnsubdiff >>
rect -2303 1831 5070 1865
rect -2303 1797 -2279 1831
rect -2245 1797 -2210 1831
rect -2176 1797 -2141 1831
rect -2107 1797 -2072 1831
rect -2038 1797 -2003 1831
rect -1969 1797 -1934 1831
rect -1900 1797 -1865 1831
rect -1831 1797 -1796 1831
rect -1762 1797 -1727 1831
rect -1693 1797 -1658 1831
rect -1624 1797 -1589 1831
rect -1555 1797 -1520 1831
rect -1486 1797 -1451 1831
rect -1417 1797 -1382 1831
rect -1348 1797 -1313 1831
rect -1279 1797 -1244 1831
rect -2303 1763 -1244 1797
rect -2303 1729 -2279 1763
rect -2245 1729 -2210 1763
rect -2176 1729 -2141 1763
rect -2107 1729 -2072 1763
rect -2038 1729 -2003 1763
rect -1969 1729 -1934 1763
rect -1900 1729 -1865 1763
rect -1831 1729 -1796 1763
rect -1762 1729 -1727 1763
rect -1693 1729 -1658 1763
rect -1624 1729 -1589 1763
rect -1555 1729 -1520 1763
rect -1486 1729 -1451 1763
rect -1417 1729 -1382 1763
rect -1348 1729 -1313 1763
rect -1279 1729 -1244 1763
rect -2303 1695 -1244 1729
rect -2303 1661 -2279 1695
rect -2245 1661 -2210 1695
rect -2176 1661 -2141 1695
rect -2107 1661 -2072 1695
rect -2038 1661 -2003 1695
rect -1969 1661 -1934 1695
rect -1900 1661 -1865 1695
rect -1831 1661 -1796 1695
rect -1762 1661 -1727 1695
rect -1693 1661 -1658 1695
rect -1624 1661 -1589 1695
rect -1555 1661 -1520 1695
rect -1486 1661 -1451 1695
rect -1417 1661 -1382 1695
rect -1348 1661 -1313 1695
rect -1279 1661 -1244 1695
rect 5046 1661 5070 1831
rect -2303 1627 -2075 1661
rect -2303 1595 -2109 1627
rect -2303 1561 -2206 1595
rect -2172 1593 -2109 1595
rect -2172 1561 -2075 1593
rect -2303 1558 -2075 1561
rect -2303 1527 -2109 1558
rect -2303 1493 -2206 1527
rect -2172 1524 -2109 1527
rect -2172 1493 -2075 1524
rect -2303 1489 -2075 1493
rect -2303 1459 -2109 1489
rect -2303 1425 -2206 1459
rect -2172 1455 -2109 1459
rect -2172 1425 -2075 1455
rect -2303 1420 -2075 1425
rect -2303 1391 -2109 1420
rect -2303 1357 -2206 1391
rect -2172 1386 -2109 1391
rect -2172 1357 -2075 1386
rect -2303 1351 -2075 1357
rect -2303 1323 -2109 1351
rect -2303 1289 -2206 1323
rect -2172 1317 -2109 1323
rect -2172 1289 -2075 1317
rect -2303 1281 -2075 1289
rect -2303 1255 -2109 1281
rect -2303 1221 -2206 1255
rect -2172 1247 -2109 1255
rect -2172 1221 -2075 1247
rect -2303 1211 -2075 1221
rect -2303 1187 -2109 1211
rect -2303 1153 -2206 1187
rect -2172 1177 -2109 1187
rect -2172 1153 -2075 1177
rect -2303 1141 -2075 1153
rect -2303 1119 -2109 1141
rect -2303 1085 -2206 1119
rect -2172 1107 -2109 1119
rect -2172 1085 -2075 1107
rect -2303 1071 -2075 1085
rect -2303 1051 -2109 1071
rect -2303 1017 -2206 1051
rect -2172 1037 -2109 1051
rect -2172 1017 -2075 1037
rect -2303 1001 -2075 1017
rect -2303 983 -2109 1001
rect -2303 949 -2206 983
rect -2172 967 -2109 983
rect -2172 949 -2075 967
rect -2303 931 -2075 949
rect -2303 915 -2109 931
rect -2303 881 -2206 915
rect -2172 897 -2109 915
rect -2172 881 -2075 897
rect -2303 861 -2075 881
rect -2303 847 -2109 861
rect -2303 813 -2206 847
rect -2172 827 -2109 847
rect -2172 813 -2075 827
rect -2303 791 -2075 813
rect -2303 779 -2109 791
rect -2303 745 -2206 779
rect -2172 757 -2109 779
rect -2172 745 -2075 757
rect -2303 721 -2075 745
rect -2303 711 -2109 721
rect -2303 677 -2206 711
rect -2172 687 -2109 711
rect -2172 677 -2075 687
rect -2303 651 -2075 677
rect -2303 643 -2109 651
rect -2303 609 -2206 643
rect -2172 617 -2109 643
rect -2172 609 -2075 617
rect -2303 581 -2075 609
rect -2303 575 -2109 581
rect -2303 541 -2206 575
rect -2172 547 -2109 575
rect -2172 541 -2075 547
rect -2303 511 -2075 541
rect -2303 507 -2109 511
rect -2303 473 -2206 507
rect -2172 477 -2109 507
rect -2172 473 -2075 477
rect -2303 441 -2075 473
rect -2303 439 -2109 441
rect -2303 405 -2206 439
rect -2172 407 -2109 439
rect -2172 405 -2075 407
rect -2303 371 -2075 405
rect -2303 337 -2206 371
rect -2172 337 -2109 371
rect -2303 303 -2075 337
rect -2303 269 -2206 303
rect -2172 301 -2075 303
rect -2172 269 -2109 301
rect -2303 267 -2109 269
rect -2303 235 -2075 267
rect 7580 1023 7614 1142
rect 7648 1108 7682 1142
rect 7716 1108 7750 1142
rect 7784 1108 7858 1142
rect 7892 1108 7926 1142
rect 7960 1108 7994 1142
rect 7580 955 7614 989
rect 8028 1023 8062 1142
rect 7580 887 7614 921
rect 7580 819 7614 853
rect 7580 751 7614 785
rect 7580 683 7614 717
rect 7580 615 7614 649
rect 7580 547 7614 581
rect 7580 479 7614 513
rect 7580 411 7614 445
rect 7580 343 7614 377
rect 7580 275 7614 309
rect -2303 201 -2206 235
rect -2172 231 -2075 235
rect -2172 201 -2109 231
rect -2303 197 -2109 201
rect -2303 167 -2075 197
rect -2303 133 -2206 167
rect -2172 161 -2075 167
rect -2172 133 -2109 161
rect -2303 127 -2109 133
rect -2303 99 -2075 127
rect -2303 65 -2206 99
rect -2172 94 -2075 99
rect 7580 207 7614 241
rect 7580 139 7614 173
rect -2172 91 -1985 94
rect -2172 65 -2109 91
rect -2303 57 -2109 65
rect -2075 60 -1985 91
rect -1951 60 -1916 94
rect -1882 60 -1847 94
rect -1813 60 -1778 94
rect -1744 60 -1709 94
rect -1675 60 -1640 94
rect -1606 60 -1571 94
rect -1537 60 -1502 94
rect -1468 60 -1433 94
rect -1399 60 -1364 94
rect -1330 60 -1295 94
rect -1261 60 -1226 94
rect -1192 60 -1158 94
rect -1124 60 -1090 94
rect -1056 60 -1022 94
rect -988 60 -954 94
rect -920 60 -886 94
rect -852 60 -818 94
rect -784 60 -750 94
rect -716 60 -682 94
rect -648 60 -614 94
rect -580 60 -546 94
rect -512 60 -478 94
rect -444 60 -410 94
rect -376 60 -342 94
rect -308 60 -274 94
rect -240 60 -206 94
rect -172 60 -138 94
rect -104 60 -70 94
rect -36 60 -2 94
rect 32 60 66 94
rect 100 60 134 94
rect 168 60 202 94
rect 236 60 270 94
rect 304 60 338 94
rect 372 60 406 94
rect 440 60 474 94
rect 508 60 542 94
rect 576 60 610 94
rect 644 60 678 94
rect 712 60 746 94
rect 780 60 814 94
rect 848 60 882 94
rect 916 60 950 94
rect 984 60 1018 94
rect 1052 60 1086 94
rect 1120 60 1154 94
rect 1188 60 1222 94
rect 1256 60 1290 94
rect 1324 60 1358 94
rect 1392 60 1426 94
rect 1460 60 1494 94
rect 1528 60 1562 94
rect 1596 60 1630 94
rect 1664 60 1698 94
rect 1732 60 1766 94
rect 1800 60 1834 94
rect 1868 60 1902 94
rect 1936 60 1970 94
rect 2004 60 2038 94
rect 2072 60 2106 94
rect 2140 60 2174 94
rect 2208 60 2242 94
rect 2276 60 2310 94
rect 2344 60 2378 94
rect 2412 60 2446 94
rect 2480 60 2514 94
rect 2548 60 2582 94
rect 2616 60 2650 94
rect 2684 60 2718 94
rect 2752 60 2786 94
rect 2820 60 2854 94
rect 2888 60 2922 94
rect 2956 60 2990 94
rect 3024 60 3058 94
rect 3092 60 3126 94
rect 3160 60 3194 94
rect 3228 60 3262 94
rect 3296 60 3330 94
rect 3364 60 3398 94
rect 3432 60 3466 94
rect 3500 60 3534 94
rect 3568 60 3602 94
rect 3636 60 3670 94
rect 3704 60 3738 94
rect 3772 60 3806 94
rect 3840 60 3874 94
rect 3908 60 3942 94
rect 3976 60 4010 94
rect 4044 60 4078 94
rect 4112 60 4146 94
rect 4180 60 4214 94
rect 4248 60 4282 94
rect 4316 60 4350 94
rect 4384 60 4418 94
rect 4452 60 4486 94
rect 4520 60 4554 94
rect 4588 60 4622 94
rect 4656 60 4690 94
rect 4724 60 4758 94
rect 4792 60 4826 94
rect 4860 60 4894 94
rect 4928 60 4962 94
rect 4996 60 5030 94
rect 5064 60 5088 94
rect -2075 57 5088 60
rect -2303 31 5088 57
rect -2303 -3 -2206 31
rect -2172 21 5088 31
rect -2172 -3 -2109 21
rect -2303 -13 -2109 -3
rect -2075 -3 5088 21
rect -2075 -13 -1975 -3
rect -2303 -37 -1975 -13
rect -1941 -37 -1907 -3
rect -1873 -37 -1839 -3
rect -1805 -37 -1771 -3
rect -1737 -37 -1703 -3
rect -1669 -37 -1635 -3
rect -1601 -37 -1567 -3
rect -1533 -37 -1499 -3
rect -1465 -37 -1431 -3
rect -1397 -37 -1363 -3
rect -1329 -37 -1295 -3
rect -1261 -37 -1227 -3
rect -1193 -37 -1159 -3
rect -1125 -37 -1091 -3
rect -1057 -37 -1023 -3
rect -989 -37 -955 -3
rect -921 -37 -887 -3
rect -853 -37 -819 -3
rect -785 -37 -751 -3
rect -717 -37 -683 -3
rect -649 -37 -615 -3
rect -581 -37 -547 -3
rect -513 -37 -479 -3
rect -445 -37 -411 -3
rect -377 -37 -343 -3
rect -309 -37 -275 -3
rect -241 -37 -207 -3
rect -173 -37 -139 -3
rect -105 -37 -71 -3
rect -37 -37 -3 -3
rect 31 -37 65 -3
rect 99 -37 133 -3
rect 167 -37 201 -3
rect 235 -37 269 -3
rect 303 -37 337 -3
rect 371 -37 405 -3
rect 439 -37 473 -3
rect 507 -37 541 -3
rect 575 -37 609 -3
rect 643 -37 677 -3
rect 711 -37 745 -3
rect 779 -37 813 -3
rect 847 -37 881 -3
rect 915 -37 949 -3
rect 983 -37 1017 -3
rect 1051 -37 1085 -3
rect 1119 -37 1153 -3
rect 1187 -37 1221 -3
rect 1255 -37 1289 -3
rect 1323 -37 1357 -3
rect 1391 -37 1425 -3
rect 1459 -37 1493 -3
rect 1527 -37 1561 -3
rect 1595 -37 1629 -3
rect 1663 -37 1697 -3
rect 1731 -37 1765 -3
rect 1799 -37 1833 -3
rect 1867 -37 1901 -3
rect 1935 -37 1969 -3
rect 2003 -37 2037 -3
rect 2071 -37 2105 -3
rect 2139 -37 2173 -3
rect 2207 -37 2241 -3
rect 2275 -37 2309 -3
rect 2343 -37 2377 -3
rect 2411 -37 2445 -3
rect 2479 -37 2513 -3
rect 2547 -37 2581 -3
rect 2615 -37 2649 -3
rect 2683 -37 2717 -3
rect 2751 -37 2785 -3
rect 2819 -37 2853 -3
rect 2887 -37 2921 -3
rect 2955 -37 2989 -3
rect 3023 -37 3057 -3
rect 3091 -37 3125 -3
rect 3159 -37 3193 -3
rect 3227 -37 3261 -3
rect 3295 -37 3329 -3
rect 3363 -37 3397 -3
rect 3431 -37 3465 -3
rect 3499 -37 3533 -3
rect 3567 -37 3601 -3
rect 3635 -37 3669 -3
rect 3703 -37 3737 -3
rect 3771 -37 3805 -3
rect 3839 -37 3873 -3
rect 3907 -37 3941 -3
rect 3975 -37 4009 -3
rect 4043 -37 4077 -3
rect 4111 -37 4145 -3
rect 4179 -37 4213 -3
rect 4247 -37 4281 -3
rect 4315 -37 4349 -3
rect 4383 -37 4417 -3
rect 4451 -37 4485 -3
rect 4519 -37 4553 -3
rect 4587 -37 4621 -3
rect 4655 -37 4689 -3
rect 4723 -37 4757 -3
rect 4791 -37 4825 -3
rect 4859 -37 4893 -3
rect 4927 -37 4961 -3
rect 4995 -37 5088 -3
rect 7580 71 7614 105
rect 7580 3 7614 37
rect 7580 -65 7614 -31
rect 8028 955 8062 989
rect 8028 887 8062 921
rect 8028 819 8062 853
rect 8028 751 8062 785
rect 8028 683 8062 717
rect 8028 615 8062 649
rect 8028 547 8062 581
rect 8028 479 8062 513
rect 8028 411 8062 445
rect 8028 343 8062 377
rect 8028 275 8062 309
rect 8028 207 8062 241
rect 8028 139 8062 173
rect 8028 71 8062 105
rect 8028 3 8062 37
rect 8028 -65 8062 -31
rect 7580 -133 7708 -99
rect 7742 -133 7776 -99
rect 7810 -133 7878 -99
rect 7912 -133 7946 -99
rect 7980 -133 8062 -99
<< mvpsubdiffcont >>
rect -1833 1474 -1799 1508
rect -1765 1474 -1731 1508
rect -1697 1474 -1663 1508
rect -1629 1474 -1595 1508
rect -1485 1474 -1451 1508
rect -1417 1474 -1383 1508
rect -1349 1474 -1315 1508
rect -1281 1474 -1247 1508
rect -1213 1474 -1179 1508
rect -1145 1474 -1111 1508
rect -1077 1474 -1043 1508
rect -1009 1474 -975 1508
rect -941 1474 -907 1508
rect -873 1474 -839 1508
rect -805 1474 -771 1508
rect -737 1474 -703 1508
rect -669 1474 -635 1508
rect -601 1474 -567 1508
rect -533 1474 -499 1508
rect -465 1474 -431 1508
rect -397 1474 -363 1508
rect -329 1474 -295 1508
rect -261 1474 -227 1508
rect -193 1474 -159 1508
rect -125 1474 -91 1508
rect -57 1474 -23 1508
rect 11 1474 45 1508
rect 79 1474 113 1508
rect 147 1474 181 1508
rect 215 1474 249 1508
rect 283 1474 317 1508
rect 351 1474 385 1508
rect 419 1474 453 1508
rect 487 1474 521 1508
rect 555 1474 589 1508
rect 623 1474 657 1508
rect 691 1474 725 1508
rect 759 1474 793 1508
rect 827 1474 861 1508
rect 895 1474 929 1508
rect 963 1474 997 1508
rect 1031 1474 1065 1508
rect 1099 1474 1133 1508
rect 1167 1474 1201 1508
rect 1235 1474 1269 1508
rect 1303 1474 1337 1508
rect 1371 1474 1405 1508
rect 1439 1474 1473 1508
rect 1507 1474 1541 1508
rect 1575 1474 1609 1508
rect 1643 1474 1677 1508
rect 1711 1474 1745 1508
rect 1779 1474 1813 1508
rect 1847 1474 1881 1508
rect 1915 1474 1949 1508
rect 1983 1474 2017 1508
rect 2051 1474 2085 1508
rect 2119 1474 2153 1508
rect 2187 1474 2221 1508
rect 2255 1474 2289 1508
rect 2323 1474 2357 1508
rect 2391 1474 2425 1508
rect 2459 1474 2493 1508
rect 2527 1474 2561 1508
rect 2595 1474 2629 1508
rect 2663 1474 2697 1508
rect 2731 1474 2765 1508
rect 2799 1474 2833 1508
rect 2867 1474 2901 1508
rect 2935 1474 2969 1508
rect 3003 1474 3037 1508
rect 3071 1474 3105 1508
rect 3139 1474 3173 1508
rect 3239 1474 3273 1508
rect 3307 1474 3341 1508
rect 3375 1474 3409 1508
rect 3443 1474 3477 1508
rect 3511 1474 3545 1508
rect 3579 1474 3613 1508
rect 3647 1474 3681 1508
rect 3715 1474 3749 1508
rect 3783 1474 3817 1508
rect 3851 1474 3885 1508
rect 3919 1474 3953 1508
rect 3987 1474 4021 1508
rect 4055 1474 4089 1508
rect 4123 1474 4157 1508
rect 4191 1474 4225 1508
rect 4259 1474 4293 1508
rect 4327 1474 4361 1508
rect 4395 1474 4429 1508
rect 4463 1474 4497 1508
rect 4531 1474 4565 1508
rect 4599 1474 4633 1508
rect 4667 1474 4701 1508
rect 4735 1474 4769 1508
rect 4803 1474 4837 1508
rect 4871 1474 4905 1508
rect 4939 1474 4973 1508
rect 5007 1474 5041 1508
rect 5075 1474 5109 1508
rect -1923 1440 -1889 1474
rect -1923 1372 -1889 1406
rect -1923 1304 -1889 1338
rect -1923 1236 -1889 1270
rect -1923 1168 -1889 1202
rect -1923 1100 -1889 1134
rect -1923 1032 -1889 1066
rect -1923 964 -1889 998
rect -1923 896 -1889 930
rect -1923 828 -1889 862
rect -1923 760 -1889 794
rect -1923 692 -1889 726
rect -1923 624 -1889 658
rect -1923 556 -1889 590
rect -1923 488 -1889 522
rect -1923 420 -1889 454
rect -1923 352 -1889 386
rect -1889 246 -1855 280
rect -1821 246 -1787 280
rect -1753 246 -1719 280
rect -1685 246 -1651 280
rect -1617 246 -1583 280
rect -1549 246 -1515 280
rect -1481 246 -1447 280
rect -1413 246 -1379 280
rect -1345 246 -1311 280
rect -1277 246 -1243 280
rect -1209 246 -1175 280
rect -1141 246 -1107 280
rect -1073 246 -1039 280
rect -1005 246 -971 280
rect -937 246 -903 280
rect -869 246 -835 280
rect -801 246 -767 280
rect -733 246 -699 280
rect -665 246 -631 280
rect -597 246 -563 280
rect -529 246 -495 280
rect -461 246 -427 280
rect -393 246 -359 280
rect -325 246 -291 280
rect -257 246 -223 280
rect -189 246 -155 280
rect -121 246 -87 280
rect -53 246 -19 280
rect 15 246 49 280
rect 83 246 117 280
rect 151 246 185 280
rect 219 246 253 280
rect 287 246 321 280
rect 355 246 389 280
rect 423 246 457 280
rect 491 246 525 280
rect 559 246 593 280
rect 627 246 661 280
rect 695 246 729 280
rect 763 246 797 280
rect 831 246 865 280
rect 899 246 933 280
rect 967 246 1001 280
rect 1035 246 1069 280
rect 1103 246 1137 280
rect 1171 246 1205 280
rect 1239 246 1273 280
rect 1307 246 1341 280
rect 1375 246 1409 280
rect 1443 246 1477 280
rect 1511 246 1545 280
rect 1579 246 1613 280
rect 1647 246 1681 280
rect 1715 246 1749 280
rect 1783 246 1817 280
rect 1851 246 1885 280
rect 1919 246 1953 280
rect 1987 246 2021 280
rect 2055 246 2089 280
rect 2123 246 2157 280
rect 2191 246 2225 280
rect 2259 246 2293 280
rect 2327 246 2361 280
rect 2395 246 2429 280
rect 2463 246 2497 280
rect 2531 246 2565 280
rect 2599 246 2633 280
rect 2667 246 2701 280
rect 2735 246 2769 280
rect 2803 246 2837 280
rect 2871 246 2905 280
rect 2939 246 2973 280
rect 3007 246 3041 280
rect 3075 246 3109 280
rect 3143 246 3177 280
rect 3211 246 3245 280
rect 3279 246 3313 280
rect 3347 246 3381 280
rect 3415 246 3449 280
rect 3483 246 3517 280
rect 3551 246 3585 280
rect 3619 246 3653 280
rect 3687 246 3721 280
rect 3755 246 3789 280
rect 3823 246 3857 280
rect 3891 246 3925 280
rect 3959 246 3993 280
rect 4027 246 4061 280
rect 4095 246 4129 280
rect 4163 246 4197 280
rect 4231 246 4265 280
rect 4299 246 4333 280
rect 4367 246 4401 280
rect 4435 246 4469 280
rect 4503 246 4537 280
rect 4571 246 4605 280
rect 4639 246 4673 280
rect 4707 246 4741 280
rect 4775 246 4809 280
rect 4843 246 4877 280
rect 4911 246 4945 280
rect 4979 246 5013 280
rect 5047 246 5081 280
<< mvnsubdiffcont >>
rect -2279 1797 -2245 1831
rect -2210 1797 -2176 1831
rect -2141 1797 -2107 1831
rect -2072 1797 -2038 1831
rect -2003 1797 -1969 1831
rect -1934 1797 -1900 1831
rect -1865 1797 -1831 1831
rect -1796 1797 -1762 1831
rect -1727 1797 -1693 1831
rect -1658 1797 -1624 1831
rect -1589 1797 -1555 1831
rect -1520 1797 -1486 1831
rect -1451 1797 -1417 1831
rect -1382 1797 -1348 1831
rect -1313 1797 -1279 1831
rect -2279 1729 -2245 1763
rect -2210 1729 -2176 1763
rect -2141 1729 -2107 1763
rect -2072 1729 -2038 1763
rect -2003 1729 -1969 1763
rect -1934 1729 -1900 1763
rect -1865 1729 -1831 1763
rect -1796 1729 -1762 1763
rect -1727 1729 -1693 1763
rect -1658 1729 -1624 1763
rect -1589 1729 -1555 1763
rect -1520 1729 -1486 1763
rect -1451 1729 -1417 1763
rect -1382 1729 -1348 1763
rect -1313 1729 -1279 1763
rect -2279 1661 -2245 1695
rect -2210 1661 -2176 1695
rect -2141 1661 -2107 1695
rect -2072 1661 -2038 1695
rect -2003 1661 -1969 1695
rect -1934 1661 -1900 1695
rect -1865 1661 -1831 1695
rect -1796 1661 -1762 1695
rect -1727 1661 -1693 1695
rect -1658 1661 -1624 1695
rect -1589 1661 -1555 1695
rect -1520 1661 -1486 1695
rect -1451 1661 -1417 1695
rect -1382 1661 -1348 1695
rect -1313 1661 -1279 1695
rect -1244 1661 5046 1831
rect -2206 1561 -2172 1595
rect -2109 1593 -2075 1627
rect -2206 1493 -2172 1527
rect -2109 1524 -2075 1558
rect -2206 1425 -2172 1459
rect -2109 1455 -2075 1489
rect -2206 1357 -2172 1391
rect -2109 1386 -2075 1420
rect -2206 1289 -2172 1323
rect -2109 1317 -2075 1351
rect -2206 1221 -2172 1255
rect -2109 1247 -2075 1281
rect -2206 1153 -2172 1187
rect -2109 1177 -2075 1211
rect -2206 1085 -2172 1119
rect -2109 1107 -2075 1141
rect -2206 1017 -2172 1051
rect -2109 1037 -2075 1071
rect -2206 949 -2172 983
rect -2109 967 -2075 1001
rect -2206 881 -2172 915
rect -2109 897 -2075 931
rect -2206 813 -2172 847
rect -2109 827 -2075 861
rect -2206 745 -2172 779
rect -2109 757 -2075 791
rect -2206 677 -2172 711
rect -2109 687 -2075 721
rect -2206 609 -2172 643
rect -2109 617 -2075 651
rect -2206 541 -2172 575
rect -2109 547 -2075 581
rect -2206 473 -2172 507
rect -2109 477 -2075 511
rect -2206 405 -2172 439
rect -2109 407 -2075 441
rect -2206 337 -2172 371
rect -2109 337 -2075 371
rect -2206 269 -2172 303
rect -2109 267 -2075 301
rect 7614 1108 7648 1142
rect 7682 1108 7716 1142
rect 7750 1108 7784 1142
rect 7858 1108 7892 1142
rect 7926 1108 7960 1142
rect 7994 1108 8028 1142
rect 7580 989 7614 1023
rect 8028 989 8062 1023
rect 7580 921 7614 955
rect 7580 853 7614 887
rect 7580 785 7614 819
rect 7580 717 7614 751
rect 7580 649 7614 683
rect 7580 581 7614 615
rect 7580 513 7614 547
rect 7580 445 7614 479
rect 7580 377 7614 411
rect 7580 309 7614 343
rect -2206 201 -2172 235
rect -2109 197 -2075 231
rect -2206 133 -2172 167
rect -2109 127 -2075 161
rect -2206 65 -2172 99
rect 7580 241 7614 275
rect 7580 173 7614 207
rect 7580 105 7614 139
rect -2109 57 -2075 91
rect -1985 60 -1951 94
rect -1916 60 -1882 94
rect -1847 60 -1813 94
rect -1778 60 -1744 94
rect -1709 60 -1675 94
rect -1640 60 -1606 94
rect -1571 60 -1537 94
rect -1502 60 -1468 94
rect -1433 60 -1399 94
rect -1364 60 -1330 94
rect -1295 60 -1261 94
rect -1226 60 -1192 94
rect -1158 60 -1124 94
rect -1090 60 -1056 94
rect -1022 60 -988 94
rect -954 60 -920 94
rect -886 60 -852 94
rect -818 60 -784 94
rect -750 60 -716 94
rect -682 60 -648 94
rect -614 60 -580 94
rect -546 60 -512 94
rect -478 60 -444 94
rect -410 60 -376 94
rect -342 60 -308 94
rect -274 60 -240 94
rect -206 60 -172 94
rect -138 60 -104 94
rect -70 60 -36 94
rect -2 60 32 94
rect 66 60 100 94
rect 134 60 168 94
rect 202 60 236 94
rect 270 60 304 94
rect 338 60 372 94
rect 406 60 440 94
rect 474 60 508 94
rect 542 60 576 94
rect 610 60 644 94
rect 678 60 712 94
rect 746 60 780 94
rect 814 60 848 94
rect 882 60 916 94
rect 950 60 984 94
rect 1018 60 1052 94
rect 1086 60 1120 94
rect 1154 60 1188 94
rect 1222 60 1256 94
rect 1290 60 1324 94
rect 1358 60 1392 94
rect 1426 60 1460 94
rect 1494 60 1528 94
rect 1562 60 1596 94
rect 1630 60 1664 94
rect 1698 60 1732 94
rect 1766 60 1800 94
rect 1834 60 1868 94
rect 1902 60 1936 94
rect 1970 60 2004 94
rect 2038 60 2072 94
rect 2106 60 2140 94
rect 2174 60 2208 94
rect 2242 60 2276 94
rect 2310 60 2344 94
rect 2378 60 2412 94
rect 2446 60 2480 94
rect 2514 60 2548 94
rect 2582 60 2616 94
rect 2650 60 2684 94
rect 2718 60 2752 94
rect 2786 60 2820 94
rect 2854 60 2888 94
rect 2922 60 2956 94
rect 2990 60 3024 94
rect 3058 60 3092 94
rect 3126 60 3160 94
rect 3194 60 3228 94
rect 3262 60 3296 94
rect 3330 60 3364 94
rect 3398 60 3432 94
rect 3466 60 3500 94
rect 3534 60 3568 94
rect 3602 60 3636 94
rect 3670 60 3704 94
rect 3738 60 3772 94
rect 3806 60 3840 94
rect 3874 60 3908 94
rect 3942 60 3976 94
rect 4010 60 4044 94
rect 4078 60 4112 94
rect 4146 60 4180 94
rect 4214 60 4248 94
rect 4282 60 4316 94
rect 4350 60 4384 94
rect 4418 60 4452 94
rect 4486 60 4520 94
rect 4554 60 4588 94
rect 4622 60 4656 94
rect 4690 60 4724 94
rect 4758 60 4792 94
rect 4826 60 4860 94
rect 4894 60 4928 94
rect 4962 60 4996 94
rect 5030 60 5064 94
rect -2206 -3 -2172 31
rect -2109 -13 -2075 21
rect -1975 -37 -1941 -3
rect -1907 -37 -1873 -3
rect -1839 -37 -1805 -3
rect -1771 -37 -1737 -3
rect -1703 -37 -1669 -3
rect -1635 -37 -1601 -3
rect -1567 -37 -1533 -3
rect -1499 -37 -1465 -3
rect -1431 -37 -1397 -3
rect -1363 -37 -1329 -3
rect -1295 -37 -1261 -3
rect -1227 -37 -1193 -3
rect -1159 -37 -1125 -3
rect -1091 -37 -1057 -3
rect -1023 -37 -989 -3
rect -955 -37 -921 -3
rect -887 -37 -853 -3
rect -819 -37 -785 -3
rect -751 -37 -717 -3
rect -683 -37 -649 -3
rect -615 -37 -581 -3
rect -547 -37 -513 -3
rect -479 -37 -445 -3
rect -411 -37 -377 -3
rect -343 -37 -309 -3
rect -275 -37 -241 -3
rect -207 -37 -173 -3
rect -139 -37 -105 -3
rect -71 -37 -37 -3
rect -3 -37 31 -3
rect 65 -37 99 -3
rect 133 -37 167 -3
rect 201 -37 235 -3
rect 269 -37 303 -3
rect 337 -37 371 -3
rect 405 -37 439 -3
rect 473 -37 507 -3
rect 541 -37 575 -3
rect 609 -37 643 -3
rect 677 -37 711 -3
rect 745 -37 779 -3
rect 813 -37 847 -3
rect 881 -37 915 -3
rect 949 -37 983 -3
rect 1017 -37 1051 -3
rect 1085 -37 1119 -3
rect 1153 -37 1187 -3
rect 1221 -37 1255 -3
rect 1289 -37 1323 -3
rect 1357 -37 1391 -3
rect 1425 -37 1459 -3
rect 1493 -37 1527 -3
rect 1561 -37 1595 -3
rect 1629 -37 1663 -3
rect 1697 -37 1731 -3
rect 1765 -37 1799 -3
rect 1833 -37 1867 -3
rect 1901 -37 1935 -3
rect 1969 -37 2003 -3
rect 2037 -37 2071 -3
rect 2105 -37 2139 -3
rect 2173 -37 2207 -3
rect 2241 -37 2275 -3
rect 2309 -37 2343 -3
rect 2377 -37 2411 -3
rect 2445 -37 2479 -3
rect 2513 -37 2547 -3
rect 2581 -37 2615 -3
rect 2649 -37 2683 -3
rect 2717 -37 2751 -3
rect 2785 -37 2819 -3
rect 2853 -37 2887 -3
rect 2921 -37 2955 -3
rect 2989 -37 3023 -3
rect 3057 -37 3091 -3
rect 3125 -37 3159 -3
rect 3193 -37 3227 -3
rect 3261 -37 3295 -3
rect 3329 -37 3363 -3
rect 3397 -37 3431 -3
rect 3465 -37 3499 -3
rect 3533 -37 3567 -3
rect 3601 -37 3635 -3
rect 3669 -37 3703 -3
rect 3737 -37 3771 -3
rect 3805 -37 3839 -3
rect 3873 -37 3907 -3
rect 3941 -37 3975 -3
rect 4009 -37 4043 -3
rect 4077 -37 4111 -3
rect 4145 -37 4179 -3
rect 4213 -37 4247 -3
rect 4281 -37 4315 -3
rect 4349 -37 4383 -3
rect 4417 -37 4451 -3
rect 4485 -37 4519 -3
rect 4553 -37 4587 -3
rect 4621 -37 4655 -3
rect 4689 -37 4723 -3
rect 4757 -37 4791 -3
rect 4825 -37 4859 -3
rect 4893 -37 4927 -3
rect 4961 -37 4995 -3
rect 7580 37 7614 71
rect 7580 -31 7614 3
rect 7580 -99 7614 -65
rect 8028 921 8062 955
rect 8028 853 8062 887
rect 8028 785 8062 819
rect 8028 717 8062 751
rect 8028 649 8062 683
rect 8028 581 8062 615
rect 8028 513 8062 547
rect 8028 445 8062 479
rect 8028 377 8062 411
rect 8028 309 8062 343
rect 8028 241 8062 275
rect 8028 173 8062 207
rect 8028 105 8062 139
rect 8028 37 8062 71
rect 8028 -31 8062 3
rect 8028 -99 8062 -65
rect 7708 -133 7742 -99
rect 7776 -133 7810 -99
rect 7878 -133 7912 -99
rect 7946 -133 7980 -99
<< poly >>
rect -1762 1426 -1562 1442
rect -1762 1392 -1722 1426
rect -1688 1392 -1626 1426
rect -1592 1392 -1562 1426
rect -1762 1380 -1562 1392
rect -1506 1426 -1306 1442
rect -1506 1392 -1466 1426
rect -1432 1392 -1370 1426
rect -1336 1392 -1306 1426
rect -1506 1380 -1306 1392
rect -1250 1426 -1050 1442
rect -1250 1392 -1210 1426
rect -1176 1392 -1114 1426
rect -1080 1392 -1050 1426
rect -1250 1380 -1050 1392
rect -994 1426 -794 1442
rect -994 1392 -954 1426
rect -920 1392 -858 1426
rect -824 1392 -794 1426
rect -994 1380 -794 1392
rect -738 1426 -538 1442
rect -738 1392 -698 1426
rect -664 1392 -602 1426
rect -568 1392 -538 1426
rect -738 1380 -538 1392
rect -482 1426 -282 1442
rect -482 1392 -442 1426
rect -408 1392 -346 1426
rect -312 1392 -282 1426
rect -482 1380 -282 1392
rect -226 1426 -26 1442
rect -226 1392 -186 1426
rect -152 1392 -90 1426
rect -56 1392 -26 1426
rect -226 1380 -26 1392
rect 30 1426 230 1442
rect 30 1392 70 1426
rect 104 1392 166 1426
rect 200 1392 230 1426
rect 30 1380 230 1392
rect 286 1426 486 1442
rect 286 1392 326 1426
rect 360 1392 422 1426
rect 456 1392 486 1426
rect 286 1380 486 1392
rect 542 1426 742 1442
rect 542 1392 582 1426
rect 616 1392 678 1426
rect 712 1392 742 1426
rect 542 1380 742 1392
rect 798 1426 998 1442
rect 798 1392 838 1426
rect 872 1392 934 1426
rect 968 1392 998 1426
rect 798 1380 998 1392
rect 1054 1426 1254 1442
rect 1054 1392 1094 1426
rect 1128 1392 1190 1426
rect 1224 1392 1254 1426
rect 1054 1380 1254 1392
rect 1310 1426 1510 1442
rect 1310 1392 1350 1426
rect 1384 1392 1446 1426
rect 1480 1392 1510 1426
rect 1310 1380 1510 1392
rect 1566 1426 1766 1442
rect 1566 1392 1606 1426
rect 1640 1392 1702 1426
rect 1736 1392 1766 1426
rect 1566 1380 1766 1392
rect 1822 1426 2022 1442
rect 1822 1392 1862 1426
rect 1896 1392 1958 1426
rect 1992 1392 2022 1426
rect 1822 1380 2022 1392
rect 2078 1426 2278 1442
rect 2078 1392 2118 1426
rect 2152 1392 2214 1426
rect 2248 1392 2278 1426
rect 2078 1380 2278 1392
rect 2334 1426 2534 1442
rect 2334 1392 2374 1426
rect 2408 1392 2470 1426
rect 2504 1392 2534 1426
rect 2334 1380 2534 1392
rect 2590 1426 2790 1442
rect 2590 1392 2630 1426
rect 2664 1392 2726 1426
rect 2760 1392 2790 1426
rect 2590 1380 2790 1392
rect 2846 1426 3046 1442
rect 2846 1392 2886 1426
rect 2920 1392 2982 1426
rect 3016 1392 3046 1426
rect 2846 1380 3046 1392
rect 3102 1426 3302 1442
rect 3102 1392 3142 1426
rect 3176 1392 3238 1426
rect 3272 1392 3302 1426
rect 3102 1380 3302 1392
rect 3358 1426 3558 1442
rect 3358 1392 3398 1426
rect 3432 1392 3494 1426
rect 3528 1392 3558 1426
rect 3358 1380 3558 1392
rect 3614 1426 3814 1442
rect 3614 1392 3654 1426
rect 3688 1392 3750 1426
rect 3784 1392 3814 1426
rect 3614 1380 3814 1392
rect 3870 1426 4070 1442
rect 3870 1392 3910 1426
rect 3944 1392 4006 1426
rect 4040 1392 4070 1426
rect 3870 1380 4070 1392
rect 4126 1426 4326 1442
rect 4126 1392 4166 1426
rect 4200 1392 4262 1426
rect 4296 1392 4326 1426
rect 4126 1380 4326 1392
rect 4492 1426 5060 1442
rect 4492 1392 4508 1426
rect 4542 1392 4580 1426
rect 4614 1392 4652 1426
rect 4686 1392 4724 1426
rect 4758 1392 4796 1426
rect 4830 1392 4868 1426
rect 4902 1392 4939 1426
rect 4973 1392 5010 1426
rect 5044 1392 5060 1426
rect -1738 1376 -1576 1380
rect -1482 1376 -1320 1380
rect -1226 1376 -1064 1380
rect -970 1376 -808 1380
rect -714 1376 -552 1380
rect -458 1376 -296 1380
rect -202 1376 -40 1380
rect 54 1376 216 1380
rect 310 1376 472 1380
rect 566 1376 728 1380
rect 822 1376 984 1380
rect 1078 1376 1240 1380
rect 1334 1376 1496 1380
rect 1590 1376 1752 1380
rect 1846 1376 2008 1380
rect 2102 1376 2264 1380
rect 2358 1376 2520 1380
rect 2614 1376 2776 1380
rect 2870 1376 3032 1380
rect 3126 1376 3288 1380
rect 3382 1376 3544 1380
rect 3638 1376 3800 1380
rect 3894 1376 4056 1380
rect 4150 1376 4312 1380
rect 4492 1376 5060 1392
rect 7721 1037 7921 1054
rect 7721 1003 7751 1037
rect 7785 1003 7847 1037
rect 7881 1003 7921 1037
rect 7721 980 7921 1003
<< polycont >>
rect -1722 1392 -1688 1426
rect -1626 1392 -1592 1426
rect -1466 1392 -1432 1426
rect -1370 1392 -1336 1426
rect -1210 1392 -1176 1426
rect -1114 1392 -1080 1426
rect -954 1392 -920 1426
rect -858 1392 -824 1426
rect -698 1392 -664 1426
rect -602 1392 -568 1426
rect -442 1392 -408 1426
rect -346 1392 -312 1426
rect -186 1392 -152 1426
rect -90 1392 -56 1426
rect 70 1392 104 1426
rect 166 1392 200 1426
rect 326 1392 360 1426
rect 422 1392 456 1426
rect 582 1392 616 1426
rect 678 1392 712 1426
rect 838 1392 872 1426
rect 934 1392 968 1426
rect 1094 1392 1128 1426
rect 1190 1392 1224 1426
rect 1350 1392 1384 1426
rect 1446 1392 1480 1426
rect 1606 1392 1640 1426
rect 1702 1392 1736 1426
rect 1862 1392 1896 1426
rect 1958 1392 1992 1426
rect 2118 1392 2152 1426
rect 2214 1392 2248 1426
rect 2374 1392 2408 1426
rect 2470 1392 2504 1426
rect 2630 1392 2664 1426
rect 2726 1392 2760 1426
rect 2886 1392 2920 1426
rect 2982 1392 3016 1426
rect 3142 1392 3176 1426
rect 3238 1392 3272 1426
rect 3398 1392 3432 1426
rect 3494 1392 3528 1426
rect 3654 1392 3688 1426
rect 3750 1392 3784 1426
rect 3910 1392 3944 1426
rect 4006 1392 4040 1426
rect 4166 1392 4200 1426
rect 4262 1392 4296 1426
rect 4508 1392 4542 1426
rect 4580 1392 4614 1426
rect 4652 1392 4686 1426
rect 4724 1392 4758 1426
rect 4796 1392 4830 1426
rect 4868 1392 4902 1426
rect 4939 1392 4973 1426
rect 5010 1392 5044 1426
rect 7751 1003 7785 1037
rect 7847 1003 7881 1037
<< locali >>
rect -2303 1831 5070 1865
rect -2303 1797 -2279 1831
rect -2245 1797 -2210 1831
rect -2176 1797 -2141 1831
rect -2107 1814 -2072 1831
rect -2038 1814 -2003 1831
rect -1969 1814 -1934 1831
rect -1900 1814 -1865 1831
rect -1831 1814 -1796 1831
rect -1762 1814 -1727 1831
rect -1693 1814 -1658 1831
rect -1624 1814 -1589 1831
rect -1555 1814 -1520 1831
rect -1486 1814 -1451 1831
rect -1417 1814 -1382 1831
rect -1348 1814 -1313 1831
rect -1279 1814 -1244 1831
rect -2303 1763 -2127 1797
rect -2303 1729 -2279 1763
rect -2245 1729 -2210 1763
rect -2176 1729 -2141 1763
rect -2303 1708 -2127 1729
rect -2303 1695 -1244 1708
rect -2303 1661 -2279 1695
rect -2245 1661 -2210 1695
rect -2176 1661 -2141 1695
rect -2107 1661 -2072 1695
rect -2038 1661 -2003 1695
rect -1969 1661 -1934 1695
rect -1900 1661 -1865 1695
rect -1831 1661 -1796 1695
rect -1762 1661 -1727 1695
rect -1693 1661 -1658 1695
rect -1624 1661 -1589 1695
rect -1555 1661 -1520 1695
rect -1486 1661 -1451 1695
rect -1417 1661 -1382 1695
rect -1348 1661 -1313 1695
rect -1279 1661 -1244 1695
rect 5046 1661 5070 1831
rect -2303 1627 -2045 1661
rect -2303 1595 -2109 1627
rect -2303 1576 -2206 1595
rect -2303 1542 -2243 1576
rect -2209 1561 -2206 1576
rect -2172 1593 -2109 1595
rect -2075 1593 -2045 1627
rect -1676 1593 -1638 1627
rect -2172 1576 -2045 1593
rect -2172 1561 -2171 1576
rect -2209 1542 -2171 1561
rect -2137 1558 -2045 1576
rect -2137 1542 -2109 1558
rect -2303 1527 -2109 1542
rect -2303 1493 -2206 1527
rect -2172 1524 -2109 1527
rect -2075 1524 -2045 1558
rect 4988 1548 5026 1582
rect -2172 1493 -2045 1524
rect -2303 1489 -2045 1493
rect -2303 1459 -2109 1489
rect -2303 1425 -2206 1459
rect -2172 1455 -2109 1459
rect -2075 1455 -2045 1489
rect -2172 1425 -2045 1455
rect -2303 1420 -2045 1425
rect -2303 1391 -2109 1420
rect -2303 1357 -2206 1391
rect -2172 1386 -2109 1391
rect -2075 1386 -2045 1420
rect -2172 1357 -2045 1386
rect -2303 1351 -2045 1357
rect -2303 1323 -2109 1351
rect -2303 1289 -2206 1323
rect -2172 1317 -2109 1323
rect -2075 1317 -2045 1351
rect -2172 1289 -2045 1317
rect -2303 1281 -2045 1289
rect -2303 1255 -2109 1281
rect -2303 1254 -2206 1255
rect -2303 1220 -2243 1254
rect -2209 1221 -2206 1254
rect -2172 1254 -2109 1255
rect -2172 1221 -2171 1254
rect -2209 1220 -2171 1221
rect -2137 1247 -2109 1254
rect -2075 1247 -2045 1281
rect -2137 1220 -2045 1247
rect -2303 1211 -2045 1220
rect -2303 1187 -2109 1211
rect -2303 1181 -2206 1187
rect -2303 1147 -2243 1181
rect -2209 1153 -2206 1181
rect -2172 1181 -2109 1187
rect -2172 1153 -2171 1181
rect -2209 1147 -2171 1153
rect -2137 1177 -2109 1181
rect -2075 1177 -2045 1211
rect -2137 1147 -2045 1177
rect -2303 1141 -2045 1147
rect -2303 1119 -2109 1141
rect -2303 1108 -2206 1119
rect -2303 1074 -2243 1108
rect -2209 1085 -2206 1108
rect -2172 1108 -2109 1119
rect -2172 1085 -2171 1108
rect -2209 1074 -2171 1085
rect -2137 1107 -2109 1108
rect -2075 1107 -2045 1141
rect -2137 1074 -2045 1107
rect -2303 1071 -2045 1074
rect -2303 1051 -2109 1071
rect -2303 1035 -2206 1051
rect -2303 1001 -2243 1035
rect -2209 1017 -2206 1035
rect -2172 1037 -2109 1051
rect -2075 1037 -2045 1071
rect -2172 1035 -2045 1037
rect -2172 1017 -2171 1035
rect -2209 1001 -2171 1017
rect -2137 1001 -2045 1035
rect -2303 983 -2109 1001
rect -2303 962 -2206 983
rect -2303 928 -2243 962
rect -2209 949 -2206 962
rect -2172 967 -2109 983
rect -2075 967 -2045 1001
rect -2172 962 -2045 967
rect -2172 949 -2171 962
rect -2209 928 -2171 949
rect -2137 931 -2045 962
rect -2137 928 -2109 931
rect -2303 915 -2109 928
rect -2303 889 -2206 915
rect -2303 855 -2243 889
rect -2209 881 -2206 889
rect -2172 897 -2109 915
rect -2075 897 -2045 931
rect -2172 889 -2045 897
rect -2172 881 -2171 889
rect -2209 855 -2171 881
rect -2137 861 -2045 889
rect -2137 855 -2109 861
rect -2303 847 -2109 855
rect -2303 816 -2206 847
rect -2303 782 -2243 816
rect -2209 813 -2206 816
rect -2172 827 -2109 847
rect -2075 827 -2045 861
rect -2172 816 -2045 827
rect -2172 813 -2171 816
rect -2209 782 -2171 813
rect -2137 791 -2045 816
rect -2137 782 -2109 791
rect -2303 779 -2109 782
rect -2303 745 -2206 779
rect -2172 757 -2109 779
rect -2075 757 -2045 791
rect -2172 745 -2045 757
rect -2303 743 -2045 745
rect -2303 709 -2243 743
rect -2209 711 -2171 743
rect -2209 709 -2206 711
rect -2303 677 -2206 709
rect -2172 709 -2171 711
rect -2137 721 -2045 743
rect -2137 709 -2109 721
rect -2172 687 -2109 709
rect -2075 687 -2045 721
rect -2172 677 -2045 687
rect -2303 670 -2045 677
rect -2303 636 -2243 670
rect -2209 643 -2171 670
rect -2209 636 -2206 643
rect -2303 609 -2206 636
rect -2172 636 -2171 643
rect -2137 651 -2045 670
rect -2137 636 -2109 651
rect -2172 617 -2109 636
rect -2075 617 -2045 651
rect -2172 609 -2045 617
rect -2303 597 -2045 609
rect -2303 275 -2243 597
rect -2137 581 -2045 597
rect -2137 547 -2109 581
rect -2075 547 -2045 581
rect -2137 511 -2045 547
rect -2137 477 -2109 511
rect -2075 477 -2045 511
rect -2137 441 -2045 477
rect -2137 407 -2109 441
rect -2075 407 -2045 441
rect -2137 371 -2045 407
rect -2137 337 -2109 371
rect -2075 337 -2045 371
rect -2137 301 -2045 337
rect -2137 275 -2109 301
rect -2303 269 -2206 275
rect -2172 269 -2109 275
rect -2303 267 -2109 269
rect -2075 267 -2045 301
rect -2303 235 -2045 267
rect -1923 1474 -1843 1508
rect -1799 1474 -1765 1508
rect -1731 1474 -1697 1508
rect -1663 1474 -1629 1508
rect -1595 1474 -1519 1508
rect -1451 1474 -1447 1508
rect -1383 1474 -1375 1508
rect -1315 1474 -1303 1508
rect -1247 1474 -1231 1508
rect -1179 1474 -1159 1508
rect -1111 1474 -1087 1508
rect -1043 1474 -1015 1508
rect -975 1474 -943 1508
rect -907 1474 -873 1508
rect -837 1474 -805 1508
rect -765 1474 -737 1508
rect -693 1474 -669 1508
rect -621 1474 -601 1508
rect -549 1474 -533 1508
rect -477 1474 -465 1508
rect -405 1474 -397 1508
rect -333 1474 -329 1508
rect -227 1474 -223 1508
rect -159 1474 -151 1508
rect -91 1474 -79 1508
rect -23 1474 -7 1508
rect 45 1474 65 1508
rect 113 1474 137 1508
rect 181 1474 209 1508
rect 249 1474 281 1508
rect 317 1474 351 1508
rect 387 1474 419 1508
rect 459 1474 487 1508
rect 531 1474 555 1508
rect 603 1474 623 1508
rect 675 1474 691 1508
rect 747 1474 759 1508
rect 819 1474 827 1508
rect 891 1474 895 1508
rect 997 1474 1001 1508
rect 1065 1474 1073 1508
rect 1133 1474 1145 1508
rect 1201 1474 1217 1508
rect 1269 1474 1289 1508
rect 1337 1474 1361 1508
rect 1405 1474 1433 1508
rect 1473 1474 1505 1508
rect 1541 1474 1575 1508
rect 1611 1474 1643 1508
rect 1683 1474 1711 1508
rect 1755 1474 1779 1508
rect 1827 1474 1847 1508
rect 1899 1474 1915 1508
rect 1971 1474 1983 1508
rect 2043 1474 2051 1508
rect 2115 1474 2119 1508
rect 2221 1474 2225 1508
rect 2289 1474 2297 1508
rect 2357 1474 2369 1508
rect 2425 1474 2442 1508
rect 2493 1474 2515 1508
rect 2561 1474 2588 1508
rect 2629 1474 2661 1508
rect 2697 1474 2731 1508
rect 2768 1474 2799 1508
rect 2841 1474 2867 1508
rect 2914 1474 2935 1508
rect 2987 1474 3003 1508
rect 3060 1474 3071 1508
rect 3133 1474 3139 1508
rect 3206 1474 3239 1508
rect 3279 1474 3307 1508
rect 3352 1474 3375 1508
rect 3425 1474 3443 1508
rect 3498 1474 3511 1508
rect 3571 1474 3579 1508
rect 3644 1474 3647 1508
rect 3681 1474 3683 1508
rect 3749 1474 3756 1508
rect 3817 1474 3829 1508
rect 3885 1474 3902 1508
rect 3953 1474 3975 1508
rect 4021 1474 4048 1508
rect 4089 1474 4121 1508
rect 4157 1474 4191 1508
rect 4228 1474 4259 1508
rect 4301 1474 4327 1508
rect 4374 1474 4395 1508
rect 4447 1474 4463 1508
rect 4520 1474 4531 1508
rect 4593 1474 4599 1508
rect 4666 1474 4667 1508
rect 4701 1474 4705 1508
rect 4769 1474 4778 1508
rect 4837 1474 4851 1508
rect 4905 1474 4939 1508
rect 4973 1474 5007 1508
rect 5041 1474 5075 1508
rect 5109 1474 5143 1508
rect -1923 1406 -1889 1440
rect -1738 1392 -1722 1426
rect -1676 1392 -1638 1426
rect -1592 1392 -1576 1426
rect -1482 1392 -1466 1426
rect -1432 1392 -1370 1426
rect -1336 1392 -1320 1426
rect -1226 1392 -1210 1426
rect -1176 1392 -1114 1426
rect -1080 1392 -1064 1426
rect -970 1392 -954 1426
rect -920 1392 -858 1426
rect -824 1392 -808 1426
rect -714 1392 -698 1426
rect -664 1392 -602 1426
rect -568 1392 -552 1426
rect -458 1392 -442 1426
rect -408 1392 -346 1426
rect -312 1392 -296 1426
rect -202 1392 -186 1426
rect -152 1392 -90 1426
rect -56 1392 -40 1426
rect 54 1392 70 1426
rect 104 1392 166 1426
rect 200 1392 216 1426
rect 310 1392 326 1426
rect 360 1392 422 1426
rect 456 1392 472 1426
rect 566 1392 582 1426
rect 616 1392 678 1426
rect 712 1392 728 1426
rect 822 1392 838 1426
rect 872 1392 934 1426
rect 968 1392 984 1426
rect 1078 1392 1094 1426
rect 1128 1392 1190 1426
rect 1224 1392 1240 1426
rect 1334 1392 1350 1426
rect 1384 1392 1446 1426
rect 1480 1392 1496 1426
rect 1590 1392 1606 1426
rect 1640 1392 1702 1426
rect 1736 1392 1752 1426
rect 1846 1392 1862 1426
rect 1896 1392 1958 1426
rect 1992 1392 2008 1426
rect 2102 1392 2118 1426
rect 2152 1392 2214 1426
rect 2248 1392 2264 1426
rect 2358 1392 2374 1426
rect 2408 1392 2470 1426
rect 2504 1392 2520 1426
rect 2614 1392 2630 1426
rect 2664 1392 2726 1426
rect 2760 1392 2776 1426
rect 2870 1392 2886 1426
rect 2920 1392 2982 1426
rect 3016 1392 3032 1426
rect 3126 1392 3142 1426
rect 3176 1392 3238 1426
rect 3272 1392 3288 1426
rect 3382 1392 3398 1426
rect 3432 1392 3494 1426
rect 3528 1392 3544 1426
rect 3638 1392 3654 1426
rect 3688 1392 3750 1426
rect 3784 1392 3800 1426
rect 3894 1392 3910 1426
rect 3944 1392 4006 1426
rect 4040 1392 4056 1426
rect 4150 1392 4166 1426
rect 4200 1392 4262 1426
rect 4296 1392 4371 1426
rect -1923 1338 -1889 1372
rect -1458 1340 -1352 1392
rect -1424 1306 -1386 1340
rect -1202 1340 -1096 1392
rect -1168 1306 -1130 1340
rect -946 1340 -840 1392
rect -912 1306 -874 1340
rect -690 1340 -584 1392
rect -656 1306 -618 1340
rect -434 1340 -328 1392
rect -400 1306 -362 1340
rect -178 1340 -72 1392
rect -144 1306 -106 1340
rect 78 1340 184 1392
rect 112 1306 150 1340
rect 334 1340 440 1392
rect 368 1306 406 1340
rect 590 1340 696 1392
rect 624 1306 662 1340
rect 846 1340 952 1392
rect 880 1306 918 1340
rect 1102 1340 1208 1392
rect 1136 1306 1174 1340
rect 1358 1340 1464 1392
rect 1392 1306 1430 1340
rect 1614 1340 1720 1392
rect 1648 1306 1686 1340
rect 1870 1340 1976 1392
rect 1904 1306 1942 1340
rect 2126 1340 2232 1392
rect 2160 1306 2198 1340
rect 2382 1340 2488 1392
rect 2416 1306 2454 1340
rect 2638 1340 2744 1392
rect 2672 1306 2710 1340
rect 2894 1340 3000 1392
rect 2928 1306 2966 1340
rect 3150 1340 3256 1392
rect 3184 1306 3222 1340
rect 3406 1340 3512 1392
rect 3440 1306 3478 1340
rect 3662 1340 3768 1392
rect 3696 1306 3734 1340
rect 3918 1340 4024 1392
rect 3952 1306 3990 1340
rect -1923 1270 -1889 1304
rect 4337 1300 4371 1392
rect 4492 1392 4508 1426
rect 4542 1392 4580 1426
rect 4614 1392 4652 1426
rect 4686 1392 4724 1426
rect 4758 1392 4796 1426
rect 4830 1392 4868 1426
rect 4902 1392 4939 1426
rect 4988 1392 5010 1426
rect 4492 1334 5060 1392
rect -1923 1202 -1889 1236
rect 4515 1260 4569 1334
rect 4515 1226 4525 1260
rect 4559 1226 4569 1260
rect 4515 1220 4569 1226
rect 4671 1260 4725 1334
rect 4671 1226 4681 1260
rect 4715 1226 4725 1260
rect 4671 1220 4725 1226
rect 4827 1260 4881 1334
rect 4827 1226 4837 1260
rect 4871 1226 4881 1260
rect 4827 1220 4881 1226
rect 4983 1333 5060 1334
rect 4983 1260 5037 1333
rect 4983 1226 4993 1260
rect 5027 1226 5037 1260
rect 4983 1220 5037 1226
rect -1923 1134 -1889 1168
rect -1923 1066 -1889 1100
rect -1923 998 -1889 1032
rect -1923 930 -1889 964
rect 4759 1104 4793 1142
rect 4759 1032 4793 1070
rect -1923 862 -1889 896
rect 3313 889 3347 927
rect -1923 794 -1889 828
rect -1923 726 -1889 760
rect -1923 658 -1889 692
rect -1923 590 -1889 624
rect -1923 522 -1889 556
rect -1923 454 -1889 488
rect -1923 386 -1889 420
rect 2033 780 2067 818
rect 2033 708 2067 746
rect 2033 636 2067 674
rect 2033 564 2067 602
rect 2033 492 2067 530
rect 2033 420 2067 458
rect 3057 780 3091 818
rect 3057 708 3091 746
rect 3057 636 3091 674
rect 3057 564 3091 602
rect 3057 492 3091 530
rect 3313 817 3347 855
rect 3313 745 3347 783
rect 3313 673 3347 711
rect 3313 601 3347 639
rect 3313 529 3347 567
rect 3825 889 3859 927
rect 3825 817 3859 855
rect 3825 745 3859 783
rect 3825 673 3859 711
rect 4759 960 4793 998
rect 4759 888 4793 926
rect 4759 816 4793 854
rect 4759 744 4793 782
rect 7580 1139 7614 1142
rect 7648 1139 7682 1142
rect 7716 1139 7750 1142
rect 7784 1139 7858 1142
rect 7892 1139 7926 1142
rect 7960 1139 7994 1142
rect 8028 1139 8062 1142
rect 7580 1105 7586 1139
rect 7648 1108 7659 1139
rect 7716 1108 7732 1139
rect 7784 1108 7805 1139
rect 7620 1105 7659 1108
rect 7693 1105 7732 1108
rect 7766 1105 7805 1108
rect 7839 1108 7858 1139
rect 7912 1108 7926 1139
rect 7984 1108 7994 1139
rect 7839 1105 7878 1108
rect 7912 1105 7950 1108
rect 7984 1105 8022 1108
rect 8056 1105 8062 1139
rect 7580 1102 8062 1105
rect 7580 1023 7614 1102
rect 7735 1003 7751 1037
rect 7805 1003 7843 1037
rect 7881 1003 7897 1037
rect 8028 1023 8062 1102
rect 7580 955 7614 989
rect 7580 887 7614 921
rect 7580 819 7614 853
rect 7580 751 7614 785
rect 3825 601 3859 639
rect 3825 529 3859 567
rect 7580 683 7614 717
rect 7580 615 7614 649
rect 7580 547 7614 581
rect 3057 420 3091 458
rect 7580 479 7614 513
rect 7580 411 7614 445
rect -1923 280 -1889 352
rect 7580 343 7614 377
rect -1923 246 -1917 280
rect -1855 246 -1845 280
rect -1787 246 -1773 280
rect -1719 246 -1701 280
rect -1651 246 -1629 280
rect -1583 246 -1557 280
rect -1515 246 -1485 280
rect -1447 246 -1413 280
rect -1379 246 -1345 280
rect -1307 246 -1277 280
rect -1235 246 -1209 280
rect -1163 246 -1141 280
rect -1091 246 -1073 280
rect -1019 246 -1005 280
rect -947 246 -937 280
rect -875 246 -869 280
rect -803 246 -801 280
rect -767 246 -765 280
rect -699 246 -693 280
rect -631 246 -621 280
rect -563 246 -549 280
rect -495 246 -477 280
rect -427 246 -405 280
rect -359 246 -333 280
rect -291 246 -261 280
rect -223 246 -189 280
rect -155 246 -121 280
rect -83 246 -53 280
rect -11 246 15 280
rect 61 246 83 280
rect 133 246 151 280
rect 205 246 219 280
rect 277 246 287 280
rect 349 246 355 280
rect 421 246 423 280
rect 457 246 460 280
rect 525 246 533 280
rect 593 246 606 280
rect 661 246 679 280
rect 729 246 752 280
rect 797 246 825 280
rect 865 246 898 280
rect 933 246 967 280
rect 1005 246 1035 280
rect 1078 246 1103 280
rect 1151 246 1171 280
rect 1224 246 1239 280
rect 1297 246 1307 280
rect 1370 246 1375 280
rect 1477 246 1482 280
rect 1545 246 1555 280
rect 1613 246 1628 280
rect 1681 246 1701 280
rect 1749 246 1774 280
rect 1817 246 1847 280
rect 1885 246 1919 280
rect 1954 246 1987 280
rect 2027 246 2055 280
rect 2100 246 2123 280
rect 2173 246 2191 280
rect 2246 246 2259 280
rect 2319 246 2327 280
rect 2392 246 2395 280
rect 2429 246 2431 280
rect 2497 246 2504 280
rect 2565 246 2577 280
rect 2633 246 2650 280
rect 2701 246 2723 280
rect 2769 246 2796 280
rect 2837 246 2869 280
rect 2905 246 2939 280
rect 2976 246 3007 280
rect 3049 246 3075 280
rect 3122 246 3143 280
rect 3195 246 3211 280
rect 3268 246 3279 280
rect 3341 246 3347 280
rect 3414 246 3415 280
rect 3449 246 3453 280
rect 3517 246 3526 280
rect 3585 246 3599 280
rect 3653 246 3672 280
rect 3721 246 3745 280
rect 3789 246 3818 280
rect 3857 246 3891 280
rect 3925 246 3959 280
rect 3998 246 4027 280
rect 4071 246 4095 280
rect 4144 246 4163 280
rect 4217 246 4231 280
rect 4290 246 4299 280
rect 4363 246 4367 280
rect 4401 246 4402 280
rect 4469 246 4475 280
rect 4537 246 4548 280
rect 4605 246 4621 280
rect 4673 246 4694 280
rect 4741 246 4767 280
rect 4809 246 4840 280
rect 4877 246 4911 280
rect 4947 246 4979 280
rect 5020 246 5047 280
rect 5093 246 5143 280
rect 7580 275 7614 309
rect -2303 201 -2206 235
rect -2172 231 -2045 235
rect -2172 201 -2109 231
rect -2303 197 -2109 201
rect -2075 197 -2045 231
rect -2303 167 -2045 197
rect -2303 133 -2206 167
rect -2172 161 -2045 167
rect -2172 133 -2109 161
rect -2303 127 -2109 133
rect -2075 127 -2045 161
rect -2303 99 -2045 127
rect -2303 65 -2206 99
rect -2172 94 -2045 99
rect 7580 207 7614 241
rect 7580 139 7614 173
rect -2172 91 -1985 94
rect -2172 65 -2109 91
rect -2303 57 -2109 65
rect -2075 60 -1985 91
rect -1951 60 -1916 94
rect -1882 60 -1847 94
rect -1813 60 -1778 94
rect -1744 60 -1709 94
rect -1675 60 -1640 94
rect -1606 60 -1571 94
rect -1537 60 -1502 94
rect -1468 60 -1433 94
rect -1399 60 -1364 94
rect -1330 60 -1295 94
rect -1261 60 -1226 94
rect -1192 60 -1158 94
rect -1124 60 -1090 94
rect -1056 60 -1022 94
rect -988 60 -954 94
rect -920 60 -886 94
rect -852 60 -818 94
rect -784 60 -750 94
rect -716 60 -682 94
rect -648 60 -614 94
rect -580 60 -546 94
rect -512 60 -478 94
rect -444 60 -410 94
rect -376 60 -342 94
rect -308 60 -274 94
rect -240 60 -206 94
rect -172 60 -138 94
rect -104 60 -70 94
rect -36 60 -2 94
rect 32 60 66 94
rect 100 60 134 94
rect 168 60 202 94
rect 236 60 270 94
rect 304 60 338 94
rect 372 60 406 94
rect 440 60 474 94
rect 508 60 542 94
rect 576 60 610 94
rect 644 60 678 94
rect 712 60 746 94
rect 780 60 814 94
rect 848 60 882 94
rect 916 60 950 94
rect 984 60 1018 94
rect 1052 60 1086 94
rect 1120 60 1154 94
rect 1188 60 1222 94
rect 1256 60 1290 94
rect 1324 60 1358 94
rect 1392 60 1426 94
rect 1460 60 1494 94
rect 1528 60 1562 94
rect 1596 60 1630 94
rect 1664 60 1698 94
rect 1732 60 1766 94
rect 1800 60 1834 94
rect 1868 60 1902 94
rect 1936 60 1970 94
rect 2004 60 2038 94
rect 2072 60 2106 94
rect 2140 60 2174 94
rect 2208 60 2242 94
rect 2276 60 2310 94
rect 2344 60 2378 94
rect 2412 60 2446 94
rect 2480 60 2514 94
rect 2548 60 2582 94
rect 2616 60 2650 94
rect 2684 60 2718 94
rect 2752 60 2786 94
rect 2820 60 2854 94
rect 2888 60 2922 94
rect 2956 60 2990 94
rect 3024 60 3058 94
rect 3092 60 3126 94
rect 3160 60 3194 94
rect 3228 60 3262 94
rect 3296 60 3330 94
rect 3364 60 3398 94
rect 3432 60 3466 94
rect 3500 60 3534 94
rect 3568 60 3602 94
rect 3636 60 3670 94
rect 3704 60 3738 94
rect 3772 60 3806 94
rect 3840 60 3874 94
rect 3908 60 3942 94
rect 3976 60 4010 94
rect 4044 60 4078 94
rect 4112 60 4146 94
rect 4180 60 4214 94
rect 4248 60 4282 94
rect 4316 60 4350 94
rect 4384 60 4418 94
rect 4452 60 4486 94
rect 4520 60 4554 94
rect 4588 60 4622 94
rect 4656 60 4690 94
rect 4724 60 4758 94
rect 4792 60 4826 94
rect 4860 60 4894 94
rect 4928 60 4962 94
rect 4996 60 5030 94
rect 5064 60 5088 94
rect -2075 57 5088 60
rect -2303 31 5088 57
rect -2303 -3 -2206 31
rect -2172 21 5088 31
rect -2172 -3 -2109 21
rect -2075 -3 5088 21
rect -2303 -37 -2194 -3
rect -2160 -37 -2122 -3
rect -2075 -13 -2050 -3
rect -2088 -37 -2050 -13
rect -2016 -37 -1978 -3
rect -1941 -37 -1907 -3
rect -1872 -37 -1839 -3
rect -1800 -37 -1771 -3
rect -1728 -37 -1703 -3
rect -1656 -37 -1635 -3
rect -1584 -37 -1567 -3
rect -1512 -37 -1499 -3
rect -1440 -37 -1431 -3
rect -1368 -37 -1363 -3
rect -1296 -37 -1295 -3
rect -1261 -37 -1258 -3
rect -1193 -37 -1186 -3
rect -1125 -37 -1114 -3
rect -1057 -37 -1042 -3
rect -989 -37 -970 -3
rect -921 -37 -898 -3
rect -853 -37 -826 -3
rect -785 -37 -754 -3
rect -717 -37 -683 -3
rect -648 -37 -615 -3
rect -576 -37 -547 -3
rect -504 -37 -479 -3
rect -432 -37 -411 -3
rect -360 -37 -343 -3
rect -288 -37 -275 -3
rect -216 -37 -207 -3
rect -144 -37 -139 -3
rect -72 -37 -71 -3
rect -37 -37 -34 -3
rect 31 -37 38 -3
rect 99 -37 110 -3
rect 167 -37 182 -3
rect 235 -37 254 -3
rect 303 -37 326 -3
rect 371 -37 398 -3
rect 439 -37 470 -3
rect 507 -37 541 -3
rect 576 -37 609 -3
rect 648 -37 677 -3
rect 720 -37 745 -3
rect 792 -37 813 -3
rect 864 -37 881 -3
rect 936 -37 949 -3
rect 1008 -37 1017 -3
rect 1080 -37 1085 -3
rect 1152 -37 1153 -3
rect 1187 -37 1190 -3
rect 1255 -37 1262 -3
rect 1323 -37 1334 -3
rect 1391 -37 1406 -3
rect 1459 -37 1478 -3
rect 1527 -37 1550 -3
rect 1595 -37 1622 -3
rect 1663 -37 1694 -3
rect 1731 -37 1765 -3
rect 1800 -37 1833 -3
rect 1872 -37 1901 -3
rect 1944 -37 1969 -3
rect 2016 -37 2037 -3
rect 2088 -37 2105 -3
rect 2160 -37 2173 -3
rect 2232 -37 2241 -3
rect 2304 -37 2309 -3
rect 2411 -37 2416 -3
rect 2479 -37 2489 -3
rect 2547 -37 2562 -3
rect 2615 -37 2635 -3
rect 2683 -37 2708 -3
rect 2751 -37 2781 -3
rect 2819 -37 2853 -3
rect 2888 -37 2921 -3
rect 2961 -37 2989 -3
rect 3034 -37 3057 -3
rect 3107 -37 3125 -3
rect 3180 -37 3193 -3
rect 3253 -37 3261 -3
rect 3326 -37 3329 -3
rect 3363 -37 3365 -3
rect 3431 -37 3438 -3
rect 3499 -37 3511 -3
rect 3567 -37 3584 -3
rect 3635 -37 3657 -3
rect 3703 -37 3730 -3
rect 3771 -37 3803 -3
rect 3839 -37 3873 -3
rect 3910 -37 3941 -3
rect 3983 -37 4009 -3
rect 4056 -37 4077 -3
rect 4129 -37 4145 -3
rect 4202 -37 4213 -3
rect 4275 -37 4281 -3
rect 4348 -37 4349 -3
rect 4383 -37 4387 -3
rect 4451 -37 4460 -3
rect 4519 -37 4533 -3
rect 4587 -37 4606 -3
rect 4655 -37 4679 -3
rect 4723 -37 4752 -3
rect 4791 -37 4825 -3
rect 4859 -37 4893 -3
rect 4932 -37 4961 -3
rect 5005 -37 5088 -3
rect 7580 71 7614 105
rect 7580 3 7614 37
rect 7580 -65 7614 -31
rect 8028 955 8062 989
rect 8028 887 8062 921
rect 8028 819 8062 853
rect 8028 751 8062 785
rect 8028 683 8062 717
rect 8028 615 8062 649
rect 8028 547 8062 581
rect 8028 479 8062 513
rect 8028 411 8062 445
rect 8028 343 8062 377
rect 8028 275 8062 309
rect 8028 207 8062 241
rect 8028 139 8062 173
rect 8028 71 8062 105
rect 8028 3 8062 37
rect 8028 -65 8062 -31
rect 7580 -133 7586 -99
rect 7620 -133 7659 -99
rect 7693 -133 7708 -99
rect 7766 -133 7776 -99
rect 7839 -133 7878 -99
rect 7912 -133 7946 -99
rect 7984 -133 8022 -99
rect 8056 -133 8062 -99
<< viali >>
rect -2127 1797 -2107 1814
rect -2107 1797 -2072 1814
rect -2072 1797 -2038 1814
rect -2038 1797 -2003 1814
rect -2003 1797 -1969 1814
rect -1969 1797 -1934 1814
rect -1934 1797 -1900 1814
rect -1900 1797 -1865 1814
rect -1865 1797 -1831 1814
rect -1831 1797 -1796 1814
rect -1796 1797 -1762 1814
rect -1762 1797 -1727 1814
rect -1727 1797 -1693 1814
rect -1693 1797 -1658 1814
rect -1658 1797 -1624 1814
rect -1624 1797 -1589 1814
rect -1589 1797 -1555 1814
rect -1555 1797 -1520 1814
rect -1520 1797 -1486 1814
rect -1486 1797 -1451 1814
rect -1451 1797 -1417 1814
rect -1417 1797 -1382 1814
rect -1382 1797 -1348 1814
rect -1348 1797 -1313 1814
rect -1313 1797 -1279 1814
rect -1279 1797 -1244 1814
rect -2127 1763 -1244 1797
rect -2127 1729 -2107 1763
rect -2107 1729 -2072 1763
rect -2072 1729 -2038 1763
rect -2038 1729 -2003 1763
rect -2003 1729 -1969 1763
rect -1969 1729 -1934 1763
rect -1934 1729 -1900 1763
rect -1900 1729 -1865 1763
rect -1865 1729 -1831 1763
rect -1831 1729 -1796 1763
rect -1796 1729 -1762 1763
rect -1762 1729 -1727 1763
rect -1727 1729 -1693 1763
rect -1693 1729 -1658 1763
rect -1658 1729 -1624 1763
rect -1624 1729 -1589 1763
rect -1589 1729 -1555 1763
rect -1555 1729 -1520 1763
rect -1520 1729 -1486 1763
rect -1486 1729 -1451 1763
rect -1451 1729 -1417 1763
rect -1417 1729 -1382 1763
rect -1382 1729 -1348 1763
rect -1348 1729 -1313 1763
rect -1313 1729 -1279 1763
rect -1279 1729 -1244 1763
rect -2127 1708 -1244 1729
rect -1244 1708 787 1814
rect 826 1780 860 1814
rect 899 1780 933 1814
rect 972 1780 1006 1814
rect 1045 1780 1079 1814
rect 1118 1780 1152 1814
rect 1191 1780 1225 1814
rect 1264 1780 1298 1814
rect 1337 1780 1371 1814
rect 1410 1780 1444 1814
rect 1483 1780 1517 1814
rect 1556 1780 1590 1814
rect 1629 1780 1663 1814
rect 1702 1780 1736 1814
rect 1775 1780 1809 1814
rect 1848 1780 1882 1814
rect 1921 1780 1955 1814
rect 1994 1780 2028 1814
rect 2067 1780 2101 1814
rect 2140 1780 2174 1814
rect 2213 1780 2247 1814
rect 2286 1780 2320 1814
rect 2359 1780 2393 1814
rect 2432 1780 2466 1814
rect 2505 1780 2539 1814
rect 2578 1780 2612 1814
rect 2651 1780 2685 1814
rect 2724 1780 2758 1814
rect 2797 1780 2831 1814
rect 2870 1780 2904 1814
rect 2943 1780 2977 1814
rect 3016 1780 3050 1814
rect 3089 1780 3123 1814
rect 3162 1780 3196 1814
rect 3235 1780 3269 1814
rect 3308 1780 3342 1814
rect 3381 1780 3415 1814
rect 3454 1780 3488 1814
rect 3527 1780 3561 1814
rect 3600 1780 3634 1814
rect 3673 1780 3707 1814
rect 3746 1780 3780 1814
rect 3819 1780 3853 1814
rect 3892 1780 3926 1814
rect 3965 1780 3999 1814
rect 4038 1780 4072 1814
rect 4111 1780 4145 1814
rect 4184 1780 4218 1814
rect 4257 1780 4291 1814
rect 4330 1780 4364 1814
rect 4403 1780 4437 1814
rect 4476 1780 4510 1814
rect 4549 1780 4583 1814
rect 4622 1780 4656 1814
rect 4695 1780 4729 1814
rect 4768 1780 4802 1814
rect 4841 1780 4875 1814
rect 4914 1780 4948 1814
rect 4987 1780 5021 1814
rect 826 1708 860 1742
rect 899 1708 933 1742
rect 972 1708 1006 1742
rect 1045 1708 1079 1742
rect 1118 1708 1152 1742
rect 1191 1708 1225 1742
rect 1264 1708 1298 1742
rect 1337 1708 1371 1742
rect 1410 1708 1444 1742
rect 1483 1708 1517 1742
rect 1556 1708 1590 1742
rect 1629 1708 1663 1742
rect 1702 1708 1736 1742
rect 1775 1708 1809 1742
rect 1848 1708 1882 1742
rect 1921 1708 1955 1742
rect 1994 1708 2028 1742
rect 2067 1708 2101 1742
rect 2140 1708 2174 1742
rect 2213 1708 2247 1742
rect 2286 1708 2320 1742
rect 2359 1708 2393 1742
rect 2432 1708 2466 1742
rect 2505 1708 2539 1742
rect 2578 1708 2612 1742
rect 2651 1708 2685 1742
rect 2724 1708 2758 1742
rect 2797 1708 2831 1742
rect 2870 1708 2904 1742
rect 2943 1708 2977 1742
rect 3016 1708 3050 1742
rect 3089 1708 3123 1742
rect 3162 1708 3196 1742
rect 3235 1708 3269 1742
rect 3308 1708 3342 1742
rect 3381 1708 3415 1742
rect 3454 1708 3488 1742
rect 3527 1708 3561 1742
rect 3600 1708 3634 1742
rect 3673 1708 3707 1742
rect 3746 1708 3780 1742
rect 3819 1708 3853 1742
rect 3892 1708 3926 1742
rect 3965 1708 3999 1742
rect 4038 1708 4072 1742
rect 4111 1708 4145 1742
rect 4184 1708 4218 1742
rect 4257 1708 4291 1742
rect 4330 1708 4364 1742
rect 4403 1708 4437 1742
rect 4476 1708 4510 1742
rect 4549 1708 4583 1742
rect 4622 1708 4656 1742
rect 4695 1708 4729 1742
rect 4768 1708 4802 1742
rect 4841 1708 4875 1742
rect 4914 1708 4948 1742
rect 4987 1708 5021 1742
rect -2243 1542 -2209 1576
rect -1710 1593 -1676 1627
rect -1638 1593 -1604 1627
rect -2171 1542 -2137 1576
rect 4954 1548 4988 1582
rect 5026 1548 5060 1582
rect -2243 1220 -2209 1254
rect -2171 1220 -2137 1254
rect -2243 1147 -2209 1181
rect -2171 1147 -2137 1181
rect -2243 1074 -2209 1108
rect -2171 1074 -2137 1108
rect -2243 1001 -2209 1035
rect -2171 1001 -2137 1035
rect -2243 928 -2209 962
rect -2171 928 -2137 962
rect -2243 855 -2209 889
rect -2171 855 -2137 889
rect -2243 782 -2209 816
rect -2171 782 -2137 816
rect -2243 709 -2209 743
rect -2171 709 -2137 743
rect -2243 636 -2209 670
rect -2171 636 -2137 670
rect -2243 575 -2137 597
rect -2243 541 -2206 575
rect -2206 541 -2172 575
rect -2172 541 -2137 575
rect -2243 507 -2137 541
rect -2243 473 -2206 507
rect -2206 473 -2172 507
rect -2172 473 -2137 507
rect -2243 439 -2137 473
rect -2243 405 -2206 439
rect -2206 405 -2172 439
rect -2172 405 -2137 439
rect -2243 371 -2137 405
rect -2243 337 -2206 371
rect -2206 337 -2172 371
rect -2172 337 -2137 371
rect -2243 303 -2137 337
rect -2243 275 -2206 303
rect -2206 275 -2172 303
rect -2172 275 -2137 303
rect -1843 1474 -1833 1508
rect -1833 1474 -1809 1508
rect -1519 1474 -1485 1508
rect -1447 1474 -1417 1508
rect -1417 1474 -1413 1508
rect -1375 1474 -1349 1508
rect -1349 1474 -1341 1508
rect -1303 1474 -1281 1508
rect -1281 1474 -1269 1508
rect -1231 1474 -1213 1508
rect -1213 1474 -1197 1508
rect -1159 1474 -1145 1508
rect -1145 1474 -1125 1508
rect -1087 1474 -1077 1508
rect -1077 1474 -1053 1508
rect -1015 1474 -1009 1508
rect -1009 1474 -981 1508
rect -943 1474 -941 1508
rect -941 1474 -909 1508
rect -871 1474 -839 1508
rect -839 1474 -837 1508
rect -799 1474 -771 1508
rect -771 1474 -765 1508
rect -727 1474 -703 1508
rect -703 1474 -693 1508
rect -655 1474 -635 1508
rect -635 1474 -621 1508
rect -583 1474 -567 1508
rect -567 1474 -549 1508
rect -511 1474 -499 1508
rect -499 1474 -477 1508
rect -439 1474 -431 1508
rect -431 1474 -405 1508
rect -367 1474 -363 1508
rect -363 1474 -333 1508
rect -295 1474 -261 1508
rect -223 1474 -193 1508
rect -193 1474 -189 1508
rect -151 1474 -125 1508
rect -125 1474 -117 1508
rect -79 1474 -57 1508
rect -57 1474 -45 1508
rect -7 1474 11 1508
rect 11 1474 27 1508
rect 65 1474 79 1508
rect 79 1474 99 1508
rect 137 1474 147 1508
rect 147 1474 171 1508
rect 209 1474 215 1508
rect 215 1474 243 1508
rect 281 1474 283 1508
rect 283 1474 315 1508
rect 353 1474 385 1508
rect 385 1474 387 1508
rect 425 1474 453 1508
rect 453 1474 459 1508
rect 497 1474 521 1508
rect 521 1474 531 1508
rect 569 1474 589 1508
rect 589 1474 603 1508
rect 641 1474 657 1508
rect 657 1474 675 1508
rect 713 1474 725 1508
rect 725 1474 747 1508
rect 785 1474 793 1508
rect 793 1474 819 1508
rect 857 1474 861 1508
rect 861 1474 891 1508
rect 929 1474 963 1508
rect 1001 1474 1031 1508
rect 1031 1474 1035 1508
rect 1073 1474 1099 1508
rect 1099 1474 1107 1508
rect 1145 1474 1167 1508
rect 1167 1474 1179 1508
rect 1217 1474 1235 1508
rect 1235 1474 1251 1508
rect 1289 1474 1303 1508
rect 1303 1474 1323 1508
rect 1361 1474 1371 1508
rect 1371 1474 1395 1508
rect 1433 1474 1439 1508
rect 1439 1474 1467 1508
rect 1505 1474 1507 1508
rect 1507 1474 1539 1508
rect 1577 1474 1609 1508
rect 1609 1474 1611 1508
rect 1649 1474 1677 1508
rect 1677 1474 1683 1508
rect 1721 1474 1745 1508
rect 1745 1474 1755 1508
rect 1793 1474 1813 1508
rect 1813 1474 1827 1508
rect 1865 1474 1881 1508
rect 1881 1474 1899 1508
rect 1937 1474 1949 1508
rect 1949 1474 1971 1508
rect 2009 1474 2017 1508
rect 2017 1474 2043 1508
rect 2081 1474 2085 1508
rect 2085 1474 2115 1508
rect 2153 1474 2187 1508
rect 2225 1474 2255 1508
rect 2255 1474 2259 1508
rect 2297 1474 2323 1508
rect 2323 1474 2331 1508
rect 2369 1474 2391 1508
rect 2391 1474 2403 1508
rect 2442 1474 2459 1508
rect 2459 1474 2476 1508
rect 2515 1474 2527 1508
rect 2527 1474 2549 1508
rect 2588 1474 2595 1508
rect 2595 1474 2622 1508
rect 2661 1474 2663 1508
rect 2663 1474 2695 1508
rect 2734 1474 2765 1508
rect 2765 1474 2768 1508
rect 2807 1474 2833 1508
rect 2833 1474 2841 1508
rect 2880 1474 2901 1508
rect 2901 1474 2914 1508
rect 2953 1474 2969 1508
rect 2969 1474 2987 1508
rect 3026 1474 3037 1508
rect 3037 1474 3060 1508
rect 3099 1474 3105 1508
rect 3105 1474 3133 1508
rect 3172 1474 3173 1508
rect 3173 1474 3206 1508
rect 3245 1474 3273 1508
rect 3273 1474 3279 1508
rect 3318 1474 3341 1508
rect 3341 1474 3352 1508
rect 3391 1474 3409 1508
rect 3409 1474 3425 1508
rect 3464 1474 3477 1508
rect 3477 1474 3498 1508
rect 3537 1474 3545 1508
rect 3545 1474 3571 1508
rect 3610 1474 3613 1508
rect 3613 1474 3644 1508
rect 3683 1474 3715 1508
rect 3715 1474 3717 1508
rect 3756 1474 3783 1508
rect 3783 1474 3790 1508
rect 3829 1474 3851 1508
rect 3851 1474 3863 1508
rect 3902 1474 3919 1508
rect 3919 1474 3936 1508
rect 3975 1474 3987 1508
rect 3987 1474 4009 1508
rect 4048 1474 4055 1508
rect 4055 1474 4082 1508
rect 4121 1474 4123 1508
rect 4123 1474 4155 1508
rect 4194 1474 4225 1508
rect 4225 1474 4228 1508
rect 4267 1474 4293 1508
rect 4293 1474 4301 1508
rect 4340 1474 4361 1508
rect 4361 1474 4374 1508
rect 4413 1474 4429 1508
rect 4429 1474 4447 1508
rect 4486 1474 4497 1508
rect 4497 1474 4520 1508
rect 4559 1474 4565 1508
rect 4565 1474 4593 1508
rect 4632 1474 4633 1508
rect 4633 1474 4666 1508
rect 4705 1474 4735 1508
rect 4735 1474 4739 1508
rect 4778 1474 4803 1508
rect 4803 1474 4812 1508
rect 4851 1474 4871 1508
rect 4871 1474 4885 1508
rect -1710 1392 -1688 1426
rect -1688 1392 -1676 1426
rect -1638 1392 -1626 1426
rect -1626 1392 -1604 1426
rect -1458 1306 -1424 1340
rect -1386 1306 -1352 1340
rect -1202 1306 -1168 1340
rect -1130 1306 -1096 1340
rect -946 1306 -912 1340
rect -874 1306 -840 1340
rect -690 1306 -656 1340
rect -618 1306 -584 1340
rect -434 1306 -400 1340
rect -362 1306 -328 1340
rect -178 1306 -144 1340
rect -106 1306 -72 1340
rect 78 1306 112 1340
rect 150 1306 184 1340
rect 334 1306 368 1340
rect 406 1306 440 1340
rect 590 1306 624 1340
rect 662 1306 696 1340
rect 846 1306 880 1340
rect 918 1306 952 1340
rect 1102 1306 1136 1340
rect 1174 1306 1208 1340
rect 1358 1306 1392 1340
rect 1430 1306 1464 1340
rect 1614 1306 1648 1340
rect 1686 1306 1720 1340
rect 1870 1306 1904 1340
rect 1942 1306 1976 1340
rect 2126 1306 2160 1340
rect 2198 1306 2232 1340
rect 2382 1306 2416 1340
rect 2454 1306 2488 1340
rect 2638 1306 2672 1340
rect 2710 1306 2744 1340
rect 2894 1306 2928 1340
rect 2966 1306 3000 1340
rect 3150 1306 3184 1340
rect 3222 1306 3256 1340
rect 3406 1306 3440 1340
rect 3478 1306 3512 1340
rect 3662 1306 3696 1340
rect 3734 1306 3768 1340
rect 3918 1306 3952 1340
rect 3990 1306 4024 1340
rect 4954 1392 4973 1426
rect 4973 1392 4988 1426
rect 5026 1392 5044 1426
rect 5044 1392 5060 1426
rect 4525 1226 4559 1260
rect 4681 1226 4715 1260
rect 4837 1226 4871 1260
rect 4993 1226 5027 1260
rect 4759 1142 4793 1176
rect 4759 1070 4793 1104
rect 4759 998 4793 1032
rect 3313 927 3347 961
rect 3313 855 3347 889
rect 2033 818 2067 852
rect 2033 746 2067 780
rect 2033 674 2067 708
rect 2033 602 2067 636
rect 2033 530 2067 564
rect 2033 458 2067 492
rect 2033 386 2067 420
rect 3057 818 3091 852
rect 3057 746 3091 780
rect 3057 674 3091 708
rect 3057 602 3091 636
rect 3057 530 3091 564
rect 3313 783 3347 817
rect 3313 711 3347 745
rect 3313 639 3347 673
rect 3313 567 3347 601
rect 3313 495 3347 529
rect 3825 927 3859 961
rect 3825 855 3859 889
rect 3825 783 3859 817
rect 3825 711 3859 745
rect 4759 926 4793 960
rect 4759 854 4793 888
rect 4759 782 4793 816
rect 4759 710 4793 744
rect 7586 1108 7614 1139
rect 7614 1108 7620 1139
rect 7659 1108 7682 1139
rect 7682 1108 7693 1139
rect 7732 1108 7750 1139
rect 7750 1108 7766 1139
rect 7586 1105 7620 1108
rect 7659 1105 7693 1108
rect 7732 1105 7766 1108
rect 7805 1105 7839 1139
rect 7878 1108 7892 1139
rect 7892 1108 7912 1139
rect 7950 1108 7960 1139
rect 7960 1108 7984 1139
rect 8022 1108 8028 1139
rect 8028 1108 8056 1139
rect 7878 1105 7912 1108
rect 7950 1105 7984 1108
rect 8022 1105 8056 1108
rect 7771 1003 7785 1037
rect 7785 1003 7805 1037
rect 7843 1003 7847 1037
rect 7847 1003 7877 1037
rect 3825 639 3859 673
rect 3825 567 3859 601
rect 3825 495 3859 529
rect 3057 458 3091 492
rect 3057 386 3091 420
rect -1917 246 -1889 280
rect -1889 246 -1883 280
rect -1845 246 -1821 280
rect -1821 246 -1811 280
rect -1773 246 -1753 280
rect -1753 246 -1739 280
rect -1701 246 -1685 280
rect -1685 246 -1667 280
rect -1629 246 -1617 280
rect -1617 246 -1595 280
rect -1557 246 -1549 280
rect -1549 246 -1523 280
rect -1485 246 -1481 280
rect -1481 246 -1451 280
rect -1413 246 -1379 280
rect -1341 246 -1311 280
rect -1311 246 -1307 280
rect -1269 246 -1243 280
rect -1243 246 -1235 280
rect -1197 246 -1175 280
rect -1175 246 -1163 280
rect -1125 246 -1107 280
rect -1107 246 -1091 280
rect -1053 246 -1039 280
rect -1039 246 -1019 280
rect -981 246 -971 280
rect -971 246 -947 280
rect -909 246 -903 280
rect -903 246 -875 280
rect -837 246 -835 280
rect -835 246 -803 280
rect -765 246 -733 280
rect -733 246 -731 280
rect -693 246 -665 280
rect -665 246 -659 280
rect -621 246 -597 280
rect -597 246 -587 280
rect -549 246 -529 280
rect -529 246 -515 280
rect -477 246 -461 280
rect -461 246 -443 280
rect -405 246 -393 280
rect -393 246 -371 280
rect -333 246 -325 280
rect -325 246 -299 280
rect -261 246 -257 280
rect -257 246 -227 280
rect -189 246 -155 280
rect -117 246 -87 280
rect -87 246 -83 280
rect -45 246 -19 280
rect -19 246 -11 280
rect 27 246 49 280
rect 49 246 61 280
rect 99 246 117 280
rect 117 246 133 280
rect 171 246 185 280
rect 185 246 205 280
rect 243 246 253 280
rect 253 246 277 280
rect 315 246 321 280
rect 321 246 349 280
rect 387 246 389 280
rect 389 246 421 280
rect 460 246 491 280
rect 491 246 494 280
rect 533 246 559 280
rect 559 246 567 280
rect 606 246 627 280
rect 627 246 640 280
rect 679 246 695 280
rect 695 246 713 280
rect 752 246 763 280
rect 763 246 786 280
rect 825 246 831 280
rect 831 246 859 280
rect 898 246 899 280
rect 899 246 932 280
rect 971 246 1001 280
rect 1001 246 1005 280
rect 1044 246 1069 280
rect 1069 246 1078 280
rect 1117 246 1137 280
rect 1137 246 1151 280
rect 1190 246 1205 280
rect 1205 246 1224 280
rect 1263 246 1273 280
rect 1273 246 1297 280
rect 1336 246 1341 280
rect 1341 246 1370 280
rect 1409 246 1443 280
rect 1482 246 1511 280
rect 1511 246 1516 280
rect 1555 246 1579 280
rect 1579 246 1589 280
rect 1628 246 1647 280
rect 1647 246 1662 280
rect 1701 246 1715 280
rect 1715 246 1735 280
rect 1774 246 1783 280
rect 1783 246 1808 280
rect 1847 246 1851 280
rect 1851 246 1881 280
rect 1920 246 1953 280
rect 1953 246 1954 280
rect 1993 246 2021 280
rect 2021 246 2027 280
rect 2066 246 2089 280
rect 2089 246 2100 280
rect 2139 246 2157 280
rect 2157 246 2173 280
rect 2212 246 2225 280
rect 2225 246 2246 280
rect 2285 246 2293 280
rect 2293 246 2319 280
rect 2358 246 2361 280
rect 2361 246 2392 280
rect 2431 246 2463 280
rect 2463 246 2465 280
rect 2504 246 2531 280
rect 2531 246 2538 280
rect 2577 246 2599 280
rect 2599 246 2611 280
rect 2650 246 2667 280
rect 2667 246 2684 280
rect 2723 246 2735 280
rect 2735 246 2757 280
rect 2796 246 2803 280
rect 2803 246 2830 280
rect 2869 246 2871 280
rect 2871 246 2903 280
rect 2942 246 2973 280
rect 2973 246 2976 280
rect 3015 246 3041 280
rect 3041 246 3049 280
rect 3088 246 3109 280
rect 3109 246 3122 280
rect 3161 246 3177 280
rect 3177 246 3195 280
rect 3234 246 3245 280
rect 3245 246 3268 280
rect 3307 246 3313 280
rect 3313 246 3341 280
rect 3380 246 3381 280
rect 3381 246 3414 280
rect 3453 246 3483 280
rect 3483 246 3487 280
rect 3526 246 3551 280
rect 3551 246 3560 280
rect 3599 246 3619 280
rect 3619 246 3633 280
rect 3672 246 3687 280
rect 3687 246 3706 280
rect 3745 246 3755 280
rect 3755 246 3779 280
rect 3818 246 3823 280
rect 3823 246 3852 280
rect 3891 246 3925 280
rect 3964 246 3993 280
rect 3993 246 3998 280
rect 4037 246 4061 280
rect 4061 246 4071 280
rect 4110 246 4129 280
rect 4129 246 4144 280
rect 4183 246 4197 280
rect 4197 246 4217 280
rect 4256 246 4265 280
rect 4265 246 4290 280
rect 4329 246 4333 280
rect 4333 246 4363 280
rect 4402 246 4435 280
rect 4435 246 4436 280
rect 4475 246 4503 280
rect 4503 246 4509 280
rect 4548 246 4571 280
rect 4571 246 4582 280
rect 4621 246 4639 280
rect 4639 246 4655 280
rect 4694 246 4707 280
rect 4707 246 4728 280
rect 4767 246 4775 280
rect 4775 246 4801 280
rect 4840 246 4843 280
rect 4843 246 4874 280
rect 4913 246 4945 280
rect 4945 246 4947 280
rect 4986 246 5013 280
rect 5013 246 5020 280
rect 5059 246 5081 280
rect 5081 246 5093 280
rect -2194 -37 -2160 -3
rect -2122 -13 -2109 -3
rect -2109 -13 -2088 -3
rect -2122 -37 -2088 -13
rect -2050 -37 -2016 -3
rect -1978 -37 -1975 -3
rect -1975 -37 -1944 -3
rect -1906 -37 -1873 -3
rect -1873 -37 -1872 -3
rect -1834 -37 -1805 -3
rect -1805 -37 -1800 -3
rect -1762 -37 -1737 -3
rect -1737 -37 -1728 -3
rect -1690 -37 -1669 -3
rect -1669 -37 -1656 -3
rect -1618 -37 -1601 -3
rect -1601 -37 -1584 -3
rect -1546 -37 -1533 -3
rect -1533 -37 -1512 -3
rect -1474 -37 -1465 -3
rect -1465 -37 -1440 -3
rect -1402 -37 -1397 -3
rect -1397 -37 -1368 -3
rect -1330 -37 -1329 -3
rect -1329 -37 -1296 -3
rect -1258 -37 -1227 -3
rect -1227 -37 -1224 -3
rect -1186 -37 -1159 -3
rect -1159 -37 -1152 -3
rect -1114 -37 -1091 -3
rect -1091 -37 -1080 -3
rect -1042 -37 -1023 -3
rect -1023 -37 -1008 -3
rect -970 -37 -955 -3
rect -955 -37 -936 -3
rect -898 -37 -887 -3
rect -887 -37 -864 -3
rect -826 -37 -819 -3
rect -819 -37 -792 -3
rect -754 -37 -751 -3
rect -751 -37 -720 -3
rect -682 -37 -649 -3
rect -649 -37 -648 -3
rect -610 -37 -581 -3
rect -581 -37 -576 -3
rect -538 -37 -513 -3
rect -513 -37 -504 -3
rect -466 -37 -445 -3
rect -445 -37 -432 -3
rect -394 -37 -377 -3
rect -377 -37 -360 -3
rect -322 -37 -309 -3
rect -309 -37 -288 -3
rect -250 -37 -241 -3
rect -241 -37 -216 -3
rect -178 -37 -173 -3
rect -173 -37 -144 -3
rect -106 -37 -105 -3
rect -105 -37 -72 -3
rect -34 -37 -3 -3
rect -3 -37 0 -3
rect 38 -37 65 -3
rect 65 -37 72 -3
rect 110 -37 133 -3
rect 133 -37 144 -3
rect 182 -37 201 -3
rect 201 -37 216 -3
rect 254 -37 269 -3
rect 269 -37 288 -3
rect 326 -37 337 -3
rect 337 -37 360 -3
rect 398 -37 405 -3
rect 405 -37 432 -3
rect 470 -37 473 -3
rect 473 -37 504 -3
rect 542 -37 575 -3
rect 575 -37 576 -3
rect 614 -37 643 -3
rect 643 -37 648 -3
rect 686 -37 711 -3
rect 711 -37 720 -3
rect 758 -37 779 -3
rect 779 -37 792 -3
rect 830 -37 847 -3
rect 847 -37 864 -3
rect 902 -37 915 -3
rect 915 -37 936 -3
rect 974 -37 983 -3
rect 983 -37 1008 -3
rect 1046 -37 1051 -3
rect 1051 -37 1080 -3
rect 1118 -37 1119 -3
rect 1119 -37 1152 -3
rect 1190 -37 1221 -3
rect 1221 -37 1224 -3
rect 1262 -37 1289 -3
rect 1289 -37 1296 -3
rect 1334 -37 1357 -3
rect 1357 -37 1368 -3
rect 1406 -37 1425 -3
rect 1425 -37 1440 -3
rect 1478 -37 1493 -3
rect 1493 -37 1512 -3
rect 1550 -37 1561 -3
rect 1561 -37 1584 -3
rect 1622 -37 1629 -3
rect 1629 -37 1656 -3
rect 1694 -37 1697 -3
rect 1697 -37 1728 -3
rect 1766 -37 1799 -3
rect 1799 -37 1800 -3
rect 1838 -37 1867 -3
rect 1867 -37 1872 -3
rect 1910 -37 1935 -3
rect 1935 -37 1944 -3
rect 1982 -37 2003 -3
rect 2003 -37 2016 -3
rect 2054 -37 2071 -3
rect 2071 -37 2088 -3
rect 2126 -37 2139 -3
rect 2139 -37 2160 -3
rect 2198 -37 2207 -3
rect 2207 -37 2232 -3
rect 2270 -37 2275 -3
rect 2275 -37 2304 -3
rect 2343 -37 2377 -3
rect 2416 -37 2445 -3
rect 2445 -37 2450 -3
rect 2489 -37 2513 -3
rect 2513 -37 2523 -3
rect 2562 -37 2581 -3
rect 2581 -37 2596 -3
rect 2635 -37 2649 -3
rect 2649 -37 2669 -3
rect 2708 -37 2717 -3
rect 2717 -37 2742 -3
rect 2781 -37 2785 -3
rect 2785 -37 2815 -3
rect 2854 -37 2887 -3
rect 2887 -37 2888 -3
rect 2927 -37 2955 -3
rect 2955 -37 2961 -3
rect 3000 -37 3023 -3
rect 3023 -37 3034 -3
rect 3073 -37 3091 -3
rect 3091 -37 3107 -3
rect 3146 -37 3159 -3
rect 3159 -37 3180 -3
rect 3219 -37 3227 -3
rect 3227 -37 3253 -3
rect 3292 -37 3295 -3
rect 3295 -37 3326 -3
rect 3365 -37 3397 -3
rect 3397 -37 3399 -3
rect 3438 -37 3465 -3
rect 3465 -37 3472 -3
rect 3511 -37 3533 -3
rect 3533 -37 3545 -3
rect 3584 -37 3601 -3
rect 3601 -37 3618 -3
rect 3657 -37 3669 -3
rect 3669 -37 3691 -3
rect 3730 -37 3737 -3
rect 3737 -37 3764 -3
rect 3803 -37 3805 -3
rect 3805 -37 3837 -3
rect 3876 -37 3907 -3
rect 3907 -37 3910 -3
rect 3949 -37 3975 -3
rect 3975 -37 3983 -3
rect 4022 -37 4043 -3
rect 4043 -37 4056 -3
rect 4095 -37 4111 -3
rect 4111 -37 4129 -3
rect 4168 -37 4179 -3
rect 4179 -37 4202 -3
rect 4241 -37 4247 -3
rect 4247 -37 4275 -3
rect 4314 -37 4315 -3
rect 4315 -37 4348 -3
rect 4387 -37 4417 -3
rect 4417 -37 4421 -3
rect 4460 -37 4485 -3
rect 4485 -37 4494 -3
rect 4533 -37 4553 -3
rect 4553 -37 4567 -3
rect 4606 -37 4621 -3
rect 4621 -37 4640 -3
rect 4679 -37 4689 -3
rect 4689 -37 4713 -3
rect 4752 -37 4757 -3
rect 4757 -37 4786 -3
rect 4825 -37 4859 -3
rect 4898 -37 4927 -3
rect 4927 -37 4932 -3
rect 4971 -37 4995 -3
rect 4995 -37 5005 -3
rect 7586 -133 7620 -99
rect 7659 -133 7693 -99
rect 7732 -133 7742 -99
rect 7742 -133 7766 -99
rect 7805 -133 7810 -99
rect 7810 -133 7839 -99
rect 7878 -133 7912 -99
rect 7950 -133 7980 -99
rect 7980 -133 7984 -99
rect 8022 -133 8056 -99
<< metal1 >>
rect -2302 1867 5070 1893
rect -2302 1865 -2131 1867
tri -2302 1820 -2257 1865 ne
rect -2257 1820 -2131 1865
tri -2257 1814 -2251 1820 ne
rect -2251 1815 -2131 1820
rect -2079 1815 -2066 1867
rect -2014 1815 5070 1867
rect -2251 1814 5070 1815
tri -2251 1746 -2183 1814 ne
rect -2183 1803 -2127 1814
rect -2183 1751 -2131 1803
rect 787 1780 826 1814
rect 860 1780 899 1814
rect 933 1780 972 1814
rect 1006 1780 1045 1814
rect 1079 1780 1118 1814
rect 1152 1780 1191 1814
rect 1225 1780 1264 1814
rect 1298 1780 1337 1814
rect 1371 1780 1410 1814
rect 1444 1780 1483 1814
rect 1517 1780 1556 1814
rect 1590 1780 1629 1814
rect 1663 1780 1702 1814
rect 1736 1780 1775 1814
rect 1809 1780 1848 1814
rect 1882 1780 1921 1814
rect 1955 1780 1994 1814
rect 2028 1780 2067 1814
rect 2101 1780 2140 1814
rect 2174 1780 2213 1814
rect 2247 1780 2286 1814
rect 2320 1780 2359 1814
rect 2393 1780 2432 1814
rect 2466 1780 2505 1814
rect 2539 1780 2578 1814
rect 2612 1780 2651 1814
rect 2685 1780 2724 1814
rect 2758 1780 2797 1814
rect 2831 1780 2870 1814
rect 2904 1780 2943 1814
rect 2977 1780 3016 1814
rect 3050 1780 3089 1814
rect 3123 1780 3162 1814
rect 3196 1780 3235 1814
rect 3269 1780 3308 1814
rect 3342 1780 3381 1814
rect 3415 1780 3454 1814
rect 3488 1780 3527 1814
rect 3561 1780 3600 1814
rect 3634 1780 3673 1814
rect 3707 1780 3746 1814
rect 3780 1780 3819 1814
rect 3853 1780 3892 1814
rect 3926 1780 3965 1814
rect 3999 1780 4038 1814
rect 4072 1780 4111 1814
rect 4145 1780 4184 1814
rect 4218 1780 4257 1814
rect 4291 1780 4330 1814
rect 4364 1780 4403 1814
rect 4437 1780 4476 1814
rect 4510 1780 4549 1814
rect 4583 1780 4622 1814
rect 4656 1780 4695 1814
rect 4729 1780 4768 1814
rect 4802 1780 4841 1814
rect 4875 1780 4914 1814
rect 4948 1780 4987 1814
rect 5021 1780 5070 1814
rect -2183 1746 -2127 1751
rect -2298 1740 -2246 1746
tri -2183 1708 -2145 1746 ne
rect -2145 1708 -2127 1746
rect 787 1742 5070 1780
rect 787 1708 826 1742
rect 860 1708 899 1742
rect 933 1708 972 1742
rect 1006 1708 1045 1742
rect 1079 1708 1118 1742
rect 1152 1708 1191 1742
rect 1225 1708 1264 1742
rect 1298 1708 1337 1742
rect 1371 1708 1410 1742
rect 1444 1708 1483 1742
rect 1517 1708 1556 1742
rect 1590 1708 1629 1742
rect 1663 1708 1702 1742
rect 1736 1708 1775 1742
rect 1809 1708 1848 1742
rect 1882 1708 1921 1742
rect 1955 1708 1994 1742
rect 2028 1708 2067 1742
rect 2101 1708 2140 1742
rect 2174 1708 2213 1742
rect 2247 1708 2286 1742
rect 2320 1708 2359 1742
rect 2393 1708 2432 1742
rect 2466 1708 2505 1742
rect 2539 1708 2578 1742
rect 2612 1708 2651 1742
rect 2685 1708 2724 1742
rect 2758 1708 2797 1742
rect 2831 1708 2870 1742
rect 2904 1708 2943 1742
rect 2977 1708 3016 1742
rect 3050 1708 3089 1742
rect 3123 1708 3162 1742
rect 3196 1708 3235 1742
rect 3269 1708 3308 1742
rect 3342 1708 3381 1742
rect 3415 1708 3454 1742
rect 3488 1708 3527 1742
rect 3561 1708 3600 1742
rect 3634 1708 3673 1742
rect 3707 1708 3746 1742
rect 3780 1708 3819 1742
rect 3853 1708 3892 1742
rect 3926 1708 3965 1742
rect 3999 1708 4038 1742
rect 4072 1708 4111 1742
rect 4145 1708 4184 1742
rect 4218 1708 4257 1742
rect 4291 1708 4330 1742
rect 4364 1708 4403 1742
rect 4437 1708 4476 1742
rect 4510 1708 4549 1742
rect 4583 1708 4622 1742
rect 4656 1708 4695 1742
rect 4729 1708 4768 1742
rect 4802 1708 4841 1742
rect 4875 1708 4914 1742
rect 4948 1708 4987 1742
rect 5021 1708 5070 1742
tri -2145 1702 -2139 1708 ne
rect -2139 1702 5070 1708
tri -2800 1675 -2790 1685 se
tri -2406 1675 -2398 1683 sw
rect -2298 1674 -2246 1688
tri -2246 1662 -2221 1687 sw
rect -2246 1656 7811 1662
rect -2246 1627 7759 1656
rect -2246 1622 -1710 1627
rect -2298 1616 -1710 1622
tri -1751 1593 -1728 1616 ne
rect -1728 1593 -1710 1616
rect -1676 1593 -1638 1627
rect -1604 1616 7759 1627
rect -1604 1593 -1591 1616
tri -1728 1588 -1723 1593 ne
rect -1723 1588 -1591 1593
tri -1591 1588 -1563 1616 nw
tri 7734 1591 7759 1616 ne
rect 7759 1592 7811 1604
rect -2249 1582 -2021 1588
tri -1723 1587 -1722 1588 ne
rect -2249 1576 -2137 1582
rect -2249 1542 -2243 1576
rect -2209 1542 -2171 1576
rect -2249 1466 -2137 1542
tri -1869 1508 -1863 1514 se
rect -1863 1508 -1771 1514
tri -1903 1474 -1869 1508 se
rect -1869 1474 -1843 1508
rect -1809 1474 -1771 1508
tri -1909 1468 -1903 1474 se
rect -1903 1468 -1771 1474
rect -2249 1460 -2021 1466
tri -1917 1460 -1909 1468 se
rect -1909 1460 -1863 1468
tri -1929 1448 -1917 1460 se
rect -1917 1448 -1863 1460
tri -1863 1448 -1843 1468 nw
rect -1929 1432 -1879 1448
tri -1879 1432 -1863 1448 nw
rect -1929 1266 -1883 1432
tri -1883 1428 -1879 1432 nw
rect -1722 1426 -1592 1588
tri -1592 1587 -1591 1588 nw
rect 4942 1582 7597 1588
rect 4942 1548 4954 1582
rect 4988 1548 5026 1582
rect 5060 1548 7597 1582
rect 4942 1542 5499 1548
tri 5499 1542 5505 1548 nw
tri 5795 1542 5801 1548 ne
rect 5801 1542 7597 1548
rect 4942 1536 5091 1542
tri 5091 1536 5097 1542 nw
tri 7585 1536 7591 1542 ne
rect 7591 1536 7597 1542
rect 7649 1536 7661 1588
rect 7713 1536 7719 1588
rect -1531 1508 -1510 1514
rect -1458 1508 -1440 1514
rect -1388 1508 -1370 1514
rect -1318 1508 -1301 1514
rect -1531 1474 -1519 1508
rect -1458 1474 -1447 1508
rect -1388 1474 -1375 1508
rect -1318 1474 -1303 1508
rect -1531 1468 -1510 1474
tri -1522 1462 -1516 1468 ne
rect -1516 1462 -1510 1468
rect -1458 1462 -1440 1474
rect -1388 1462 -1370 1474
rect -1318 1462 -1301 1474
rect -1249 1462 -1232 1514
rect -1180 1462 -1163 1514
rect -1111 1462 -1094 1514
rect -1042 1462 -1025 1514
rect -973 1462 -956 1514
rect -904 1462 -887 1514
rect -835 1462 -818 1514
rect -766 1508 -749 1514
rect -697 1508 4897 1514
rect -765 1474 -749 1508
rect -693 1474 -655 1508
rect -621 1474 -583 1508
rect -549 1474 -511 1508
rect -477 1474 -439 1508
rect -405 1474 -367 1508
rect -333 1474 -295 1508
rect -261 1474 -223 1508
rect -189 1474 -151 1508
rect -117 1474 -79 1508
rect -45 1474 -7 1508
rect 27 1474 65 1508
rect 99 1474 137 1508
rect 171 1474 209 1508
rect 243 1474 281 1508
rect 315 1474 353 1508
rect 387 1474 425 1508
rect 459 1474 497 1508
rect 531 1474 569 1508
rect 603 1474 641 1508
rect 675 1474 713 1508
rect 747 1474 785 1508
rect 819 1474 857 1508
rect 891 1474 929 1508
rect 963 1474 1001 1508
rect 1035 1474 1073 1508
rect 1107 1474 1145 1508
rect 1179 1474 1217 1508
rect 1251 1474 1289 1508
rect 1323 1474 1361 1508
rect 1395 1474 1433 1508
rect 1467 1474 1505 1508
rect 1539 1474 1577 1508
rect 1611 1474 1649 1508
rect 1683 1474 1721 1508
rect 1755 1474 1793 1508
rect 1827 1474 1865 1508
rect 1899 1474 1937 1508
rect 1971 1474 2009 1508
rect 2043 1474 2081 1508
rect 2115 1474 2153 1508
rect 2187 1474 2225 1508
rect 2259 1474 2297 1508
rect 2331 1474 2369 1508
rect 2403 1474 2442 1508
rect 2476 1474 2515 1508
rect 2549 1474 2588 1508
rect 2622 1474 2661 1508
rect 2695 1474 2734 1508
rect 2768 1474 2807 1508
rect 2841 1474 2880 1508
rect 2914 1474 2953 1508
rect 2987 1474 3026 1508
rect 3060 1474 3099 1508
rect 3133 1474 3172 1508
rect 3206 1474 3245 1508
rect 3279 1474 3318 1508
rect 3352 1474 3391 1508
rect 3425 1474 3464 1508
rect 3498 1474 3537 1508
rect 3571 1474 3610 1508
rect 3644 1474 3683 1508
rect 3717 1474 3756 1508
rect 3790 1474 3829 1508
rect 3863 1474 3902 1508
rect 3936 1474 3975 1508
rect 4009 1474 4048 1508
rect 4082 1474 4121 1508
rect 4155 1474 4194 1508
rect 4228 1474 4267 1508
rect 4301 1474 4340 1508
rect 4374 1474 4413 1508
rect 4447 1474 4486 1508
rect 4520 1474 4559 1508
rect 4593 1474 4632 1508
rect 4666 1474 4705 1508
rect 4739 1474 4778 1508
rect 4812 1474 4851 1508
rect 4885 1474 4897 1508
rect -766 1462 -749 1474
rect -697 1468 4897 1474
rect -697 1462 -691 1468
tri -691 1462 -685 1468 nw
rect -1722 1392 -1710 1426
rect -1676 1392 -1638 1426
rect -1604 1392 -1592 1426
rect -1722 1386 -1592 1392
rect 4942 1426 5072 1536
tri 5072 1517 5091 1536 nw
rect 7759 1534 7811 1540
rect 4942 1392 4954 1426
rect 4988 1392 5026 1426
rect 5060 1392 5072 1426
rect 4942 1386 5072 1392
rect -1470 1340 5143 1346
rect -1470 1306 -1458 1340
rect -1424 1306 -1386 1340
rect -1352 1306 -1202 1340
rect -1168 1306 -1130 1340
rect -1096 1306 -946 1340
rect -912 1306 -874 1340
rect -840 1306 -690 1340
rect -656 1306 -618 1340
rect -584 1306 -434 1340
rect -400 1306 -362 1340
rect -328 1306 -178 1340
rect -144 1306 -106 1340
rect -72 1306 78 1340
rect 112 1306 150 1340
rect 184 1306 334 1340
rect 368 1306 406 1340
rect 440 1306 590 1340
rect 624 1306 662 1340
rect 696 1306 846 1340
rect 880 1306 918 1340
rect 952 1306 1102 1340
rect 1136 1306 1174 1340
rect 1208 1306 1358 1340
rect 1392 1306 1430 1340
rect 1464 1306 1614 1340
rect 1648 1306 1686 1340
rect 1720 1306 1870 1340
rect 1904 1306 1942 1340
rect 1976 1306 2126 1340
rect 2160 1306 2198 1340
rect 2232 1306 2382 1340
rect 2416 1306 2454 1340
rect 2488 1306 2638 1340
rect 2672 1306 2710 1340
rect 2744 1306 2894 1340
rect 2928 1306 2966 1340
rect 3000 1306 3150 1340
rect 3184 1306 3222 1340
rect 3256 1306 3406 1340
rect 3440 1306 3478 1340
rect 3512 1306 3662 1340
rect 3696 1306 3734 1340
rect 3768 1306 3918 1340
rect 3952 1306 3990 1340
rect 4024 1306 5143 1340
rect -1470 1294 5143 1306
rect -2249 1260 -2021 1266
rect -2249 1254 -2137 1260
rect -2902 1183 -2450 1235
rect -2398 1183 -2384 1235
rect -2332 1183 -2326 1235
rect -2249 1220 -2243 1254
rect -2209 1220 -2171 1254
rect -2249 1208 -2137 1220
rect -2085 1208 -2073 1260
rect -2249 1193 -2021 1208
rect -1767 1260 5039 1266
rect -1767 1226 4525 1260
rect 4559 1226 4681 1260
rect 4715 1226 4837 1260
rect 4871 1226 4993 1260
rect 5027 1226 5039 1260
rect -1767 1220 5039 1226
rect -1767 1200 -1762 1220
tri -1762 1200 -1742 1220 nw
tri -1767 1195 -1762 1200 nw
rect -2249 1181 -2137 1193
rect -2249 1147 -2243 1181
rect -2209 1147 -2171 1181
rect -2249 1141 -2137 1147
rect -2085 1141 -2073 1193
rect -2249 1126 -2021 1141
rect -2902 1069 -2450 1121
rect -2398 1069 -2384 1121
rect -2332 1069 -2326 1121
rect -2249 1108 -2137 1126
rect -2249 1074 -2243 1108
rect -2209 1074 -2171 1108
rect -2085 1074 -2073 1126
rect -1301 1092 -179 1192
rect -177 1191 -141 1192
rect -178 1093 -140 1191
rect -139 1176 5111 1192
rect -139 1142 4759 1176
rect 4793 1142 5111 1176
rect -139 1104 5111 1142
rect -177 1092 -141 1093
rect -139 1092 4759 1104
rect -2249 1059 -2021 1074
rect -1255 1070 -1252 1092
tri -1252 1070 -1230 1092 nw
tri -814 1070 -792 1092 ne
rect -792 1070 -789 1092
rect -1255 1069 -1253 1070
tri -1253 1069 -1252 1070 nw
tri -792 1069 -791 1070 ne
rect -791 1069 -789 1070
tri -1255 1067 -1253 1069 nw
tri -791 1067 -789 1069 ne
rect -743 1070 -740 1092
tri -740 1070 -718 1092 nw
tri -302 1070 -280 1092 ne
rect -280 1070 -277 1092
tri -743 1067 -740 1070 nw
tri -280 1067 -277 1070 ne
rect -231 1070 -228 1092
tri -228 1070 -206 1092 nw
tri 2025 1070 2047 1092 ne
rect 2047 1070 2153 1092
tri 2153 1070 2175 1092 nw
tri 3049 1070 3071 1092 ne
rect 3071 1070 3177 1092
tri 3177 1070 3199 1092 nw
tri 3282 1070 3304 1092 ne
rect 3304 1070 3356 1092
tri 3356 1070 3378 1092 nw
tri 3794 1070 3816 1092 ne
rect 3816 1070 3868 1092
tri 3868 1070 3890 1092 nw
tri 4414 1070 4436 1092 ne
rect 4436 1070 4439 1092
tri -231 1067 -228 1070 nw
tri 2047 1067 2050 1070 ne
rect -2249 1035 -2137 1059
rect -2249 1001 -2243 1035
rect -2209 1001 -2171 1035
rect -2085 1007 -2073 1059
rect -2137 1001 -2021 1007
rect -2902 944 -2450 996
rect -2398 944 -2384 996
rect -2332 944 -2326 996
rect -2249 992 -2021 1001
rect -2249 962 -2137 992
rect -2249 928 -2243 962
rect -2209 928 -2171 962
rect -2085 940 -2073 992
rect 235 964 1842 1064
rect 1843 965 1844 1063
rect 1880 965 1881 1063
rect 1882 1037 1934 1064
tri 1934 1037 1961 1064 sw
rect 1882 1032 1961 1037
tri 1961 1032 1966 1037 sw
rect 1882 1007 1966 1032
tri 1966 1007 1991 1032 sw
tri 2025 1007 2050 1032 se
rect 2050 1007 2150 1070
tri 2150 1067 2153 1070 nw
tri 3071 1067 3074 1070 ne
rect 1882 977 2150 1007
rect 1882 964 2137 977
tri 2137 964 2150 977 nw
rect 2283 964 2866 1064
rect 2867 965 2868 1063
rect 2906 1063 2958 1064
tri 2958 1063 2959 1064 sw
rect 2904 965 2905 1063
rect 2906 1037 2959 1063
tri 2959 1037 2985 1063 sw
rect 2906 1032 2985 1037
tri 2985 1032 2990 1037 sw
rect 2906 1027 2990 1032
tri 2990 1027 2995 1032 sw
tri 3069 1027 3074 1032 se
rect 3074 1027 3174 1070
tri 3174 1067 3177 1070 nw
tri 3304 1067 3307 1070 ne
rect 3307 1065 3353 1070
tri 3353 1067 3356 1070 nw
tri 3816 1067 3819 1070 ne
rect 3308 1063 3352 1064
rect 3819 1065 3865 1070
tri 3865 1067 3868 1070 nw
tri 4436 1067 4439 1070 ne
rect 4485 1070 4488 1092
tri 4488 1070 4510 1092 nw
tri 4728 1070 4750 1092 ne
rect 4750 1070 4759 1092
rect 4793 1092 5111 1104
rect 6944 1139 8068 1200
rect 6944 1105 7586 1139
rect 7620 1105 7659 1139
rect 7693 1105 7732 1139
rect 7766 1105 7805 1139
rect 7839 1105 7878 1139
rect 7912 1105 7950 1139
rect 7984 1105 8022 1139
rect 8056 1105 8068 1139
rect 6944 1096 8068 1105
rect 4793 1070 4799 1092
tri 4485 1067 4488 1070 nw
tri 4750 1067 4753 1070 ne
rect 3820 1063 3864 1064
rect 3819 1027 3865 1063
rect 2906 1007 2995 1027
tri 2995 1007 3015 1027 sw
tri 3049 1007 3069 1027 se
rect 3069 1007 3174 1027
rect 2906 977 3174 1007
rect 2906 964 3161 977
tri 3161 964 3174 977 nw
rect 3308 1026 3352 1027
rect -2137 928 -2021 940
rect 281 961 303 964
tri 303 961 306 964 nw
tri 722 961 725 964 ne
rect 725 961 747 964
tri 281 939 303 961 nw
tri 725 939 747 961 ne
rect 793 961 815 964
tri 815 961 818 964 nw
tri 1234 961 1237 964 ne
rect 1237 961 1259 964
tri 793 939 815 961 nw
tri 1237 939 1259 961 ne
rect 1305 961 1327 964
tri 1327 961 1330 964 nw
tri 1746 961 1749 964 ne
rect 1749 961 1771 964
tri 1305 939 1327 961 nw
tri 1749 939 1771 961 ne
rect 1817 961 1839 964
tri 1839 961 1842 964 nw
tri 1892 961 1895 964 ne
rect 1895 961 2134 964
tri 2134 961 2137 964 nw
rect 2329 961 2351 964
tri 2351 961 2354 964 nw
tri 2770 961 2773 964 ne
rect 2773 961 2795 964
rect 1817 944 1822 961
tri 1822 944 1839 961 nw
tri 1895 944 1912 961 ne
rect 1912 944 2112 961
tri 1817 939 1822 944 nw
tri 1912 939 1917 944 ne
rect 1917 939 2112 944
tri 2112 939 2134 961 nw
tri 2329 939 2351 961 nw
tri 2773 939 2795 961 ne
rect 2841 961 2863 964
tri 2863 961 2866 964 nw
tri 2916 961 2919 964 ne
rect 2919 961 3158 964
tri 3158 961 3161 964 nw
rect 3307 961 3353 1025
rect 2841 944 2846 961
tri 2846 944 2863 961 nw
tri 2919 944 2936 961 ne
rect 2936 944 3124 961
tri 2841 939 2846 944 nw
tri 2936 939 2941 944 ne
rect 2941 939 3124 944
rect -2249 925 -2021 928
tri 1917 927 1929 939 ne
rect 1929 927 2100 939
tri 2100 927 2112 939 nw
tri 2941 927 2953 939 ne
rect 2953 927 3124 939
tri 3124 927 3158 961 nw
rect 3307 927 3313 961
rect 3347 927 3353 961
tri 1929 926 1930 927 ne
rect 1930 926 2099 927
tri 2099 926 2100 927 nw
tri 2953 926 2954 927 ne
rect 2954 926 3123 927
tri 3123 926 3124 927 nw
rect -2249 889 -2137 925
rect -2249 855 -2243 889
rect -2209 855 -2171 889
rect -2085 873 -2073 925
tri 1930 907 1949 926 ne
rect 1949 907 2080 926
tri 2080 907 2099 926 nw
tri 2954 907 2973 926 ne
rect 2973 907 3104 926
tri 3104 907 3123 926 nw
rect -2137 858 -2021 873
rect 3307 889 3353 927
rect -2249 816 -2137 855
rect -2249 782 -2243 816
rect -2209 782 -2171 816
rect -2085 806 -2073 858
rect -2137 791 -2021 806
rect -2249 743 -2137 782
rect -2249 709 -2243 743
rect -2209 709 -2171 743
rect -2085 739 -2073 791
rect -2137 724 -2021 739
rect -2249 672 -2137 709
rect -2085 672 -2073 724
rect -2249 670 -2021 672
rect -2249 636 -2243 670
rect -2209 636 -2171 670
rect -2137 657 -2021 670
rect -2249 605 -2137 636
rect -2085 605 -2073 657
rect -2249 597 -2021 605
tri -2406 275 -2405 276 sw
rect -2249 275 -2243 597
rect -2137 590 -2021 597
rect -2085 538 -2073 590
rect -2137 523 -2021 538
rect -2085 471 -2073 523
rect -2137 456 -2021 471
rect 2027 852 2073 864
rect 2027 818 2033 852
rect 2067 818 2073 852
rect 2027 780 2073 818
rect 2027 746 2033 780
rect 2067 746 2073 780
rect 2027 708 2073 746
rect 2027 674 2033 708
rect 2067 674 2073 708
rect 2027 636 2073 674
rect 2027 602 2033 636
rect 2067 602 2073 636
rect 2027 564 2073 602
rect 2027 530 2033 564
rect 2067 530 2073 564
rect 2027 492 2073 530
rect -2085 404 -2073 456
rect -2137 389 -2021 404
rect -2085 337 -2073 389
tri -1883 458 -1876 465 sw
tri -1564 458 -1557 465 se
rect -1883 440 -1876 458
tri -1876 440 -1858 458 sw
tri -1582 440 -1564 458 se
rect -1564 440 -1557 458
tri -1511 458 -1504 465 sw
tri -1052 458 -1045 465 se
rect -1511 440 -1504 458
tri -1504 440 -1486 458 sw
tri -1070 440 -1052 458 se
rect -1052 440 -1045 458
tri -999 458 -992 465 sw
tri -540 458 -533 465 se
rect -999 440 -992 458
tri -992 440 -974 458 sw
tri -558 440 -540 458 se
rect -540 440 -533 458
tri -487 458 -480 465 sw
tri -28 458 -21 465 se
rect -487 440 -480 458
tri -480 440 -462 458 sw
tri -46 440 -28 458 se
rect -28 440 -21 458
tri 25 458 32 465 sw
tri 484 458 491 465 se
rect 25 440 32 458
tri 32 440 50 458 sw
tri 466 440 484 458 se
rect 484 440 491 458
tri 537 458 544 465 sw
tri 996 458 1003 465 se
rect 537 440 544 458
tri 544 440 562 458 sw
tri 978 440 996 458 se
rect 996 440 1003 458
tri 1049 458 1056 465 sw
tri 1508 458 1515 465 se
rect 1049 440 1056 458
tri 1056 440 1074 458 sw
tri 1490 440 1508 458 se
rect 1508 440 1515 458
tri 1561 458 1568 465 sw
tri 2020 458 2027 465 se
rect 2027 458 2033 492
rect 2067 458 2073 492
rect 3051 852 3097 864
rect 3051 818 3057 852
rect 3091 818 3097 852
rect 3051 780 3097 818
rect 3051 746 3057 780
rect 3091 746 3097 780
rect 3051 708 3097 746
rect 3051 674 3057 708
rect 3091 674 3097 708
rect 3051 636 3097 674
rect 3051 602 3057 636
rect 3091 602 3097 636
rect 3051 564 3097 602
rect 3051 530 3057 564
rect 3091 530 3097 564
rect 3051 492 3097 530
tri 2073 458 2080 465 sw
tri 2532 458 2539 465 se
rect 1561 440 1568 458
tri 1568 440 1586 458 sw
tri 2002 440 2020 458 se
rect 2020 440 2080 458
tri 2080 440 2098 458 sw
tri 2514 440 2532 458 se
rect 2532 440 2539 458
tri 2585 458 2592 465 sw
tri 3044 458 3051 465 se
rect 3051 458 3057 492
rect 3091 458 3097 492
rect 3307 855 3313 889
rect 3347 855 3353 889
rect 3307 817 3353 855
rect 3307 783 3313 817
rect 3347 783 3353 817
rect 3307 745 3353 783
rect 3307 711 3313 745
rect 3347 711 3353 745
rect 3307 673 3353 711
rect 3307 639 3313 673
rect 3347 639 3353 673
rect 3307 601 3353 639
rect 3307 567 3313 601
rect 3347 567 3353 601
rect 3307 529 3353 567
rect 3307 495 3313 529
rect 3347 495 3353 529
rect 3307 483 3353 495
rect 3820 1026 3864 1027
rect 3819 961 3865 1025
rect 3819 927 3825 961
rect 3859 927 3865 961
rect 3819 889 3865 927
rect 3819 855 3825 889
rect 3859 855 3865 889
rect 3819 817 3865 855
rect 3819 783 3825 817
rect 3859 783 3865 817
rect 3819 745 3865 783
rect 3819 711 3825 745
rect 3859 711 3865 745
rect 3819 673 3865 711
rect 4753 1032 4799 1070
tri 4799 1067 4824 1092 nw
tri 5040 1067 5065 1092 ne
rect 4753 998 4759 1032
rect 4793 998 4799 1032
rect 4753 960 4799 998
rect 6944 1065 7620 1096
tri 7620 1071 7645 1096 nw
tri 7901 1071 7926 1096 ne
rect 7926 1065 8068 1096
rect 6944 1000 7574 1065
rect 6944 975 6972 1000
tri 6972 975 6997 1000 nw
tri 7549 975 7574 1000 ne
rect 7759 1037 7889 1043
rect 7811 1003 7843 1037
rect 7877 1003 7889 1037
rect 7811 997 7889 1003
rect 4753 926 4759 960
rect 4793 926 4799 960
rect 4753 888 4799 926
rect 7759 973 7811 985
rect 7759 915 7811 921
tri 7811 919 7889 997 nw
rect 4753 854 4759 888
rect 4793 854 4799 888
rect 4753 816 4799 854
rect 4753 782 4759 816
rect 4793 782 4799 816
rect 4753 744 4799 782
rect 7667 895 7719 901
rect 7667 831 7719 843
rect 7667 773 7719 779
tri 7667 770 7670 773 ne
tri 7716 770 7719 773 nw
rect 4753 710 4759 744
rect 4793 710 4799 744
rect 4753 698 4799 710
rect 3819 639 3825 673
rect 3859 639 3865 673
tri 4643 670 4668 695 sw
tri 4884 670 4909 695 se
rect 3819 601 3865 639
rect 3819 567 3825 601
rect 3859 567 3865 601
rect 3819 529 3865 567
rect 3819 495 3825 529
rect 3859 495 3865 529
rect 3819 483 3865 495
rect 4597 468 4909 670
rect 2585 440 2592 458
tri 2592 440 2610 458 sw
tri 3026 440 3044 458 se
rect 3044 440 3097 458
tri 3097 440 3122 465 sw
tri 3538 440 3563 465 se
tri 3609 440 3634 465 sw
tri 4050 440 4075 465 se
tri 4121 440 4146 465 sw
tri 4306 440 4331 465 se
tri 4377 440 4402 465 sw
rect -1883 420 5127 440
rect -1883 368 -1510 420
rect -1458 368 -1440 420
rect -1388 368 -1370 420
rect -1318 368 -1301 420
rect -1249 368 -1232 420
rect -1180 368 -1163 420
rect -1111 368 -1094 420
rect -1042 368 -1025 420
rect -973 368 -956 420
rect -904 368 -887 420
rect -835 368 -818 420
rect -766 368 -749 420
rect -697 386 2033 420
rect 2067 386 3057 420
rect 3091 386 5127 420
rect -697 368 5127 386
rect -1883 356 5127 368
rect -1883 344 -1510 356
rect -2137 321 -2021 337
rect -2406 246 -2405 275
tri -2405 246 -2376 275 sw
rect -2249 269 -2137 275
rect -2085 269 -2073 321
rect -2249 263 -2021 269
rect -1929 304 -1510 344
rect -1458 304 -1440 356
rect -1388 304 -1370 356
rect -1318 304 -1301 356
rect -1249 304 -1232 356
rect -1180 304 -1163 356
rect -1111 304 -1094 356
rect -1042 304 -1025 356
rect -973 304 -956 356
rect -904 304 -887 356
rect -835 304 -818 356
rect -766 304 -749 356
rect -697 304 5127 356
rect -1929 292 5127 304
rect -1929 280 -1510 292
rect -1458 280 -1440 292
rect -1388 280 -1370 292
rect -1318 280 -1301 292
rect -1249 280 -1232 292
rect -1180 280 -1163 292
rect -1111 280 -1094 292
rect -1042 280 -1025 292
rect -973 280 -956 292
rect -904 280 -887 292
rect -835 280 -818 292
rect -766 280 -749 292
rect -697 286 5127 292
tri 5127 286 5143 302 sw
rect -697 280 5143 286
rect -1929 246 -1917 280
rect -1883 246 -1845 280
rect -1811 246 -1773 280
rect -1739 246 -1701 280
rect -1667 246 -1629 280
rect -1595 246 -1557 280
rect -1523 246 -1510 280
rect -1451 246 -1440 280
rect -1379 246 -1370 280
rect -1307 246 -1301 280
rect -1235 246 -1232 280
rect -766 246 -765 280
rect -697 246 -693 280
rect -659 246 -621 280
rect -587 246 -549 280
rect -515 246 -477 280
rect -443 246 -405 280
rect -371 246 -333 280
rect -299 246 -261 280
rect -227 246 -189 280
rect -155 246 -117 280
rect -83 246 -45 280
rect -11 246 27 280
rect 61 246 99 280
rect 133 246 171 280
rect 205 246 243 280
rect 277 246 315 280
rect 349 246 387 280
rect 421 246 460 280
rect 494 246 533 280
rect 567 246 606 280
rect 640 246 679 280
rect 713 246 752 280
rect 786 246 825 280
rect 859 246 898 280
rect 932 246 971 280
rect 1005 246 1044 280
rect 1078 246 1117 280
rect 1151 246 1190 280
rect 1224 246 1263 280
rect 1297 246 1336 280
rect 1370 246 1409 280
rect 1443 246 1482 280
rect 1516 246 1555 280
rect 1589 246 1628 280
rect 1662 246 1701 280
rect 1735 246 1774 280
rect 1808 246 1847 280
rect 1881 246 1920 280
rect 1954 246 1993 280
rect 2027 246 2066 280
rect 2100 246 2139 280
rect 2173 246 2212 280
rect 2246 246 2285 280
rect 2319 246 2358 280
rect 2392 246 2431 280
rect 2465 246 2504 280
rect 2538 246 2577 280
rect 2611 246 2650 280
rect 2684 246 2723 280
rect 2757 246 2796 280
rect 2830 246 2869 280
rect 2903 246 2942 280
rect 2976 246 3015 280
rect 3049 246 3088 280
rect 3122 246 3161 280
rect 3195 246 3234 280
rect 3268 246 3307 280
rect 3341 246 3380 280
rect 3414 246 3453 280
rect 3487 246 3526 280
rect 3560 246 3599 280
rect 3633 246 3672 280
rect 3706 246 3745 280
rect 3779 246 3818 280
rect 3852 246 3891 280
rect 3925 246 3964 280
rect 3998 246 4037 280
rect 4071 246 4110 280
rect 4144 246 4183 280
rect 4217 246 4256 280
rect 4290 246 4329 280
rect 4363 246 4402 280
rect 4436 246 4475 280
rect 4509 246 4548 280
rect 4582 246 4621 280
rect 4655 246 4694 280
rect 4728 246 4767 280
rect 4801 246 4840 280
rect 4874 246 4913 280
rect 4947 246 4986 280
rect 5020 246 5059 280
rect 5093 246 5143 280
rect -2406 240 -2376 246
tri -2376 240 -2370 246 sw
rect -1929 240 -1510 246
rect -1458 240 -1440 246
rect -1388 240 -1370 246
rect -1318 240 -1301 246
rect -1249 240 -1232 246
rect -1180 240 -1163 246
rect -1111 240 -1094 246
rect -1042 240 -1025 246
rect -973 240 -956 246
rect -904 240 -887 246
rect -835 240 -818 246
rect -766 240 -749 246
rect -697 240 5143 246
rect -2406 212 -2370 240
tri -2370 212 -2342 240 sw
rect -2406 49 4877 212
rect -2406 32 -2184 49
tri -2184 32 -2167 49 nw
tri -1980 32 -1963 49 ne
rect -1963 32 4877 49
rect 6944 157 6972 182
tri 6972 157 6997 182 sw
tri 7549 157 7574 182 se
tri -2143 4 -2138 9 se
rect -2138 4 -2131 9
rect -2902 3 -2299 4
tri -2299 3 -2298 4 sw
tri -2144 3 -2143 4 se
rect -2143 3 -2131 4
rect -2902 -3 -2298 3
tri -2298 -3 -2292 3 sw
rect -2206 -3 -2131 3
rect -2902 -28 -2292 -3
tri -2292 -28 -2267 -3 sw
rect -2902 -37 -2267 -28
tri -2267 -37 -2258 -28 sw
rect -2206 -37 -2194 -3
rect -2160 -37 -2131 -3
rect -2902 -43 -2258 -37
tri -2258 -43 -2252 -37 sw
rect -2206 -43 -2131 -37
rect -2079 -43 -2066 9
rect -2014 3 -2008 9
tri -2008 3 -2003 8 sw
rect -2014 -3 5017 3
rect -2014 -37 -1978 -3
rect -1944 -37 -1906 -3
rect -1872 -37 -1834 -3
rect -1800 -37 -1762 -3
rect -1728 -37 -1690 -3
rect -1656 -37 -1618 -3
rect -1584 -37 -1546 -3
rect -1512 -37 -1474 -3
rect -1440 -37 -1402 -3
rect -1368 -37 -1330 -3
rect -1296 -37 -1258 -3
rect -1224 -37 -1186 -3
rect -1152 -37 -1114 -3
rect -1080 -37 -1042 -3
rect -1008 -37 -970 -3
rect -936 -37 -898 -3
rect -864 -37 -826 -3
rect -792 -37 -754 -3
rect -720 -37 -682 -3
rect -648 -37 -610 -3
rect -576 -37 -538 -3
rect -504 -37 -466 -3
rect -432 -37 -394 -3
rect -360 -37 -322 -3
rect -288 -37 -250 -3
rect -216 -37 -178 -3
rect -144 -37 -106 -3
rect -72 -37 -34 -3
rect 0 -37 38 -3
rect 72 -37 110 -3
rect 144 -37 182 -3
rect 216 -37 254 -3
rect 288 -37 326 -3
rect 360 -37 398 -3
rect 432 -37 470 -3
rect 504 -37 542 -3
rect 576 -37 614 -3
rect 648 -37 686 -3
rect 720 -37 758 -3
rect 792 -37 830 -3
rect 864 -37 902 -3
rect 936 -37 974 -3
rect 1008 -37 1046 -3
rect 1080 -37 1118 -3
rect 1152 -37 1190 -3
rect 1224 -37 1262 -3
rect 1296 -37 1334 -3
rect 1368 -37 1406 -3
rect 1440 -37 1478 -3
rect 1512 -37 1550 -3
rect 1584 -37 1622 -3
rect 1656 -37 1694 -3
rect 1728 -37 1766 -3
rect 1800 -37 1838 -3
rect 1872 -37 1910 -3
rect 1944 -37 1982 -3
rect 2016 -37 2054 -3
rect 2088 -37 2126 -3
rect 2160 -37 2198 -3
rect 2232 -37 2270 -3
rect 2304 -37 2343 -3
rect 2377 -37 2416 -3
rect 2450 -37 2489 -3
rect 2523 -37 2562 -3
rect 2596 -37 2635 -3
rect 2669 -37 2708 -3
rect 2742 -37 2781 -3
rect 2815 -37 2854 -3
rect 2888 -37 2927 -3
rect 2961 -37 3000 -3
rect 3034 -37 3073 -3
rect 3107 -37 3146 -3
rect 3180 -37 3219 -3
rect 3253 -37 3292 -3
rect 3326 -37 3365 -3
rect 3399 -37 3438 -3
rect 3472 -37 3511 -3
rect 3545 -37 3584 -3
rect 3618 -37 3657 -3
rect 3691 -37 3730 -3
rect 3764 -37 3803 -3
rect 3837 -37 3876 -3
rect 3910 -37 3949 -3
rect 3983 -37 4022 -3
rect 4056 -37 4095 -3
rect 4129 -37 4168 -3
rect 4202 -37 4241 -3
rect 4275 -37 4314 -3
rect 4348 -37 4387 -3
rect 4421 -37 4460 -3
rect 4494 -37 4533 -3
rect 4567 -37 4606 -3
rect 4640 -37 4679 -3
rect 4713 -37 4752 -3
rect 4786 -37 4825 -3
rect 4859 -37 4898 -3
rect 4932 -37 4971 -3
rect 5005 -37 5017 -3
rect -2014 -43 5017 -37
rect 6944 -43 7574 157
rect -2902 -48 -2252 -43
tri -2321 -88 -2281 -48 ne
rect -2281 -68 -2252 -48
tri -2252 -68 -2227 -43 sw
tri 7478 -68 7503 -43 ne
rect 7503 -68 7574 -43
rect -2281 -88 -2227 -68
tri -2227 -88 -2207 -68 sw
tri 7503 -88 7523 -68 ne
rect 7523 -73 7574 -68
tri 7620 -73 7625 -68 sw
tri 7921 -73 7926 -68 se
rect 7926 -73 8022 1065
rect 7523 -88 7625 -73
tri 7625 -88 7640 -73 sw
tri 7906 -88 7921 -73 se
rect 7921 -88 8068 -73
rect -2902 -140 -2829 -88
rect -2745 -99 -2321 -88
tri -2321 -99 -2310 -88 sw
tri -2281 -99 -2270 -88 ne
rect -2270 -93 -2207 -88
tri -2207 -93 -2202 -88 sw
tri 7523 -93 7528 -88 ne
rect 7528 -93 7640 -88
tri 7640 -93 7645 -88 sw
tri 7901 -93 7906 -88 se
rect 7906 -93 8068 -88
rect -2270 -99 -2202 -93
tri -2202 -99 -2196 -93 sw
tri 7528 -99 7534 -93 ne
rect 7534 -99 8068 -93
rect -2745 -102 -2310 -99
tri -2310 -102 -2307 -99 sw
tri -2270 -102 -2267 -99 ne
rect -2267 -102 -2196 -99
tri -2196 -102 -2193 -99 sw
tri 7534 -102 7537 -99 ne
rect 7537 -102 7586 -99
rect -2745 -120 -2307 -102
tri -2307 -120 -2289 -102 sw
tri -2267 -120 -2249 -102 ne
rect -2249 -120 5127 -102
rect -2745 -133 -2289 -120
tri -2289 -133 -2276 -120 sw
tri -2249 -133 -2236 -120 ne
rect -2236 -133 5127 -120
tri 7537 -133 7568 -102 ne
rect 7568 -133 7586 -102
rect 7620 -133 7659 -99
rect 7693 -133 7732 -99
rect 7766 -133 7805 -99
rect 7839 -133 7878 -99
rect 7912 -133 7950 -99
rect 7984 -133 8022 -99
rect 8056 -133 8068 -99
rect -2745 -139 -2276 -133
tri -2276 -139 -2270 -133 sw
tri -2236 -139 -2230 -133 ne
rect -2230 -139 5127 -133
tri 7568 -139 7574 -133 ne
rect 7574 -139 8068 -133
rect -2745 -140 -2270 -139
tri -2270 -140 -2269 -139 sw
tri -2230 -140 -2229 -139 ne
rect -2229 -140 5127 -139
tri -2745 -165 -2720 -140 ne
rect -2720 -165 -2590 -140
tri -2590 -165 -2565 -140 nw
tri -2343 -165 -2318 -140 ne
rect -2318 -154 -2269 -140
tri -2269 -154 -2255 -140 sw
tri -2229 -154 -2215 -140 ne
rect -2215 -154 5127 -140
rect -2318 -165 -2255 -154
tri -2318 -194 -2289 -165 ne
rect -2289 -194 -2255 -165
tri -2255 -194 -2215 -154 sw
tri -2289 -203 -2280 -194 ne
rect -2280 -203 5127 -194
tri -2745 -228 -2720 -203 se
rect -2720 -228 -2590 -203
tri -2590 -228 -2565 -203 sw
tri -2280 -228 -2255 -203 ne
rect -2255 -228 5127 -203
rect -2902 -246 -2301 -228
tri -2301 -246 -2283 -228 sw
tri -2255 -246 -2237 -228 ne
rect -2237 -246 5127 -228
rect -2902 -254 -2283 -246
tri -2283 -254 -2275 -246 sw
rect -2902 -280 -2275 -254
tri -2323 -308 -2295 -280 ne
rect -2295 -308 -2275 -280
rect -2902 -328 -2335 -308
tri -2335 -328 -2315 -308 sw
tri -2295 -328 -2275 -308 ne
tri -2275 -328 -2201 -254 sw
rect -2902 -334 -2315 -328
tri -2315 -334 -2309 -328 sw
tri -2275 -334 -2269 -328 ne
rect -2269 -334 5127 -328
rect -2902 -360 -2309 -334
tri -2357 -408 -2309 -360 ne
tri -2309 -368 -2275 -334 sw
tri -2269 -368 -2235 -334 ne
rect -2235 -368 5127 -334
rect -2309 -380 -2275 -368
tri -2275 -380 -2263 -368 sw
tri -2235 -380 -2223 -368 ne
rect -2223 -380 5127 -368
rect -2309 -408 -2263 -380
tri -2263 -408 -2235 -380 sw
tri -2309 -460 -2257 -408 ne
rect -2257 -460 5127 -408
rect -2800 -626 -2398 -595
tri -2800 -636 -2790 -626 ne
rect -2790 -636 -2398 -626
<< rmetal1 >>
rect -179 1191 -177 1192
rect -141 1191 -139 1192
rect -179 1093 -178 1191
rect -140 1093 -139 1191
rect -179 1092 -177 1093
rect -141 1092 -139 1093
rect 1842 1063 1844 1064
rect 1842 965 1843 1063
rect 1842 964 1844 965
rect 1880 1063 1882 1064
rect 1881 965 1882 1063
rect 1880 964 1882 965
rect 2866 1063 2868 1064
rect 2866 965 2867 1063
rect 2866 964 2868 965
rect 2904 1063 2906 1064
rect 2905 965 2906 1063
rect 3307 1064 3353 1065
rect 3307 1063 3308 1064
rect 3352 1063 3353 1064
rect 3819 1064 3865 1065
rect 3819 1063 3820 1064
rect 3864 1063 3865 1064
rect 2904 964 2906 965
rect 3307 1026 3308 1027
rect 3352 1026 3353 1027
rect 3307 1025 3353 1026
rect 3819 1026 3820 1027
rect 3864 1026 3865 1027
rect 3819 1025 3865 1026
<< via1 >>
rect -2131 1815 -2079 1867
rect -2066 1815 -2014 1867
rect -2131 1751 -2127 1803
rect -2127 1751 -2079 1803
rect -2066 1751 -2014 1803
rect -2298 1688 -2246 1740
rect -2298 1622 -2246 1674
rect 7759 1604 7811 1656
rect -2137 1466 -2021 1582
rect 7597 1536 7649 1588
rect 7661 1536 7713 1588
rect 7759 1540 7811 1592
rect -1510 1508 -1458 1514
rect -1440 1508 -1388 1514
rect -1370 1508 -1318 1514
rect -1301 1508 -1249 1514
rect -1510 1474 -1485 1508
rect -1485 1474 -1458 1508
rect -1440 1474 -1413 1508
rect -1413 1474 -1388 1508
rect -1370 1474 -1341 1508
rect -1341 1474 -1318 1508
rect -1301 1474 -1269 1508
rect -1269 1474 -1249 1508
rect -1510 1462 -1458 1474
rect -1440 1462 -1388 1474
rect -1370 1462 -1318 1474
rect -1301 1462 -1249 1474
rect -1232 1508 -1180 1514
rect -1232 1474 -1231 1508
rect -1231 1474 -1197 1508
rect -1197 1474 -1180 1508
rect -1232 1462 -1180 1474
rect -1163 1508 -1111 1514
rect -1163 1474 -1159 1508
rect -1159 1474 -1125 1508
rect -1125 1474 -1111 1508
rect -1163 1462 -1111 1474
rect -1094 1508 -1042 1514
rect -1094 1474 -1087 1508
rect -1087 1474 -1053 1508
rect -1053 1474 -1042 1508
rect -1094 1462 -1042 1474
rect -1025 1508 -973 1514
rect -1025 1474 -1015 1508
rect -1015 1474 -981 1508
rect -981 1474 -973 1508
rect -1025 1462 -973 1474
rect -956 1508 -904 1514
rect -956 1474 -943 1508
rect -943 1474 -909 1508
rect -909 1474 -904 1508
rect -956 1462 -904 1474
rect -887 1508 -835 1514
rect -887 1474 -871 1508
rect -871 1474 -837 1508
rect -837 1474 -835 1508
rect -887 1462 -835 1474
rect -818 1508 -766 1514
rect -749 1508 -697 1514
rect -818 1474 -799 1508
rect -799 1474 -766 1508
rect -749 1474 -727 1508
rect -727 1474 -697 1508
rect -818 1462 -766 1474
rect -749 1462 -697 1474
rect -2450 1183 -2398 1235
rect -2384 1183 -2332 1235
rect -2137 1208 -2085 1260
rect -2073 1208 -2021 1260
rect -2137 1141 -2085 1193
rect -2073 1141 -2021 1193
rect -2450 1069 -2398 1121
rect -2384 1069 -2332 1121
rect -2137 1074 -2085 1126
rect -2073 1074 -2021 1126
rect -2137 1007 -2085 1059
rect -2073 1007 -2021 1059
rect -2450 944 -2398 996
rect -2384 944 -2332 996
rect -2137 940 -2085 992
rect -2073 940 -2021 992
rect -2137 873 -2085 925
rect -2073 873 -2021 925
rect -2137 806 -2085 858
rect -2073 806 -2021 858
rect -2137 739 -2085 791
rect -2073 739 -2021 791
rect -2137 672 -2085 724
rect -2073 672 -2021 724
rect -2137 605 -2085 657
rect -2073 605 -2021 657
rect -2137 538 -2085 590
rect -2073 538 -2021 590
rect -2137 471 -2085 523
rect -2073 471 -2021 523
rect -2137 404 -2085 456
rect -2073 404 -2021 456
rect -2137 337 -2085 389
rect -2073 337 -2021 389
rect 7759 1003 7771 1037
rect 7771 1003 7805 1037
rect 7805 1003 7811 1037
rect 7759 985 7811 1003
rect 7759 921 7811 973
rect 7667 843 7719 895
rect 7667 779 7719 831
rect -1510 368 -1458 420
rect -1440 368 -1388 420
rect -1370 368 -1318 420
rect -1301 368 -1249 420
rect -1232 368 -1180 420
rect -1163 368 -1111 420
rect -1094 368 -1042 420
rect -1025 368 -973 420
rect -956 368 -904 420
rect -887 368 -835 420
rect -818 368 -766 420
rect -749 368 -697 420
rect -2137 269 -2085 321
rect -2073 269 -2021 321
rect -1510 304 -1458 356
rect -1440 304 -1388 356
rect -1370 304 -1318 356
rect -1301 304 -1249 356
rect -1232 304 -1180 356
rect -1163 304 -1111 356
rect -1094 304 -1042 356
rect -1025 304 -973 356
rect -956 304 -904 356
rect -887 304 -835 356
rect -818 304 -766 356
rect -749 304 -697 356
rect -1510 280 -1458 292
rect -1440 280 -1388 292
rect -1370 280 -1318 292
rect -1301 280 -1249 292
rect -1232 280 -1180 292
rect -1163 280 -1111 292
rect -1094 280 -1042 292
rect -1025 280 -973 292
rect -956 280 -904 292
rect -887 280 -835 292
rect -818 280 -766 292
rect -749 280 -697 292
rect -1510 246 -1485 280
rect -1485 246 -1458 280
rect -1440 246 -1413 280
rect -1413 246 -1388 280
rect -1370 246 -1341 280
rect -1341 246 -1318 280
rect -1301 246 -1269 280
rect -1269 246 -1249 280
rect -1232 246 -1197 280
rect -1197 246 -1180 280
rect -1163 246 -1125 280
rect -1125 246 -1111 280
rect -1094 246 -1091 280
rect -1091 246 -1053 280
rect -1053 246 -1042 280
rect -1025 246 -1019 280
rect -1019 246 -981 280
rect -981 246 -973 280
rect -956 246 -947 280
rect -947 246 -909 280
rect -909 246 -904 280
rect -887 246 -875 280
rect -875 246 -837 280
rect -837 246 -835 280
rect -818 246 -803 280
rect -803 246 -766 280
rect -749 246 -731 280
rect -731 246 -697 280
rect -1510 240 -1458 246
rect -1440 240 -1388 246
rect -1370 240 -1318 246
rect -1301 240 -1249 246
rect -1232 240 -1180 246
rect -1163 240 -1111 246
rect -1094 240 -1042 246
rect -1025 240 -973 246
rect -956 240 -904 246
rect -887 240 -835 246
rect -818 240 -766 246
rect -749 240 -697 246
rect -2131 -3 -2079 9
rect -2131 -37 -2122 -3
rect -2122 -37 -2088 -3
rect -2088 -37 -2079 -3
rect -2131 -43 -2079 -37
rect -2066 -3 -2014 9
rect -2066 -37 -2050 -3
rect -2050 -37 -2016 -3
rect -2016 -37 -2014 -3
rect -2066 -43 -2014 -37
<< metal2 >>
rect -3052 1815 -2732 1867
tri -2732 1815 -2680 1867 sw
rect -3052 1803 -2680 1815
tri -2680 1803 -2668 1815 sw
rect -3052 1751 -2668 1803
tri -2668 1751 -2616 1803 sw
rect -3052 1740 -2616 1751
tri -2616 1740 -2605 1751 sw
rect -3052 1715 -2605 1740
tri -2605 1715 -2580 1740 sw
rect -3052 1599 -2580 1715
rect -3052 1592 -2587 1599
tri -2587 1592 -2580 1599 nw
rect -3052 1588 -2591 1592
tri -2591 1588 -2587 1592 nw
rect -3052 1582 -2597 1588
tri -2597 1582 -2591 1588 nw
rect -3052 1466 -2713 1582
tri -2713 1466 -2597 1582 nw
rect -3052 1462 -2717 1466
tri -2717 1462 -2713 1466 nw
rect -3052 -223 -2732 1462
tri -2732 1447 -2717 1462 nw
tri -2403 1235 -2378 1260 se
rect -2378 1235 -2326 1867
rect -2456 1183 -2450 1235
rect -2398 1183 -2384 1235
rect -2332 1183 -2326 1235
rect -2298 1740 -2246 1867
rect -2298 1674 -2246 1688
tri -2303 1141 -2298 1146 se
rect -2298 1141 -2246 1622
tri -2318 1126 -2303 1141 se
rect -2303 1126 -2246 1141
tri -2323 1121 -2318 1126 se
rect -2318 1121 -2246 1126
rect -2456 1069 -2450 1121
rect -2398 1069 -2384 1121
rect -2332 1069 -2246 1121
tri -2232 1007 -2218 1021 se
rect -2218 1007 -2166 1867
tri -2243 996 -2232 1007 se
rect -2232 996 -2166 1007
rect -2456 944 -2450 996
rect -2398 944 -2384 996
rect -2332 944 -2166 996
rect -2137 1815 -2131 1867
rect -2079 1815 -2066 1867
rect -2014 1815 -2008 1867
rect -2137 1803 -2008 1815
rect -2137 1751 -2131 1803
rect -2079 1751 -2066 1803
rect -2014 1751 -2008 1803
rect -2137 1582 -2008 1751
rect -2021 1466 -2008 1582
rect -2137 1260 -2008 1466
rect -2085 1208 -2073 1260
rect -2021 1208 -2008 1260
rect -2137 1193 -2008 1208
rect -2085 1141 -2073 1193
rect -2021 1141 -2008 1193
rect -2137 1126 -2008 1141
rect -2085 1074 -2073 1126
rect -2021 1074 -2008 1126
rect -2137 1059 -2008 1074
rect -2085 1007 -2073 1059
rect -2021 1007 -2008 1059
rect -2137 992 -2008 1007
rect -2085 940 -2073 992
rect -2021 940 -2008 992
rect -2137 925 -2008 940
rect -2085 873 -2073 925
rect -2021 873 -2008 925
rect -2137 858 -2008 873
rect -2085 806 -2073 858
rect -2021 806 -2008 858
rect -2137 791 -2008 806
rect -2085 739 -2073 791
rect -2021 739 -2008 791
rect -2137 724 -2008 739
rect -2085 672 -2073 724
rect -2021 672 -2008 724
rect -2137 657 -2008 672
rect -2085 605 -2073 657
rect -2021 605 -2008 657
rect -2137 590 -2008 605
rect -2085 538 -2073 590
rect -2021 538 -2008 590
rect -2137 523 -2008 538
rect -2085 471 -2073 523
rect -2021 471 -2008 523
rect -2137 456 -2008 471
rect -2085 404 -2073 456
rect -2021 404 -2008 456
rect -2137 389 -2008 404
rect -2085 337 -2073 389
rect -2021 337 -2008 389
rect -2137 321 -2008 337
rect -2085 269 -2073 321
rect -2021 269 -2008 321
rect -2662 -520 -2406 32
rect -2137 9 -2008 269
rect -2137 -43 -2131 9
rect -2079 -43 -2066 9
rect -2014 -43 -2008 9
tri -2241 -520 -2137 -416 se
rect -2137 -520 -2008 -43
rect -1516 1514 -691 1867
rect -1516 1462 -1510 1514
rect -1458 1462 -1440 1514
rect -1388 1462 -1370 1514
rect -1318 1462 -1301 1514
rect -1249 1462 -1232 1514
rect -1180 1462 -1163 1514
rect -1111 1462 -1094 1514
rect -1042 1462 -1025 1514
rect -973 1462 -956 1514
rect -904 1462 -887 1514
rect -835 1462 -818 1514
rect -766 1462 -749 1514
rect -697 1462 -691 1514
rect -1516 420 -691 1462
rect -1516 368 -1510 420
rect -1458 368 -1440 420
rect -1388 368 -1370 420
rect -1318 368 -1301 420
rect -1249 368 -1232 420
rect -1180 368 -1163 420
rect -1111 368 -1094 420
rect -1042 368 -1025 420
rect -973 368 -956 420
rect -904 368 -887 420
rect -835 368 -818 420
rect -766 368 -749 420
rect -697 368 -691 420
rect -1516 356 -691 368
rect -1516 304 -1510 356
rect -1458 304 -1440 356
rect -1388 304 -1370 356
rect -1318 304 -1301 356
rect -1249 304 -1232 356
rect -1180 304 -1163 356
rect -1111 304 -1094 356
rect -1042 304 -1025 356
rect -973 304 -956 356
rect -904 304 -887 356
rect -835 304 -818 356
rect -766 304 -749 356
rect -697 304 -691 356
rect -1516 292 -691 304
rect -1516 240 -1510 292
rect -1458 240 -1440 292
rect -1388 240 -1370 292
rect -1318 240 -1301 292
rect -1249 240 -1232 292
rect -1180 240 -1163 292
rect -1111 240 -1094 292
rect -1042 240 -1025 292
rect -973 240 -956 292
rect -904 240 -887 292
rect -835 240 -818 292
rect -766 240 -749 292
rect -697 240 -691 292
tri -2008 -520 -1649 -161 sw
rect -1516 -223 -691 240
rect 1254 -519 1446 1865
rect 1993 -519 2123 1865
rect 2689 -519 2881 1865
rect 3177 -519 3229 1898
rect 3269 -519 3321 1898
rect 3870 -519 4062 1865
rect 4392 -519 4584 1865
rect 7759 1656 7811 1662
rect 7759 1592 7811 1604
rect 7591 1536 7597 1588
rect 7649 1536 7661 1588
rect 7713 1536 7719 1588
tri 7642 1534 7644 1536 ne
rect 7644 1534 7719 1536
tri 7644 1511 7667 1534 ne
rect 7667 895 7719 1534
rect 7759 1037 7811 1540
rect 7759 973 7811 985
rect 7759 915 7811 921
rect 7667 831 7719 843
rect 7667 773 7719 779
rect 4685 212 4877 468
tri -2350 -629 -2241 -520 se
rect -2241 -629 -1649 -520
tri -1649 -629 -1540 -520 sw
rect -2350 -657 -1540 -629
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 -1352 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 -1096 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 -840 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 -584 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 -328 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 -72 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 184 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 440 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 696 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 952 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 1208 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 1464 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 1720 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 1976 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform -1 0 2232 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform -1 0 2488 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform -1 0 2744 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform -1 0 3000 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform -1 0 3256 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform -1 0 3512 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform -1 0 3768 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform -1 0 4024 0 -1 1340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform -1 0 -1604 0 -1 1627
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform -1 0 -1604 0 -1 1426
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 4954 0 -1 1426
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 7771 0 -1 1037
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 4954 0 -1 1582
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform 0 -1 -1517 -1 0 1140
box -12 -6 766 40
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_1
timestamp 1707688321
transform 0 1 -1807 -1 0 1254
box -12 -6 766 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1707688321
transform 0 -1 1043 -1 0 924
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1707688321
transform 0 -1 531 -1 0 924
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_2
timestamp 1707688321
transform 0 -1 1555 -1 0 924
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_3
timestamp 1707688321
transform 0 -1 2835 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_4
timestamp 1707688321
transform 0 -1 2579 -1 0 924
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_5
timestamp 1707688321
transform 0 -1 1811 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_6
timestamp 1707688321
transform 0 -1 275 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_7
timestamp 1707688321
transform 0 -1 787 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_8
timestamp 1707688321
transform 0 -1 1299 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_9
timestamp 1707688321
transform 0 -1 2323 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_10
timestamp 1707688321
transform 0 -1 4637 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_11
timestamp 1707688321
transform 0 -1 4949 -1 0 1018
box -12 -6 550 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1707688321
transform 0 -1 -1005 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_1
timestamp 1707688321
transform 0 -1 19 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_2
timestamp 1707688321
transform 0 -1 -493 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_3
timestamp 1707688321
transform 0 -1 4371 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_4
timestamp 1707688321
transform 0 -1 4115 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_5
timestamp 1707688321
transform 0 -1 3603 -1 0 996
box -12 -6 622 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1707688321
transform 0 -1 5105 -1 0 1162
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_1
timestamp 1707688321
transform 0 -1 4479 -1 0 1162
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_2
timestamp 1707688321
transform 0 -1 -749 1 0 480
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_3
timestamp 1707688321
transform 0 -1 -237 1 0 480
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_4
timestamp 1707688321
transform 0 -1 -1261 1 0 480
box -12 -6 694 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform 0 -1 7614 1 0 -61
box -12 -6 1126 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_1
timestamp 1707688321
transform 0 -1 8062 1 0 -61
box -12 -6 1126 40
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1707688321
transform 0 -1 2067 -1 0 852
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_1
timestamp 1707688321
transform 0 -1 3091 -1 0 852
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_2
timestamp 1707688321
transform 0 -1 3347 -1 0 961
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_3
timestamp 1707688321
transform 0 -1 3859 -1 0 961
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_4
timestamp 1707688321
transform 0 -1 4793 -1 0 1176
box 0 0 1 1
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1707688321
transform 0 -1 7710 -1 0 889
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1707688321
transform 0 -1 7966 -1 0 889
box -12 -6 910 40
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 5027 0 -1 1260
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform -1 0 4559 0 -1 1260
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1707688321
transform -1 0 4715 0 -1 1260
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1707688321
transform -1 0 4871 0 -1 1260
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1707688321
transform 1 0 -1843 0 1 1474
box 0 0 1 1
use L1M1_CDNS_524688791851040  L1M1_CDNS_524688791851040_0
timestamp 1707688321
transform 0 1 -1923 1 0 344
box -12 -6 1054 40
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1707688321
transform -1 0 -2406 0 -1 -520
box 0 0 256 116
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 1 0 4685 0 1 468
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 1 0 4685 0 1 32
box 0 0 192 180
use M1M2_CDNS_524688791851150  M1M2_CDNS_524688791851150_0
timestamp 1707688321
transform -1 0 -2406 0 1 32
box 0 0 256 244
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 -2790 0 -1 1715
box 0 0 384 116
use nfet_CDNS_52468879185994  nfet_CDNS_52468879185994_0
timestamp 1707688321
transform -1 0 -1562 0 1 354
box -79 -26 279 1026
use nfet_CDNS_52468879185994  nfet_CDNS_52468879185994_1
timestamp 1707688321
transform 1 0 4126 0 1 354
box -79 -26 279 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_0
timestamp 1707688321
transform 1 0 3614 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_1
timestamp 1707688321
transform 1 0 -482 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_2
timestamp 1707688321
transform 1 0 -994 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_3
timestamp 1707688321
transform 1 0 -1506 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_4
timestamp 1707688321
transform 1 0 1566 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_5
timestamp 1707688321
transform 1 0 1054 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_6
timestamp 1707688321
transform 1 0 542 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_7
timestamp 1707688321
transform 1 0 30 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_8
timestamp 1707688321
transform 1 0 2590 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_9
timestamp 1707688321
transform 1 0 2078 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_10
timestamp 1707688321
transform 1 0 3102 0 1 354
box -79 -26 535 1026
use nfet_CDNS_524688791851618  nfet_CDNS_524688791851618_0
timestamp 1707688321
transform 1 0 4492 0 1 354
box -79 -26 647 1026
use pfet_CDNS_524688791851619  pfet_CDNS_524688791851619_0
timestamp 1707688321
transform -1 0 7921 0 1 -45
box -119 -66 319 1066
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1707688321
transform 0 1 -2801 -1 0 1675
box 0 0 2270 404
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1707688321
transform 0 -1 3353 1 0 973
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851477  sky130_fd_io__tk_em1o_CDNS_524688791851477_0
timestamp 1707688321
transform 1 0 1790 0 -1 1064
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851477  sky130_fd_io__tk_em1o_CDNS_524688791851477_1
timestamp 1707688321
transform 1 0 2814 0 -1 1064
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1707688321
transform 0 -1 3865 1 0 973
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851617  sky130_fd_io__tk_em1s_CDNS_524688791851617_0
timestamp 1707688321
transform 1 0 -231 0 1 1092
box 0 0 1 1
<< labels >>
flabel comment s -2777 970 -2777 970 3 FreeSans 200 0 0 0 en_hicc
flabel comment s -2777 1209 -2777 1209 3 FreeSans 200 0 0 0 pu_h_n<0>
flabel comment s -2777 1095 -2777 1095 3 FreeSans 200 0 0 0 pu_h_n<1>
flabel comment s -2352 1849 -2352 1849 3 FreeSans 200 270 0 0 pu_h_n<0>
flabel comment s -2273 1851 -2273 1851 3 FreeSans 200 270 0 0 pu_h_n<1>
flabel comment s -2193 1847 -2193 1847 3 FreeSans 200 270 0 0 en_hicc
flabel comment s -1101 1847 -1101 1847 3 FreeSans 200 270 0 0 vgnd
flabel comment s 1343 1847 1343 1847 3 FreeSans 200 270 0 0 vgnd
flabel comment s 2056 1847 2056 1847 3 FreeSans 200 270 0 0 vcc_io
flabel comment s 2782 1847 2782 1847 3 FreeSans 200 270 0 0 vgnd
flabel comment s 3962 1847 3962 1847 3 FreeSans 200 270 0 0 vgnd
flabel comment s 4476 1847 4476 1847 3 FreeSans 200 270 0 0 vgnd
flabel comment s 4476 -498 4476 -498 3 FreeSans 200 90 0 0 vgnd
flabel comment s 3962 -498 3962 -498 3 FreeSans 200 90 0 0 vgnd
flabel comment s 2782 -498 2782 -498 3 FreeSans 200 90 0 0 vgnd
flabel comment s 2056 -498 2056 -498 3 FreeSans 200 90 0 0 vcc_io
flabel comment s 1343 -498 1343 -498 3 FreeSans 200 90 0 0 vgnd
flabel comment s -1101 -498 -1101 -498 3 FreeSans 200 90 0 0 vgnd
flabel comment s -2864 -329 -2864 -329 3 FreeSans 200 0 0 0 drvhi_h
flabel comment s -2866 -20 -2866 -20 3 FreeSans 200 0 0 0 slow_h_n
flabel comment s -2864 -251 -2864 -251 3 FreeSans 200 0 0 0 puen_reg_h
flabel comment s -2866 -114 -2866 -114 3 FreeSans 200 0 0 0 vreg_en_h
flabel comment s 3203 1883 3203 1883 3 FreeSans 200 270 0 0 od_h
flabel comment s 3293 1883 3293 1883 3 FreeSans 200 270 0 0 oe_hs_h
flabel comment s 3203 -498 3203 -498 3 FreeSans 200 90 0 0 od_h
flabel comment s 3293 -498 3293 -498 3 FreeSans 200 90 0 0 oe_hs_h
flabel comment s 4205 802 4205 802 0 FreeSans 1000 90 0 0 dummy
flabel metal1 s 6944 975 6972 1200 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 6944 -43 6972 182 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s -2298 1616 -2246 1687 0 FreeSans 200 0 0 0 pu_h_n
port 3 nsew
flabel metal1 s 5067 1294 5143 1346 0 FreeSans 200 0 0 0 refleak_bias
port 4 nsew
flabel metal2 s -2529 -616 -2529 -616 0 FreeSans 200 0 0 0 pad_esd
flabel metal2 s -1516 1820 -691 1867 0 FreeSans 200 0 0 0 vgnd_io
port 5 nsew
flabel metal2 s -3052 -223 -2732 -185 0 FreeSans 200 0 0 0 pad
port 6 nsew
flabel metal2 s -3052 1829 -2732 1867 0 FreeSans 200 0 0 0 pad
port 6 nsew
flabel metal2 s -1516 -43 -691 3 0 FreeSans 200 0 0 0 vgnd_io
port 5 nsew
<< properties >>
string GDS_END 97473514
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97346642
string path -50.225 -0.500 127.200 -0.500 
<< end >>
