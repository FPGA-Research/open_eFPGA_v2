magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 538 414 1177
<< poly >>
rect 114 303 144 819
rect 214 551 244 819
rect 196 535 262 551
rect 196 501 212 535
rect 246 501 262 535
rect 196 485 262 501
rect 96 287 162 303
rect 96 253 112 287
rect 146 253 162 287
rect 96 237 162 253
rect 114 225 144 237
rect 214 225 244 485
<< polycont >>
rect 212 501 246 535
rect 112 253 146 287
<< locali >>
rect 0 1103 378 1137
rect 62 924 96 1103
rect 262 924 296 1103
rect 162 874 196 924
rect 162 840 364 874
rect 212 535 246 551
rect 212 485 246 501
rect 112 287 146 303
rect 112 237 146 253
rect 330 243 364 840
rect 262 209 364 243
rect 262 158 296 209
rect 62 17 96 92
rect 0 -17 378 17
use contact_12  contact_12_0
timestamp 1707688321
transform 1 0 196 0 1 485
box 0 0 1 1
use contact_12  contact_12_1
timestamp 1707688321
transform 1 0 96 0 1 237
box 0 0 1 1
use nmos_m1_w0_740_sactive_dli  nmos_m1_w0_740_sactive_dli_0
timestamp 1707688321
transform 1 0 154 0 1 51
box -26 -26 176 174
use nmos_m1_w0_740_sli_dactive  nmos_m1_w0_740_sli_dactive_0
timestamp 1707688321
transform 1 0 54 0 1 51
box -26 -26 176 174
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_0
timestamp 1707688321
transform 1 0 154 0 1 845
box -59 -54 209 278
use pmos_m1_w1_120_sli_dli  pmos_m1_w1_120_sli_dli_1
timestamp 1707688321
transform 1 0 54 0 1 845
box -59 -54 209 278
<< labels >>
rlabel locali s 347 857 347 857 4 Z
port 3 nsew
rlabel locali s 189 0 189 0 4 gnd
port 5 nsew
rlabel locali s 189 1120 189 1120 4 vdd
port 4 nsew
rlabel locali s 229 518 229 518 4 B
port 2 nsew
rlabel locali s 129 270 129 270 4 A
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 378 1120
string GDS_END 31830
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 29490
<< end >>
