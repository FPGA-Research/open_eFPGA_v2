magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 203
rect 30 -17 64 21
<< locali >>
rect 932 383 1001 417
rect 932 349 998 383
rect 932 336 1001 349
rect 852 315 1001 336
rect 852 302 998 315
rect 27 199 160 265
rect 211 199 361 265
rect 400 199 623 265
rect 679 199 811 265
rect 852 165 895 302
rect 1035 259 1082 325
rect 946 215 1082 259
rect 459 131 1069 165
rect 647 51 681 131
rect 817 51 851 131
rect 1035 51 1069 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 19 299 69 527
rect 119 349 153 493
rect 187 383 253 527
rect 287 349 321 493
rect 357 383 427 527
rect 461 349 495 493
rect 529 383 595 527
rect 822 485 888 493
rect 1035 485 1069 493
rect 629 451 1069 485
rect 717 349 783 417
rect 822 383 888 451
rect 119 315 783 349
rect 1035 359 1069 451
rect 35 131 421 165
rect 35 51 69 131
rect 103 17 169 93
rect 203 51 237 131
rect 271 61 609 95
rect 717 17 783 93
rect 935 17 1001 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 400 199 623 265 6 A1
port 1 nsew signal input
rlabel locali s 211 199 361 265 6 A2
port 2 nsew signal input
rlabel locali s 27 199 160 265 6 A3
port 3 nsew signal input
rlabel locali s 679 199 811 265 6 B1
port 4 nsew signal input
rlabel locali s 946 215 1082 259 6 C1
port 5 nsew signal input
rlabel locali s 1035 259 1082 325 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1103 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1035 51 1069 131 6 Y
port 10 nsew signal output
rlabel locali s 817 51 851 131 6 Y
port 10 nsew signal output
rlabel locali s 647 51 681 131 6 Y
port 10 nsew signal output
rlabel locali s 459 131 1069 165 6 Y
port 10 nsew signal output
rlabel locali s 852 165 895 302 6 Y
port 10 nsew signal output
rlabel locali s 852 302 998 315 6 Y
port 10 nsew signal output
rlabel locali s 852 315 1001 336 6 Y
port 10 nsew signal output
rlabel locali s 932 336 1001 349 6 Y
port 10 nsew signal output
rlabel locali s 932 349 998 383 6 Y
port 10 nsew signal output
rlabel locali s 932 383 1001 417 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3717714
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3707396
<< end >>
