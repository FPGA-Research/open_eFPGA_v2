magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 545 1736 554
rect 0 0 1736 9
<< via2 >>
rect 0 9 1736 545
<< metal3 >>
rect -5 545 1741 550
rect -5 9 0 545
rect 1736 9 1741 545
rect -5 4 1741 9
<< properties >>
string GDS_END 94891838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94881850
<< end >>
