magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 3386
rect 285 0 288 3386
<< via1 >>
rect 3 0 285 3386
<< metal2 >>
rect 0 0 3 3386
rect 285 0 288 3386
<< properties >>
string GDS_END 93718824
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93657636
<< end >>
