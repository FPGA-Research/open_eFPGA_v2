magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 11 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 113 47 143 177
rect 197 47 227 177
rect 281 47 311 177
rect 365 47 395 177
rect 449 47 479 177
rect 533 47 563 177
<< scpmoshvt >>
rect 113 297 143 497
rect 197 297 227 497
rect 281 297 311 497
rect 365 297 395 497
rect 449 297 479 497
rect 533 297 563 497
<< ndiff >>
rect 37 93 113 177
rect 37 59 45 93
rect 79 59 113 93
rect 37 47 113 59
rect 143 101 197 177
rect 143 67 153 101
rect 187 67 197 101
rect 143 47 197 67
rect 227 93 281 177
rect 227 59 237 93
rect 271 59 281 93
rect 227 47 281 59
rect 311 101 365 177
rect 311 67 321 101
rect 355 67 365 101
rect 311 47 365 67
rect 395 93 449 177
rect 395 59 405 93
rect 439 59 449 93
rect 395 47 449 59
rect 479 101 533 177
rect 479 67 489 101
rect 523 67 533 101
rect 479 47 533 67
rect 563 94 617 177
rect 563 60 573 94
rect 607 60 617 94
rect 563 47 617 60
<< pdiff >>
rect 27 485 113 497
rect 27 451 35 485
rect 69 451 113 485
rect 27 417 113 451
rect 27 383 35 417
rect 69 383 113 417
rect 27 349 113 383
rect 27 315 35 349
rect 69 315 113 349
rect 27 297 113 315
rect 143 485 197 497
rect 143 451 153 485
rect 187 451 197 485
rect 143 417 197 451
rect 143 383 153 417
rect 187 383 197 417
rect 143 349 197 383
rect 143 315 153 349
rect 187 315 197 349
rect 143 297 197 315
rect 227 485 281 497
rect 227 451 237 485
rect 271 451 281 485
rect 227 417 281 451
rect 227 383 237 417
rect 271 383 281 417
rect 227 297 281 383
rect 311 485 365 497
rect 311 451 321 485
rect 355 451 365 485
rect 311 417 365 451
rect 311 383 321 417
rect 355 383 365 417
rect 311 349 365 383
rect 311 315 321 349
rect 355 315 365 349
rect 311 297 365 315
rect 395 485 449 497
rect 395 451 405 485
rect 439 451 449 485
rect 395 417 449 451
rect 395 383 405 417
rect 439 383 449 417
rect 395 297 449 383
rect 479 485 533 497
rect 479 451 489 485
rect 523 451 533 485
rect 479 417 533 451
rect 479 383 489 417
rect 523 383 533 417
rect 479 349 533 383
rect 479 315 489 349
rect 523 315 533 349
rect 479 297 533 315
rect 563 485 617 497
rect 563 451 573 485
rect 607 451 617 485
rect 563 297 617 451
<< ndiffc >>
rect 45 59 79 93
rect 153 67 187 101
rect 237 59 271 93
rect 321 67 355 101
rect 405 59 439 93
rect 489 67 523 101
rect 573 60 607 94
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 153 451 187 485
rect 153 383 187 417
rect 153 315 187 349
rect 237 451 271 485
rect 237 383 271 417
rect 321 451 355 485
rect 321 383 355 417
rect 321 315 355 349
rect 405 451 439 485
rect 405 383 439 417
rect 489 451 523 485
rect 489 383 523 417
rect 489 315 523 349
rect 573 451 607 485
<< poly >>
rect 113 497 143 523
rect 197 497 227 523
rect 281 497 311 523
rect 365 497 395 523
rect 449 497 479 523
rect 533 497 563 523
rect 113 265 143 297
rect 197 265 227 297
rect 281 265 311 297
rect 365 265 395 297
rect 449 265 479 297
rect 533 265 563 297
rect 21 249 563 265
rect 21 215 37 249
rect 71 215 305 249
rect 339 215 389 249
rect 423 215 473 249
rect 507 215 563 249
rect 21 199 563 215
rect 113 177 143 199
rect 197 177 227 199
rect 281 177 311 199
rect 365 177 395 199
rect 449 177 479 199
rect 533 177 563 199
rect 113 21 143 47
rect 197 21 227 47
rect 281 21 311 47
rect 365 21 395 47
rect 449 21 479 47
rect 533 21 563 47
<< polycont >>
rect 37 215 71 249
rect 305 215 339 249
rect 389 215 423 249
rect 473 215 507 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 26 485 85 527
rect 26 451 35 485
rect 69 451 85 485
rect 26 417 85 451
rect 26 383 35 417
rect 69 383 85 417
rect 26 349 85 383
rect 26 315 35 349
rect 69 315 85 349
rect 26 299 85 315
rect 137 485 203 493
rect 137 451 153 485
rect 187 451 203 485
rect 137 417 203 451
rect 137 383 153 417
rect 187 383 203 417
rect 137 349 203 383
rect 237 485 271 527
rect 237 417 271 451
rect 237 367 271 383
rect 305 485 371 493
rect 305 451 321 485
rect 355 451 371 485
rect 305 417 371 451
rect 305 383 321 417
rect 355 383 371 417
rect 137 315 153 349
rect 187 333 203 349
rect 305 349 371 383
rect 405 485 439 527
rect 405 417 439 451
rect 405 367 439 383
rect 473 485 539 493
rect 473 451 489 485
rect 523 451 539 485
rect 473 417 539 451
rect 573 485 607 527
rect 573 435 607 451
rect 473 383 489 417
rect 523 383 539 417
rect 305 333 321 349
rect 187 315 321 333
rect 355 333 371 349
rect 473 349 539 383
rect 473 333 489 349
rect 355 315 489 333
rect 523 337 539 349
rect 523 315 627 337
rect 137 299 627 315
rect 21 249 523 265
rect 21 215 37 249
rect 71 215 305 249
rect 339 215 389 249
rect 423 215 473 249
rect 507 215 523 249
rect 557 181 627 299
rect 153 145 627 181
rect 26 93 79 109
rect 26 59 45 93
rect 26 17 79 59
rect 153 101 187 145
rect 153 51 187 67
rect 237 93 271 109
rect 237 17 271 59
rect 321 101 355 145
rect 321 51 355 67
rect 405 93 439 109
rect 405 17 439 59
rect 489 101 523 145
rect 489 51 523 67
rect 557 94 607 110
rect 557 60 573 94
rect 557 17 607 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 573 153 607 187 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 573 221 607 255 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 573 289 607 323 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 297 221 331 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 389 221 423 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 481 221 515 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 inv_6
rlabel metal1 s 0 -48 644 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 2229860
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2223910
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
