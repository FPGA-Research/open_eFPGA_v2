magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 222 582
<< pwell >>
rect 3 38 181 195
<< locali >>
rect 17 294 167 491
rect 17 53 167 162
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 29 -17 63 17
rect 121 -17 155 17
<< metal1 >>
rect 0 561 184 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 184 561
rect 0 496 184 527
rect 0 17 184 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 184 17
rect 0 -48 184 -17
<< labels >>
rlabel metal1 s 0 -48 184 48 8 VGND
port 1 nsew ground bidirectional abutment
rlabel locali s 17 53 167 162 6 VNB
port 2 nsew ground bidirectional
rlabel pwell s 3 38 181 195 6 VNB
port 2 nsew ground bidirectional
rlabel locali s 17 294 167 491 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -38 261 222 582 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 496 184 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 184 544
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 561584
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 559332
<< end >>
