magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -26 -26 286 3026
<< psubdiff >>
rect 0 2970 60 3000
rect 0 2936 11 2970
rect 45 2936 60 2970
rect 0 2902 60 2936
rect 0 2868 11 2902
rect 45 2868 60 2902
rect 0 2834 60 2868
rect 0 2800 11 2834
rect 45 2800 60 2834
rect 0 2766 60 2800
rect 0 2732 11 2766
rect 45 2732 60 2766
rect 0 2698 60 2732
rect 0 2664 11 2698
rect 45 2664 60 2698
rect 0 2630 60 2664
rect 0 2596 11 2630
rect 45 2596 60 2630
rect 0 2562 60 2596
rect 0 2528 11 2562
rect 45 2528 60 2562
rect 0 2494 60 2528
rect 0 2460 11 2494
rect 45 2460 60 2494
rect 0 2426 60 2460
rect 0 2392 11 2426
rect 45 2392 60 2426
rect 0 2358 60 2392
rect 0 2324 11 2358
rect 45 2324 60 2358
rect 0 2290 60 2324
rect 0 2256 11 2290
rect 45 2256 60 2290
rect 0 2222 60 2256
rect 0 2188 11 2222
rect 45 2188 60 2222
rect 0 2154 60 2188
rect 0 2120 11 2154
rect 45 2120 60 2154
rect 0 2086 60 2120
rect 0 2052 11 2086
rect 45 2052 60 2086
rect 0 2018 60 2052
rect 0 1984 11 2018
rect 45 1984 60 2018
rect 0 1950 60 1984
rect 0 1916 11 1950
rect 45 1916 60 1950
rect 0 1882 60 1916
rect 0 1848 11 1882
rect 45 1848 60 1882
rect 0 1814 60 1848
rect 0 1780 11 1814
rect 45 1780 60 1814
rect 0 1746 60 1780
rect 0 1712 11 1746
rect 45 1712 60 1746
rect 0 1678 60 1712
rect 0 1644 11 1678
rect 45 1644 60 1678
rect 0 1610 60 1644
rect 0 1576 11 1610
rect 45 1576 60 1610
rect 0 1542 60 1576
rect 0 1508 11 1542
rect 45 1508 60 1542
rect 0 1474 60 1508
rect 0 1440 11 1474
rect 45 1440 60 1474
rect 0 1406 60 1440
rect 0 1372 11 1406
rect 45 1372 60 1406
rect 0 1338 60 1372
rect 0 1304 11 1338
rect 45 1304 60 1338
rect 0 1270 60 1304
rect 0 1236 11 1270
rect 45 1236 60 1270
rect 0 1202 60 1236
rect 0 1168 11 1202
rect 45 1168 60 1202
rect 0 1134 60 1168
rect 0 1100 11 1134
rect 45 1100 60 1134
rect 0 1066 60 1100
rect 0 1032 11 1066
rect 45 1032 60 1066
rect 0 998 60 1032
rect 0 964 11 998
rect 45 964 60 998
rect 0 930 60 964
rect 0 896 11 930
rect 45 896 60 930
rect 0 862 60 896
rect 0 828 11 862
rect 45 828 60 862
rect 0 794 60 828
rect 0 760 11 794
rect 45 760 60 794
rect 0 726 60 760
rect 0 692 11 726
rect 45 692 60 726
rect 0 658 60 692
rect 0 624 11 658
rect 45 624 60 658
rect 0 590 60 624
rect 0 556 11 590
rect 45 556 60 590
rect 0 522 60 556
rect 0 488 11 522
rect 45 488 60 522
rect 0 454 60 488
rect 0 420 11 454
rect 45 420 60 454
rect 0 386 60 420
rect 0 352 11 386
rect 45 352 60 386
rect 0 318 60 352
rect 0 284 11 318
rect 45 284 60 318
rect 0 250 60 284
rect 0 216 11 250
rect 45 216 60 250
rect 0 182 60 216
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
rect 200 2970 260 3000
rect 200 2936 215 2970
rect 249 2936 260 2970
rect 200 2902 260 2936
rect 200 2868 215 2902
rect 249 2868 260 2902
rect 200 2834 260 2868
rect 200 2800 215 2834
rect 249 2800 260 2834
rect 200 2766 260 2800
rect 200 2732 215 2766
rect 249 2732 260 2766
rect 200 2698 260 2732
rect 200 2664 215 2698
rect 249 2664 260 2698
rect 200 2630 260 2664
rect 200 2596 215 2630
rect 249 2596 260 2630
rect 200 2562 260 2596
rect 200 2528 215 2562
rect 249 2528 260 2562
rect 200 2494 260 2528
rect 200 2460 215 2494
rect 249 2460 260 2494
rect 200 2426 260 2460
rect 200 2392 215 2426
rect 249 2392 260 2426
rect 200 2358 260 2392
rect 200 2324 215 2358
rect 249 2324 260 2358
rect 200 2290 260 2324
rect 200 2256 215 2290
rect 249 2256 260 2290
rect 200 2222 260 2256
rect 200 2188 215 2222
rect 249 2188 260 2222
rect 200 2154 260 2188
rect 200 2120 215 2154
rect 249 2120 260 2154
rect 200 2086 260 2120
rect 200 2052 215 2086
rect 249 2052 260 2086
rect 200 2018 260 2052
rect 200 1984 215 2018
rect 249 1984 260 2018
rect 200 1950 260 1984
rect 200 1916 215 1950
rect 249 1916 260 1950
rect 200 1882 260 1916
rect 200 1848 215 1882
rect 249 1848 260 1882
rect 200 1814 260 1848
rect 200 1780 215 1814
rect 249 1780 260 1814
rect 200 1746 260 1780
rect 200 1712 215 1746
rect 249 1712 260 1746
rect 200 1678 260 1712
rect 200 1644 215 1678
rect 249 1644 260 1678
rect 200 1610 260 1644
rect 200 1576 215 1610
rect 249 1576 260 1610
rect 200 1542 260 1576
rect 200 1508 215 1542
rect 249 1508 260 1542
rect 200 1474 260 1508
rect 200 1440 215 1474
rect 249 1440 260 1474
rect 200 1406 260 1440
rect 200 1372 215 1406
rect 249 1372 260 1406
rect 200 1338 260 1372
rect 200 1304 215 1338
rect 249 1304 260 1338
rect 200 1270 260 1304
rect 200 1236 215 1270
rect 249 1236 260 1270
rect 200 1202 260 1236
rect 200 1168 215 1202
rect 249 1168 260 1202
rect 200 1134 260 1168
rect 200 1100 215 1134
rect 249 1100 260 1134
rect 200 1066 260 1100
rect 200 1032 215 1066
rect 249 1032 260 1066
rect 200 998 260 1032
rect 200 964 215 998
rect 249 964 260 998
rect 200 930 260 964
rect 200 896 215 930
rect 249 896 260 930
rect 200 862 260 896
rect 200 828 215 862
rect 249 828 260 862
rect 200 794 260 828
rect 200 760 215 794
rect 249 760 260 794
rect 200 726 260 760
rect 200 692 215 726
rect 249 692 260 726
rect 200 658 260 692
rect 200 624 215 658
rect 249 624 260 658
rect 200 590 260 624
rect 200 556 215 590
rect 249 556 260 590
rect 200 522 260 556
rect 200 488 215 522
rect 249 488 260 522
rect 200 454 260 488
rect 200 420 215 454
rect 249 420 260 454
rect 200 386 260 420
rect 200 352 215 386
rect 249 352 260 386
rect 200 318 260 352
rect 200 284 215 318
rect 249 284 260 318
rect 200 250 260 284
rect 200 216 215 250
rect 249 216 260 250
rect 200 182 260 216
rect 200 148 215 182
rect 249 148 260 182
rect 200 114 260 148
rect 200 80 215 114
rect 249 80 260 114
rect 200 46 260 80
rect 200 12 215 46
rect 249 12 260 46
rect 200 0 260 12
<< nsubdiff >>
rect 60 0 200 3000
<< psubdiffcont >>
rect 11 2936 45 2970
rect 11 2868 45 2902
rect 11 2800 45 2834
rect 11 2732 45 2766
rect 11 2664 45 2698
rect 11 2596 45 2630
rect 11 2528 45 2562
rect 11 2460 45 2494
rect 11 2392 45 2426
rect 11 2324 45 2358
rect 11 2256 45 2290
rect 11 2188 45 2222
rect 11 2120 45 2154
rect 11 2052 45 2086
rect 11 1984 45 2018
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
rect 215 2936 249 2970
rect 215 2868 249 2902
rect 215 2800 249 2834
rect 215 2732 249 2766
rect 215 2664 249 2698
rect 215 2596 249 2630
rect 215 2528 249 2562
rect 215 2460 249 2494
rect 215 2392 249 2426
rect 215 2324 249 2358
rect 215 2256 249 2290
rect 215 2188 249 2222
rect 215 2120 249 2154
rect 215 2052 249 2086
rect 215 1984 249 2018
rect 215 1916 249 1950
rect 215 1848 249 1882
rect 215 1780 249 1814
rect 215 1712 249 1746
rect 215 1644 249 1678
rect 215 1576 249 1610
rect 215 1508 249 1542
rect 215 1440 249 1474
rect 215 1372 249 1406
rect 215 1304 249 1338
rect 215 1236 249 1270
rect 215 1168 249 1202
rect 215 1100 249 1134
rect 215 1032 249 1066
rect 215 964 249 998
rect 215 896 249 930
rect 215 828 249 862
rect 215 760 249 794
rect 215 692 249 726
rect 215 624 249 658
rect 215 556 249 590
rect 215 488 249 522
rect 215 420 249 454
rect 215 352 249 386
rect 215 284 249 318
rect 215 216 249 250
rect 215 148 249 182
rect 215 80 249 114
rect 215 12 249 46
<< locali >>
rect 11 2970 249 2986
rect 45 2936 215 2970
rect 11 2902 249 2936
rect 45 2868 215 2902
rect 11 2834 249 2868
rect 45 2800 215 2834
rect 11 2766 249 2800
rect 45 2732 215 2766
rect 11 2698 249 2732
rect 45 2664 215 2698
rect 11 2630 249 2664
rect 45 2596 215 2630
rect 11 2562 249 2596
rect 45 2528 215 2562
rect 11 2494 249 2528
rect 45 2460 215 2494
rect 11 2426 249 2460
rect 45 2392 215 2426
rect 11 2358 249 2392
rect 45 2324 215 2358
rect 11 2290 249 2324
rect 45 2256 215 2290
rect 11 2222 249 2256
rect 45 2188 215 2222
rect 11 2154 249 2188
rect 45 2120 215 2154
rect 11 2086 249 2120
rect 45 2052 215 2086
rect 11 2018 249 2052
rect 45 1984 215 2018
rect 11 1950 249 1984
rect 45 1916 215 1950
rect 11 1882 249 1916
rect 45 1848 215 1882
rect 11 1814 249 1848
rect 45 1780 215 1814
rect 11 1746 249 1780
rect 45 1712 215 1746
rect 11 1678 249 1712
rect 45 1644 215 1678
rect 11 1610 249 1644
rect 45 1576 215 1610
rect 11 1542 249 1576
rect 45 1508 215 1542
rect 11 1474 249 1508
rect 45 1440 215 1474
rect 11 1406 249 1440
rect 45 1372 215 1406
rect 11 1338 249 1372
rect 45 1304 215 1338
rect 11 1270 249 1304
rect 45 1236 215 1270
rect 11 1202 249 1236
rect 45 1168 215 1202
rect 11 1134 249 1168
rect 45 1100 215 1134
rect 11 1066 249 1100
rect 45 1032 215 1066
rect 11 998 249 1032
rect 45 964 215 998
rect 11 930 249 964
rect 45 896 215 930
rect 11 862 249 896
rect 45 828 215 862
rect 11 794 249 828
rect 45 760 215 794
rect 11 726 249 760
rect 45 692 215 726
rect 11 658 249 692
rect 45 624 215 658
rect 11 590 249 624
rect 45 556 215 590
rect 11 522 249 556
rect 45 488 215 522
rect 11 454 249 488
rect 45 420 215 454
rect 11 386 249 420
rect 45 352 215 386
rect 11 318 249 352
rect 45 284 215 318
rect 11 250 249 284
rect 45 216 215 250
rect 11 182 249 216
rect 45 148 215 182
rect 11 114 249 148
rect 45 80 215 114
rect 11 46 249 80
rect 45 12 215 46
rect 11 -4 249 12
<< properties >>
string GDS_END 89385734
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89376706
<< end >>
