magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 2152 1591 2424
rect 0 272 272 2152
rect 1319 272 1591 2152
rect 0 0 1591 272
<< pwell >>
rect 332 332 1259 2092
<< mvnmosesd >>
tri 695 1712 735 1752 ne
tri 695 672 735 712 se
rect 735 672 855 1752
tri 855 1712 895 1752 nw
tri 855 672 895 712 sw
<< mvndiff >>
rect 594 1712 695 1752
tri 695 1712 735 1752 sw
rect 594 712 735 1712
rect 594 672 695 712
tri 695 672 735 712 nw
tri 855 1712 895 1752 se
rect 895 1712 996 1752
rect 855 712 996 1712
tri 855 672 895 712 ne
rect 895 672 996 712
<< mvpsubdiff >>
rect 358 1926 1233 2066
rect 358 498 462 1926
rect 1129 498 1233 1926
rect 358 358 1233 498
<< mvnsubdiff >>
rect 66 2218 1525 2358
rect 66 206 206 2218
rect 1385 206 1525 2218
rect 66 66 1525 206
<< poly >>
rect 655 1846 935 1866
rect 655 1812 676 1846
rect 710 1812 744 1846
rect 778 1812 812 1846
rect 846 1812 880 1846
rect 914 1812 935 1846
rect 655 1792 935 1812
tri 655 1752 695 1792 ne
rect 695 1752 895 1792
tri 895 1752 935 1792 nw
tri 655 632 695 672 se
rect 695 632 895 672
tri 895 632 935 672 sw
rect 655 558 935 632
<< polycont >>
rect 676 1812 710 1846
rect 744 1812 778 1846
rect 812 1812 846 1846
rect 880 1812 914 1846
<< locali >>
rect 66 2305 1525 2358
rect 66 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1525 2305
rect 66 2218 1525 2271
rect 66 206 206 2218
rect 358 2003 1233 2066
rect 358 1969 454 2003
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 1969 1233 2003
rect 358 1924 1233 1969
rect 358 498 498 1924
rect 662 1847 927 1867
rect 662 1846 725 1847
rect 759 1846 797 1847
rect 831 1846 927 1847
rect 662 1812 676 1846
rect 710 1813 725 1846
rect 778 1813 797 1846
rect 710 1812 744 1813
rect 778 1812 812 1813
rect 846 1812 880 1846
rect 914 1812 927 1846
rect 662 1785 927 1812
rect 593 672 701 1751
rect 888 672 996 1751
rect 1093 498 1233 1924
rect 358 358 1233 498
rect 1385 206 1525 2218
rect 66 142 1525 206
rect 66 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1525 142
rect 66 66 1525 108
<< viali >>
rect 307 2271 341 2305
rect 379 2271 413 2305
rect 451 2271 485 2305
rect 523 2271 557 2305
rect 595 2271 629 2305
rect 959 2271 993 2305
rect 1031 2271 1065 2305
rect 1103 2271 1137 2305
rect 1175 2271 1209 2305
rect 1247 2271 1281 2305
rect 454 1969 488 2003
rect 526 1969 560 2003
rect 598 1969 632 2003
rect 928 1969 962 2003
rect 1000 1969 1034 2003
rect 1072 1969 1106 2003
rect 725 1846 759 1847
rect 797 1846 831 1847
rect 725 1813 744 1846
rect 744 1813 759 1846
rect 797 1813 812 1846
rect 812 1813 831 1846
rect 1118 108 1152 142
rect 1190 108 1224 142
rect 1262 108 1296 142
<< metal1 >>
tri 161 2311 208 2358 se
rect 208 2311 669 2358
tri 155 2305 161 2311 se
rect 161 2305 669 2311
tri 121 2271 155 2305 se
rect 155 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 669 2305
tri 115 2265 121 2271 se
rect 121 2265 669 2271
tri 66 2216 115 2265 se
rect 115 2218 669 2265
rect 115 2216 286 2218
tri 286 2216 288 2218 nw
rect 66 69 206 2216
tri 206 2136 286 2216 nw
tri 367 2009 424 2066 se
rect 424 2009 669 2066
tri 361 2003 367 2009 se
rect 367 2003 669 2009
rect 66 66 203 69
rect 204 67 205 68
tri 358 2000 361 2003 se
rect 361 2000 454 2003
rect 358 1969 454 2000
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 669 2003
rect 358 1901 669 1969
rect 358 1853 563 1901
tri 563 1853 611 1901 nw
rect 358 1847 557 1853
tri 557 1847 563 1853 nw
rect 703 1847 852 2359
rect 886 2311 1383 2358
tri 1383 2311 1430 2358 sw
rect 886 2305 1430 2311
rect 886 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1430 2305
rect 886 2265 1430 2271
tri 1430 2265 1476 2311 sw
rect 886 2218 1476 2265
tri 1289 2216 1291 2218 ne
rect 1291 2216 1476 2218
tri 1476 2216 1525 2265 sw
tri 1291 2124 1383 2216 ne
rect 1383 2124 1525 2216
tri 1383 2122 1385 2124 ne
rect 886 2009 1167 2066
tri 1167 2009 1224 2066 sw
rect 886 2003 1224 2009
rect 886 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 2000 1224 2003
tri 1224 2000 1233 2009 sw
rect 1106 1969 1233 2000
rect 886 1901 1233 1969
rect 358 69 536 1847
tri 536 1826 557 1847 nw
rect 703 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 852 1847
tri 1012 1820 1093 1901 ne
rect 703 1791 852 1813
rect 358 66 533 69
rect 534 67 535 68
rect 572 66 772 1709
rect 831 66 1031 1752
rect 1093 358 1233 1901
tri 1289 206 1385 302 se
rect 1385 208 1525 2124
rect 1385 206 1523 208
tri 1523 206 1525 208 nw
rect 1070 148 1465 206
tri 1465 148 1523 206 nw
rect 1070 142 1419 148
rect 1070 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1419 142
rect 1070 102 1419 108
tri 1419 102 1465 148 nw
rect 1070 66 1383 102
tri 1383 66 1419 102 nw
<< rmetal1 >>
rect 203 68 206 69
rect 203 67 204 68
rect 205 67 206 68
rect 203 66 206 67
rect 533 68 536 69
rect 533 67 534 68
rect 535 67 536 68
rect 533 66 536 67
use DFL1_CDNS_52468879185222  DFL1_CDNS_52468879185222_0
timestamp 1707688321
transform 1 0 594 0 1 705
box -26 -26 76 968
use DFL1_CDNS_52468879185222  DFL1_CDNS_52468879185222_1
timestamp 1707688321
transform 1 0 938 0 1 705
box -26 -26 76 968
use L1M1_CDNS_52468879185216  L1M1_CDNS_52468879185216_0
timestamp 1707688321
transform 1 0 928 0 1 1969
box 0 0 1 1
use L1M1_CDNS_52468879185216  L1M1_CDNS_52468879185216_1
timestamp 1707688321
transform 1 0 454 0 1 1969
box 0 0 1 1
use L1M1_CDNS_52468879185216  L1M1_CDNS_52468879185216_2
timestamp 1707688321
transform 1 0 1118 0 1 108
box 0 0 1 1
use L1M1_CDNS_52468879185217  L1M1_CDNS_52468879185217_0
timestamp 1707688321
transform 1 0 1438 0 1 273
box -12 -6 46 1768
use L1M1_CDNS_52468879185217  L1M1_CDNS_52468879185217_1
timestamp 1707688321
transform 1 0 119 0 1 273
box -12 -6 46 1768
use L1M1_CDNS_52468879185218  L1M1_CDNS_52468879185218_0
timestamp 1707688321
transform 1 0 395 0 1 401
box -12 -6 46 1408
use L1M1_CDNS_52468879185218  L1M1_CDNS_52468879185218_1
timestamp 1707688321
transform 1 0 1146 0 1 401
box -12 -6 46 1408
use L1M1_CDNS_52468879185219  L1M1_CDNS_52468879185219_0
timestamp 1707688321
transform 1 0 621 0 1 757
box -12 -6 46 832
use L1M1_CDNS_52468879185219  L1M1_CDNS_52468879185219_1
timestamp 1707688321
transform 1 0 915 0 1 757
box -12 -6 46 832
use L1M1_CDNS_52468879185220  L1M1_CDNS_52468879185220_0
timestamp 1707688321
transform 1 0 307 0 1 2271
box 0 0 1 1
use L1M1_CDNS_52468879185220  L1M1_CDNS_52468879185220_1
timestamp 1707688321
transform 1 0 959 0 1 2271
box 0 0 1 1
use L1M1_CDNS_52468879185221  L1M1_CDNS_52468879185221_0
timestamp 1707688321
transform 1 0 725 0 1 1813
box 0 0 1 1
use PYL1_CDNS_52468879185211  PYL1_CDNS_52468879185211_0
timestamp 1707688321
transform 1 0 660 0 1 1796
box 0 0 1 1
use TPL1_CDNS_52468879185212  TPL1_CDNS_52468879185212_0
timestamp 1707688321
transform 1 0 279 0 1 2247
box -36 -36 1070 118
use TPL1_CDNS_52468879185212  TPL1_CDNS_52468879185212_1
timestamp 1707688321
transform 1 0 279 0 1 95
box -36 -36 1070 118
use TPL1_CDNS_52468879185213  TPL1_CDNS_52468879185213_0
timestamp 1707688321
transform 1 0 449 0 1 387
box -26 -26 720 108
use TPL1_CDNS_52468879185213  TPL1_CDNS_52468879185213_1
timestamp 1707688321
transform 1 0 449 0 1 1955
box -26 -26 720 108
use TPL1_CDNS_52468879185214  TPL1_CDNS_52468879185214_0
timestamp 1707688321
transform 1 0 1132 0 1 509
box -26 -26 108 1332
use TPL1_CDNS_52468879185214  TPL1_CDNS_52468879185214_1
timestamp 1707688321
transform 1 0 380 0 1 509
box -26 -26 108 1332
use TPL1_CDNS_52468879185215  TPL1_CDNS_52468879185215_0
timestamp 1707688321
transform 1 0 1414 0 1 198
box -36 -36 118 1954
use TPL1_CDNS_52468879185215  TPL1_CDNS_52468879185215_1
timestamp 1707688321
transform 1 0 95 0 1 198
box -36 -36 118 1954
<< labels >>
flabel comment s 783 2298 783 2298 0 FreeSans 500 0 0 0 Do not merge with PFET NWELL
flabel comment s 129 1085 129 1085 0 FreeSans 500 90 0 0 Do not merge with PFET NWELL
flabel comment s 1452 1103 1452 1103 0 FreeSans 500 270 0 0 Do not merge with PFET NWELL
flabel metal1 s 888 70 996 103 0 FreeSans 400 0 0 0 in
port 1 nsew
flabel metal1 s 387 82 514 122 0 FreeSans 300 0 0 0 nbody
port 2 nsew
flabel metal1 s 628 78 721 118 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 68 77 204 117 0 FreeSans 200 0 0 0 nwellRing
port 4 nsew
flabel metal1 s 703 2259 852 2359 0 FreeSans 300 0 0 0 gate
port 5 nsew
<< properties >>
string GDS_END 85841866
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85837568
<< end >>
