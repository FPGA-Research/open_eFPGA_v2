magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 154
rect 61 0 64 154
<< via1 >>
rect 3 0 61 154
<< metal2 >>
rect 0 0 3 154
rect 61 0 64 154
<< properties >>
string GDS_END 85244614
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85243842
<< end >>
