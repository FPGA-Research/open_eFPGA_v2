magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -53 50677 162 50743
rect -53 34928 261 50677
rect -2967 34747 261 34928
rect -2867 34614 261 34747
rect 2 9740 584 9871
rect 1754 9740 2560 9864
rect 3730 9763 4788 9871
rect 5958 9740 6452 9864
<< pwell >>
rect -2995 34994 -127 50674
rect -2992 7396 -240 17977
rect 18255 14234 29695 14510
rect 15805 14058 29695 14234
rect 15805 13782 18707 14058
rect 4395 10040 6265 11960
rect 13198 10203 15910 12147
rect 12454 9969 15910 10203
rect 12454 9932 15220 9969
rect 32002 8322 32087 8568
<< pdiff >>
rect 28582 15752 30572 15812
rect 1513 5830 2218 5881
rect 3194 5830 3770 5881
rect 1513 5778 3770 5830
<< psubdiff >>
rect 4421 11910 6239 11934
rect 4421 11332 4429 11910
rect 6231 11332 6239 11910
rect 4421 11297 6239 11332
rect 4421 11263 4429 11297
rect 4463 11263 4497 11297
rect 4531 11263 4565 11297
rect 4599 11263 4633 11297
rect 4667 11263 4701 11297
rect 4735 11263 4769 11297
rect 4803 11263 4837 11297
rect 4871 11263 4905 11297
rect 4939 11263 4973 11297
rect 5007 11263 5041 11297
rect 5075 11263 5109 11297
rect 5143 11263 5177 11297
rect 5211 11263 5245 11297
rect 5279 11263 5313 11297
rect 5347 11263 5381 11297
rect 5415 11263 5449 11297
rect 5483 11263 5517 11297
rect 5551 11263 5585 11297
rect 5619 11263 5653 11297
rect 5687 11263 5721 11297
rect 5755 11263 5789 11297
rect 5823 11263 5857 11297
rect 5891 11263 5925 11297
rect 5959 11263 5993 11297
rect 6027 11263 6061 11297
rect 6095 11263 6129 11297
rect 6163 11263 6197 11297
rect 6231 11263 6239 11297
rect 4421 11228 6239 11263
rect 4421 11194 4429 11228
rect 4463 11194 4497 11228
rect 4531 11194 4565 11228
rect 4599 11194 4633 11228
rect 4667 11194 4701 11228
rect 4735 11194 4769 11228
rect 4803 11194 4837 11228
rect 4871 11194 4905 11228
rect 4939 11194 4973 11228
rect 5007 11194 5041 11228
rect 5075 11194 5109 11228
rect 5143 11194 5177 11228
rect 5211 11194 5245 11228
rect 5279 11194 5313 11228
rect 5347 11194 5381 11228
rect 5415 11194 5449 11228
rect 5483 11194 5517 11228
rect 5551 11194 5585 11228
rect 5619 11194 5653 11228
rect 5687 11194 5721 11228
rect 5755 11194 5789 11228
rect 5823 11194 5857 11228
rect 5891 11194 5925 11228
rect 5959 11194 5993 11228
rect 6027 11194 6061 11228
rect 6095 11194 6129 11228
rect 6163 11194 6197 11228
rect 6231 11194 6239 11228
rect 4421 11159 6239 11194
rect 4421 11125 4429 11159
rect 4463 11125 4497 11159
rect 4531 11125 4565 11159
rect 4599 11125 4633 11159
rect 4667 11125 4701 11159
rect 4735 11125 4769 11159
rect 4803 11125 4837 11159
rect 4871 11125 4905 11159
rect 4939 11125 4973 11159
rect 5007 11125 5041 11159
rect 5075 11125 5109 11159
rect 5143 11125 5177 11159
rect 5211 11125 5245 11159
rect 5279 11125 5313 11159
rect 5347 11125 5381 11159
rect 5415 11125 5449 11159
rect 5483 11125 5517 11159
rect 5551 11125 5585 11159
rect 5619 11125 5653 11159
rect 5687 11125 5721 11159
rect 5755 11125 5789 11159
rect 5823 11125 5857 11159
rect 5891 11125 5925 11159
rect 5959 11125 5993 11159
rect 6027 11125 6061 11159
rect 6095 11125 6129 11159
rect 6163 11125 6197 11159
rect 6231 11125 6239 11159
rect 4421 11090 6239 11125
rect 4421 11056 4429 11090
rect 4463 11056 4497 11090
rect 4531 11056 4565 11090
rect 4599 11056 4633 11090
rect 4667 11056 4701 11090
rect 4735 11056 4769 11090
rect 4803 11056 4837 11090
rect 4871 11056 4905 11090
rect 4939 11056 4973 11090
rect 5007 11056 5041 11090
rect 5075 11056 5109 11090
rect 5143 11056 5177 11090
rect 5211 11056 5245 11090
rect 5279 11056 5313 11090
rect 5347 11056 5381 11090
rect 5415 11056 5449 11090
rect 5483 11056 5517 11090
rect 5551 11056 5585 11090
rect 5619 11056 5653 11090
rect 5687 11056 5721 11090
rect 5755 11056 5789 11090
rect 5823 11056 5857 11090
rect 5891 11056 5925 11090
rect 5959 11056 5993 11090
rect 6027 11056 6061 11090
rect 6095 11056 6129 11090
rect 6163 11056 6197 11090
rect 6231 11056 6239 11090
rect 4421 11021 6239 11056
rect 4421 10987 4429 11021
rect 4463 10987 4497 11021
rect 4531 10987 4565 11021
rect 4599 10987 4633 11021
rect 4667 10987 4701 11021
rect 4735 10987 4769 11021
rect 4803 10987 4837 11021
rect 4871 10987 4905 11021
rect 4939 10987 4973 11021
rect 5007 10987 5041 11021
rect 5075 10987 5109 11021
rect 5143 10987 5177 11021
rect 5211 10987 5245 11021
rect 5279 10987 5313 11021
rect 5347 10987 5381 11021
rect 5415 10987 5449 11021
rect 5483 10987 5517 11021
rect 5551 10987 5585 11021
rect 5619 10987 5653 11021
rect 5687 10987 5721 11021
rect 5755 10987 5789 11021
rect 5823 10987 5857 11021
rect 5891 10987 5925 11021
rect 5959 10987 5993 11021
rect 6027 10987 6061 11021
rect 6095 10987 6129 11021
rect 6163 10987 6197 11021
rect 6231 10987 6239 11021
rect 4421 10952 6239 10987
rect 4421 10918 4429 10952
rect 4463 10918 4497 10952
rect 4531 10918 4565 10952
rect 4599 10918 4633 10952
rect 4667 10918 4701 10952
rect 4735 10918 4769 10952
rect 4803 10918 4837 10952
rect 4871 10918 4905 10952
rect 4939 10918 4973 10952
rect 5007 10918 5041 10952
rect 5075 10918 5109 10952
rect 5143 10918 5177 10952
rect 5211 10918 5245 10952
rect 5279 10918 5313 10952
rect 5347 10918 5381 10952
rect 5415 10918 5449 10952
rect 5483 10918 5517 10952
rect 5551 10918 5585 10952
rect 5619 10918 5653 10952
rect 5687 10918 5721 10952
rect 5755 10918 5789 10952
rect 5823 10918 5857 10952
rect 5891 10918 5925 10952
rect 5959 10918 5993 10952
rect 6027 10918 6061 10952
rect 6095 10918 6129 10952
rect 6163 10918 6197 10952
rect 6231 10918 6239 10952
rect 4421 10883 6239 10918
rect 4421 10849 4429 10883
rect 4463 10849 4497 10883
rect 4531 10849 4565 10883
rect 4599 10849 4633 10883
rect 4667 10849 4701 10883
rect 4735 10849 4769 10883
rect 4803 10849 4837 10883
rect 4871 10849 4905 10883
rect 4939 10849 4973 10883
rect 5007 10849 5041 10883
rect 5075 10849 5109 10883
rect 5143 10849 5177 10883
rect 5211 10849 5245 10883
rect 5279 10849 5313 10883
rect 5347 10849 5381 10883
rect 5415 10849 5449 10883
rect 5483 10849 5517 10883
rect 5551 10849 5585 10883
rect 5619 10849 5653 10883
rect 5687 10849 5721 10883
rect 5755 10849 5789 10883
rect 5823 10849 5857 10883
rect 5891 10849 5925 10883
rect 5959 10849 5993 10883
rect 6027 10849 6061 10883
rect 6095 10849 6129 10883
rect 6163 10849 6197 10883
rect 6231 10849 6239 10883
rect 4421 10814 6239 10849
rect 4421 10780 4429 10814
rect 4463 10780 4497 10814
rect 4531 10780 4565 10814
rect 4599 10780 4633 10814
rect 4667 10780 4701 10814
rect 4735 10780 4769 10814
rect 4803 10780 4837 10814
rect 4871 10780 4905 10814
rect 4939 10780 4973 10814
rect 5007 10780 5041 10814
rect 5075 10780 5109 10814
rect 5143 10780 5177 10814
rect 5211 10780 5245 10814
rect 5279 10780 5313 10814
rect 5347 10780 5381 10814
rect 5415 10780 5449 10814
rect 5483 10780 5517 10814
rect 5551 10780 5585 10814
rect 5619 10780 5653 10814
rect 5687 10780 5721 10814
rect 5755 10780 5789 10814
rect 5823 10780 5857 10814
rect 5891 10780 5925 10814
rect 5959 10780 5993 10814
rect 6027 10780 6061 10814
rect 6095 10780 6129 10814
rect 6163 10780 6197 10814
rect 6231 10780 6239 10814
rect 4421 10745 6239 10780
rect 4421 10711 4429 10745
rect 4463 10711 4497 10745
rect 4531 10711 4565 10745
rect 4599 10711 4633 10745
rect 4667 10711 4701 10745
rect 4735 10711 4769 10745
rect 4803 10711 4837 10745
rect 4871 10711 4905 10745
rect 4939 10711 4973 10745
rect 5007 10711 5041 10745
rect 5075 10711 5109 10745
rect 5143 10711 5177 10745
rect 5211 10711 5245 10745
rect 5279 10711 5313 10745
rect 5347 10711 5381 10745
rect 5415 10711 5449 10745
rect 5483 10711 5517 10745
rect 5551 10711 5585 10745
rect 5619 10711 5653 10745
rect 5687 10711 5721 10745
rect 5755 10711 5789 10745
rect 5823 10711 5857 10745
rect 5891 10711 5925 10745
rect 5959 10711 5993 10745
rect 6027 10711 6061 10745
rect 6095 10711 6129 10745
rect 6163 10711 6197 10745
rect 6231 10711 6239 10745
rect 4421 10676 6239 10711
rect 4421 10642 4429 10676
rect 4463 10642 4497 10676
rect 4531 10642 4565 10676
rect 4599 10642 4633 10676
rect 4667 10642 4701 10676
rect 4735 10642 4769 10676
rect 4803 10642 4837 10676
rect 4871 10642 4905 10676
rect 4939 10642 4973 10676
rect 5007 10642 5041 10676
rect 5075 10642 5109 10676
rect 5143 10642 5177 10676
rect 5211 10642 5245 10676
rect 5279 10642 5313 10676
rect 5347 10642 5381 10676
rect 5415 10642 5449 10676
rect 5483 10642 5517 10676
rect 5551 10642 5585 10676
rect 5619 10642 5653 10676
rect 5687 10642 5721 10676
rect 5755 10642 5789 10676
rect 5823 10642 5857 10676
rect 5891 10642 5925 10676
rect 5959 10642 5993 10676
rect 6027 10642 6061 10676
rect 6095 10642 6129 10676
rect 6163 10642 6197 10676
rect 6231 10642 6239 10676
rect 4421 10607 6239 10642
rect 4421 10573 4429 10607
rect 4463 10573 4497 10607
rect 4531 10573 4565 10607
rect 4599 10573 4633 10607
rect 4667 10573 4701 10607
rect 4735 10573 4769 10607
rect 4803 10573 4837 10607
rect 4871 10573 4905 10607
rect 4939 10573 4973 10607
rect 5007 10573 5041 10607
rect 5075 10573 5109 10607
rect 5143 10573 5177 10607
rect 5211 10573 5245 10607
rect 5279 10573 5313 10607
rect 5347 10573 5381 10607
rect 5415 10573 5449 10607
rect 5483 10573 5517 10607
rect 5551 10573 5585 10607
rect 5619 10573 5653 10607
rect 5687 10573 5721 10607
rect 5755 10573 5789 10607
rect 5823 10573 5857 10607
rect 5891 10573 5925 10607
rect 5959 10573 5993 10607
rect 6027 10573 6061 10607
rect 6095 10573 6129 10607
rect 6163 10573 6197 10607
rect 6231 10573 6239 10607
rect 4421 10538 6239 10573
rect 4421 10504 4429 10538
rect 4463 10504 4497 10538
rect 4531 10504 4565 10538
rect 4599 10504 4633 10538
rect 4667 10504 4701 10538
rect 4735 10504 4769 10538
rect 4803 10504 4837 10538
rect 4871 10504 4905 10538
rect 4939 10504 4973 10538
rect 5007 10504 5041 10538
rect 5075 10504 5109 10538
rect 5143 10504 5177 10538
rect 5211 10504 5245 10538
rect 5279 10504 5313 10538
rect 5347 10504 5381 10538
rect 5415 10504 5449 10538
rect 5483 10504 5517 10538
rect 5551 10504 5585 10538
rect 5619 10504 5653 10538
rect 5687 10504 5721 10538
rect 5755 10504 5789 10538
rect 5823 10504 5857 10538
rect 5891 10504 5925 10538
rect 5959 10504 5993 10538
rect 6027 10504 6061 10538
rect 6095 10504 6129 10538
rect 6163 10504 6197 10538
rect 6231 10504 6239 10538
rect 4421 10469 6239 10504
rect 4421 10435 4429 10469
rect 4463 10435 4497 10469
rect 4531 10435 4565 10469
rect 4599 10435 4633 10469
rect 4667 10435 4701 10469
rect 4735 10435 4769 10469
rect 4803 10435 4837 10469
rect 4871 10435 4905 10469
rect 4939 10435 4973 10469
rect 5007 10435 5041 10469
rect 5075 10435 5109 10469
rect 5143 10435 5177 10469
rect 5211 10435 5245 10469
rect 5279 10435 5313 10469
rect 5347 10435 5381 10469
rect 5415 10435 5449 10469
rect 5483 10435 5517 10469
rect 5551 10435 5585 10469
rect 5619 10435 5653 10469
rect 5687 10435 5721 10469
rect 5755 10435 5789 10469
rect 5823 10435 5857 10469
rect 5891 10435 5925 10469
rect 5959 10435 5993 10469
rect 6027 10435 6061 10469
rect 6095 10435 6129 10469
rect 6163 10435 6197 10469
rect 6231 10435 6239 10469
rect 4421 10400 6239 10435
rect 4421 10366 4429 10400
rect 4463 10366 4497 10400
rect 4531 10366 4565 10400
rect 4599 10366 4633 10400
rect 4667 10366 4701 10400
rect 4735 10366 4769 10400
rect 4803 10366 4837 10400
rect 4871 10366 4905 10400
rect 4939 10366 4973 10400
rect 5007 10366 5041 10400
rect 5075 10366 5109 10400
rect 5143 10366 5177 10400
rect 5211 10366 5245 10400
rect 5279 10366 5313 10400
rect 5347 10366 5381 10400
rect 5415 10366 5449 10400
rect 5483 10366 5517 10400
rect 5551 10366 5585 10400
rect 5619 10366 5653 10400
rect 5687 10366 5721 10400
rect 5755 10366 5789 10400
rect 5823 10366 5857 10400
rect 5891 10366 5925 10400
rect 5959 10366 5993 10400
rect 6027 10366 6061 10400
rect 6095 10366 6129 10400
rect 6163 10366 6197 10400
rect 6231 10366 6239 10400
rect 4421 10331 6239 10366
rect 4421 10297 4429 10331
rect 4463 10297 4497 10331
rect 4531 10297 4565 10331
rect 4599 10297 4633 10331
rect 4667 10297 4701 10331
rect 4735 10297 4769 10331
rect 4803 10297 4837 10331
rect 4871 10297 4905 10331
rect 4939 10297 4973 10331
rect 5007 10297 5041 10331
rect 5075 10297 5109 10331
rect 5143 10297 5177 10331
rect 5211 10297 5245 10331
rect 5279 10297 5313 10331
rect 5347 10297 5381 10331
rect 5415 10297 5449 10331
rect 5483 10297 5517 10331
rect 5551 10297 5585 10331
rect 5619 10297 5653 10331
rect 5687 10297 5721 10331
rect 5755 10297 5789 10331
rect 5823 10297 5857 10331
rect 5891 10297 5925 10331
rect 5959 10297 5993 10331
rect 6027 10297 6061 10331
rect 6095 10297 6129 10331
rect 6163 10297 6197 10331
rect 6231 10297 6239 10331
rect 4421 10262 6239 10297
rect 4421 10228 4429 10262
rect 4463 10228 4497 10262
rect 4531 10228 4565 10262
rect 4599 10228 4633 10262
rect 4667 10228 4701 10262
rect 4735 10228 4769 10262
rect 4803 10228 4837 10262
rect 4871 10228 4905 10262
rect 4939 10228 4973 10262
rect 5007 10228 5041 10262
rect 5075 10228 5109 10262
rect 5143 10228 5177 10262
rect 5211 10228 5245 10262
rect 5279 10228 5313 10262
rect 5347 10228 5381 10262
rect 5415 10228 5449 10262
rect 5483 10228 5517 10262
rect 5551 10228 5585 10262
rect 5619 10228 5653 10262
rect 5687 10228 5721 10262
rect 5755 10228 5789 10262
rect 5823 10228 5857 10262
rect 5891 10228 5925 10262
rect 5959 10228 5993 10262
rect 6027 10228 6061 10262
rect 6095 10228 6129 10262
rect 6163 10228 6197 10262
rect 6231 10228 6239 10262
rect 4421 10193 6239 10228
rect 4421 10159 4429 10193
rect 4463 10159 4497 10193
rect 4531 10159 4565 10193
rect 4599 10159 4633 10193
rect 4667 10159 4701 10193
rect 4735 10159 4769 10193
rect 4803 10159 4837 10193
rect 4871 10159 4905 10193
rect 4939 10159 4973 10193
rect 5007 10159 5041 10193
rect 5075 10159 5109 10193
rect 5143 10159 5177 10193
rect 5211 10159 5245 10193
rect 5279 10159 5313 10193
rect 5347 10159 5381 10193
rect 5415 10159 5449 10193
rect 5483 10159 5517 10193
rect 5551 10159 5585 10193
rect 5619 10159 5653 10193
rect 5687 10159 5721 10193
rect 5755 10159 5789 10193
rect 5823 10159 5857 10193
rect 5891 10159 5925 10193
rect 5959 10159 5993 10193
rect 6027 10159 6061 10193
rect 6095 10159 6129 10193
rect 6163 10159 6197 10193
rect 6231 10159 6239 10193
rect 4421 10124 6239 10159
rect 4421 10090 4429 10124
rect 4463 10090 4497 10124
rect 4531 10090 4565 10124
rect 4599 10090 4633 10124
rect 4667 10090 4701 10124
rect 4735 10090 4769 10124
rect 4803 10090 4837 10124
rect 4871 10090 4905 10124
rect 4939 10090 4973 10124
rect 5007 10090 5041 10124
rect 5075 10090 5109 10124
rect 5143 10090 5177 10124
rect 5211 10090 5245 10124
rect 5279 10090 5313 10124
rect 5347 10090 5381 10124
rect 5415 10090 5449 10124
rect 5483 10090 5517 10124
rect 5551 10090 5585 10124
rect 5619 10090 5653 10124
rect 5687 10090 5721 10124
rect 5755 10090 5789 10124
rect 5823 10090 5857 10124
rect 5891 10090 5925 10124
rect 5959 10090 5993 10124
rect 6027 10090 6061 10124
rect 6095 10090 6129 10124
rect 6163 10090 6197 10124
rect 6231 10090 6239 10124
rect 4421 10066 6239 10090
<< mvpsubdiff >>
rect -2969 50624 -153 50648
rect -2969 37942 -2938 50624
rect -184 37942 -153 50624
rect -2969 37907 -153 37942
rect -2969 37873 -2938 37907
rect -2904 37873 -2870 37907
rect -2836 37873 -2802 37907
rect -2768 37873 -2734 37907
rect -2700 37873 -2666 37907
rect -2632 37873 -2598 37907
rect -2564 37873 -2530 37907
rect -2496 37873 -2462 37907
rect -2428 37873 -2394 37907
rect -2360 37873 -2326 37907
rect -2292 37873 -2258 37907
rect -2224 37873 -2190 37907
rect -2156 37873 -2122 37907
rect -2088 37873 -2054 37907
rect -2020 37873 -1986 37907
rect -1952 37873 -1918 37907
rect -1884 37873 -1850 37907
rect -1816 37873 -1782 37907
rect -1748 37873 -1714 37907
rect -1680 37873 -1646 37907
rect -1612 37873 -1578 37907
rect -1544 37873 -1510 37907
rect -1476 37873 -1442 37907
rect -1408 37873 -1374 37907
rect -1340 37873 -1306 37907
rect -1272 37873 -1238 37907
rect -1204 37873 -1170 37907
rect -1136 37873 -1102 37907
rect -1068 37873 -1034 37907
rect -1000 37873 -966 37907
rect -932 37873 -898 37907
rect -864 37873 -830 37907
rect -796 37873 -762 37907
rect -728 37873 -694 37907
rect -660 37873 -626 37907
rect -592 37873 -558 37907
rect -524 37873 -490 37907
rect -456 37873 -422 37907
rect -388 37873 -354 37907
rect -320 37873 -286 37907
rect -252 37873 -218 37907
rect -184 37873 -153 37907
rect -2969 37838 -153 37873
rect -2969 37804 -2938 37838
rect -2904 37804 -2870 37838
rect -2836 37804 -2802 37838
rect -2768 37804 -2734 37838
rect -2700 37804 -2666 37838
rect -2632 37804 -2598 37838
rect -2564 37804 -2530 37838
rect -2496 37804 -2462 37838
rect -2428 37804 -2394 37838
rect -2360 37804 -2326 37838
rect -2292 37804 -2258 37838
rect -2224 37804 -2190 37838
rect -2156 37804 -2122 37838
rect -2088 37804 -2054 37838
rect -2020 37804 -1986 37838
rect -1952 37804 -1918 37838
rect -1884 37804 -1850 37838
rect -1816 37804 -1782 37838
rect -1748 37804 -1714 37838
rect -1680 37804 -1646 37838
rect -1612 37804 -1578 37838
rect -1544 37804 -1510 37838
rect -1476 37804 -1442 37838
rect -1408 37804 -1374 37838
rect -1340 37804 -1306 37838
rect -1272 37804 -1238 37838
rect -1204 37804 -1170 37838
rect -1136 37804 -1102 37838
rect -1068 37804 -1034 37838
rect -1000 37804 -966 37838
rect -932 37804 -898 37838
rect -864 37804 -830 37838
rect -796 37804 -762 37838
rect -728 37804 -694 37838
rect -660 37804 -626 37838
rect -592 37804 -558 37838
rect -524 37804 -490 37838
rect -456 37804 -422 37838
rect -388 37804 -354 37838
rect -320 37804 -286 37838
rect -252 37804 -218 37838
rect -184 37804 -153 37838
rect -2969 37769 -153 37804
rect -2969 37735 -2938 37769
rect -2904 37735 -2870 37769
rect -2836 37735 -2802 37769
rect -2768 37735 -2734 37769
rect -2700 37735 -2666 37769
rect -2632 37735 -2598 37769
rect -2564 37735 -2530 37769
rect -2496 37735 -2462 37769
rect -2428 37735 -2394 37769
rect -2360 37735 -2326 37769
rect -2292 37735 -2258 37769
rect -2224 37735 -2190 37769
rect -2156 37735 -2122 37769
rect -2088 37735 -2054 37769
rect -2020 37735 -1986 37769
rect -1952 37735 -1918 37769
rect -1884 37735 -1850 37769
rect -1816 37735 -1782 37769
rect -1748 37735 -1714 37769
rect -1680 37735 -1646 37769
rect -1612 37735 -1578 37769
rect -1544 37735 -1510 37769
rect -1476 37735 -1442 37769
rect -1408 37735 -1374 37769
rect -1340 37735 -1306 37769
rect -1272 37735 -1238 37769
rect -1204 37735 -1170 37769
rect -1136 37735 -1102 37769
rect -1068 37735 -1034 37769
rect -1000 37735 -966 37769
rect -932 37735 -898 37769
rect -864 37735 -830 37769
rect -796 37735 -762 37769
rect -728 37735 -694 37769
rect -660 37735 -626 37769
rect -592 37735 -558 37769
rect -524 37735 -490 37769
rect -456 37735 -422 37769
rect -388 37735 -354 37769
rect -320 37735 -286 37769
rect -252 37735 -218 37769
rect -184 37735 -153 37769
rect -2969 37700 -153 37735
rect -2969 37666 -2938 37700
rect -2904 37666 -2870 37700
rect -2836 37666 -2802 37700
rect -2768 37666 -2734 37700
rect -2700 37666 -2666 37700
rect -2632 37666 -2598 37700
rect -2564 37666 -2530 37700
rect -2496 37666 -2462 37700
rect -2428 37666 -2394 37700
rect -2360 37666 -2326 37700
rect -2292 37666 -2258 37700
rect -2224 37666 -2190 37700
rect -2156 37666 -2122 37700
rect -2088 37666 -2054 37700
rect -2020 37666 -1986 37700
rect -1952 37666 -1918 37700
rect -1884 37666 -1850 37700
rect -1816 37666 -1782 37700
rect -1748 37666 -1714 37700
rect -1680 37666 -1646 37700
rect -1612 37666 -1578 37700
rect -1544 37666 -1510 37700
rect -1476 37666 -1442 37700
rect -1408 37666 -1374 37700
rect -1340 37666 -1306 37700
rect -1272 37666 -1238 37700
rect -1204 37666 -1170 37700
rect -1136 37666 -1102 37700
rect -1068 37666 -1034 37700
rect -1000 37666 -966 37700
rect -932 37666 -898 37700
rect -864 37666 -830 37700
rect -796 37666 -762 37700
rect -728 37666 -694 37700
rect -660 37666 -626 37700
rect -592 37666 -558 37700
rect -524 37666 -490 37700
rect -456 37666 -422 37700
rect -388 37666 -354 37700
rect -320 37666 -286 37700
rect -252 37666 -218 37700
rect -184 37666 -153 37700
rect -2969 37631 -153 37666
rect -2969 37597 -2938 37631
rect -2904 37597 -2870 37631
rect -2836 37597 -2802 37631
rect -2768 37597 -2734 37631
rect -2700 37597 -2666 37631
rect -2632 37597 -2598 37631
rect -2564 37597 -2530 37631
rect -2496 37597 -2462 37631
rect -2428 37597 -2394 37631
rect -2360 37597 -2326 37631
rect -2292 37597 -2258 37631
rect -2224 37597 -2190 37631
rect -2156 37597 -2122 37631
rect -2088 37597 -2054 37631
rect -2020 37597 -1986 37631
rect -1952 37597 -1918 37631
rect -1884 37597 -1850 37631
rect -1816 37597 -1782 37631
rect -1748 37597 -1714 37631
rect -1680 37597 -1646 37631
rect -1612 37597 -1578 37631
rect -1544 37597 -1510 37631
rect -1476 37597 -1442 37631
rect -1408 37597 -1374 37631
rect -1340 37597 -1306 37631
rect -1272 37597 -1238 37631
rect -1204 37597 -1170 37631
rect -1136 37597 -1102 37631
rect -1068 37597 -1034 37631
rect -1000 37597 -966 37631
rect -932 37597 -898 37631
rect -864 37597 -830 37631
rect -796 37597 -762 37631
rect -728 37597 -694 37631
rect -660 37597 -626 37631
rect -592 37597 -558 37631
rect -524 37597 -490 37631
rect -456 37597 -422 37631
rect -388 37597 -354 37631
rect -320 37597 -286 37631
rect -252 37597 -218 37631
rect -184 37597 -153 37631
rect -2969 37562 -153 37597
rect -2969 37528 -2938 37562
rect -2904 37528 -2870 37562
rect -2836 37528 -2802 37562
rect -2768 37528 -2734 37562
rect -2700 37528 -2666 37562
rect -2632 37528 -2598 37562
rect -2564 37528 -2530 37562
rect -2496 37528 -2462 37562
rect -2428 37528 -2394 37562
rect -2360 37528 -2326 37562
rect -2292 37528 -2258 37562
rect -2224 37528 -2190 37562
rect -2156 37528 -2122 37562
rect -2088 37528 -2054 37562
rect -2020 37528 -1986 37562
rect -1952 37528 -1918 37562
rect -1884 37528 -1850 37562
rect -1816 37528 -1782 37562
rect -1748 37528 -1714 37562
rect -1680 37528 -1646 37562
rect -1612 37528 -1578 37562
rect -1544 37528 -1510 37562
rect -1476 37528 -1442 37562
rect -1408 37528 -1374 37562
rect -1340 37528 -1306 37562
rect -1272 37528 -1238 37562
rect -1204 37528 -1170 37562
rect -1136 37528 -1102 37562
rect -1068 37528 -1034 37562
rect -1000 37528 -966 37562
rect -932 37528 -898 37562
rect -864 37528 -830 37562
rect -796 37528 -762 37562
rect -728 37528 -694 37562
rect -660 37528 -626 37562
rect -592 37528 -558 37562
rect -524 37528 -490 37562
rect -456 37528 -422 37562
rect -388 37528 -354 37562
rect -320 37528 -286 37562
rect -252 37528 -218 37562
rect -184 37528 -153 37562
rect -2969 37493 -153 37528
rect -2969 37459 -2938 37493
rect -2904 37459 -2870 37493
rect -2836 37459 -2802 37493
rect -2768 37459 -2734 37493
rect -2700 37459 -2666 37493
rect -2632 37459 -2598 37493
rect -2564 37459 -2530 37493
rect -2496 37459 -2462 37493
rect -2428 37459 -2394 37493
rect -2360 37459 -2326 37493
rect -2292 37459 -2258 37493
rect -2224 37459 -2190 37493
rect -2156 37459 -2122 37493
rect -2088 37459 -2054 37493
rect -2020 37459 -1986 37493
rect -1952 37459 -1918 37493
rect -1884 37459 -1850 37493
rect -1816 37459 -1782 37493
rect -1748 37459 -1714 37493
rect -1680 37459 -1646 37493
rect -1612 37459 -1578 37493
rect -1544 37459 -1510 37493
rect -1476 37459 -1442 37493
rect -1408 37459 -1374 37493
rect -1340 37459 -1306 37493
rect -1272 37459 -1238 37493
rect -1204 37459 -1170 37493
rect -1136 37459 -1102 37493
rect -1068 37459 -1034 37493
rect -1000 37459 -966 37493
rect -932 37459 -898 37493
rect -864 37459 -830 37493
rect -796 37459 -762 37493
rect -728 37459 -694 37493
rect -660 37459 -626 37493
rect -592 37459 -558 37493
rect -524 37459 -490 37493
rect -456 37459 -422 37493
rect -388 37459 -354 37493
rect -320 37459 -286 37493
rect -252 37459 -218 37493
rect -184 37459 -153 37493
rect -2969 37424 -153 37459
rect -2969 37390 -2938 37424
rect -2904 37390 -2870 37424
rect -2836 37390 -2802 37424
rect -2768 37390 -2734 37424
rect -2700 37390 -2666 37424
rect -2632 37390 -2598 37424
rect -2564 37390 -2530 37424
rect -2496 37390 -2462 37424
rect -2428 37390 -2394 37424
rect -2360 37390 -2326 37424
rect -2292 37390 -2258 37424
rect -2224 37390 -2190 37424
rect -2156 37390 -2122 37424
rect -2088 37390 -2054 37424
rect -2020 37390 -1986 37424
rect -1952 37390 -1918 37424
rect -1884 37390 -1850 37424
rect -1816 37390 -1782 37424
rect -1748 37390 -1714 37424
rect -1680 37390 -1646 37424
rect -1612 37390 -1578 37424
rect -1544 37390 -1510 37424
rect -1476 37390 -1442 37424
rect -1408 37390 -1374 37424
rect -1340 37390 -1306 37424
rect -1272 37390 -1238 37424
rect -1204 37390 -1170 37424
rect -1136 37390 -1102 37424
rect -1068 37390 -1034 37424
rect -1000 37390 -966 37424
rect -932 37390 -898 37424
rect -864 37390 -830 37424
rect -796 37390 -762 37424
rect -728 37390 -694 37424
rect -660 37390 -626 37424
rect -592 37390 -558 37424
rect -524 37390 -490 37424
rect -456 37390 -422 37424
rect -388 37390 -354 37424
rect -320 37390 -286 37424
rect -252 37390 -218 37424
rect -184 37390 -153 37424
rect -2969 37355 -153 37390
rect -2969 37321 -2938 37355
rect -2904 37321 -2870 37355
rect -2836 37321 -2802 37355
rect -2768 37321 -2734 37355
rect -2700 37321 -2666 37355
rect -2632 37321 -2598 37355
rect -2564 37321 -2530 37355
rect -2496 37321 -2462 37355
rect -2428 37321 -2394 37355
rect -2360 37321 -2326 37355
rect -2292 37321 -2258 37355
rect -2224 37321 -2190 37355
rect -2156 37321 -2122 37355
rect -2088 37321 -2054 37355
rect -2020 37321 -1986 37355
rect -1952 37321 -1918 37355
rect -1884 37321 -1850 37355
rect -1816 37321 -1782 37355
rect -1748 37321 -1714 37355
rect -1680 37321 -1646 37355
rect -1612 37321 -1578 37355
rect -1544 37321 -1510 37355
rect -1476 37321 -1442 37355
rect -1408 37321 -1374 37355
rect -1340 37321 -1306 37355
rect -1272 37321 -1238 37355
rect -1204 37321 -1170 37355
rect -1136 37321 -1102 37355
rect -1068 37321 -1034 37355
rect -1000 37321 -966 37355
rect -932 37321 -898 37355
rect -864 37321 -830 37355
rect -796 37321 -762 37355
rect -728 37321 -694 37355
rect -660 37321 -626 37355
rect -592 37321 -558 37355
rect -524 37321 -490 37355
rect -456 37321 -422 37355
rect -388 37321 -354 37355
rect -320 37321 -286 37355
rect -252 37321 -218 37355
rect -184 37321 -153 37355
rect -2969 37286 -153 37321
rect -2969 37252 -2938 37286
rect -2904 37252 -2870 37286
rect -2836 37252 -2802 37286
rect -2768 37252 -2734 37286
rect -2700 37252 -2666 37286
rect -2632 37252 -2598 37286
rect -2564 37252 -2530 37286
rect -2496 37252 -2462 37286
rect -2428 37252 -2394 37286
rect -2360 37252 -2326 37286
rect -2292 37252 -2258 37286
rect -2224 37252 -2190 37286
rect -2156 37252 -2122 37286
rect -2088 37252 -2054 37286
rect -2020 37252 -1986 37286
rect -1952 37252 -1918 37286
rect -1884 37252 -1850 37286
rect -1816 37252 -1782 37286
rect -1748 37252 -1714 37286
rect -1680 37252 -1646 37286
rect -1612 37252 -1578 37286
rect -1544 37252 -1510 37286
rect -1476 37252 -1442 37286
rect -1408 37252 -1374 37286
rect -1340 37252 -1306 37286
rect -1272 37252 -1238 37286
rect -1204 37252 -1170 37286
rect -1136 37252 -1102 37286
rect -1068 37252 -1034 37286
rect -1000 37252 -966 37286
rect -932 37252 -898 37286
rect -864 37252 -830 37286
rect -796 37252 -762 37286
rect -728 37252 -694 37286
rect -660 37252 -626 37286
rect -592 37252 -558 37286
rect -524 37252 -490 37286
rect -456 37252 -422 37286
rect -388 37252 -354 37286
rect -320 37252 -286 37286
rect -252 37252 -218 37286
rect -184 37252 -153 37286
rect -2969 37217 -153 37252
rect -2969 37183 -2938 37217
rect -2904 37183 -2870 37217
rect -2836 37183 -2802 37217
rect -2768 37183 -2734 37217
rect -2700 37183 -2666 37217
rect -2632 37183 -2598 37217
rect -2564 37183 -2530 37217
rect -2496 37183 -2462 37217
rect -2428 37183 -2394 37217
rect -2360 37183 -2326 37217
rect -2292 37183 -2258 37217
rect -2224 37183 -2190 37217
rect -2156 37183 -2122 37217
rect -2088 37183 -2054 37217
rect -2020 37183 -1986 37217
rect -1952 37183 -1918 37217
rect -1884 37183 -1850 37217
rect -1816 37183 -1782 37217
rect -1748 37183 -1714 37217
rect -1680 37183 -1646 37217
rect -1612 37183 -1578 37217
rect -1544 37183 -1510 37217
rect -1476 37183 -1442 37217
rect -1408 37183 -1374 37217
rect -1340 37183 -1306 37217
rect -1272 37183 -1238 37217
rect -1204 37183 -1170 37217
rect -1136 37183 -1102 37217
rect -1068 37183 -1034 37217
rect -1000 37183 -966 37217
rect -932 37183 -898 37217
rect -864 37183 -830 37217
rect -796 37183 -762 37217
rect -728 37183 -694 37217
rect -660 37183 -626 37217
rect -592 37183 -558 37217
rect -524 37183 -490 37217
rect -456 37183 -422 37217
rect -388 37183 -354 37217
rect -320 37183 -286 37217
rect -252 37183 -218 37217
rect -184 37183 -153 37217
rect -2969 37148 -153 37183
rect -2969 37114 -2938 37148
rect -2904 37114 -2870 37148
rect -2836 37114 -2802 37148
rect -2768 37114 -2734 37148
rect -2700 37114 -2666 37148
rect -2632 37114 -2598 37148
rect -2564 37114 -2530 37148
rect -2496 37114 -2462 37148
rect -2428 37114 -2394 37148
rect -2360 37114 -2326 37148
rect -2292 37114 -2258 37148
rect -2224 37114 -2190 37148
rect -2156 37114 -2122 37148
rect -2088 37114 -2054 37148
rect -2020 37114 -1986 37148
rect -1952 37114 -1918 37148
rect -1884 37114 -1850 37148
rect -1816 37114 -1782 37148
rect -1748 37114 -1714 37148
rect -1680 37114 -1646 37148
rect -1612 37114 -1578 37148
rect -1544 37114 -1510 37148
rect -1476 37114 -1442 37148
rect -1408 37114 -1374 37148
rect -1340 37114 -1306 37148
rect -1272 37114 -1238 37148
rect -1204 37114 -1170 37148
rect -1136 37114 -1102 37148
rect -1068 37114 -1034 37148
rect -1000 37114 -966 37148
rect -932 37114 -898 37148
rect -864 37114 -830 37148
rect -796 37114 -762 37148
rect -728 37114 -694 37148
rect -660 37114 -626 37148
rect -592 37114 -558 37148
rect -524 37114 -490 37148
rect -456 37114 -422 37148
rect -388 37114 -354 37148
rect -320 37114 -286 37148
rect -252 37114 -218 37148
rect -184 37114 -153 37148
rect -2969 37079 -153 37114
rect -2969 37045 -2938 37079
rect -2904 37045 -2870 37079
rect -2836 37045 -2802 37079
rect -2768 37045 -2734 37079
rect -2700 37045 -2666 37079
rect -2632 37045 -2598 37079
rect -2564 37045 -2530 37079
rect -2496 37045 -2462 37079
rect -2428 37045 -2394 37079
rect -2360 37045 -2326 37079
rect -2292 37045 -2258 37079
rect -2224 37045 -2190 37079
rect -2156 37045 -2122 37079
rect -2088 37045 -2054 37079
rect -2020 37045 -1986 37079
rect -1952 37045 -1918 37079
rect -1884 37045 -1850 37079
rect -1816 37045 -1782 37079
rect -1748 37045 -1714 37079
rect -1680 37045 -1646 37079
rect -1612 37045 -1578 37079
rect -1544 37045 -1510 37079
rect -1476 37045 -1442 37079
rect -1408 37045 -1374 37079
rect -1340 37045 -1306 37079
rect -1272 37045 -1238 37079
rect -1204 37045 -1170 37079
rect -1136 37045 -1102 37079
rect -1068 37045 -1034 37079
rect -1000 37045 -966 37079
rect -932 37045 -898 37079
rect -864 37045 -830 37079
rect -796 37045 -762 37079
rect -728 37045 -694 37079
rect -660 37045 -626 37079
rect -592 37045 -558 37079
rect -524 37045 -490 37079
rect -456 37045 -422 37079
rect -388 37045 -354 37079
rect -320 37045 -286 37079
rect -252 37045 -218 37079
rect -184 37045 -153 37079
rect -2969 37010 -153 37045
rect -2969 36976 -2938 37010
rect -2904 36976 -2870 37010
rect -2836 36976 -2802 37010
rect -2768 36976 -2734 37010
rect -2700 36976 -2666 37010
rect -2632 36976 -2598 37010
rect -2564 36976 -2530 37010
rect -2496 36976 -2462 37010
rect -2428 36976 -2394 37010
rect -2360 36976 -2326 37010
rect -2292 36976 -2258 37010
rect -2224 36976 -2190 37010
rect -2156 36976 -2122 37010
rect -2088 36976 -2054 37010
rect -2020 36976 -1986 37010
rect -1952 36976 -1918 37010
rect -1884 36976 -1850 37010
rect -1816 36976 -1782 37010
rect -1748 36976 -1714 37010
rect -1680 36976 -1646 37010
rect -1612 36976 -1578 37010
rect -1544 36976 -1510 37010
rect -1476 36976 -1442 37010
rect -1408 36976 -1374 37010
rect -1340 36976 -1306 37010
rect -1272 36976 -1238 37010
rect -1204 36976 -1170 37010
rect -1136 36976 -1102 37010
rect -1068 36976 -1034 37010
rect -1000 36976 -966 37010
rect -932 36976 -898 37010
rect -864 36976 -830 37010
rect -796 36976 -762 37010
rect -728 36976 -694 37010
rect -660 36976 -626 37010
rect -592 36976 -558 37010
rect -524 36976 -490 37010
rect -456 36976 -422 37010
rect -388 36976 -354 37010
rect -320 36976 -286 37010
rect -252 36976 -218 37010
rect -184 36976 -153 37010
rect -2969 36941 -153 36976
rect -2969 36907 -2938 36941
rect -2904 36907 -2870 36941
rect -2836 36907 -2802 36941
rect -2768 36907 -2734 36941
rect -2700 36907 -2666 36941
rect -2632 36907 -2598 36941
rect -2564 36907 -2530 36941
rect -2496 36907 -2462 36941
rect -2428 36907 -2394 36941
rect -2360 36907 -2326 36941
rect -2292 36907 -2258 36941
rect -2224 36907 -2190 36941
rect -2156 36907 -2122 36941
rect -2088 36907 -2054 36941
rect -2020 36907 -1986 36941
rect -1952 36907 -1918 36941
rect -1884 36907 -1850 36941
rect -1816 36907 -1782 36941
rect -1748 36907 -1714 36941
rect -1680 36907 -1646 36941
rect -1612 36907 -1578 36941
rect -1544 36907 -1510 36941
rect -1476 36907 -1442 36941
rect -1408 36907 -1374 36941
rect -1340 36907 -1306 36941
rect -1272 36907 -1238 36941
rect -1204 36907 -1170 36941
rect -1136 36907 -1102 36941
rect -1068 36907 -1034 36941
rect -1000 36907 -966 36941
rect -932 36907 -898 36941
rect -864 36907 -830 36941
rect -796 36907 -762 36941
rect -728 36907 -694 36941
rect -660 36907 -626 36941
rect -592 36907 -558 36941
rect -524 36907 -490 36941
rect -456 36907 -422 36941
rect -388 36907 -354 36941
rect -320 36907 -286 36941
rect -252 36907 -218 36941
rect -184 36907 -153 36941
rect -2969 36872 -153 36907
rect -2969 36838 -2938 36872
rect -2904 36838 -2870 36872
rect -2836 36838 -2802 36872
rect -2768 36838 -2734 36872
rect -2700 36838 -2666 36872
rect -2632 36838 -2598 36872
rect -2564 36838 -2530 36872
rect -2496 36838 -2462 36872
rect -2428 36838 -2394 36872
rect -2360 36838 -2326 36872
rect -2292 36838 -2258 36872
rect -2224 36838 -2190 36872
rect -2156 36838 -2122 36872
rect -2088 36838 -2054 36872
rect -2020 36838 -1986 36872
rect -1952 36838 -1918 36872
rect -1884 36838 -1850 36872
rect -1816 36838 -1782 36872
rect -1748 36838 -1714 36872
rect -1680 36838 -1646 36872
rect -1612 36838 -1578 36872
rect -1544 36838 -1510 36872
rect -1476 36838 -1442 36872
rect -1408 36838 -1374 36872
rect -1340 36838 -1306 36872
rect -1272 36838 -1238 36872
rect -1204 36838 -1170 36872
rect -1136 36838 -1102 36872
rect -1068 36838 -1034 36872
rect -1000 36838 -966 36872
rect -932 36838 -898 36872
rect -864 36838 -830 36872
rect -796 36838 -762 36872
rect -728 36838 -694 36872
rect -660 36838 -626 36872
rect -592 36838 -558 36872
rect -524 36838 -490 36872
rect -456 36838 -422 36872
rect -388 36838 -354 36872
rect -320 36838 -286 36872
rect -252 36838 -218 36872
rect -184 36838 -153 36872
rect -2969 36803 -153 36838
rect -2969 36769 -2938 36803
rect -2904 36769 -2870 36803
rect -2836 36769 -2802 36803
rect -2768 36769 -2734 36803
rect -2700 36769 -2666 36803
rect -2632 36769 -2598 36803
rect -2564 36769 -2530 36803
rect -2496 36769 -2462 36803
rect -2428 36769 -2394 36803
rect -2360 36769 -2326 36803
rect -2292 36769 -2258 36803
rect -2224 36769 -2190 36803
rect -2156 36769 -2122 36803
rect -2088 36769 -2054 36803
rect -2020 36769 -1986 36803
rect -1952 36769 -1918 36803
rect -1884 36769 -1850 36803
rect -1816 36769 -1782 36803
rect -1748 36769 -1714 36803
rect -1680 36769 -1646 36803
rect -1612 36769 -1578 36803
rect -1544 36769 -1510 36803
rect -1476 36769 -1442 36803
rect -1408 36769 -1374 36803
rect -1340 36769 -1306 36803
rect -1272 36769 -1238 36803
rect -1204 36769 -1170 36803
rect -1136 36769 -1102 36803
rect -1068 36769 -1034 36803
rect -1000 36769 -966 36803
rect -932 36769 -898 36803
rect -864 36769 -830 36803
rect -796 36769 -762 36803
rect -728 36769 -694 36803
rect -660 36769 -626 36803
rect -592 36769 -558 36803
rect -524 36769 -490 36803
rect -456 36769 -422 36803
rect -388 36769 -354 36803
rect -320 36769 -286 36803
rect -252 36769 -218 36803
rect -184 36769 -153 36803
rect -2969 36734 -153 36769
rect -2969 36700 -2938 36734
rect -2904 36700 -2870 36734
rect -2836 36700 -2802 36734
rect -2768 36700 -2734 36734
rect -2700 36700 -2666 36734
rect -2632 36700 -2598 36734
rect -2564 36700 -2530 36734
rect -2496 36700 -2462 36734
rect -2428 36700 -2394 36734
rect -2360 36700 -2326 36734
rect -2292 36700 -2258 36734
rect -2224 36700 -2190 36734
rect -2156 36700 -2122 36734
rect -2088 36700 -2054 36734
rect -2020 36700 -1986 36734
rect -1952 36700 -1918 36734
rect -1884 36700 -1850 36734
rect -1816 36700 -1782 36734
rect -1748 36700 -1714 36734
rect -1680 36700 -1646 36734
rect -1612 36700 -1578 36734
rect -1544 36700 -1510 36734
rect -1476 36700 -1442 36734
rect -1408 36700 -1374 36734
rect -1340 36700 -1306 36734
rect -1272 36700 -1238 36734
rect -1204 36700 -1170 36734
rect -1136 36700 -1102 36734
rect -1068 36700 -1034 36734
rect -1000 36700 -966 36734
rect -932 36700 -898 36734
rect -864 36700 -830 36734
rect -796 36700 -762 36734
rect -728 36700 -694 36734
rect -660 36700 -626 36734
rect -592 36700 -558 36734
rect -524 36700 -490 36734
rect -456 36700 -422 36734
rect -388 36700 -354 36734
rect -320 36700 -286 36734
rect -252 36700 -218 36734
rect -184 36700 -153 36734
rect -2969 36665 -153 36700
rect -2969 36631 -2938 36665
rect -2904 36631 -2870 36665
rect -2836 36631 -2802 36665
rect -2768 36631 -2734 36665
rect -2700 36631 -2666 36665
rect -2632 36631 -2598 36665
rect -2564 36631 -2530 36665
rect -2496 36631 -2462 36665
rect -2428 36631 -2394 36665
rect -2360 36631 -2326 36665
rect -2292 36631 -2258 36665
rect -2224 36631 -2190 36665
rect -2156 36631 -2122 36665
rect -2088 36631 -2054 36665
rect -2020 36631 -1986 36665
rect -1952 36631 -1918 36665
rect -1884 36631 -1850 36665
rect -1816 36631 -1782 36665
rect -1748 36631 -1714 36665
rect -1680 36631 -1646 36665
rect -1612 36631 -1578 36665
rect -1544 36631 -1510 36665
rect -1476 36631 -1442 36665
rect -1408 36631 -1374 36665
rect -1340 36631 -1306 36665
rect -1272 36631 -1238 36665
rect -1204 36631 -1170 36665
rect -1136 36631 -1102 36665
rect -1068 36631 -1034 36665
rect -1000 36631 -966 36665
rect -932 36631 -898 36665
rect -864 36631 -830 36665
rect -796 36631 -762 36665
rect -728 36631 -694 36665
rect -660 36631 -626 36665
rect -592 36631 -558 36665
rect -524 36631 -490 36665
rect -456 36631 -422 36665
rect -388 36631 -354 36665
rect -320 36631 -286 36665
rect -252 36631 -218 36665
rect -184 36631 -153 36665
rect -2969 36596 -153 36631
rect -2969 36562 -2938 36596
rect -2904 36562 -2870 36596
rect -2836 36562 -2802 36596
rect -2768 36562 -2734 36596
rect -2700 36562 -2666 36596
rect -2632 36562 -2598 36596
rect -2564 36562 -2530 36596
rect -2496 36562 -2462 36596
rect -2428 36562 -2394 36596
rect -2360 36562 -2326 36596
rect -2292 36562 -2258 36596
rect -2224 36562 -2190 36596
rect -2156 36562 -2122 36596
rect -2088 36562 -2054 36596
rect -2020 36562 -1986 36596
rect -1952 36562 -1918 36596
rect -1884 36562 -1850 36596
rect -1816 36562 -1782 36596
rect -1748 36562 -1714 36596
rect -1680 36562 -1646 36596
rect -1612 36562 -1578 36596
rect -1544 36562 -1510 36596
rect -1476 36562 -1442 36596
rect -1408 36562 -1374 36596
rect -1340 36562 -1306 36596
rect -1272 36562 -1238 36596
rect -1204 36562 -1170 36596
rect -1136 36562 -1102 36596
rect -1068 36562 -1034 36596
rect -1000 36562 -966 36596
rect -932 36562 -898 36596
rect -864 36562 -830 36596
rect -796 36562 -762 36596
rect -728 36562 -694 36596
rect -660 36562 -626 36596
rect -592 36562 -558 36596
rect -524 36562 -490 36596
rect -456 36562 -422 36596
rect -388 36562 -354 36596
rect -320 36562 -286 36596
rect -252 36562 -218 36596
rect -184 36562 -153 36596
rect -2969 36527 -153 36562
rect -2969 36493 -2938 36527
rect -2904 36493 -2870 36527
rect -2836 36493 -2802 36527
rect -2768 36493 -2734 36527
rect -2700 36493 -2666 36527
rect -2632 36493 -2598 36527
rect -2564 36493 -2530 36527
rect -2496 36493 -2462 36527
rect -2428 36493 -2394 36527
rect -2360 36493 -2326 36527
rect -2292 36493 -2258 36527
rect -2224 36493 -2190 36527
rect -2156 36493 -2122 36527
rect -2088 36493 -2054 36527
rect -2020 36493 -1986 36527
rect -1952 36493 -1918 36527
rect -1884 36493 -1850 36527
rect -1816 36493 -1782 36527
rect -1748 36493 -1714 36527
rect -1680 36493 -1646 36527
rect -1612 36493 -1578 36527
rect -1544 36493 -1510 36527
rect -1476 36493 -1442 36527
rect -1408 36493 -1374 36527
rect -1340 36493 -1306 36527
rect -1272 36493 -1238 36527
rect -1204 36493 -1170 36527
rect -1136 36493 -1102 36527
rect -1068 36493 -1034 36527
rect -1000 36493 -966 36527
rect -932 36493 -898 36527
rect -864 36493 -830 36527
rect -796 36493 -762 36527
rect -728 36493 -694 36527
rect -660 36493 -626 36527
rect -592 36493 -558 36527
rect -524 36493 -490 36527
rect -456 36493 -422 36527
rect -388 36493 -354 36527
rect -320 36493 -286 36527
rect -252 36493 -218 36527
rect -184 36493 -153 36527
rect -2969 36458 -153 36493
rect -2969 36424 -2938 36458
rect -2904 36424 -2870 36458
rect -2836 36424 -2802 36458
rect -2768 36424 -2734 36458
rect -2700 36424 -2666 36458
rect -2632 36424 -2598 36458
rect -2564 36424 -2530 36458
rect -2496 36424 -2462 36458
rect -2428 36424 -2394 36458
rect -2360 36424 -2326 36458
rect -2292 36424 -2258 36458
rect -2224 36424 -2190 36458
rect -2156 36424 -2122 36458
rect -2088 36424 -2054 36458
rect -2020 36424 -1986 36458
rect -1952 36424 -1918 36458
rect -1884 36424 -1850 36458
rect -1816 36424 -1782 36458
rect -1748 36424 -1714 36458
rect -1680 36424 -1646 36458
rect -1612 36424 -1578 36458
rect -1544 36424 -1510 36458
rect -1476 36424 -1442 36458
rect -1408 36424 -1374 36458
rect -1340 36424 -1306 36458
rect -1272 36424 -1238 36458
rect -1204 36424 -1170 36458
rect -1136 36424 -1102 36458
rect -1068 36424 -1034 36458
rect -1000 36424 -966 36458
rect -932 36424 -898 36458
rect -864 36424 -830 36458
rect -796 36424 -762 36458
rect -728 36424 -694 36458
rect -660 36424 -626 36458
rect -592 36424 -558 36458
rect -524 36424 -490 36458
rect -456 36424 -422 36458
rect -388 36424 -354 36458
rect -320 36424 -286 36458
rect -252 36424 -218 36458
rect -184 36424 -153 36458
rect -2969 36389 -153 36424
rect -2969 36355 -2938 36389
rect -2904 36355 -2870 36389
rect -2836 36355 -2802 36389
rect -2768 36355 -2734 36389
rect -2700 36355 -2666 36389
rect -2632 36355 -2598 36389
rect -2564 36355 -2530 36389
rect -2496 36355 -2462 36389
rect -2428 36355 -2394 36389
rect -2360 36355 -2326 36389
rect -2292 36355 -2258 36389
rect -2224 36355 -2190 36389
rect -2156 36355 -2122 36389
rect -2088 36355 -2054 36389
rect -2020 36355 -1986 36389
rect -1952 36355 -1918 36389
rect -1884 36355 -1850 36389
rect -1816 36355 -1782 36389
rect -1748 36355 -1714 36389
rect -1680 36355 -1646 36389
rect -1612 36355 -1578 36389
rect -1544 36355 -1510 36389
rect -1476 36355 -1442 36389
rect -1408 36355 -1374 36389
rect -1340 36355 -1306 36389
rect -1272 36355 -1238 36389
rect -1204 36355 -1170 36389
rect -1136 36355 -1102 36389
rect -1068 36355 -1034 36389
rect -1000 36355 -966 36389
rect -932 36355 -898 36389
rect -864 36355 -830 36389
rect -796 36355 -762 36389
rect -728 36355 -694 36389
rect -660 36355 -626 36389
rect -592 36355 -558 36389
rect -524 36355 -490 36389
rect -456 36355 -422 36389
rect -388 36355 -354 36389
rect -320 36355 -286 36389
rect -252 36355 -218 36389
rect -184 36355 -153 36389
rect -2969 36320 -153 36355
rect -2969 36286 -2938 36320
rect -2904 36286 -2870 36320
rect -2836 36286 -2802 36320
rect -2768 36286 -2734 36320
rect -2700 36286 -2666 36320
rect -2632 36286 -2598 36320
rect -2564 36286 -2530 36320
rect -2496 36286 -2462 36320
rect -2428 36286 -2394 36320
rect -2360 36286 -2326 36320
rect -2292 36286 -2258 36320
rect -2224 36286 -2190 36320
rect -2156 36286 -2122 36320
rect -2088 36286 -2054 36320
rect -2020 36286 -1986 36320
rect -1952 36286 -1918 36320
rect -1884 36286 -1850 36320
rect -1816 36286 -1782 36320
rect -1748 36286 -1714 36320
rect -1680 36286 -1646 36320
rect -1612 36286 -1578 36320
rect -1544 36286 -1510 36320
rect -1476 36286 -1442 36320
rect -1408 36286 -1374 36320
rect -1340 36286 -1306 36320
rect -1272 36286 -1238 36320
rect -1204 36286 -1170 36320
rect -1136 36286 -1102 36320
rect -1068 36286 -1034 36320
rect -1000 36286 -966 36320
rect -932 36286 -898 36320
rect -864 36286 -830 36320
rect -796 36286 -762 36320
rect -728 36286 -694 36320
rect -660 36286 -626 36320
rect -592 36286 -558 36320
rect -524 36286 -490 36320
rect -456 36286 -422 36320
rect -388 36286 -354 36320
rect -320 36286 -286 36320
rect -252 36286 -218 36320
rect -184 36286 -153 36320
rect -2969 36251 -153 36286
rect -2969 36217 -2938 36251
rect -2904 36217 -2870 36251
rect -2836 36217 -2802 36251
rect -2768 36217 -2734 36251
rect -2700 36217 -2666 36251
rect -2632 36217 -2598 36251
rect -2564 36217 -2530 36251
rect -2496 36217 -2462 36251
rect -2428 36217 -2394 36251
rect -2360 36217 -2326 36251
rect -2292 36217 -2258 36251
rect -2224 36217 -2190 36251
rect -2156 36217 -2122 36251
rect -2088 36217 -2054 36251
rect -2020 36217 -1986 36251
rect -1952 36217 -1918 36251
rect -1884 36217 -1850 36251
rect -1816 36217 -1782 36251
rect -1748 36217 -1714 36251
rect -1680 36217 -1646 36251
rect -1612 36217 -1578 36251
rect -1544 36217 -1510 36251
rect -1476 36217 -1442 36251
rect -1408 36217 -1374 36251
rect -1340 36217 -1306 36251
rect -1272 36217 -1238 36251
rect -1204 36217 -1170 36251
rect -1136 36217 -1102 36251
rect -1068 36217 -1034 36251
rect -1000 36217 -966 36251
rect -932 36217 -898 36251
rect -864 36217 -830 36251
rect -796 36217 -762 36251
rect -728 36217 -694 36251
rect -660 36217 -626 36251
rect -592 36217 -558 36251
rect -524 36217 -490 36251
rect -456 36217 -422 36251
rect -388 36217 -354 36251
rect -320 36217 -286 36251
rect -252 36217 -218 36251
rect -184 36217 -153 36251
rect -2969 36182 -153 36217
rect -2969 36148 -2938 36182
rect -2904 36148 -2870 36182
rect -2836 36148 -2802 36182
rect -2768 36148 -2734 36182
rect -2700 36148 -2666 36182
rect -2632 36148 -2598 36182
rect -2564 36148 -2530 36182
rect -2496 36148 -2462 36182
rect -2428 36148 -2394 36182
rect -2360 36148 -2326 36182
rect -2292 36148 -2258 36182
rect -2224 36148 -2190 36182
rect -2156 36148 -2122 36182
rect -2088 36148 -2054 36182
rect -2020 36148 -1986 36182
rect -1952 36148 -1918 36182
rect -1884 36148 -1850 36182
rect -1816 36148 -1782 36182
rect -1748 36148 -1714 36182
rect -1680 36148 -1646 36182
rect -1612 36148 -1578 36182
rect -1544 36148 -1510 36182
rect -1476 36148 -1442 36182
rect -1408 36148 -1374 36182
rect -1340 36148 -1306 36182
rect -1272 36148 -1238 36182
rect -1204 36148 -1170 36182
rect -1136 36148 -1102 36182
rect -1068 36148 -1034 36182
rect -1000 36148 -966 36182
rect -932 36148 -898 36182
rect -864 36148 -830 36182
rect -796 36148 -762 36182
rect -728 36148 -694 36182
rect -660 36148 -626 36182
rect -592 36148 -558 36182
rect -524 36148 -490 36182
rect -456 36148 -422 36182
rect -388 36148 -354 36182
rect -320 36148 -286 36182
rect -252 36148 -218 36182
rect -184 36148 -153 36182
rect -2969 36113 -153 36148
rect -2969 36079 -2938 36113
rect -2904 36079 -2870 36113
rect -2836 36079 -2802 36113
rect -2768 36079 -2734 36113
rect -2700 36079 -2666 36113
rect -2632 36079 -2598 36113
rect -2564 36079 -2530 36113
rect -2496 36079 -2462 36113
rect -2428 36079 -2394 36113
rect -2360 36079 -2326 36113
rect -2292 36079 -2258 36113
rect -2224 36079 -2190 36113
rect -2156 36079 -2122 36113
rect -2088 36079 -2054 36113
rect -2020 36079 -1986 36113
rect -1952 36079 -1918 36113
rect -1884 36079 -1850 36113
rect -1816 36079 -1782 36113
rect -1748 36079 -1714 36113
rect -1680 36079 -1646 36113
rect -1612 36079 -1578 36113
rect -1544 36079 -1510 36113
rect -1476 36079 -1442 36113
rect -1408 36079 -1374 36113
rect -1340 36079 -1306 36113
rect -1272 36079 -1238 36113
rect -1204 36079 -1170 36113
rect -1136 36079 -1102 36113
rect -1068 36079 -1034 36113
rect -1000 36079 -966 36113
rect -932 36079 -898 36113
rect -864 36079 -830 36113
rect -796 36079 -762 36113
rect -728 36079 -694 36113
rect -660 36079 -626 36113
rect -592 36079 -558 36113
rect -524 36079 -490 36113
rect -456 36079 -422 36113
rect -388 36079 -354 36113
rect -320 36079 -286 36113
rect -252 36079 -218 36113
rect -184 36079 -153 36113
rect -2969 36044 -153 36079
rect -2969 36010 -2938 36044
rect -2904 36010 -2870 36044
rect -2836 36010 -2802 36044
rect -2768 36010 -2734 36044
rect -2700 36010 -2666 36044
rect -2632 36010 -2598 36044
rect -2564 36010 -2530 36044
rect -2496 36010 -2462 36044
rect -2428 36010 -2394 36044
rect -2360 36010 -2326 36044
rect -2292 36010 -2258 36044
rect -2224 36010 -2190 36044
rect -2156 36010 -2122 36044
rect -2088 36010 -2054 36044
rect -2020 36010 -1986 36044
rect -1952 36010 -1918 36044
rect -1884 36010 -1850 36044
rect -1816 36010 -1782 36044
rect -1748 36010 -1714 36044
rect -1680 36010 -1646 36044
rect -1612 36010 -1578 36044
rect -1544 36010 -1510 36044
rect -1476 36010 -1442 36044
rect -1408 36010 -1374 36044
rect -1340 36010 -1306 36044
rect -1272 36010 -1238 36044
rect -1204 36010 -1170 36044
rect -1136 36010 -1102 36044
rect -1068 36010 -1034 36044
rect -1000 36010 -966 36044
rect -932 36010 -898 36044
rect -864 36010 -830 36044
rect -796 36010 -762 36044
rect -728 36010 -694 36044
rect -660 36010 -626 36044
rect -592 36010 -558 36044
rect -524 36010 -490 36044
rect -456 36010 -422 36044
rect -388 36010 -354 36044
rect -320 36010 -286 36044
rect -252 36010 -218 36044
rect -184 36010 -153 36044
rect -2969 35975 -153 36010
rect -2969 35941 -2938 35975
rect -2904 35941 -2870 35975
rect -2836 35941 -2802 35975
rect -2768 35941 -2734 35975
rect -2700 35941 -2666 35975
rect -2632 35941 -2598 35975
rect -2564 35941 -2530 35975
rect -2496 35941 -2462 35975
rect -2428 35941 -2394 35975
rect -2360 35941 -2326 35975
rect -2292 35941 -2258 35975
rect -2224 35941 -2190 35975
rect -2156 35941 -2122 35975
rect -2088 35941 -2054 35975
rect -2020 35941 -1986 35975
rect -1952 35941 -1918 35975
rect -1884 35941 -1850 35975
rect -1816 35941 -1782 35975
rect -1748 35941 -1714 35975
rect -1680 35941 -1646 35975
rect -1612 35941 -1578 35975
rect -1544 35941 -1510 35975
rect -1476 35941 -1442 35975
rect -1408 35941 -1374 35975
rect -1340 35941 -1306 35975
rect -1272 35941 -1238 35975
rect -1204 35941 -1170 35975
rect -1136 35941 -1102 35975
rect -1068 35941 -1034 35975
rect -1000 35941 -966 35975
rect -932 35941 -898 35975
rect -864 35941 -830 35975
rect -796 35941 -762 35975
rect -728 35941 -694 35975
rect -660 35941 -626 35975
rect -592 35941 -558 35975
rect -524 35941 -490 35975
rect -456 35941 -422 35975
rect -388 35941 -354 35975
rect -320 35941 -286 35975
rect -252 35941 -218 35975
rect -184 35941 -153 35975
rect -2969 35906 -153 35941
rect -2969 35872 -2938 35906
rect -2904 35872 -2870 35906
rect -2836 35872 -2802 35906
rect -2768 35872 -2734 35906
rect -2700 35872 -2666 35906
rect -2632 35872 -2598 35906
rect -2564 35872 -2530 35906
rect -2496 35872 -2462 35906
rect -2428 35872 -2394 35906
rect -2360 35872 -2326 35906
rect -2292 35872 -2258 35906
rect -2224 35872 -2190 35906
rect -2156 35872 -2122 35906
rect -2088 35872 -2054 35906
rect -2020 35872 -1986 35906
rect -1952 35872 -1918 35906
rect -1884 35872 -1850 35906
rect -1816 35872 -1782 35906
rect -1748 35872 -1714 35906
rect -1680 35872 -1646 35906
rect -1612 35872 -1578 35906
rect -1544 35872 -1510 35906
rect -1476 35872 -1442 35906
rect -1408 35872 -1374 35906
rect -1340 35872 -1306 35906
rect -1272 35872 -1238 35906
rect -1204 35872 -1170 35906
rect -1136 35872 -1102 35906
rect -1068 35872 -1034 35906
rect -1000 35872 -966 35906
rect -932 35872 -898 35906
rect -864 35872 -830 35906
rect -796 35872 -762 35906
rect -728 35872 -694 35906
rect -660 35872 -626 35906
rect -592 35872 -558 35906
rect -524 35872 -490 35906
rect -456 35872 -422 35906
rect -388 35872 -354 35906
rect -320 35872 -286 35906
rect -252 35872 -218 35906
rect -184 35872 -153 35906
rect -2969 35837 -153 35872
rect -2969 35803 -2938 35837
rect -2904 35803 -2870 35837
rect -2836 35803 -2802 35837
rect -2768 35803 -2734 35837
rect -2700 35803 -2666 35837
rect -2632 35803 -2598 35837
rect -2564 35803 -2530 35837
rect -2496 35803 -2462 35837
rect -2428 35803 -2394 35837
rect -2360 35803 -2326 35837
rect -2292 35803 -2258 35837
rect -2224 35803 -2190 35837
rect -2156 35803 -2122 35837
rect -2088 35803 -2054 35837
rect -2020 35803 -1986 35837
rect -1952 35803 -1918 35837
rect -1884 35803 -1850 35837
rect -1816 35803 -1782 35837
rect -1748 35803 -1714 35837
rect -1680 35803 -1646 35837
rect -1612 35803 -1578 35837
rect -1544 35803 -1510 35837
rect -1476 35803 -1442 35837
rect -1408 35803 -1374 35837
rect -1340 35803 -1306 35837
rect -1272 35803 -1238 35837
rect -1204 35803 -1170 35837
rect -1136 35803 -1102 35837
rect -1068 35803 -1034 35837
rect -1000 35803 -966 35837
rect -932 35803 -898 35837
rect -864 35803 -830 35837
rect -796 35803 -762 35837
rect -728 35803 -694 35837
rect -660 35803 -626 35837
rect -592 35803 -558 35837
rect -524 35803 -490 35837
rect -456 35803 -422 35837
rect -388 35803 -354 35837
rect -320 35803 -286 35837
rect -252 35803 -218 35837
rect -184 35803 -153 35837
rect -2969 35768 -153 35803
rect -2969 35734 -2938 35768
rect -2904 35734 -2870 35768
rect -2836 35734 -2802 35768
rect -2768 35734 -2734 35768
rect -2700 35734 -2666 35768
rect -2632 35734 -2598 35768
rect -2564 35734 -2530 35768
rect -2496 35734 -2462 35768
rect -2428 35734 -2394 35768
rect -2360 35734 -2326 35768
rect -2292 35734 -2258 35768
rect -2224 35734 -2190 35768
rect -2156 35734 -2122 35768
rect -2088 35734 -2054 35768
rect -2020 35734 -1986 35768
rect -1952 35734 -1918 35768
rect -1884 35734 -1850 35768
rect -1816 35734 -1782 35768
rect -1748 35734 -1714 35768
rect -1680 35734 -1646 35768
rect -1612 35734 -1578 35768
rect -1544 35734 -1510 35768
rect -1476 35734 -1442 35768
rect -1408 35734 -1374 35768
rect -1340 35734 -1306 35768
rect -1272 35734 -1238 35768
rect -1204 35734 -1170 35768
rect -1136 35734 -1102 35768
rect -1068 35734 -1034 35768
rect -1000 35734 -966 35768
rect -932 35734 -898 35768
rect -864 35734 -830 35768
rect -796 35734 -762 35768
rect -728 35734 -694 35768
rect -660 35734 -626 35768
rect -592 35734 -558 35768
rect -524 35734 -490 35768
rect -456 35734 -422 35768
rect -388 35734 -354 35768
rect -320 35734 -286 35768
rect -252 35734 -218 35768
rect -184 35734 -153 35768
rect -2969 35699 -153 35734
rect -2969 35665 -2938 35699
rect -2904 35665 -2870 35699
rect -2836 35665 -2802 35699
rect -2768 35665 -2734 35699
rect -2700 35665 -2666 35699
rect -2632 35665 -2598 35699
rect -2564 35665 -2530 35699
rect -2496 35665 -2462 35699
rect -2428 35665 -2394 35699
rect -2360 35665 -2326 35699
rect -2292 35665 -2258 35699
rect -2224 35665 -2190 35699
rect -2156 35665 -2122 35699
rect -2088 35665 -2054 35699
rect -2020 35665 -1986 35699
rect -1952 35665 -1918 35699
rect -1884 35665 -1850 35699
rect -1816 35665 -1782 35699
rect -1748 35665 -1714 35699
rect -1680 35665 -1646 35699
rect -1612 35665 -1578 35699
rect -1544 35665 -1510 35699
rect -1476 35665 -1442 35699
rect -1408 35665 -1374 35699
rect -1340 35665 -1306 35699
rect -1272 35665 -1238 35699
rect -1204 35665 -1170 35699
rect -1136 35665 -1102 35699
rect -1068 35665 -1034 35699
rect -1000 35665 -966 35699
rect -932 35665 -898 35699
rect -864 35665 -830 35699
rect -796 35665 -762 35699
rect -728 35665 -694 35699
rect -660 35665 -626 35699
rect -592 35665 -558 35699
rect -524 35665 -490 35699
rect -456 35665 -422 35699
rect -388 35665 -354 35699
rect -320 35665 -286 35699
rect -252 35665 -218 35699
rect -184 35665 -153 35699
rect -2969 35630 -153 35665
rect -2969 35596 -2938 35630
rect -2904 35596 -2870 35630
rect -2836 35596 -2802 35630
rect -2768 35596 -2734 35630
rect -2700 35596 -2666 35630
rect -2632 35596 -2598 35630
rect -2564 35596 -2530 35630
rect -2496 35596 -2462 35630
rect -2428 35596 -2394 35630
rect -2360 35596 -2326 35630
rect -2292 35596 -2258 35630
rect -2224 35596 -2190 35630
rect -2156 35596 -2122 35630
rect -2088 35596 -2054 35630
rect -2020 35596 -1986 35630
rect -1952 35596 -1918 35630
rect -1884 35596 -1850 35630
rect -1816 35596 -1782 35630
rect -1748 35596 -1714 35630
rect -1680 35596 -1646 35630
rect -1612 35596 -1578 35630
rect -1544 35596 -1510 35630
rect -1476 35596 -1442 35630
rect -1408 35596 -1374 35630
rect -1340 35596 -1306 35630
rect -1272 35596 -1238 35630
rect -1204 35596 -1170 35630
rect -1136 35596 -1102 35630
rect -1068 35596 -1034 35630
rect -1000 35596 -966 35630
rect -932 35596 -898 35630
rect -864 35596 -830 35630
rect -796 35596 -762 35630
rect -728 35596 -694 35630
rect -660 35596 -626 35630
rect -592 35596 -558 35630
rect -524 35596 -490 35630
rect -456 35596 -422 35630
rect -388 35596 -354 35630
rect -320 35596 -286 35630
rect -252 35596 -218 35630
rect -184 35596 -153 35630
rect -2969 35561 -153 35596
rect -2969 35527 -2938 35561
rect -2904 35527 -2870 35561
rect -2836 35527 -2802 35561
rect -2768 35527 -2734 35561
rect -2700 35527 -2666 35561
rect -2632 35527 -2598 35561
rect -2564 35527 -2530 35561
rect -2496 35527 -2462 35561
rect -2428 35527 -2394 35561
rect -2360 35527 -2326 35561
rect -2292 35527 -2258 35561
rect -2224 35527 -2190 35561
rect -2156 35527 -2122 35561
rect -2088 35527 -2054 35561
rect -2020 35527 -1986 35561
rect -1952 35527 -1918 35561
rect -1884 35527 -1850 35561
rect -1816 35527 -1782 35561
rect -1748 35527 -1714 35561
rect -1680 35527 -1646 35561
rect -1612 35527 -1578 35561
rect -1544 35527 -1510 35561
rect -1476 35527 -1442 35561
rect -1408 35527 -1374 35561
rect -1340 35527 -1306 35561
rect -1272 35527 -1238 35561
rect -1204 35527 -1170 35561
rect -1136 35527 -1102 35561
rect -1068 35527 -1034 35561
rect -1000 35527 -966 35561
rect -932 35527 -898 35561
rect -864 35527 -830 35561
rect -796 35527 -762 35561
rect -728 35527 -694 35561
rect -660 35527 -626 35561
rect -592 35527 -558 35561
rect -524 35527 -490 35561
rect -456 35527 -422 35561
rect -388 35527 -354 35561
rect -320 35527 -286 35561
rect -252 35527 -218 35561
rect -184 35527 -153 35561
rect -2969 35492 -153 35527
rect -2969 35458 -2938 35492
rect -2904 35458 -2870 35492
rect -2836 35458 -2802 35492
rect -2768 35458 -2734 35492
rect -2700 35458 -2666 35492
rect -2632 35458 -2598 35492
rect -2564 35458 -2530 35492
rect -2496 35458 -2462 35492
rect -2428 35458 -2394 35492
rect -2360 35458 -2326 35492
rect -2292 35458 -2258 35492
rect -2224 35458 -2190 35492
rect -2156 35458 -2122 35492
rect -2088 35458 -2054 35492
rect -2020 35458 -1986 35492
rect -1952 35458 -1918 35492
rect -1884 35458 -1850 35492
rect -1816 35458 -1782 35492
rect -1748 35458 -1714 35492
rect -1680 35458 -1646 35492
rect -1612 35458 -1578 35492
rect -1544 35458 -1510 35492
rect -1476 35458 -1442 35492
rect -1408 35458 -1374 35492
rect -1340 35458 -1306 35492
rect -1272 35458 -1238 35492
rect -1204 35458 -1170 35492
rect -1136 35458 -1102 35492
rect -1068 35458 -1034 35492
rect -1000 35458 -966 35492
rect -932 35458 -898 35492
rect -864 35458 -830 35492
rect -796 35458 -762 35492
rect -728 35458 -694 35492
rect -660 35458 -626 35492
rect -592 35458 -558 35492
rect -524 35458 -490 35492
rect -456 35458 -422 35492
rect -388 35458 -354 35492
rect -320 35458 -286 35492
rect -252 35458 -218 35492
rect -184 35458 -153 35492
rect -2969 35423 -153 35458
rect -2969 35389 -2938 35423
rect -2904 35389 -2870 35423
rect -2836 35389 -2802 35423
rect -2768 35389 -2734 35423
rect -2700 35389 -2666 35423
rect -2632 35389 -2598 35423
rect -2564 35389 -2530 35423
rect -2496 35389 -2462 35423
rect -2428 35389 -2394 35423
rect -2360 35389 -2326 35423
rect -2292 35389 -2258 35423
rect -2224 35389 -2190 35423
rect -2156 35389 -2122 35423
rect -2088 35389 -2054 35423
rect -2020 35389 -1986 35423
rect -1952 35389 -1918 35423
rect -1884 35389 -1850 35423
rect -1816 35389 -1782 35423
rect -1748 35389 -1714 35423
rect -1680 35389 -1646 35423
rect -1612 35389 -1578 35423
rect -1544 35389 -1510 35423
rect -1476 35389 -1442 35423
rect -1408 35389 -1374 35423
rect -1340 35389 -1306 35423
rect -1272 35389 -1238 35423
rect -1204 35389 -1170 35423
rect -1136 35389 -1102 35423
rect -1068 35389 -1034 35423
rect -1000 35389 -966 35423
rect -932 35389 -898 35423
rect -864 35389 -830 35423
rect -796 35389 -762 35423
rect -728 35389 -694 35423
rect -660 35389 -626 35423
rect -592 35389 -558 35423
rect -524 35389 -490 35423
rect -456 35389 -422 35423
rect -388 35389 -354 35423
rect -320 35389 -286 35423
rect -252 35389 -218 35423
rect -184 35389 -153 35423
rect -2969 35354 -153 35389
rect -2969 35320 -2938 35354
rect -2904 35320 -2870 35354
rect -2836 35320 -2802 35354
rect -2768 35320 -2734 35354
rect -2700 35320 -2666 35354
rect -2632 35320 -2598 35354
rect -2564 35320 -2530 35354
rect -2496 35320 -2462 35354
rect -2428 35320 -2394 35354
rect -2360 35320 -2326 35354
rect -2292 35320 -2258 35354
rect -2224 35320 -2190 35354
rect -2156 35320 -2122 35354
rect -2088 35320 -2054 35354
rect -2020 35320 -1986 35354
rect -1952 35320 -1918 35354
rect -1884 35320 -1850 35354
rect -1816 35320 -1782 35354
rect -1748 35320 -1714 35354
rect -1680 35320 -1646 35354
rect -1612 35320 -1578 35354
rect -1544 35320 -1510 35354
rect -1476 35320 -1442 35354
rect -1408 35320 -1374 35354
rect -1340 35320 -1306 35354
rect -1272 35320 -1238 35354
rect -1204 35320 -1170 35354
rect -1136 35320 -1102 35354
rect -1068 35320 -1034 35354
rect -1000 35320 -966 35354
rect -932 35320 -898 35354
rect -864 35320 -830 35354
rect -796 35320 -762 35354
rect -728 35320 -694 35354
rect -660 35320 -626 35354
rect -592 35320 -558 35354
rect -524 35320 -490 35354
rect -456 35320 -422 35354
rect -388 35320 -354 35354
rect -320 35320 -286 35354
rect -252 35320 -218 35354
rect -184 35320 -153 35354
rect -2969 35285 -153 35320
rect -2969 35251 -2938 35285
rect -2904 35251 -2870 35285
rect -2836 35251 -2802 35285
rect -2768 35251 -2734 35285
rect -2700 35251 -2666 35285
rect -2632 35251 -2598 35285
rect -2564 35251 -2530 35285
rect -2496 35251 -2462 35285
rect -2428 35251 -2394 35285
rect -2360 35251 -2326 35285
rect -2292 35251 -2258 35285
rect -2224 35251 -2190 35285
rect -2156 35251 -2122 35285
rect -2088 35251 -2054 35285
rect -2020 35251 -1986 35285
rect -1952 35251 -1918 35285
rect -1884 35251 -1850 35285
rect -1816 35251 -1782 35285
rect -1748 35251 -1714 35285
rect -1680 35251 -1646 35285
rect -1612 35251 -1578 35285
rect -1544 35251 -1510 35285
rect -1476 35251 -1442 35285
rect -1408 35251 -1374 35285
rect -1340 35251 -1306 35285
rect -1272 35251 -1238 35285
rect -1204 35251 -1170 35285
rect -1136 35251 -1102 35285
rect -1068 35251 -1034 35285
rect -1000 35251 -966 35285
rect -932 35251 -898 35285
rect -864 35251 -830 35285
rect -796 35251 -762 35285
rect -728 35251 -694 35285
rect -660 35251 -626 35285
rect -592 35251 -558 35285
rect -524 35251 -490 35285
rect -456 35251 -422 35285
rect -388 35251 -354 35285
rect -320 35251 -286 35285
rect -252 35251 -218 35285
rect -184 35251 -153 35285
rect -2969 35216 -153 35251
rect -2969 35182 -2938 35216
rect -2904 35182 -2870 35216
rect -2836 35182 -2802 35216
rect -2768 35182 -2734 35216
rect -2700 35182 -2666 35216
rect -2632 35182 -2598 35216
rect -2564 35182 -2530 35216
rect -2496 35182 -2462 35216
rect -2428 35182 -2394 35216
rect -2360 35182 -2326 35216
rect -2292 35182 -2258 35216
rect -2224 35182 -2190 35216
rect -2156 35182 -2122 35216
rect -2088 35182 -2054 35216
rect -2020 35182 -1986 35216
rect -1952 35182 -1918 35216
rect -1884 35182 -1850 35216
rect -1816 35182 -1782 35216
rect -1748 35182 -1714 35216
rect -1680 35182 -1646 35216
rect -1612 35182 -1578 35216
rect -1544 35182 -1510 35216
rect -1476 35182 -1442 35216
rect -1408 35182 -1374 35216
rect -1340 35182 -1306 35216
rect -1272 35182 -1238 35216
rect -1204 35182 -1170 35216
rect -1136 35182 -1102 35216
rect -1068 35182 -1034 35216
rect -1000 35182 -966 35216
rect -932 35182 -898 35216
rect -864 35182 -830 35216
rect -796 35182 -762 35216
rect -728 35182 -694 35216
rect -660 35182 -626 35216
rect -592 35182 -558 35216
rect -524 35182 -490 35216
rect -456 35182 -422 35216
rect -388 35182 -354 35216
rect -320 35182 -286 35216
rect -252 35182 -218 35216
rect -184 35182 -153 35216
rect -2969 35147 -153 35182
rect -2969 35113 -2938 35147
rect -2904 35113 -2870 35147
rect -2836 35113 -2802 35147
rect -2768 35113 -2734 35147
rect -2700 35113 -2666 35147
rect -2632 35113 -2598 35147
rect -2564 35113 -2530 35147
rect -2496 35113 -2462 35147
rect -2428 35113 -2394 35147
rect -2360 35113 -2326 35147
rect -2292 35113 -2258 35147
rect -2224 35113 -2190 35147
rect -2156 35113 -2122 35147
rect -2088 35113 -2054 35147
rect -2020 35113 -1986 35147
rect -1952 35113 -1918 35147
rect -1884 35113 -1850 35147
rect -1816 35113 -1782 35147
rect -1748 35113 -1714 35147
rect -1680 35113 -1646 35147
rect -1612 35113 -1578 35147
rect -1544 35113 -1510 35147
rect -1476 35113 -1442 35147
rect -1408 35113 -1374 35147
rect -1340 35113 -1306 35147
rect -1272 35113 -1238 35147
rect -1204 35113 -1170 35147
rect -1136 35113 -1102 35147
rect -1068 35113 -1034 35147
rect -1000 35113 -966 35147
rect -932 35113 -898 35147
rect -864 35113 -830 35147
rect -796 35113 -762 35147
rect -728 35113 -694 35147
rect -660 35113 -626 35147
rect -592 35113 -558 35147
rect -524 35113 -490 35147
rect -456 35113 -422 35147
rect -388 35113 -354 35147
rect -320 35113 -286 35147
rect -252 35113 -218 35147
rect -184 35113 -153 35147
rect -2969 35078 -153 35113
rect -2969 35044 -2938 35078
rect -2904 35044 -2870 35078
rect -2836 35044 -2802 35078
rect -2768 35044 -2734 35078
rect -2700 35044 -2666 35078
rect -2632 35044 -2598 35078
rect -2564 35044 -2530 35078
rect -2496 35044 -2462 35078
rect -2428 35044 -2394 35078
rect -2360 35044 -2326 35078
rect -2292 35044 -2258 35078
rect -2224 35044 -2190 35078
rect -2156 35044 -2122 35078
rect -2088 35044 -2054 35078
rect -2020 35044 -1986 35078
rect -1952 35044 -1918 35078
rect -1884 35044 -1850 35078
rect -1816 35044 -1782 35078
rect -1748 35044 -1714 35078
rect -1680 35044 -1646 35078
rect -1612 35044 -1578 35078
rect -1544 35044 -1510 35078
rect -1476 35044 -1442 35078
rect -1408 35044 -1374 35078
rect -1340 35044 -1306 35078
rect -1272 35044 -1238 35078
rect -1204 35044 -1170 35078
rect -1136 35044 -1102 35078
rect -1068 35044 -1034 35078
rect -1000 35044 -966 35078
rect -932 35044 -898 35078
rect -864 35044 -830 35078
rect -796 35044 -762 35078
rect -728 35044 -694 35078
rect -660 35044 -626 35078
rect -592 35044 -558 35078
rect -524 35044 -490 35078
rect -456 35044 -422 35078
rect -388 35044 -354 35078
rect -320 35044 -286 35078
rect -252 35044 -218 35078
rect -184 35044 -153 35078
rect -2969 35020 -153 35044
rect -2966 17927 -266 17951
rect -2966 10413 -2959 17927
rect -273 10413 -266 17927
rect 18281 14481 29669 14484
rect 18281 14447 18349 14481
rect 18383 14447 18418 14481
rect 18452 14447 18487 14481
rect 18521 14447 18556 14481
rect 18590 14447 18625 14481
rect 18659 14447 18694 14481
rect 18728 14447 18763 14481
rect 18797 14447 18832 14481
rect 18866 14447 18901 14481
rect 18935 14447 18970 14481
rect 19004 14447 19039 14481
rect 19073 14447 19108 14481
rect 19142 14447 19177 14481
rect 19211 14447 19246 14481
rect 19280 14447 19315 14481
rect 19349 14447 19384 14481
rect 19418 14447 19453 14481
rect 19487 14447 19522 14481
rect 19556 14447 19591 14481
rect 19625 14447 19660 14481
rect 19694 14447 19729 14481
rect 19763 14447 19798 14481
rect 19832 14447 19867 14481
rect 19901 14447 19936 14481
rect 19970 14447 20005 14481
rect 20039 14447 20074 14481
rect 20108 14447 20143 14481
rect 20177 14447 20212 14481
rect 20246 14447 20281 14481
rect 20315 14447 20350 14481
rect 20384 14447 20419 14481
rect 20453 14447 20488 14481
rect 20522 14447 20557 14481
rect 20591 14447 20626 14481
rect 20660 14447 20695 14481
rect 20729 14447 20764 14481
rect 20798 14447 20833 14481
rect 20867 14447 20902 14481
rect 20936 14447 20971 14481
rect 21005 14447 21040 14481
rect 21074 14447 21109 14481
rect 21143 14447 21178 14481
rect 21212 14447 21247 14481
rect 21281 14447 21315 14481
rect 21349 14447 21383 14481
rect 21417 14447 21451 14481
rect 21485 14447 21519 14481
rect 21553 14447 21587 14481
rect 21621 14447 21655 14481
rect 21689 14447 21723 14481
rect 21757 14447 21791 14481
rect 21825 14447 21859 14481
rect 21893 14447 21927 14481
rect 21961 14447 21995 14481
rect 22029 14447 22063 14481
rect 22097 14447 22131 14481
rect 22165 14447 22199 14481
rect 22233 14447 22267 14481
rect 22301 14447 22335 14481
rect 22369 14447 22403 14481
rect 22437 14447 22471 14481
rect 22505 14447 22539 14481
rect 22573 14447 22607 14481
rect 22641 14447 22675 14481
rect 22709 14447 22743 14481
rect 22777 14447 22811 14481
rect 22845 14447 22879 14481
rect 22913 14447 22947 14481
rect 22981 14447 23015 14481
rect 23049 14447 23083 14481
rect 23117 14447 23151 14481
rect 23185 14447 23219 14481
rect 23253 14447 23287 14481
rect 23321 14447 23355 14481
rect 23389 14447 23423 14481
rect 23457 14447 23491 14481
rect 23525 14447 23559 14481
rect 23593 14447 23627 14481
rect 23661 14447 23695 14481
rect 23729 14447 23763 14481
rect 23797 14447 23831 14481
rect 23865 14447 23899 14481
rect 23933 14447 23967 14481
rect 24001 14447 24035 14481
rect 24069 14447 24103 14481
rect 24137 14447 24171 14481
rect 24205 14447 24239 14481
rect 24273 14447 24307 14481
rect 24341 14447 24375 14481
rect 24409 14447 24443 14481
rect 24477 14447 24511 14481
rect 24545 14447 24579 14481
rect 24613 14447 24647 14481
rect 24681 14447 24715 14481
rect 24749 14447 24783 14481
rect 24817 14447 24851 14481
rect 24885 14447 24919 14481
rect 24953 14447 24987 14481
rect 25021 14447 25055 14481
rect 25089 14447 25123 14481
rect 25157 14447 25191 14481
rect 25225 14447 25259 14481
rect 25293 14447 25327 14481
rect 25361 14447 25395 14481
rect 25429 14447 25463 14481
rect 25497 14447 25531 14481
rect 25565 14447 25599 14481
rect 25633 14447 25667 14481
rect 25701 14447 25735 14481
rect 25769 14447 25803 14481
rect 25837 14447 25871 14481
rect 25905 14447 25939 14481
rect 25973 14447 26007 14481
rect 26041 14447 26075 14481
rect 26109 14447 26143 14481
rect 26177 14447 26211 14481
rect 26245 14447 26279 14481
rect 26313 14447 26347 14481
rect 26381 14447 26415 14481
rect 26449 14447 26483 14481
rect 26517 14447 26551 14481
rect 26585 14447 26619 14481
rect 26653 14447 26687 14481
rect 26721 14447 26755 14481
rect 26789 14447 26823 14481
rect 26857 14447 26891 14481
rect 26925 14447 26959 14481
rect 26993 14447 27027 14481
rect 27061 14447 27095 14481
rect 27129 14447 27163 14481
rect 27197 14447 27231 14481
rect 27265 14447 27299 14481
rect 27333 14447 27367 14481
rect 27401 14447 27435 14481
rect 27469 14447 27503 14481
rect 27537 14447 27571 14481
rect 27605 14447 27639 14481
rect 27673 14447 27707 14481
rect 27741 14447 27775 14481
rect 27809 14447 27843 14481
rect 27877 14447 27911 14481
rect 27945 14447 27979 14481
rect 28013 14447 28047 14481
rect 28081 14447 28115 14481
rect 28149 14447 28183 14481
rect 28217 14447 28251 14481
rect 28285 14447 28319 14481
rect 28353 14447 28387 14481
rect 28421 14447 28455 14481
rect 28489 14447 28523 14481
rect 28557 14447 28591 14481
rect 28625 14447 28659 14481
rect 28693 14447 28727 14481
rect 28761 14447 28795 14481
rect 28829 14447 28863 14481
rect 28897 14447 28931 14481
rect 28965 14447 28999 14481
rect 29033 14447 29067 14481
rect 29101 14447 29135 14481
rect 29169 14447 29203 14481
rect 29237 14447 29271 14481
rect 29305 14447 29339 14481
rect 29373 14447 29407 14481
rect 29441 14447 29475 14481
rect 29509 14447 29543 14481
rect 29577 14447 29611 14481
rect 29645 14447 29669 14481
rect 18281 14415 29669 14447
rect 18281 14381 18284 14415
rect 18318 14409 29669 14415
rect 18318 14381 18356 14409
rect 18281 14375 18356 14381
rect 18390 14375 18425 14409
rect 18459 14375 18494 14409
rect 18528 14375 18563 14409
rect 18597 14375 18632 14409
rect 18666 14375 18701 14409
rect 18735 14375 18770 14409
rect 18804 14375 18839 14409
rect 18873 14375 18908 14409
rect 18942 14375 18977 14409
rect 19011 14375 19046 14409
rect 19080 14375 19115 14409
rect 19149 14375 19184 14409
rect 19218 14375 19253 14409
rect 19287 14375 19322 14409
rect 19356 14375 19391 14409
rect 19425 14375 19460 14409
rect 19494 14375 19529 14409
rect 19563 14375 19598 14409
rect 19632 14375 19667 14409
rect 19701 14375 19736 14409
rect 19770 14375 19805 14409
rect 19839 14375 19874 14409
rect 19908 14375 19943 14409
rect 19977 14375 20012 14409
rect 20046 14375 20081 14409
rect 20115 14375 20150 14409
rect 20184 14375 20219 14409
rect 20253 14375 20288 14409
rect 20322 14375 20357 14409
rect 20391 14375 20426 14409
rect 20460 14375 20495 14409
rect 20529 14375 20564 14409
rect 20598 14375 20633 14409
rect 20667 14375 20702 14409
rect 20736 14375 20771 14409
rect 20805 14375 20839 14409
rect 20873 14375 20907 14409
rect 20941 14375 20975 14409
rect 21009 14375 21043 14409
rect 21077 14375 21111 14409
rect 21145 14375 21179 14409
rect 21213 14375 21247 14409
rect 21281 14375 21315 14409
rect 21349 14375 21383 14409
rect 21417 14375 21451 14409
rect 21485 14375 21519 14409
rect 21553 14375 21587 14409
rect 21621 14375 21655 14409
rect 21689 14375 21723 14409
rect 21757 14375 21791 14409
rect 21825 14375 21859 14409
rect 21893 14375 21927 14409
rect 21961 14375 21995 14409
rect 22029 14375 22063 14409
rect 22097 14375 22131 14409
rect 22165 14375 22199 14409
rect 22233 14375 22267 14409
rect 22301 14375 22335 14409
rect 22369 14375 22403 14409
rect 22437 14375 22471 14409
rect 22505 14375 22539 14409
rect 22573 14375 22607 14409
rect 22641 14375 22675 14409
rect 22709 14375 22743 14409
rect 22777 14375 22811 14409
rect 22845 14375 22879 14409
rect 22913 14375 22947 14409
rect 22981 14375 23015 14409
rect 23049 14375 23083 14409
rect 23117 14375 23151 14409
rect 23185 14375 23219 14409
rect 23253 14375 23287 14409
rect 23321 14375 23355 14409
rect 23389 14375 23423 14409
rect 23457 14375 23491 14409
rect 23525 14375 23559 14409
rect 23593 14375 23627 14409
rect 23661 14375 23695 14409
rect 23729 14375 23763 14409
rect 23797 14375 23831 14409
rect 23865 14375 23899 14409
rect 23933 14375 23967 14409
rect 24001 14375 24035 14409
rect 24069 14375 24103 14409
rect 24137 14375 24171 14409
rect 24205 14375 24239 14409
rect 24273 14375 24307 14409
rect 24341 14375 24375 14409
rect 24409 14375 24443 14409
rect 24477 14375 24511 14409
rect 24545 14375 24579 14409
rect 24613 14375 24647 14409
rect 24681 14375 24715 14409
rect 24749 14375 24783 14409
rect 24817 14375 24851 14409
rect 24885 14375 24919 14409
rect 24953 14375 24987 14409
rect 25021 14375 25055 14409
rect 25089 14375 25123 14409
rect 25157 14375 25191 14409
rect 25225 14375 25259 14409
rect 25293 14375 25327 14409
rect 25361 14375 25395 14409
rect 25429 14375 25463 14409
rect 25497 14375 25531 14409
rect 25565 14375 25599 14409
rect 25633 14375 25667 14409
rect 25701 14375 25735 14409
rect 25769 14375 25803 14409
rect 25837 14375 25871 14409
rect 25905 14375 25939 14409
rect 25973 14375 26007 14409
rect 26041 14375 26075 14409
rect 26109 14375 26143 14409
rect 26177 14375 26211 14409
rect 26245 14375 26279 14409
rect 26313 14375 26347 14409
rect 26381 14375 26415 14409
rect 26449 14375 26483 14409
rect 26517 14375 26551 14409
rect 26585 14375 26619 14409
rect 26653 14375 26687 14409
rect 26721 14375 26755 14409
rect 26789 14375 26823 14409
rect 26857 14375 26891 14409
rect 26925 14375 26959 14409
rect 26993 14375 27027 14409
rect 27061 14375 27095 14409
rect 27129 14375 27163 14409
rect 27197 14375 27231 14409
rect 27265 14375 27299 14409
rect 27333 14375 27367 14409
rect 27401 14375 27435 14409
rect 27469 14375 27503 14409
rect 27537 14375 27571 14409
rect 27605 14375 27639 14409
rect 27673 14375 27707 14409
rect 27741 14375 27775 14409
rect 27809 14375 27843 14409
rect 27877 14375 27911 14409
rect 27945 14375 27979 14409
rect 28013 14375 28047 14409
rect 28081 14375 28115 14409
rect 28149 14375 28183 14409
rect 28217 14375 28251 14409
rect 28285 14375 28319 14409
rect 28353 14375 28387 14409
rect 28421 14375 28455 14409
rect 28489 14375 28523 14409
rect 28557 14375 28591 14409
rect 28625 14375 28659 14409
rect 28693 14375 28727 14409
rect 28761 14375 28795 14409
rect 28829 14375 28863 14409
rect 28897 14375 28931 14409
rect 28965 14375 28999 14409
rect 29033 14375 29067 14409
rect 29101 14375 29135 14409
rect 29169 14375 29203 14409
rect 29237 14375 29271 14409
rect 29305 14375 29339 14409
rect 29373 14375 29407 14409
rect 29441 14375 29475 14409
rect 29509 14375 29543 14409
rect 29577 14375 29611 14409
rect 29645 14375 29669 14409
rect 18281 14345 29669 14375
rect 18281 14311 18284 14345
rect 18318 14340 29669 14345
rect 18318 14311 18356 14340
rect 18281 14306 18356 14311
rect 18390 14337 29669 14340
rect 18390 14306 18428 14337
rect 18281 14303 18428 14306
rect 18462 14303 18497 14337
rect 18531 14303 18566 14337
rect 18600 14303 18635 14337
rect 18669 14303 18704 14337
rect 18738 14303 18773 14337
rect 18807 14303 18842 14337
rect 18876 14303 18911 14337
rect 18945 14303 18980 14337
rect 19014 14303 19049 14337
rect 19083 14303 19118 14337
rect 19152 14303 19187 14337
rect 19221 14303 19256 14337
rect 19290 14303 19325 14337
rect 19359 14303 19394 14337
rect 19428 14303 19463 14337
rect 19497 14303 19532 14337
rect 19566 14303 19601 14337
rect 19635 14303 19670 14337
rect 19704 14303 19739 14337
rect 19773 14303 19808 14337
rect 19842 14303 19877 14337
rect 19911 14303 19946 14337
rect 19980 14303 20015 14337
rect 20049 14303 20084 14337
rect 20118 14303 20153 14337
rect 20187 14303 20222 14337
rect 20256 14303 20291 14337
rect 20325 14303 20360 14337
rect 20394 14303 20429 14337
rect 20463 14303 20498 14337
rect 20532 14303 20567 14337
rect 20601 14303 20635 14337
rect 20669 14303 20703 14337
rect 20737 14303 20771 14337
rect 20805 14303 20839 14337
rect 20873 14303 20907 14337
rect 20941 14303 20975 14337
rect 21009 14303 21043 14337
rect 21077 14303 21111 14337
rect 21145 14303 21179 14337
rect 21213 14303 21247 14337
rect 21281 14303 21315 14337
rect 21349 14303 21383 14337
rect 21417 14303 21451 14337
rect 21485 14303 21519 14337
rect 21553 14303 21587 14337
rect 21621 14303 21655 14337
rect 21689 14303 21723 14337
rect 21757 14303 21791 14337
rect 21825 14303 21859 14337
rect 21893 14303 21927 14337
rect 21961 14303 21995 14337
rect 22029 14303 22063 14337
rect 22097 14303 22131 14337
rect 22165 14303 22199 14337
rect 22233 14303 22267 14337
rect 22301 14303 22335 14337
rect 22369 14303 22403 14337
rect 22437 14303 22471 14337
rect 22505 14303 22539 14337
rect 22573 14303 22607 14337
rect 22641 14303 22675 14337
rect 22709 14303 22743 14337
rect 22777 14303 22811 14337
rect 22845 14303 22879 14337
rect 22913 14303 22947 14337
rect 22981 14303 23015 14337
rect 23049 14303 23083 14337
rect 23117 14303 23151 14337
rect 23185 14303 23219 14337
rect 23253 14303 23287 14337
rect 23321 14303 23355 14337
rect 23389 14303 23423 14337
rect 23457 14303 23491 14337
rect 23525 14303 23559 14337
rect 23593 14303 23627 14337
rect 23661 14303 23695 14337
rect 23729 14303 23763 14337
rect 23797 14303 23831 14337
rect 23865 14303 23899 14337
rect 23933 14303 23967 14337
rect 24001 14303 24035 14337
rect 24069 14303 24103 14337
rect 24137 14303 24171 14337
rect 24205 14303 24239 14337
rect 24273 14303 24307 14337
rect 24341 14303 24375 14337
rect 24409 14303 24443 14337
rect 24477 14303 24511 14337
rect 24545 14303 24579 14337
rect 24613 14303 24647 14337
rect 24681 14303 24715 14337
rect 24749 14303 24783 14337
rect 24817 14303 24851 14337
rect 24885 14303 24919 14337
rect 24953 14303 24987 14337
rect 25021 14303 25055 14337
rect 25089 14303 25123 14337
rect 25157 14303 25191 14337
rect 25225 14303 25259 14337
rect 25293 14303 25327 14337
rect 25361 14303 25395 14337
rect 25429 14303 25463 14337
rect 25497 14303 25531 14337
rect 25565 14303 25599 14337
rect 25633 14303 25667 14337
rect 25701 14303 25735 14337
rect 25769 14303 25803 14337
rect 25837 14303 25871 14337
rect 25905 14303 25939 14337
rect 25973 14303 26007 14337
rect 26041 14303 26075 14337
rect 26109 14303 26143 14337
rect 26177 14303 26211 14337
rect 26245 14303 26279 14337
rect 26313 14303 26347 14337
rect 26381 14303 26415 14337
rect 26449 14303 26483 14337
rect 26517 14303 26551 14337
rect 26585 14303 26619 14337
rect 26653 14303 26687 14337
rect 26721 14303 26755 14337
rect 26789 14303 26823 14337
rect 26857 14303 26891 14337
rect 26925 14303 26959 14337
rect 26993 14303 27027 14337
rect 27061 14303 27095 14337
rect 27129 14303 27163 14337
rect 27197 14303 27231 14337
rect 27265 14303 27299 14337
rect 27333 14303 27367 14337
rect 27401 14303 27435 14337
rect 27469 14303 27503 14337
rect 27537 14303 27571 14337
rect 27605 14303 27639 14337
rect 27673 14303 27707 14337
rect 27741 14303 27775 14337
rect 27809 14303 27843 14337
rect 27877 14303 27911 14337
rect 27945 14303 27979 14337
rect 28013 14303 28047 14337
rect 28081 14303 28115 14337
rect 28149 14303 28183 14337
rect 28217 14303 28251 14337
rect 28285 14303 28319 14337
rect 28353 14303 28387 14337
rect 28421 14303 28455 14337
rect 28489 14303 28523 14337
rect 28557 14303 28591 14337
rect 28625 14303 28659 14337
rect 28693 14303 28727 14337
rect 28761 14303 28795 14337
rect 28829 14303 28863 14337
rect 28897 14303 28931 14337
rect 28965 14303 28999 14337
rect 29033 14303 29067 14337
rect 29101 14303 29135 14337
rect 29169 14303 29203 14337
rect 29237 14303 29271 14337
rect 29305 14303 29339 14337
rect 29373 14303 29407 14337
rect 29441 14303 29475 14337
rect 29509 14303 29543 14337
rect 29577 14303 29611 14337
rect 29645 14303 29669 14337
rect 18281 14275 29669 14303
rect 18281 14241 18284 14275
rect 18318 14271 29669 14275
rect 18318 14241 18356 14271
rect 18281 14237 18356 14241
rect 18390 14268 29669 14271
rect 18390 14237 18428 14268
rect 18281 14234 18428 14237
rect 18462 14265 29669 14268
rect 18462 14234 18500 14265
rect 18281 14231 18500 14234
rect 18534 14231 18569 14265
rect 18603 14231 18638 14265
rect 18672 14231 18707 14265
rect 18741 14231 18776 14265
rect 18810 14231 18845 14265
rect 18879 14231 18914 14265
rect 18948 14231 18983 14265
rect 19017 14231 19052 14265
rect 19086 14231 19121 14265
rect 19155 14231 19190 14265
rect 19224 14231 19259 14265
rect 19293 14231 19328 14265
rect 19362 14231 19397 14265
rect 19431 14231 19466 14265
rect 19500 14231 19535 14265
rect 19569 14231 19604 14265
rect 19638 14231 19673 14265
rect 19707 14231 19742 14265
rect 19776 14231 19811 14265
rect 19845 14231 19880 14265
rect 19914 14231 19949 14265
rect 19983 14231 20018 14265
rect 20052 14231 20087 14265
rect 20121 14231 20156 14265
rect 20190 14231 20225 14265
rect 20259 14231 20294 14265
rect 20328 14231 20363 14265
rect 20397 14231 20431 14265
rect 20465 14231 20499 14265
rect 20533 14231 20567 14265
rect 20601 14231 20635 14265
rect 20669 14231 20703 14265
rect 20737 14231 20771 14265
rect 20805 14231 20839 14265
rect 20873 14231 20907 14265
rect 20941 14231 20975 14265
rect 21009 14231 21043 14265
rect 21077 14231 21111 14265
rect 21145 14231 21179 14265
rect 21213 14231 21247 14265
rect 21281 14231 21315 14265
rect 21349 14231 21383 14265
rect 21417 14231 21451 14265
rect 21485 14231 21519 14265
rect 21553 14231 21587 14265
rect 21621 14231 21655 14265
rect 21689 14231 21723 14265
rect 21757 14231 21791 14265
rect 21825 14231 21859 14265
rect 21893 14231 21927 14265
rect 21961 14231 21995 14265
rect 22029 14231 22063 14265
rect 22097 14231 22131 14265
rect 22165 14231 22199 14265
rect 22233 14231 22267 14265
rect 22301 14231 22335 14265
rect 22369 14231 22403 14265
rect 22437 14231 22471 14265
rect 22505 14231 22539 14265
rect 22573 14231 22607 14265
rect 22641 14231 22675 14265
rect 22709 14231 22743 14265
rect 22777 14231 22811 14265
rect 22845 14231 22879 14265
rect 22913 14231 22947 14265
rect 22981 14231 23015 14265
rect 23049 14231 23083 14265
rect 23117 14231 23151 14265
rect 23185 14231 23219 14265
rect 23253 14231 23287 14265
rect 23321 14231 23355 14265
rect 23389 14231 23423 14265
rect 23457 14231 23491 14265
rect 23525 14231 23559 14265
rect 23593 14231 23627 14265
rect 23661 14231 23695 14265
rect 23729 14231 23763 14265
rect 23797 14231 23831 14265
rect 23865 14231 23899 14265
rect 23933 14231 23967 14265
rect 24001 14231 24035 14265
rect 24069 14231 24103 14265
rect 24137 14231 24171 14265
rect 24205 14231 24239 14265
rect 24273 14231 24307 14265
rect 24341 14231 24375 14265
rect 24409 14231 24443 14265
rect 24477 14231 24511 14265
rect 24545 14231 24579 14265
rect 24613 14231 24647 14265
rect 24681 14231 24715 14265
rect 24749 14231 24783 14265
rect 24817 14231 24851 14265
rect 24885 14231 24919 14265
rect 24953 14231 24987 14265
rect 25021 14231 25055 14265
rect 25089 14231 25123 14265
rect 25157 14231 25191 14265
rect 25225 14231 25259 14265
rect 25293 14231 25327 14265
rect 25361 14231 25395 14265
rect 25429 14231 25463 14265
rect 25497 14231 25531 14265
rect 25565 14231 25599 14265
rect 25633 14231 25667 14265
rect 25701 14231 25735 14265
rect 25769 14231 25803 14265
rect 25837 14231 25871 14265
rect 25905 14231 25939 14265
rect 25973 14231 26007 14265
rect 26041 14231 26075 14265
rect 26109 14231 26143 14265
rect 26177 14231 26211 14265
rect 26245 14231 26279 14265
rect 26313 14231 26347 14265
rect 26381 14231 26415 14265
rect 26449 14231 26483 14265
rect 26517 14231 26551 14265
rect 26585 14231 26619 14265
rect 26653 14231 26687 14265
rect 26721 14231 26755 14265
rect 26789 14231 26823 14265
rect 26857 14231 26891 14265
rect 26925 14231 26959 14265
rect 26993 14231 27027 14265
rect 27061 14231 27095 14265
rect 27129 14231 27163 14265
rect 27197 14231 27231 14265
rect 27265 14231 27299 14265
rect 27333 14231 27367 14265
rect 27401 14231 27435 14265
rect 27469 14231 27503 14265
rect 27537 14231 27571 14265
rect 27605 14231 27639 14265
rect 27673 14231 27707 14265
rect 27741 14231 27775 14265
rect 27809 14231 27843 14265
rect 27877 14231 27911 14265
rect 27945 14231 27979 14265
rect 28013 14231 28047 14265
rect 28081 14231 28115 14265
rect 28149 14231 28183 14265
rect 28217 14231 28251 14265
rect 28285 14231 28319 14265
rect 28353 14231 28387 14265
rect 28421 14231 28455 14265
rect 28489 14231 28523 14265
rect 28557 14231 28591 14265
rect 28625 14231 28659 14265
rect 28693 14231 28727 14265
rect 28761 14231 28795 14265
rect 28829 14231 28863 14265
rect 28897 14231 28931 14265
rect 28965 14231 28999 14265
rect 29033 14231 29067 14265
rect 29101 14231 29135 14265
rect 29169 14231 29203 14265
rect 29237 14231 29271 14265
rect 29305 14231 29339 14265
rect 29373 14231 29407 14265
rect 29441 14231 29475 14265
rect 29509 14231 29543 14265
rect 29577 14231 29611 14265
rect 29645 14231 29669 14265
rect 18281 14208 29669 14231
rect 15831 14205 29669 14208
rect 15831 14171 15855 14205
rect 15889 14171 15925 14205
rect 15959 14171 15995 14205
rect 16029 14171 16065 14205
rect 16099 14171 16135 14205
rect 16169 14171 16205 14205
rect 16239 14171 16275 14205
rect 16309 14171 16345 14205
rect 16379 14171 16415 14205
rect 16449 14171 16485 14205
rect 16519 14171 16555 14205
rect 16589 14171 16625 14205
rect 16659 14171 16695 14205
rect 16729 14171 16765 14205
rect 16799 14171 16835 14205
rect 16869 14171 16904 14205
rect 16938 14171 16973 14205
rect 17007 14171 17042 14205
rect 17076 14171 17111 14205
rect 17145 14171 17180 14205
rect 17214 14171 17249 14205
rect 17283 14171 17318 14205
rect 17352 14171 17387 14205
rect 17421 14171 17456 14205
rect 17490 14171 17525 14205
rect 17559 14171 17594 14205
rect 17628 14171 17663 14205
rect 17697 14171 17732 14205
rect 17766 14171 17801 14205
rect 17835 14171 17870 14205
rect 17904 14171 17939 14205
rect 17973 14171 18008 14205
rect 18042 14171 18077 14205
rect 18111 14171 18146 14205
rect 18180 14171 18215 14205
rect 18249 14171 18284 14205
rect 18318 14202 29669 14205
rect 18318 14171 18356 14202
rect 15831 14168 18356 14171
rect 18390 14199 29669 14202
rect 18390 14168 18428 14199
rect 15831 14165 18428 14168
rect 18462 14196 29669 14199
rect 18462 14165 18500 14196
rect 15831 14162 18500 14165
rect 18534 14193 29669 14196
rect 18534 14162 18572 14193
rect 15831 14159 18572 14162
rect 18606 14159 18641 14193
rect 18675 14159 18710 14193
rect 18744 14159 18779 14193
rect 18813 14159 18848 14193
rect 18882 14159 18917 14193
rect 18951 14159 18986 14193
rect 19020 14159 19055 14193
rect 19089 14159 19124 14193
rect 19158 14159 19193 14193
rect 19227 14159 19262 14193
rect 19296 14159 19331 14193
rect 19365 14159 19400 14193
rect 19434 14159 19469 14193
rect 19503 14159 19538 14193
rect 19572 14159 19607 14193
rect 19641 14159 19676 14193
rect 19710 14159 19745 14193
rect 19779 14159 19814 14193
rect 19848 14159 19883 14193
rect 19917 14159 19952 14193
rect 19986 14159 20021 14193
rect 20055 14159 20090 14193
rect 20124 14159 20159 14193
rect 20193 14159 20227 14193
rect 20261 14159 20295 14193
rect 20329 14159 20363 14193
rect 20397 14159 20431 14193
rect 20465 14159 20499 14193
rect 20533 14159 20567 14193
rect 20601 14159 20635 14193
rect 20669 14159 20703 14193
rect 20737 14159 20771 14193
rect 20805 14159 20839 14193
rect 20873 14159 20907 14193
rect 20941 14159 20975 14193
rect 21009 14159 21043 14193
rect 21077 14159 21111 14193
rect 21145 14159 21179 14193
rect 21213 14159 21247 14193
rect 21281 14159 21315 14193
rect 21349 14159 21383 14193
rect 21417 14159 21451 14193
rect 21485 14159 21519 14193
rect 21553 14159 21587 14193
rect 21621 14159 21655 14193
rect 21689 14159 21723 14193
rect 21757 14159 21791 14193
rect 21825 14159 21859 14193
rect 21893 14159 21927 14193
rect 21961 14159 21995 14193
rect 22029 14159 22063 14193
rect 22097 14159 22131 14193
rect 22165 14159 22199 14193
rect 22233 14159 22267 14193
rect 22301 14159 22335 14193
rect 22369 14159 22403 14193
rect 22437 14159 22471 14193
rect 22505 14159 22539 14193
rect 22573 14159 22607 14193
rect 22641 14159 22675 14193
rect 22709 14159 22743 14193
rect 22777 14159 22811 14193
rect 22845 14159 22879 14193
rect 22913 14159 22947 14193
rect 22981 14159 23015 14193
rect 23049 14159 23083 14193
rect 23117 14159 23151 14193
rect 23185 14159 23219 14193
rect 23253 14159 23287 14193
rect 23321 14159 23355 14193
rect 23389 14159 23423 14193
rect 23457 14159 23491 14193
rect 23525 14159 23559 14193
rect 23593 14159 23627 14193
rect 23661 14159 23695 14193
rect 23729 14159 23763 14193
rect 23797 14159 23831 14193
rect 23865 14159 23899 14193
rect 23933 14159 23967 14193
rect 24001 14159 24035 14193
rect 24069 14159 24103 14193
rect 24137 14159 24171 14193
rect 24205 14159 24239 14193
rect 24273 14159 24307 14193
rect 24341 14159 24375 14193
rect 24409 14159 24443 14193
rect 24477 14159 24511 14193
rect 24545 14159 24579 14193
rect 24613 14159 24647 14193
rect 24681 14159 24715 14193
rect 24749 14159 24783 14193
rect 24817 14159 24851 14193
rect 24885 14159 24919 14193
rect 24953 14159 24987 14193
rect 25021 14159 25055 14193
rect 25089 14159 25123 14193
rect 25157 14159 25191 14193
rect 25225 14159 25259 14193
rect 25293 14159 25327 14193
rect 25361 14159 25395 14193
rect 25429 14159 25463 14193
rect 25497 14159 25531 14193
rect 25565 14159 25599 14193
rect 25633 14159 25667 14193
rect 25701 14159 25735 14193
rect 25769 14159 25803 14193
rect 25837 14159 25871 14193
rect 25905 14159 25939 14193
rect 25973 14159 26007 14193
rect 26041 14159 26075 14193
rect 26109 14159 26143 14193
rect 26177 14159 26211 14193
rect 26245 14159 26279 14193
rect 26313 14159 26347 14193
rect 26381 14159 26415 14193
rect 26449 14159 26483 14193
rect 26517 14159 26551 14193
rect 26585 14159 26619 14193
rect 26653 14159 26687 14193
rect 26721 14159 26755 14193
rect 26789 14159 26823 14193
rect 26857 14159 26891 14193
rect 26925 14159 26959 14193
rect 26993 14159 27027 14193
rect 27061 14159 27095 14193
rect 27129 14159 27163 14193
rect 27197 14159 27231 14193
rect 27265 14159 27299 14193
rect 27333 14159 27367 14193
rect 27401 14159 27435 14193
rect 27469 14159 27503 14193
rect 27537 14159 27571 14193
rect 27605 14159 27639 14193
rect 27673 14159 27707 14193
rect 27741 14159 27775 14193
rect 27809 14159 27843 14193
rect 27877 14159 27911 14193
rect 27945 14159 27979 14193
rect 28013 14159 28047 14193
rect 28081 14159 28115 14193
rect 28149 14159 28183 14193
rect 28217 14159 28251 14193
rect 28285 14159 28319 14193
rect 28353 14159 28387 14193
rect 28421 14159 28455 14193
rect 28489 14159 28523 14193
rect 28557 14159 28591 14193
rect 28625 14159 28659 14193
rect 28693 14159 28727 14193
rect 28761 14159 28795 14193
rect 28829 14159 28863 14193
rect 28897 14159 28931 14193
rect 28965 14159 28999 14193
rect 29033 14159 29067 14193
rect 29101 14159 29135 14193
rect 29169 14159 29203 14193
rect 29237 14159 29271 14193
rect 29305 14159 29339 14193
rect 29373 14159 29407 14193
rect 29441 14159 29475 14193
rect 29509 14159 29543 14193
rect 29577 14159 29611 14193
rect 29645 14159 29669 14193
rect 15831 14133 29669 14159
rect 15831 14099 15855 14133
rect 15889 14099 15925 14133
rect 15959 14099 15995 14133
rect 16029 14099 16065 14133
rect 16099 14099 16135 14133
rect 16169 14099 16205 14133
rect 16239 14099 16275 14133
rect 16309 14099 16345 14133
rect 16379 14099 16415 14133
rect 16449 14099 16485 14133
rect 16519 14099 16555 14133
rect 16589 14099 16625 14133
rect 16659 14099 16695 14133
rect 16729 14099 16765 14133
rect 16799 14099 16835 14133
rect 16869 14099 16905 14133
rect 16939 14099 16975 14133
rect 17009 14099 17045 14133
rect 17079 14099 17114 14133
rect 17148 14099 17183 14133
rect 17217 14099 17252 14133
rect 17286 14099 17321 14133
rect 17355 14099 17390 14133
rect 17424 14099 17459 14133
rect 17493 14099 17528 14133
rect 17562 14099 17597 14133
rect 17631 14099 17666 14133
rect 17700 14099 17735 14133
rect 17769 14099 17804 14133
rect 17838 14099 17873 14133
rect 17907 14099 17942 14133
rect 17976 14099 18011 14133
rect 18045 14099 18080 14133
rect 18114 14099 18149 14133
rect 18183 14099 18218 14133
rect 18252 14099 18287 14133
rect 18321 14099 18356 14133
rect 18390 14130 29669 14133
rect 18390 14099 18428 14130
rect 15831 14096 18428 14099
rect 18462 14127 29669 14130
rect 18462 14096 18500 14127
rect 15831 14093 18500 14096
rect 18534 14124 29669 14127
rect 18534 14093 18572 14124
rect 15831 14090 18572 14093
rect 18606 14121 29669 14124
rect 18606 14090 18644 14121
rect 15831 14087 18644 14090
rect 18678 14087 18713 14121
rect 18747 14087 18782 14121
rect 18816 14087 18851 14121
rect 18885 14087 18920 14121
rect 18954 14087 18989 14121
rect 19023 14087 19058 14121
rect 19092 14087 19127 14121
rect 19161 14087 19196 14121
rect 19230 14087 19265 14121
rect 19299 14087 19334 14121
rect 19368 14087 19403 14121
rect 19437 14087 19472 14121
rect 19506 14087 19541 14121
rect 19575 14087 19610 14121
rect 19644 14087 19679 14121
rect 19713 14087 19748 14121
rect 19782 14087 19817 14121
rect 19851 14087 19886 14121
rect 19920 14087 19955 14121
rect 19989 14087 20023 14121
rect 20057 14087 20091 14121
rect 20125 14087 20159 14121
rect 20193 14087 20227 14121
rect 20261 14087 20295 14121
rect 20329 14087 20363 14121
rect 20397 14087 20431 14121
rect 20465 14087 20499 14121
rect 20533 14087 20567 14121
rect 20601 14087 20635 14121
rect 20669 14087 20703 14121
rect 20737 14087 20771 14121
rect 20805 14087 20839 14121
rect 20873 14087 20907 14121
rect 20941 14087 20975 14121
rect 21009 14087 21043 14121
rect 21077 14087 21111 14121
rect 21145 14087 21179 14121
rect 21213 14087 21247 14121
rect 21281 14087 21315 14121
rect 21349 14087 21383 14121
rect 21417 14087 21451 14121
rect 21485 14087 21519 14121
rect 21553 14087 21587 14121
rect 21621 14087 21655 14121
rect 21689 14087 21723 14121
rect 21757 14087 21791 14121
rect 21825 14087 21859 14121
rect 21893 14087 21927 14121
rect 21961 14087 21995 14121
rect 22029 14087 22063 14121
rect 22097 14087 22131 14121
rect 22165 14087 22199 14121
rect 22233 14087 22267 14121
rect 22301 14087 22335 14121
rect 22369 14087 22403 14121
rect 22437 14087 22471 14121
rect 22505 14087 22539 14121
rect 22573 14087 22607 14121
rect 22641 14087 22675 14121
rect 22709 14087 22743 14121
rect 22777 14087 22811 14121
rect 22845 14087 22879 14121
rect 22913 14087 22947 14121
rect 22981 14087 23015 14121
rect 23049 14087 23083 14121
rect 23117 14087 23151 14121
rect 23185 14087 23219 14121
rect 23253 14087 23287 14121
rect 23321 14087 23355 14121
rect 23389 14087 23423 14121
rect 23457 14087 23491 14121
rect 23525 14087 23559 14121
rect 23593 14087 23627 14121
rect 23661 14087 23695 14121
rect 23729 14087 23763 14121
rect 23797 14087 23831 14121
rect 23865 14087 23899 14121
rect 23933 14087 23967 14121
rect 24001 14087 24035 14121
rect 24069 14087 24103 14121
rect 24137 14087 24171 14121
rect 24205 14087 24239 14121
rect 24273 14087 24307 14121
rect 24341 14087 24375 14121
rect 24409 14087 24443 14121
rect 24477 14087 24511 14121
rect 24545 14087 24579 14121
rect 24613 14087 24647 14121
rect 24681 14087 24715 14121
rect 24749 14087 24783 14121
rect 24817 14087 24851 14121
rect 24885 14087 24919 14121
rect 24953 14087 24987 14121
rect 25021 14087 25055 14121
rect 25089 14087 25123 14121
rect 25157 14087 25191 14121
rect 25225 14087 25259 14121
rect 25293 14087 25327 14121
rect 25361 14087 25395 14121
rect 25429 14087 25463 14121
rect 25497 14087 25531 14121
rect 25565 14087 25599 14121
rect 25633 14087 25667 14121
rect 25701 14087 25735 14121
rect 25769 14087 25803 14121
rect 25837 14087 25871 14121
rect 25905 14087 25939 14121
rect 25973 14087 26007 14121
rect 26041 14087 26075 14121
rect 26109 14087 26143 14121
rect 26177 14087 26211 14121
rect 26245 14087 26279 14121
rect 26313 14087 26347 14121
rect 26381 14087 26415 14121
rect 26449 14087 26483 14121
rect 26517 14087 26551 14121
rect 26585 14087 26619 14121
rect 26653 14087 26687 14121
rect 26721 14087 26755 14121
rect 26789 14087 26823 14121
rect 26857 14087 26891 14121
rect 26925 14087 26959 14121
rect 26993 14087 27027 14121
rect 27061 14087 27095 14121
rect 27129 14087 27163 14121
rect 27197 14087 27231 14121
rect 27265 14087 27299 14121
rect 27333 14087 27367 14121
rect 27401 14087 27435 14121
rect 27469 14087 27503 14121
rect 27537 14087 27571 14121
rect 27605 14087 27639 14121
rect 27673 14087 27707 14121
rect 27741 14087 27775 14121
rect 27809 14087 27843 14121
rect 27877 14087 27911 14121
rect 27945 14087 27979 14121
rect 28013 14087 28047 14121
rect 28081 14087 28115 14121
rect 28149 14087 28183 14121
rect 28217 14087 28251 14121
rect 28285 14087 28319 14121
rect 28353 14087 28387 14121
rect 28421 14087 28455 14121
rect 28489 14087 28523 14121
rect 28557 14087 28591 14121
rect 28625 14087 28659 14121
rect 28693 14087 28727 14121
rect 28761 14087 28795 14121
rect 28829 14087 28863 14121
rect 28897 14087 28931 14121
rect 28965 14087 28999 14121
rect 29033 14087 29067 14121
rect 29101 14087 29135 14121
rect 29169 14087 29203 14121
rect 29237 14087 29271 14121
rect 29305 14087 29339 14121
rect 29373 14087 29407 14121
rect 29441 14087 29475 14121
rect 29509 14087 29543 14121
rect 29577 14087 29611 14121
rect 29645 14087 29669 14121
rect 15831 14084 29669 14087
rect 15831 14061 18681 14084
rect 15831 14027 15855 14061
rect 15889 14027 15925 14061
rect 15959 14027 15995 14061
rect 16029 14027 16065 14061
rect 16099 14027 16135 14061
rect 16169 14027 16205 14061
rect 16239 14027 16275 14061
rect 16309 14027 16345 14061
rect 16379 14027 16415 14061
rect 16449 14027 16485 14061
rect 16519 14027 16555 14061
rect 16589 14027 16625 14061
rect 16659 14027 16695 14061
rect 16729 14027 16765 14061
rect 16799 14027 16835 14061
rect 16869 14027 16905 14061
rect 16939 14027 16975 14061
rect 17009 14027 17045 14061
rect 17079 14027 17115 14061
rect 17149 14027 17185 14061
rect 17219 14027 17255 14061
rect 17289 14027 17324 14061
rect 17358 14027 17393 14061
rect 17427 14027 17462 14061
rect 17496 14027 17531 14061
rect 17565 14027 17600 14061
rect 17634 14027 17669 14061
rect 17703 14027 17738 14061
rect 17772 14027 17807 14061
rect 17841 14027 17876 14061
rect 17910 14027 17945 14061
rect 17979 14027 18014 14061
rect 18048 14027 18083 14061
rect 18117 14027 18152 14061
rect 18186 14027 18221 14061
rect 18255 14027 18290 14061
rect 18324 14027 18359 14061
rect 18393 14027 18428 14061
rect 18462 14058 18681 14061
rect 18462 14027 18500 14058
rect 15831 14024 18500 14027
rect 18534 14055 18681 14058
rect 18534 14024 18572 14055
rect 15831 14021 18572 14024
rect 18606 14051 18681 14055
rect 18606 14021 18644 14051
rect 15831 14017 18644 14021
rect 18678 14017 18681 14051
rect 15831 13989 18681 14017
rect 15831 13955 15855 13989
rect 15889 13955 15925 13989
rect 15959 13955 15995 13989
rect 16029 13955 16065 13989
rect 16099 13955 16135 13989
rect 16169 13955 16205 13989
rect 16239 13955 16275 13989
rect 16309 13955 16345 13989
rect 16379 13955 16415 13989
rect 16449 13955 16485 13989
rect 16519 13955 16555 13989
rect 16589 13955 16625 13989
rect 16659 13955 16695 13989
rect 16729 13955 16765 13989
rect 16799 13955 16835 13989
rect 16869 13955 16905 13989
rect 16939 13955 16975 13989
rect 17009 13955 17045 13989
rect 17079 13955 17115 13989
rect 17149 13955 17185 13989
rect 17219 13955 17255 13989
rect 17289 13955 17325 13989
rect 17359 13955 17395 13989
rect 17429 13955 17465 13989
rect 17499 13955 17534 13989
rect 17568 13955 17603 13989
rect 17637 13955 17672 13989
rect 17706 13955 17741 13989
rect 17775 13955 17810 13989
rect 17844 13955 17879 13989
rect 17913 13955 17948 13989
rect 17982 13955 18017 13989
rect 18051 13955 18086 13989
rect 18120 13955 18155 13989
rect 18189 13955 18224 13989
rect 18258 13955 18293 13989
rect 18327 13955 18362 13989
rect 18396 13955 18431 13989
rect 18465 13955 18500 13989
rect 18534 13986 18681 13989
rect 18534 13955 18572 13986
rect 15831 13952 18572 13955
rect 18606 13981 18681 13986
rect 18606 13952 18644 13981
rect 15831 13947 18644 13952
rect 18678 13947 18681 13981
rect 15831 13917 18681 13947
rect 15831 13883 15855 13917
rect 15889 13883 15925 13917
rect 15959 13883 15995 13917
rect 16029 13883 16065 13917
rect 16099 13883 16135 13917
rect 16169 13883 16205 13917
rect 16239 13883 16275 13917
rect 16309 13883 16345 13917
rect 16379 13883 16415 13917
rect 16449 13883 16485 13917
rect 16519 13883 16555 13917
rect 16589 13883 16625 13917
rect 16659 13883 16695 13917
rect 16729 13883 16765 13917
rect 16799 13883 16835 13917
rect 16869 13883 16905 13917
rect 16939 13883 16975 13917
rect 17009 13883 17045 13917
rect 17079 13883 17115 13917
rect 17149 13883 17185 13917
rect 17219 13883 17255 13917
rect 17289 13883 17325 13917
rect 17359 13883 17395 13917
rect 17429 13883 17465 13917
rect 17499 13883 17535 13917
rect 17569 13883 17605 13917
rect 17639 13883 17675 13917
rect 17709 13883 17744 13917
rect 17778 13883 17813 13917
rect 17847 13883 17882 13917
rect 17916 13883 17951 13917
rect 17985 13883 18020 13917
rect 18054 13883 18089 13917
rect 18123 13883 18158 13917
rect 18192 13883 18227 13917
rect 18261 13883 18296 13917
rect 18330 13883 18365 13917
rect 18399 13883 18434 13917
rect 18468 13883 18503 13917
rect 18537 13883 18572 13917
rect 18606 13910 18681 13917
rect 18606 13883 18644 13910
rect 15831 13876 18644 13883
rect 18678 13876 18681 13910
rect 15831 13845 18681 13876
rect 15831 13811 15855 13845
rect 15889 13811 15924 13845
rect 15958 13811 15993 13845
rect 16027 13811 16062 13845
rect 16096 13811 16131 13845
rect 16165 13811 16199 13845
rect 16233 13811 16267 13845
rect 16301 13811 16335 13845
rect 16369 13811 16403 13845
rect 16437 13811 16471 13845
rect 16505 13811 16539 13845
rect 16573 13811 16607 13845
rect 16641 13811 16675 13845
rect 16709 13811 16743 13845
rect 16777 13811 16811 13845
rect 16845 13811 16879 13845
rect 16913 13811 16947 13845
rect 16981 13811 17015 13845
rect 17049 13811 17083 13845
rect 17117 13811 17151 13845
rect 17185 13811 17219 13845
rect 17253 13811 17287 13845
rect 17321 13811 17355 13845
rect 17389 13811 17423 13845
rect 17457 13811 17491 13845
rect 17525 13811 17559 13845
rect 17593 13811 17627 13845
rect 17661 13811 17695 13845
rect 17729 13811 17763 13845
rect 17797 13811 17831 13845
rect 17865 13811 17899 13845
rect 17933 13811 17967 13845
rect 18001 13811 18035 13845
rect 18069 13811 18103 13845
rect 18137 13811 18171 13845
rect 18205 13811 18239 13845
rect 18273 13811 18307 13845
rect 18341 13811 18375 13845
rect 18409 13811 18443 13845
rect 18477 13811 18511 13845
rect 18545 13811 18579 13845
rect 18613 13811 18681 13845
rect 15831 13808 18681 13811
rect 13224 12087 13279 12121
rect 13313 12087 13347 12121
rect 13381 12087 13415 12121
rect 13449 12087 13483 12121
rect 13517 12087 13551 12121
rect 13585 12087 13619 12121
rect 13653 12087 13687 12121
rect 13721 12087 13755 12121
rect 13789 12087 13823 12121
rect 13857 12087 13891 12121
rect 13925 12087 13959 12121
rect 13993 12087 14027 12121
rect 14061 12087 14095 12121
rect 14129 12087 14163 12121
rect 14197 12087 14231 12121
rect 14265 12087 14299 12121
rect 14333 12087 14367 12121
rect 14401 12087 14435 12121
rect 14469 12087 14503 12121
rect 14537 12087 14571 12121
rect 14605 12087 14639 12121
rect 14673 12087 14707 12121
rect 14741 12087 14775 12121
rect 14809 12087 14843 12121
rect 14877 12087 14911 12121
rect 14945 12087 14979 12121
rect 15013 12087 15047 12121
rect 15081 12087 15115 12121
rect 15149 12087 15183 12121
rect 15217 12087 15251 12121
rect 15285 12087 15319 12121
rect 15353 12087 15387 12121
rect 15421 12087 15455 12121
rect 15489 12087 15523 12121
rect 15557 12087 15591 12121
rect 15625 12087 15659 12121
rect 15693 12087 15727 12121
rect 15761 12087 15795 12121
rect 15829 12087 15884 12121
rect 13224 12052 15884 12087
rect 13224 12018 13279 12052
rect 13313 12018 13347 12052
rect 13381 12018 13415 12052
rect 13449 12018 13483 12052
rect 13517 12018 13551 12052
rect 13585 12018 13619 12052
rect 13653 12018 13687 12052
rect 13721 12018 13755 12052
rect 13789 12018 13823 12052
rect 13857 12018 13891 12052
rect 13925 12018 13959 12052
rect 13993 12018 14027 12052
rect 14061 12018 14095 12052
rect 14129 12018 14163 12052
rect 14197 12018 14231 12052
rect 14265 12018 14299 12052
rect 14333 12018 14367 12052
rect 14401 12018 14435 12052
rect 14469 12018 14503 12052
rect 14537 12018 14571 12052
rect 14605 12018 14639 12052
rect 14673 12018 14707 12052
rect 14741 12018 14775 12052
rect 14809 12018 14843 12052
rect 14877 12018 14911 12052
rect 14945 12018 14979 12052
rect 15013 12018 15047 12052
rect 15081 12018 15115 12052
rect 15149 12018 15183 12052
rect 15217 12018 15251 12052
rect 15285 12018 15319 12052
rect 15353 12018 15387 12052
rect 15421 12018 15455 12052
rect 15489 12018 15523 12052
rect 15557 12018 15591 12052
rect 15625 12018 15659 12052
rect 15693 12018 15727 12052
rect 15761 12018 15795 12052
rect 15829 12018 15884 12052
rect 13224 11983 15884 12018
rect 13224 11949 13279 11983
rect 13313 11949 13347 11983
rect 13381 11949 13415 11983
rect 13449 11949 13483 11983
rect 13517 11949 13551 11983
rect 13585 11949 13619 11983
rect 13653 11949 13687 11983
rect 13721 11949 13755 11983
rect 13789 11949 13823 11983
rect 13857 11949 13891 11983
rect 13925 11949 13959 11983
rect 13993 11949 14027 11983
rect 14061 11949 14095 11983
rect 14129 11949 14163 11983
rect 14197 11949 14231 11983
rect 14265 11949 14299 11983
rect 14333 11949 14367 11983
rect 14401 11949 14435 11983
rect 14469 11949 14503 11983
rect 14537 11949 14571 11983
rect 14605 11949 14639 11983
rect 14673 11949 14707 11983
rect 14741 11949 14775 11983
rect 14809 11949 14843 11983
rect 14877 11949 14911 11983
rect 14945 11949 14979 11983
rect 15013 11949 15047 11983
rect 15081 11949 15115 11983
rect 15149 11949 15183 11983
rect 15217 11949 15251 11983
rect 15285 11949 15319 11983
rect 15353 11949 15387 11983
rect 15421 11949 15455 11983
rect 15489 11949 15523 11983
rect 15557 11949 15591 11983
rect 15625 11949 15659 11983
rect 15693 11949 15727 11983
rect 15761 11949 15795 11983
rect 15829 11949 15884 11983
rect -2966 10378 -266 10413
rect -2966 10344 -2959 10378
rect -2925 10344 -2891 10378
rect -2857 10344 -2823 10378
rect -2789 10344 -2755 10378
rect -2721 10344 -2687 10378
rect -2653 10344 -2619 10378
rect -2585 10344 -2551 10378
rect -2517 10344 -2483 10378
rect -2449 10344 -2415 10378
rect -2381 10344 -2347 10378
rect -2313 10344 -2279 10378
rect -2245 10344 -2211 10378
rect -2177 10344 -2143 10378
rect -2109 10344 -2075 10378
rect -2041 10344 -2007 10378
rect -1973 10344 -1939 10378
rect -1905 10344 -1871 10378
rect -1837 10344 -1803 10378
rect -1769 10344 -1735 10378
rect -1701 10344 -1667 10378
rect -1633 10344 -1599 10378
rect -1565 10344 -1531 10378
rect -1497 10344 -1463 10378
rect -1429 10344 -1395 10378
rect -1361 10344 -1327 10378
rect -1293 10344 -1259 10378
rect -1225 10344 -1191 10378
rect -1157 10344 -1123 10378
rect -1089 10344 -1055 10378
rect -1021 10344 -987 10378
rect -953 10344 -919 10378
rect -885 10344 -851 10378
rect -817 10344 -783 10378
rect -749 10344 -715 10378
rect -681 10344 -647 10378
rect -613 10344 -579 10378
rect -545 10344 -511 10378
rect -477 10344 -443 10378
rect -409 10344 -375 10378
rect -341 10344 -307 10378
rect -273 10344 -266 10378
rect -2966 10309 -266 10344
rect -2966 10275 -2959 10309
rect -2925 10275 -2891 10309
rect -2857 10275 -2823 10309
rect -2789 10275 -2755 10309
rect -2721 10275 -2687 10309
rect -2653 10275 -2619 10309
rect -2585 10275 -2551 10309
rect -2517 10275 -2483 10309
rect -2449 10275 -2415 10309
rect -2381 10275 -2347 10309
rect -2313 10275 -2279 10309
rect -2245 10275 -2211 10309
rect -2177 10275 -2143 10309
rect -2109 10275 -2075 10309
rect -2041 10275 -2007 10309
rect -1973 10275 -1939 10309
rect -1905 10275 -1871 10309
rect -1837 10275 -1803 10309
rect -1769 10275 -1735 10309
rect -1701 10275 -1667 10309
rect -1633 10275 -1599 10309
rect -1565 10275 -1531 10309
rect -1497 10275 -1463 10309
rect -1429 10275 -1395 10309
rect -1361 10275 -1327 10309
rect -1293 10275 -1259 10309
rect -1225 10275 -1191 10309
rect -1157 10275 -1123 10309
rect -1089 10275 -1055 10309
rect -1021 10275 -987 10309
rect -953 10275 -919 10309
rect -885 10275 -851 10309
rect -817 10275 -783 10309
rect -749 10275 -715 10309
rect -681 10275 -647 10309
rect -613 10275 -579 10309
rect -545 10275 -511 10309
rect -477 10275 -443 10309
rect -409 10275 -375 10309
rect -341 10275 -307 10309
rect -273 10275 -266 10309
rect -2966 10240 -266 10275
rect -2966 10206 -2959 10240
rect -2925 10206 -2891 10240
rect -2857 10206 -2823 10240
rect -2789 10206 -2755 10240
rect -2721 10206 -2687 10240
rect -2653 10206 -2619 10240
rect -2585 10206 -2551 10240
rect -2517 10206 -2483 10240
rect -2449 10206 -2415 10240
rect -2381 10206 -2347 10240
rect -2313 10206 -2279 10240
rect -2245 10206 -2211 10240
rect -2177 10206 -2143 10240
rect -2109 10206 -2075 10240
rect -2041 10206 -2007 10240
rect -1973 10206 -1939 10240
rect -1905 10206 -1871 10240
rect -1837 10206 -1803 10240
rect -1769 10206 -1735 10240
rect -1701 10206 -1667 10240
rect -1633 10206 -1599 10240
rect -1565 10206 -1531 10240
rect -1497 10206 -1463 10240
rect -1429 10206 -1395 10240
rect -1361 10206 -1327 10240
rect -1293 10206 -1259 10240
rect -1225 10206 -1191 10240
rect -1157 10206 -1123 10240
rect -1089 10206 -1055 10240
rect -1021 10206 -987 10240
rect -953 10206 -919 10240
rect -885 10206 -851 10240
rect -817 10206 -783 10240
rect -749 10206 -715 10240
rect -681 10206 -647 10240
rect -613 10206 -579 10240
rect -545 10206 -511 10240
rect -477 10206 -443 10240
rect -409 10206 -375 10240
rect -341 10206 -307 10240
rect -273 10206 -266 10240
rect -2966 10171 -266 10206
rect -2966 10137 -2959 10171
rect -2925 10137 -2891 10171
rect -2857 10137 -2823 10171
rect -2789 10137 -2755 10171
rect -2721 10137 -2687 10171
rect -2653 10137 -2619 10171
rect -2585 10137 -2551 10171
rect -2517 10137 -2483 10171
rect -2449 10137 -2415 10171
rect -2381 10137 -2347 10171
rect -2313 10137 -2279 10171
rect -2245 10137 -2211 10171
rect -2177 10137 -2143 10171
rect -2109 10137 -2075 10171
rect -2041 10137 -2007 10171
rect -1973 10137 -1939 10171
rect -1905 10137 -1871 10171
rect -1837 10137 -1803 10171
rect -1769 10137 -1735 10171
rect -1701 10137 -1667 10171
rect -1633 10137 -1599 10171
rect -1565 10137 -1531 10171
rect -1497 10137 -1463 10171
rect -1429 10137 -1395 10171
rect -1361 10137 -1327 10171
rect -1293 10137 -1259 10171
rect -1225 10137 -1191 10171
rect -1157 10137 -1123 10171
rect -1089 10137 -1055 10171
rect -1021 10137 -987 10171
rect -953 10137 -919 10171
rect -885 10137 -851 10171
rect -817 10137 -783 10171
rect -749 10137 -715 10171
rect -681 10137 -647 10171
rect -613 10137 -579 10171
rect -545 10137 -511 10171
rect -477 10137 -443 10171
rect -409 10137 -375 10171
rect -341 10137 -307 10171
rect -273 10137 -266 10171
rect -2966 10102 -266 10137
rect -2966 10068 -2959 10102
rect -2925 10068 -2891 10102
rect -2857 10068 -2823 10102
rect -2789 10068 -2755 10102
rect -2721 10068 -2687 10102
rect -2653 10068 -2619 10102
rect -2585 10068 -2551 10102
rect -2517 10068 -2483 10102
rect -2449 10068 -2415 10102
rect -2381 10068 -2347 10102
rect -2313 10068 -2279 10102
rect -2245 10068 -2211 10102
rect -2177 10068 -2143 10102
rect -2109 10068 -2075 10102
rect -2041 10068 -2007 10102
rect -1973 10068 -1939 10102
rect -1905 10068 -1871 10102
rect -1837 10068 -1803 10102
rect -1769 10068 -1735 10102
rect -1701 10068 -1667 10102
rect -1633 10068 -1599 10102
rect -1565 10068 -1531 10102
rect -1497 10068 -1463 10102
rect -1429 10068 -1395 10102
rect -1361 10068 -1327 10102
rect -1293 10068 -1259 10102
rect -1225 10068 -1191 10102
rect -1157 10068 -1123 10102
rect -1089 10068 -1055 10102
rect -1021 10068 -987 10102
rect -953 10068 -919 10102
rect -885 10068 -851 10102
rect -817 10068 -783 10102
rect -749 10068 -715 10102
rect -681 10068 -647 10102
rect -613 10068 -579 10102
rect -545 10068 -511 10102
rect -477 10068 -443 10102
rect -409 10068 -375 10102
rect -341 10068 -307 10102
rect -273 10068 -266 10102
rect -2966 10033 -266 10068
rect 13224 11914 15884 11949
rect 13224 11880 13279 11914
rect 13313 11880 13347 11914
rect 13381 11880 13415 11914
rect 13449 11880 13483 11914
rect 13517 11880 13551 11914
rect 13585 11880 13619 11914
rect 13653 11880 13687 11914
rect 13721 11880 13755 11914
rect 13789 11880 13823 11914
rect 13857 11880 13891 11914
rect 13925 11880 13959 11914
rect 13993 11880 14027 11914
rect 14061 11880 14095 11914
rect 14129 11880 14163 11914
rect 14197 11880 14231 11914
rect 14265 11880 14299 11914
rect 14333 11880 14367 11914
rect 14401 11880 14435 11914
rect 14469 11880 14503 11914
rect 14537 11880 14571 11914
rect 14605 11880 14639 11914
rect 14673 11880 14707 11914
rect 14741 11880 14775 11914
rect 14809 11880 14843 11914
rect 14877 11880 14911 11914
rect 14945 11880 14979 11914
rect 15013 11880 15047 11914
rect 15081 11880 15115 11914
rect 15149 11880 15183 11914
rect 15217 11880 15251 11914
rect 15285 11880 15319 11914
rect 15353 11880 15387 11914
rect 15421 11880 15455 11914
rect 15489 11880 15523 11914
rect 15557 11880 15591 11914
rect 15625 11880 15659 11914
rect 15693 11880 15727 11914
rect 15761 11880 15795 11914
rect 15829 11880 15884 11914
rect 13224 11845 15884 11880
rect 13224 11811 13279 11845
rect 13313 11811 13347 11845
rect 13381 11811 13415 11845
rect 13449 11811 13483 11845
rect 13517 11811 13551 11845
rect 13585 11811 13619 11845
rect 13653 11811 13687 11845
rect 13721 11811 13755 11845
rect 13789 11811 13823 11845
rect 13857 11811 13891 11845
rect 13925 11811 13959 11845
rect 13993 11811 14027 11845
rect 14061 11811 14095 11845
rect 14129 11811 14163 11845
rect 14197 11811 14231 11845
rect 14265 11811 14299 11845
rect 14333 11811 14367 11845
rect 14401 11811 14435 11845
rect 14469 11811 14503 11845
rect 14537 11811 14571 11845
rect 14605 11811 14639 11845
rect 14673 11811 14707 11845
rect 14741 11811 14775 11845
rect 14809 11811 14843 11845
rect 14877 11811 14911 11845
rect 14945 11811 14979 11845
rect 15013 11811 15047 11845
rect 15081 11811 15115 11845
rect 15149 11811 15183 11845
rect 15217 11811 15251 11845
rect 15285 11811 15319 11845
rect 15353 11811 15387 11845
rect 15421 11811 15455 11845
rect 15489 11811 15523 11845
rect 15557 11811 15591 11845
rect 15625 11811 15659 11845
rect 15693 11811 15727 11845
rect 15761 11811 15795 11845
rect 15829 11811 15884 11845
rect 13224 11776 15884 11811
rect 13224 11742 13279 11776
rect 13313 11742 13347 11776
rect 13381 11742 13415 11776
rect 13449 11742 13483 11776
rect 13517 11742 13551 11776
rect 13585 11742 13619 11776
rect 13653 11742 13687 11776
rect 13721 11742 13755 11776
rect 13789 11742 13823 11776
rect 13857 11742 13891 11776
rect 13925 11742 13959 11776
rect 13993 11742 14027 11776
rect 14061 11742 14095 11776
rect 14129 11742 14163 11776
rect 14197 11742 14231 11776
rect 14265 11742 14299 11776
rect 14333 11742 14367 11776
rect 14401 11742 14435 11776
rect 14469 11742 14503 11776
rect 14537 11742 14571 11776
rect 14605 11742 14639 11776
rect 14673 11742 14707 11776
rect 14741 11742 14775 11776
rect 14809 11742 14843 11776
rect 14877 11742 14911 11776
rect 14945 11742 14979 11776
rect 15013 11742 15047 11776
rect 15081 11742 15115 11776
rect 15149 11742 15183 11776
rect 15217 11742 15251 11776
rect 15285 11742 15319 11776
rect 15353 11742 15387 11776
rect 15421 11742 15455 11776
rect 15489 11742 15523 11776
rect 15557 11742 15591 11776
rect 15625 11742 15659 11776
rect 15693 11742 15727 11776
rect 15761 11742 15795 11776
rect 15829 11742 15884 11776
rect 13224 11707 15884 11742
rect 13224 11673 13279 11707
rect 13313 11673 13347 11707
rect 13381 11673 13415 11707
rect 13449 11673 13483 11707
rect 13517 11673 13551 11707
rect 13585 11673 13619 11707
rect 13653 11673 13687 11707
rect 13721 11673 13755 11707
rect 13789 11673 13823 11707
rect 13857 11673 13891 11707
rect 13925 11673 13959 11707
rect 13993 11673 14027 11707
rect 14061 11673 14095 11707
rect 14129 11673 14163 11707
rect 14197 11673 14231 11707
rect 14265 11673 14299 11707
rect 14333 11673 14367 11707
rect 14401 11673 14435 11707
rect 14469 11673 14503 11707
rect 14537 11673 14571 11707
rect 14605 11673 14639 11707
rect 14673 11673 14707 11707
rect 14741 11673 14775 11707
rect 14809 11673 14843 11707
rect 14877 11673 14911 11707
rect 14945 11673 14979 11707
rect 15013 11673 15047 11707
rect 15081 11673 15115 11707
rect 15149 11673 15183 11707
rect 15217 11673 15251 11707
rect 15285 11673 15319 11707
rect 15353 11673 15387 11707
rect 15421 11673 15455 11707
rect 15489 11673 15523 11707
rect 15557 11673 15591 11707
rect 15625 11673 15659 11707
rect 15693 11673 15727 11707
rect 15761 11673 15795 11707
rect 15829 11673 15884 11707
rect 13224 11638 15884 11673
rect 13224 11604 13279 11638
rect 13313 11604 13347 11638
rect 13381 11604 13415 11638
rect 13449 11604 13483 11638
rect 13517 11604 13551 11638
rect 13585 11604 13619 11638
rect 13653 11604 13687 11638
rect 13721 11604 13755 11638
rect 13789 11604 13823 11638
rect 13857 11604 13891 11638
rect 13925 11604 13959 11638
rect 13993 11604 14027 11638
rect 14061 11604 14095 11638
rect 14129 11604 14163 11638
rect 14197 11604 14231 11638
rect 14265 11604 14299 11638
rect 14333 11604 14367 11638
rect 14401 11604 14435 11638
rect 14469 11604 14503 11638
rect 14537 11604 14571 11638
rect 14605 11604 14639 11638
rect 14673 11604 14707 11638
rect 14741 11604 14775 11638
rect 14809 11604 14843 11638
rect 14877 11604 14911 11638
rect 14945 11604 14979 11638
rect 15013 11604 15047 11638
rect 15081 11604 15115 11638
rect 15149 11604 15183 11638
rect 15217 11604 15251 11638
rect 15285 11604 15319 11638
rect 15353 11604 15387 11638
rect 15421 11604 15455 11638
rect 15489 11604 15523 11638
rect 15557 11604 15591 11638
rect 15625 11604 15659 11638
rect 15693 11604 15727 11638
rect 15761 11604 15795 11638
rect 15829 11604 15884 11638
rect 13224 11569 15884 11604
rect 13224 11535 13279 11569
rect 13313 11535 13347 11569
rect 13381 11535 13415 11569
rect 13449 11535 13483 11569
rect 13517 11535 13551 11569
rect 13585 11535 13619 11569
rect 13653 11535 13687 11569
rect 13721 11535 13755 11569
rect 13789 11535 13823 11569
rect 13857 11535 13891 11569
rect 13925 11535 13959 11569
rect 13993 11535 14027 11569
rect 14061 11535 14095 11569
rect 14129 11535 14163 11569
rect 14197 11535 14231 11569
rect 14265 11535 14299 11569
rect 14333 11535 14367 11569
rect 14401 11535 14435 11569
rect 14469 11535 14503 11569
rect 14537 11535 14571 11569
rect 14605 11535 14639 11569
rect 14673 11535 14707 11569
rect 14741 11535 14775 11569
rect 14809 11535 14843 11569
rect 14877 11535 14911 11569
rect 14945 11535 14979 11569
rect 15013 11535 15047 11569
rect 15081 11535 15115 11569
rect 15149 11535 15183 11569
rect 15217 11535 15251 11569
rect 15285 11535 15319 11569
rect 15353 11535 15387 11569
rect 15421 11535 15455 11569
rect 15489 11535 15523 11569
rect 15557 11535 15591 11569
rect 15625 11535 15659 11569
rect 15693 11535 15727 11569
rect 15761 11535 15795 11569
rect 15829 11535 15884 11569
rect 13224 11499 15884 11535
rect 13224 11465 13279 11499
rect 13313 11465 13347 11499
rect 13381 11465 13415 11499
rect 13449 11465 13483 11499
rect 13517 11465 13551 11499
rect 13585 11465 13619 11499
rect 13653 11465 13687 11499
rect 13721 11465 13755 11499
rect 13789 11465 13823 11499
rect 13857 11465 13891 11499
rect 13925 11465 13959 11499
rect 13993 11465 14027 11499
rect 14061 11465 14095 11499
rect 14129 11465 14163 11499
rect 14197 11465 14231 11499
rect 14265 11465 14299 11499
rect 14333 11465 14367 11499
rect 14401 11465 14435 11499
rect 14469 11465 14503 11499
rect 14537 11465 14571 11499
rect 14605 11465 14639 11499
rect 14673 11465 14707 11499
rect 14741 11465 14775 11499
rect 14809 11465 14843 11499
rect 14877 11465 14911 11499
rect 14945 11465 14979 11499
rect 15013 11465 15047 11499
rect 15081 11465 15115 11499
rect 15149 11465 15183 11499
rect 15217 11465 15251 11499
rect 15285 11465 15319 11499
rect 15353 11465 15387 11499
rect 15421 11465 15455 11499
rect 15489 11465 15523 11499
rect 15557 11465 15591 11499
rect 15625 11465 15659 11499
rect 15693 11465 15727 11499
rect 15761 11465 15795 11499
rect 15829 11465 15884 11499
rect 13224 11429 15884 11465
rect 13224 11395 13279 11429
rect 13313 11395 13347 11429
rect 13381 11395 13415 11429
rect 13449 11395 13483 11429
rect 13517 11395 13551 11429
rect 13585 11395 13619 11429
rect 13653 11395 13687 11429
rect 13721 11395 13755 11429
rect 13789 11395 13823 11429
rect 13857 11395 13891 11429
rect 13925 11395 13959 11429
rect 13993 11395 14027 11429
rect 14061 11395 14095 11429
rect 14129 11395 14163 11429
rect 14197 11395 14231 11429
rect 14265 11395 14299 11429
rect 14333 11395 14367 11429
rect 14401 11395 14435 11429
rect 14469 11395 14503 11429
rect 14537 11395 14571 11429
rect 14605 11395 14639 11429
rect 14673 11395 14707 11429
rect 14741 11395 14775 11429
rect 14809 11395 14843 11429
rect 14877 11395 14911 11429
rect 14945 11395 14979 11429
rect 15013 11395 15047 11429
rect 15081 11395 15115 11429
rect 15149 11395 15183 11429
rect 15217 11395 15251 11429
rect 15285 11395 15319 11429
rect 15353 11395 15387 11429
rect 15421 11395 15455 11429
rect 15489 11395 15523 11429
rect 15557 11395 15591 11429
rect 15625 11395 15659 11429
rect 15693 11395 15727 11429
rect 15761 11395 15795 11429
rect 15829 11395 15884 11429
rect 13224 11359 15884 11395
rect 13224 11325 13279 11359
rect 13313 11325 13347 11359
rect 13381 11325 13415 11359
rect 13449 11325 13483 11359
rect 13517 11325 13551 11359
rect 13585 11325 13619 11359
rect 13653 11325 13687 11359
rect 13721 11325 13755 11359
rect 13789 11325 13823 11359
rect 13857 11325 13891 11359
rect 13925 11325 13959 11359
rect 13993 11325 14027 11359
rect 14061 11325 14095 11359
rect 14129 11325 14163 11359
rect 14197 11325 14231 11359
rect 14265 11325 14299 11359
rect 14333 11325 14367 11359
rect 14401 11325 14435 11359
rect 14469 11325 14503 11359
rect 14537 11325 14571 11359
rect 14605 11325 14639 11359
rect 14673 11325 14707 11359
rect 14741 11325 14775 11359
rect 14809 11325 14843 11359
rect 14877 11325 14911 11359
rect 14945 11325 14979 11359
rect 15013 11325 15047 11359
rect 15081 11325 15115 11359
rect 15149 11325 15183 11359
rect 15217 11325 15251 11359
rect 15285 11325 15319 11359
rect 15353 11325 15387 11359
rect 15421 11325 15455 11359
rect 15489 11325 15523 11359
rect 15557 11325 15591 11359
rect 15625 11325 15659 11359
rect 15693 11325 15727 11359
rect 15761 11325 15795 11359
rect 15829 11325 15884 11359
rect 13224 11289 15884 11325
rect 13224 11255 13279 11289
rect 13313 11255 13347 11289
rect 13381 11255 13415 11289
rect 13449 11255 13483 11289
rect 13517 11255 13551 11289
rect 13585 11255 13619 11289
rect 13653 11255 13687 11289
rect 13721 11255 13755 11289
rect 13789 11255 13823 11289
rect 13857 11255 13891 11289
rect 13925 11255 13959 11289
rect 13993 11255 14027 11289
rect 14061 11255 14095 11289
rect 14129 11255 14163 11289
rect 14197 11255 14231 11289
rect 14265 11255 14299 11289
rect 14333 11255 14367 11289
rect 14401 11255 14435 11289
rect 14469 11255 14503 11289
rect 14537 11255 14571 11289
rect 14605 11255 14639 11289
rect 14673 11255 14707 11289
rect 14741 11255 14775 11289
rect 14809 11255 14843 11289
rect 14877 11255 14911 11289
rect 14945 11255 14979 11289
rect 15013 11255 15047 11289
rect 15081 11255 15115 11289
rect 15149 11255 15183 11289
rect 15217 11255 15251 11289
rect 15285 11255 15319 11289
rect 15353 11255 15387 11289
rect 15421 11255 15455 11289
rect 15489 11255 15523 11289
rect 15557 11255 15591 11289
rect 15625 11255 15659 11289
rect 15693 11255 15727 11289
rect 15761 11255 15795 11289
rect 15829 11255 15884 11289
rect 13224 11219 15884 11255
rect 13224 11185 13279 11219
rect 13313 11185 13347 11219
rect 13381 11185 13415 11219
rect 13449 11185 13483 11219
rect 13517 11185 13551 11219
rect 13585 11185 13619 11219
rect 13653 11185 13687 11219
rect 13721 11185 13755 11219
rect 13789 11185 13823 11219
rect 13857 11185 13891 11219
rect 13925 11185 13959 11219
rect 13993 11185 14027 11219
rect 14061 11185 14095 11219
rect 14129 11185 14163 11219
rect 14197 11185 14231 11219
rect 14265 11185 14299 11219
rect 14333 11185 14367 11219
rect 14401 11185 14435 11219
rect 14469 11185 14503 11219
rect 14537 11185 14571 11219
rect 14605 11185 14639 11219
rect 14673 11185 14707 11219
rect 14741 11185 14775 11219
rect 14809 11185 14843 11219
rect 14877 11185 14911 11219
rect 14945 11185 14979 11219
rect 15013 11185 15047 11219
rect 15081 11185 15115 11219
rect 15149 11185 15183 11219
rect 15217 11185 15251 11219
rect 15285 11185 15319 11219
rect 15353 11185 15387 11219
rect 15421 11185 15455 11219
rect 15489 11185 15523 11219
rect 15557 11185 15591 11219
rect 15625 11185 15659 11219
rect 15693 11185 15727 11219
rect 15761 11185 15795 11219
rect 15829 11185 15884 11219
rect 13224 11149 15884 11185
rect 13224 11115 13279 11149
rect 13313 11115 13347 11149
rect 13381 11115 13415 11149
rect 13449 11115 13483 11149
rect 13517 11115 13551 11149
rect 13585 11115 13619 11149
rect 13653 11115 13687 11149
rect 13721 11115 13755 11149
rect 13789 11115 13823 11149
rect 13857 11115 13891 11149
rect 13925 11115 13959 11149
rect 13993 11115 14027 11149
rect 14061 11115 14095 11149
rect 14129 11115 14163 11149
rect 14197 11115 14231 11149
rect 14265 11115 14299 11149
rect 14333 11115 14367 11149
rect 14401 11115 14435 11149
rect 14469 11115 14503 11149
rect 14537 11115 14571 11149
rect 14605 11115 14639 11149
rect 14673 11115 14707 11149
rect 14741 11115 14775 11149
rect 14809 11115 14843 11149
rect 14877 11115 14911 11149
rect 14945 11115 14979 11149
rect 15013 11115 15047 11149
rect 15081 11115 15115 11149
rect 15149 11115 15183 11149
rect 15217 11115 15251 11149
rect 15285 11115 15319 11149
rect 15353 11115 15387 11149
rect 15421 11115 15455 11149
rect 15489 11115 15523 11149
rect 15557 11115 15591 11149
rect 15625 11115 15659 11149
rect 15693 11115 15727 11149
rect 15761 11115 15795 11149
rect 15829 11115 15884 11149
rect 13224 11079 15884 11115
rect 13224 11045 13279 11079
rect 13313 11045 13347 11079
rect 13381 11045 13415 11079
rect 13449 11045 13483 11079
rect 13517 11045 13551 11079
rect 13585 11045 13619 11079
rect 13653 11045 13687 11079
rect 13721 11045 13755 11079
rect 13789 11045 13823 11079
rect 13857 11045 13891 11079
rect 13925 11045 13959 11079
rect 13993 11045 14027 11079
rect 14061 11045 14095 11079
rect 14129 11045 14163 11079
rect 14197 11045 14231 11079
rect 14265 11045 14299 11079
rect 14333 11045 14367 11079
rect 14401 11045 14435 11079
rect 14469 11045 14503 11079
rect 14537 11045 14571 11079
rect 14605 11045 14639 11079
rect 14673 11045 14707 11079
rect 14741 11045 14775 11079
rect 14809 11045 14843 11079
rect 14877 11045 14911 11079
rect 14945 11045 14979 11079
rect 15013 11045 15047 11079
rect 15081 11045 15115 11079
rect 15149 11045 15183 11079
rect 15217 11045 15251 11079
rect 15285 11045 15319 11079
rect 15353 11045 15387 11079
rect 15421 11045 15455 11079
rect 15489 11045 15523 11079
rect 15557 11045 15591 11079
rect 15625 11045 15659 11079
rect 15693 11045 15727 11079
rect 15761 11045 15795 11079
rect 15829 11045 15884 11079
rect 13224 11009 15884 11045
rect 13224 10975 13279 11009
rect 13313 10975 13347 11009
rect 13381 10975 13415 11009
rect 13449 10975 13483 11009
rect 13517 10975 13551 11009
rect 13585 10975 13619 11009
rect 13653 10975 13687 11009
rect 13721 10975 13755 11009
rect 13789 10975 13823 11009
rect 13857 10975 13891 11009
rect 13925 10975 13959 11009
rect 13993 10975 14027 11009
rect 14061 10975 14095 11009
rect 14129 10975 14163 11009
rect 14197 10975 14231 11009
rect 14265 10975 14299 11009
rect 14333 10975 14367 11009
rect 14401 10975 14435 11009
rect 14469 10975 14503 11009
rect 14537 10975 14571 11009
rect 14605 10975 14639 11009
rect 14673 10975 14707 11009
rect 14741 10975 14775 11009
rect 14809 10975 14843 11009
rect 14877 10975 14911 11009
rect 14945 10975 14979 11009
rect 15013 10975 15047 11009
rect 15081 10975 15115 11009
rect 15149 10975 15183 11009
rect 15217 10975 15251 11009
rect 15285 10975 15319 11009
rect 15353 10975 15387 11009
rect 15421 10975 15455 11009
rect 15489 10975 15523 11009
rect 15557 10975 15591 11009
rect 15625 10975 15659 11009
rect 15693 10975 15727 11009
rect 15761 10975 15795 11009
rect 15829 10975 15884 11009
rect 13224 10939 15884 10975
rect 13224 10905 13279 10939
rect 13313 10905 13347 10939
rect 13381 10905 13415 10939
rect 13449 10905 13483 10939
rect 13517 10905 13551 10939
rect 13585 10905 13619 10939
rect 13653 10905 13687 10939
rect 13721 10905 13755 10939
rect 13789 10905 13823 10939
rect 13857 10905 13891 10939
rect 13925 10905 13959 10939
rect 13993 10905 14027 10939
rect 14061 10905 14095 10939
rect 14129 10905 14163 10939
rect 14197 10905 14231 10939
rect 14265 10905 14299 10939
rect 14333 10905 14367 10939
rect 14401 10905 14435 10939
rect 14469 10905 14503 10939
rect 14537 10905 14571 10939
rect 14605 10905 14639 10939
rect 14673 10905 14707 10939
rect 14741 10905 14775 10939
rect 14809 10905 14843 10939
rect 14877 10905 14911 10939
rect 14945 10905 14979 10939
rect 15013 10905 15047 10939
rect 15081 10905 15115 10939
rect 15149 10905 15183 10939
rect 15217 10905 15251 10939
rect 15285 10905 15319 10939
rect 15353 10905 15387 10939
rect 15421 10905 15455 10939
rect 15489 10905 15523 10939
rect 15557 10905 15591 10939
rect 15625 10905 15659 10939
rect 15693 10905 15727 10939
rect 15761 10905 15795 10939
rect 15829 10905 15884 10939
rect 13224 10869 15884 10905
rect 13224 10835 13279 10869
rect 13313 10835 13347 10869
rect 13381 10835 13415 10869
rect 13449 10835 13483 10869
rect 13517 10835 13551 10869
rect 13585 10835 13619 10869
rect 13653 10835 13687 10869
rect 13721 10835 13755 10869
rect 13789 10835 13823 10869
rect 13857 10835 13891 10869
rect 13925 10835 13959 10869
rect 13993 10835 14027 10869
rect 14061 10835 14095 10869
rect 14129 10835 14163 10869
rect 14197 10835 14231 10869
rect 14265 10835 14299 10869
rect 14333 10835 14367 10869
rect 14401 10835 14435 10869
rect 14469 10835 14503 10869
rect 14537 10835 14571 10869
rect 14605 10835 14639 10869
rect 14673 10835 14707 10869
rect 14741 10835 14775 10869
rect 14809 10835 14843 10869
rect 14877 10835 14911 10869
rect 14945 10835 14979 10869
rect 15013 10835 15047 10869
rect 15081 10835 15115 10869
rect 15149 10835 15183 10869
rect 15217 10835 15251 10869
rect 15285 10835 15319 10869
rect 15353 10835 15387 10869
rect 15421 10835 15455 10869
rect 15489 10835 15523 10869
rect 15557 10835 15591 10869
rect 15625 10835 15659 10869
rect 15693 10835 15727 10869
rect 15761 10835 15795 10869
rect 15829 10835 15884 10869
rect 13224 10799 15884 10835
rect 13224 10765 13279 10799
rect 13313 10765 13347 10799
rect 13381 10765 13415 10799
rect 13449 10765 13483 10799
rect 13517 10765 13551 10799
rect 13585 10765 13619 10799
rect 13653 10765 13687 10799
rect 13721 10765 13755 10799
rect 13789 10765 13823 10799
rect 13857 10765 13891 10799
rect 13925 10765 13959 10799
rect 13993 10765 14027 10799
rect 14061 10765 14095 10799
rect 14129 10765 14163 10799
rect 14197 10765 14231 10799
rect 14265 10765 14299 10799
rect 14333 10765 14367 10799
rect 14401 10765 14435 10799
rect 14469 10765 14503 10799
rect 14537 10765 14571 10799
rect 14605 10765 14639 10799
rect 14673 10765 14707 10799
rect 14741 10765 14775 10799
rect 14809 10765 14843 10799
rect 14877 10765 14911 10799
rect 14945 10765 14979 10799
rect 15013 10765 15047 10799
rect 15081 10765 15115 10799
rect 15149 10765 15183 10799
rect 15217 10765 15251 10799
rect 15285 10765 15319 10799
rect 15353 10765 15387 10799
rect 15421 10765 15455 10799
rect 15489 10765 15523 10799
rect 15557 10765 15591 10799
rect 15625 10765 15659 10799
rect 15693 10765 15727 10799
rect 15761 10765 15795 10799
rect 15829 10765 15884 10799
rect 13224 10729 15884 10765
rect 13224 10695 13279 10729
rect 13313 10695 13347 10729
rect 13381 10695 13415 10729
rect 13449 10695 13483 10729
rect 13517 10695 13551 10729
rect 13585 10695 13619 10729
rect 13653 10695 13687 10729
rect 13721 10695 13755 10729
rect 13789 10695 13823 10729
rect 13857 10695 13891 10729
rect 13925 10695 13959 10729
rect 13993 10695 14027 10729
rect 14061 10695 14095 10729
rect 14129 10695 14163 10729
rect 14197 10695 14231 10729
rect 14265 10695 14299 10729
rect 14333 10695 14367 10729
rect 14401 10695 14435 10729
rect 14469 10695 14503 10729
rect 14537 10695 14571 10729
rect 14605 10695 14639 10729
rect 14673 10695 14707 10729
rect 14741 10695 14775 10729
rect 14809 10695 14843 10729
rect 14877 10695 14911 10729
rect 14945 10695 14979 10729
rect 15013 10695 15047 10729
rect 15081 10695 15115 10729
rect 15149 10695 15183 10729
rect 15217 10695 15251 10729
rect 15285 10695 15319 10729
rect 15353 10695 15387 10729
rect 15421 10695 15455 10729
rect 15489 10695 15523 10729
rect 15557 10695 15591 10729
rect 15625 10695 15659 10729
rect 15693 10695 15727 10729
rect 15761 10695 15795 10729
rect 15829 10695 15884 10729
rect 13224 10659 15884 10695
rect 13224 10625 13279 10659
rect 13313 10625 13347 10659
rect 13381 10625 13415 10659
rect 13449 10625 13483 10659
rect 13517 10625 13551 10659
rect 13585 10625 13619 10659
rect 13653 10625 13687 10659
rect 13721 10625 13755 10659
rect 13789 10625 13823 10659
rect 13857 10625 13891 10659
rect 13925 10625 13959 10659
rect 13993 10625 14027 10659
rect 14061 10625 14095 10659
rect 14129 10625 14163 10659
rect 14197 10625 14231 10659
rect 14265 10625 14299 10659
rect 14333 10625 14367 10659
rect 14401 10625 14435 10659
rect 14469 10625 14503 10659
rect 14537 10625 14571 10659
rect 14605 10625 14639 10659
rect 14673 10625 14707 10659
rect 14741 10625 14775 10659
rect 14809 10625 14843 10659
rect 14877 10625 14911 10659
rect 14945 10625 14979 10659
rect 15013 10625 15047 10659
rect 15081 10625 15115 10659
rect 15149 10625 15183 10659
rect 15217 10625 15251 10659
rect 15285 10625 15319 10659
rect 15353 10625 15387 10659
rect 15421 10625 15455 10659
rect 15489 10625 15523 10659
rect 15557 10625 15591 10659
rect 15625 10625 15659 10659
rect 15693 10625 15727 10659
rect 15761 10625 15795 10659
rect 15829 10625 15884 10659
rect 13224 10589 15884 10625
rect 13224 10555 13279 10589
rect 13313 10555 13347 10589
rect 13381 10555 13415 10589
rect 13449 10555 13483 10589
rect 13517 10555 13551 10589
rect 13585 10555 13619 10589
rect 13653 10555 13687 10589
rect 13721 10555 13755 10589
rect 13789 10555 13823 10589
rect 13857 10555 13891 10589
rect 13925 10555 13959 10589
rect 13993 10555 14027 10589
rect 14061 10555 14095 10589
rect 14129 10555 14163 10589
rect 14197 10555 14231 10589
rect 14265 10555 14299 10589
rect 14333 10555 14367 10589
rect 14401 10555 14435 10589
rect 14469 10555 14503 10589
rect 14537 10555 14571 10589
rect 14605 10555 14639 10589
rect 14673 10555 14707 10589
rect 14741 10555 14775 10589
rect 14809 10555 14843 10589
rect 14877 10555 14911 10589
rect 14945 10555 14979 10589
rect 15013 10555 15047 10589
rect 15081 10555 15115 10589
rect 15149 10555 15183 10589
rect 15217 10555 15251 10589
rect 15285 10555 15319 10589
rect 15353 10555 15387 10589
rect 15421 10555 15455 10589
rect 15489 10555 15523 10589
rect 15557 10555 15591 10589
rect 15625 10555 15659 10589
rect 15693 10555 15727 10589
rect 15761 10555 15795 10589
rect 15829 10555 15884 10589
rect 13224 10519 15884 10555
rect 13224 10485 13279 10519
rect 13313 10485 13347 10519
rect 13381 10485 13415 10519
rect 13449 10485 13483 10519
rect 13517 10485 13551 10519
rect 13585 10485 13619 10519
rect 13653 10485 13687 10519
rect 13721 10485 13755 10519
rect 13789 10485 13823 10519
rect 13857 10485 13891 10519
rect 13925 10485 13959 10519
rect 13993 10485 14027 10519
rect 14061 10485 14095 10519
rect 14129 10485 14163 10519
rect 14197 10485 14231 10519
rect 14265 10485 14299 10519
rect 14333 10485 14367 10519
rect 14401 10485 14435 10519
rect 14469 10485 14503 10519
rect 14537 10485 14571 10519
rect 14605 10485 14639 10519
rect 14673 10485 14707 10519
rect 14741 10485 14775 10519
rect 14809 10485 14843 10519
rect 14877 10485 14911 10519
rect 14945 10485 14979 10519
rect 15013 10485 15047 10519
rect 15081 10485 15115 10519
rect 15149 10485 15183 10519
rect 15217 10485 15251 10519
rect 15285 10485 15319 10519
rect 15353 10485 15387 10519
rect 15421 10485 15455 10519
rect 15489 10485 15523 10519
rect 15557 10485 15591 10519
rect 15625 10485 15659 10519
rect 15693 10485 15727 10519
rect 15761 10485 15795 10519
rect 15829 10485 15884 10519
rect 13224 10449 15884 10485
rect 13224 10415 13279 10449
rect 13313 10415 13347 10449
rect 13381 10415 13415 10449
rect 13449 10415 13483 10449
rect 13517 10415 13551 10449
rect 13585 10415 13619 10449
rect 13653 10415 13687 10449
rect 13721 10415 13755 10449
rect 13789 10415 13823 10449
rect 13857 10415 13891 10449
rect 13925 10415 13959 10449
rect 13993 10415 14027 10449
rect 14061 10415 14095 10449
rect 14129 10415 14163 10449
rect 14197 10415 14231 10449
rect 14265 10415 14299 10449
rect 14333 10415 14367 10449
rect 14401 10415 14435 10449
rect 14469 10415 14503 10449
rect 14537 10415 14571 10449
rect 14605 10415 14639 10449
rect 14673 10415 14707 10449
rect 14741 10415 14775 10449
rect 14809 10415 14843 10449
rect 14877 10415 14911 10449
rect 14945 10415 14979 10449
rect 15013 10415 15047 10449
rect 15081 10415 15115 10449
rect 15149 10415 15183 10449
rect 15217 10415 15251 10449
rect 15285 10415 15319 10449
rect 15353 10415 15387 10449
rect 15421 10415 15455 10449
rect 15489 10415 15523 10449
rect 15557 10415 15591 10449
rect 15625 10415 15659 10449
rect 15693 10415 15727 10449
rect 15761 10415 15795 10449
rect 15829 10415 15884 10449
rect 13224 10379 15884 10415
rect 13224 10345 13279 10379
rect 13313 10345 13347 10379
rect 13381 10345 13415 10379
rect 13449 10345 13483 10379
rect 13517 10345 13551 10379
rect 13585 10345 13619 10379
rect 13653 10345 13687 10379
rect 13721 10345 13755 10379
rect 13789 10345 13823 10379
rect 13857 10345 13891 10379
rect 13925 10345 13959 10379
rect 13993 10345 14027 10379
rect 14061 10345 14095 10379
rect 14129 10345 14163 10379
rect 14197 10345 14231 10379
rect 14265 10345 14299 10379
rect 14333 10345 14367 10379
rect 14401 10345 14435 10379
rect 14469 10345 14503 10379
rect 14537 10345 14571 10379
rect 14605 10345 14639 10379
rect 14673 10345 14707 10379
rect 14741 10345 14775 10379
rect 14809 10345 14843 10379
rect 14877 10345 14911 10379
rect 14945 10345 14979 10379
rect 15013 10345 15047 10379
rect 15081 10345 15115 10379
rect 15149 10345 15183 10379
rect 15217 10345 15251 10379
rect 15285 10345 15319 10379
rect 15353 10345 15387 10379
rect 15421 10345 15455 10379
rect 15489 10345 15523 10379
rect 15557 10345 15591 10379
rect 15625 10345 15659 10379
rect 15693 10345 15727 10379
rect 15761 10345 15795 10379
rect 15829 10345 15884 10379
rect 13224 10309 15884 10345
rect 13224 10275 13279 10309
rect 13313 10275 13347 10309
rect 13381 10275 13415 10309
rect 13449 10275 13483 10309
rect 13517 10275 13551 10309
rect 13585 10275 13619 10309
rect 13653 10275 13687 10309
rect 13721 10275 13755 10309
rect 13789 10275 13823 10309
rect 13857 10275 13891 10309
rect 13925 10275 13959 10309
rect 13993 10275 14027 10309
rect 14061 10275 14095 10309
rect 14129 10275 14163 10309
rect 14197 10275 14231 10309
rect 14265 10275 14299 10309
rect 14333 10275 14367 10309
rect 14401 10275 14435 10309
rect 14469 10275 14503 10309
rect 14537 10275 14571 10309
rect 14605 10275 14639 10309
rect 14673 10275 14707 10309
rect 14741 10275 14775 10309
rect 14809 10275 14843 10309
rect 14877 10275 14911 10309
rect 14945 10275 14979 10309
rect 15013 10275 15047 10309
rect 15081 10275 15115 10309
rect 15149 10275 15183 10309
rect 15217 10275 15251 10309
rect 15285 10275 15319 10309
rect 15353 10275 15387 10309
rect 15421 10275 15455 10309
rect 15489 10275 15523 10309
rect 15557 10275 15591 10309
rect 15625 10275 15659 10309
rect 15693 10275 15727 10309
rect 15761 10275 15795 10309
rect 15829 10275 15884 10309
rect 13224 10239 15884 10275
rect 13224 10205 13279 10239
rect 13313 10205 13347 10239
rect 13381 10205 13415 10239
rect 13449 10205 13483 10239
rect 13517 10205 13551 10239
rect 13585 10205 13619 10239
rect 13653 10205 13687 10239
rect 13721 10205 13755 10239
rect 13789 10205 13823 10239
rect 13857 10205 13891 10239
rect 13925 10205 13959 10239
rect 13993 10205 14027 10239
rect 14061 10205 14095 10239
rect 14129 10205 14163 10239
rect 14197 10205 14231 10239
rect 14265 10205 14299 10239
rect 14333 10205 14367 10239
rect 14401 10205 14435 10239
rect 14469 10205 14503 10239
rect 14537 10205 14571 10239
rect 14605 10205 14639 10239
rect 14673 10205 14707 10239
rect 14741 10205 14775 10239
rect 14809 10205 14843 10239
rect 14877 10205 14911 10239
rect 14945 10205 14979 10239
rect 15013 10205 15047 10239
rect 15081 10205 15115 10239
rect 15149 10205 15183 10239
rect 15217 10205 15251 10239
rect 15285 10205 15319 10239
rect 15353 10205 15387 10239
rect 15421 10205 15455 10239
rect 15489 10205 15523 10239
rect 15557 10205 15591 10239
rect 15625 10205 15659 10239
rect 15693 10205 15727 10239
rect 15761 10205 15795 10239
rect 15829 10205 15884 10239
rect 13224 10177 15884 10205
rect 12480 10169 15884 10177
rect 12480 10162 13279 10169
rect 12480 10128 12504 10162
rect 12538 10128 12599 10162
rect 12633 10128 12694 10162
rect 12728 10128 12788 10162
rect 12822 10128 12882 10162
rect 12916 10128 12976 10162
rect 13010 10135 13279 10162
rect 13313 10135 13347 10169
rect 13381 10135 13415 10169
rect 13449 10135 13483 10169
rect 13517 10135 13551 10169
rect 13585 10135 13619 10169
rect 13653 10135 13687 10169
rect 13721 10135 13755 10169
rect 13789 10135 13823 10169
rect 13857 10135 13891 10169
rect 13925 10135 13959 10169
rect 13993 10135 14027 10169
rect 14061 10135 14095 10169
rect 14129 10135 14163 10169
rect 14197 10135 14231 10169
rect 14265 10135 14299 10169
rect 14333 10135 14367 10169
rect 14401 10135 14435 10169
rect 14469 10135 14503 10169
rect 14537 10135 14571 10169
rect 14605 10135 14639 10169
rect 14673 10135 14707 10169
rect 14741 10135 14775 10169
rect 14809 10135 14843 10169
rect 14877 10135 14911 10169
rect 14945 10135 14979 10169
rect 15013 10135 15047 10169
rect 15081 10135 15115 10169
rect 15149 10135 15183 10169
rect 15217 10135 15251 10169
rect 15285 10135 15319 10169
rect 15353 10135 15387 10169
rect 15421 10135 15455 10169
rect 15489 10135 15523 10169
rect 15557 10135 15591 10169
rect 15625 10135 15659 10169
rect 15693 10135 15727 10169
rect 15761 10135 15795 10169
rect 15829 10135 15884 10169
rect 13010 10128 15884 10135
rect 12480 10099 15884 10128
rect 12480 10094 13279 10099
rect -2966 9999 -2959 10033
rect -2925 9999 -2891 10033
rect -2857 9999 -2823 10033
rect -2789 9999 -2755 10033
rect -2721 9999 -2687 10033
rect -2653 9999 -2619 10033
rect -2585 9999 -2551 10033
rect -2517 9999 -2483 10033
rect -2449 9999 -2415 10033
rect -2381 9999 -2347 10033
rect -2313 9999 -2279 10033
rect -2245 9999 -2211 10033
rect -2177 9999 -2143 10033
rect -2109 9999 -2075 10033
rect -2041 9999 -2007 10033
rect -1973 9999 -1939 10033
rect -1905 9999 -1871 10033
rect -1837 9999 -1803 10033
rect -1769 9999 -1735 10033
rect -1701 9999 -1667 10033
rect -1633 9999 -1599 10033
rect -1565 9999 -1531 10033
rect -1497 9999 -1463 10033
rect -1429 9999 -1395 10033
rect -1361 9999 -1327 10033
rect -1293 9999 -1259 10033
rect -1225 9999 -1191 10033
rect -1157 9999 -1123 10033
rect -1089 9999 -1055 10033
rect -1021 9999 -987 10033
rect -953 9999 -919 10033
rect -885 9999 -851 10033
rect -817 9999 -783 10033
rect -749 9999 -715 10033
rect -681 9999 -647 10033
rect -613 9999 -579 10033
rect -545 9999 -511 10033
rect -477 9999 -443 10033
rect -409 9999 -375 10033
rect -341 9999 -307 10033
rect -273 9999 -266 10033
rect -2966 9964 -266 9999
rect -2966 9930 -2959 9964
rect -2925 9930 -2891 9964
rect -2857 9930 -2823 9964
rect -2789 9930 -2755 9964
rect -2721 9930 -2687 9964
rect -2653 9930 -2619 9964
rect -2585 9930 -2551 9964
rect -2517 9930 -2483 9964
rect -2449 9930 -2415 9964
rect -2381 9930 -2347 9964
rect -2313 9930 -2279 9964
rect -2245 9930 -2211 9964
rect -2177 9930 -2143 9964
rect -2109 9930 -2075 9964
rect -2041 9930 -2007 9964
rect -1973 9930 -1939 9964
rect -1905 9930 -1871 9964
rect -1837 9930 -1803 9964
rect -1769 9930 -1735 9964
rect -1701 9930 -1667 9964
rect -1633 9930 -1599 9964
rect -1565 9930 -1531 9964
rect -1497 9930 -1463 9964
rect -1429 9930 -1395 9964
rect -1361 9930 -1327 9964
rect -1293 9930 -1259 9964
rect -1225 9930 -1191 9964
rect -1157 9930 -1123 9964
rect -1089 9930 -1055 9964
rect -1021 9930 -987 9964
rect -953 9930 -919 9964
rect -885 9930 -851 9964
rect -817 9930 -783 9964
rect -749 9930 -715 9964
rect -681 9930 -647 9964
rect -613 9930 -579 9964
rect -545 9930 -511 9964
rect -477 9930 -443 9964
rect -409 9930 -375 9964
rect -341 9930 -307 9964
rect -273 9930 -266 9964
rect 12480 10060 12504 10094
rect 12538 10060 12599 10094
rect 12633 10060 12694 10094
rect 12728 10060 12788 10094
rect 12822 10060 12882 10094
rect 12916 10060 12976 10094
rect 13010 10065 13279 10094
rect 13313 10065 13347 10099
rect 13381 10065 13415 10099
rect 13449 10065 13483 10099
rect 13517 10065 13551 10099
rect 13585 10065 13619 10099
rect 13653 10065 13687 10099
rect 13721 10065 13755 10099
rect 13789 10065 13823 10099
rect 13857 10065 13891 10099
rect 13925 10065 13959 10099
rect 13993 10065 14027 10099
rect 14061 10065 14095 10099
rect 14129 10065 14163 10099
rect 14197 10065 14231 10099
rect 14265 10065 14299 10099
rect 14333 10065 14367 10099
rect 14401 10065 14435 10099
rect 14469 10065 14503 10099
rect 14537 10065 14571 10099
rect 14605 10065 14639 10099
rect 14673 10065 14707 10099
rect 14741 10065 14775 10099
rect 14809 10065 14843 10099
rect 14877 10065 14911 10099
rect 14945 10065 14979 10099
rect 15013 10065 15047 10099
rect 15081 10065 15115 10099
rect 15149 10065 15183 10099
rect 15217 10065 15251 10099
rect 15285 10065 15319 10099
rect 15353 10065 15387 10099
rect 15421 10065 15455 10099
rect 15489 10065 15523 10099
rect 15557 10065 15591 10099
rect 15625 10065 15659 10099
rect 15693 10065 15727 10099
rect 15761 10065 15795 10099
rect 15829 10065 15884 10099
rect 13010 10060 15884 10065
rect 12480 10056 15884 10060
rect 12480 10026 13077 10056
rect 12480 9992 12504 10026
rect 12538 9992 12599 10026
rect 12633 9992 12694 10026
rect 12728 9992 12788 10026
rect 12822 9992 12882 10026
rect 12916 9992 12976 10026
rect 13010 10022 13077 10026
rect 13111 10022 13160 10056
rect 13194 10029 15884 10056
rect 13194 10022 13279 10029
rect 13010 9995 13279 10022
rect 13313 9995 13347 10029
rect 13381 9995 13415 10029
rect 13449 9995 13483 10029
rect 13517 9995 13551 10029
rect 13585 9995 13619 10029
rect 13653 9995 13687 10029
rect 13721 9995 13755 10029
rect 13789 9995 13823 10029
rect 13857 9995 13891 10029
rect 13925 9995 13959 10029
rect 13993 9995 14027 10029
rect 14061 9995 14095 10029
rect 14129 9995 14163 10029
rect 14197 9995 14231 10029
rect 14265 9995 14299 10029
rect 14333 9995 14367 10029
rect 14401 9995 14435 10029
rect 14469 9995 14503 10029
rect 14537 9995 14571 10029
rect 14605 9995 14639 10029
rect 14673 9995 14707 10029
rect 14741 9995 14775 10029
rect 14809 9995 14843 10029
rect 14877 9995 14911 10029
rect 14945 9995 14979 10029
rect 15013 9995 15047 10029
rect 15081 9995 15115 10029
rect 15149 9995 15183 10029
rect 15217 9995 15251 10029
rect 15285 9995 15319 10029
rect 15353 9995 15387 10029
rect 15421 9995 15455 10029
rect 15489 9995 15523 10029
rect 15557 9995 15591 10029
rect 15625 9995 15659 10029
rect 15693 9995 15727 10029
rect 15761 9995 15795 10029
rect 15829 9995 15884 10029
rect 13010 9992 15194 9995
rect 12480 9958 15194 9992
rect -2966 9895 -266 9930
rect -2966 9861 -2959 9895
rect -2925 9861 -2891 9895
rect -2857 9861 -2823 9895
rect -2789 9861 -2755 9895
rect -2721 9861 -2687 9895
rect -2653 9861 -2619 9895
rect -2585 9861 -2551 9895
rect -2517 9861 -2483 9895
rect -2449 9861 -2415 9895
rect -2381 9861 -2347 9895
rect -2313 9861 -2279 9895
rect -2245 9861 -2211 9895
rect -2177 9861 -2143 9895
rect -2109 9861 -2075 9895
rect -2041 9861 -2007 9895
rect -1973 9861 -1939 9895
rect -1905 9861 -1871 9895
rect -1837 9861 -1803 9895
rect -1769 9861 -1735 9895
rect -1701 9861 -1667 9895
rect -1633 9861 -1599 9895
rect -1565 9861 -1531 9895
rect -1497 9861 -1463 9895
rect -1429 9861 -1395 9895
rect -1361 9861 -1327 9895
rect -1293 9861 -1259 9895
rect -1225 9861 -1191 9895
rect -1157 9861 -1123 9895
rect -1089 9861 -1055 9895
rect -1021 9861 -987 9895
rect -953 9861 -919 9895
rect -885 9861 -851 9895
rect -817 9861 -783 9895
rect -749 9861 -715 9895
rect -681 9861 -647 9895
rect -613 9861 -579 9895
rect -545 9861 -511 9895
rect -477 9861 -443 9895
rect -409 9861 -375 9895
rect -341 9861 -307 9895
rect -273 9861 -266 9895
rect -2966 9826 -266 9861
rect -2966 9792 -2959 9826
rect -2925 9792 -2891 9826
rect -2857 9792 -2823 9826
rect -2789 9792 -2755 9826
rect -2721 9792 -2687 9826
rect -2653 9792 -2619 9826
rect -2585 9792 -2551 9826
rect -2517 9792 -2483 9826
rect -2449 9792 -2415 9826
rect -2381 9792 -2347 9826
rect -2313 9792 -2279 9826
rect -2245 9792 -2211 9826
rect -2177 9792 -2143 9826
rect -2109 9792 -2075 9826
rect -2041 9792 -2007 9826
rect -1973 9792 -1939 9826
rect -1905 9792 -1871 9826
rect -1837 9792 -1803 9826
rect -1769 9792 -1735 9826
rect -1701 9792 -1667 9826
rect -1633 9792 -1599 9826
rect -1565 9792 -1531 9826
rect -1497 9792 -1463 9826
rect -1429 9792 -1395 9826
rect -1361 9792 -1327 9826
rect -1293 9792 -1259 9826
rect -1225 9792 -1191 9826
rect -1157 9792 -1123 9826
rect -1089 9792 -1055 9826
rect -1021 9792 -987 9826
rect -953 9792 -919 9826
rect -885 9792 -851 9826
rect -817 9792 -783 9826
rect -749 9792 -715 9826
rect -681 9792 -647 9826
rect -613 9792 -579 9826
rect -545 9792 -511 9826
rect -477 9792 -443 9826
rect -409 9792 -375 9826
rect -341 9792 -307 9826
rect -273 9792 -266 9826
rect -2966 9757 -266 9792
rect -2966 9723 -2959 9757
rect -2925 9723 -2891 9757
rect -2857 9723 -2823 9757
rect -2789 9723 -2755 9757
rect -2721 9723 -2687 9757
rect -2653 9723 -2619 9757
rect -2585 9723 -2551 9757
rect -2517 9723 -2483 9757
rect -2449 9723 -2415 9757
rect -2381 9723 -2347 9757
rect -2313 9723 -2279 9757
rect -2245 9723 -2211 9757
rect -2177 9723 -2143 9757
rect -2109 9723 -2075 9757
rect -2041 9723 -2007 9757
rect -1973 9723 -1939 9757
rect -1905 9723 -1871 9757
rect -1837 9723 -1803 9757
rect -1769 9723 -1735 9757
rect -1701 9723 -1667 9757
rect -1633 9723 -1599 9757
rect -1565 9723 -1531 9757
rect -1497 9723 -1463 9757
rect -1429 9723 -1395 9757
rect -1361 9723 -1327 9757
rect -1293 9723 -1259 9757
rect -1225 9723 -1191 9757
rect -1157 9723 -1123 9757
rect -1089 9723 -1055 9757
rect -1021 9723 -987 9757
rect -953 9723 -919 9757
rect -885 9723 -851 9757
rect -817 9723 -783 9757
rect -749 9723 -715 9757
rect -681 9723 -647 9757
rect -613 9723 -579 9757
rect -545 9723 -511 9757
rect -477 9723 -443 9757
rect -409 9723 -375 9757
rect -341 9723 -307 9757
rect -273 9723 -266 9757
rect -2966 9688 -266 9723
rect -2966 9654 -2959 9688
rect -2925 9654 -2891 9688
rect -2857 9654 -2823 9688
rect -2789 9654 -2755 9688
rect -2721 9654 -2687 9688
rect -2653 9654 -2619 9688
rect -2585 9654 -2551 9688
rect -2517 9654 -2483 9688
rect -2449 9654 -2415 9688
rect -2381 9654 -2347 9688
rect -2313 9654 -2279 9688
rect -2245 9654 -2211 9688
rect -2177 9654 -2143 9688
rect -2109 9654 -2075 9688
rect -2041 9654 -2007 9688
rect -1973 9654 -1939 9688
rect -1905 9654 -1871 9688
rect -1837 9654 -1803 9688
rect -1769 9654 -1735 9688
rect -1701 9654 -1667 9688
rect -1633 9654 -1599 9688
rect -1565 9654 -1531 9688
rect -1497 9654 -1463 9688
rect -1429 9654 -1395 9688
rect -1361 9654 -1327 9688
rect -1293 9654 -1259 9688
rect -1225 9654 -1191 9688
rect -1157 9654 -1123 9688
rect -1089 9654 -1055 9688
rect -1021 9654 -987 9688
rect -953 9654 -919 9688
rect -885 9654 -851 9688
rect -817 9654 -783 9688
rect -749 9654 -715 9688
rect -681 9654 -647 9688
rect -613 9654 -579 9688
rect -545 9654 -511 9688
rect -477 9654 -443 9688
rect -409 9654 -375 9688
rect -341 9654 -307 9688
rect -273 9654 -266 9688
rect -2966 9619 -266 9654
rect -2966 9585 -2959 9619
rect -2925 9585 -2891 9619
rect -2857 9585 -2823 9619
rect -2789 9585 -2755 9619
rect -2721 9585 -2687 9619
rect -2653 9585 -2619 9619
rect -2585 9585 -2551 9619
rect -2517 9585 -2483 9619
rect -2449 9585 -2415 9619
rect -2381 9585 -2347 9619
rect -2313 9585 -2279 9619
rect -2245 9585 -2211 9619
rect -2177 9585 -2143 9619
rect -2109 9585 -2075 9619
rect -2041 9585 -2007 9619
rect -1973 9585 -1939 9619
rect -1905 9585 -1871 9619
rect -1837 9585 -1803 9619
rect -1769 9585 -1735 9619
rect -1701 9585 -1667 9619
rect -1633 9585 -1599 9619
rect -1565 9585 -1531 9619
rect -1497 9585 -1463 9619
rect -1429 9585 -1395 9619
rect -1361 9585 -1327 9619
rect -1293 9585 -1259 9619
rect -1225 9585 -1191 9619
rect -1157 9585 -1123 9619
rect -1089 9585 -1055 9619
rect -1021 9585 -987 9619
rect -953 9585 -919 9619
rect -885 9585 -851 9619
rect -817 9585 -783 9619
rect -749 9585 -715 9619
rect -681 9585 -647 9619
rect -613 9585 -579 9619
rect -545 9585 -511 9619
rect -477 9585 -443 9619
rect -409 9585 -375 9619
rect -341 9585 -307 9619
rect -273 9585 -266 9619
rect -2966 9550 -266 9585
rect -2966 9516 -2959 9550
rect -2925 9516 -2891 9550
rect -2857 9516 -2823 9550
rect -2789 9516 -2755 9550
rect -2721 9516 -2687 9550
rect -2653 9516 -2619 9550
rect -2585 9516 -2551 9550
rect -2517 9516 -2483 9550
rect -2449 9516 -2415 9550
rect -2381 9516 -2347 9550
rect -2313 9516 -2279 9550
rect -2245 9516 -2211 9550
rect -2177 9516 -2143 9550
rect -2109 9516 -2075 9550
rect -2041 9516 -2007 9550
rect -1973 9516 -1939 9550
rect -1905 9516 -1871 9550
rect -1837 9516 -1803 9550
rect -1769 9516 -1735 9550
rect -1701 9516 -1667 9550
rect -1633 9516 -1599 9550
rect -1565 9516 -1531 9550
rect -1497 9516 -1463 9550
rect -1429 9516 -1395 9550
rect -1361 9516 -1327 9550
rect -1293 9516 -1259 9550
rect -1225 9516 -1191 9550
rect -1157 9516 -1123 9550
rect -1089 9516 -1055 9550
rect -1021 9516 -987 9550
rect -953 9516 -919 9550
rect -885 9516 -851 9550
rect -817 9516 -783 9550
rect -749 9516 -715 9550
rect -681 9516 -647 9550
rect -613 9516 -579 9550
rect -545 9516 -511 9550
rect -477 9516 -443 9550
rect -409 9516 -375 9550
rect -341 9516 -307 9550
rect -273 9516 -266 9550
rect -2966 9481 -266 9516
rect -2966 9447 -2959 9481
rect -2925 9447 -2891 9481
rect -2857 9447 -2823 9481
rect -2789 9447 -2755 9481
rect -2721 9447 -2687 9481
rect -2653 9447 -2619 9481
rect -2585 9447 -2551 9481
rect -2517 9447 -2483 9481
rect -2449 9447 -2415 9481
rect -2381 9447 -2347 9481
rect -2313 9447 -2279 9481
rect -2245 9447 -2211 9481
rect -2177 9447 -2143 9481
rect -2109 9447 -2075 9481
rect -2041 9447 -2007 9481
rect -1973 9447 -1939 9481
rect -1905 9447 -1871 9481
rect -1837 9447 -1803 9481
rect -1769 9447 -1735 9481
rect -1701 9447 -1667 9481
rect -1633 9447 -1599 9481
rect -1565 9447 -1531 9481
rect -1497 9447 -1463 9481
rect -1429 9447 -1395 9481
rect -1361 9447 -1327 9481
rect -1293 9447 -1259 9481
rect -1225 9447 -1191 9481
rect -1157 9447 -1123 9481
rect -1089 9447 -1055 9481
rect -1021 9447 -987 9481
rect -953 9447 -919 9481
rect -885 9447 -851 9481
rect -817 9447 -783 9481
rect -749 9447 -715 9481
rect -681 9447 -647 9481
rect -613 9447 -579 9481
rect -545 9447 -511 9481
rect -477 9447 -443 9481
rect -409 9447 -375 9481
rect -341 9447 -307 9481
rect -273 9447 -266 9481
rect -2966 9412 -266 9447
rect -2966 9378 -2959 9412
rect -2925 9378 -2891 9412
rect -2857 9378 -2823 9412
rect -2789 9378 -2755 9412
rect -2721 9378 -2687 9412
rect -2653 9378 -2619 9412
rect -2585 9378 -2551 9412
rect -2517 9378 -2483 9412
rect -2449 9378 -2415 9412
rect -2381 9378 -2347 9412
rect -2313 9378 -2279 9412
rect -2245 9378 -2211 9412
rect -2177 9378 -2143 9412
rect -2109 9378 -2075 9412
rect -2041 9378 -2007 9412
rect -1973 9378 -1939 9412
rect -1905 9378 -1871 9412
rect -1837 9378 -1803 9412
rect -1769 9378 -1735 9412
rect -1701 9378 -1667 9412
rect -1633 9378 -1599 9412
rect -1565 9378 -1531 9412
rect -1497 9378 -1463 9412
rect -1429 9378 -1395 9412
rect -1361 9378 -1327 9412
rect -1293 9378 -1259 9412
rect -1225 9378 -1191 9412
rect -1157 9378 -1123 9412
rect -1089 9378 -1055 9412
rect -1021 9378 -987 9412
rect -953 9378 -919 9412
rect -885 9378 -851 9412
rect -817 9378 -783 9412
rect -749 9378 -715 9412
rect -681 9378 -647 9412
rect -613 9378 -579 9412
rect -545 9378 -511 9412
rect -477 9378 -443 9412
rect -409 9378 -375 9412
rect -341 9378 -307 9412
rect -273 9378 -266 9412
rect -2966 9343 -266 9378
rect -2966 9309 -2959 9343
rect -2925 9309 -2891 9343
rect -2857 9309 -2823 9343
rect -2789 9309 -2755 9343
rect -2721 9309 -2687 9343
rect -2653 9309 -2619 9343
rect -2585 9309 -2551 9343
rect -2517 9309 -2483 9343
rect -2449 9309 -2415 9343
rect -2381 9309 -2347 9343
rect -2313 9309 -2279 9343
rect -2245 9309 -2211 9343
rect -2177 9309 -2143 9343
rect -2109 9309 -2075 9343
rect -2041 9309 -2007 9343
rect -1973 9309 -1939 9343
rect -1905 9309 -1871 9343
rect -1837 9309 -1803 9343
rect -1769 9309 -1735 9343
rect -1701 9309 -1667 9343
rect -1633 9309 -1599 9343
rect -1565 9309 -1531 9343
rect -1497 9309 -1463 9343
rect -1429 9309 -1395 9343
rect -1361 9309 -1327 9343
rect -1293 9309 -1259 9343
rect -1225 9309 -1191 9343
rect -1157 9309 -1123 9343
rect -1089 9309 -1055 9343
rect -1021 9309 -987 9343
rect -953 9309 -919 9343
rect -885 9309 -851 9343
rect -817 9309 -783 9343
rect -749 9309 -715 9343
rect -681 9309 -647 9343
rect -613 9309 -579 9343
rect -545 9309 -511 9343
rect -477 9309 -443 9343
rect -409 9309 -375 9343
rect -341 9309 -307 9343
rect -273 9309 -266 9343
rect -2966 9274 -266 9309
rect -2966 9240 -2959 9274
rect -2925 9240 -2891 9274
rect -2857 9240 -2823 9274
rect -2789 9240 -2755 9274
rect -2721 9240 -2687 9274
rect -2653 9240 -2619 9274
rect -2585 9240 -2551 9274
rect -2517 9240 -2483 9274
rect -2449 9240 -2415 9274
rect -2381 9240 -2347 9274
rect -2313 9240 -2279 9274
rect -2245 9240 -2211 9274
rect -2177 9240 -2143 9274
rect -2109 9240 -2075 9274
rect -2041 9240 -2007 9274
rect -1973 9240 -1939 9274
rect -1905 9240 -1871 9274
rect -1837 9240 -1803 9274
rect -1769 9240 -1735 9274
rect -1701 9240 -1667 9274
rect -1633 9240 -1599 9274
rect -1565 9240 -1531 9274
rect -1497 9240 -1463 9274
rect -1429 9240 -1395 9274
rect -1361 9240 -1327 9274
rect -1293 9240 -1259 9274
rect -1225 9240 -1191 9274
rect -1157 9240 -1123 9274
rect -1089 9240 -1055 9274
rect -1021 9240 -987 9274
rect -953 9240 -919 9274
rect -885 9240 -851 9274
rect -817 9240 -783 9274
rect -749 9240 -715 9274
rect -681 9240 -647 9274
rect -613 9240 -579 9274
rect -545 9240 -511 9274
rect -477 9240 -443 9274
rect -409 9240 -375 9274
rect -341 9240 -307 9274
rect -273 9240 -266 9274
rect -2966 9205 -266 9240
rect -2966 9171 -2959 9205
rect -2925 9171 -2891 9205
rect -2857 9171 -2823 9205
rect -2789 9171 -2755 9205
rect -2721 9171 -2687 9205
rect -2653 9171 -2619 9205
rect -2585 9171 -2551 9205
rect -2517 9171 -2483 9205
rect -2449 9171 -2415 9205
rect -2381 9171 -2347 9205
rect -2313 9171 -2279 9205
rect -2245 9171 -2211 9205
rect -2177 9171 -2143 9205
rect -2109 9171 -2075 9205
rect -2041 9171 -2007 9205
rect -1973 9171 -1939 9205
rect -1905 9171 -1871 9205
rect -1837 9171 -1803 9205
rect -1769 9171 -1735 9205
rect -1701 9171 -1667 9205
rect -1633 9171 -1599 9205
rect -1565 9171 -1531 9205
rect -1497 9171 -1463 9205
rect -1429 9171 -1395 9205
rect -1361 9171 -1327 9205
rect -1293 9171 -1259 9205
rect -1225 9171 -1191 9205
rect -1157 9171 -1123 9205
rect -1089 9171 -1055 9205
rect -1021 9171 -987 9205
rect -953 9171 -919 9205
rect -885 9171 -851 9205
rect -817 9171 -783 9205
rect -749 9171 -715 9205
rect -681 9171 -647 9205
rect -613 9171 -579 9205
rect -545 9171 -511 9205
rect -477 9171 -443 9205
rect -409 9171 -375 9205
rect -341 9171 -307 9205
rect -273 9171 -266 9205
rect -2966 9136 -266 9171
rect -2966 9102 -2959 9136
rect -2925 9102 -2891 9136
rect -2857 9102 -2823 9136
rect -2789 9102 -2755 9136
rect -2721 9102 -2687 9136
rect -2653 9102 -2619 9136
rect -2585 9102 -2551 9136
rect -2517 9102 -2483 9136
rect -2449 9102 -2415 9136
rect -2381 9102 -2347 9136
rect -2313 9102 -2279 9136
rect -2245 9102 -2211 9136
rect -2177 9102 -2143 9136
rect -2109 9102 -2075 9136
rect -2041 9102 -2007 9136
rect -1973 9102 -1939 9136
rect -1905 9102 -1871 9136
rect -1837 9102 -1803 9136
rect -1769 9102 -1735 9136
rect -1701 9102 -1667 9136
rect -1633 9102 -1599 9136
rect -1565 9102 -1531 9136
rect -1497 9102 -1463 9136
rect -1429 9102 -1395 9136
rect -1361 9102 -1327 9136
rect -1293 9102 -1259 9136
rect -1225 9102 -1191 9136
rect -1157 9102 -1123 9136
rect -1089 9102 -1055 9136
rect -1021 9102 -987 9136
rect -953 9102 -919 9136
rect -885 9102 -851 9136
rect -817 9102 -783 9136
rect -749 9102 -715 9136
rect -681 9102 -647 9136
rect -613 9102 -579 9136
rect -545 9102 -511 9136
rect -477 9102 -443 9136
rect -409 9102 -375 9136
rect -341 9102 -307 9136
rect -273 9102 -266 9136
rect -2966 9067 -266 9102
rect -2966 9033 -2959 9067
rect -2925 9033 -2891 9067
rect -2857 9033 -2823 9067
rect -2789 9033 -2755 9067
rect -2721 9033 -2687 9067
rect -2653 9033 -2619 9067
rect -2585 9033 -2551 9067
rect -2517 9033 -2483 9067
rect -2449 9033 -2415 9067
rect -2381 9033 -2347 9067
rect -2313 9033 -2279 9067
rect -2245 9033 -2211 9067
rect -2177 9033 -2143 9067
rect -2109 9033 -2075 9067
rect -2041 9033 -2007 9067
rect -1973 9033 -1939 9067
rect -1905 9033 -1871 9067
rect -1837 9033 -1803 9067
rect -1769 9033 -1735 9067
rect -1701 9033 -1667 9067
rect -1633 9033 -1599 9067
rect -1565 9033 -1531 9067
rect -1497 9033 -1463 9067
rect -1429 9033 -1395 9067
rect -1361 9033 -1327 9067
rect -1293 9033 -1259 9067
rect -1225 9033 -1191 9067
rect -1157 9033 -1123 9067
rect -1089 9033 -1055 9067
rect -1021 9033 -987 9067
rect -953 9033 -919 9067
rect -885 9033 -851 9067
rect -817 9033 -783 9067
rect -749 9033 -715 9067
rect -681 9033 -647 9067
rect -613 9033 -579 9067
rect -545 9033 -511 9067
rect -477 9033 -443 9067
rect -409 9033 -375 9067
rect -341 9033 -307 9067
rect -273 9033 -266 9067
rect -2966 8998 -266 9033
rect -2966 8964 -2959 8998
rect -2925 8964 -2891 8998
rect -2857 8964 -2823 8998
rect -2789 8964 -2755 8998
rect -2721 8964 -2687 8998
rect -2653 8964 -2619 8998
rect -2585 8964 -2551 8998
rect -2517 8964 -2483 8998
rect -2449 8964 -2415 8998
rect -2381 8964 -2347 8998
rect -2313 8964 -2279 8998
rect -2245 8964 -2211 8998
rect -2177 8964 -2143 8998
rect -2109 8964 -2075 8998
rect -2041 8964 -2007 8998
rect -1973 8964 -1939 8998
rect -1905 8964 -1871 8998
rect -1837 8964 -1803 8998
rect -1769 8964 -1735 8998
rect -1701 8964 -1667 8998
rect -1633 8964 -1599 8998
rect -1565 8964 -1531 8998
rect -1497 8964 -1463 8998
rect -1429 8964 -1395 8998
rect -1361 8964 -1327 8998
rect -1293 8964 -1259 8998
rect -1225 8964 -1191 8998
rect -1157 8964 -1123 8998
rect -1089 8964 -1055 8998
rect -1021 8964 -987 8998
rect -953 8964 -919 8998
rect -885 8964 -851 8998
rect -817 8964 -783 8998
rect -749 8964 -715 8998
rect -681 8964 -647 8998
rect -613 8964 -579 8998
rect -545 8964 -511 8998
rect -477 8964 -443 8998
rect -409 8964 -375 8998
rect -341 8964 -307 8998
rect -273 8964 -266 8998
rect -2966 8929 -266 8964
rect -2966 8895 -2959 8929
rect -2925 8895 -2891 8929
rect -2857 8895 -2823 8929
rect -2789 8895 -2755 8929
rect -2721 8895 -2687 8929
rect -2653 8895 -2619 8929
rect -2585 8895 -2551 8929
rect -2517 8895 -2483 8929
rect -2449 8895 -2415 8929
rect -2381 8895 -2347 8929
rect -2313 8895 -2279 8929
rect -2245 8895 -2211 8929
rect -2177 8895 -2143 8929
rect -2109 8895 -2075 8929
rect -2041 8895 -2007 8929
rect -1973 8895 -1939 8929
rect -1905 8895 -1871 8929
rect -1837 8895 -1803 8929
rect -1769 8895 -1735 8929
rect -1701 8895 -1667 8929
rect -1633 8895 -1599 8929
rect -1565 8895 -1531 8929
rect -1497 8895 -1463 8929
rect -1429 8895 -1395 8929
rect -1361 8895 -1327 8929
rect -1293 8895 -1259 8929
rect -1225 8895 -1191 8929
rect -1157 8895 -1123 8929
rect -1089 8895 -1055 8929
rect -1021 8895 -987 8929
rect -953 8895 -919 8929
rect -885 8895 -851 8929
rect -817 8895 -783 8929
rect -749 8895 -715 8929
rect -681 8895 -647 8929
rect -613 8895 -579 8929
rect -545 8895 -511 8929
rect -477 8895 -443 8929
rect -409 8895 -375 8929
rect -341 8895 -307 8929
rect -273 8895 -266 8929
rect -2966 8860 -266 8895
rect -2966 8826 -2959 8860
rect -2925 8826 -2891 8860
rect -2857 8826 -2823 8860
rect -2789 8826 -2755 8860
rect -2721 8826 -2687 8860
rect -2653 8826 -2619 8860
rect -2585 8826 -2551 8860
rect -2517 8826 -2483 8860
rect -2449 8826 -2415 8860
rect -2381 8826 -2347 8860
rect -2313 8826 -2279 8860
rect -2245 8826 -2211 8860
rect -2177 8826 -2143 8860
rect -2109 8826 -2075 8860
rect -2041 8826 -2007 8860
rect -1973 8826 -1939 8860
rect -1905 8826 -1871 8860
rect -1837 8826 -1803 8860
rect -1769 8826 -1735 8860
rect -1701 8826 -1667 8860
rect -1633 8826 -1599 8860
rect -1565 8826 -1531 8860
rect -1497 8826 -1463 8860
rect -1429 8826 -1395 8860
rect -1361 8826 -1327 8860
rect -1293 8826 -1259 8860
rect -1225 8826 -1191 8860
rect -1157 8826 -1123 8860
rect -1089 8826 -1055 8860
rect -1021 8826 -987 8860
rect -953 8826 -919 8860
rect -885 8826 -851 8860
rect -817 8826 -783 8860
rect -749 8826 -715 8860
rect -681 8826 -647 8860
rect -613 8826 -579 8860
rect -545 8826 -511 8860
rect -477 8826 -443 8860
rect -409 8826 -375 8860
rect -341 8826 -307 8860
rect -273 8826 -266 8860
rect -2966 8791 -266 8826
rect -2966 8757 -2959 8791
rect -2925 8757 -2891 8791
rect -2857 8757 -2823 8791
rect -2789 8757 -2755 8791
rect -2721 8757 -2687 8791
rect -2653 8757 -2619 8791
rect -2585 8757 -2551 8791
rect -2517 8757 -2483 8791
rect -2449 8757 -2415 8791
rect -2381 8757 -2347 8791
rect -2313 8757 -2279 8791
rect -2245 8757 -2211 8791
rect -2177 8757 -2143 8791
rect -2109 8757 -2075 8791
rect -2041 8757 -2007 8791
rect -1973 8757 -1939 8791
rect -1905 8757 -1871 8791
rect -1837 8757 -1803 8791
rect -1769 8757 -1735 8791
rect -1701 8757 -1667 8791
rect -1633 8757 -1599 8791
rect -1565 8757 -1531 8791
rect -1497 8757 -1463 8791
rect -1429 8757 -1395 8791
rect -1361 8757 -1327 8791
rect -1293 8757 -1259 8791
rect -1225 8757 -1191 8791
rect -1157 8757 -1123 8791
rect -1089 8757 -1055 8791
rect -1021 8757 -987 8791
rect -953 8757 -919 8791
rect -885 8757 -851 8791
rect -817 8757 -783 8791
rect -749 8757 -715 8791
rect -681 8757 -647 8791
rect -613 8757 -579 8791
rect -545 8757 -511 8791
rect -477 8757 -443 8791
rect -409 8757 -375 8791
rect -341 8757 -307 8791
rect -273 8757 -266 8791
rect -2966 8722 -266 8757
rect -2966 8688 -2959 8722
rect -2925 8688 -2891 8722
rect -2857 8688 -2823 8722
rect -2789 8688 -2755 8722
rect -2721 8688 -2687 8722
rect -2653 8688 -2619 8722
rect -2585 8688 -2551 8722
rect -2517 8688 -2483 8722
rect -2449 8688 -2415 8722
rect -2381 8688 -2347 8722
rect -2313 8688 -2279 8722
rect -2245 8688 -2211 8722
rect -2177 8688 -2143 8722
rect -2109 8688 -2075 8722
rect -2041 8688 -2007 8722
rect -1973 8688 -1939 8722
rect -1905 8688 -1871 8722
rect -1837 8688 -1803 8722
rect -1769 8688 -1735 8722
rect -1701 8688 -1667 8722
rect -1633 8688 -1599 8722
rect -1565 8688 -1531 8722
rect -1497 8688 -1463 8722
rect -1429 8688 -1395 8722
rect -1361 8688 -1327 8722
rect -1293 8688 -1259 8722
rect -1225 8688 -1191 8722
rect -1157 8688 -1123 8722
rect -1089 8688 -1055 8722
rect -1021 8688 -987 8722
rect -953 8688 -919 8722
rect -885 8688 -851 8722
rect -817 8688 -783 8722
rect -749 8688 -715 8722
rect -681 8688 -647 8722
rect -613 8688 -579 8722
rect -545 8688 -511 8722
rect -477 8688 -443 8722
rect -409 8688 -375 8722
rect -341 8688 -307 8722
rect -273 8688 -266 8722
rect -2966 8653 -266 8688
rect -2966 8619 -2959 8653
rect -2925 8619 -2891 8653
rect -2857 8619 -2823 8653
rect -2789 8619 -2755 8653
rect -2721 8619 -2687 8653
rect -2653 8619 -2619 8653
rect -2585 8619 -2551 8653
rect -2517 8619 -2483 8653
rect -2449 8619 -2415 8653
rect -2381 8619 -2347 8653
rect -2313 8619 -2279 8653
rect -2245 8619 -2211 8653
rect -2177 8619 -2143 8653
rect -2109 8619 -2075 8653
rect -2041 8619 -2007 8653
rect -1973 8619 -1939 8653
rect -1905 8619 -1871 8653
rect -1837 8619 -1803 8653
rect -1769 8619 -1735 8653
rect -1701 8619 -1667 8653
rect -1633 8619 -1599 8653
rect -1565 8619 -1531 8653
rect -1497 8619 -1463 8653
rect -1429 8619 -1395 8653
rect -1361 8619 -1327 8653
rect -1293 8619 -1259 8653
rect -1225 8619 -1191 8653
rect -1157 8619 -1123 8653
rect -1089 8619 -1055 8653
rect -1021 8619 -987 8653
rect -953 8619 -919 8653
rect -885 8619 -851 8653
rect -817 8619 -783 8653
rect -749 8619 -715 8653
rect -681 8619 -647 8653
rect -613 8619 -579 8653
rect -545 8619 -511 8653
rect -477 8619 -443 8653
rect -409 8619 -375 8653
rect -341 8619 -307 8653
rect -273 8619 -266 8653
rect -2966 8584 -266 8619
rect -2966 8550 -2959 8584
rect -2925 8550 -2891 8584
rect -2857 8550 -2823 8584
rect -2789 8550 -2755 8584
rect -2721 8550 -2687 8584
rect -2653 8550 -2619 8584
rect -2585 8550 -2551 8584
rect -2517 8550 -2483 8584
rect -2449 8550 -2415 8584
rect -2381 8550 -2347 8584
rect -2313 8550 -2279 8584
rect -2245 8550 -2211 8584
rect -2177 8550 -2143 8584
rect -2109 8550 -2075 8584
rect -2041 8550 -2007 8584
rect -1973 8550 -1939 8584
rect -1905 8550 -1871 8584
rect -1837 8550 -1803 8584
rect -1769 8550 -1735 8584
rect -1701 8550 -1667 8584
rect -1633 8550 -1599 8584
rect -1565 8550 -1531 8584
rect -1497 8550 -1463 8584
rect -1429 8550 -1395 8584
rect -1361 8550 -1327 8584
rect -1293 8550 -1259 8584
rect -1225 8550 -1191 8584
rect -1157 8550 -1123 8584
rect -1089 8550 -1055 8584
rect -1021 8550 -987 8584
rect -953 8550 -919 8584
rect -885 8550 -851 8584
rect -817 8550 -783 8584
rect -749 8550 -715 8584
rect -681 8550 -647 8584
rect -613 8550 -579 8584
rect -545 8550 -511 8584
rect -477 8550 -443 8584
rect -409 8550 -375 8584
rect -341 8550 -307 8584
rect -273 8550 -266 8584
rect -2966 8515 -266 8550
rect -2966 8481 -2959 8515
rect -2925 8481 -2891 8515
rect -2857 8481 -2823 8515
rect -2789 8481 -2755 8515
rect -2721 8481 -2687 8515
rect -2653 8481 -2619 8515
rect -2585 8481 -2551 8515
rect -2517 8481 -2483 8515
rect -2449 8481 -2415 8515
rect -2381 8481 -2347 8515
rect -2313 8481 -2279 8515
rect -2245 8481 -2211 8515
rect -2177 8481 -2143 8515
rect -2109 8481 -2075 8515
rect -2041 8481 -2007 8515
rect -1973 8481 -1939 8515
rect -1905 8481 -1871 8515
rect -1837 8481 -1803 8515
rect -1769 8481 -1735 8515
rect -1701 8481 -1667 8515
rect -1633 8481 -1599 8515
rect -1565 8481 -1531 8515
rect -1497 8481 -1463 8515
rect -1429 8481 -1395 8515
rect -1361 8481 -1327 8515
rect -1293 8481 -1259 8515
rect -1225 8481 -1191 8515
rect -1157 8481 -1123 8515
rect -1089 8481 -1055 8515
rect -1021 8481 -987 8515
rect -953 8481 -919 8515
rect -885 8481 -851 8515
rect -817 8481 -783 8515
rect -749 8481 -715 8515
rect -681 8481 -647 8515
rect -613 8481 -579 8515
rect -545 8481 -511 8515
rect -477 8481 -443 8515
rect -409 8481 -375 8515
rect -341 8481 -307 8515
rect -273 8481 -266 8515
rect -2966 8446 -266 8481
rect -2966 8412 -2959 8446
rect -2925 8412 -2891 8446
rect -2857 8412 -2823 8446
rect -2789 8412 -2755 8446
rect -2721 8412 -2687 8446
rect -2653 8412 -2619 8446
rect -2585 8412 -2551 8446
rect -2517 8412 -2483 8446
rect -2449 8412 -2415 8446
rect -2381 8412 -2347 8446
rect -2313 8412 -2279 8446
rect -2245 8412 -2211 8446
rect -2177 8412 -2143 8446
rect -2109 8412 -2075 8446
rect -2041 8412 -2007 8446
rect -1973 8412 -1939 8446
rect -1905 8412 -1871 8446
rect -1837 8412 -1803 8446
rect -1769 8412 -1735 8446
rect -1701 8412 -1667 8446
rect -1633 8412 -1599 8446
rect -1565 8412 -1531 8446
rect -1497 8412 -1463 8446
rect -1429 8412 -1395 8446
rect -1361 8412 -1327 8446
rect -1293 8412 -1259 8446
rect -1225 8412 -1191 8446
rect -1157 8412 -1123 8446
rect -1089 8412 -1055 8446
rect -1021 8412 -987 8446
rect -953 8412 -919 8446
rect -885 8412 -851 8446
rect -817 8412 -783 8446
rect -749 8412 -715 8446
rect -681 8412 -647 8446
rect -613 8412 -579 8446
rect -545 8412 -511 8446
rect -477 8412 -443 8446
rect -409 8412 -375 8446
rect -341 8412 -307 8446
rect -273 8412 -266 8446
rect -2966 8377 -266 8412
rect -2966 8343 -2959 8377
rect -2925 8343 -2891 8377
rect -2857 8343 -2823 8377
rect -2789 8343 -2755 8377
rect -2721 8343 -2687 8377
rect -2653 8343 -2619 8377
rect -2585 8343 -2551 8377
rect -2517 8343 -2483 8377
rect -2449 8343 -2415 8377
rect -2381 8343 -2347 8377
rect -2313 8343 -2279 8377
rect -2245 8343 -2211 8377
rect -2177 8343 -2143 8377
rect -2109 8343 -2075 8377
rect -2041 8343 -2007 8377
rect -1973 8343 -1939 8377
rect -1905 8343 -1871 8377
rect -1837 8343 -1803 8377
rect -1769 8343 -1735 8377
rect -1701 8343 -1667 8377
rect -1633 8343 -1599 8377
rect -1565 8343 -1531 8377
rect -1497 8343 -1463 8377
rect -1429 8343 -1395 8377
rect -1361 8343 -1327 8377
rect -1293 8343 -1259 8377
rect -1225 8343 -1191 8377
rect -1157 8343 -1123 8377
rect -1089 8343 -1055 8377
rect -1021 8343 -987 8377
rect -953 8343 -919 8377
rect -885 8343 -851 8377
rect -817 8343 -783 8377
rect -749 8343 -715 8377
rect -681 8343 -647 8377
rect -613 8343 -579 8377
rect -545 8343 -511 8377
rect -477 8343 -443 8377
rect -409 8343 -375 8377
rect -341 8343 -307 8377
rect -273 8343 -266 8377
rect 32028 8348 32061 8542
rect -2966 8308 -266 8343
rect -2966 8274 -2959 8308
rect -2925 8274 -2891 8308
rect -2857 8274 -2823 8308
rect -2789 8274 -2755 8308
rect -2721 8274 -2687 8308
rect -2653 8274 -2619 8308
rect -2585 8274 -2551 8308
rect -2517 8274 -2483 8308
rect -2449 8274 -2415 8308
rect -2381 8274 -2347 8308
rect -2313 8274 -2279 8308
rect -2245 8274 -2211 8308
rect -2177 8274 -2143 8308
rect -2109 8274 -2075 8308
rect -2041 8274 -2007 8308
rect -1973 8274 -1939 8308
rect -1905 8274 -1871 8308
rect -1837 8274 -1803 8308
rect -1769 8274 -1735 8308
rect -1701 8274 -1667 8308
rect -1633 8274 -1599 8308
rect -1565 8274 -1531 8308
rect -1497 8274 -1463 8308
rect -1429 8274 -1395 8308
rect -1361 8274 -1327 8308
rect -1293 8274 -1259 8308
rect -1225 8274 -1191 8308
rect -1157 8274 -1123 8308
rect -1089 8274 -1055 8308
rect -1021 8274 -987 8308
rect -953 8274 -919 8308
rect -885 8274 -851 8308
rect -817 8274 -783 8308
rect -749 8274 -715 8308
rect -681 8274 -647 8308
rect -613 8274 -579 8308
rect -545 8274 -511 8308
rect -477 8274 -443 8308
rect -409 8274 -375 8308
rect -341 8274 -307 8308
rect -273 8274 -266 8308
rect -2966 8239 -266 8274
rect -2966 8205 -2959 8239
rect -2925 8205 -2891 8239
rect -2857 8205 -2823 8239
rect -2789 8205 -2755 8239
rect -2721 8205 -2687 8239
rect -2653 8205 -2619 8239
rect -2585 8205 -2551 8239
rect -2517 8205 -2483 8239
rect -2449 8205 -2415 8239
rect -2381 8205 -2347 8239
rect -2313 8205 -2279 8239
rect -2245 8205 -2211 8239
rect -2177 8205 -2143 8239
rect -2109 8205 -2075 8239
rect -2041 8205 -2007 8239
rect -1973 8205 -1939 8239
rect -1905 8205 -1871 8239
rect -1837 8205 -1803 8239
rect -1769 8205 -1735 8239
rect -1701 8205 -1667 8239
rect -1633 8205 -1599 8239
rect -1565 8205 -1531 8239
rect -1497 8205 -1463 8239
rect -1429 8205 -1395 8239
rect -1361 8205 -1327 8239
rect -1293 8205 -1259 8239
rect -1225 8205 -1191 8239
rect -1157 8205 -1123 8239
rect -1089 8205 -1055 8239
rect -1021 8205 -987 8239
rect -953 8205 -919 8239
rect -885 8205 -851 8239
rect -817 8205 -783 8239
rect -749 8205 -715 8239
rect -681 8205 -647 8239
rect -613 8205 -579 8239
rect -545 8205 -511 8239
rect -477 8205 -443 8239
rect -409 8205 -375 8239
rect -341 8205 -307 8239
rect -273 8205 -266 8239
rect -2966 8170 -266 8205
rect -2966 8136 -2959 8170
rect -2925 8136 -2891 8170
rect -2857 8136 -2823 8170
rect -2789 8136 -2755 8170
rect -2721 8136 -2687 8170
rect -2653 8136 -2619 8170
rect -2585 8136 -2551 8170
rect -2517 8136 -2483 8170
rect -2449 8136 -2415 8170
rect -2381 8136 -2347 8170
rect -2313 8136 -2279 8170
rect -2245 8136 -2211 8170
rect -2177 8136 -2143 8170
rect -2109 8136 -2075 8170
rect -2041 8136 -2007 8170
rect -1973 8136 -1939 8170
rect -1905 8136 -1871 8170
rect -1837 8136 -1803 8170
rect -1769 8136 -1735 8170
rect -1701 8136 -1667 8170
rect -1633 8136 -1599 8170
rect -1565 8136 -1531 8170
rect -1497 8136 -1463 8170
rect -1429 8136 -1395 8170
rect -1361 8136 -1327 8170
rect -1293 8136 -1259 8170
rect -1225 8136 -1191 8170
rect -1157 8136 -1123 8170
rect -1089 8136 -1055 8170
rect -1021 8136 -987 8170
rect -953 8136 -919 8170
rect -885 8136 -851 8170
rect -817 8136 -783 8170
rect -749 8136 -715 8170
rect -681 8136 -647 8170
rect -613 8136 -579 8170
rect -545 8136 -511 8170
rect -477 8136 -443 8170
rect -409 8136 -375 8170
rect -341 8136 -307 8170
rect -273 8136 -266 8170
rect -2966 8101 -266 8136
rect -2966 8067 -2959 8101
rect -2925 8067 -2891 8101
rect -2857 8067 -2823 8101
rect -2789 8067 -2755 8101
rect -2721 8067 -2687 8101
rect -2653 8067 -2619 8101
rect -2585 8067 -2551 8101
rect -2517 8067 -2483 8101
rect -2449 8067 -2415 8101
rect -2381 8067 -2347 8101
rect -2313 8067 -2279 8101
rect -2245 8067 -2211 8101
rect -2177 8067 -2143 8101
rect -2109 8067 -2075 8101
rect -2041 8067 -2007 8101
rect -1973 8067 -1939 8101
rect -1905 8067 -1871 8101
rect -1837 8067 -1803 8101
rect -1769 8067 -1735 8101
rect -1701 8067 -1667 8101
rect -1633 8067 -1599 8101
rect -1565 8067 -1531 8101
rect -1497 8067 -1463 8101
rect -1429 8067 -1395 8101
rect -1361 8067 -1327 8101
rect -1293 8067 -1259 8101
rect -1225 8067 -1191 8101
rect -1157 8067 -1123 8101
rect -1089 8067 -1055 8101
rect -1021 8067 -987 8101
rect -953 8067 -919 8101
rect -885 8067 -851 8101
rect -817 8067 -783 8101
rect -749 8067 -715 8101
rect -681 8067 -647 8101
rect -613 8067 -579 8101
rect -545 8067 -511 8101
rect -477 8067 -443 8101
rect -409 8067 -375 8101
rect -341 8067 -307 8101
rect -273 8067 -266 8101
rect -2966 8032 -266 8067
rect -2966 7998 -2959 8032
rect -2925 7998 -2891 8032
rect -2857 7998 -2823 8032
rect -2789 7998 -2755 8032
rect -2721 7998 -2687 8032
rect -2653 7998 -2619 8032
rect -2585 7998 -2551 8032
rect -2517 7998 -2483 8032
rect -2449 7998 -2415 8032
rect -2381 7998 -2347 8032
rect -2313 7998 -2279 8032
rect -2245 7998 -2211 8032
rect -2177 7998 -2143 8032
rect -2109 7998 -2075 8032
rect -2041 7998 -2007 8032
rect -1973 7998 -1939 8032
rect -1905 7998 -1871 8032
rect -1837 7998 -1803 8032
rect -1769 7998 -1735 8032
rect -1701 7998 -1667 8032
rect -1633 7998 -1599 8032
rect -1565 7998 -1531 8032
rect -1497 7998 -1463 8032
rect -1429 7998 -1395 8032
rect -1361 7998 -1327 8032
rect -1293 7998 -1259 8032
rect -1225 7998 -1191 8032
rect -1157 7998 -1123 8032
rect -1089 7998 -1055 8032
rect -1021 7998 -987 8032
rect -953 7998 -919 8032
rect -885 7998 -851 8032
rect -817 7998 -783 8032
rect -749 7998 -715 8032
rect -681 7998 -647 8032
rect -613 7998 -579 8032
rect -545 7998 -511 8032
rect -477 7998 -443 8032
rect -409 7998 -375 8032
rect -341 7998 -307 8032
rect -273 7998 -266 8032
rect -2966 7963 -266 7998
rect -2966 7929 -2959 7963
rect -2925 7929 -2891 7963
rect -2857 7929 -2823 7963
rect -2789 7929 -2755 7963
rect -2721 7929 -2687 7963
rect -2653 7929 -2619 7963
rect -2585 7929 -2551 7963
rect -2517 7929 -2483 7963
rect -2449 7929 -2415 7963
rect -2381 7929 -2347 7963
rect -2313 7929 -2279 7963
rect -2245 7929 -2211 7963
rect -2177 7929 -2143 7963
rect -2109 7929 -2075 7963
rect -2041 7929 -2007 7963
rect -1973 7929 -1939 7963
rect -1905 7929 -1871 7963
rect -1837 7929 -1803 7963
rect -1769 7929 -1735 7963
rect -1701 7929 -1667 7963
rect -1633 7929 -1599 7963
rect -1565 7929 -1531 7963
rect -1497 7929 -1463 7963
rect -1429 7929 -1395 7963
rect -1361 7929 -1327 7963
rect -1293 7929 -1259 7963
rect -1225 7929 -1191 7963
rect -1157 7929 -1123 7963
rect -1089 7929 -1055 7963
rect -1021 7929 -987 7963
rect -953 7929 -919 7963
rect -885 7929 -851 7963
rect -817 7929 -783 7963
rect -749 7929 -715 7963
rect -681 7929 -647 7963
rect -613 7929 -579 7963
rect -545 7929 -511 7963
rect -477 7929 -443 7963
rect -409 7929 -375 7963
rect -341 7929 -307 7963
rect -273 7929 -266 7963
rect -2966 7894 -266 7929
rect -2966 7860 -2959 7894
rect -2925 7860 -2891 7894
rect -2857 7860 -2823 7894
rect -2789 7860 -2755 7894
rect -2721 7860 -2687 7894
rect -2653 7860 -2619 7894
rect -2585 7860 -2551 7894
rect -2517 7860 -2483 7894
rect -2449 7860 -2415 7894
rect -2381 7860 -2347 7894
rect -2313 7860 -2279 7894
rect -2245 7860 -2211 7894
rect -2177 7860 -2143 7894
rect -2109 7860 -2075 7894
rect -2041 7860 -2007 7894
rect -1973 7860 -1939 7894
rect -1905 7860 -1871 7894
rect -1837 7860 -1803 7894
rect -1769 7860 -1735 7894
rect -1701 7860 -1667 7894
rect -1633 7860 -1599 7894
rect -1565 7860 -1531 7894
rect -1497 7860 -1463 7894
rect -1429 7860 -1395 7894
rect -1361 7860 -1327 7894
rect -1293 7860 -1259 7894
rect -1225 7860 -1191 7894
rect -1157 7860 -1123 7894
rect -1089 7860 -1055 7894
rect -1021 7860 -987 7894
rect -953 7860 -919 7894
rect -885 7860 -851 7894
rect -817 7860 -783 7894
rect -749 7860 -715 7894
rect -681 7860 -647 7894
rect -613 7860 -579 7894
rect -545 7860 -511 7894
rect -477 7860 -443 7894
rect -409 7860 -375 7894
rect -341 7860 -307 7894
rect -273 7860 -266 7894
rect -2966 7825 -266 7860
rect -2966 7791 -2959 7825
rect -2925 7791 -2891 7825
rect -2857 7791 -2823 7825
rect -2789 7791 -2755 7825
rect -2721 7791 -2687 7825
rect -2653 7791 -2619 7825
rect -2585 7791 -2551 7825
rect -2517 7791 -2483 7825
rect -2449 7791 -2415 7825
rect -2381 7791 -2347 7825
rect -2313 7791 -2279 7825
rect -2245 7791 -2211 7825
rect -2177 7791 -2143 7825
rect -2109 7791 -2075 7825
rect -2041 7791 -2007 7825
rect -1973 7791 -1939 7825
rect -1905 7791 -1871 7825
rect -1837 7791 -1803 7825
rect -1769 7791 -1735 7825
rect -1701 7791 -1667 7825
rect -1633 7791 -1599 7825
rect -1565 7791 -1531 7825
rect -1497 7791 -1463 7825
rect -1429 7791 -1395 7825
rect -1361 7791 -1327 7825
rect -1293 7791 -1259 7825
rect -1225 7791 -1191 7825
rect -1157 7791 -1123 7825
rect -1089 7791 -1055 7825
rect -1021 7791 -987 7825
rect -953 7791 -919 7825
rect -885 7791 -851 7825
rect -817 7791 -783 7825
rect -749 7791 -715 7825
rect -681 7791 -647 7825
rect -613 7791 -579 7825
rect -545 7791 -511 7825
rect -477 7791 -443 7825
rect -409 7791 -375 7825
rect -341 7791 -307 7825
rect -273 7791 -266 7825
rect -2966 7756 -266 7791
rect -2966 7722 -2959 7756
rect -2925 7722 -2891 7756
rect -2857 7722 -2823 7756
rect -2789 7722 -2755 7756
rect -2721 7722 -2687 7756
rect -2653 7722 -2619 7756
rect -2585 7722 -2551 7756
rect -2517 7722 -2483 7756
rect -2449 7722 -2415 7756
rect -2381 7722 -2347 7756
rect -2313 7722 -2279 7756
rect -2245 7722 -2211 7756
rect -2177 7722 -2143 7756
rect -2109 7722 -2075 7756
rect -2041 7722 -2007 7756
rect -1973 7722 -1939 7756
rect -1905 7722 -1871 7756
rect -1837 7722 -1803 7756
rect -1769 7722 -1735 7756
rect -1701 7722 -1667 7756
rect -1633 7722 -1599 7756
rect -1565 7722 -1531 7756
rect -1497 7722 -1463 7756
rect -1429 7722 -1395 7756
rect -1361 7722 -1327 7756
rect -1293 7722 -1259 7756
rect -1225 7722 -1191 7756
rect -1157 7722 -1123 7756
rect -1089 7722 -1055 7756
rect -1021 7722 -987 7756
rect -953 7722 -919 7756
rect -885 7722 -851 7756
rect -817 7722 -783 7756
rect -749 7722 -715 7756
rect -681 7722 -647 7756
rect -613 7722 -579 7756
rect -545 7722 -511 7756
rect -477 7722 -443 7756
rect -409 7722 -375 7756
rect -341 7722 -307 7756
rect -273 7722 -266 7756
rect -2966 7687 -266 7722
rect -2966 7653 -2959 7687
rect -2925 7653 -2891 7687
rect -2857 7653 -2823 7687
rect -2789 7653 -2755 7687
rect -2721 7653 -2687 7687
rect -2653 7653 -2619 7687
rect -2585 7653 -2551 7687
rect -2517 7653 -2483 7687
rect -2449 7653 -2415 7687
rect -2381 7653 -2347 7687
rect -2313 7653 -2279 7687
rect -2245 7653 -2211 7687
rect -2177 7653 -2143 7687
rect -2109 7653 -2075 7687
rect -2041 7653 -2007 7687
rect -1973 7653 -1939 7687
rect -1905 7653 -1871 7687
rect -1837 7653 -1803 7687
rect -1769 7653 -1735 7687
rect -1701 7653 -1667 7687
rect -1633 7653 -1599 7687
rect -1565 7653 -1531 7687
rect -1497 7653 -1463 7687
rect -1429 7653 -1395 7687
rect -1361 7653 -1327 7687
rect -1293 7653 -1259 7687
rect -1225 7653 -1191 7687
rect -1157 7653 -1123 7687
rect -1089 7653 -1055 7687
rect -1021 7653 -987 7687
rect -953 7653 -919 7687
rect -885 7653 -851 7687
rect -817 7653 -783 7687
rect -749 7653 -715 7687
rect -681 7653 -647 7687
rect -613 7653 -579 7687
rect -545 7653 -511 7687
rect -477 7653 -443 7687
rect -409 7653 -375 7687
rect -341 7653 -307 7687
rect -273 7653 -266 7687
rect -2966 7618 -266 7653
rect -2966 7584 -2959 7618
rect -2925 7584 -2891 7618
rect -2857 7584 -2823 7618
rect -2789 7584 -2755 7618
rect -2721 7584 -2687 7618
rect -2653 7584 -2619 7618
rect -2585 7584 -2551 7618
rect -2517 7584 -2483 7618
rect -2449 7584 -2415 7618
rect -2381 7584 -2347 7618
rect -2313 7584 -2279 7618
rect -2245 7584 -2211 7618
rect -2177 7584 -2143 7618
rect -2109 7584 -2075 7618
rect -2041 7584 -2007 7618
rect -1973 7584 -1939 7618
rect -1905 7584 -1871 7618
rect -1837 7584 -1803 7618
rect -1769 7584 -1735 7618
rect -1701 7584 -1667 7618
rect -1633 7584 -1599 7618
rect -1565 7584 -1531 7618
rect -1497 7584 -1463 7618
rect -1429 7584 -1395 7618
rect -1361 7584 -1327 7618
rect -1293 7584 -1259 7618
rect -1225 7584 -1191 7618
rect -1157 7584 -1123 7618
rect -1089 7584 -1055 7618
rect -1021 7584 -987 7618
rect -953 7584 -919 7618
rect -885 7584 -851 7618
rect -817 7584 -783 7618
rect -749 7584 -715 7618
rect -681 7584 -647 7618
rect -613 7584 -579 7618
rect -545 7584 -511 7618
rect -477 7584 -443 7618
rect -409 7584 -375 7618
rect -341 7584 -307 7618
rect -273 7584 -266 7618
rect -2966 7549 -266 7584
rect -2966 7515 -2959 7549
rect -2925 7515 -2891 7549
rect -2857 7515 -2823 7549
rect -2789 7515 -2755 7549
rect -2721 7515 -2687 7549
rect -2653 7515 -2619 7549
rect -2585 7515 -2551 7549
rect -2517 7515 -2483 7549
rect -2449 7515 -2415 7549
rect -2381 7515 -2347 7549
rect -2313 7515 -2279 7549
rect -2245 7515 -2211 7549
rect -2177 7515 -2143 7549
rect -2109 7515 -2075 7549
rect -2041 7515 -2007 7549
rect -1973 7515 -1939 7549
rect -1905 7515 -1871 7549
rect -1837 7515 -1803 7549
rect -1769 7515 -1735 7549
rect -1701 7515 -1667 7549
rect -1633 7515 -1599 7549
rect -1565 7515 -1531 7549
rect -1497 7515 -1463 7549
rect -1429 7515 -1395 7549
rect -1361 7515 -1327 7549
rect -1293 7515 -1259 7549
rect -1225 7515 -1191 7549
rect -1157 7515 -1123 7549
rect -1089 7515 -1055 7549
rect -1021 7515 -987 7549
rect -953 7515 -919 7549
rect -885 7515 -851 7549
rect -817 7515 -783 7549
rect -749 7515 -715 7549
rect -681 7515 -647 7549
rect -613 7515 -579 7549
rect -545 7515 -511 7549
rect -477 7515 -443 7549
rect -409 7515 -375 7549
rect -341 7515 -307 7549
rect -273 7515 -266 7549
rect -2966 7480 -266 7515
rect -2966 7446 -2959 7480
rect -2925 7446 -2891 7480
rect -2857 7446 -2823 7480
rect -2789 7446 -2755 7480
rect -2721 7446 -2687 7480
rect -2653 7446 -2619 7480
rect -2585 7446 -2551 7480
rect -2517 7446 -2483 7480
rect -2449 7446 -2415 7480
rect -2381 7446 -2347 7480
rect -2313 7446 -2279 7480
rect -2245 7446 -2211 7480
rect -2177 7446 -2143 7480
rect -2109 7446 -2075 7480
rect -2041 7446 -2007 7480
rect -1973 7446 -1939 7480
rect -1905 7446 -1871 7480
rect -1837 7446 -1803 7480
rect -1769 7446 -1735 7480
rect -1701 7446 -1667 7480
rect -1633 7446 -1599 7480
rect -1565 7446 -1531 7480
rect -1497 7446 -1463 7480
rect -1429 7446 -1395 7480
rect -1361 7446 -1327 7480
rect -1293 7446 -1259 7480
rect -1225 7446 -1191 7480
rect -1157 7446 -1123 7480
rect -1089 7446 -1055 7480
rect -1021 7446 -987 7480
rect -953 7446 -919 7480
rect -885 7446 -851 7480
rect -817 7446 -783 7480
rect -749 7446 -715 7480
rect -681 7446 -647 7480
rect -613 7446 -579 7480
rect -545 7446 -511 7480
rect -477 7446 -443 7480
rect -409 7446 -375 7480
rect -341 7446 -307 7480
rect -273 7446 -266 7480
rect -2966 7422 -266 7446
<< mvnsubdiff >>
rect 14 50636 228 50677
rect 14 50602 15 50636
rect 49 50632 228 50636
rect 49 50602 87 50632
rect 14 50598 87 50602
rect 121 50627 228 50632
rect 121 50598 159 50627
rect 14 50593 159 50598
rect 193 50593 228 50627
rect 14 50568 228 50593
rect 14 50534 15 50568
rect 49 50564 228 50568
rect 49 50534 87 50564
rect 14 50530 87 50534
rect 121 50559 228 50564
rect 121 50530 159 50559
rect 14 50525 159 50530
rect 193 50525 228 50559
rect 14 50500 228 50525
rect 14 50466 15 50500
rect 49 50496 228 50500
rect 49 50466 87 50496
rect 14 50462 87 50466
rect 121 50491 228 50496
rect 121 50462 159 50491
rect 14 50457 159 50462
rect 193 50457 228 50491
rect 14 50432 228 50457
rect 14 50398 15 50432
rect 49 50428 228 50432
rect 49 50398 87 50428
rect 14 50394 87 50398
rect 121 50423 228 50428
rect 121 50394 159 50423
rect 14 50389 159 50394
rect 193 50389 228 50423
rect 14 50364 228 50389
rect 14 50330 15 50364
rect 49 50360 228 50364
rect 49 50330 87 50360
rect 14 50326 87 50330
rect 121 50355 228 50360
rect 121 50326 159 50355
rect 14 50321 159 50326
rect 193 50321 228 50355
rect 14 50296 228 50321
rect 14 50262 15 50296
rect 49 50292 228 50296
rect 49 50262 87 50292
rect 14 50258 87 50262
rect 121 50287 228 50292
rect 121 50258 159 50287
rect 14 50253 159 50258
rect 193 50253 228 50287
rect 14 50228 228 50253
rect 14 50194 15 50228
rect 49 50224 228 50228
rect 49 50194 87 50224
rect 14 50190 87 50194
rect 121 50219 228 50224
rect 121 50190 159 50219
rect 14 50185 159 50190
rect 193 50185 228 50219
rect 14 50160 228 50185
rect 14 50126 15 50160
rect 49 50156 228 50160
rect 49 50126 87 50156
rect 14 50122 87 50126
rect 121 50151 228 50156
rect 121 50122 159 50151
rect 14 50117 159 50122
rect 193 50117 228 50151
rect 14 50092 228 50117
rect 14 50058 15 50092
rect 49 50088 228 50092
rect 49 50058 87 50088
rect 14 50054 87 50058
rect 121 50083 228 50088
rect 121 50054 159 50083
rect 14 50049 159 50054
rect 193 50049 228 50083
rect 14 50024 228 50049
rect 14 49990 15 50024
rect 49 50020 228 50024
rect 49 49990 87 50020
rect 14 49986 87 49990
rect 121 50015 228 50020
rect 121 49986 159 50015
rect 14 49981 159 49986
rect 193 49981 228 50015
rect 14 49956 228 49981
rect 14 49922 15 49956
rect 49 49952 228 49956
rect 49 49922 87 49952
rect 14 49918 87 49922
rect 121 49947 228 49952
rect 121 49918 159 49947
rect 14 49913 159 49918
rect 193 49913 228 49947
rect 14 49888 228 49913
rect 14 49854 15 49888
rect 49 49884 228 49888
rect 49 49854 87 49884
rect 14 49850 87 49854
rect 121 49879 228 49884
rect 121 49850 159 49879
rect 14 49845 159 49850
rect 193 49845 228 49879
rect 14 49820 228 49845
rect 14 49786 15 49820
rect 49 49816 228 49820
rect 49 49786 87 49816
rect 14 49782 87 49786
rect 121 49811 228 49816
rect 121 49782 159 49811
rect 14 49777 159 49782
rect 193 49777 228 49811
rect 14 49752 228 49777
rect 14 49718 15 49752
rect 49 49748 228 49752
rect 49 49718 87 49748
rect 14 49714 87 49718
rect 121 49743 228 49748
rect 121 49714 159 49743
rect 14 49709 159 49714
rect 193 49709 228 49743
rect 14 49684 228 49709
rect 14 49650 15 49684
rect 49 49680 228 49684
rect 49 49650 87 49680
rect 14 49646 87 49650
rect 121 49675 228 49680
rect 121 49646 159 49675
rect 14 49641 159 49646
rect 193 49641 228 49675
rect 14 49616 228 49641
rect 14 49582 15 49616
rect 49 49612 228 49616
rect 49 49582 87 49612
rect 14 49578 87 49582
rect 121 49607 228 49612
rect 121 49578 159 49607
rect 14 49573 159 49578
rect 193 49573 228 49607
rect 14 49548 228 49573
rect 14 49514 15 49548
rect 49 49544 228 49548
rect 49 49514 87 49544
rect 14 49510 87 49514
rect 121 49539 228 49544
rect 121 49510 159 49539
rect 14 49505 159 49510
rect 193 49505 228 49539
rect 14 49480 228 49505
rect 14 49446 15 49480
rect 49 49476 228 49480
rect 49 49446 87 49476
rect 14 49442 87 49446
rect 121 49471 228 49476
rect 121 49442 159 49471
rect 14 49437 159 49442
rect 193 49437 228 49471
rect 14 49412 228 49437
rect 14 49378 15 49412
rect 49 49408 228 49412
rect 49 49378 87 49408
rect 14 49374 87 49378
rect 121 49403 228 49408
rect 121 49374 159 49403
rect 14 49369 159 49374
rect 193 49369 228 49403
rect 14 49344 228 49369
rect 14 49310 15 49344
rect 49 49340 228 49344
rect 49 49310 87 49340
rect 14 49306 87 49310
rect 121 49335 228 49340
rect 121 49306 159 49335
rect 14 49301 159 49306
rect 193 49301 228 49335
rect 14 49276 228 49301
rect 14 49242 15 49276
rect 49 49272 228 49276
rect 49 49242 87 49272
rect 14 49238 87 49242
rect 121 49267 228 49272
rect 121 49238 159 49267
rect 14 49233 159 49238
rect 193 49233 228 49267
rect 14 49208 228 49233
rect 14 49174 15 49208
rect 49 49204 228 49208
rect 49 49174 87 49204
rect 14 49170 87 49174
rect 121 49199 228 49204
rect 121 49170 159 49199
rect 14 49165 159 49170
rect 193 49165 228 49199
rect 14 49140 228 49165
rect 14 49106 15 49140
rect 49 49136 228 49140
rect 49 49106 87 49136
rect 14 49102 87 49106
rect 121 49131 228 49136
rect 121 49102 159 49131
rect 14 49097 159 49102
rect 193 49097 228 49131
rect 14 49072 228 49097
rect 14 49038 15 49072
rect 49 49068 228 49072
rect 49 49038 87 49068
rect 14 49034 87 49038
rect 121 49063 228 49068
rect 121 49034 159 49063
rect 14 49029 159 49034
rect 193 49029 228 49063
rect 14 49004 228 49029
rect 14 48970 15 49004
rect 49 49000 228 49004
rect 49 48970 87 49000
rect 14 48966 87 48970
rect 121 48995 228 49000
rect 121 48966 159 48995
rect 14 48961 159 48966
rect 193 48961 228 48995
rect 14 48936 228 48961
rect 14 48902 15 48936
rect 49 48932 228 48936
rect 49 48902 87 48932
rect 14 48898 87 48902
rect 121 48927 228 48932
rect 121 48898 159 48927
rect 14 48893 159 48898
rect 193 48893 228 48927
rect 14 48868 228 48893
rect 14 48834 15 48868
rect 49 48864 228 48868
rect 49 48834 87 48864
rect 14 48830 87 48834
rect 121 48859 228 48864
rect 121 48830 159 48859
rect 14 48825 159 48830
rect 193 48825 228 48859
rect 14 48800 228 48825
rect 14 48766 15 48800
rect 49 48796 228 48800
rect 49 48766 87 48796
rect 14 48762 87 48766
rect 121 48791 228 48796
rect 121 48762 159 48791
rect 14 48757 159 48762
rect 193 48757 228 48791
rect 14 48732 228 48757
rect 14 48698 15 48732
rect 49 48728 228 48732
rect 49 48698 87 48728
rect 14 48694 87 48698
rect 121 48723 228 48728
rect 121 48694 159 48723
rect 14 48689 159 48694
rect 193 48689 228 48723
rect 14 48664 228 48689
rect 14 48630 15 48664
rect 49 48660 228 48664
rect 49 48630 87 48660
rect 14 48626 87 48630
rect 121 48655 228 48660
rect 121 48626 159 48655
rect 14 48621 159 48626
rect 193 48621 228 48655
rect 14 48596 228 48621
rect 14 48562 15 48596
rect 49 48592 228 48596
rect 49 48562 87 48592
rect 14 48558 87 48562
rect 121 48587 228 48592
rect 121 48558 159 48587
rect 14 48553 159 48558
rect 193 48553 228 48587
rect 14 48528 228 48553
rect 14 48494 15 48528
rect 49 48524 228 48528
rect 49 48494 87 48524
rect 14 48490 87 48494
rect 121 48519 228 48524
rect 121 48490 159 48519
rect 14 48485 159 48490
rect 193 48485 228 48519
rect 14 48460 228 48485
rect 14 48426 15 48460
rect 49 48456 228 48460
rect 49 48426 87 48456
rect 14 48422 87 48426
rect 121 48451 228 48456
rect 121 48422 159 48451
rect 14 48417 159 48422
rect 193 48417 228 48451
rect 14 48392 228 48417
rect 14 48358 15 48392
rect 49 48388 228 48392
rect 49 48358 87 48388
rect 14 48354 87 48358
rect 121 48383 228 48388
rect 121 48354 159 48383
rect 14 48349 159 48354
rect 193 48349 228 48383
rect 14 48324 228 48349
rect 14 48290 15 48324
rect 49 48320 228 48324
rect 49 48290 87 48320
rect 14 48286 87 48290
rect 121 48315 228 48320
rect 121 48286 159 48315
rect 14 48281 159 48286
rect 193 48281 228 48315
rect 14 48256 228 48281
rect 14 48222 15 48256
rect 49 48252 228 48256
rect 49 48222 87 48252
rect 14 48218 87 48222
rect 121 48247 228 48252
rect 121 48218 159 48247
rect 14 48213 159 48218
rect 193 48213 228 48247
rect 14 48188 228 48213
rect 14 48154 15 48188
rect 49 48184 228 48188
rect 49 48154 87 48184
rect 14 48150 87 48154
rect 121 48179 228 48184
rect 121 48150 159 48179
rect 14 48145 159 48150
rect 193 48145 228 48179
rect 14 48120 228 48145
rect 14 48086 15 48120
rect 49 48116 228 48120
rect 49 48086 87 48116
rect 14 48082 87 48086
rect 121 48111 228 48116
rect 121 48082 159 48111
rect 14 48077 159 48082
rect 193 48077 228 48111
rect 14 48052 228 48077
rect 14 48018 15 48052
rect 49 48048 228 48052
rect 49 48018 87 48048
rect 14 48014 87 48018
rect 121 48043 228 48048
rect 121 48014 159 48043
rect 14 48009 159 48014
rect 193 48009 228 48043
rect 14 47984 228 48009
rect 14 47950 15 47984
rect 49 47980 228 47984
rect 49 47950 87 47980
rect 14 47946 87 47950
rect 121 47975 228 47980
rect 121 47946 159 47975
rect 14 47941 159 47946
rect 193 47941 228 47975
rect 14 47916 228 47941
rect 14 47882 15 47916
rect 49 47912 228 47916
rect 49 47882 87 47912
rect 14 47878 87 47882
rect 121 47907 228 47912
rect 121 47878 159 47907
rect 14 47873 159 47878
rect 193 47873 228 47907
rect 14 47848 228 47873
rect 14 47814 15 47848
rect 49 47844 228 47848
rect 49 47814 87 47844
rect 14 47810 87 47814
rect 121 47839 228 47844
rect 121 47810 159 47839
rect 14 47805 159 47810
rect 193 47805 228 47839
rect 14 47780 228 47805
rect 14 47746 15 47780
rect 49 47776 228 47780
rect 49 47746 87 47776
rect 14 47742 87 47746
rect 121 47771 228 47776
rect 121 47742 159 47771
rect 14 47737 159 47742
rect 193 47737 228 47771
rect 14 47712 228 47737
rect 14 47678 15 47712
rect 49 47708 228 47712
rect 49 47678 87 47708
rect 14 47674 87 47678
rect 121 47703 228 47708
rect 121 47674 159 47703
rect 14 47669 159 47674
rect 193 47669 228 47703
rect 14 47644 228 47669
rect 14 47610 15 47644
rect 49 47640 228 47644
rect 49 47610 87 47640
rect 14 47606 87 47610
rect 121 47635 228 47640
rect 121 47606 159 47635
rect 14 47601 159 47606
rect 193 47601 228 47635
rect 14 47576 228 47601
rect 14 47542 15 47576
rect 49 47572 228 47576
rect 49 47542 87 47572
rect 14 47538 87 47542
rect 121 47567 228 47572
rect 121 47538 159 47567
rect 14 47533 159 47538
rect 193 47533 228 47567
rect 14 47508 228 47533
rect 14 47474 15 47508
rect 49 47504 228 47508
rect 49 47474 87 47504
rect 14 47470 87 47474
rect 121 47499 228 47504
rect 121 47470 159 47499
rect 14 47465 159 47470
rect 193 47465 228 47499
rect 14 47440 228 47465
rect 14 47406 15 47440
rect 49 47436 228 47440
rect 49 47406 87 47436
rect 14 47402 87 47406
rect 121 47431 228 47436
rect 121 47402 159 47431
rect 14 47397 159 47402
rect 193 47397 228 47431
rect 14 47372 228 47397
rect 14 47338 15 47372
rect 49 47368 228 47372
rect 49 47338 87 47368
rect 14 47334 87 47338
rect 121 47363 228 47368
rect 121 47334 159 47363
rect 14 47329 159 47334
rect 193 47329 228 47363
rect 14 47304 228 47329
rect 14 47270 15 47304
rect 49 47300 228 47304
rect 49 47270 87 47300
rect 14 47266 87 47270
rect 121 47295 228 47300
rect 121 47266 159 47295
rect 14 47261 159 47266
rect 193 47261 228 47295
rect 14 47236 228 47261
rect 14 47202 15 47236
rect 49 47232 228 47236
rect 49 47202 87 47232
rect 14 47198 87 47202
rect 121 47227 228 47232
rect 121 47198 159 47227
rect 14 47193 159 47198
rect 193 47193 228 47227
rect 14 47168 228 47193
rect 14 47134 15 47168
rect 49 47164 228 47168
rect 49 47134 87 47164
rect 14 47130 87 47134
rect 121 47159 228 47164
rect 121 47130 159 47159
rect 14 47125 159 47130
rect 193 47125 228 47159
rect 14 47100 228 47125
rect 14 47066 15 47100
rect 49 47096 228 47100
rect 49 47066 87 47096
rect 14 47062 87 47066
rect 121 47091 228 47096
rect 121 47062 159 47091
rect 14 47057 159 47062
rect 193 47057 228 47091
rect 14 47032 228 47057
rect 14 46998 15 47032
rect 49 47028 228 47032
rect 49 46998 87 47028
rect 14 46994 87 46998
rect 121 47023 228 47028
rect 121 46994 159 47023
rect 14 46989 159 46994
rect 193 46989 228 47023
rect 14 46964 228 46989
rect 14 46930 15 46964
rect 49 46960 228 46964
rect 49 46930 87 46960
rect 14 46926 87 46930
rect 121 46955 228 46960
rect 121 46926 159 46955
rect 14 46921 159 46926
rect 193 46921 228 46955
rect 14 46896 228 46921
rect 14 46862 15 46896
rect 49 46892 228 46896
rect 49 46862 87 46892
rect 14 46858 87 46862
rect 121 46887 228 46892
rect 121 46858 159 46887
rect 14 46853 159 46858
rect 193 46853 228 46887
rect 14 46828 228 46853
rect 14 46794 15 46828
rect 49 46824 228 46828
rect 49 46794 87 46824
rect 14 46790 87 46794
rect 121 46819 228 46824
rect 121 46790 159 46819
rect 14 46785 159 46790
rect 193 46785 228 46819
rect 14 46760 228 46785
rect 14 46726 15 46760
rect 49 46756 228 46760
rect 49 46726 87 46756
rect 14 46722 87 46726
rect 121 46751 228 46756
rect 121 46722 159 46751
rect 14 46717 159 46722
rect 193 46717 228 46751
rect 14 46692 228 46717
rect 14 46658 15 46692
rect 49 46688 228 46692
rect 49 46658 87 46688
rect 14 46654 87 46658
rect 121 46683 228 46688
rect 121 46654 159 46683
rect 14 46649 159 46654
rect 193 46649 228 46683
rect 14 46624 228 46649
rect 14 46590 15 46624
rect 49 46620 228 46624
rect 49 46590 87 46620
rect 14 46586 87 46590
rect 121 46615 228 46620
rect 121 46586 159 46615
rect 14 46581 159 46586
rect 193 46581 228 46615
rect 14 46556 228 46581
rect 14 46522 15 46556
rect 49 46552 228 46556
rect 49 46522 87 46552
rect 14 46518 87 46522
rect 121 46547 228 46552
rect 121 46518 159 46547
rect 14 46513 159 46518
rect 193 46513 228 46547
rect 14 46488 228 46513
rect 14 46454 15 46488
rect 49 46484 228 46488
rect 49 46454 87 46484
rect 14 46450 87 46454
rect 121 46479 228 46484
rect 121 46450 159 46479
rect 14 46445 159 46450
rect 193 46445 228 46479
rect 14 46420 228 46445
rect 14 46386 15 46420
rect 49 46416 228 46420
rect 49 46386 87 46416
rect 14 46382 87 46386
rect 121 46411 228 46416
rect 121 46382 159 46411
rect 14 46377 159 46382
rect 193 46377 228 46411
rect 14 46352 228 46377
rect 14 46318 15 46352
rect 49 46348 228 46352
rect 49 46318 87 46348
rect 14 46314 87 46318
rect 121 46343 228 46348
rect 121 46314 159 46343
rect 14 46309 159 46314
rect 193 46309 228 46343
rect 14 46284 228 46309
rect 14 46250 15 46284
rect 49 46280 228 46284
rect 49 46250 87 46280
rect 14 46246 87 46250
rect 121 46275 228 46280
rect 121 46246 159 46275
rect 14 46241 159 46246
rect 193 46241 228 46275
rect 14 46216 228 46241
rect 14 46182 15 46216
rect 49 46212 228 46216
rect 49 46182 87 46212
rect 14 46178 87 46182
rect 121 46207 228 46212
rect 121 46178 159 46207
rect 14 46173 159 46178
rect 193 46173 228 46207
rect 14 46148 228 46173
rect 14 46114 15 46148
rect 49 46144 228 46148
rect 49 46114 87 46144
rect 14 46110 87 46114
rect 121 46139 228 46144
rect 121 46110 159 46139
rect 14 46105 159 46110
rect 193 46105 228 46139
rect 14 46080 228 46105
rect 14 46046 15 46080
rect 49 46076 228 46080
rect 49 46046 87 46076
rect 14 46042 87 46046
rect 121 46071 228 46076
rect 121 46042 159 46071
rect 14 46037 159 46042
rect 193 46037 228 46071
rect 14 46012 228 46037
rect 14 45978 15 46012
rect 49 46008 228 46012
rect 49 45978 87 46008
rect 14 45974 87 45978
rect 121 46003 228 46008
rect 121 45974 159 46003
rect 14 45969 159 45974
rect 193 45969 228 46003
rect 14 45944 228 45969
rect 14 45910 15 45944
rect 49 45940 228 45944
rect 49 45910 87 45940
rect 14 45906 87 45910
rect 121 45935 228 45940
rect 121 45906 159 45935
rect 14 45901 159 45906
rect 193 45901 228 45935
rect 14 45876 228 45901
rect 14 45842 15 45876
rect 49 45872 228 45876
rect 49 45842 87 45872
rect 14 45838 87 45842
rect 121 45867 228 45872
rect 121 45838 159 45867
rect 14 45833 159 45838
rect 193 45833 228 45867
rect 14 45808 228 45833
rect 14 45774 15 45808
rect 49 45804 228 45808
rect 49 45774 87 45804
rect 14 45770 87 45774
rect 121 45799 228 45804
rect 121 45770 159 45799
rect 14 45765 159 45770
rect 193 45765 228 45799
rect 14 45740 228 45765
rect 14 45706 15 45740
rect 49 45736 228 45740
rect 49 45706 87 45736
rect 14 45702 87 45706
rect 121 45731 228 45736
rect 121 45702 159 45731
rect 14 45697 159 45702
rect 193 45697 228 45731
rect 14 45672 228 45697
rect 14 45638 15 45672
rect 49 45668 228 45672
rect 49 45638 87 45668
rect 14 45634 87 45638
rect 121 45663 228 45668
rect 121 45634 159 45663
rect 14 45629 159 45634
rect 193 45629 228 45663
rect 14 45604 228 45629
rect 14 45570 15 45604
rect 49 45600 228 45604
rect 49 45570 87 45600
rect 14 45566 87 45570
rect 121 45595 228 45600
rect 121 45566 159 45595
rect 14 45561 159 45566
rect 193 45561 228 45595
rect 14 45536 228 45561
rect 14 45502 15 45536
rect 49 45532 228 45536
rect 49 45502 87 45532
rect 14 45498 87 45502
rect 121 45527 228 45532
rect 121 45498 159 45527
rect 14 45493 159 45498
rect 193 45493 228 45527
rect 14 45468 228 45493
rect 14 45434 15 45468
rect 49 45464 228 45468
rect 49 45434 87 45464
rect 14 45430 87 45434
rect 121 45459 228 45464
rect 121 45430 159 45459
rect 14 45425 159 45430
rect 193 45425 228 45459
rect 14 45400 228 45425
rect 14 45366 15 45400
rect 49 45396 228 45400
rect 49 45366 87 45396
rect 14 45362 87 45366
rect 121 45391 228 45396
rect 121 45362 159 45391
rect 14 45357 159 45362
rect 193 45357 228 45391
rect 14 45332 228 45357
rect 14 45298 15 45332
rect 49 45328 228 45332
rect 49 45298 87 45328
rect 14 45294 87 45298
rect 121 45323 228 45328
rect 121 45294 159 45323
rect 14 45289 159 45294
rect 193 45289 228 45323
rect 14 45264 228 45289
rect 14 45230 15 45264
rect 49 45260 228 45264
rect 49 45230 87 45260
rect 14 45226 87 45230
rect 121 45255 228 45260
rect 121 45226 159 45255
rect 14 45221 159 45226
rect 193 45221 228 45255
rect 14 45196 228 45221
rect 14 45162 15 45196
rect 49 45192 228 45196
rect 49 45162 87 45192
rect 14 45158 87 45162
rect 121 45187 228 45192
rect 121 45158 159 45187
rect 14 45153 159 45158
rect 193 45153 228 45187
rect 14 45128 228 45153
rect 14 45094 15 45128
rect 49 45124 228 45128
rect 49 45094 87 45124
rect 14 45090 87 45094
rect 121 45119 228 45124
rect 121 45090 159 45119
rect 14 45085 159 45090
rect 193 45085 228 45119
rect 14 45060 228 45085
rect 14 45026 15 45060
rect 49 45056 228 45060
rect 49 45026 87 45056
rect 14 45022 87 45026
rect 121 45051 228 45056
rect 121 45022 159 45051
rect 14 45017 159 45022
rect 193 45017 228 45051
rect 14 44992 228 45017
rect 14 44958 15 44992
rect 49 44988 228 44992
rect 49 44958 87 44988
rect 14 44954 87 44958
rect 121 44983 228 44988
rect 121 44954 159 44983
rect 14 44949 159 44954
rect 193 44949 228 44983
rect 14 44924 228 44949
rect 14 44890 15 44924
rect 49 44920 228 44924
rect 49 44890 87 44920
rect 14 44886 87 44890
rect 121 44915 228 44920
rect 121 44886 159 44915
rect 14 44881 159 44886
rect 193 44881 228 44915
rect 14 44856 228 44881
rect 14 44822 15 44856
rect 49 44852 228 44856
rect 49 44822 87 44852
rect 14 44818 87 44822
rect 121 44847 228 44852
rect 121 44818 159 44847
rect 14 44813 159 44818
rect 193 44813 228 44847
rect 14 44788 228 44813
rect 14 44754 15 44788
rect 49 44784 228 44788
rect 49 44754 87 44784
rect 14 44750 87 44754
rect 121 44779 228 44784
rect 121 44750 159 44779
rect 14 44745 159 44750
rect 193 44745 228 44779
rect 14 44720 228 44745
rect 14 44686 15 44720
rect 49 44716 228 44720
rect 49 44686 87 44716
rect 14 44682 87 44686
rect 121 44711 228 44716
rect 121 44682 159 44711
rect 14 44677 159 44682
rect 193 44677 228 44711
rect 14 44652 228 44677
rect 14 44618 15 44652
rect 49 44648 228 44652
rect 49 44618 87 44648
rect 14 44614 87 44618
rect 121 44643 228 44648
rect 121 44614 159 44643
rect 14 44609 159 44614
rect 193 44609 228 44643
rect 14 44584 228 44609
rect 14 44550 15 44584
rect 49 44580 228 44584
rect 49 44550 87 44580
rect 14 44546 87 44550
rect 121 44575 228 44580
rect 121 44546 159 44575
rect 14 44541 159 44546
rect 193 44541 228 44575
rect 14 44516 228 44541
rect 14 44482 15 44516
rect 49 44512 228 44516
rect 49 44482 87 44512
rect 14 44478 87 44482
rect 121 44507 228 44512
rect 121 44478 159 44507
rect 14 44473 159 44478
rect 193 44473 228 44507
rect 14 44448 228 44473
rect 14 44414 15 44448
rect 49 44444 228 44448
rect 49 44414 87 44444
rect 14 44410 87 44414
rect 121 44439 228 44444
rect 121 44410 159 44439
rect 14 44405 159 44410
rect 193 44405 228 44439
rect 14 44380 228 44405
rect 14 44346 15 44380
rect 49 44376 228 44380
rect 49 44346 87 44376
rect 14 44342 87 44346
rect 121 44371 228 44376
rect 121 44342 159 44371
rect 14 44337 159 44342
rect 193 44337 228 44371
rect 14 44312 228 44337
rect 14 44278 15 44312
rect 49 44308 228 44312
rect 49 44278 87 44308
rect 14 44274 87 44278
rect 121 44303 228 44308
rect 121 44274 159 44303
rect 14 44269 159 44274
rect 193 44269 228 44303
rect 14 44244 228 44269
rect 14 44210 15 44244
rect 49 44240 228 44244
rect 49 44210 87 44240
rect 14 44206 87 44210
rect 121 44235 228 44240
rect 121 44206 159 44235
rect 14 44201 159 44206
rect 193 44201 228 44235
rect 14 44176 228 44201
rect 14 44142 15 44176
rect 49 44172 228 44176
rect 49 44142 87 44172
rect 14 44138 87 44142
rect 121 44167 228 44172
rect 121 44138 159 44167
rect 14 44133 159 44138
rect 193 44133 228 44167
rect 14 44108 228 44133
rect 14 44074 15 44108
rect 49 44104 228 44108
rect 49 44074 87 44104
rect 14 44070 87 44074
rect 121 44099 228 44104
rect 121 44070 159 44099
rect 14 44065 159 44070
rect 193 44065 228 44099
rect 14 44040 228 44065
rect 14 44006 15 44040
rect 49 44036 228 44040
rect 49 44006 87 44036
rect 14 44002 87 44006
rect 121 44031 228 44036
rect 121 44002 159 44031
rect 14 43997 159 44002
rect 193 43997 228 44031
rect 14 43972 228 43997
rect 14 43938 15 43972
rect 49 43968 228 43972
rect 49 43938 87 43968
rect 14 43934 87 43938
rect 121 43963 228 43968
rect 121 43934 159 43963
rect 14 43929 159 43934
rect 193 43929 228 43963
rect 14 43904 228 43929
rect 14 43870 15 43904
rect 49 43900 228 43904
rect 49 43870 87 43900
rect 14 43866 87 43870
rect 121 43895 228 43900
rect 121 43866 159 43895
rect 14 43861 159 43866
rect 193 43861 228 43895
rect 14 43836 228 43861
rect 14 43802 15 43836
rect 49 43832 228 43836
rect 49 43802 87 43832
rect 14 43798 87 43802
rect 121 43827 228 43832
rect 121 43798 159 43827
rect 14 43793 159 43798
rect 193 43793 228 43827
rect 14 43768 228 43793
rect 14 43734 15 43768
rect 49 43764 228 43768
rect 49 43734 87 43764
rect 14 43730 87 43734
rect 121 43759 228 43764
rect 121 43730 159 43759
rect 14 43725 159 43730
rect 193 43725 228 43759
rect 14 43700 228 43725
rect 14 43666 15 43700
rect 49 43696 228 43700
rect 49 43666 87 43696
rect 14 43662 87 43666
rect 121 43691 228 43696
rect 121 43662 159 43691
rect 14 43657 159 43662
rect 193 43657 228 43691
rect 14 43632 228 43657
rect 14 43598 15 43632
rect 49 43628 228 43632
rect 49 43598 87 43628
rect 14 43594 87 43598
rect 121 43623 228 43628
rect 121 43594 159 43623
rect 14 43589 159 43594
rect 193 43589 228 43623
rect 14 43564 228 43589
rect 14 43530 15 43564
rect 49 43560 228 43564
rect 49 43530 87 43560
rect 14 43526 87 43530
rect 121 43555 228 43560
rect 121 43526 159 43555
rect 14 43521 159 43526
rect 193 43521 228 43555
rect 14 43496 228 43521
rect 14 43462 15 43496
rect 49 43492 228 43496
rect 49 43462 87 43492
rect 14 43458 87 43462
rect 121 43487 228 43492
rect 121 43458 159 43487
rect 14 43453 159 43458
rect 193 43453 228 43487
rect 14 43428 228 43453
rect 14 43394 15 43428
rect 49 43424 228 43428
rect 49 43394 87 43424
rect 14 43390 87 43394
rect 121 43419 228 43424
rect 121 43390 159 43419
rect 14 43385 159 43390
rect 193 43385 228 43419
rect 14 43360 228 43385
rect 14 43326 15 43360
rect 49 43356 228 43360
rect 49 43326 87 43356
rect 14 43322 87 43326
rect 121 43351 228 43356
rect 121 43322 159 43351
rect 14 43317 159 43322
rect 193 43317 228 43351
rect 14 43292 228 43317
rect 14 43258 15 43292
rect 49 43288 228 43292
rect 49 43258 87 43288
rect 14 43254 87 43258
rect 121 43283 228 43288
rect 121 43254 159 43283
rect 14 43249 159 43254
rect 193 43249 228 43283
rect 14 43224 228 43249
rect 14 43190 15 43224
rect 49 43220 228 43224
rect 49 43190 87 43220
rect 14 43186 87 43190
rect 121 43215 228 43220
rect 121 43186 159 43215
rect 14 43181 159 43186
rect 193 43181 228 43215
rect 14 43156 228 43181
rect 14 43122 15 43156
rect 49 43152 228 43156
rect 49 43122 87 43152
rect 14 43118 87 43122
rect 121 43147 228 43152
rect 121 43118 159 43147
rect 14 43113 159 43118
rect 193 43113 228 43147
rect 14 43088 228 43113
rect 14 43054 15 43088
rect 49 43084 228 43088
rect 49 43054 87 43084
rect 14 43050 87 43054
rect 121 43079 228 43084
rect 121 43050 159 43079
rect 14 43045 159 43050
rect 193 43045 228 43079
rect 14 43020 228 43045
rect 14 42986 15 43020
rect 49 43016 228 43020
rect 49 42986 87 43016
rect 14 42982 87 42986
rect 121 43011 228 43016
rect 121 42982 159 43011
rect 14 42977 159 42982
rect 193 42977 228 43011
rect 14 42952 228 42977
rect 14 42918 15 42952
rect 49 42948 228 42952
rect 49 42918 87 42948
rect 14 42914 87 42918
rect 121 42943 228 42948
rect 121 42914 159 42943
rect 14 42909 159 42914
rect 193 42909 228 42943
rect 14 42884 228 42909
rect 14 42850 15 42884
rect 49 42880 228 42884
rect 49 42850 87 42880
rect 14 42846 87 42850
rect 121 42875 228 42880
rect 121 42846 159 42875
rect 14 42841 159 42846
rect 193 42841 228 42875
rect 14 42816 228 42841
rect 14 42782 15 42816
rect 49 42812 228 42816
rect 49 42782 87 42812
rect 14 42778 87 42782
rect 121 42807 228 42812
rect 121 42778 159 42807
rect 14 42773 159 42778
rect 193 42773 228 42807
rect 14 42748 228 42773
rect 14 42714 15 42748
rect 49 42744 228 42748
rect 49 42714 87 42744
rect 14 42710 87 42714
rect 121 42739 228 42744
rect 121 42710 159 42739
rect 14 42705 159 42710
rect 193 42705 228 42739
rect 14 42680 228 42705
rect 14 42646 15 42680
rect 49 42676 228 42680
rect 49 42646 87 42676
rect 14 42642 87 42646
rect 121 42671 228 42676
rect 121 42642 159 42671
rect 14 42637 159 42642
rect 193 42637 228 42671
rect 14 42612 228 42637
rect 14 42578 15 42612
rect 49 42608 228 42612
rect 49 42578 87 42608
rect 14 42574 87 42578
rect 121 42603 228 42608
rect 121 42574 159 42603
rect 14 42569 159 42574
rect 193 42569 228 42603
rect 14 42544 228 42569
rect 14 42510 15 42544
rect 49 42540 228 42544
rect 49 42510 87 42540
rect 14 42506 87 42510
rect 121 42535 228 42540
rect 121 42506 159 42535
rect 14 42501 159 42506
rect 193 42501 228 42535
rect 14 42476 228 42501
rect 14 42442 15 42476
rect 49 42472 228 42476
rect 49 42442 87 42472
rect 14 42438 87 42442
rect 121 42467 228 42472
rect 121 42438 159 42467
rect 14 42433 159 42438
rect 193 42433 228 42467
rect 14 42408 228 42433
rect 14 42374 15 42408
rect 49 42404 228 42408
rect 49 42374 87 42404
rect 14 42370 87 42374
rect 121 42399 228 42404
rect 121 42370 159 42399
rect 14 42365 159 42370
rect 193 42365 228 42399
rect 14 42340 228 42365
rect 14 42306 15 42340
rect 49 42336 228 42340
rect 49 42306 87 42336
rect 14 42302 87 42306
rect 121 42331 228 42336
rect 121 42302 159 42331
rect 14 42297 159 42302
rect 193 42297 228 42331
rect 14 42272 228 42297
rect 14 42238 15 42272
rect 49 42268 228 42272
rect 49 42238 87 42268
rect 14 42234 87 42238
rect 121 42263 228 42268
rect 121 42234 159 42263
rect 14 42229 159 42234
rect 193 42229 228 42263
rect 14 42204 228 42229
rect 14 42170 15 42204
rect 49 42200 228 42204
rect 49 42170 87 42200
rect 14 42166 87 42170
rect 121 42195 228 42200
rect 121 42166 159 42195
rect 14 42161 159 42166
rect 193 42161 228 42195
rect 14 42136 228 42161
rect 14 42102 15 42136
rect 49 42132 228 42136
rect 49 42102 87 42132
rect 14 42098 87 42102
rect 121 42127 228 42132
rect 121 42098 159 42127
rect 14 42093 159 42098
rect 193 42093 228 42127
rect 14 42068 228 42093
rect 14 42034 15 42068
rect 49 42064 228 42068
rect 49 42034 87 42064
rect 14 42030 87 42034
rect 121 42059 228 42064
rect 121 42030 159 42059
rect 14 42025 159 42030
rect 193 42025 228 42059
rect 14 42000 228 42025
rect 14 41966 15 42000
rect 49 41996 228 42000
rect 49 41966 87 41996
rect 14 41962 87 41966
rect 121 41991 228 41996
rect 121 41962 159 41991
rect 14 41957 159 41962
rect 193 41957 228 41991
rect 14 41932 228 41957
rect 14 41898 15 41932
rect 49 41928 228 41932
rect 49 41898 87 41928
rect 14 41894 87 41898
rect 121 41923 228 41928
rect 121 41894 159 41923
rect 14 41889 159 41894
rect 193 41889 228 41923
rect 14 41864 228 41889
rect 14 41830 15 41864
rect 49 41860 228 41864
rect 49 41830 87 41860
rect 14 41826 87 41830
rect 121 41855 228 41860
rect 121 41826 159 41855
rect 14 41821 159 41826
rect 193 41821 228 41855
rect 14 41796 228 41821
rect 14 41762 15 41796
rect 49 41792 228 41796
rect 49 41762 87 41792
rect 14 41758 87 41762
rect 121 41787 228 41792
rect 121 41758 159 41787
rect 14 41753 159 41758
rect 193 41753 228 41787
rect 14 41728 228 41753
rect 14 41694 15 41728
rect 49 41724 228 41728
rect 49 41694 87 41724
rect 14 41690 87 41694
rect 121 41719 228 41724
rect 121 41690 159 41719
rect 14 41685 159 41690
rect 193 41685 228 41719
rect 14 41660 228 41685
rect 14 41626 15 41660
rect 49 41656 228 41660
rect 49 41626 87 41656
rect 14 41622 87 41626
rect 121 41651 228 41656
rect 121 41622 159 41651
rect 14 41617 159 41622
rect 193 41617 228 41651
rect 14 41592 228 41617
rect 14 41558 15 41592
rect 49 41588 228 41592
rect 49 41558 87 41588
rect 14 41554 87 41558
rect 121 41583 228 41588
rect 121 41554 159 41583
rect 14 41549 159 41554
rect 193 41549 228 41583
rect 14 41524 228 41549
rect 14 41490 15 41524
rect 49 41520 228 41524
rect 49 41490 87 41520
rect 14 41486 87 41490
rect 121 41515 228 41520
rect 121 41486 159 41515
rect 14 41481 159 41486
rect 193 41481 228 41515
rect 14 41456 228 41481
rect 14 41422 15 41456
rect 49 41452 228 41456
rect 49 41422 87 41452
rect 14 41418 87 41422
rect 121 41447 228 41452
rect 121 41418 159 41447
rect 14 41413 159 41418
rect 193 41413 228 41447
rect 14 41388 228 41413
rect 14 41354 15 41388
rect 49 41384 228 41388
rect 49 41354 87 41384
rect 14 41350 87 41354
rect 121 41379 228 41384
rect 121 41350 159 41379
rect 14 41345 159 41350
rect 193 41345 228 41379
rect 14 41320 228 41345
rect 14 41286 15 41320
rect 49 41316 228 41320
rect 49 41286 87 41316
rect 14 41282 87 41286
rect 121 41311 228 41316
rect 121 41282 159 41311
rect 14 41277 159 41282
rect 193 41277 228 41311
rect 14 41252 228 41277
rect 14 41218 15 41252
rect 49 41248 228 41252
rect 49 41218 87 41248
rect 14 41214 87 41218
rect 121 41243 228 41248
rect 121 41214 159 41243
rect 14 41209 159 41214
rect 193 41209 228 41243
rect 14 41184 228 41209
rect 14 41150 15 41184
rect 49 41180 228 41184
rect 49 41150 87 41180
rect 14 41146 87 41150
rect 121 41175 228 41180
rect 121 41146 159 41175
rect 14 41141 159 41146
rect 193 41141 228 41175
rect 14 41116 228 41141
rect 14 41082 15 41116
rect 49 41112 228 41116
rect 49 41082 87 41112
rect 14 41078 87 41082
rect 121 41107 228 41112
rect 121 41078 159 41107
rect 14 41073 159 41078
rect 193 41073 228 41107
rect 14 41048 228 41073
rect 14 41014 15 41048
rect 49 41044 228 41048
rect 49 41014 87 41044
rect 14 41010 87 41014
rect 121 41039 228 41044
rect 121 41010 159 41039
rect 14 41005 159 41010
rect 193 41005 228 41039
rect 14 40980 228 41005
rect 14 40946 15 40980
rect 49 40976 228 40980
rect 49 40946 87 40976
rect 14 40942 87 40946
rect 121 40971 228 40976
rect 121 40942 159 40971
rect 14 40937 159 40942
rect 193 40937 228 40971
rect 14 40912 228 40937
rect 14 40878 15 40912
rect 49 40908 228 40912
rect 49 40878 87 40908
rect 14 40874 87 40878
rect 121 40903 228 40908
rect 121 40874 159 40903
rect 14 40869 159 40874
rect 193 40869 228 40903
rect 14 40844 228 40869
rect 14 40810 15 40844
rect 49 40840 228 40844
rect 49 40810 87 40840
rect 14 40806 87 40810
rect 121 40835 228 40840
rect 121 40806 159 40835
rect 14 40801 159 40806
rect 193 40801 228 40835
rect 14 40776 228 40801
rect 14 40742 15 40776
rect 49 40772 228 40776
rect 49 40742 87 40772
rect 14 40738 87 40742
rect 121 40767 228 40772
rect 121 40738 159 40767
rect 14 40733 159 40738
rect 193 40733 228 40767
rect 14 40708 228 40733
rect 14 40674 15 40708
rect 49 40704 228 40708
rect 49 40674 87 40704
rect 14 40670 87 40674
rect 121 40699 228 40704
rect 121 40670 159 40699
rect 14 40665 159 40670
rect 193 40665 228 40699
rect 14 40640 228 40665
rect 14 40606 15 40640
rect 49 40636 228 40640
rect 49 40606 87 40636
rect 14 40602 87 40606
rect 121 40631 228 40636
rect 121 40602 159 40631
rect 14 40597 159 40602
rect 193 40597 228 40631
rect 14 40572 228 40597
rect 14 40538 15 40572
rect 49 40568 228 40572
rect 49 40538 87 40568
rect 14 40534 87 40538
rect 121 40563 228 40568
rect 121 40534 159 40563
rect 14 40529 159 40534
rect 193 40529 228 40563
rect 14 40504 228 40529
rect 14 40470 15 40504
rect 49 40500 228 40504
rect 49 40470 87 40500
rect 14 40466 87 40470
rect 121 40495 228 40500
rect 121 40466 159 40495
rect 14 40461 159 40466
rect 193 40461 228 40495
rect 14 40436 228 40461
rect 14 40402 15 40436
rect 49 40432 228 40436
rect 49 40402 87 40432
rect 14 40398 87 40402
rect 121 40427 228 40432
rect 121 40398 159 40427
rect 14 40393 159 40398
rect 193 40393 228 40427
rect 14 40368 228 40393
rect 14 40334 15 40368
rect 49 40364 228 40368
rect 49 40334 87 40364
rect 14 40330 87 40334
rect 121 40359 228 40364
rect 121 40330 159 40359
rect 14 40325 159 40330
rect 193 40325 228 40359
rect 14 40300 228 40325
rect 14 40266 15 40300
rect 49 40296 228 40300
rect 49 40266 87 40296
rect 14 40262 87 40266
rect 121 40291 228 40296
rect 121 40262 159 40291
rect 14 40257 159 40262
rect 193 40257 228 40291
rect 14 40232 228 40257
rect 14 40198 15 40232
rect 49 40228 228 40232
rect 49 40198 87 40228
rect 14 40194 87 40198
rect 121 40223 228 40228
rect 121 40194 159 40223
rect 14 40189 159 40194
rect 193 40189 228 40223
rect 14 40164 228 40189
rect 14 40130 15 40164
rect 49 40160 228 40164
rect 49 40130 87 40160
rect 14 40126 87 40130
rect 121 40155 228 40160
rect 121 40126 159 40155
rect 14 40121 159 40126
rect 193 40121 228 40155
rect 14 40096 228 40121
rect 14 40062 15 40096
rect 49 40092 228 40096
rect 49 40062 87 40092
rect 14 40058 87 40062
rect 121 40087 228 40092
rect 121 40058 159 40087
rect 14 40053 159 40058
rect 193 40053 228 40087
rect 14 40028 228 40053
rect 14 39994 15 40028
rect 49 40024 228 40028
rect 49 39994 87 40024
rect 14 39990 87 39994
rect 121 40019 228 40024
rect 121 39990 159 40019
rect 14 39985 159 39990
rect 193 39985 228 40019
rect 14 39960 228 39985
rect 14 39926 15 39960
rect 49 39956 228 39960
rect 49 39926 87 39956
rect 14 39922 87 39926
rect 121 39951 228 39956
rect 121 39922 159 39951
rect 14 39917 159 39922
rect 193 39917 228 39951
rect 14 39892 228 39917
rect 14 39858 15 39892
rect 49 39888 228 39892
rect 49 39858 87 39888
rect 14 39854 87 39858
rect 121 39883 228 39888
rect 121 39854 159 39883
rect 14 39849 159 39854
rect 193 39849 228 39883
rect 14 39824 228 39849
rect 14 39790 15 39824
rect 49 39820 228 39824
rect 49 39790 87 39820
rect 14 39786 87 39790
rect 121 39815 228 39820
rect 121 39786 159 39815
rect 14 39781 159 39786
rect 193 39781 228 39815
rect 14 39756 228 39781
rect 14 39722 15 39756
rect 49 39752 228 39756
rect 49 39722 87 39752
rect 14 39718 87 39722
rect 121 39747 228 39752
rect 121 39718 159 39747
rect 14 39713 159 39718
rect 193 39713 228 39747
rect 14 39688 228 39713
rect 14 39654 15 39688
rect 49 39684 228 39688
rect 49 39654 87 39684
rect 14 39650 87 39654
rect 121 39679 228 39684
rect 121 39650 159 39679
rect 14 39645 159 39650
rect 193 39645 228 39679
rect 14 39620 228 39645
rect 14 39586 15 39620
rect 49 39616 228 39620
rect 49 39586 87 39616
rect 14 39582 87 39586
rect 121 39611 228 39616
rect 121 39582 159 39611
rect 14 39577 159 39582
rect 193 39577 228 39611
rect 14 39552 228 39577
rect 14 39518 15 39552
rect 49 39548 228 39552
rect 49 39518 87 39548
rect 14 39514 87 39518
rect 121 39543 228 39548
rect 121 39514 159 39543
rect 14 39509 159 39514
rect 193 39509 228 39543
rect 14 39484 228 39509
rect 14 39450 15 39484
rect 49 39480 228 39484
rect 49 39450 87 39480
rect 14 39446 87 39450
rect 121 39475 228 39480
rect 121 39446 159 39475
rect 14 39441 159 39446
rect 193 39441 228 39475
rect 14 39416 228 39441
rect 14 39382 15 39416
rect 49 39412 228 39416
rect 49 39382 87 39412
rect 14 39378 87 39382
rect 121 39407 228 39412
rect 121 39378 159 39407
rect 14 39373 159 39378
rect 193 39373 228 39407
rect 14 39348 228 39373
rect 14 39314 15 39348
rect 49 39344 228 39348
rect 49 39314 87 39344
rect 14 39310 87 39314
rect 121 39339 228 39344
rect 121 39310 159 39339
rect 14 39305 159 39310
rect 193 39305 228 39339
rect 14 39280 228 39305
rect 14 39246 15 39280
rect 49 39276 228 39280
rect 49 39246 87 39276
rect 14 39242 87 39246
rect 121 39271 228 39276
rect 121 39242 159 39271
rect 14 39237 159 39242
rect 193 39237 228 39271
rect 14 39212 228 39237
rect 14 39178 15 39212
rect 49 39208 228 39212
rect 49 39178 87 39208
rect 14 39174 87 39178
rect 121 39203 228 39208
rect 121 39174 159 39203
rect 14 39169 159 39174
rect 193 39169 228 39203
rect 14 39144 228 39169
rect 14 39110 15 39144
rect 49 39140 228 39144
rect 49 39110 87 39140
rect 14 39106 87 39110
rect 121 39135 228 39140
rect 121 39106 159 39135
rect 14 39101 159 39106
rect 193 39101 228 39135
rect 14 39076 228 39101
rect 14 39042 15 39076
rect 49 39072 228 39076
rect 49 39042 87 39072
rect 14 39038 87 39042
rect 121 39067 228 39072
rect 121 39038 159 39067
rect 14 39033 159 39038
rect 193 39033 228 39067
rect 14 39008 228 39033
rect 14 38974 15 39008
rect 49 39004 228 39008
rect 49 38974 87 39004
rect 14 38970 87 38974
rect 121 38999 228 39004
rect 121 38970 159 38999
rect 14 38965 159 38970
rect 193 38965 228 38999
rect 14 38940 228 38965
rect 14 38906 15 38940
rect 49 38936 228 38940
rect 49 38906 87 38936
rect 14 38902 87 38906
rect 121 38931 228 38936
rect 121 38902 159 38931
rect 14 38897 159 38902
rect 193 38897 228 38931
rect 14 38872 228 38897
rect 14 38838 15 38872
rect 49 38868 228 38872
rect 49 38838 87 38868
rect 14 38834 87 38838
rect 121 38863 228 38868
rect 121 38834 159 38863
rect 14 38829 159 38834
rect 193 38861 228 38863
rect 193 38829 194 38861
rect 14 38804 194 38829
rect 14 38770 15 38804
rect 49 38800 194 38804
rect 49 38770 87 38800
rect 14 38766 87 38770
rect 121 38795 194 38800
rect 121 38766 159 38795
rect 14 38761 159 38766
rect 193 38761 194 38795
rect 14 38736 194 38761
rect 14 38702 15 38736
rect 49 38732 194 38736
rect 49 38702 87 38732
rect 14 38698 87 38702
rect 121 38727 194 38732
rect 121 38698 159 38727
rect 14 38693 159 38698
rect 193 38693 194 38727
rect 14 38668 194 38693
rect 14 38634 15 38668
rect 49 38664 194 38668
rect 49 38634 87 38664
rect 14 38630 87 38634
rect 121 38659 194 38664
rect 121 38630 159 38659
rect 14 38625 159 38630
rect 193 38625 194 38659
rect 14 38600 194 38625
rect 14 38566 15 38600
rect 49 38596 194 38600
rect 49 38566 87 38596
rect 14 38562 87 38566
rect 121 38591 194 38596
rect 121 38562 159 38591
rect 14 38557 159 38562
rect 193 38557 194 38591
rect 14 38532 194 38557
rect 14 38498 15 38532
rect 49 38528 194 38532
rect 49 38498 87 38528
rect 14 38494 87 38498
rect 121 38523 194 38528
rect 121 38494 159 38523
rect 14 38489 159 38494
rect 193 38489 194 38523
rect 14 38464 194 38489
rect 14 38430 15 38464
rect 49 38460 194 38464
rect 49 38430 87 38460
rect 14 38426 87 38430
rect 121 38455 194 38460
rect 121 38426 159 38455
rect 14 38421 159 38426
rect 193 38421 194 38455
rect 14 38396 194 38421
rect 14 38362 15 38396
rect 49 38392 194 38396
rect 49 38362 87 38392
rect 14 38358 87 38362
rect 121 38387 194 38392
rect 121 38358 159 38387
rect 14 38353 159 38358
rect 193 38353 194 38387
rect 14 38328 194 38353
rect 14 38294 15 38328
rect 49 38324 194 38328
rect 49 38294 87 38324
rect 14 38290 87 38294
rect 121 38319 194 38324
rect 121 38290 159 38319
rect 14 38285 159 38290
rect 193 38285 194 38319
rect 14 38260 194 38285
rect 14 38226 15 38260
rect 49 38256 194 38260
rect 49 38226 87 38256
rect 14 38222 87 38226
rect 121 38251 194 38256
rect 121 38222 159 38251
rect 14 38217 159 38222
rect 193 38217 194 38251
rect 14 38192 194 38217
rect 14 38158 15 38192
rect 49 38188 194 38192
rect 49 38158 87 38188
rect 14 38154 87 38158
rect 121 38183 194 38188
rect 121 38154 159 38183
rect 14 38149 159 38154
rect 193 38149 194 38183
rect 14 38124 194 38149
rect 14 38090 15 38124
rect 49 38120 194 38124
rect 49 38090 87 38120
rect 14 38086 87 38090
rect 121 38115 194 38120
rect 121 38086 159 38115
rect 14 38081 159 38086
rect 193 38081 194 38115
rect 14 38056 194 38081
rect 14 38022 15 38056
rect 49 38052 194 38056
rect 49 38022 87 38052
rect 14 38018 87 38022
rect 121 38047 194 38052
rect 121 38018 159 38047
rect 14 38013 159 38018
rect 193 38013 194 38047
rect 14 37988 194 38013
rect 14 37954 15 37988
rect 49 37984 194 37988
rect 49 37954 87 37984
rect 14 37950 87 37954
rect 121 37979 194 37984
rect 121 37950 159 37979
rect 14 37945 159 37950
rect 193 37945 194 37979
rect 14 37920 194 37945
rect 14 37886 15 37920
rect 49 37916 194 37920
rect 49 37886 87 37916
rect 14 37882 87 37886
rect 121 37911 194 37916
rect 121 37882 159 37911
rect 14 37877 159 37882
rect 193 37877 194 37911
rect 14 37852 194 37877
rect 14 37818 15 37852
rect 49 37848 194 37852
rect 49 37818 87 37848
rect 14 37814 87 37818
rect 121 37843 194 37848
rect 121 37814 159 37843
rect 14 37809 159 37814
rect 193 37809 194 37843
rect 14 37784 194 37809
rect 14 37750 15 37784
rect 49 37780 194 37784
rect 49 37750 87 37780
rect 14 37746 87 37750
rect 121 37775 194 37780
rect 121 37746 159 37775
rect 14 37741 159 37746
rect 193 37741 194 37775
rect 14 37716 194 37741
rect 14 37682 15 37716
rect 49 37712 194 37716
rect 49 37682 87 37712
rect 14 37678 87 37682
rect 121 37707 194 37712
rect 121 37678 159 37707
rect 14 37673 159 37678
rect 193 37673 194 37707
rect 14 37648 194 37673
rect 14 37614 15 37648
rect 49 37644 194 37648
rect 49 37614 87 37644
rect 14 37610 87 37614
rect 121 37639 194 37644
rect 121 37610 159 37639
rect 14 37605 159 37610
rect 193 37605 194 37639
rect 14 37580 194 37605
rect 14 37546 15 37580
rect 49 37576 194 37580
rect 49 37546 87 37576
rect 14 37542 87 37546
rect 121 37571 194 37576
rect 121 37542 159 37571
rect 14 37537 159 37542
rect 193 37537 194 37571
rect 14 37512 194 37537
rect 14 37478 15 37512
rect 49 37508 194 37512
rect 49 37478 87 37508
rect 14 37474 87 37478
rect 121 37503 194 37508
rect 121 37474 159 37503
rect 14 37469 159 37474
rect 193 37469 194 37503
rect 14 37444 194 37469
rect 14 37410 15 37444
rect 49 37440 194 37444
rect 49 37410 87 37440
rect 14 37406 87 37410
rect 121 37435 194 37440
rect 121 37406 159 37435
rect 14 37401 159 37406
rect 193 37401 194 37435
rect 14 37376 194 37401
rect 14 37342 15 37376
rect 49 37372 194 37376
rect 49 37342 87 37372
rect 14 37338 87 37342
rect 121 37367 194 37372
rect 121 37338 159 37367
rect 14 37333 159 37338
rect 193 37333 194 37367
rect 14 37308 194 37333
rect 14 37274 15 37308
rect 49 37304 194 37308
rect 49 37274 87 37304
rect 14 37270 87 37274
rect 121 37299 194 37304
rect 121 37270 159 37299
rect 14 37265 159 37270
rect 193 37265 194 37299
rect 14 37240 194 37265
rect 14 37206 15 37240
rect 49 37236 194 37240
rect 49 37206 87 37236
rect 14 37202 87 37206
rect 121 37231 194 37236
rect 121 37202 159 37231
rect 14 37197 159 37202
rect 193 37197 194 37231
rect 14 37172 194 37197
rect 14 37138 15 37172
rect 49 37168 194 37172
rect 49 37138 87 37168
rect 14 37134 87 37138
rect 121 37163 194 37168
rect 121 37134 159 37163
rect 14 37129 159 37134
rect 193 37129 194 37163
rect 14 37104 194 37129
rect 14 37070 15 37104
rect 49 37100 194 37104
rect 49 37070 87 37100
rect 14 37066 87 37070
rect 121 37095 194 37100
rect 121 37066 159 37095
rect 14 37061 159 37066
rect 193 37061 194 37095
rect 14 37036 194 37061
rect 14 37002 15 37036
rect 49 37032 194 37036
rect 49 37002 87 37032
rect 14 36998 87 37002
rect 121 37027 194 37032
rect 121 36998 159 37027
rect 14 36993 159 36998
rect 193 36993 194 37027
rect 14 36968 194 36993
rect 14 36934 15 36968
rect 49 36964 194 36968
rect 49 36934 87 36964
rect 14 36930 87 36934
rect 121 36959 194 36964
rect 121 36930 159 36959
rect 14 36925 159 36930
rect 193 36925 194 36959
rect 14 36900 194 36925
rect 14 36866 15 36900
rect 49 36896 194 36900
rect 49 36866 87 36896
rect 14 36862 87 36866
rect 121 36891 194 36896
rect 121 36862 159 36891
rect 14 36857 159 36862
rect 193 36857 194 36891
rect 14 36832 194 36857
rect 14 36798 15 36832
rect 49 36828 194 36832
rect 49 36798 87 36828
rect 14 36794 87 36798
rect 121 36823 194 36828
rect 121 36794 159 36823
rect 14 36789 159 36794
rect 193 36789 194 36823
rect 14 36764 194 36789
rect 14 36730 15 36764
rect 49 36760 194 36764
rect 49 36730 87 36760
rect 14 36726 87 36730
rect 121 36755 194 36760
rect 121 36726 159 36755
rect 14 36721 159 36726
rect 193 36721 194 36755
rect 14 36696 194 36721
rect 14 36662 15 36696
rect 49 36692 194 36696
rect 49 36662 87 36692
rect 14 36658 87 36662
rect 121 36687 194 36692
rect 121 36658 159 36687
rect 14 36653 159 36658
rect 193 36653 194 36687
rect 14 36628 194 36653
rect 14 36594 15 36628
rect 49 36624 194 36628
rect 49 36594 87 36624
rect 14 36590 87 36594
rect 121 36619 194 36624
rect 121 36590 159 36619
rect 14 36585 159 36590
rect 193 36585 194 36619
rect 14 36560 194 36585
rect 14 36526 15 36560
rect 49 36556 194 36560
rect 49 36526 87 36556
rect 14 36522 87 36526
rect 121 36551 194 36556
rect 121 36522 159 36551
rect 14 36517 159 36522
rect 193 36517 194 36551
rect 14 36492 194 36517
rect 14 36458 15 36492
rect 49 36488 194 36492
rect 49 36458 87 36488
rect 14 36454 87 36458
rect 121 36483 194 36488
rect 121 36454 159 36483
rect 14 36449 159 36454
rect 193 36449 194 36483
rect 14 36424 194 36449
rect 14 36390 15 36424
rect 49 36420 194 36424
rect 49 36390 87 36420
rect 14 36386 87 36390
rect 121 36415 194 36420
rect 121 36386 159 36415
rect 14 36381 159 36386
rect 193 36381 194 36415
rect 14 36356 194 36381
rect 14 36322 15 36356
rect 49 36352 194 36356
rect 49 36322 87 36352
rect 14 36318 87 36322
rect 121 36347 194 36352
rect 121 36318 159 36347
rect 14 36313 159 36318
rect 193 36313 194 36347
rect 14 36288 194 36313
rect 14 36254 15 36288
rect 49 36284 194 36288
rect 49 36254 87 36284
rect 14 36250 87 36254
rect 121 36279 194 36284
rect 121 36250 159 36279
rect 14 36245 159 36250
rect 193 36245 194 36279
rect 14 36220 194 36245
rect 14 36186 15 36220
rect 49 36216 194 36220
rect 49 36186 87 36216
rect 14 36182 87 36186
rect 121 36211 194 36216
rect 121 36182 159 36211
rect 14 36177 159 36182
rect 193 36177 194 36211
rect 14 36152 194 36177
rect 14 36118 15 36152
rect 49 36148 194 36152
rect 49 36118 87 36148
rect 14 36114 87 36118
rect 121 36143 194 36148
rect 121 36114 159 36143
rect 14 36109 159 36114
rect 193 36109 194 36143
rect 14 36084 194 36109
rect 14 36050 15 36084
rect 49 36080 194 36084
rect 49 36050 87 36080
rect 14 36046 87 36050
rect 121 36075 194 36080
rect 121 36046 159 36075
rect 14 36041 159 36046
rect 193 36041 194 36075
rect 14 36016 194 36041
rect 14 35982 15 36016
rect 49 36012 194 36016
rect 49 35982 87 36012
rect 14 35978 87 35982
rect 121 36007 194 36012
rect 121 35978 159 36007
rect 14 35973 159 35978
rect 193 35973 194 36007
rect 14 35948 194 35973
rect 14 35914 15 35948
rect 49 35944 194 35948
rect 49 35914 87 35944
rect 14 35910 87 35914
rect 121 35939 194 35944
rect 121 35910 159 35939
rect 14 35905 159 35910
rect 193 35905 194 35939
rect 14 35880 194 35905
rect 14 35846 15 35880
rect 49 35876 194 35880
rect 49 35846 87 35876
rect 14 35842 87 35846
rect 121 35871 194 35876
rect 121 35842 159 35871
rect 14 35837 159 35842
rect 193 35837 194 35871
rect 14 35812 194 35837
rect 14 35778 15 35812
rect 49 35808 194 35812
rect 49 35778 87 35808
rect 14 35774 87 35778
rect 121 35803 194 35808
rect 121 35774 159 35803
rect 14 35769 159 35774
rect 193 35769 194 35803
rect 14 35744 194 35769
rect 14 35710 15 35744
rect 49 35740 194 35744
rect 49 35710 87 35740
rect 14 35706 87 35710
rect 121 35735 194 35740
rect 121 35706 159 35735
rect 14 35701 159 35706
rect 193 35701 194 35735
rect 14 35676 194 35701
rect 14 35642 15 35676
rect 49 35672 194 35676
rect 49 35642 87 35672
rect 14 35638 87 35642
rect 121 35667 194 35672
rect 121 35638 159 35667
rect 14 35633 159 35638
rect 193 35633 194 35667
rect 14 35608 194 35633
rect 14 35574 15 35608
rect 49 35604 194 35608
rect 49 35574 87 35604
rect 14 35570 87 35574
rect 121 35599 194 35604
rect 121 35570 159 35599
rect 14 35565 159 35570
rect 193 35565 194 35599
rect 14 35540 194 35565
rect 14 35506 15 35540
rect 49 35536 194 35540
rect 49 35506 87 35536
rect 14 35502 87 35506
rect 121 35531 194 35536
rect 121 35502 159 35531
rect 14 35497 159 35502
rect 193 35497 194 35531
rect 14 35472 194 35497
rect 14 35438 15 35472
rect 49 35468 194 35472
rect 49 35438 87 35468
rect 14 35434 87 35438
rect 121 35463 194 35468
rect 121 35434 159 35463
rect 14 35429 159 35434
rect 193 35429 194 35463
rect 14 35404 194 35429
rect 14 35370 15 35404
rect 49 35400 194 35404
rect 49 35370 87 35400
rect 14 35366 87 35370
rect 121 35395 194 35400
rect 121 35366 159 35395
rect 14 35361 159 35366
rect 193 35361 194 35395
rect 14 35336 194 35361
rect 14 35302 15 35336
rect 49 35332 194 35336
rect 49 35302 87 35332
rect 14 35298 87 35302
rect 121 35327 194 35332
rect 121 35298 159 35327
rect 14 35293 159 35298
rect 193 35293 194 35327
rect 14 35268 194 35293
rect 14 35234 15 35268
rect 49 35264 194 35268
rect 49 35234 87 35264
rect 14 35230 87 35234
rect 121 35259 194 35264
rect 121 35230 159 35259
rect 14 35225 159 35230
rect 193 35225 194 35259
rect 14 35200 194 35225
rect 14 35166 15 35200
rect 49 35196 194 35200
rect 49 35166 87 35196
rect 14 35162 87 35166
rect 121 35191 194 35196
rect 121 35162 159 35191
rect 14 35157 159 35162
rect 193 35157 194 35191
rect 14 35132 194 35157
rect 14 35098 15 35132
rect 49 35128 194 35132
rect 49 35098 87 35128
rect 14 35094 87 35098
rect 121 35123 194 35128
rect 121 35094 159 35123
rect 14 35089 159 35094
rect 193 35089 194 35123
rect 14 35064 194 35089
rect 14 35030 15 35064
rect 49 35060 194 35064
rect 49 35030 87 35060
rect 14 35026 87 35030
rect 121 35055 194 35060
rect 121 35026 159 35055
rect 14 35021 159 35026
rect 193 35021 194 35055
rect 14 34996 194 35021
rect 14 34962 15 34996
rect 49 34992 194 34996
rect 49 34962 87 34992
rect 14 34958 87 34962
rect 121 34987 194 34992
rect 121 34958 159 34987
rect 14 34953 159 34958
rect 193 34953 194 34987
rect 14 34928 194 34953
rect 14 34894 15 34928
rect 49 34924 194 34928
rect 49 34894 87 34924
rect 14 34890 87 34894
rect 121 34919 194 34924
rect 121 34890 159 34919
rect 14 34885 159 34890
rect 193 34885 194 34919
rect 14 34861 194 34885
rect -2867 34860 194 34861
rect -2867 34826 -2833 34860
rect -2799 34826 -2765 34860
rect -2731 34826 -2697 34860
rect -2663 34826 -2629 34860
rect -2595 34826 -2561 34860
rect -2527 34826 -2493 34860
rect -2459 34826 -2425 34860
rect -2391 34826 -2357 34860
rect -2323 34826 -2289 34860
rect -2255 34826 -2221 34860
rect -2187 34826 -2153 34860
rect -2119 34826 -2085 34860
rect -2051 34826 -2017 34860
rect -1983 34826 -1949 34860
rect -1915 34826 -1881 34860
rect -1847 34826 -1813 34860
rect -1779 34826 -1745 34860
rect -1711 34826 -1677 34860
rect -1643 34826 -1609 34860
rect -1575 34826 -1541 34860
rect -1507 34826 -1473 34860
rect -1439 34826 -1405 34860
rect -1371 34826 -1337 34860
rect -1303 34826 -1269 34860
rect -1235 34826 -1201 34860
rect -1167 34826 -1133 34860
rect -1099 34826 -1065 34860
rect -1031 34826 -997 34860
rect -963 34826 -929 34860
rect -895 34826 -861 34860
rect -827 34826 -793 34860
rect -759 34826 -725 34860
rect -691 34826 -657 34860
rect -623 34826 -589 34860
rect -555 34826 -521 34860
rect -487 34826 -453 34860
rect -419 34826 -385 34860
rect -351 34826 -317 34860
rect -283 34826 -249 34860
rect -215 34826 -181 34860
rect -147 34826 -113 34860
rect -79 34826 15 34860
rect 49 34856 194 34860
rect 49 34826 87 34856
rect -2867 34822 87 34826
rect 121 34851 194 34856
rect 121 34822 159 34851
rect -2867 34817 159 34822
rect 193 34817 194 34851
rect -2867 34788 194 34817
rect -2867 34754 -2833 34788
rect -2799 34754 -2765 34788
rect -2731 34754 -2697 34788
rect -2663 34754 -2629 34788
rect -2595 34754 -2561 34788
rect -2527 34754 -2493 34788
rect -2459 34754 -2425 34788
rect -2391 34754 -2357 34788
rect -2323 34754 -2289 34788
rect -2255 34754 -2221 34788
rect -2187 34754 -2153 34788
rect -2119 34754 -2085 34788
rect -2051 34754 -2017 34788
rect -1983 34754 -1949 34788
rect -1915 34754 -1881 34788
rect -1847 34754 -1813 34788
rect -1779 34754 -1745 34788
rect -1711 34754 -1677 34788
rect -1643 34754 -1609 34788
rect -1575 34754 -1541 34788
rect -1507 34754 -1473 34788
rect -1439 34754 -1405 34788
rect -1371 34754 -1337 34788
rect -1303 34754 -1269 34788
rect -1235 34754 -1201 34788
rect -1167 34754 -1133 34788
rect -1099 34754 -1065 34788
rect -1031 34754 -997 34788
rect -963 34754 -929 34788
rect -895 34754 -861 34788
rect -827 34754 -793 34788
rect -759 34754 -725 34788
rect -691 34754 -657 34788
rect -623 34754 -589 34788
rect -555 34754 -521 34788
rect -487 34754 -453 34788
rect -419 34754 -385 34788
rect -351 34754 -317 34788
rect -283 34754 -249 34788
rect -215 34754 -181 34788
rect -147 34754 -113 34788
rect -79 34754 -45 34788
rect -11 34754 87 34788
rect 121 34783 194 34788
rect 121 34754 159 34783
rect -2867 34749 159 34754
rect 193 34749 194 34783
rect -2867 34716 194 34749
rect -2867 34682 -2833 34716
rect -2799 34682 -2765 34716
rect -2731 34682 -2697 34716
rect -2663 34682 -2629 34716
rect -2595 34682 -2561 34716
rect -2527 34682 -2493 34716
rect -2459 34682 -2425 34716
rect -2391 34682 -2357 34716
rect -2323 34682 -2289 34716
rect -2255 34682 -2221 34716
rect -2187 34682 -2153 34716
rect -2119 34682 -2085 34716
rect -2051 34682 -2017 34716
rect -1983 34682 -1949 34716
rect -1915 34682 -1881 34716
rect -1847 34682 -1813 34716
rect -1779 34682 -1745 34716
rect -1711 34682 -1677 34716
rect -1643 34682 -1609 34716
rect -1575 34682 -1541 34716
rect -1507 34682 -1473 34716
rect -1439 34682 -1405 34716
rect -1371 34682 -1337 34716
rect -1303 34682 -1269 34716
rect -1235 34682 -1201 34716
rect -1167 34682 -1133 34716
rect -1099 34682 -1065 34716
rect -1031 34682 -997 34716
rect -963 34682 -929 34716
rect -895 34682 -861 34716
rect -827 34682 -793 34716
rect -759 34682 -725 34716
rect -691 34682 -657 34716
rect -623 34682 -589 34716
rect -555 34682 -521 34716
rect -487 34682 -453 34716
rect -419 34682 -385 34716
rect -351 34682 -317 34716
rect -283 34682 -249 34716
rect -215 34682 -181 34716
rect -147 34682 -113 34716
rect -79 34682 -45 34716
rect -11 34682 23 34716
rect 57 34682 91 34716
rect 125 34682 194 34716
rect -2867 34647 194 34682
<< psubdiffcont >>
rect 4429 11332 6231 11910
rect 4429 11263 4463 11297
rect 4497 11263 4531 11297
rect 4565 11263 4599 11297
rect 4633 11263 4667 11297
rect 4701 11263 4735 11297
rect 4769 11263 4803 11297
rect 4837 11263 4871 11297
rect 4905 11263 4939 11297
rect 4973 11263 5007 11297
rect 5041 11263 5075 11297
rect 5109 11263 5143 11297
rect 5177 11263 5211 11297
rect 5245 11263 5279 11297
rect 5313 11263 5347 11297
rect 5381 11263 5415 11297
rect 5449 11263 5483 11297
rect 5517 11263 5551 11297
rect 5585 11263 5619 11297
rect 5653 11263 5687 11297
rect 5721 11263 5755 11297
rect 5789 11263 5823 11297
rect 5857 11263 5891 11297
rect 5925 11263 5959 11297
rect 5993 11263 6027 11297
rect 6061 11263 6095 11297
rect 6129 11263 6163 11297
rect 6197 11263 6231 11297
rect 4429 11194 4463 11228
rect 4497 11194 4531 11228
rect 4565 11194 4599 11228
rect 4633 11194 4667 11228
rect 4701 11194 4735 11228
rect 4769 11194 4803 11228
rect 4837 11194 4871 11228
rect 4905 11194 4939 11228
rect 4973 11194 5007 11228
rect 5041 11194 5075 11228
rect 5109 11194 5143 11228
rect 5177 11194 5211 11228
rect 5245 11194 5279 11228
rect 5313 11194 5347 11228
rect 5381 11194 5415 11228
rect 5449 11194 5483 11228
rect 5517 11194 5551 11228
rect 5585 11194 5619 11228
rect 5653 11194 5687 11228
rect 5721 11194 5755 11228
rect 5789 11194 5823 11228
rect 5857 11194 5891 11228
rect 5925 11194 5959 11228
rect 5993 11194 6027 11228
rect 6061 11194 6095 11228
rect 6129 11194 6163 11228
rect 6197 11194 6231 11228
rect 4429 11125 4463 11159
rect 4497 11125 4531 11159
rect 4565 11125 4599 11159
rect 4633 11125 4667 11159
rect 4701 11125 4735 11159
rect 4769 11125 4803 11159
rect 4837 11125 4871 11159
rect 4905 11125 4939 11159
rect 4973 11125 5007 11159
rect 5041 11125 5075 11159
rect 5109 11125 5143 11159
rect 5177 11125 5211 11159
rect 5245 11125 5279 11159
rect 5313 11125 5347 11159
rect 5381 11125 5415 11159
rect 5449 11125 5483 11159
rect 5517 11125 5551 11159
rect 5585 11125 5619 11159
rect 5653 11125 5687 11159
rect 5721 11125 5755 11159
rect 5789 11125 5823 11159
rect 5857 11125 5891 11159
rect 5925 11125 5959 11159
rect 5993 11125 6027 11159
rect 6061 11125 6095 11159
rect 6129 11125 6163 11159
rect 6197 11125 6231 11159
rect 4429 11056 4463 11090
rect 4497 11056 4531 11090
rect 4565 11056 4599 11090
rect 4633 11056 4667 11090
rect 4701 11056 4735 11090
rect 4769 11056 4803 11090
rect 4837 11056 4871 11090
rect 4905 11056 4939 11090
rect 4973 11056 5007 11090
rect 5041 11056 5075 11090
rect 5109 11056 5143 11090
rect 5177 11056 5211 11090
rect 5245 11056 5279 11090
rect 5313 11056 5347 11090
rect 5381 11056 5415 11090
rect 5449 11056 5483 11090
rect 5517 11056 5551 11090
rect 5585 11056 5619 11090
rect 5653 11056 5687 11090
rect 5721 11056 5755 11090
rect 5789 11056 5823 11090
rect 5857 11056 5891 11090
rect 5925 11056 5959 11090
rect 5993 11056 6027 11090
rect 6061 11056 6095 11090
rect 6129 11056 6163 11090
rect 6197 11056 6231 11090
rect 4429 10987 4463 11021
rect 4497 10987 4531 11021
rect 4565 10987 4599 11021
rect 4633 10987 4667 11021
rect 4701 10987 4735 11021
rect 4769 10987 4803 11021
rect 4837 10987 4871 11021
rect 4905 10987 4939 11021
rect 4973 10987 5007 11021
rect 5041 10987 5075 11021
rect 5109 10987 5143 11021
rect 5177 10987 5211 11021
rect 5245 10987 5279 11021
rect 5313 10987 5347 11021
rect 5381 10987 5415 11021
rect 5449 10987 5483 11021
rect 5517 10987 5551 11021
rect 5585 10987 5619 11021
rect 5653 10987 5687 11021
rect 5721 10987 5755 11021
rect 5789 10987 5823 11021
rect 5857 10987 5891 11021
rect 5925 10987 5959 11021
rect 5993 10987 6027 11021
rect 6061 10987 6095 11021
rect 6129 10987 6163 11021
rect 6197 10987 6231 11021
rect 4429 10918 4463 10952
rect 4497 10918 4531 10952
rect 4565 10918 4599 10952
rect 4633 10918 4667 10952
rect 4701 10918 4735 10952
rect 4769 10918 4803 10952
rect 4837 10918 4871 10952
rect 4905 10918 4939 10952
rect 4973 10918 5007 10952
rect 5041 10918 5075 10952
rect 5109 10918 5143 10952
rect 5177 10918 5211 10952
rect 5245 10918 5279 10952
rect 5313 10918 5347 10952
rect 5381 10918 5415 10952
rect 5449 10918 5483 10952
rect 5517 10918 5551 10952
rect 5585 10918 5619 10952
rect 5653 10918 5687 10952
rect 5721 10918 5755 10952
rect 5789 10918 5823 10952
rect 5857 10918 5891 10952
rect 5925 10918 5959 10952
rect 5993 10918 6027 10952
rect 6061 10918 6095 10952
rect 6129 10918 6163 10952
rect 6197 10918 6231 10952
rect 4429 10849 4463 10883
rect 4497 10849 4531 10883
rect 4565 10849 4599 10883
rect 4633 10849 4667 10883
rect 4701 10849 4735 10883
rect 4769 10849 4803 10883
rect 4837 10849 4871 10883
rect 4905 10849 4939 10883
rect 4973 10849 5007 10883
rect 5041 10849 5075 10883
rect 5109 10849 5143 10883
rect 5177 10849 5211 10883
rect 5245 10849 5279 10883
rect 5313 10849 5347 10883
rect 5381 10849 5415 10883
rect 5449 10849 5483 10883
rect 5517 10849 5551 10883
rect 5585 10849 5619 10883
rect 5653 10849 5687 10883
rect 5721 10849 5755 10883
rect 5789 10849 5823 10883
rect 5857 10849 5891 10883
rect 5925 10849 5959 10883
rect 5993 10849 6027 10883
rect 6061 10849 6095 10883
rect 6129 10849 6163 10883
rect 6197 10849 6231 10883
rect 4429 10780 4463 10814
rect 4497 10780 4531 10814
rect 4565 10780 4599 10814
rect 4633 10780 4667 10814
rect 4701 10780 4735 10814
rect 4769 10780 4803 10814
rect 4837 10780 4871 10814
rect 4905 10780 4939 10814
rect 4973 10780 5007 10814
rect 5041 10780 5075 10814
rect 5109 10780 5143 10814
rect 5177 10780 5211 10814
rect 5245 10780 5279 10814
rect 5313 10780 5347 10814
rect 5381 10780 5415 10814
rect 5449 10780 5483 10814
rect 5517 10780 5551 10814
rect 5585 10780 5619 10814
rect 5653 10780 5687 10814
rect 5721 10780 5755 10814
rect 5789 10780 5823 10814
rect 5857 10780 5891 10814
rect 5925 10780 5959 10814
rect 5993 10780 6027 10814
rect 6061 10780 6095 10814
rect 6129 10780 6163 10814
rect 6197 10780 6231 10814
rect 4429 10711 4463 10745
rect 4497 10711 4531 10745
rect 4565 10711 4599 10745
rect 4633 10711 4667 10745
rect 4701 10711 4735 10745
rect 4769 10711 4803 10745
rect 4837 10711 4871 10745
rect 4905 10711 4939 10745
rect 4973 10711 5007 10745
rect 5041 10711 5075 10745
rect 5109 10711 5143 10745
rect 5177 10711 5211 10745
rect 5245 10711 5279 10745
rect 5313 10711 5347 10745
rect 5381 10711 5415 10745
rect 5449 10711 5483 10745
rect 5517 10711 5551 10745
rect 5585 10711 5619 10745
rect 5653 10711 5687 10745
rect 5721 10711 5755 10745
rect 5789 10711 5823 10745
rect 5857 10711 5891 10745
rect 5925 10711 5959 10745
rect 5993 10711 6027 10745
rect 6061 10711 6095 10745
rect 6129 10711 6163 10745
rect 6197 10711 6231 10745
rect 4429 10642 4463 10676
rect 4497 10642 4531 10676
rect 4565 10642 4599 10676
rect 4633 10642 4667 10676
rect 4701 10642 4735 10676
rect 4769 10642 4803 10676
rect 4837 10642 4871 10676
rect 4905 10642 4939 10676
rect 4973 10642 5007 10676
rect 5041 10642 5075 10676
rect 5109 10642 5143 10676
rect 5177 10642 5211 10676
rect 5245 10642 5279 10676
rect 5313 10642 5347 10676
rect 5381 10642 5415 10676
rect 5449 10642 5483 10676
rect 5517 10642 5551 10676
rect 5585 10642 5619 10676
rect 5653 10642 5687 10676
rect 5721 10642 5755 10676
rect 5789 10642 5823 10676
rect 5857 10642 5891 10676
rect 5925 10642 5959 10676
rect 5993 10642 6027 10676
rect 6061 10642 6095 10676
rect 6129 10642 6163 10676
rect 6197 10642 6231 10676
rect 4429 10573 4463 10607
rect 4497 10573 4531 10607
rect 4565 10573 4599 10607
rect 4633 10573 4667 10607
rect 4701 10573 4735 10607
rect 4769 10573 4803 10607
rect 4837 10573 4871 10607
rect 4905 10573 4939 10607
rect 4973 10573 5007 10607
rect 5041 10573 5075 10607
rect 5109 10573 5143 10607
rect 5177 10573 5211 10607
rect 5245 10573 5279 10607
rect 5313 10573 5347 10607
rect 5381 10573 5415 10607
rect 5449 10573 5483 10607
rect 5517 10573 5551 10607
rect 5585 10573 5619 10607
rect 5653 10573 5687 10607
rect 5721 10573 5755 10607
rect 5789 10573 5823 10607
rect 5857 10573 5891 10607
rect 5925 10573 5959 10607
rect 5993 10573 6027 10607
rect 6061 10573 6095 10607
rect 6129 10573 6163 10607
rect 6197 10573 6231 10607
rect 4429 10504 4463 10538
rect 4497 10504 4531 10538
rect 4565 10504 4599 10538
rect 4633 10504 4667 10538
rect 4701 10504 4735 10538
rect 4769 10504 4803 10538
rect 4837 10504 4871 10538
rect 4905 10504 4939 10538
rect 4973 10504 5007 10538
rect 5041 10504 5075 10538
rect 5109 10504 5143 10538
rect 5177 10504 5211 10538
rect 5245 10504 5279 10538
rect 5313 10504 5347 10538
rect 5381 10504 5415 10538
rect 5449 10504 5483 10538
rect 5517 10504 5551 10538
rect 5585 10504 5619 10538
rect 5653 10504 5687 10538
rect 5721 10504 5755 10538
rect 5789 10504 5823 10538
rect 5857 10504 5891 10538
rect 5925 10504 5959 10538
rect 5993 10504 6027 10538
rect 6061 10504 6095 10538
rect 6129 10504 6163 10538
rect 6197 10504 6231 10538
rect 4429 10435 4463 10469
rect 4497 10435 4531 10469
rect 4565 10435 4599 10469
rect 4633 10435 4667 10469
rect 4701 10435 4735 10469
rect 4769 10435 4803 10469
rect 4837 10435 4871 10469
rect 4905 10435 4939 10469
rect 4973 10435 5007 10469
rect 5041 10435 5075 10469
rect 5109 10435 5143 10469
rect 5177 10435 5211 10469
rect 5245 10435 5279 10469
rect 5313 10435 5347 10469
rect 5381 10435 5415 10469
rect 5449 10435 5483 10469
rect 5517 10435 5551 10469
rect 5585 10435 5619 10469
rect 5653 10435 5687 10469
rect 5721 10435 5755 10469
rect 5789 10435 5823 10469
rect 5857 10435 5891 10469
rect 5925 10435 5959 10469
rect 5993 10435 6027 10469
rect 6061 10435 6095 10469
rect 6129 10435 6163 10469
rect 6197 10435 6231 10469
rect 4429 10366 4463 10400
rect 4497 10366 4531 10400
rect 4565 10366 4599 10400
rect 4633 10366 4667 10400
rect 4701 10366 4735 10400
rect 4769 10366 4803 10400
rect 4837 10366 4871 10400
rect 4905 10366 4939 10400
rect 4973 10366 5007 10400
rect 5041 10366 5075 10400
rect 5109 10366 5143 10400
rect 5177 10366 5211 10400
rect 5245 10366 5279 10400
rect 5313 10366 5347 10400
rect 5381 10366 5415 10400
rect 5449 10366 5483 10400
rect 5517 10366 5551 10400
rect 5585 10366 5619 10400
rect 5653 10366 5687 10400
rect 5721 10366 5755 10400
rect 5789 10366 5823 10400
rect 5857 10366 5891 10400
rect 5925 10366 5959 10400
rect 5993 10366 6027 10400
rect 6061 10366 6095 10400
rect 6129 10366 6163 10400
rect 6197 10366 6231 10400
rect 4429 10297 4463 10331
rect 4497 10297 4531 10331
rect 4565 10297 4599 10331
rect 4633 10297 4667 10331
rect 4701 10297 4735 10331
rect 4769 10297 4803 10331
rect 4837 10297 4871 10331
rect 4905 10297 4939 10331
rect 4973 10297 5007 10331
rect 5041 10297 5075 10331
rect 5109 10297 5143 10331
rect 5177 10297 5211 10331
rect 5245 10297 5279 10331
rect 5313 10297 5347 10331
rect 5381 10297 5415 10331
rect 5449 10297 5483 10331
rect 5517 10297 5551 10331
rect 5585 10297 5619 10331
rect 5653 10297 5687 10331
rect 5721 10297 5755 10331
rect 5789 10297 5823 10331
rect 5857 10297 5891 10331
rect 5925 10297 5959 10331
rect 5993 10297 6027 10331
rect 6061 10297 6095 10331
rect 6129 10297 6163 10331
rect 6197 10297 6231 10331
rect 4429 10228 4463 10262
rect 4497 10228 4531 10262
rect 4565 10228 4599 10262
rect 4633 10228 4667 10262
rect 4701 10228 4735 10262
rect 4769 10228 4803 10262
rect 4837 10228 4871 10262
rect 4905 10228 4939 10262
rect 4973 10228 5007 10262
rect 5041 10228 5075 10262
rect 5109 10228 5143 10262
rect 5177 10228 5211 10262
rect 5245 10228 5279 10262
rect 5313 10228 5347 10262
rect 5381 10228 5415 10262
rect 5449 10228 5483 10262
rect 5517 10228 5551 10262
rect 5585 10228 5619 10262
rect 5653 10228 5687 10262
rect 5721 10228 5755 10262
rect 5789 10228 5823 10262
rect 5857 10228 5891 10262
rect 5925 10228 5959 10262
rect 5993 10228 6027 10262
rect 6061 10228 6095 10262
rect 6129 10228 6163 10262
rect 6197 10228 6231 10262
rect 4429 10159 4463 10193
rect 4497 10159 4531 10193
rect 4565 10159 4599 10193
rect 4633 10159 4667 10193
rect 4701 10159 4735 10193
rect 4769 10159 4803 10193
rect 4837 10159 4871 10193
rect 4905 10159 4939 10193
rect 4973 10159 5007 10193
rect 5041 10159 5075 10193
rect 5109 10159 5143 10193
rect 5177 10159 5211 10193
rect 5245 10159 5279 10193
rect 5313 10159 5347 10193
rect 5381 10159 5415 10193
rect 5449 10159 5483 10193
rect 5517 10159 5551 10193
rect 5585 10159 5619 10193
rect 5653 10159 5687 10193
rect 5721 10159 5755 10193
rect 5789 10159 5823 10193
rect 5857 10159 5891 10193
rect 5925 10159 5959 10193
rect 5993 10159 6027 10193
rect 6061 10159 6095 10193
rect 6129 10159 6163 10193
rect 6197 10159 6231 10193
rect 4429 10090 4463 10124
rect 4497 10090 4531 10124
rect 4565 10090 4599 10124
rect 4633 10090 4667 10124
rect 4701 10090 4735 10124
rect 4769 10090 4803 10124
rect 4837 10090 4871 10124
rect 4905 10090 4939 10124
rect 4973 10090 5007 10124
rect 5041 10090 5075 10124
rect 5109 10090 5143 10124
rect 5177 10090 5211 10124
rect 5245 10090 5279 10124
rect 5313 10090 5347 10124
rect 5381 10090 5415 10124
rect 5449 10090 5483 10124
rect 5517 10090 5551 10124
rect 5585 10090 5619 10124
rect 5653 10090 5687 10124
rect 5721 10090 5755 10124
rect 5789 10090 5823 10124
rect 5857 10090 5891 10124
rect 5925 10090 5959 10124
rect 5993 10090 6027 10124
rect 6061 10090 6095 10124
rect 6129 10090 6163 10124
rect 6197 10090 6231 10124
<< mvpsubdiffcont >>
rect -2938 37942 -184 50624
rect -2938 37873 -2904 37907
rect -2870 37873 -2836 37907
rect -2802 37873 -2768 37907
rect -2734 37873 -2700 37907
rect -2666 37873 -2632 37907
rect -2598 37873 -2564 37907
rect -2530 37873 -2496 37907
rect -2462 37873 -2428 37907
rect -2394 37873 -2360 37907
rect -2326 37873 -2292 37907
rect -2258 37873 -2224 37907
rect -2190 37873 -2156 37907
rect -2122 37873 -2088 37907
rect -2054 37873 -2020 37907
rect -1986 37873 -1952 37907
rect -1918 37873 -1884 37907
rect -1850 37873 -1816 37907
rect -1782 37873 -1748 37907
rect -1714 37873 -1680 37907
rect -1646 37873 -1612 37907
rect -1578 37873 -1544 37907
rect -1510 37873 -1476 37907
rect -1442 37873 -1408 37907
rect -1374 37873 -1340 37907
rect -1306 37873 -1272 37907
rect -1238 37873 -1204 37907
rect -1170 37873 -1136 37907
rect -1102 37873 -1068 37907
rect -1034 37873 -1000 37907
rect -966 37873 -932 37907
rect -898 37873 -864 37907
rect -830 37873 -796 37907
rect -762 37873 -728 37907
rect -694 37873 -660 37907
rect -626 37873 -592 37907
rect -558 37873 -524 37907
rect -490 37873 -456 37907
rect -422 37873 -388 37907
rect -354 37873 -320 37907
rect -286 37873 -252 37907
rect -218 37873 -184 37907
rect -2938 37804 -2904 37838
rect -2870 37804 -2836 37838
rect -2802 37804 -2768 37838
rect -2734 37804 -2700 37838
rect -2666 37804 -2632 37838
rect -2598 37804 -2564 37838
rect -2530 37804 -2496 37838
rect -2462 37804 -2428 37838
rect -2394 37804 -2360 37838
rect -2326 37804 -2292 37838
rect -2258 37804 -2224 37838
rect -2190 37804 -2156 37838
rect -2122 37804 -2088 37838
rect -2054 37804 -2020 37838
rect -1986 37804 -1952 37838
rect -1918 37804 -1884 37838
rect -1850 37804 -1816 37838
rect -1782 37804 -1748 37838
rect -1714 37804 -1680 37838
rect -1646 37804 -1612 37838
rect -1578 37804 -1544 37838
rect -1510 37804 -1476 37838
rect -1442 37804 -1408 37838
rect -1374 37804 -1340 37838
rect -1306 37804 -1272 37838
rect -1238 37804 -1204 37838
rect -1170 37804 -1136 37838
rect -1102 37804 -1068 37838
rect -1034 37804 -1000 37838
rect -966 37804 -932 37838
rect -898 37804 -864 37838
rect -830 37804 -796 37838
rect -762 37804 -728 37838
rect -694 37804 -660 37838
rect -626 37804 -592 37838
rect -558 37804 -524 37838
rect -490 37804 -456 37838
rect -422 37804 -388 37838
rect -354 37804 -320 37838
rect -286 37804 -252 37838
rect -218 37804 -184 37838
rect -2938 37735 -2904 37769
rect -2870 37735 -2836 37769
rect -2802 37735 -2768 37769
rect -2734 37735 -2700 37769
rect -2666 37735 -2632 37769
rect -2598 37735 -2564 37769
rect -2530 37735 -2496 37769
rect -2462 37735 -2428 37769
rect -2394 37735 -2360 37769
rect -2326 37735 -2292 37769
rect -2258 37735 -2224 37769
rect -2190 37735 -2156 37769
rect -2122 37735 -2088 37769
rect -2054 37735 -2020 37769
rect -1986 37735 -1952 37769
rect -1918 37735 -1884 37769
rect -1850 37735 -1816 37769
rect -1782 37735 -1748 37769
rect -1714 37735 -1680 37769
rect -1646 37735 -1612 37769
rect -1578 37735 -1544 37769
rect -1510 37735 -1476 37769
rect -1442 37735 -1408 37769
rect -1374 37735 -1340 37769
rect -1306 37735 -1272 37769
rect -1238 37735 -1204 37769
rect -1170 37735 -1136 37769
rect -1102 37735 -1068 37769
rect -1034 37735 -1000 37769
rect -966 37735 -932 37769
rect -898 37735 -864 37769
rect -830 37735 -796 37769
rect -762 37735 -728 37769
rect -694 37735 -660 37769
rect -626 37735 -592 37769
rect -558 37735 -524 37769
rect -490 37735 -456 37769
rect -422 37735 -388 37769
rect -354 37735 -320 37769
rect -286 37735 -252 37769
rect -218 37735 -184 37769
rect -2938 37666 -2904 37700
rect -2870 37666 -2836 37700
rect -2802 37666 -2768 37700
rect -2734 37666 -2700 37700
rect -2666 37666 -2632 37700
rect -2598 37666 -2564 37700
rect -2530 37666 -2496 37700
rect -2462 37666 -2428 37700
rect -2394 37666 -2360 37700
rect -2326 37666 -2292 37700
rect -2258 37666 -2224 37700
rect -2190 37666 -2156 37700
rect -2122 37666 -2088 37700
rect -2054 37666 -2020 37700
rect -1986 37666 -1952 37700
rect -1918 37666 -1884 37700
rect -1850 37666 -1816 37700
rect -1782 37666 -1748 37700
rect -1714 37666 -1680 37700
rect -1646 37666 -1612 37700
rect -1578 37666 -1544 37700
rect -1510 37666 -1476 37700
rect -1442 37666 -1408 37700
rect -1374 37666 -1340 37700
rect -1306 37666 -1272 37700
rect -1238 37666 -1204 37700
rect -1170 37666 -1136 37700
rect -1102 37666 -1068 37700
rect -1034 37666 -1000 37700
rect -966 37666 -932 37700
rect -898 37666 -864 37700
rect -830 37666 -796 37700
rect -762 37666 -728 37700
rect -694 37666 -660 37700
rect -626 37666 -592 37700
rect -558 37666 -524 37700
rect -490 37666 -456 37700
rect -422 37666 -388 37700
rect -354 37666 -320 37700
rect -286 37666 -252 37700
rect -218 37666 -184 37700
rect -2938 37597 -2904 37631
rect -2870 37597 -2836 37631
rect -2802 37597 -2768 37631
rect -2734 37597 -2700 37631
rect -2666 37597 -2632 37631
rect -2598 37597 -2564 37631
rect -2530 37597 -2496 37631
rect -2462 37597 -2428 37631
rect -2394 37597 -2360 37631
rect -2326 37597 -2292 37631
rect -2258 37597 -2224 37631
rect -2190 37597 -2156 37631
rect -2122 37597 -2088 37631
rect -2054 37597 -2020 37631
rect -1986 37597 -1952 37631
rect -1918 37597 -1884 37631
rect -1850 37597 -1816 37631
rect -1782 37597 -1748 37631
rect -1714 37597 -1680 37631
rect -1646 37597 -1612 37631
rect -1578 37597 -1544 37631
rect -1510 37597 -1476 37631
rect -1442 37597 -1408 37631
rect -1374 37597 -1340 37631
rect -1306 37597 -1272 37631
rect -1238 37597 -1204 37631
rect -1170 37597 -1136 37631
rect -1102 37597 -1068 37631
rect -1034 37597 -1000 37631
rect -966 37597 -932 37631
rect -898 37597 -864 37631
rect -830 37597 -796 37631
rect -762 37597 -728 37631
rect -694 37597 -660 37631
rect -626 37597 -592 37631
rect -558 37597 -524 37631
rect -490 37597 -456 37631
rect -422 37597 -388 37631
rect -354 37597 -320 37631
rect -286 37597 -252 37631
rect -218 37597 -184 37631
rect -2938 37528 -2904 37562
rect -2870 37528 -2836 37562
rect -2802 37528 -2768 37562
rect -2734 37528 -2700 37562
rect -2666 37528 -2632 37562
rect -2598 37528 -2564 37562
rect -2530 37528 -2496 37562
rect -2462 37528 -2428 37562
rect -2394 37528 -2360 37562
rect -2326 37528 -2292 37562
rect -2258 37528 -2224 37562
rect -2190 37528 -2156 37562
rect -2122 37528 -2088 37562
rect -2054 37528 -2020 37562
rect -1986 37528 -1952 37562
rect -1918 37528 -1884 37562
rect -1850 37528 -1816 37562
rect -1782 37528 -1748 37562
rect -1714 37528 -1680 37562
rect -1646 37528 -1612 37562
rect -1578 37528 -1544 37562
rect -1510 37528 -1476 37562
rect -1442 37528 -1408 37562
rect -1374 37528 -1340 37562
rect -1306 37528 -1272 37562
rect -1238 37528 -1204 37562
rect -1170 37528 -1136 37562
rect -1102 37528 -1068 37562
rect -1034 37528 -1000 37562
rect -966 37528 -932 37562
rect -898 37528 -864 37562
rect -830 37528 -796 37562
rect -762 37528 -728 37562
rect -694 37528 -660 37562
rect -626 37528 -592 37562
rect -558 37528 -524 37562
rect -490 37528 -456 37562
rect -422 37528 -388 37562
rect -354 37528 -320 37562
rect -286 37528 -252 37562
rect -218 37528 -184 37562
rect -2938 37459 -2904 37493
rect -2870 37459 -2836 37493
rect -2802 37459 -2768 37493
rect -2734 37459 -2700 37493
rect -2666 37459 -2632 37493
rect -2598 37459 -2564 37493
rect -2530 37459 -2496 37493
rect -2462 37459 -2428 37493
rect -2394 37459 -2360 37493
rect -2326 37459 -2292 37493
rect -2258 37459 -2224 37493
rect -2190 37459 -2156 37493
rect -2122 37459 -2088 37493
rect -2054 37459 -2020 37493
rect -1986 37459 -1952 37493
rect -1918 37459 -1884 37493
rect -1850 37459 -1816 37493
rect -1782 37459 -1748 37493
rect -1714 37459 -1680 37493
rect -1646 37459 -1612 37493
rect -1578 37459 -1544 37493
rect -1510 37459 -1476 37493
rect -1442 37459 -1408 37493
rect -1374 37459 -1340 37493
rect -1306 37459 -1272 37493
rect -1238 37459 -1204 37493
rect -1170 37459 -1136 37493
rect -1102 37459 -1068 37493
rect -1034 37459 -1000 37493
rect -966 37459 -932 37493
rect -898 37459 -864 37493
rect -830 37459 -796 37493
rect -762 37459 -728 37493
rect -694 37459 -660 37493
rect -626 37459 -592 37493
rect -558 37459 -524 37493
rect -490 37459 -456 37493
rect -422 37459 -388 37493
rect -354 37459 -320 37493
rect -286 37459 -252 37493
rect -218 37459 -184 37493
rect -2938 37390 -2904 37424
rect -2870 37390 -2836 37424
rect -2802 37390 -2768 37424
rect -2734 37390 -2700 37424
rect -2666 37390 -2632 37424
rect -2598 37390 -2564 37424
rect -2530 37390 -2496 37424
rect -2462 37390 -2428 37424
rect -2394 37390 -2360 37424
rect -2326 37390 -2292 37424
rect -2258 37390 -2224 37424
rect -2190 37390 -2156 37424
rect -2122 37390 -2088 37424
rect -2054 37390 -2020 37424
rect -1986 37390 -1952 37424
rect -1918 37390 -1884 37424
rect -1850 37390 -1816 37424
rect -1782 37390 -1748 37424
rect -1714 37390 -1680 37424
rect -1646 37390 -1612 37424
rect -1578 37390 -1544 37424
rect -1510 37390 -1476 37424
rect -1442 37390 -1408 37424
rect -1374 37390 -1340 37424
rect -1306 37390 -1272 37424
rect -1238 37390 -1204 37424
rect -1170 37390 -1136 37424
rect -1102 37390 -1068 37424
rect -1034 37390 -1000 37424
rect -966 37390 -932 37424
rect -898 37390 -864 37424
rect -830 37390 -796 37424
rect -762 37390 -728 37424
rect -694 37390 -660 37424
rect -626 37390 -592 37424
rect -558 37390 -524 37424
rect -490 37390 -456 37424
rect -422 37390 -388 37424
rect -354 37390 -320 37424
rect -286 37390 -252 37424
rect -218 37390 -184 37424
rect -2938 37321 -2904 37355
rect -2870 37321 -2836 37355
rect -2802 37321 -2768 37355
rect -2734 37321 -2700 37355
rect -2666 37321 -2632 37355
rect -2598 37321 -2564 37355
rect -2530 37321 -2496 37355
rect -2462 37321 -2428 37355
rect -2394 37321 -2360 37355
rect -2326 37321 -2292 37355
rect -2258 37321 -2224 37355
rect -2190 37321 -2156 37355
rect -2122 37321 -2088 37355
rect -2054 37321 -2020 37355
rect -1986 37321 -1952 37355
rect -1918 37321 -1884 37355
rect -1850 37321 -1816 37355
rect -1782 37321 -1748 37355
rect -1714 37321 -1680 37355
rect -1646 37321 -1612 37355
rect -1578 37321 -1544 37355
rect -1510 37321 -1476 37355
rect -1442 37321 -1408 37355
rect -1374 37321 -1340 37355
rect -1306 37321 -1272 37355
rect -1238 37321 -1204 37355
rect -1170 37321 -1136 37355
rect -1102 37321 -1068 37355
rect -1034 37321 -1000 37355
rect -966 37321 -932 37355
rect -898 37321 -864 37355
rect -830 37321 -796 37355
rect -762 37321 -728 37355
rect -694 37321 -660 37355
rect -626 37321 -592 37355
rect -558 37321 -524 37355
rect -490 37321 -456 37355
rect -422 37321 -388 37355
rect -354 37321 -320 37355
rect -286 37321 -252 37355
rect -218 37321 -184 37355
rect -2938 37252 -2904 37286
rect -2870 37252 -2836 37286
rect -2802 37252 -2768 37286
rect -2734 37252 -2700 37286
rect -2666 37252 -2632 37286
rect -2598 37252 -2564 37286
rect -2530 37252 -2496 37286
rect -2462 37252 -2428 37286
rect -2394 37252 -2360 37286
rect -2326 37252 -2292 37286
rect -2258 37252 -2224 37286
rect -2190 37252 -2156 37286
rect -2122 37252 -2088 37286
rect -2054 37252 -2020 37286
rect -1986 37252 -1952 37286
rect -1918 37252 -1884 37286
rect -1850 37252 -1816 37286
rect -1782 37252 -1748 37286
rect -1714 37252 -1680 37286
rect -1646 37252 -1612 37286
rect -1578 37252 -1544 37286
rect -1510 37252 -1476 37286
rect -1442 37252 -1408 37286
rect -1374 37252 -1340 37286
rect -1306 37252 -1272 37286
rect -1238 37252 -1204 37286
rect -1170 37252 -1136 37286
rect -1102 37252 -1068 37286
rect -1034 37252 -1000 37286
rect -966 37252 -932 37286
rect -898 37252 -864 37286
rect -830 37252 -796 37286
rect -762 37252 -728 37286
rect -694 37252 -660 37286
rect -626 37252 -592 37286
rect -558 37252 -524 37286
rect -490 37252 -456 37286
rect -422 37252 -388 37286
rect -354 37252 -320 37286
rect -286 37252 -252 37286
rect -218 37252 -184 37286
rect -2938 37183 -2904 37217
rect -2870 37183 -2836 37217
rect -2802 37183 -2768 37217
rect -2734 37183 -2700 37217
rect -2666 37183 -2632 37217
rect -2598 37183 -2564 37217
rect -2530 37183 -2496 37217
rect -2462 37183 -2428 37217
rect -2394 37183 -2360 37217
rect -2326 37183 -2292 37217
rect -2258 37183 -2224 37217
rect -2190 37183 -2156 37217
rect -2122 37183 -2088 37217
rect -2054 37183 -2020 37217
rect -1986 37183 -1952 37217
rect -1918 37183 -1884 37217
rect -1850 37183 -1816 37217
rect -1782 37183 -1748 37217
rect -1714 37183 -1680 37217
rect -1646 37183 -1612 37217
rect -1578 37183 -1544 37217
rect -1510 37183 -1476 37217
rect -1442 37183 -1408 37217
rect -1374 37183 -1340 37217
rect -1306 37183 -1272 37217
rect -1238 37183 -1204 37217
rect -1170 37183 -1136 37217
rect -1102 37183 -1068 37217
rect -1034 37183 -1000 37217
rect -966 37183 -932 37217
rect -898 37183 -864 37217
rect -830 37183 -796 37217
rect -762 37183 -728 37217
rect -694 37183 -660 37217
rect -626 37183 -592 37217
rect -558 37183 -524 37217
rect -490 37183 -456 37217
rect -422 37183 -388 37217
rect -354 37183 -320 37217
rect -286 37183 -252 37217
rect -218 37183 -184 37217
rect -2938 37114 -2904 37148
rect -2870 37114 -2836 37148
rect -2802 37114 -2768 37148
rect -2734 37114 -2700 37148
rect -2666 37114 -2632 37148
rect -2598 37114 -2564 37148
rect -2530 37114 -2496 37148
rect -2462 37114 -2428 37148
rect -2394 37114 -2360 37148
rect -2326 37114 -2292 37148
rect -2258 37114 -2224 37148
rect -2190 37114 -2156 37148
rect -2122 37114 -2088 37148
rect -2054 37114 -2020 37148
rect -1986 37114 -1952 37148
rect -1918 37114 -1884 37148
rect -1850 37114 -1816 37148
rect -1782 37114 -1748 37148
rect -1714 37114 -1680 37148
rect -1646 37114 -1612 37148
rect -1578 37114 -1544 37148
rect -1510 37114 -1476 37148
rect -1442 37114 -1408 37148
rect -1374 37114 -1340 37148
rect -1306 37114 -1272 37148
rect -1238 37114 -1204 37148
rect -1170 37114 -1136 37148
rect -1102 37114 -1068 37148
rect -1034 37114 -1000 37148
rect -966 37114 -932 37148
rect -898 37114 -864 37148
rect -830 37114 -796 37148
rect -762 37114 -728 37148
rect -694 37114 -660 37148
rect -626 37114 -592 37148
rect -558 37114 -524 37148
rect -490 37114 -456 37148
rect -422 37114 -388 37148
rect -354 37114 -320 37148
rect -286 37114 -252 37148
rect -218 37114 -184 37148
rect -2938 37045 -2904 37079
rect -2870 37045 -2836 37079
rect -2802 37045 -2768 37079
rect -2734 37045 -2700 37079
rect -2666 37045 -2632 37079
rect -2598 37045 -2564 37079
rect -2530 37045 -2496 37079
rect -2462 37045 -2428 37079
rect -2394 37045 -2360 37079
rect -2326 37045 -2292 37079
rect -2258 37045 -2224 37079
rect -2190 37045 -2156 37079
rect -2122 37045 -2088 37079
rect -2054 37045 -2020 37079
rect -1986 37045 -1952 37079
rect -1918 37045 -1884 37079
rect -1850 37045 -1816 37079
rect -1782 37045 -1748 37079
rect -1714 37045 -1680 37079
rect -1646 37045 -1612 37079
rect -1578 37045 -1544 37079
rect -1510 37045 -1476 37079
rect -1442 37045 -1408 37079
rect -1374 37045 -1340 37079
rect -1306 37045 -1272 37079
rect -1238 37045 -1204 37079
rect -1170 37045 -1136 37079
rect -1102 37045 -1068 37079
rect -1034 37045 -1000 37079
rect -966 37045 -932 37079
rect -898 37045 -864 37079
rect -830 37045 -796 37079
rect -762 37045 -728 37079
rect -694 37045 -660 37079
rect -626 37045 -592 37079
rect -558 37045 -524 37079
rect -490 37045 -456 37079
rect -422 37045 -388 37079
rect -354 37045 -320 37079
rect -286 37045 -252 37079
rect -218 37045 -184 37079
rect -2938 36976 -2904 37010
rect -2870 36976 -2836 37010
rect -2802 36976 -2768 37010
rect -2734 36976 -2700 37010
rect -2666 36976 -2632 37010
rect -2598 36976 -2564 37010
rect -2530 36976 -2496 37010
rect -2462 36976 -2428 37010
rect -2394 36976 -2360 37010
rect -2326 36976 -2292 37010
rect -2258 36976 -2224 37010
rect -2190 36976 -2156 37010
rect -2122 36976 -2088 37010
rect -2054 36976 -2020 37010
rect -1986 36976 -1952 37010
rect -1918 36976 -1884 37010
rect -1850 36976 -1816 37010
rect -1782 36976 -1748 37010
rect -1714 36976 -1680 37010
rect -1646 36976 -1612 37010
rect -1578 36976 -1544 37010
rect -1510 36976 -1476 37010
rect -1442 36976 -1408 37010
rect -1374 36976 -1340 37010
rect -1306 36976 -1272 37010
rect -1238 36976 -1204 37010
rect -1170 36976 -1136 37010
rect -1102 36976 -1068 37010
rect -1034 36976 -1000 37010
rect -966 36976 -932 37010
rect -898 36976 -864 37010
rect -830 36976 -796 37010
rect -762 36976 -728 37010
rect -694 36976 -660 37010
rect -626 36976 -592 37010
rect -558 36976 -524 37010
rect -490 36976 -456 37010
rect -422 36976 -388 37010
rect -354 36976 -320 37010
rect -286 36976 -252 37010
rect -218 36976 -184 37010
rect -2938 36907 -2904 36941
rect -2870 36907 -2836 36941
rect -2802 36907 -2768 36941
rect -2734 36907 -2700 36941
rect -2666 36907 -2632 36941
rect -2598 36907 -2564 36941
rect -2530 36907 -2496 36941
rect -2462 36907 -2428 36941
rect -2394 36907 -2360 36941
rect -2326 36907 -2292 36941
rect -2258 36907 -2224 36941
rect -2190 36907 -2156 36941
rect -2122 36907 -2088 36941
rect -2054 36907 -2020 36941
rect -1986 36907 -1952 36941
rect -1918 36907 -1884 36941
rect -1850 36907 -1816 36941
rect -1782 36907 -1748 36941
rect -1714 36907 -1680 36941
rect -1646 36907 -1612 36941
rect -1578 36907 -1544 36941
rect -1510 36907 -1476 36941
rect -1442 36907 -1408 36941
rect -1374 36907 -1340 36941
rect -1306 36907 -1272 36941
rect -1238 36907 -1204 36941
rect -1170 36907 -1136 36941
rect -1102 36907 -1068 36941
rect -1034 36907 -1000 36941
rect -966 36907 -932 36941
rect -898 36907 -864 36941
rect -830 36907 -796 36941
rect -762 36907 -728 36941
rect -694 36907 -660 36941
rect -626 36907 -592 36941
rect -558 36907 -524 36941
rect -490 36907 -456 36941
rect -422 36907 -388 36941
rect -354 36907 -320 36941
rect -286 36907 -252 36941
rect -218 36907 -184 36941
rect -2938 36838 -2904 36872
rect -2870 36838 -2836 36872
rect -2802 36838 -2768 36872
rect -2734 36838 -2700 36872
rect -2666 36838 -2632 36872
rect -2598 36838 -2564 36872
rect -2530 36838 -2496 36872
rect -2462 36838 -2428 36872
rect -2394 36838 -2360 36872
rect -2326 36838 -2292 36872
rect -2258 36838 -2224 36872
rect -2190 36838 -2156 36872
rect -2122 36838 -2088 36872
rect -2054 36838 -2020 36872
rect -1986 36838 -1952 36872
rect -1918 36838 -1884 36872
rect -1850 36838 -1816 36872
rect -1782 36838 -1748 36872
rect -1714 36838 -1680 36872
rect -1646 36838 -1612 36872
rect -1578 36838 -1544 36872
rect -1510 36838 -1476 36872
rect -1442 36838 -1408 36872
rect -1374 36838 -1340 36872
rect -1306 36838 -1272 36872
rect -1238 36838 -1204 36872
rect -1170 36838 -1136 36872
rect -1102 36838 -1068 36872
rect -1034 36838 -1000 36872
rect -966 36838 -932 36872
rect -898 36838 -864 36872
rect -830 36838 -796 36872
rect -762 36838 -728 36872
rect -694 36838 -660 36872
rect -626 36838 -592 36872
rect -558 36838 -524 36872
rect -490 36838 -456 36872
rect -422 36838 -388 36872
rect -354 36838 -320 36872
rect -286 36838 -252 36872
rect -218 36838 -184 36872
rect -2938 36769 -2904 36803
rect -2870 36769 -2836 36803
rect -2802 36769 -2768 36803
rect -2734 36769 -2700 36803
rect -2666 36769 -2632 36803
rect -2598 36769 -2564 36803
rect -2530 36769 -2496 36803
rect -2462 36769 -2428 36803
rect -2394 36769 -2360 36803
rect -2326 36769 -2292 36803
rect -2258 36769 -2224 36803
rect -2190 36769 -2156 36803
rect -2122 36769 -2088 36803
rect -2054 36769 -2020 36803
rect -1986 36769 -1952 36803
rect -1918 36769 -1884 36803
rect -1850 36769 -1816 36803
rect -1782 36769 -1748 36803
rect -1714 36769 -1680 36803
rect -1646 36769 -1612 36803
rect -1578 36769 -1544 36803
rect -1510 36769 -1476 36803
rect -1442 36769 -1408 36803
rect -1374 36769 -1340 36803
rect -1306 36769 -1272 36803
rect -1238 36769 -1204 36803
rect -1170 36769 -1136 36803
rect -1102 36769 -1068 36803
rect -1034 36769 -1000 36803
rect -966 36769 -932 36803
rect -898 36769 -864 36803
rect -830 36769 -796 36803
rect -762 36769 -728 36803
rect -694 36769 -660 36803
rect -626 36769 -592 36803
rect -558 36769 -524 36803
rect -490 36769 -456 36803
rect -422 36769 -388 36803
rect -354 36769 -320 36803
rect -286 36769 -252 36803
rect -218 36769 -184 36803
rect -2938 36700 -2904 36734
rect -2870 36700 -2836 36734
rect -2802 36700 -2768 36734
rect -2734 36700 -2700 36734
rect -2666 36700 -2632 36734
rect -2598 36700 -2564 36734
rect -2530 36700 -2496 36734
rect -2462 36700 -2428 36734
rect -2394 36700 -2360 36734
rect -2326 36700 -2292 36734
rect -2258 36700 -2224 36734
rect -2190 36700 -2156 36734
rect -2122 36700 -2088 36734
rect -2054 36700 -2020 36734
rect -1986 36700 -1952 36734
rect -1918 36700 -1884 36734
rect -1850 36700 -1816 36734
rect -1782 36700 -1748 36734
rect -1714 36700 -1680 36734
rect -1646 36700 -1612 36734
rect -1578 36700 -1544 36734
rect -1510 36700 -1476 36734
rect -1442 36700 -1408 36734
rect -1374 36700 -1340 36734
rect -1306 36700 -1272 36734
rect -1238 36700 -1204 36734
rect -1170 36700 -1136 36734
rect -1102 36700 -1068 36734
rect -1034 36700 -1000 36734
rect -966 36700 -932 36734
rect -898 36700 -864 36734
rect -830 36700 -796 36734
rect -762 36700 -728 36734
rect -694 36700 -660 36734
rect -626 36700 -592 36734
rect -558 36700 -524 36734
rect -490 36700 -456 36734
rect -422 36700 -388 36734
rect -354 36700 -320 36734
rect -286 36700 -252 36734
rect -218 36700 -184 36734
rect -2938 36631 -2904 36665
rect -2870 36631 -2836 36665
rect -2802 36631 -2768 36665
rect -2734 36631 -2700 36665
rect -2666 36631 -2632 36665
rect -2598 36631 -2564 36665
rect -2530 36631 -2496 36665
rect -2462 36631 -2428 36665
rect -2394 36631 -2360 36665
rect -2326 36631 -2292 36665
rect -2258 36631 -2224 36665
rect -2190 36631 -2156 36665
rect -2122 36631 -2088 36665
rect -2054 36631 -2020 36665
rect -1986 36631 -1952 36665
rect -1918 36631 -1884 36665
rect -1850 36631 -1816 36665
rect -1782 36631 -1748 36665
rect -1714 36631 -1680 36665
rect -1646 36631 -1612 36665
rect -1578 36631 -1544 36665
rect -1510 36631 -1476 36665
rect -1442 36631 -1408 36665
rect -1374 36631 -1340 36665
rect -1306 36631 -1272 36665
rect -1238 36631 -1204 36665
rect -1170 36631 -1136 36665
rect -1102 36631 -1068 36665
rect -1034 36631 -1000 36665
rect -966 36631 -932 36665
rect -898 36631 -864 36665
rect -830 36631 -796 36665
rect -762 36631 -728 36665
rect -694 36631 -660 36665
rect -626 36631 -592 36665
rect -558 36631 -524 36665
rect -490 36631 -456 36665
rect -422 36631 -388 36665
rect -354 36631 -320 36665
rect -286 36631 -252 36665
rect -218 36631 -184 36665
rect -2938 36562 -2904 36596
rect -2870 36562 -2836 36596
rect -2802 36562 -2768 36596
rect -2734 36562 -2700 36596
rect -2666 36562 -2632 36596
rect -2598 36562 -2564 36596
rect -2530 36562 -2496 36596
rect -2462 36562 -2428 36596
rect -2394 36562 -2360 36596
rect -2326 36562 -2292 36596
rect -2258 36562 -2224 36596
rect -2190 36562 -2156 36596
rect -2122 36562 -2088 36596
rect -2054 36562 -2020 36596
rect -1986 36562 -1952 36596
rect -1918 36562 -1884 36596
rect -1850 36562 -1816 36596
rect -1782 36562 -1748 36596
rect -1714 36562 -1680 36596
rect -1646 36562 -1612 36596
rect -1578 36562 -1544 36596
rect -1510 36562 -1476 36596
rect -1442 36562 -1408 36596
rect -1374 36562 -1340 36596
rect -1306 36562 -1272 36596
rect -1238 36562 -1204 36596
rect -1170 36562 -1136 36596
rect -1102 36562 -1068 36596
rect -1034 36562 -1000 36596
rect -966 36562 -932 36596
rect -898 36562 -864 36596
rect -830 36562 -796 36596
rect -762 36562 -728 36596
rect -694 36562 -660 36596
rect -626 36562 -592 36596
rect -558 36562 -524 36596
rect -490 36562 -456 36596
rect -422 36562 -388 36596
rect -354 36562 -320 36596
rect -286 36562 -252 36596
rect -218 36562 -184 36596
rect -2938 36493 -2904 36527
rect -2870 36493 -2836 36527
rect -2802 36493 -2768 36527
rect -2734 36493 -2700 36527
rect -2666 36493 -2632 36527
rect -2598 36493 -2564 36527
rect -2530 36493 -2496 36527
rect -2462 36493 -2428 36527
rect -2394 36493 -2360 36527
rect -2326 36493 -2292 36527
rect -2258 36493 -2224 36527
rect -2190 36493 -2156 36527
rect -2122 36493 -2088 36527
rect -2054 36493 -2020 36527
rect -1986 36493 -1952 36527
rect -1918 36493 -1884 36527
rect -1850 36493 -1816 36527
rect -1782 36493 -1748 36527
rect -1714 36493 -1680 36527
rect -1646 36493 -1612 36527
rect -1578 36493 -1544 36527
rect -1510 36493 -1476 36527
rect -1442 36493 -1408 36527
rect -1374 36493 -1340 36527
rect -1306 36493 -1272 36527
rect -1238 36493 -1204 36527
rect -1170 36493 -1136 36527
rect -1102 36493 -1068 36527
rect -1034 36493 -1000 36527
rect -966 36493 -932 36527
rect -898 36493 -864 36527
rect -830 36493 -796 36527
rect -762 36493 -728 36527
rect -694 36493 -660 36527
rect -626 36493 -592 36527
rect -558 36493 -524 36527
rect -490 36493 -456 36527
rect -422 36493 -388 36527
rect -354 36493 -320 36527
rect -286 36493 -252 36527
rect -218 36493 -184 36527
rect -2938 36424 -2904 36458
rect -2870 36424 -2836 36458
rect -2802 36424 -2768 36458
rect -2734 36424 -2700 36458
rect -2666 36424 -2632 36458
rect -2598 36424 -2564 36458
rect -2530 36424 -2496 36458
rect -2462 36424 -2428 36458
rect -2394 36424 -2360 36458
rect -2326 36424 -2292 36458
rect -2258 36424 -2224 36458
rect -2190 36424 -2156 36458
rect -2122 36424 -2088 36458
rect -2054 36424 -2020 36458
rect -1986 36424 -1952 36458
rect -1918 36424 -1884 36458
rect -1850 36424 -1816 36458
rect -1782 36424 -1748 36458
rect -1714 36424 -1680 36458
rect -1646 36424 -1612 36458
rect -1578 36424 -1544 36458
rect -1510 36424 -1476 36458
rect -1442 36424 -1408 36458
rect -1374 36424 -1340 36458
rect -1306 36424 -1272 36458
rect -1238 36424 -1204 36458
rect -1170 36424 -1136 36458
rect -1102 36424 -1068 36458
rect -1034 36424 -1000 36458
rect -966 36424 -932 36458
rect -898 36424 -864 36458
rect -830 36424 -796 36458
rect -762 36424 -728 36458
rect -694 36424 -660 36458
rect -626 36424 -592 36458
rect -558 36424 -524 36458
rect -490 36424 -456 36458
rect -422 36424 -388 36458
rect -354 36424 -320 36458
rect -286 36424 -252 36458
rect -218 36424 -184 36458
rect -2938 36355 -2904 36389
rect -2870 36355 -2836 36389
rect -2802 36355 -2768 36389
rect -2734 36355 -2700 36389
rect -2666 36355 -2632 36389
rect -2598 36355 -2564 36389
rect -2530 36355 -2496 36389
rect -2462 36355 -2428 36389
rect -2394 36355 -2360 36389
rect -2326 36355 -2292 36389
rect -2258 36355 -2224 36389
rect -2190 36355 -2156 36389
rect -2122 36355 -2088 36389
rect -2054 36355 -2020 36389
rect -1986 36355 -1952 36389
rect -1918 36355 -1884 36389
rect -1850 36355 -1816 36389
rect -1782 36355 -1748 36389
rect -1714 36355 -1680 36389
rect -1646 36355 -1612 36389
rect -1578 36355 -1544 36389
rect -1510 36355 -1476 36389
rect -1442 36355 -1408 36389
rect -1374 36355 -1340 36389
rect -1306 36355 -1272 36389
rect -1238 36355 -1204 36389
rect -1170 36355 -1136 36389
rect -1102 36355 -1068 36389
rect -1034 36355 -1000 36389
rect -966 36355 -932 36389
rect -898 36355 -864 36389
rect -830 36355 -796 36389
rect -762 36355 -728 36389
rect -694 36355 -660 36389
rect -626 36355 -592 36389
rect -558 36355 -524 36389
rect -490 36355 -456 36389
rect -422 36355 -388 36389
rect -354 36355 -320 36389
rect -286 36355 -252 36389
rect -218 36355 -184 36389
rect -2938 36286 -2904 36320
rect -2870 36286 -2836 36320
rect -2802 36286 -2768 36320
rect -2734 36286 -2700 36320
rect -2666 36286 -2632 36320
rect -2598 36286 -2564 36320
rect -2530 36286 -2496 36320
rect -2462 36286 -2428 36320
rect -2394 36286 -2360 36320
rect -2326 36286 -2292 36320
rect -2258 36286 -2224 36320
rect -2190 36286 -2156 36320
rect -2122 36286 -2088 36320
rect -2054 36286 -2020 36320
rect -1986 36286 -1952 36320
rect -1918 36286 -1884 36320
rect -1850 36286 -1816 36320
rect -1782 36286 -1748 36320
rect -1714 36286 -1680 36320
rect -1646 36286 -1612 36320
rect -1578 36286 -1544 36320
rect -1510 36286 -1476 36320
rect -1442 36286 -1408 36320
rect -1374 36286 -1340 36320
rect -1306 36286 -1272 36320
rect -1238 36286 -1204 36320
rect -1170 36286 -1136 36320
rect -1102 36286 -1068 36320
rect -1034 36286 -1000 36320
rect -966 36286 -932 36320
rect -898 36286 -864 36320
rect -830 36286 -796 36320
rect -762 36286 -728 36320
rect -694 36286 -660 36320
rect -626 36286 -592 36320
rect -558 36286 -524 36320
rect -490 36286 -456 36320
rect -422 36286 -388 36320
rect -354 36286 -320 36320
rect -286 36286 -252 36320
rect -218 36286 -184 36320
rect -2938 36217 -2904 36251
rect -2870 36217 -2836 36251
rect -2802 36217 -2768 36251
rect -2734 36217 -2700 36251
rect -2666 36217 -2632 36251
rect -2598 36217 -2564 36251
rect -2530 36217 -2496 36251
rect -2462 36217 -2428 36251
rect -2394 36217 -2360 36251
rect -2326 36217 -2292 36251
rect -2258 36217 -2224 36251
rect -2190 36217 -2156 36251
rect -2122 36217 -2088 36251
rect -2054 36217 -2020 36251
rect -1986 36217 -1952 36251
rect -1918 36217 -1884 36251
rect -1850 36217 -1816 36251
rect -1782 36217 -1748 36251
rect -1714 36217 -1680 36251
rect -1646 36217 -1612 36251
rect -1578 36217 -1544 36251
rect -1510 36217 -1476 36251
rect -1442 36217 -1408 36251
rect -1374 36217 -1340 36251
rect -1306 36217 -1272 36251
rect -1238 36217 -1204 36251
rect -1170 36217 -1136 36251
rect -1102 36217 -1068 36251
rect -1034 36217 -1000 36251
rect -966 36217 -932 36251
rect -898 36217 -864 36251
rect -830 36217 -796 36251
rect -762 36217 -728 36251
rect -694 36217 -660 36251
rect -626 36217 -592 36251
rect -558 36217 -524 36251
rect -490 36217 -456 36251
rect -422 36217 -388 36251
rect -354 36217 -320 36251
rect -286 36217 -252 36251
rect -218 36217 -184 36251
rect -2938 36148 -2904 36182
rect -2870 36148 -2836 36182
rect -2802 36148 -2768 36182
rect -2734 36148 -2700 36182
rect -2666 36148 -2632 36182
rect -2598 36148 -2564 36182
rect -2530 36148 -2496 36182
rect -2462 36148 -2428 36182
rect -2394 36148 -2360 36182
rect -2326 36148 -2292 36182
rect -2258 36148 -2224 36182
rect -2190 36148 -2156 36182
rect -2122 36148 -2088 36182
rect -2054 36148 -2020 36182
rect -1986 36148 -1952 36182
rect -1918 36148 -1884 36182
rect -1850 36148 -1816 36182
rect -1782 36148 -1748 36182
rect -1714 36148 -1680 36182
rect -1646 36148 -1612 36182
rect -1578 36148 -1544 36182
rect -1510 36148 -1476 36182
rect -1442 36148 -1408 36182
rect -1374 36148 -1340 36182
rect -1306 36148 -1272 36182
rect -1238 36148 -1204 36182
rect -1170 36148 -1136 36182
rect -1102 36148 -1068 36182
rect -1034 36148 -1000 36182
rect -966 36148 -932 36182
rect -898 36148 -864 36182
rect -830 36148 -796 36182
rect -762 36148 -728 36182
rect -694 36148 -660 36182
rect -626 36148 -592 36182
rect -558 36148 -524 36182
rect -490 36148 -456 36182
rect -422 36148 -388 36182
rect -354 36148 -320 36182
rect -286 36148 -252 36182
rect -218 36148 -184 36182
rect -2938 36079 -2904 36113
rect -2870 36079 -2836 36113
rect -2802 36079 -2768 36113
rect -2734 36079 -2700 36113
rect -2666 36079 -2632 36113
rect -2598 36079 -2564 36113
rect -2530 36079 -2496 36113
rect -2462 36079 -2428 36113
rect -2394 36079 -2360 36113
rect -2326 36079 -2292 36113
rect -2258 36079 -2224 36113
rect -2190 36079 -2156 36113
rect -2122 36079 -2088 36113
rect -2054 36079 -2020 36113
rect -1986 36079 -1952 36113
rect -1918 36079 -1884 36113
rect -1850 36079 -1816 36113
rect -1782 36079 -1748 36113
rect -1714 36079 -1680 36113
rect -1646 36079 -1612 36113
rect -1578 36079 -1544 36113
rect -1510 36079 -1476 36113
rect -1442 36079 -1408 36113
rect -1374 36079 -1340 36113
rect -1306 36079 -1272 36113
rect -1238 36079 -1204 36113
rect -1170 36079 -1136 36113
rect -1102 36079 -1068 36113
rect -1034 36079 -1000 36113
rect -966 36079 -932 36113
rect -898 36079 -864 36113
rect -830 36079 -796 36113
rect -762 36079 -728 36113
rect -694 36079 -660 36113
rect -626 36079 -592 36113
rect -558 36079 -524 36113
rect -490 36079 -456 36113
rect -422 36079 -388 36113
rect -354 36079 -320 36113
rect -286 36079 -252 36113
rect -218 36079 -184 36113
rect -2938 36010 -2904 36044
rect -2870 36010 -2836 36044
rect -2802 36010 -2768 36044
rect -2734 36010 -2700 36044
rect -2666 36010 -2632 36044
rect -2598 36010 -2564 36044
rect -2530 36010 -2496 36044
rect -2462 36010 -2428 36044
rect -2394 36010 -2360 36044
rect -2326 36010 -2292 36044
rect -2258 36010 -2224 36044
rect -2190 36010 -2156 36044
rect -2122 36010 -2088 36044
rect -2054 36010 -2020 36044
rect -1986 36010 -1952 36044
rect -1918 36010 -1884 36044
rect -1850 36010 -1816 36044
rect -1782 36010 -1748 36044
rect -1714 36010 -1680 36044
rect -1646 36010 -1612 36044
rect -1578 36010 -1544 36044
rect -1510 36010 -1476 36044
rect -1442 36010 -1408 36044
rect -1374 36010 -1340 36044
rect -1306 36010 -1272 36044
rect -1238 36010 -1204 36044
rect -1170 36010 -1136 36044
rect -1102 36010 -1068 36044
rect -1034 36010 -1000 36044
rect -966 36010 -932 36044
rect -898 36010 -864 36044
rect -830 36010 -796 36044
rect -762 36010 -728 36044
rect -694 36010 -660 36044
rect -626 36010 -592 36044
rect -558 36010 -524 36044
rect -490 36010 -456 36044
rect -422 36010 -388 36044
rect -354 36010 -320 36044
rect -286 36010 -252 36044
rect -218 36010 -184 36044
rect -2938 35941 -2904 35975
rect -2870 35941 -2836 35975
rect -2802 35941 -2768 35975
rect -2734 35941 -2700 35975
rect -2666 35941 -2632 35975
rect -2598 35941 -2564 35975
rect -2530 35941 -2496 35975
rect -2462 35941 -2428 35975
rect -2394 35941 -2360 35975
rect -2326 35941 -2292 35975
rect -2258 35941 -2224 35975
rect -2190 35941 -2156 35975
rect -2122 35941 -2088 35975
rect -2054 35941 -2020 35975
rect -1986 35941 -1952 35975
rect -1918 35941 -1884 35975
rect -1850 35941 -1816 35975
rect -1782 35941 -1748 35975
rect -1714 35941 -1680 35975
rect -1646 35941 -1612 35975
rect -1578 35941 -1544 35975
rect -1510 35941 -1476 35975
rect -1442 35941 -1408 35975
rect -1374 35941 -1340 35975
rect -1306 35941 -1272 35975
rect -1238 35941 -1204 35975
rect -1170 35941 -1136 35975
rect -1102 35941 -1068 35975
rect -1034 35941 -1000 35975
rect -966 35941 -932 35975
rect -898 35941 -864 35975
rect -830 35941 -796 35975
rect -762 35941 -728 35975
rect -694 35941 -660 35975
rect -626 35941 -592 35975
rect -558 35941 -524 35975
rect -490 35941 -456 35975
rect -422 35941 -388 35975
rect -354 35941 -320 35975
rect -286 35941 -252 35975
rect -218 35941 -184 35975
rect -2938 35872 -2904 35906
rect -2870 35872 -2836 35906
rect -2802 35872 -2768 35906
rect -2734 35872 -2700 35906
rect -2666 35872 -2632 35906
rect -2598 35872 -2564 35906
rect -2530 35872 -2496 35906
rect -2462 35872 -2428 35906
rect -2394 35872 -2360 35906
rect -2326 35872 -2292 35906
rect -2258 35872 -2224 35906
rect -2190 35872 -2156 35906
rect -2122 35872 -2088 35906
rect -2054 35872 -2020 35906
rect -1986 35872 -1952 35906
rect -1918 35872 -1884 35906
rect -1850 35872 -1816 35906
rect -1782 35872 -1748 35906
rect -1714 35872 -1680 35906
rect -1646 35872 -1612 35906
rect -1578 35872 -1544 35906
rect -1510 35872 -1476 35906
rect -1442 35872 -1408 35906
rect -1374 35872 -1340 35906
rect -1306 35872 -1272 35906
rect -1238 35872 -1204 35906
rect -1170 35872 -1136 35906
rect -1102 35872 -1068 35906
rect -1034 35872 -1000 35906
rect -966 35872 -932 35906
rect -898 35872 -864 35906
rect -830 35872 -796 35906
rect -762 35872 -728 35906
rect -694 35872 -660 35906
rect -626 35872 -592 35906
rect -558 35872 -524 35906
rect -490 35872 -456 35906
rect -422 35872 -388 35906
rect -354 35872 -320 35906
rect -286 35872 -252 35906
rect -218 35872 -184 35906
rect -2938 35803 -2904 35837
rect -2870 35803 -2836 35837
rect -2802 35803 -2768 35837
rect -2734 35803 -2700 35837
rect -2666 35803 -2632 35837
rect -2598 35803 -2564 35837
rect -2530 35803 -2496 35837
rect -2462 35803 -2428 35837
rect -2394 35803 -2360 35837
rect -2326 35803 -2292 35837
rect -2258 35803 -2224 35837
rect -2190 35803 -2156 35837
rect -2122 35803 -2088 35837
rect -2054 35803 -2020 35837
rect -1986 35803 -1952 35837
rect -1918 35803 -1884 35837
rect -1850 35803 -1816 35837
rect -1782 35803 -1748 35837
rect -1714 35803 -1680 35837
rect -1646 35803 -1612 35837
rect -1578 35803 -1544 35837
rect -1510 35803 -1476 35837
rect -1442 35803 -1408 35837
rect -1374 35803 -1340 35837
rect -1306 35803 -1272 35837
rect -1238 35803 -1204 35837
rect -1170 35803 -1136 35837
rect -1102 35803 -1068 35837
rect -1034 35803 -1000 35837
rect -966 35803 -932 35837
rect -898 35803 -864 35837
rect -830 35803 -796 35837
rect -762 35803 -728 35837
rect -694 35803 -660 35837
rect -626 35803 -592 35837
rect -558 35803 -524 35837
rect -490 35803 -456 35837
rect -422 35803 -388 35837
rect -354 35803 -320 35837
rect -286 35803 -252 35837
rect -218 35803 -184 35837
rect -2938 35734 -2904 35768
rect -2870 35734 -2836 35768
rect -2802 35734 -2768 35768
rect -2734 35734 -2700 35768
rect -2666 35734 -2632 35768
rect -2598 35734 -2564 35768
rect -2530 35734 -2496 35768
rect -2462 35734 -2428 35768
rect -2394 35734 -2360 35768
rect -2326 35734 -2292 35768
rect -2258 35734 -2224 35768
rect -2190 35734 -2156 35768
rect -2122 35734 -2088 35768
rect -2054 35734 -2020 35768
rect -1986 35734 -1952 35768
rect -1918 35734 -1884 35768
rect -1850 35734 -1816 35768
rect -1782 35734 -1748 35768
rect -1714 35734 -1680 35768
rect -1646 35734 -1612 35768
rect -1578 35734 -1544 35768
rect -1510 35734 -1476 35768
rect -1442 35734 -1408 35768
rect -1374 35734 -1340 35768
rect -1306 35734 -1272 35768
rect -1238 35734 -1204 35768
rect -1170 35734 -1136 35768
rect -1102 35734 -1068 35768
rect -1034 35734 -1000 35768
rect -966 35734 -932 35768
rect -898 35734 -864 35768
rect -830 35734 -796 35768
rect -762 35734 -728 35768
rect -694 35734 -660 35768
rect -626 35734 -592 35768
rect -558 35734 -524 35768
rect -490 35734 -456 35768
rect -422 35734 -388 35768
rect -354 35734 -320 35768
rect -286 35734 -252 35768
rect -218 35734 -184 35768
rect -2938 35665 -2904 35699
rect -2870 35665 -2836 35699
rect -2802 35665 -2768 35699
rect -2734 35665 -2700 35699
rect -2666 35665 -2632 35699
rect -2598 35665 -2564 35699
rect -2530 35665 -2496 35699
rect -2462 35665 -2428 35699
rect -2394 35665 -2360 35699
rect -2326 35665 -2292 35699
rect -2258 35665 -2224 35699
rect -2190 35665 -2156 35699
rect -2122 35665 -2088 35699
rect -2054 35665 -2020 35699
rect -1986 35665 -1952 35699
rect -1918 35665 -1884 35699
rect -1850 35665 -1816 35699
rect -1782 35665 -1748 35699
rect -1714 35665 -1680 35699
rect -1646 35665 -1612 35699
rect -1578 35665 -1544 35699
rect -1510 35665 -1476 35699
rect -1442 35665 -1408 35699
rect -1374 35665 -1340 35699
rect -1306 35665 -1272 35699
rect -1238 35665 -1204 35699
rect -1170 35665 -1136 35699
rect -1102 35665 -1068 35699
rect -1034 35665 -1000 35699
rect -966 35665 -932 35699
rect -898 35665 -864 35699
rect -830 35665 -796 35699
rect -762 35665 -728 35699
rect -694 35665 -660 35699
rect -626 35665 -592 35699
rect -558 35665 -524 35699
rect -490 35665 -456 35699
rect -422 35665 -388 35699
rect -354 35665 -320 35699
rect -286 35665 -252 35699
rect -218 35665 -184 35699
rect -2938 35596 -2904 35630
rect -2870 35596 -2836 35630
rect -2802 35596 -2768 35630
rect -2734 35596 -2700 35630
rect -2666 35596 -2632 35630
rect -2598 35596 -2564 35630
rect -2530 35596 -2496 35630
rect -2462 35596 -2428 35630
rect -2394 35596 -2360 35630
rect -2326 35596 -2292 35630
rect -2258 35596 -2224 35630
rect -2190 35596 -2156 35630
rect -2122 35596 -2088 35630
rect -2054 35596 -2020 35630
rect -1986 35596 -1952 35630
rect -1918 35596 -1884 35630
rect -1850 35596 -1816 35630
rect -1782 35596 -1748 35630
rect -1714 35596 -1680 35630
rect -1646 35596 -1612 35630
rect -1578 35596 -1544 35630
rect -1510 35596 -1476 35630
rect -1442 35596 -1408 35630
rect -1374 35596 -1340 35630
rect -1306 35596 -1272 35630
rect -1238 35596 -1204 35630
rect -1170 35596 -1136 35630
rect -1102 35596 -1068 35630
rect -1034 35596 -1000 35630
rect -966 35596 -932 35630
rect -898 35596 -864 35630
rect -830 35596 -796 35630
rect -762 35596 -728 35630
rect -694 35596 -660 35630
rect -626 35596 -592 35630
rect -558 35596 -524 35630
rect -490 35596 -456 35630
rect -422 35596 -388 35630
rect -354 35596 -320 35630
rect -286 35596 -252 35630
rect -218 35596 -184 35630
rect -2938 35527 -2904 35561
rect -2870 35527 -2836 35561
rect -2802 35527 -2768 35561
rect -2734 35527 -2700 35561
rect -2666 35527 -2632 35561
rect -2598 35527 -2564 35561
rect -2530 35527 -2496 35561
rect -2462 35527 -2428 35561
rect -2394 35527 -2360 35561
rect -2326 35527 -2292 35561
rect -2258 35527 -2224 35561
rect -2190 35527 -2156 35561
rect -2122 35527 -2088 35561
rect -2054 35527 -2020 35561
rect -1986 35527 -1952 35561
rect -1918 35527 -1884 35561
rect -1850 35527 -1816 35561
rect -1782 35527 -1748 35561
rect -1714 35527 -1680 35561
rect -1646 35527 -1612 35561
rect -1578 35527 -1544 35561
rect -1510 35527 -1476 35561
rect -1442 35527 -1408 35561
rect -1374 35527 -1340 35561
rect -1306 35527 -1272 35561
rect -1238 35527 -1204 35561
rect -1170 35527 -1136 35561
rect -1102 35527 -1068 35561
rect -1034 35527 -1000 35561
rect -966 35527 -932 35561
rect -898 35527 -864 35561
rect -830 35527 -796 35561
rect -762 35527 -728 35561
rect -694 35527 -660 35561
rect -626 35527 -592 35561
rect -558 35527 -524 35561
rect -490 35527 -456 35561
rect -422 35527 -388 35561
rect -354 35527 -320 35561
rect -286 35527 -252 35561
rect -218 35527 -184 35561
rect -2938 35458 -2904 35492
rect -2870 35458 -2836 35492
rect -2802 35458 -2768 35492
rect -2734 35458 -2700 35492
rect -2666 35458 -2632 35492
rect -2598 35458 -2564 35492
rect -2530 35458 -2496 35492
rect -2462 35458 -2428 35492
rect -2394 35458 -2360 35492
rect -2326 35458 -2292 35492
rect -2258 35458 -2224 35492
rect -2190 35458 -2156 35492
rect -2122 35458 -2088 35492
rect -2054 35458 -2020 35492
rect -1986 35458 -1952 35492
rect -1918 35458 -1884 35492
rect -1850 35458 -1816 35492
rect -1782 35458 -1748 35492
rect -1714 35458 -1680 35492
rect -1646 35458 -1612 35492
rect -1578 35458 -1544 35492
rect -1510 35458 -1476 35492
rect -1442 35458 -1408 35492
rect -1374 35458 -1340 35492
rect -1306 35458 -1272 35492
rect -1238 35458 -1204 35492
rect -1170 35458 -1136 35492
rect -1102 35458 -1068 35492
rect -1034 35458 -1000 35492
rect -966 35458 -932 35492
rect -898 35458 -864 35492
rect -830 35458 -796 35492
rect -762 35458 -728 35492
rect -694 35458 -660 35492
rect -626 35458 -592 35492
rect -558 35458 -524 35492
rect -490 35458 -456 35492
rect -422 35458 -388 35492
rect -354 35458 -320 35492
rect -286 35458 -252 35492
rect -218 35458 -184 35492
rect -2938 35389 -2904 35423
rect -2870 35389 -2836 35423
rect -2802 35389 -2768 35423
rect -2734 35389 -2700 35423
rect -2666 35389 -2632 35423
rect -2598 35389 -2564 35423
rect -2530 35389 -2496 35423
rect -2462 35389 -2428 35423
rect -2394 35389 -2360 35423
rect -2326 35389 -2292 35423
rect -2258 35389 -2224 35423
rect -2190 35389 -2156 35423
rect -2122 35389 -2088 35423
rect -2054 35389 -2020 35423
rect -1986 35389 -1952 35423
rect -1918 35389 -1884 35423
rect -1850 35389 -1816 35423
rect -1782 35389 -1748 35423
rect -1714 35389 -1680 35423
rect -1646 35389 -1612 35423
rect -1578 35389 -1544 35423
rect -1510 35389 -1476 35423
rect -1442 35389 -1408 35423
rect -1374 35389 -1340 35423
rect -1306 35389 -1272 35423
rect -1238 35389 -1204 35423
rect -1170 35389 -1136 35423
rect -1102 35389 -1068 35423
rect -1034 35389 -1000 35423
rect -966 35389 -932 35423
rect -898 35389 -864 35423
rect -830 35389 -796 35423
rect -762 35389 -728 35423
rect -694 35389 -660 35423
rect -626 35389 -592 35423
rect -558 35389 -524 35423
rect -490 35389 -456 35423
rect -422 35389 -388 35423
rect -354 35389 -320 35423
rect -286 35389 -252 35423
rect -218 35389 -184 35423
rect -2938 35320 -2904 35354
rect -2870 35320 -2836 35354
rect -2802 35320 -2768 35354
rect -2734 35320 -2700 35354
rect -2666 35320 -2632 35354
rect -2598 35320 -2564 35354
rect -2530 35320 -2496 35354
rect -2462 35320 -2428 35354
rect -2394 35320 -2360 35354
rect -2326 35320 -2292 35354
rect -2258 35320 -2224 35354
rect -2190 35320 -2156 35354
rect -2122 35320 -2088 35354
rect -2054 35320 -2020 35354
rect -1986 35320 -1952 35354
rect -1918 35320 -1884 35354
rect -1850 35320 -1816 35354
rect -1782 35320 -1748 35354
rect -1714 35320 -1680 35354
rect -1646 35320 -1612 35354
rect -1578 35320 -1544 35354
rect -1510 35320 -1476 35354
rect -1442 35320 -1408 35354
rect -1374 35320 -1340 35354
rect -1306 35320 -1272 35354
rect -1238 35320 -1204 35354
rect -1170 35320 -1136 35354
rect -1102 35320 -1068 35354
rect -1034 35320 -1000 35354
rect -966 35320 -932 35354
rect -898 35320 -864 35354
rect -830 35320 -796 35354
rect -762 35320 -728 35354
rect -694 35320 -660 35354
rect -626 35320 -592 35354
rect -558 35320 -524 35354
rect -490 35320 -456 35354
rect -422 35320 -388 35354
rect -354 35320 -320 35354
rect -286 35320 -252 35354
rect -218 35320 -184 35354
rect -2938 35251 -2904 35285
rect -2870 35251 -2836 35285
rect -2802 35251 -2768 35285
rect -2734 35251 -2700 35285
rect -2666 35251 -2632 35285
rect -2598 35251 -2564 35285
rect -2530 35251 -2496 35285
rect -2462 35251 -2428 35285
rect -2394 35251 -2360 35285
rect -2326 35251 -2292 35285
rect -2258 35251 -2224 35285
rect -2190 35251 -2156 35285
rect -2122 35251 -2088 35285
rect -2054 35251 -2020 35285
rect -1986 35251 -1952 35285
rect -1918 35251 -1884 35285
rect -1850 35251 -1816 35285
rect -1782 35251 -1748 35285
rect -1714 35251 -1680 35285
rect -1646 35251 -1612 35285
rect -1578 35251 -1544 35285
rect -1510 35251 -1476 35285
rect -1442 35251 -1408 35285
rect -1374 35251 -1340 35285
rect -1306 35251 -1272 35285
rect -1238 35251 -1204 35285
rect -1170 35251 -1136 35285
rect -1102 35251 -1068 35285
rect -1034 35251 -1000 35285
rect -966 35251 -932 35285
rect -898 35251 -864 35285
rect -830 35251 -796 35285
rect -762 35251 -728 35285
rect -694 35251 -660 35285
rect -626 35251 -592 35285
rect -558 35251 -524 35285
rect -490 35251 -456 35285
rect -422 35251 -388 35285
rect -354 35251 -320 35285
rect -286 35251 -252 35285
rect -218 35251 -184 35285
rect -2938 35182 -2904 35216
rect -2870 35182 -2836 35216
rect -2802 35182 -2768 35216
rect -2734 35182 -2700 35216
rect -2666 35182 -2632 35216
rect -2598 35182 -2564 35216
rect -2530 35182 -2496 35216
rect -2462 35182 -2428 35216
rect -2394 35182 -2360 35216
rect -2326 35182 -2292 35216
rect -2258 35182 -2224 35216
rect -2190 35182 -2156 35216
rect -2122 35182 -2088 35216
rect -2054 35182 -2020 35216
rect -1986 35182 -1952 35216
rect -1918 35182 -1884 35216
rect -1850 35182 -1816 35216
rect -1782 35182 -1748 35216
rect -1714 35182 -1680 35216
rect -1646 35182 -1612 35216
rect -1578 35182 -1544 35216
rect -1510 35182 -1476 35216
rect -1442 35182 -1408 35216
rect -1374 35182 -1340 35216
rect -1306 35182 -1272 35216
rect -1238 35182 -1204 35216
rect -1170 35182 -1136 35216
rect -1102 35182 -1068 35216
rect -1034 35182 -1000 35216
rect -966 35182 -932 35216
rect -898 35182 -864 35216
rect -830 35182 -796 35216
rect -762 35182 -728 35216
rect -694 35182 -660 35216
rect -626 35182 -592 35216
rect -558 35182 -524 35216
rect -490 35182 -456 35216
rect -422 35182 -388 35216
rect -354 35182 -320 35216
rect -286 35182 -252 35216
rect -218 35182 -184 35216
rect -2938 35113 -2904 35147
rect -2870 35113 -2836 35147
rect -2802 35113 -2768 35147
rect -2734 35113 -2700 35147
rect -2666 35113 -2632 35147
rect -2598 35113 -2564 35147
rect -2530 35113 -2496 35147
rect -2462 35113 -2428 35147
rect -2394 35113 -2360 35147
rect -2326 35113 -2292 35147
rect -2258 35113 -2224 35147
rect -2190 35113 -2156 35147
rect -2122 35113 -2088 35147
rect -2054 35113 -2020 35147
rect -1986 35113 -1952 35147
rect -1918 35113 -1884 35147
rect -1850 35113 -1816 35147
rect -1782 35113 -1748 35147
rect -1714 35113 -1680 35147
rect -1646 35113 -1612 35147
rect -1578 35113 -1544 35147
rect -1510 35113 -1476 35147
rect -1442 35113 -1408 35147
rect -1374 35113 -1340 35147
rect -1306 35113 -1272 35147
rect -1238 35113 -1204 35147
rect -1170 35113 -1136 35147
rect -1102 35113 -1068 35147
rect -1034 35113 -1000 35147
rect -966 35113 -932 35147
rect -898 35113 -864 35147
rect -830 35113 -796 35147
rect -762 35113 -728 35147
rect -694 35113 -660 35147
rect -626 35113 -592 35147
rect -558 35113 -524 35147
rect -490 35113 -456 35147
rect -422 35113 -388 35147
rect -354 35113 -320 35147
rect -286 35113 -252 35147
rect -218 35113 -184 35147
rect -2938 35044 -2904 35078
rect -2870 35044 -2836 35078
rect -2802 35044 -2768 35078
rect -2734 35044 -2700 35078
rect -2666 35044 -2632 35078
rect -2598 35044 -2564 35078
rect -2530 35044 -2496 35078
rect -2462 35044 -2428 35078
rect -2394 35044 -2360 35078
rect -2326 35044 -2292 35078
rect -2258 35044 -2224 35078
rect -2190 35044 -2156 35078
rect -2122 35044 -2088 35078
rect -2054 35044 -2020 35078
rect -1986 35044 -1952 35078
rect -1918 35044 -1884 35078
rect -1850 35044 -1816 35078
rect -1782 35044 -1748 35078
rect -1714 35044 -1680 35078
rect -1646 35044 -1612 35078
rect -1578 35044 -1544 35078
rect -1510 35044 -1476 35078
rect -1442 35044 -1408 35078
rect -1374 35044 -1340 35078
rect -1306 35044 -1272 35078
rect -1238 35044 -1204 35078
rect -1170 35044 -1136 35078
rect -1102 35044 -1068 35078
rect -1034 35044 -1000 35078
rect -966 35044 -932 35078
rect -898 35044 -864 35078
rect -830 35044 -796 35078
rect -762 35044 -728 35078
rect -694 35044 -660 35078
rect -626 35044 -592 35078
rect -558 35044 -524 35078
rect -490 35044 -456 35078
rect -422 35044 -388 35078
rect -354 35044 -320 35078
rect -286 35044 -252 35078
rect -218 35044 -184 35078
rect -2959 10413 -273 17927
rect 18349 14447 18383 14481
rect 18418 14447 18452 14481
rect 18487 14447 18521 14481
rect 18556 14447 18590 14481
rect 18625 14447 18659 14481
rect 18694 14447 18728 14481
rect 18763 14447 18797 14481
rect 18832 14447 18866 14481
rect 18901 14447 18935 14481
rect 18970 14447 19004 14481
rect 19039 14447 19073 14481
rect 19108 14447 19142 14481
rect 19177 14447 19211 14481
rect 19246 14447 19280 14481
rect 19315 14447 19349 14481
rect 19384 14447 19418 14481
rect 19453 14447 19487 14481
rect 19522 14447 19556 14481
rect 19591 14447 19625 14481
rect 19660 14447 19694 14481
rect 19729 14447 19763 14481
rect 19798 14447 19832 14481
rect 19867 14447 19901 14481
rect 19936 14447 19970 14481
rect 20005 14447 20039 14481
rect 20074 14447 20108 14481
rect 20143 14447 20177 14481
rect 20212 14447 20246 14481
rect 20281 14447 20315 14481
rect 20350 14447 20384 14481
rect 20419 14447 20453 14481
rect 20488 14447 20522 14481
rect 20557 14447 20591 14481
rect 20626 14447 20660 14481
rect 20695 14447 20729 14481
rect 20764 14447 20798 14481
rect 20833 14447 20867 14481
rect 20902 14447 20936 14481
rect 20971 14447 21005 14481
rect 21040 14447 21074 14481
rect 21109 14447 21143 14481
rect 21178 14447 21212 14481
rect 21247 14447 21281 14481
rect 21315 14447 21349 14481
rect 21383 14447 21417 14481
rect 21451 14447 21485 14481
rect 21519 14447 21553 14481
rect 21587 14447 21621 14481
rect 21655 14447 21689 14481
rect 21723 14447 21757 14481
rect 21791 14447 21825 14481
rect 21859 14447 21893 14481
rect 21927 14447 21961 14481
rect 21995 14447 22029 14481
rect 22063 14447 22097 14481
rect 22131 14447 22165 14481
rect 22199 14447 22233 14481
rect 22267 14447 22301 14481
rect 22335 14447 22369 14481
rect 22403 14447 22437 14481
rect 22471 14447 22505 14481
rect 22539 14447 22573 14481
rect 22607 14447 22641 14481
rect 22675 14447 22709 14481
rect 22743 14447 22777 14481
rect 22811 14447 22845 14481
rect 22879 14447 22913 14481
rect 22947 14447 22981 14481
rect 23015 14447 23049 14481
rect 23083 14447 23117 14481
rect 23151 14447 23185 14481
rect 23219 14447 23253 14481
rect 23287 14447 23321 14481
rect 23355 14447 23389 14481
rect 23423 14447 23457 14481
rect 23491 14447 23525 14481
rect 23559 14447 23593 14481
rect 23627 14447 23661 14481
rect 23695 14447 23729 14481
rect 23763 14447 23797 14481
rect 23831 14447 23865 14481
rect 23899 14447 23933 14481
rect 23967 14447 24001 14481
rect 24035 14447 24069 14481
rect 24103 14447 24137 14481
rect 24171 14447 24205 14481
rect 24239 14447 24273 14481
rect 24307 14447 24341 14481
rect 24375 14447 24409 14481
rect 24443 14447 24477 14481
rect 24511 14447 24545 14481
rect 24579 14447 24613 14481
rect 24647 14447 24681 14481
rect 24715 14447 24749 14481
rect 24783 14447 24817 14481
rect 24851 14447 24885 14481
rect 24919 14447 24953 14481
rect 24987 14447 25021 14481
rect 25055 14447 25089 14481
rect 25123 14447 25157 14481
rect 25191 14447 25225 14481
rect 25259 14447 25293 14481
rect 25327 14447 25361 14481
rect 25395 14447 25429 14481
rect 25463 14447 25497 14481
rect 25531 14447 25565 14481
rect 25599 14447 25633 14481
rect 25667 14447 25701 14481
rect 25735 14447 25769 14481
rect 25803 14447 25837 14481
rect 25871 14447 25905 14481
rect 25939 14447 25973 14481
rect 26007 14447 26041 14481
rect 26075 14447 26109 14481
rect 26143 14447 26177 14481
rect 26211 14447 26245 14481
rect 26279 14447 26313 14481
rect 26347 14447 26381 14481
rect 26415 14447 26449 14481
rect 26483 14447 26517 14481
rect 26551 14447 26585 14481
rect 26619 14447 26653 14481
rect 26687 14447 26721 14481
rect 26755 14447 26789 14481
rect 26823 14447 26857 14481
rect 26891 14447 26925 14481
rect 26959 14447 26993 14481
rect 27027 14447 27061 14481
rect 27095 14447 27129 14481
rect 27163 14447 27197 14481
rect 27231 14447 27265 14481
rect 27299 14447 27333 14481
rect 27367 14447 27401 14481
rect 27435 14447 27469 14481
rect 27503 14447 27537 14481
rect 27571 14447 27605 14481
rect 27639 14447 27673 14481
rect 27707 14447 27741 14481
rect 27775 14447 27809 14481
rect 27843 14447 27877 14481
rect 27911 14447 27945 14481
rect 27979 14447 28013 14481
rect 28047 14447 28081 14481
rect 28115 14447 28149 14481
rect 28183 14447 28217 14481
rect 28251 14447 28285 14481
rect 28319 14447 28353 14481
rect 28387 14447 28421 14481
rect 28455 14447 28489 14481
rect 28523 14447 28557 14481
rect 28591 14447 28625 14481
rect 28659 14447 28693 14481
rect 28727 14447 28761 14481
rect 28795 14447 28829 14481
rect 28863 14447 28897 14481
rect 28931 14447 28965 14481
rect 28999 14447 29033 14481
rect 29067 14447 29101 14481
rect 29135 14447 29169 14481
rect 29203 14447 29237 14481
rect 29271 14447 29305 14481
rect 29339 14447 29373 14481
rect 29407 14447 29441 14481
rect 29475 14447 29509 14481
rect 29543 14447 29577 14481
rect 29611 14447 29645 14481
rect 18284 14381 18318 14415
rect 18356 14375 18390 14409
rect 18425 14375 18459 14409
rect 18494 14375 18528 14409
rect 18563 14375 18597 14409
rect 18632 14375 18666 14409
rect 18701 14375 18735 14409
rect 18770 14375 18804 14409
rect 18839 14375 18873 14409
rect 18908 14375 18942 14409
rect 18977 14375 19011 14409
rect 19046 14375 19080 14409
rect 19115 14375 19149 14409
rect 19184 14375 19218 14409
rect 19253 14375 19287 14409
rect 19322 14375 19356 14409
rect 19391 14375 19425 14409
rect 19460 14375 19494 14409
rect 19529 14375 19563 14409
rect 19598 14375 19632 14409
rect 19667 14375 19701 14409
rect 19736 14375 19770 14409
rect 19805 14375 19839 14409
rect 19874 14375 19908 14409
rect 19943 14375 19977 14409
rect 20012 14375 20046 14409
rect 20081 14375 20115 14409
rect 20150 14375 20184 14409
rect 20219 14375 20253 14409
rect 20288 14375 20322 14409
rect 20357 14375 20391 14409
rect 20426 14375 20460 14409
rect 20495 14375 20529 14409
rect 20564 14375 20598 14409
rect 20633 14375 20667 14409
rect 20702 14375 20736 14409
rect 20771 14375 20805 14409
rect 20839 14375 20873 14409
rect 20907 14375 20941 14409
rect 20975 14375 21009 14409
rect 21043 14375 21077 14409
rect 21111 14375 21145 14409
rect 21179 14375 21213 14409
rect 21247 14375 21281 14409
rect 21315 14375 21349 14409
rect 21383 14375 21417 14409
rect 21451 14375 21485 14409
rect 21519 14375 21553 14409
rect 21587 14375 21621 14409
rect 21655 14375 21689 14409
rect 21723 14375 21757 14409
rect 21791 14375 21825 14409
rect 21859 14375 21893 14409
rect 21927 14375 21961 14409
rect 21995 14375 22029 14409
rect 22063 14375 22097 14409
rect 22131 14375 22165 14409
rect 22199 14375 22233 14409
rect 22267 14375 22301 14409
rect 22335 14375 22369 14409
rect 22403 14375 22437 14409
rect 22471 14375 22505 14409
rect 22539 14375 22573 14409
rect 22607 14375 22641 14409
rect 22675 14375 22709 14409
rect 22743 14375 22777 14409
rect 22811 14375 22845 14409
rect 22879 14375 22913 14409
rect 22947 14375 22981 14409
rect 23015 14375 23049 14409
rect 23083 14375 23117 14409
rect 23151 14375 23185 14409
rect 23219 14375 23253 14409
rect 23287 14375 23321 14409
rect 23355 14375 23389 14409
rect 23423 14375 23457 14409
rect 23491 14375 23525 14409
rect 23559 14375 23593 14409
rect 23627 14375 23661 14409
rect 23695 14375 23729 14409
rect 23763 14375 23797 14409
rect 23831 14375 23865 14409
rect 23899 14375 23933 14409
rect 23967 14375 24001 14409
rect 24035 14375 24069 14409
rect 24103 14375 24137 14409
rect 24171 14375 24205 14409
rect 24239 14375 24273 14409
rect 24307 14375 24341 14409
rect 24375 14375 24409 14409
rect 24443 14375 24477 14409
rect 24511 14375 24545 14409
rect 24579 14375 24613 14409
rect 24647 14375 24681 14409
rect 24715 14375 24749 14409
rect 24783 14375 24817 14409
rect 24851 14375 24885 14409
rect 24919 14375 24953 14409
rect 24987 14375 25021 14409
rect 25055 14375 25089 14409
rect 25123 14375 25157 14409
rect 25191 14375 25225 14409
rect 25259 14375 25293 14409
rect 25327 14375 25361 14409
rect 25395 14375 25429 14409
rect 25463 14375 25497 14409
rect 25531 14375 25565 14409
rect 25599 14375 25633 14409
rect 25667 14375 25701 14409
rect 25735 14375 25769 14409
rect 25803 14375 25837 14409
rect 25871 14375 25905 14409
rect 25939 14375 25973 14409
rect 26007 14375 26041 14409
rect 26075 14375 26109 14409
rect 26143 14375 26177 14409
rect 26211 14375 26245 14409
rect 26279 14375 26313 14409
rect 26347 14375 26381 14409
rect 26415 14375 26449 14409
rect 26483 14375 26517 14409
rect 26551 14375 26585 14409
rect 26619 14375 26653 14409
rect 26687 14375 26721 14409
rect 26755 14375 26789 14409
rect 26823 14375 26857 14409
rect 26891 14375 26925 14409
rect 26959 14375 26993 14409
rect 27027 14375 27061 14409
rect 27095 14375 27129 14409
rect 27163 14375 27197 14409
rect 27231 14375 27265 14409
rect 27299 14375 27333 14409
rect 27367 14375 27401 14409
rect 27435 14375 27469 14409
rect 27503 14375 27537 14409
rect 27571 14375 27605 14409
rect 27639 14375 27673 14409
rect 27707 14375 27741 14409
rect 27775 14375 27809 14409
rect 27843 14375 27877 14409
rect 27911 14375 27945 14409
rect 27979 14375 28013 14409
rect 28047 14375 28081 14409
rect 28115 14375 28149 14409
rect 28183 14375 28217 14409
rect 28251 14375 28285 14409
rect 28319 14375 28353 14409
rect 28387 14375 28421 14409
rect 28455 14375 28489 14409
rect 28523 14375 28557 14409
rect 28591 14375 28625 14409
rect 28659 14375 28693 14409
rect 28727 14375 28761 14409
rect 28795 14375 28829 14409
rect 28863 14375 28897 14409
rect 28931 14375 28965 14409
rect 28999 14375 29033 14409
rect 29067 14375 29101 14409
rect 29135 14375 29169 14409
rect 29203 14375 29237 14409
rect 29271 14375 29305 14409
rect 29339 14375 29373 14409
rect 29407 14375 29441 14409
rect 29475 14375 29509 14409
rect 29543 14375 29577 14409
rect 29611 14375 29645 14409
rect 18284 14311 18318 14345
rect 18356 14306 18390 14340
rect 18428 14303 18462 14337
rect 18497 14303 18531 14337
rect 18566 14303 18600 14337
rect 18635 14303 18669 14337
rect 18704 14303 18738 14337
rect 18773 14303 18807 14337
rect 18842 14303 18876 14337
rect 18911 14303 18945 14337
rect 18980 14303 19014 14337
rect 19049 14303 19083 14337
rect 19118 14303 19152 14337
rect 19187 14303 19221 14337
rect 19256 14303 19290 14337
rect 19325 14303 19359 14337
rect 19394 14303 19428 14337
rect 19463 14303 19497 14337
rect 19532 14303 19566 14337
rect 19601 14303 19635 14337
rect 19670 14303 19704 14337
rect 19739 14303 19773 14337
rect 19808 14303 19842 14337
rect 19877 14303 19911 14337
rect 19946 14303 19980 14337
rect 20015 14303 20049 14337
rect 20084 14303 20118 14337
rect 20153 14303 20187 14337
rect 20222 14303 20256 14337
rect 20291 14303 20325 14337
rect 20360 14303 20394 14337
rect 20429 14303 20463 14337
rect 20498 14303 20532 14337
rect 20567 14303 20601 14337
rect 20635 14303 20669 14337
rect 20703 14303 20737 14337
rect 20771 14303 20805 14337
rect 20839 14303 20873 14337
rect 20907 14303 20941 14337
rect 20975 14303 21009 14337
rect 21043 14303 21077 14337
rect 21111 14303 21145 14337
rect 21179 14303 21213 14337
rect 21247 14303 21281 14337
rect 21315 14303 21349 14337
rect 21383 14303 21417 14337
rect 21451 14303 21485 14337
rect 21519 14303 21553 14337
rect 21587 14303 21621 14337
rect 21655 14303 21689 14337
rect 21723 14303 21757 14337
rect 21791 14303 21825 14337
rect 21859 14303 21893 14337
rect 21927 14303 21961 14337
rect 21995 14303 22029 14337
rect 22063 14303 22097 14337
rect 22131 14303 22165 14337
rect 22199 14303 22233 14337
rect 22267 14303 22301 14337
rect 22335 14303 22369 14337
rect 22403 14303 22437 14337
rect 22471 14303 22505 14337
rect 22539 14303 22573 14337
rect 22607 14303 22641 14337
rect 22675 14303 22709 14337
rect 22743 14303 22777 14337
rect 22811 14303 22845 14337
rect 22879 14303 22913 14337
rect 22947 14303 22981 14337
rect 23015 14303 23049 14337
rect 23083 14303 23117 14337
rect 23151 14303 23185 14337
rect 23219 14303 23253 14337
rect 23287 14303 23321 14337
rect 23355 14303 23389 14337
rect 23423 14303 23457 14337
rect 23491 14303 23525 14337
rect 23559 14303 23593 14337
rect 23627 14303 23661 14337
rect 23695 14303 23729 14337
rect 23763 14303 23797 14337
rect 23831 14303 23865 14337
rect 23899 14303 23933 14337
rect 23967 14303 24001 14337
rect 24035 14303 24069 14337
rect 24103 14303 24137 14337
rect 24171 14303 24205 14337
rect 24239 14303 24273 14337
rect 24307 14303 24341 14337
rect 24375 14303 24409 14337
rect 24443 14303 24477 14337
rect 24511 14303 24545 14337
rect 24579 14303 24613 14337
rect 24647 14303 24681 14337
rect 24715 14303 24749 14337
rect 24783 14303 24817 14337
rect 24851 14303 24885 14337
rect 24919 14303 24953 14337
rect 24987 14303 25021 14337
rect 25055 14303 25089 14337
rect 25123 14303 25157 14337
rect 25191 14303 25225 14337
rect 25259 14303 25293 14337
rect 25327 14303 25361 14337
rect 25395 14303 25429 14337
rect 25463 14303 25497 14337
rect 25531 14303 25565 14337
rect 25599 14303 25633 14337
rect 25667 14303 25701 14337
rect 25735 14303 25769 14337
rect 25803 14303 25837 14337
rect 25871 14303 25905 14337
rect 25939 14303 25973 14337
rect 26007 14303 26041 14337
rect 26075 14303 26109 14337
rect 26143 14303 26177 14337
rect 26211 14303 26245 14337
rect 26279 14303 26313 14337
rect 26347 14303 26381 14337
rect 26415 14303 26449 14337
rect 26483 14303 26517 14337
rect 26551 14303 26585 14337
rect 26619 14303 26653 14337
rect 26687 14303 26721 14337
rect 26755 14303 26789 14337
rect 26823 14303 26857 14337
rect 26891 14303 26925 14337
rect 26959 14303 26993 14337
rect 27027 14303 27061 14337
rect 27095 14303 27129 14337
rect 27163 14303 27197 14337
rect 27231 14303 27265 14337
rect 27299 14303 27333 14337
rect 27367 14303 27401 14337
rect 27435 14303 27469 14337
rect 27503 14303 27537 14337
rect 27571 14303 27605 14337
rect 27639 14303 27673 14337
rect 27707 14303 27741 14337
rect 27775 14303 27809 14337
rect 27843 14303 27877 14337
rect 27911 14303 27945 14337
rect 27979 14303 28013 14337
rect 28047 14303 28081 14337
rect 28115 14303 28149 14337
rect 28183 14303 28217 14337
rect 28251 14303 28285 14337
rect 28319 14303 28353 14337
rect 28387 14303 28421 14337
rect 28455 14303 28489 14337
rect 28523 14303 28557 14337
rect 28591 14303 28625 14337
rect 28659 14303 28693 14337
rect 28727 14303 28761 14337
rect 28795 14303 28829 14337
rect 28863 14303 28897 14337
rect 28931 14303 28965 14337
rect 28999 14303 29033 14337
rect 29067 14303 29101 14337
rect 29135 14303 29169 14337
rect 29203 14303 29237 14337
rect 29271 14303 29305 14337
rect 29339 14303 29373 14337
rect 29407 14303 29441 14337
rect 29475 14303 29509 14337
rect 29543 14303 29577 14337
rect 29611 14303 29645 14337
rect 18284 14241 18318 14275
rect 18356 14237 18390 14271
rect 18428 14234 18462 14268
rect 18500 14231 18534 14265
rect 18569 14231 18603 14265
rect 18638 14231 18672 14265
rect 18707 14231 18741 14265
rect 18776 14231 18810 14265
rect 18845 14231 18879 14265
rect 18914 14231 18948 14265
rect 18983 14231 19017 14265
rect 19052 14231 19086 14265
rect 19121 14231 19155 14265
rect 19190 14231 19224 14265
rect 19259 14231 19293 14265
rect 19328 14231 19362 14265
rect 19397 14231 19431 14265
rect 19466 14231 19500 14265
rect 19535 14231 19569 14265
rect 19604 14231 19638 14265
rect 19673 14231 19707 14265
rect 19742 14231 19776 14265
rect 19811 14231 19845 14265
rect 19880 14231 19914 14265
rect 19949 14231 19983 14265
rect 20018 14231 20052 14265
rect 20087 14231 20121 14265
rect 20156 14231 20190 14265
rect 20225 14231 20259 14265
rect 20294 14231 20328 14265
rect 20363 14231 20397 14265
rect 20431 14231 20465 14265
rect 20499 14231 20533 14265
rect 20567 14231 20601 14265
rect 20635 14231 20669 14265
rect 20703 14231 20737 14265
rect 20771 14231 20805 14265
rect 20839 14231 20873 14265
rect 20907 14231 20941 14265
rect 20975 14231 21009 14265
rect 21043 14231 21077 14265
rect 21111 14231 21145 14265
rect 21179 14231 21213 14265
rect 21247 14231 21281 14265
rect 21315 14231 21349 14265
rect 21383 14231 21417 14265
rect 21451 14231 21485 14265
rect 21519 14231 21553 14265
rect 21587 14231 21621 14265
rect 21655 14231 21689 14265
rect 21723 14231 21757 14265
rect 21791 14231 21825 14265
rect 21859 14231 21893 14265
rect 21927 14231 21961 14265
rect 21995 14231 22029 14265
rect 22063 14231 22097 14265
rect 22131 14231 22165 14265
rect 22199 14231 22233 14265
rect 22267 14231 22301 14265
rect 22335 14231 22369 14265
rect 22403 14231 22437 14265
rect 22471 14231 22505 14265
rect 22539 14231 22573 14265
rect 22607 14231 22641 14265
rect 22675 14231 22709 14265
rect 22743 14231 22777 14265
rect 22811 14231 22845 14265
rect 22879 14231 22913 14265
rect 22947 14231 22981 14265
rect 23015 14231 23049 14265
rect 23083 14231 23117 14265
rect 23151 14231 23185 14265
rect 23219 14231 23253 14265
rect 23287 14231 23321 14265
rect 23355 14231 23389 14265
rect 23423 14231 23457 14265
rect 23491 14231 23525 14265
rect 23559 14231 23593 14265
rect 23627 14231 23661 14265
rect 23695 14231 23729 14265
rect 23763 14231 23797 14265
rect 23831 14231 23865 14265
rect 23899 14231 23933 14265
rect 23967 14231 24001 14265
rect 24035 14231 24069 14265
rect 24103 14231 24137 14265
rect 24171 14231 24205 14265
rect 24239 14231 24273 14265
rect 24307 14231 24341 14265
rect 24375 14231 24409 14265
rect 24443 14231 24477 14265
rect 24511 14231 24545 14265
rect 24579 14231 24613 14265
rect 24647 14231 24681 14265
rect 24715 14231 24749 14265
rect 24783 14231 24817 14265
rect 24851 14231 24885 14265
rect 24919 14231 24953 14265
rect 24987 14231 25021 14265
rect 25055 14231 25089 14265
rect 25123 14231 25157 14265
rect 25191 14231 25225 14265
rect 25259 14231 25293 14265
rect 25327 14231 25361 14265
rect 25395 14231 25429 14265
rect 25463 14231 25497 14265
rect 25531 14231 25565 14265
rect 25599 14231 25633 14265
rect 25667 14231 25701 14265
rect 25735 14231 25769 14265
rect 25803 14231 25837 14265
rect 25871 14231 25905 14265
rect 25939 14231 25973 14265
rect 26007 14231 26041 14265
rect 26075 14231 26109 14265
rect 26143 14231 26177 14265
rect 26211 14231 26245 14265
rect 26279 14231 26313 14265
rect 26347 14231 26381 14265
rect 26415 14231 26449 14265
rect 26483 14231 26517 14265
rect 26551 14231 26585 14265
rect 26619 14231 26653 14265
rect 26687 14231 26721 14265
rect 26755 14231 26789 14265
rect 26823 14231 26857 14265
rect 26891 14231 26925 14265
rect 26959 14231 26993 14265
rect 27027 14231 27061 14265
rect 27095 14231 27129 14265
rect 27163 14231 27197 14265
rect 27231 14231 27265 14265
rect 27299 14231 27333 14265
rect 27367 14231 27401 14265
rect 27435 14231 27469 14265
rect 27503 14231 27537 14265
rect 27571 14231 27605 14265
rect 27639 14231 27673 14265
rect 27707 14231 27741 14265
rect 27775 14231 27809 14265
rect 27843 14231 27877 14265
rect 27911 14231 27945 14265
rect 27979 14231 28013 14265
rect 28047 14231 28081 14265
rect 28115 14231 28149 14265
rect 28183 14231 28217 14265
rect 28251 14231 28285 14265
rect 28319 14231 28353 14265
rect 28387 14231 28421 14265
rect 28455 14231 28489 14265
rect 28523 14231 28557 14265
rect 28591 14231 28625 14265
rect 28659 14231 28693 14265
rect 28727 14231 28761 14265
rect 28795 14231 28829 14265
rect 28863 14231 28897 14265
rect 28931 14231 28965 14265
rect 28999 14231 29033 14265
rect 29067 14231 29101 14265
rect 29135 14231 29169 14265
rect 29203 14231 29237 14265
rect 29271 14231 29305 14265
rect 29339 14231 29373 14265
rect 29407 14231 29441 14265
rect 29475 14231 29509 14265
rect 29543 14231 29577 14265
rect 29611 14231 29645 14265
rect 15855 14171 15889 14205
rect 15925 14171 15959 14205
rect 15995 14171 16029 14205
rect 16065 14171 16099 14205
rect 16135 14171 16169 14205
rect 16205 14171 16239 14205
rect 16275 14171 16309 14205
rect 16345 14171 16379 14205
rect 16415 14171 16449 14205
rect 16485 14171 16519 14205
rect 16555 14171 16589 14205
rect 16625 14171 16659 14205
rect 16695 14171 16729 14205
rect 16765 14171 16799 14205
rect 16835 14171 16869 14205
rect 16904 14171 16938 14205
rect 16973 14171 17007 14205
rect 17042 14171 17076 14205
rect 17111 14171 17145 14205
rect 17180 14171 17214 14205
rect 17249 14171 17283 14205
rect 17318 14171 17352 14205
rect 17387 14171 17421 14205
rect 17456 14171 17490 14205
rect 17525 14171 17559 14205
rect 17594 14171 17628 14205
rect 17663 14171 17697 14205
rect 17732 14171 17766 14205
rect 17801 14171 17835 14205
rect 17870 14171 17904 14205
rect 17939 14171 17973 14205
rect 18008 14171 18042 14205
rect 18077 14171 18111 14205
rect 18146 14171 18180 14205
rect 18215 14171 18249 14205
rect 18284 14171 18318 14205
rect 18356 14168 18390 14202
rect 18428 14165 18462 14199
rect 18500 14162 18534 14196
rect 18572 14159 18606 14193
rect 18641 14159 18675 14193
rect 18710 14159 18744 14193
rect 18779 14159 18813 14193
rect 18848 14159 18882 14193
rect 18917 14159 18951 14193
rect 18986 14159 19020 14193
rect 19055 14159 19089 14193
rect 19124 14159 19158 14193
rect 19193 14159 19227 14193
rect 19262 14159 19296 14193
rect 19331 14159 19365 14193
rect 19400 14159 19434 14193
rect 19469 14159 19503 14193
rect 19538 14159 19572 14193
rect 19607 14159 19641 14193
rect 19676 14159 19710 14193
rect 19745 14159 19779 14193
rect 19814 14159 19848 14193
rect 19883 14159 19917 14193
rect 19952 14159 19986 14193
rect 20021 14159 20055 14193
rect 20090 14159 20124 14193
rect 20159 14159 20193 14193
rect 20227 14159 20261 14193
rect 20295 14159 20329 14193
rect 20363 14159 20397 14193
rect 20431 14159 20465 14193
rect 20499 14159 20533 14193
rect 20567 14159 20601 14193
rect 20635 14159 20669 14193
rect 20703 14159 20737 14193
rect 20771 14159 20805 14193
rect 20839 14159 20873 14193
rect 20907 14159 20941 14193
rect 20975 14159 21009 14193
rect 21043 14159 21077 14193
rect 21111 14159 21145 14193
rect 21179 14159 21213 14193
rect 21247 14159 21281 14193
rect 21315 14159 21349 14193
rect 21383 14159 21417 14193
rect 21451 14159 21485 14193
rect 21519 14159 21553 14193
rect 21587 14159 21621 14193
rect 21655 14159 21689 14193
rect 21723 14159 21757 14193
rect 21791 14159 21825 14193
rect 21859 14159 21893 14193
rect 21927 14159 21961 14193
rect 21995 14159 22029 14193
rect 22063 14159 22097 14193
rect 22131 14159 22165 14193
rect 22199 14159 22233 14193
rect 22267 14159 22301 14193
rect 22335 14159 22369 14193
rect 22403 14159 22437 14193
rect 22471 14159 22505 14193
rect 22539 14159 22573 14193
rect 22607 14159 22641 14193
rect 22675 14159 22709 14193
rect 22743 14159 22777 14193
rect 22811 14159 22845 14193
rect 22879 14159 22913 14193
rect 22947 14159 22981 14193
rect 23015 14159 23049 14193
rect 23083 14159 23117 14193
rect 23151 14159 23185 14193
rect 23219 14159 23253 14193
rect 23287 14159 23321 14193
rect 23355 14159 23389 14193
rect 23423 14159 23457 14193
rect 23491 14159 23525 14193
rect 23559 14159 23593 14193
rect 23627 14159 23661 14193
rect 23695 14159 23729 14193
rect 23763 14159 23797 14193
rect 23831 14159 23865 14193
rect 23899 14159 23933 14193
rect 23967 14159 24001 14193
rect 24035 14159 24069 14193
rect 24103 14159 24137 14193
rect 24171 14159 24205 14193
rect 24239 14159 24273 14193
rect 24307 14159 24341 14193
rect 24375 14159 24409 14193
rect 24443 14159 24477 14193
rect 24511 14159 24545 14193
rect 24579 14159 24613 14193
rect 24647 14159 24681 14193
rect 24715 14159 24749 14193
rect 24783 14159 24817 14193
rect 24851 14159 24885 14193
rect 24919 14159 24953 14193
rect 24987 14159 25021 14193
rect 25055 14159 25089 14193
rect 25123 14159 25157 14193
rect 25191 14159 25225 14193
rect 25259 14159 25293 14193
rect 25327 14159 25361 14193
rect 25395 14159 25429 14193
rect 25463 14159 25497 14193
rect 25531 14159 25565 14193
rect 25599 14159 25633 14193
rect 25667 14159 25701 14193
rect 25735 14159 25769 14193
rect 25803 14159 25837 14193
rect 25871 14159 25905 14193
rect 25939 14159 25973 14193
rect 26007 14159 26041 14193
rect 26075 14159 26109 14193
rect 26143 14159 26177 14193
rect 26211 14159 26245 14193
rect 26279 14159 26313 14193
rect 26347 14159 26381 14193
rect 26415 14159 26449 14193
rect 26483 14159 26517 14193
rect 26551 14159 26585 14193
rect 26619 14159 26653 14193
rect 26687 14159 26721 14193
rect 26755 14159 26789 14193
rect 26823 14159 26857 14193
rect 26891 14159 26925 14193
rect 26959 14159 26993 14193
rect 27027 14159 27061 14193
rect 27095 14159 27129 14193
rect 27163 14159 27197 14193
rect 27231 14159 27265 14193
rect 27299 14159 27333 14193
rect 27367 14159 27401 14193
rect 27435 14159 27469 14193
rect 27503 14159 27537 14193
rect 27571 14159 27605 14193
rect 27639 14159 27673 14193
rect 27707 14159 27741 14193
rect 27775 14159 27809 14193
rect 27843 14159 27877 14193
rect 27911 14159 27945 14193
rect 27979 14159 28013 14193
rect 28047 14159 28081 14193
rect 28115 14159 28149 14193
rect 28183 14159 28217 14193
rect 28251 14159 28285 14193
rect 28319 14159 28353 14193
rect 28387 14159 28421 14193
rect 28455 14159 28489 14193
rect 28523 14159 28557 14193
rect 28591 14159 28625 14193
rect 28659 14159 28693 14193
rect 28727 14159 28761 14193
rect 28795 14159 28829 14193
rect 28863 14159 28897 14193
rect 28931 14159 28965 14193
rect 28999 14159 29033 14193
rect 29067 14159 29101 14193
rect 29135 14159 29169 14193
rect 29203 14159 29237 14193
rect 29271 14159 29305 14193
rect 29339 14159 29373 14193
rect 29407 14159 29441 14193
rect 29475 14159 29509 14193
rect 29543 14159 29577 14193
rect 29611 14159 29645 14193
rect 15855 14099 15889 14133
rect 15925 14099 15959 14133
rect 15995 14099 16029 14133
rect 16065 14099 16099 14133
rect 16135 14099 16169 14133
rect 16205 14099 16239 14133
rect 16275 14099 16309 14133
rect 16345 14099 16379 14133
rect 16415 14099 16449 14133
rect 16485 14099 16519 14133
rect 16555 14099 16589 14133
rect 16625 14099 16659 14133
rect 16695 14099 16729 14133
rect 16765 14099 16799 14133
rect 16835 14099 16869 14133
rect 16905 14099 16939 14133
rect 16975 14099 17009 14133
rect 17045 14099 17079 14133
rect 17114 14099 17148 14133
rect 17183 14099 17217 14133
rect 17252 14099 17286 14133
rect 17321 14099 17355 14133
rect 17390 14099 17424 14133
rect 17459 14099 17493 14133
rect 17528 14099 17562 14133
rect 17597 14099 17631 14133
rect 17666 14099 17700 14133
rect 17735 14099 17769 14133
rect 17804 14099 17838 14133
rect 17873 14099 17907 14133
rect 17942 14099 17976 14133
rect 18011 14099 18045 14133
rect 18080 14099 18114 14133
rect 18149 14099 18183 14133
rect 18218 14099 18252 14133
rect 18287 14099 18321 14133
rect 18356 14099 18390 14133
rect 18428 14096 18462 14130
rect 18500 14093 18534 14127
rect 18572 14090 18606 14124
rect 18644 14087 18678 14121
rect 18713 14087 18747 14121
rect 18782 14087 18816 14121
rect 18851 14087 18885 14121
rect 18920 14087 18954 14121
rect 18989 14087 19023 14121
rect 19058 14087 19092 14121
rect 19127 14087 19161 14121
rect 19196 14087 19230 14121
rect 19265 14087 19299 14121
rect 19334 14087 19368 14121
rect 19403 14087 19437 14121
rect 19472 14087 19506 14121
rect 19541 14087 19575 14121
rect 19610 14087 19644 14121
rect 19679 14087 19713 14121
rect 19748 14087 19782 14121
rect 19817 14087 19851 14121
rect 19886 14087 19920 14121
rect 19955 14087 19989 14121
rect 20023 14087 20057 14121
rect 20091 14087 20125 14121
rect 20159 14087 20193 14121
rect 20227 14087 20261 14121
rect 20295 14087 20329 14121
rect 20363 14087 20397 14121
rect 20431 14087 20465 14121
rect 20499 14087 20533 14121
rect 20567 14087 20601 14121
rect 20635 14087 20669 14121
rect 20703 14087 20737 14121
rect 20771 14087 20805 14121
rect 20839 14087 20873 14121
rect 20907 14087 20941 14121
rect 20975 14087 21009 14121
rect 21043 14087 21077 14121
rect 21111 14087 21145 14121
rect 21179 14087 21213 14121
rect 21247 14087 21281 14121
rect 21315 14087 21349 14121
rect 21383 14087 21417 14121
rect 21451 14087 21485 14121
rect 21519 14087 21553 14121
rect 21587 14087 21621 14121
rect 21655 14087 21689 14121
rect 21723 14087 21757 14121
rect 21791 14087 21825 14121
rect 21859 14087 21893 14121
rect 21927 14087 21961 14121
rect 21995 14087 22029 14121
rect 22063 14087 22097 14121
rect 22131 14087 22165 14121
rect 22199 14087 22233 14121
rect 22267 14087 22301 14121
rect 22335 14087 22369 14121
rect 22403 14087 22437 14121
rect 22471 14087 22505 14121
rect 22539 14087 22573 14121
rect 22607 14087 22641 14121
rect 22675 14087 22709 14121
rect 22743 14087 22777 14121
rect 22811 14087 22845 14121
rect 22879 14087 22913 14121
rect 22947 14087 22981 14121
rect 23015 14087 23049 14121
rect 23083 14087 23117 14121
rect 23151 14087 23185 14121
rect 23219 14087 23253 14121
rect 23287 14087 23321 14121
rect 23355 14087 23389 14121
rect 23423 14087 23457 14121
rect 23491 14087 23525 14121
rect 23559 14087 23593 14121
rect 23627 14087 23661 14121
rect 23695 14087 23729 14121
rect 23763 14087 23797 14121
rect 23831 14087 23865 14121
rect 23899 14087 23933 14121
rect 23967 14087 24001 14121
rect 24035 14087 24069 14121
rect 24103 14087 24137 14121
rect 24171 14087 24205 14121
rect 24239 14087 24273 14121
rect 24307 14087 24341 14121
rect 24375 14087 24409 14121
rect 24443 14087 24477 14121
rect 24511 14087 24545 14121
rect 24579 14087 24613 14121
rect 24647 14087 24681 14121
rect 24715 14087 24749 14121
rect 24783 14087 24817 14121
rect 24851 14087 24885 14121
rect 24919 14087 24953 14121
rect 24987 14087 25021 14121
rect 25055 14087 25089 14121
rect 25123 14087 25157 14121
rect 25191 14087 25225 14121
rect 25259 14087 25293 14121
rect 25327 14087 25361 14121
rect 25395 14087 25429 14121
rect 25463 14087 25497 14121
rect 25531 14087 25565 14121
rect 25599 14087 25633 14121
rect 25667 14087 25701 14121
rect 25735 14087 25769 14121
rect 25803 14087 25837 14121
rect 25871 14087 25905 14121
rect 25939 14087 25973 14121
rect 26007 14087 26041 14121
rect 26075 14087 26109 14121
rect 26143 14087 26177 14121
rect 26211 14087 26245 14121
rect 26279 14087 26313 14121
rect 26347 14087 26381 14121
rect 26415 14087 26449 14121
rect 26483 14087 26517 14121
rect 26551 14087 26585 14121
rect 26619 14087 26653 14121
rect 26687 14087 26721 14121
rect 26755 14087 26789 14121
rect 26823 14087 26857 14121
rect 26891 14087 26925 14121
rect 26959 14087 26993 14121
rect 27027 14087 27061 14121
rect 27095 14087 27129 14121
rect 27163 14087 27197 14121
rect 27231 14087 27265 14121
rect 27299 14087 27333 14121
rect 27367 14087 27401 14121
rect 27435 14087 27469 14121
rect 27503 14087 27537 14121
rect 27571 14087 27605 14121
rect 27639 14087 27673 14121
rect 27707 14087 27741 14121
rect 27775 14087 27809 14121
rect 27843 14087 27877 14121
rect 27911 14087 27945 14121
rect 27979 14087 28013 14121
rect 28047 14087 28081 14121
rect 28115 14087 28149 14121
rect 28183 14087 28217 14121
rect 28251 14087 28285 14121
rect 28319 14087 28353 14121
rect 28387 14087 28421 14121
rect 28455 14087 28489 14121
rect 28523 14087 28557 14121
rect 28591 14087 28625 14121
rect 28659 14087 28693 14121
rect 28727 14087 28761 14121
rect 28795 14087 28829 14121
rect 28863 14087 28897 14121
rect 28931 14087 28965 14121
rect 28999 14087 29033 14121
rect 29067 14087 29101 14121
rect 29135 14087 29169 14121
rect 29203 14087 29237 14121
rect 29271 14087 29305 14121
rect 29339 14087 29373 14121
rect 29407 14087 29441 14121
rect 29475 14087 29509 14121
rect 29543 14087 29577 14121
rect 29611 14087 29645 14121
rect 15855 14027 15889 14061
rect 15925 14027 15959 14061
rect 15995 14027 16029 14061
rect 16065 14027 16099 14061
rect 16135 14027 16169 14061
rect 16205 14027 16239 14061
rect 16275 14027 16309 14061
rect 16345 14027 16379 14061
rect 16415 14027 16449 14061
rect 16485 14027 16519 14061
rect 16555 14027 16589 14061
rect 16625 14027 16659 14061
rect 16695 14027 16729 14061
rect 16765 14027 16799 14061
rect 16835 14027 16869 14061
rect 16905 14027 16939 14061
rect 16975 14027 17009 14061
rect 17045 14027 17079 14061
rect 17115 14027 17149 14061
rect 17185 14027 17219 14061
rect 17255 14027 17289 14061
rect 17324 14027 17358 14061
rect 17393 14027 17427 14061
rect 17462 14027 17496 14061
rect 17531 14027 17565 14061
rect 17600 14027 17634 14061
rect 17669 14027 17703 14061
rect 17738 14027 17772 14061
rect 17807 14027 17841 14061
rect 17876 14027 17910 14061
rect 17945 14027 17979 14061
rect 18014 14027 18048 14061
rect 18083 14027 18117 14061
rect 18152 14027 18186 14061
rect 18221 14027 18255 14061
rect 18290 14027 18324 14061
rect 18359 14027 18393 14061
rect 18428 14027 18462 14061
rect 18500 14024 18534 14058
rect 18572 14021 18606 14055
rect 18644 14017 18678 14051
rect 15855 13955 15889 13989
rect 15925 13955 15959 13989
rect 15995 13955 16029 13989
rect 16065 13955 16099 13989
rect 16135 13955 16169 13989
rect 16205 13955 16239 13989
rect 16275 13955 16309 13989
rect 16345 13955 16379 13989
rect 16415 13955 16449 13989
rect 16485 13955 16519 13989
rect 16555 13955 16589 13989
rect 16625 13955 16659 13989
rect 16695 13955 16729 13989
rect 16765 13955 16799 13989
rect 16835 13955 16869 13989
rect 16905 13955 16939 13989
rect 16975 13955 17009 13989
rect 17045 13955 17079 13989
rect 17115 13955 17149 13989
rect 17185 13955 17219 13989
rect 17255 13955 17289 13989
rect 17325 13955 17359 13989
rect 17395 13955 17429 13989
rect 17465 13955 17499 13989
rect 17534 13955 17568 13989
rect 17603 13955 17637 13989
rect 17672 13955 17706 13989
rect 17741 13955 17775 13989
rect 17810 13955 17844 13989
rect 17879 13955 17913 13989
rect 17948 13955 17982 13989
rect 18017 13955 18051 13989
rect 18086 13955 18120 13989
rect 18155 13955 18189 13989
rect 18224 13955 18258 13989
rect 18293 13955 18327 13989
rect 18362 13955 18396 13989
rect 18431 13955 18465 13989
rect 18500 13955 18534 13989
rect 18572 13952 18606 13986
rect 18644 13947 18678 13981
rect 15855 13883 15889 13917
rect 15925 13883 15959 13917
rect 15995 13883 16029 13917
rect 16065 13883 16099 13917
rect 16135 13883 16169 13917
rect 16205 13883 16239 13917
rect 16275 13883 16309 13917
rect 16345 13883 16379 13917
rect 16415 13883 16449 13917
rect 16485 13883 16519 13917
rect 16555 13883 16589 13917
rect 16625 13883 16659 13917
rect 16695 13883 16729 13917
rect 16765 13883 16799 13917
rect 16835 13883 16869 13917
rect 16905 13883 16939 13917
rect 16975 13883 17009 13917
rect 17045 13883 17079 13917
rect 17115 13883 17149 13917
rect 17185 13883 17219 13917
rect 17255 13883 17289 13917
rect 17325 13883 17359 13917
rect 17395 13883 17429 13917
rect 17465 13883 17499 13917
rect 17535 13883 17569 13917
rect 17605 13883 17639 13917
rect 17675 13883 17709 13917
rect 17744 13883 17778 13917
rect 17813 13883 17847 13917
rect 17882 13883 17916 13917
rect 17951 13883 17985 13917
rect 18020 13883 18054 13917
rect 18089 13883 18123 13917
rect 18158 13883 18192 13917
rect 18227 13883 18261 13917
rect 18296 13883 18330 13917
rect 18365 13883 18399 13917
rect 18434 13883 18468 13917
rect 18503 13883 18537 13917
rect 18572 13883 18606 13917
rect 18644 13876 18678 13910
rect 15855 13811 15889 13845
rect 15924 13811 15958 13845
rect 15993 13811 16027 13845
rect 16062 13811 16096 13845
rect 16131 13811 16165 13845
rect 16199 13811 16233 13845
rect 16267 13811 16301 13845
rect 16335 13811 16369 13845
rect 16403 13811 16437 13845
rect 16471 13811 16505 13845
rect 16539 13811 16573 13845
rect 16607 13811 16641 13845
rect 16675 13811 16709 13845
rect 16743 13811 16777 13845
rect 16811 13811 16845 13845
rect 16879 13811 16913 13845
rect 16947 13811 16981 13845
rect 17015 13811 17049 13845
rect 17083 13811 17117 13845
rect 17151 13811 17185 13845
rect 17219 13811 17253 13845
rect 17287 13811 17321 13845
rect 17355 13811 17389 13845
rect 17423 13811 17457 13845
rect 17491 13811 17525 13845
rect 17559 13811 17593 13845
rect 17627 13811 17661 13845
rect 17695 13811 17729 13845
rect 17763 13811 17797 13845
rect 17831 13811 17865 13845
rect 17899 13811 17933 13845
rect 17967 13811 18001 13845
rect 18035 13811 18069 13845
rect 18103 13811 18137 13845
rect 18171 13811 18205 13845
rect 18239 13811 18273 13845
rect 18307 13811 18341 13845
rect 18375 13811 18409 13845
rect 18443 13811 18477 13845
rect 18511 13811 18545 13845
rect 18579 13811 18613 13845
rect 13279 12087 13313 12121
rect 13347 12087 13381 12121
rect 13415 12087 13449 12121
rect 13483 12087 13517 12121
rect 13551 12087 13585 12121
rect 13619 12087 13653 12121
rect 13687 12087 13721 12121
rect 13755 12087 13789 12121
rect 13823 12087 13857 12121
rect 13891 12087 13925 12121
rect 13959 12087 13993 12121
rect 14027 12087 14061 12121
rect 14095 12087 14129 12121
rect 14163 12087 14197 12121
rect 14231 12087 14265 12121
rect 14299 12087 14333 12121
rect 14367 12087 14401 12121
rect 14435 12087 14469 12121
rect 14503 12087 14537 12121
rect 14571 12087 14605 12121
rect 14639 12087 14673 12121
rect 14707 12087 14741 12121
rect 14775 12087 14809 12121
rect 14843 12087 14877 12121
rect 14911 12087 14945 12121
rect 14979 12087 15013 12121
rect 15047 12087 15081 12121
rect 15115 12087 15149 12121
rect 15183 12087 15217 12121
rect 15251 12087 15285 12121
rect 15319 12087 15353 12121
rect 15387 12087 15421 12121
rect 15455 12087 15489 12121
rect 15523 12087 15557 12121
rect 15591 12087 15625 12121
rect 15659 12087 15693 12121
rect 15727 12087 15761 12121
rect 15795 12087 15829 12121
rect 13279 12018 13313 12052
rect 13347 12018 13381 12052
rect 13415 12018 13449 12052
rect 13483 12018 13517 12052
rect 13551 12018 13585 12052
rect 13619 12018 13653 12052
rect 13687 12018 13721 12052
rect 13755 12018 13789 12052
rect 13823 12018 13857 12052
rect 13891 12018 13925 12052
rect 13959 12018 13993 12052
rect 14027 12018 14061 12052
rect 14095 12018 14129 12052
rect 14163 12018 14197 12052
rect 14231 12018 14265 12052
rect 14299 12018 14333 12052
rect 14367 12018 14401 12052
rect 14435 12018 14469 12052
rect 14503 12018 14537 12052
rect 14571 12018 14605 12052
rect 14639 12018 14673 12052
rect 14707 12018 14741 12052
rect 14775 12018 14809 12052
rect 14843 12018 14877 12052
rect 14911 12018 14945 12052
rect 14979 12018 15013 12052
rect 15047 12018 15081 12052
rect 15115 12018 15149 12052
rect 15183 12018 15217 12052
rect 15251 12018 15285 12052
rect 15319 12018 15353 12052
rect 15387 12018 15421 12052
rect 15455 12018 15489 12052
rect 15523 12018 15557 12052
rect 15591 12018 15625 12052
rect 15659 12018 15693 12052
rect 15727 12018 15761 12052
rect 15795 12018 15829 12052
rect 13279 11949 13313 11983
rect 13347 11949 13381 11983
rect 13415 11949 13449 11983
rect 13483 11949 13517 11983
rect 13551 11949 13585 11983
rect 13619 11949 13653 11983
rect 13687 11949 13721 11983
rect 13755 11949 13789 11983
rect 13823 11949 13857 11983
rect 13891 11949 13925 11983
rect 13959 11949 13993 11983
rect 14027 11949 14061 11983
rect 14095 11949 14129 11983
rect 14163 11949 14197 11983
rect 14231 11949 14265 11983
rect 14299 11949 14333 11983
rect 14367 11949 14401 11983
rect 14435 11949 14469 11983
rect 14503 11949 14537 11983
rect 14571 11949 14605 11983
rect 14639 11949 14673 11983
rect 14707 11949 14741 11983
rect 14775 11949 14809 11983
rect 14843 11949 14877 11983
rect 14911 11949 14945 11983
rect 14979 11949 15013 11983
rect 15047 11949 15081 11983
rect 15115 11949 15149 11983
rect 15183 11949 15217 11983
rect 15251 11949 15285 11983
rect 15319 11949 15353 11983
rect 15387 11949 15421 11983
rect 15455 11949 15489 11983
rect 15523 11949 15557 11983
rect 15591 11949 15625 11983
rect 15659 11949 15693 11983
rect 15727 11949 15761 11983
rect 15795 11949 15829 11983
rect -2959 10344 -2925 10378
rect -2891 10344 -2857 10378
rect -2823 10344 -2789 10378
rect -2755 10344 -2721 10378
rect -2687 10344 -2653 10378
rect -2619 10344 -2585 10378
rect -2551 10344 -2517 10378
rect -2483 10344 -2449 10378
rect -2415 10344 -2381 10378
rect -2347 10344 -2313 10378
rect -2279 10344 -2245 10378
rect -2211 10344 -2177 10378
rect -2143 10344 -2109 10378
rect -2075 10344 -2041 10378
rect -2007 10344 -1973 10378
rect -1939 10344 -1905 10378
rect -1871 10344 -1837 10378
rect -1803 10344 -1769 10378
rect -1735 10344 -1701 10378
rect -1667 10344 -1633 10378
rect -1599 10344 -1565 10378
rect -1531 10344 -1497 10378
rect -1463 10344 -1429 10378
rect -1395 10344 -1361 10378
rect -1327 10344 -1293 10378
rect -1259 10344 -1225 10378
rect -1191 10344 -1157 10378
rect -1123 10344 -1089 10378
rect -1055 10344 -1021 10378
rect -987 10344 -953 10378
rect -919 10344 -885 10378
rect -851 10344 -817 10378
rect -783 10344 -749 10378
rect -715 10344 -681 10378
rect -647 10344 -613 10378
rect -579 10344 -545 10378
rect -511 10344 -477 10378
rect -443 10344 -409 10378
rect -375 10344 -341 10378
rect -307 10344 -273 10378
rect -2959 10275 -2925 10309
rect -2891 10275 -2857 10309
rect -2823 10275 -2789 10309
rect -2755 10275 -2721 10309
rect -2687 10275 -2653 10309
rect -2619 10275 -2585 10309
rect -2551 10275 -2517 10309
rect -2483 10275 -2449 10309
rect -2415 10275 -2381 10309
rect -2347 10275 -2313 10309
rect -2279 10275 -2245 10309
rect -2211 10275 -2177 10309
rect -2143 10275 -2109 10309
rect -2075 10275 -2041 10309
rect -2007 10275 -1973 10309
rect -1939 10275 -1905 10309
rect -1871 10275 -1837 10309
rect -1803 10275 -1769 10309
rect -1735 10275 -1701 10309
rect -1667 10275 -1633 10309
rect -1599 10275 -1565 10309
rect -1531 10275 -1497 10309
rect -1463 10275 -1429 10309
rect -1395 10275 -1361 10309
rect -1327 10275 -1293 10309
rect -1259 10275 -1225 10309
rect -1191 10275 -1157 10309
rect -1123 10275 -1089 10309
rect -1055 10275 -1021 10309
rect -987 10275 -953 10309
rect -919 10275 -885 10309
rect -851 10275 -817 10309
rect -783 10275 -749 10309
rect -715 10275 -681 10309
rect -647 10275 -613 10309
rect -579 10275 -545 10309
rect -511 10275 -477 10309
rect -443 10275 -409 10309
rect -375 10275 -341 10309
rect -307 10275 -273 10309
rect -2959 10206 -2925 10240
rect -2891 10206 -2857 10240
rect -2823 10206 -2789 10240
rect -2755 10206 -2721 10240
rect -2687 10206 -2653 10240
rect -2619 10206 -2585 10240
rect -2551 10206 -2517 10240
rect -2483 10206 -2449 10240
rect -2415 10206 -2381 10240
rect -2347 10206 -2313 10240
rect -2279 10206 -2245 10240
rect -2211 10206 -2177 10240
rect -2143 10206 -2109 10240
rect -2075 10206 -2041 10240
rect -2007 10206 -1973 10240
rect -1939 10206 -1905 10240
rect -1871 10206 -1837 10240
rect -1803 10206 -1769 10240
rect -1735 10206 -1701 10240
rect -1667 10206 -1633 10240
rect -1599 10206 -1565 10240
rect -1531 10206 -1497 10240
rect -1463 10206 -1429 10240
rect -1395 10206 -1361 10240
rect -1327 10206 -1293 10240
rect -1259 10206 -1225 10240
rect -1191 10206 -1157 10240
rect -1123 10206 -1089 10240
rect -1055 10206 -1021 10240
rect -987 10206 -953 10240
rect -919 10206 -885 10240
rect -851 10206 -817 10240
rect -783 10206 -749 10240
rect -715 10206 -681 10240
rect -647 10206 -613 10240
rect -579 10206 -545 10240
rect -511 10206 -477 10240
rect -443 10206 -409 10240
rect -375 10206 -341 10240
rect -307 10206 -273 10240
rect -2959 10137 -2925 10171
rect -2891 10137 -2857 10171
rect -2823 10137 -2789 10171
rect -2755 10137 -2721 10171
rect -2687 10137 -2653 10171
rect -2619 10137 -2585 10171
rect -2551 10137 -2517 10171
rect -2483 10137 -2449 10171
rect -2415 10137 -2381 10171
rect -2347 10137 -2313 10171
rect -2279 10137 -2245 10171
rect -2211 10137 -2177 10171
rect -2143 10137 -2109 10171
rect -2075 10137 -2041 10171
rect -2007 10137 -1973 10171
rect -1939 10137 -1905 10171
rect -1871 10137 -1837 10171
rect -1803 10137 -1769 10171
rect -1735 10137 -1701 10171
rect -1667 10137 -1633 10171
rect -1599 10137 -1565 10171
rect -1531 10137 -1497 10171
rect -1463 10137 -1429 10171
rect -1395 10137 -1361 10171
rect -1327 10137 -1293 10171
rect -1259 10137 -1225 10171
rect -1191 10137 -1157 10171
rect -1123 10137 -1089 10171
rect -1055 10137 -1021 10171
rect -987 10137 -953 10171
rect -919 10137 -885 10171
rect -851 10137 -817 10171
rect -783 10137 -749 10171
rect -715 10137 -681 10171
rect -647 10137 -613 10171
rect -579 10137 -545 10171
rect -511 10137 -477 10171
rect -443 10137 -409 10171
rect -375 10137 -341 10171
rect -307 10137 -273 10171
rect -2959 10068 -2925 10102
rect -2891 10068 -2857 10102
rect -2823 10068 -2789 10102
rect -2755 10068 -2721 10102
rect -2687 10068 -2653 10102
rect -2619 10068 -2585 10102
rect -2551 10068 -2517 10102
rect -2483 10068 -2449 10102
rect -2415 10068 -2381 10102
rect -2347 10068 -2313 10102
rect -2279 10068 -2245 10102
rect -2211 10068 -2177 10102
rect -2143 10068 -2109 10102
rect -2075 10068 -2041 10102
rect -2007 10068 -1973 10102
rect -1939 10068 -1905 10102
rect -1871 10068 -1837 10102
rect -1803 10068 -1769 10102
rect -1735 10068 -1701 10102
rect -1667 10068 -1633 10102
rect -1599 10068 -1565 10102
rect -1531 10068 -1497 10102
rect -1463 10068 -1429 10102
rect -1395 10068 -1361 10102
rect -1327 10068 -1293 10102
rect -1259 10068 -1225 10102
rect -1191 10068 -1157 10102
rect -1123 10068 -1089 10102
rect -1055 10068 -1021 10102
rect -987 10068 -953 10102
rect -919 10068 -885 10102
rect -851 10068 -817 10102
rect -783 10068 -749 10102
rect -715 10068 -681 10102
rect -647 10068 -613 10102
rect -579 10068 -545 10102
rect -511 10068 -477 10102
rect -443 10068 -409 10102
rect -375 10068 -341 10102
rect -307 10068 -273 10102
rect 13279 11880 13313 11914
rect 13347 11880 13381 11914
rect 13415 11880 13449 11914
rect 13483 11880 13517 11914
rect 13551 11880 13585 11914
rect 13619 11880 13653 11914
rect 13687 11880 13721 11914
rect 13755 11880 13789 11914
rect 13823 11880 13857 11914
rect 13891 11880 13925 11914
rect 13959 11880 13993 11914
rect 14027 11880 14061 11914
rect 14095 11880 14129 11914
rect 14163 11880 14197 11914
rect 14231 11880 14265 11914
rect 14299 11880 14333 11914
rect 14367 11880 14401 11914
rect 14435 11880 14469 11914
rect 14503 11880 14537 11914
rect 14571 11880 14605 11914
rect 14639 11880 14673 11914
rect 14707 11880 14741 11914
rect 14775 11880 14809 11914
rect 14843 11880 14877 11914
rect 14911 11880 14945 11914
rect 14979 11880 15013 11914
rect 15047 11880 15081 11914
rect 15115 11880 15149 11914
rect 15183 11880 15217 11914
rect 15251 11880 15285 11914
rect 15319 11880 15353 11914
rect 15387 11880 15421 11914
rect 15455 11880 15489 11914
rect 15523 11880 15557 11914
rect 15591 11880 15625 11914
rect 15659 11880 15693 11914
rect 15727 11880 15761 11914
rect 15795 11880 15829 11914
rect 13279 11811 13313 11845
rect 13347 11811 13381 11845
rect 13415 11811 13449 11845
rect 13483 11811 13517 11845
rect 13551 11811 13585 11845
rect 13619 11811 13653 11845
rect 13687 11811 13721 11845
rect 13755 11811 13789 11845
rect 13823 11811 13857 11845
rect 13891 11811 13925 11845
rect 13959 11811 13993 11845
rect 14027 11811 14061 11845
rect 14095 11811 14129 11845
rect 14163 11811 14197 11845
rect 14231 11811 14265 11845
rect 14299 11811 14333 11845
rect 14367 11811 14401 11845
rect 14435 11811 14469 11845
rect 14503 11811 14537 11845
rect 14571 11811 14605 11845
rect 14639 11811 14673 11845
rect 14707 11811 14741 11845
rect 14775 11811 14809 11845
rect 14843 11811 14877 11845
rect 14911 11811 14945 11845
rect 14979 11811 15013 11845
rect 15047 11811 15081 11845
rect 15115 11811 15149 11845
rect 15183 11811 15217 11845
rect 15251 11811 15285 11845
rect 15319 11811 15353 11845
rect 15387 11811 15421 11845
rect 15455 11811 15489 11845
rect 15523 11811 15557 11845
rect 15591 11811 15625 11845
rect 15659 11811 15693 11845
rect 15727 11811 15761 11845
rect 15795 11811 15829 11845
rect 13279 11742 13313 11776
rect 13347 11742 13381 11776
rect 13415 11742 13449 11776
rect 13483 11742 13517 11776
rect 13551 11742 13585 11776
rect 13619 11742 13653 11776
rect 13687 11742 13721 11776
rect 13755 11742 13789 11776
rect 13823 11742 13857 11776
rect 13891 11742 13925 11776
rect 13959 11742 13993 11776
rect 14027 11742 14061 11776
rect 14095 11742 14129 11776
rect 14163 11742 14197 11776
rect 14231 11742 14265 11776
rect 14299 11742 14333 11776
rect 14367 11742 14401 11776
rect 14435 11742 14469 11776
rect 14503 11742 14537 11776
rect 14571 11742 14605 11776
rect 14639 11742 14673 11776
rect 14707 11742 14741 11776
rect 14775 11742 14809 11776
rect 14843 11742 14877 11776
rect 14911 11742 14945 11776
rect 14979 11742 15013 11776
rect 15047 11742 15081 11776
rect 15115 11742 15149 11776
rect 15183 11742 15217 11776
rect 15251 11742 15285 11776
rect 15319 11742 15353 11776
rect 15387 11742 15421 11776
rect 15455 11742 15489 11776
rect 15523 11742 15557 11776
rect 15591 11742 15625 11776
rect 15659 11742 15693 11776
rect 15727 11742 15761 11776
rect 15795 11742 15829 11776
rect 13279 11673 13313 11707
rect 13347 11673 13381 11707
rect 13415 11673 13449 11707
rect 13483 11673 13517 11707
rect 13551 11673 13585 11707
rect 13619 11673 13653 11707
rect 13687 11673 13721 11707
rect 13755 11673 13789 11707
rect 13823 11673 13857 11707
rect 13891 11673 13925 11707
rect 13959 11673 13993 11707
rect 14027 11673 14061 11707
rect 14095 11673 14129 11707
rect 14163 11673 14197 11707
rect 14231 11673 14265 11707
rect 14299 11673 14333 11707
rect 14367 11673 14401 11707
rect 14435 11673 14469 11707
rect 14503 11673 14537 11707
rect 14571 11673 14605 11707
rect 14639 11673 14673 11707
rect 14707 11673 14741 11707
rect 14775 11673 14809 11707
rect 14843 11673 14877 11707
rect 14911 11673 14945 11707
rect 14979 11673 15013 11707
rect 15047 11673 15081 11707
rect 15115 11673 15149 11707
rect 15183 11673 15217 11707
rect 15251 11673 15285 11707
rect 15319 11673 15353 11707
rect 15387 11673 15421 11707
rect 15455 11673 15489 11707
rect 15523 11673 15557 11707
rect 15591 11673 15625 11707
rect 15659 11673 15693 11707
rect 15727 11673 15761 11707
rect 15795 11673 15829 11707
rect 13279 11604 13313 11638
rect 13347 11604 13381 11638
rect 13415 11604 13449 11638
rect 13483 11604 13517 11638
rect 13551 11604 13585 11638
rect 13619 11604 13653 11638
rect 13687 11604 13721 11638
rect 13755 11604 13789 11638
rect 13823 11604 13857 11638
rect 13891 11604 13925 11638
rect 13959 11604 13993 11638
rect 14027 11604 14061 11638
rect 14095 11604 14129 11638
rect 14163 11604 14197 11638
rect 14231 11604 14265 11638
rect 14299 11604 14333 11638
rect 14367 11604 14401 11638
rect 14435 11604 14469 11638
rect 14503 11604 14537 11638
rect 14571 11604 14605 11638
rect 14639 11604 14673 11638
rect 14707 11604 14741 11638
rect 14775 11604 14809 11638
rect 14843 11604 14877 11638
rect 14911 11604 14945 11638
rect 14979 11604 15013 11638
rect 15047 11604 15081 11638
rect 15115 11604 15149 11638
rect 15183 11604 15217 11638
rect 15251 11604 15285 11638
rect 15319 11604 15353 11638
rect 15387 11604 15421 11638
rect 15455 11604 15489 11638
rect 15523 11604 15557 11638
rect 15591 11604 15625 11638
rect 15659 11604 15693 11638
rect 15727 11604 15761 11638
rect 15795 11604 15829 11638
rect 13279 11535 13313 11569
rect 13347 11535 13381 11569
rect 13415 11535 13449 11569
rect 13483 11535 13517 11569
rect 13551 11535 13585 11569
rect 13619 11535 13653 11569
rect 13687 11535 13721 11569
rect 13755 11535 13789 11569
rect 13823 11535 13857 11569
rect 13891 11535 13925 11569
rect 13959 11535 13993 11569
rect 14027 11535 14061 11569
rect 14095 11535 14129 11569
rect 14163 11535 14197 11569
rect 14231 11535 14265 11569
rect 14299 11535 14333 11569
rect 14367 11535 14401 11569
rect 14435 11535 14469 11569
rect 14503 11535 14537 11569
rect 14571 11535 14605 11569
rect 14639 11535 14673 11569
rect 14707 11535 14741 11569
rect 14775 11535 14809 11569
rect 14843 11535 14877 11569
rect 14911 11535 14945 11569
rect 14979 11535 15013 11569
rect 15047 11535 15081 11569
rect 15115 11535 15149 11569
rect 15183 11535 15217 11569
rect 15251 11535 15285 11569
rect 15319 11535 15353 11569
rect 15387 11535 15421 11569
rect 15455 11535 15489 11569
rect 15523 11535 15557 11569
rect 15591 11535 15625 11569
rect 15659 11535 15693 11569
rect 15727 11535 15761 11569
rect 15795 11535 15829 11569
rect 13279 11465 13313 11499
rect 13347 11465 13381 11499
rect 13415 11465 13449 11499
rect 13483 11465 13517 11499
rect 13551 11465 13585 11499
rect 13619 11465 13653 11499
rect 13687 11465 13721 11499
rect 13755 11465 13789 11499
rect 13823 11465 13857 11499
rect 13891 11465 13925 11499
rect 13959 11465 13993 11499
rect 14027 11465 14061 11499
rect 14095 11465 14129 11499
rect 14163 11465 14197 11499
rect 14231 11465 14265 11499
rect 14299 11465 14333 11499
rect 14367 11465 14401 11499
rect 14435 11465 14469 11499
rect 14503 11465 14537 11499
rect 14571 11465 14605 11499
rect 14639 11465 14673 11499
rect 14707 11465 14741 11499
rect 14775 11465 14809 11499
rect 14843 11465 14877 11499
rect 14911 11465 14945 11499
rect 14979 11465 15013 11499
rect 15047 11465 15081 11499
rect 15115 11465 15149 11499
rect 15183 11465 15217 11499
rect 15251 11465 15285 11499
rect 15319 11465 15353 11499
rect 15387 11465 15421 11499
rect 15455 11465 15489 11499
rect 15523 11465 15557 11499
rect 15591 11465 15625 11499
rect 15659 11465 15693 11499
rect 15727 11465 15761 11499
rect 15795 11465 15829 11499
rect 13279 11395 13313 11429
rect 13347 11395 13381 11429
rect 13415 11395 13449 11429
rect 13483 11395 13517 11429
rect 13551 11395 13585 11429
rect 13619 11395 13653 11429
rect 13687 11395 13721 11429
rect 13755 11395 13789 11429
rect 13823 11395 13857 11429
rect 13891 11395 13925 11429
rect 13959 11395 13993 11429
rect 14027 11395 14061 11429
rect 14095 11395 14129 11429
rect 14163 11395 14197 11429
rect 14231 11395 14265 11429
rect 14299 11395 14333 11429
rect 14367 11395 14401 11429
rect 14435 11395 14469 11429
rect 14503 11395 14537 11429
rect 14571 11395 14605 11429
rect 14639 11395 14673 11429
rect 14707 11395 14741 11429
rect 14775 11395 14809 11429
rect 14843 11395 14877 11429
rect 14911 11395 14945 11429
rect 14979 11395 15013 11429
rect 15047 11395 15081 11429
rect 15115 11395 15149 11429
rect 15183 11395 15217 11429
rect 15251 11395 15285 11429
rect 15319 11395 15353 11429
rect 15387 11395 15421 11429
rect 15455 11395 15489 11429
rect 15523 11395 15557 11429
rect 15591 11395 15625 11429
rect 15659 11395 15693 11429
rect 15727 11395 15761 11429
rect 15795 11395 15829 11429
rect 13279 11325 13313 11359
rect 13347 11325 13381 11359
rect 13415 11325 13449 11359
rect 13483 11325 13517 11359
rect 13551 11325 13585 11359
rect 13619 11325 13653 11359
rect 13687 11325 13721 11359
rect 13755 11325 13789 11359
rect 13823 11325 13857 11359
rect 13891 11325 13925 11359
rect 13959 11325 13993 11359
rect 14027 11325 14061 11359
rect 14095 11325 14129 11359
rect 14163 11325 14197 11359
rect 14231 11325 14265 11359
rect 14299 11325 14333 11359
rect 14367 11325 14401 11359
rect 14435 11325 14469 11359
rect 14503 11325 14537 11359
rect 14571 11325 14605 11359
rect 14639 11325 14673 11359
rect 14707 11325 14741 11359
rect 14775 11325 14809 11359
rect 14843 11325 14877 11359
rect 14911 11325 14945 11359
rect 14979 11325 15013 11359
rect 15047 11325 15081 11359
rect 15115 11325 15149 11359
rect 15183 11325 15217 11359
rect 15251 11325 15285 11359
rect 15319 11325 15353 11359
rect 15387 11325 15421 11359
rect 15455 11325 15489 11359
rect 15523 11325 15557 11359
rect 15591 11325 15625 11359
rect 15659 11325 15693 11359
rect 15727 11325 15761 11359
rect 15795 11325 15829 11359
rect 13279 11255 13313 11289
rect 13347 11255 13381 11289
rect 13415 11255 13449 11289
rect 13483 11255 13517 11289
rect 13551 11255 13585 11289
rect 13619 11255 13653 11289
rect 13687 11255 13721 11289
rect 13755 11255 13789 11289
rect 13823 11255 13857 11289
rect 13891 11255 13925 11289
rect 13959 11255 13993 11289
rect 14027 11255 14061 11289
rect 14095 11255 14129 11289
rect 14163 11255 14197 11289
rect 14231 11255 14265 11289
rect 14299 11255 14333 11289
rect 14367 11255 14401 11289
rect 14435 11255 14469 11289
rect 14503 11255 14537 11289
rect 14571 11255 14605 11289
rect 14639 11255 14673 11289
rect 14707 11255 14741 11289
rect 14775 11255 14809 11289
rect 14843 11255 14877 11289
rect 14911 11255 14945 11289
rect 14979 11255 15013 11289
rect 15047 11255 15081 11289
rect 15115 11255 15149 11289
rect 15183 11255 15217 11289
rect 15251 11255 15285 11289
rect 15319 11255 15353 11289
rect 15387 11255 15421 11289
rect 15455 11255 15489 11289
rect 15523 11255 15557 11289
rect 15591 11255 15625 11289
rect 15659 11255 15693 11289
rect 15727 11255 15761 11289
rect 15795 11255 15829 11289
rect 13279 11185 13313 11219
rect 13347 11185 13381 11219
rect 13415 11185 13449 11219
rect 13483 11185 13517 11219
rect 13551 11185 13585 11219
rect 13619 11185 13653 11219
rect 13687 11185 13721 11219
rect 13755 11185 13789 11219
rect 13823 11185 13857 11219
rect 13891 11185 13925 11219
rect 13959 11185 13993 11219
rect 14027 11185 14061 11219
rect 14095 11185 14129 11219
rect 14163 11185 14197 11219
rect 14231 11185 14265 11219
rect 14299 11185 14333 11219
rect 14367 11185 14401 11219
rect 14435 11185 14469 11219
rect 14503 11185 14537 11219
rect 14571 11185 14605 11219
rect 14639 11185 14673 11219
rect 14707 11185 14741 11219
rect 14775 11185 14809 11219
rect 14843 11185 14877 11219
rect 14911 11185 14945 11219
rect 14979 11185 15013 11219
rect 15047 11185 15081 11219
rect 15115 11185 15149 11219
rect 15183 11185 15217 11219
rect 15251 11185 15285 11219
rect 15319 11185 15353 11219
rect 15387 11185 15421 11219
rect 15455 11185 15489 11219
rect 15523 11185 15557 11219
rect 15591 11185 15625 11219
rect 15659 11185 15693 11219
rect 15727 11185 15761 11219
rect 15795 11185 15829 11219
rect 13279 11115 13313 11149
rect 13347 11115 13381 11149
rect 13415 11115 13449 11149
rect 13483 11115 13517 11149
rect 13551 11115 13585 11149
rect 13619 11115 13653 11149
rect 13687 11115 13721 11149
rect 13755 11115 13789 11149
rect 13823 11115 13857 11149
rect 13891 11115 13925 11149
rect 13959 11115 13993 11149
rect 14027 11115 14061 11149
rect 14095 11115 14129 11149
rect 14163 11115 14197 11149
rect 14231 11115 14265 11149
rect 14299 11115 14333 11149
rect 14367 11115 14401 11149
rect 14435 11115 14469 11149
rect 14503 11115 14537 11149
rect 14571 11115 14605 11149
rect 14639 11115 14673 11149
rect 14707 11115 14741 11149
rect 14775 11115 14809 11149
rect 14843 11115 14877 11149
rect 14911 11115 14945 11149
rect 14979 11115 15013 11149
rect 15047 11115 15081 11149
rect 15115 11115 15149 11149
rect 15183 11115 15217 11149
rect 15251 11115 15285 11149
rect 15319 11115 15353 11149
rect 15387 11115 15421 11149
rect 15455 11115 15489 11149
rect 15523 11115 15557 11149
rect 15591 11115 15625 11149
rect 15659 11115 15693 11149
rect 15727 11115 15761 11149
rect 15795 11115 15829 11149
rect 13279 11045 13313 11079
rect 13347 11045 13381 11079
rect 13415 11045 13449 11079
rect 13483 11045 13517 11079
rect 13551 11045 13585 11079
rect 13619 11045 13653 11079
rect 13687 11045 13721 11079
rect 13755 11045 13789 11079
rect 13823 11045 13857 11079
rect 13891 11045 13925 11079
rect 13959 11045 13993 11079
rect 14027 11045 14061 11079
rect 14095 11045 14129 11079
rect 14163 11045 14197 11079
rect 14231 11045 14265 11079
rect 14299 11045 14333 11079
rect 14367 11045 14401 11079
rect 14435 11045 14469 11079
rect 14503 11045 14537 11079
rect 14571 11045 14605 11079
rect 14639 11045 14673 11079
rect 14707 11045 14741 11079
rect 14775 11045 14809 11079
rect 14843 11045 14877 11079
rect 14911 11045 14945 11079
rect 14979 11045 15013 11079
rect 15047 11045 15081 11079
rect 15115 11045 15149 11079
rect 15183 11045 15217 11079
rect 15251 11045 15285 11079
rect 15319 11045 15353 11079
rect 15387 11045 15421 11079
rect 15455 11045 15489 11079
rect 15523 11045 15557 11079
rect 15591 11045 15625 11079
rect 15659 11045 15693 11079
rect 15727 11045 15761 11079
rect 15795 11045 15829 11079
rect 13279 10975 13313 11009
rect 13347 10975 13381 11009
rect 13415 10975 13449 11009
rect 13483 10975 13517 11009
rect 13551 10975 13585 11009
rect 13619 10975 13653 11009
rect 13687 10975 13721 11009
rect 13755 10975 13789 11009
rect 13823 10975 13857 11009
rect 13891 10975 13925 11009
rect 13959 10975 13993 11009
rect 14027 10975 14061 11009
rect 14095 10975 14129 11009
rect 14163 10975 14197 11009
rect 14231 10975 14265 11009
rect 14299 10975 14333 11009
rect 14367 10975 14401 11009
rect 14435 10975 14469 11009
rect 14503 10975 14537 11009
rect 14571 10975 14605 11009
rect 14639 10975 14673 11009
rect 14707 10975 14741 11009
rect 14775 10975 14809 11009
rect 14843 10975 14877 11009
rect 14911 10975 14945 11009
rect 14979 10975 15013 11009
rect 15047 10975 15081 11009
rect 15115 10975 15149 11009
rect 15183 10975 15217 11009
rect 15251 10975 15285 11009
rect 15319 10975 15353 11009
rect 15387 10975 15421 11009
rect 15455 10975 15489 11009
rect 15523 10975 15557 11009
rect 15591 10975 15625 11009
rect 15659 10975 15693 11009
rect 15727 10975 15761 11009
rect 15795 10975 15829 11009
rect 13279 10905 13313 10939
rect 13347 10905 13381 10939
rect 13415 10905 13449 10939
rect 13483 10905 13517 10939
rect 13551 10905 13585 10939
rect 13619 10905 13653 10939
rect 13687 10905 13721 10939
rect 13755 10905 13789 10939
rect 13823 10905 13857 10939
rect 13891 10905 13925 10939
rect 13959 10905 13993 10939
rect 14027 10905 14061 10939
rect 14095 10905 14129 10939
rect 14163 10905 14197 10939
rect 14231 10905 14265 10939
rect 14299 10905 14333 10939
rect 14367 10905 14401 10939
rect 14435 10905 14469 10939
rect 14503 10905 14537 10939
rect 14571 10905 14605 10939
rect 14639 10905 14673 10939
rect 14707 10905 14741 10939
rect 14775 10905 14809 10939
rect 14843 10905 14877 10939
rect 14911 10905 14945 10939
rect 14979 10905 15013 10939
rect 15047 10905 15081 10939
rect 15115 10905 15149 10939
rect 15183 10905 15217 10939
rect 15251 10905 15285 10939
rect 15319 10905 15353 10939
rect 15387 10905 15421 10939
rect 15455 10905 15489 10939
rect 15523 10905 15557 10939
rect 15591 10905 15625 10939
rect 15659 10905 15693 10939
rect 15727 10905 15761 10939
rect 15795 10905 15829 10939
rect 13279 10835 13313 10869
rect 13347 10835 13381 10869
rect 13415 10835 13449 10869
rect 13483 10835 13517 10869
rect 13551 10835 13585 10869
rect 13619 10835 13653 10869
rect 13687 10835 13721 10869
rect 13755 10835 13789 10869
rect 13823 10835 13857 10869
rect 13891 10835 13925 10869
rect 13959 10835 13993 10869
rect 14027 10835 14061 10869
rect 14095 10835 14129 10869
rect 14163 10835 14197 10869
rect 14231 10835 14265 10869
rect 14299 10835 14333 10869
rect 14367 10835 14401 10869
rect 14435 10835 14469 10869
rect 14503 10835 14537 10869
rect 14571 10835 14605 10869
rect 14639 10835 14673 10869
rect 14707 10835 14741 10869
rect 14775 10835 14809 10869
rect 14843 10835 14877 10869
rect 14911 10835 14945 10869
rect 14979 10835 15013 10869
rect 15047 10835 15081 10869
rect 15115 10835 15149 10869
rect 15183 10835 15217 10869
rect 15251 10835 15285 10869
rect 15319 10835 15353 10869
rect 15387 10835 15421 10869
rect 15455 10835 15489 10869
rect 15523 10835 15557 10869
rect 15591 10835 15625 10869
rect 15659 10835 15693 10869
rect 15727 10835 15761 10869
rect 15795 10835 15829 10869
rect 13279 10765 13313 10799
rect 13347 10765 13381 10799
rect 13415 10765 13449 10799
rect 13483 10765 13517 10799
rect 13551 10765 13585 10799
rect 13619 10765 13653 10799
rect 13687 10765 13721 10799
rect 13755 10765 13789 10799
rect 13823 10765 13857 10799
rect 13891 10765 13925 10799
rect 13959 10765 13993 10799
rect 14027 10765 14061 10799
rect 14095 10765 14129 10799
rect 14163 10765 14197 10799
rect 14231 10765 14265 10799
rect 14299 10765 14333 10799
rect 14367 10765 14401 10799
rect 14435 10765 14469 10799
rect 14503 10765 14537 10799
rect 14571 10765 14605 10799
rect 14639 10765 14673 10799
rect 14707 10765 14741 10799
rect 14775 10765 14809 10799
rect 14843 10765 14877 10799
rect 14911 10765 14945 10799
rect 14979 10765 15013 10799
rect 15047 10765 15081 10799
rect 15115 10765 15149 10799
rect 15183 10765 15217 10799
rect 15251 10765 15285 10799
rect 15319 10765 15353 10799
rect 15387 10765 15421 10799
rect 15455 10765 15489 10799
rect 15523 10765 15557 10799
rect 15591 10765 15625 10799
rect 15659 10765 15693 10799
rect 15727 10765 15761 10799
rect 15795 10765 15829 10799
rect 13279 10695 13313 10729
rect 13347 10695 13381 10729
rect 13415 10695 13449 10729
rect 13483 10695 13517 10729
rect 13551 10695 13585 10729
rect 13619 10695 13653 10729
rect 13687 10695 13721 10729
rect 13755 10695 13789 10729
rect 13823 10695 13857 10729
rect 13891 10695 13925 10729
rect 13959 10695 13993 10729
rect 14027 10695 14061 10729
rect 14095 10695 14129 10729
rect 14163 10695 14197 10729
rect 14231 10695 14265 10729
rect 14299 10695 14333 10729
rect 14367 10695 14401 10729
rect 14435 10695 14469 10729
rect 14503 10695 14537 10729
rect 14571 10695 14605 10729
rect 14639 10695 14673 10729
rect 14707 10695 14741 10729
rect 14775 10695 14809 10729
rect 14843 10695 14877 10729
rect 14911 10695 14945 10729
rect 14979 10695 15013 10729
rect 15047 10695 15081 10729
rect 15115 10695 15149 10729
rect 15183 10695 15217 10729
rect 15251 10695 15285 10729
rect 15319 10695 15353 10729
rect 15387 10695 15421 10729
rect 15455 10695 15489 10729
rect 15523 10695 15557 10729
rect 15591 10695 15625 10729
rect 15659 10695 15693 10729
rect 15727 10695 15761 10729
rect 15795 10695 15829 10729
rect 13279 10625 13313 10659
rect 13347 10625 13381 10659
rect 13415 10625 13449 10659
rect 13483 10625 13517 10659
rect 13551 10625 13585 10659
rect 13619 10625 13653 10659
rect 13687 10625 13721 10659
rect 13755 10625 13789 10659
rect 13823 10625 13857 10659
rect 13891 10625 13925 10659
rect 13959 10625 13993 10659
rect 14027 10625 14061 10659
rect 14095 10625 14129 10659
rect 14163 10625 14197 10659
rect 14231 10625 14265 10659
rect 14299 10625 14333 10659
rect 14367 10625 14401 10659
rect 14435 10625 14469 10659
rect 14503 10625 14537 10659
rect 14571 10625 14605 10659
rect 14639 10625 14673 10659
rect 14707 10625 14741 10659
rect 14775 10625 14809 10659
rect 14843 10625 14877 10659
rect 14911 10625 14945 10659
rect 14979 10625 15013 10659
rect 15047 10625 15081 10659
rect 15115 10625 15149 10659
rect 15183 10625 15217 10659
rect 15251 10625 15285 10659
rect 15319 10625 15353 10659
rect 15387 10625 15421 10659
rect 15455 10625 15489 10659
rect 15523 10625 15557 10659
rect 15591 10625 15625 10659
rect 15659 10625 15693 10659
rect 15727 10625 15761 10659
rect 15795 10625 15829 10659
rect 13279 10555 13313 10589
rect 13347 10555 13381 10589
rect 13415 10555 13449 10589
rect 13483 10555 13517 10589
rect 13551 10555 13585 10589
rect 13619 10555 13653 10589
rect 13687 10555 13721 10589
rect 13755 10555 13789 10589
rect 13823 10555 13857 10589
rect 13891 10555 13925 10589
rect 13959 10555 13993 10589
rect 14027 10555 14061 10589
rect 14095 10555 14129 10589
rect 14163 10555 14197 10589
rect 14231 10555 14265 10589
rect 14299 10555 14333 10589
rect 14367 10555 14401 10589
rect 14435 10555 14469 10589
rect 14503 10555 14537 10589
rect 14571 10555 14605 10589
rect 14639 10555 14673 10589
rect 14707 10555 14741 10589
rect 14775 10555 14809 10589
rect 14843 10555 14877 10589
rect 14911 10555 14945 10589
rect 14979 10555 15013 10589
rect 15047 10555 15081 10589
rect 15115 10555 15149 10589
rect 15183 10555 15217 10589
rect 15251 10555 15285 10589
rect 15319 10555 15353 10589
rect 15387 10555 15421 10589
rect 15455 10555 15489 10589
rect 15523 10555 15557 10589
rect 15591 10555 15625 10589
rect 15659 10555 15693 10589
rect 15727 10555 15761 10589
rect 15795 10555 15829 10589
rect 13279 10485 13313 10519
rect 13347 10485 13381 10519
rect 13415 10485 13449 10519
rect 13483 10485 13517 10519
rect 13551 10485 13585 10519
rect 13619 10485 13653 10519
rect 13687 10485 13721 10519
rect 13755 10485 13789 10519
rect 13823 10485 13857 10519
rect 13891 10485 13925 10519
rect 13959 10485 13993 10519
rect 14027 10485 14061 10519
rect 14095 10485 14129 10519
rect 14163 10485 14197 10519
rect 14231 10485 14265 10519
rect 14299 10485 14333 10519
rect 14367 10485 14401 10519
rect 14435 10485 14469 10519
rect 14503 10485 14537 10519
rect 14571 10485 14605 10519
rect 14639 10485 14673 10519
rect 14707 10485 14741 10519
rect 14775 10485 14809 10519
rect 14843 10485 14877 10519
rect 14911 10485 14945 10519
rect 14979 10485 15013 10519
rect 15047 10485 15081 10519
rect 15115 10485 15149 10519
rect 15183 10485 15217 10519
rect 15251 10485 15285 10519
rect 15319 10485 15353 10519
rect 15387 10485 15421 10519
rect 15455 10485 15489 10519
rect 15523 10485 15557 10519
rect 15591 10485 15625 10519
rect 15659 10485 15693 10519
rect 15727 10485 15761 10519
rect 15795 10485 15829 10519
rect 13279 10415 13313 10449
rect 13347 10415 13381 10449
rect 13415 10415 13449 10449
rect 13483 10415 13517 10449
rect 13551 10415 13585 10449
rect 13619 10415 13653 10449
rect 13687 10415 13721 10449
rect 13755 10415 13789 10449
rect 13823 10415 13857 10449
rect 13891 10415 13925 10449
rect 13959 10415 13993 10449
rect 14027 10415 14061 10449
rect 14095 10415 14129 10449
rect 14163 10415 14197 10449
rect 14231 10415 14265 10449
rect 14299 10415 14333 10449
rect 14367 10415 14401 10449
rect 14435 10415 14469 10449
rect 14503 10415 14537 10449
rect 14571 10415 14605 10449
rect 14639 10415 14673 10449
rect 14707 10415 14741 10449
rect 14775 10415 14809 10449
rect 14843 10415 14877 10449
rect 14911 10415 14945 10449
rect 14979 10415 15013 10449
rect 15047 10415 15081 10449
rect 15115 10415 15149 10449
rect 15183 10415 15217 10449
rect 15251 10415 15285 10449
rect 15319 10415 15353 10449
rect 15387 10415 15421 10449
rect 15455 10415 15489 10449
rect 15523 10415 15557 10449
rect 15591 10415 15625 10449
rect 15659 10415 15693 10449
rect 15727 10415 15761 10449
rect 15795 10415 15829 10449
rect 13279 10345 13313 10379
rect 13347 10345 13381 10379
rect 13415 10345 13449 10379
rect 13483 10345 13517 10379
rect 13551 10345 13585 10379
rect 13619 10345 13653 10379
rect 13687 10345 13721 10379
rect 13755 10345 13789 10379
rect 13823 10345 13857 10379
rect 13891 10345 13925 10379
rect 13959 10345 13993 10379
rect 14027 10345 14061 10379
rect 14095 10345 14129 10379
rect 14163 10345 14197 10379
rect 14231 10345 14265 10379
rect 14299 10345 14333 10379
rect 14367 10345 14401 10379
rect 14435 10345 14469 10379
rect 14503 10345 14537 10379
rect 14571 10345 14605 10379
rect 14639 10345 14673 10379
rect 14707 10345 14741 10379
rect 14775 10345 14809 10379
rect 14843 10345 14877 10379
rect 14911 10345 14945 10379
rect 14979 10345 15013 10379
rect 15047 10345 15081 10379
rect 15115 10345 15149 10379
rect 15183 10345 15217 10379
rect 15251 10345 15285 10379
rect 15319 10345 15353 10379
rect 15387 10345 15421 10379
rect 15455 10345 15489 10379
rect 15523 10345 15557 10379
rect 15591 10345 15625 10379
rect 15659 10345 15693 10379
rect 15727 10345 15761 10379
rect 15795 10345 15829 10379
rect 13279 10275 13313 10309
rect 13347 10275 13381 10309
rect 13415 10275 13449 10309
rect 13483 10275 13517 10309
rect 13551 10275 13585 10309
rect 13619 10275 13653 10309
rect 13687 10275 13721 10309
rect 13755 10275 13789 10309
rect 13823 10275 13857 10309
rect 13891 10275 13925 10309
rect 13959 10275 13993 10309
rect 14027 10275 14061 10309
rect 14095 10275 14129 10309
rect 14163 10275 14197 10309
rect 14231 10275 14265 10309
rect 14299 10275 14333 10309
rect 14367 10275 14401 10309
rect 14435 10275 14469 10309
rect 14503 10275 14537 10309
rect 14571 10275 14605 10309
rect 14639 10275 14673 10309
rect 14707 10275 14741 10309
rect 14775 10275 14809 10309
rect 14843 10275 14877 10309
rect 14911 10275 14945 10309
rect 14979 10275 15013 10309
rect 15047 10275 15081 10309
rect 15115 10275 15149 10309
rect 15183 10275 15217 10309
rect 15251 10275 15285 10309
rect 15319 10275 15353 10309
rect 15387 10275 15421 10309
rect 15455 10275 15489 10309
rect 15523 10275 15557 10309
rect 15591 10275 15625 10309
rect 15659 10275 15693 10309
rect 15727 10275 15761 10309
rect 15795 10275 15829 10309
rect 13279 10205 13313 10239
rect 13347 10205 13381 10239
rect 13415 10205 13449 10239
rect 13483 10205 13517 10239
rect 13551 10205 13585 10239
rect 13619 10205 13653 10239
rect 13687 10205 13721 10239
rect 13755 10205 13789 10239
rect 13823 10205 13857 10239
rect 13891 10205 13925 10239
rect 13959 10205 13993 10239
rect 14027 10205 14061 10239
rect 14095 10205 14129 10239
rect 14163 10205 14197 10239
rect 14231 10205 14265 10239
rect 14299 10205 14333 10239
rect 14367 10205 14401 10239
rect 14435 10205 14469 10239
rect 14503 10205 14537 10239
rect 14571 10205 14605 10239
rect 14639 10205 14673 10239
rect 14707 10205 14741 10239
rect 14775 10205 14809 10239
rect 14843 10205 14877 10239
rect 14911 10205 14945 10239
rect 14979 10205 15013 10239
rect 15047 10205 15081 10239
rect 15115 10205 15149 10239
rect 15183 10205 15217 10239
rect 15251 10205 15285 10239
rect 15319 10205 15353 10239
rect 15387 10205 15421 10239
rect 15455 10205 15489 10239
rect 15523 10205 15557 10239
rect 15591 10205 15625 10239
rect 15659 10205 15693 10239
rect 15727 10205 15761 10239
rect 15795 10205 15829 10239
rect 12504 10128 12538 10162
rect 12599 10128 12633 10162
rect 12694 10128 12728 10162
rect 12788 10128 12822 10162
rect 12882 10128 12916 10162
rect 12976 10128 13010 10162
rect 13279 10135 13313 10169
rect 13347 10135 13381 10169
rect 13415 10135 13449 10169
rect 13483 10135 13517 10169
rect 13551 10135 13585 10169
rect 13619 10135 13653 10169
rect 13687 10135 13721 10169
rect 13755 10135 13789 10169
rect 13823 10135 13857 10169
rect 13891 10135 13925 10169
rect 13959 10135 13993 10169
rect 14027 10135 14061 10169
rect 14095 10135 14129 10169
rect 14163 10135 14197 10169
rect 14231 10135 14265 10169
rect 14299 10135 14333 10169
rect 14367 10135 14401 10169
rect 14435 10135 14469 10169
rect 14503 10135 14537 10169
rect 14571 10135 14605 10169
rect 14639 10135 14673 10169
rect 14707 10135 14741 10169
rect 14775 10135 14809 10169
rect 14843 10135 14877 10169
rect 14911 10135 14945 10169
rect 14979 10135 15013 10169
rect 15047 10135 15081 10169
rect 15115 10135 15149 10169
rect 15183 10135 15217 10169
rect 15251 10135 15285 10169
rect 15319 10135 15353 10169
rect 15387 10135 15421 10169
rect 15455 10135 15489 10169
rect 15523 10135 15557 10169
rect 15591 10135 15625 10169
rect 15659 10135 15693 10169
rect 15727 10135 15761 10169
rect 15795 10135 15829 10169
rect -2959 9999 -2925 10033
rect -2891 9999 -2857 10033
rect -2823 9999 -2789 10033
rect -2755 9999 -2721 10033
rect -2687 9999 -2653 10033
rect -2619 9999 -2585 10033
rect -2551 9999 -2517 10033
rect -2483 9999 -2449 10033
rect -2415 9999 -2381 10033
rect -2347 9999 -2313 10033
rect -2279 9999 -2245 10033
rect -2211 9999 -2177 10033
rect -2143 9999 -2109 10033
rect -2075 9999 -2041 10033
rect -2007 9999 -1973 10033
rect -1939 9999 -1905 10033
rect -1871 9999 -1837 10033
rect -1803 9999 -1769 10033
rect -1735 9999 -1701 10033
rect -1667 9999 -1633 10033
rect -1599 9999 -1565 10033
rect -1531 9999 -1497 10033
rect -1463 9999 -1429 10033
rect -1395 9999 -1361 10033
rect -1327 9999 -1293 10033
rect -1259 9999 -1225 10033
rect -1191 9999 -1157 10033
rect -1123 9999 -1089 10033
rect -1055 9999 -1021 10033
rect -987 9999 -953 10033
rect -919 9999 -885 10033
rect -851 9999 -817 10033
rect -783 9999 -749 10033
rect -715 9999 -681 10033
rect -647 9999 -613 10033
rect -579 9999 -545 10033
rect -511 9999 -477 10033
rect -443 9999 -409 10033
rect -375 9999 -341 10033
rect -307 9999 -273 10033
rect -2959 9930 -2925 9964
rect -2891 9930 -2857 9964
rect -2823 9930 -2789 9964
rect -2755 9930 -2721 9964
rect -2687 9930 -2653 9964
rect -2619 9930 -2585 9964
rect -2551 9930 -2517 9964
rect -2483 9930 -2449 9964
rect -2415 9930 -2381 9964
rect -2347 9930 -2313 9964
rect -2279 9930 -2245 9964
rect -2211 9930 -2177 9964
rect -2143 9930 -2109 9964
rect -2075 9930 -2041 9964
rect -2007 9930 -1973 9964
rect -1939 9930 -1905 9964
rect -1871 9930 -1837 9964
rect -1803 9930 -1769 9964
rect -1735 9930 -1701 9964
rect -1667 9930 -1633 9964
rect -1599 9930 -1565 9964
rect -1531 9930 -1497 9964
rect -1463 9930 -1429 9964
rect -1395 9930 -1361 9964
rect -1327 9930 -1293 9964
rect -1259 9930 -1225 9964
rect -1191 9930 -1157 9964
rect -1123 9930 -1089 9964
rect -1055 9930 -1021 9964
rect -987 9930 -953 9964
rect -919 9930 -885 9964
rect -851 9930 -817 9964
rect -783 9930 -749 9964
rect -715 9930 -681 9964
rect -647 9930 -613 9964
rect -579 9930 -545 9964
rect -511 9930 -477 9964
rect -443 9930 -409 9964
rect -375 9930 -341 9964
rect -307 9930 -273 9964
rect 12504 10060 12538 10094
rect 12599 10060 12633 10094
rect 12694 10060 12728 10094
rect 12788 10060 12822 10094
rect 12882 10060 12916 10094
rect 12976 10060 13010 10094
rect 13279 10065 13313 10099
rect 13347 10065 13381 10099
rect 13415 10065 13449 10099
rect 13483 10065 13517 10099
rect 13551 10065 13585 10099
rect 13619 10065 13653 10099
rect 13687 10065 13721 10099
rect 13755 10065 13789 10099
rect 13823 10065 13857 10099
rect 13891 10065 13925 10099
rect 13959 10065 13993 10099
rect 14027 10065 14061 10099
rect 14095 10065 14129 10099
rect 14163 10065 14197 10099
rect 14231 10065 14265 10099
rect 14299 10065 14333 10099
rect 14367 10065 14401 10099
rect 14435 10065 14469 10099
rect 14503 10065 14537 10099
rect 14571 10065 14605 10099
rect 14639 10065 14673 10099
rect 14707 10065 14741 10099
rect 14775 10065 14809 10099
rect 14843 10065 14877 10099
rect 14911 10065 14945 10099
rect 14979 10065 15013 10099
rect 15047 10065 15081 10099
rect 15115 10065 15149 10099
rect 15183 10065 15217 10099
rect 15251 10065 15285 10099
rect 15319 10065 15353 10099
rect 15387 10065 15421 10099
rect 15455 10065 15489 10099
rect 15523 10065 15557 10099
rect 15591 10065 15625 10099
rect 15659 10065 15693 10099
rect 15727 10065 15761 10099
rect 15795 10065 15829 10099
rect 12504 9992 12538 10026
rect 12599 9992 12633 10026
rect 12694 9992 12728 10026
rect 12788 9992 12822 10026
rect 12882 9992 12916 10026
rect 12976 9992 13010 10026
rect 13077 10022 13111 10056
rect 13160 10022 13194 10056
rect 13279 9995 13313 10029
rect 13347 9995 13381 10029
rect 13415 9995 13449 10029
rect 13483 9995 13517 10029
rect 13551 9995 13585 10029
rect 13619 9995 13653 10029
rect 13687 9995 13721 10029
rect 13755 9995 13789 10029
rect 13823 9995 13857 10029
rect 13891 9995 13925 10029
rect 13959 9995 13993 10029
rect 14027 9995 14061 10029
rect 14095 9995 14129 10029
rect 14163 9995 14197 10029
rect 14231 9995 14265 10029
rect 14299 9995 14333 10029
rect 14367 9995 14401 10029
rect 14435 9995 14469 10029
rect 14503 9995 14537 10029
rect 14571 9995 14605 10029
rect 14639 9995 14673 10029
rect 14707 9995 14741 10029
rect 14775 9995 14809 10029
rect 14843 9995 14877 10029
rect 14911 9995 14945 10029
rect 14979 9995 15013 10029
rect 15047 9995 15081 10029
rect 15115 9995 15149 10029
rect 15183 9995 15217 10029
rect 15251 9995 15285 10029
rect 15319 9995 15353 10029
rect 15387 9995 15421 10029
rect 15455 9995 15489 10029
rect 15523 9995 15557 10029
rect 15591 9995 15625 10029
rect 15659 9995 15693 10029
rect 15727 9995 15761 10029
rect 15795 9995 15829 10029
rect -2959 9861 -2925 9895
rect -2891 9861 -2857 9895
rect -2823 9861 -2789 9895
rect -2755 9861 -2721 9895
rect -2687 9861 -2653 9895
rect -2619 9861 -2585 9895
rect -2551 9861 -2517 9895
rect -2483 9861 -2449 9895
rect -2415 9861 -2381 9895
rect -2347 9861 -2313 9895
rect -2279 9861 -2245 9895
rect -2211 9861 -2177 9895
rect -2143 9861 -2109 9895
rect -2075 9861 -2041 9895
rect -2007 9861 -1973 9895
rect -1939 9861 -1905 9895
rect -1871 9861 -1837 9895
rect -1803 9861 -1769 9895
rect -1735 9861 -1701 9895
rect -1667 9861 -1633 9895
rect -1599 9861 -1565 9895
rect -1531 9861 -1497 9895
rect -1463 9861 -1429 9895
rect -1395 9861 -1361 9895
rect -1327 9861 -1293 9895
rect -1259 9861 -1225 9895
rect -1191 9861 -1157 9895
rect -1123 9861 -1089 9895
rect -1055 9861 -1021 9895
rect -987 9861 -953 9895
rect -919 9861 -885 9895
rect -851 9861 -817 9895
rect -783 9861 -749 9895
rect -715 9861 -681 9895
rect -647 9861 -613 9895
rect -579 9861 -545 9895
rect -511 9861 -477 9895
rect -443 9861 -409 9895
rect -375 9861 -341 9895
rect -307 9861 -273 9895
rect -2959 9792 -2925 9826
rect -2891 9792 -2857 9826
rect -2823 9792 -2789 9826
rect -2755 9792 -2721 9826
rect -2687 9792 -2653 9826
rect -2619 9792 -2585 9826
rect -2551 9792 -2517 9826
rect -2483 9792 -2449 9826
rect -2415 9792 -2381 9826
rect -2347 9792 -2313 9826
rect -2279 9792 -2245 9826
rect -2211 9792 -2177 9826
rect -2143 9792 -2109 9826
rect -2075 9792 -2041 9826
rect -2007 9792 -1973 9826
rect -1939 9792 -1905 9826
rect -1871 9792 -1837 9826
rect -1803 9792 -1769 9826
rect -1735 9792 -1701 9826
rect -1667 9792 -1633 9826
rect -1599 9792 -1565 9826
rect -1531 9792 -1497 9826
rect -1463 9792 -1429 9826
rect -1395 9792 -1361 9826
rect -1327 9792 -1293 9826
rect -1259 9792 -1225 9826
rect -1191 9792 -1157 9826
rect -1123 9792 -1089 9826
rect -1055 9792 -1021 9826
rect -987 9792 -953 9826
rect -919 9792 -885 9826
rect -851 9792 -817 9826
rect -783 9792 -749 9826
rect -715 9792 -681 9826
rect -647 9792 -613 9826
rect -579 9792 -545 9826
rect -511 9792 -477 9826
rect -443 9792 -409 9826
rect -375 9792 -341 9826
rect -307 9792 -273 9826
rect -2959 9723 -2925 9757
rect -2891 9723 -2857 9757
rect -2823 9723 -2789 9757
rect -2755 9723 -2721 9757
rect -2687 9723 -2653 9757
rect -2619 9723 -2585 9757
rect -2551 9723 -2517 9757
rect -2483 9723 -2449 9757
rect -2415 9723 -2381 9757
rect -2347 9723 -2313 9757
rect -2279 9723 -2245 9757
rect -2211 9723 -2177 9757
rect -2143 9723 -2109 9757
rect -2075 9723 -2041 9757
rect -2007 9723 -1973 9757
rect -1939 9723 -1905 9757
rect -1871 9723 -1837 9757
rect -1803 9723 -1769 9757
rect -1735 9723 -1701 9757
rect -1667 9723 -1633 9757
rect -1599 9723 -1565 9757
rect -1531 9723 -1497 9757
rect -1463 9723 -1429 9757
rect -1395 9723 -1361 9757
rect -1327 9723 -1293 9757
rect -1259 9723 -1225 9757
rect -1191 9723 -1157 9757
rect -1123 9723 -1089 9757
rect -1055 9723 -1021 9757
rect -987 9723 -953 9757
rect -919 9723 -885 9757
rect -851 9723 -817 9757
rect -783 9723 -749 9757
rect -715 9723 -681 9757
rect -647 9723 -613 9757
rect -579 9723 -545 9757
rect -511 9723 -477 9757
rect -443 9723 -409 9757
rect -375 9723 -341 9757
rect -307 9723 -273 9757
rect -2959 9654 -2925 9688
rect -2891 9654 -2857 9688
rect -2823 9654 -2789 9688
rect -2755 9654 -2721 9688
rect -2687 9654 -2653 9688
rect -2619 9654 -2585 9688
rect -2551 9654 -2517 9688
rect -2483 9654 -2449 9688
rect -2415 9654 -2381 9688
rect -2347 9654 -2313 9688
rect -2279 9654 -2245 9688
rect -2211 9654 -2177 9688
rect -2143 9654 -2109 9688
rect -2075 9654 -2041 9688
rect -2007 9654 -1973 9688
rect -1939 9654 -1905 9688
rect -1871 9654 -1837 9688
rect -1803 9654 -1769 9688
rect -1735 9654 -1701 9688
rect -1667 9654 -1633 9688
rect -1599 9654 -1565 9688
rect -1531 9654 -1497 9688
rect -1463 9654 -1429 9688
rect -1395 9654 -1361 9688
rect -1327 9654 -1293 9688
rect -1259 9654 -1225 9688
rect -1191 9654 -1157 9688
rect -1123 9654 -1089 9688
rect -1055 9654 -1021 9688
rect -987 9654 -953 9688
rect -919 9654 -885 9688
rect -851 9654 -817 9688
rect -783 9654 -749 9688
rect -715 9654 -681 9688
rect -647 9654 -613 9688
rect -579 9654 -545 9688
rect -511 9654 -477 9688
rect -443 9654 -409 9688
rect -375 9654 -341 9688
rect -307 9654 -273 9688
rect -2959 9585 -2925 9619
rect -2891 9585 -2857 9619
rect -2823 9585 -2789 9619
rect -2755 9585 -2721 9619
rect -2687 9585 -2653 9619
rect -2619 9585 -2585 9619
rect -2551 9585 -2517 9619
rect -2483 9585 -2449 9619
rect -2415 9585 -2381 9619
rect -2347 9585 -2313 9619
rect -2279 9585 -2245 9619
rect -2211 9585 -2177 9619
rect -2143 9585 -2109 9619
rect -2075 9585 -2041 9619
rect -2007 9585 -1973 9619
rect -1939 9585 -1905 9619
rect -1871 9585 -1837 9619
rect -1803 9585 -1769 9619
rect -1735 9585 -1701 9619
rect -1667 9585 -1633 9619
rect -1599 9585 -1565 9619
rect -1531 9585 -1497 9619
rect -1463 9585 -1429 9619
rect -1395 9585 -1361 9619
rect -1327 9585 -1293 9619
rect -1259 9585 -1225 9619
rect -1191 9585 -1157 9619
rect -1123 9585 -1089 9619
rect -1055 9585 -1021 9619
rect -987 9585 -953 9619
rect -919 9585 -885 9619
rect -851 9585 -817 9619
rect -783 9585 -749 9619
rect -715 9585 -681 9619
rect -647 9585 -613 9619
rect -579 9585 -545 9619
rect -511 9585 -477 9619
rect -443 9585 -409 9619
rect -375 9585 -341 9619
rect -307 9585 -273 9619
rect -2959 9516 -2925 9550
rect -2891 9516 -2857 9550
rect -2823 9516 -2789 9550
rect -2755 9516 -2721 9550
rect -2687 9516 -2653 9550
rect -2619 9516 -2585 9550
rect -2551 9516 -2517 9550
rect -2483 9516 -2449 9550
rect -2415 9516 -2381 9550
rect -2347 9516 -2313 9550
rect -2279 9516 -2245 9550
rect -2211 9516 -2177 9550
rect -2143 9516 -2109 9550
rect -2075 9516 -2041 9550
rect -2007 9516 -1973 9550
rect -1939 9516 -1905 9550
rect -1871 9516 -1837 9550
rect -1803 9516 -1769 9550
rect -1735 9516 -1701 9550
rect -1667 9516 -1633 9550
rect -1599 9516 -1565 9550
rect -1531 9516 -1497 9550
rect -1463 9516 -1429 9550
rect -1395 9516 -1361 9550
rect -1327 9516 -1293 9550
rect -1259 9516 -1225 9550
rect -1191 9516 -1157 9550
rect -1123 9516 -1089 9550
rect -1055 9516 -1021 9550
rect -987 9516 -953 9550
rect -919 9516 -885 9550
rect -851 9516 -817 9550
rect -783 9516 -749 9550
rect -715 9516 -681 9550
rect -647 9516 -613 9550
rect -579 9516 -545 9550
rect -511 9516 -477 9550
rect -443 9516 -409 9550
rect -375 9516 -341 9550
rect -307 9516 -273 9550
rect -2959 9447 -2925 9481
rect -2891 9447 -2857 9481
rect -2823 9447 -2789 9481
rect -2755 9447 -2721 9481
rect -2687 9447 -2653 9481
rect -2619 9447 -2585 9481
rect -2551 9447 -2517 9481
rect -2483 9447 -2449 9481
rect -2415 9447 -2381 9481
rect -2347 9447 -2313 9481
rect -2279 9447 -2245 9481
rect -2211 9447 -2177 9481
rect -2143 9447 -2109 9481
rect -2075 9447 -2041 9481
rect -2007 9447 -1973 9481
rect -1939 9447 -1905 9481
rect -1871 9447 -1837 9481
rect -1803 9447 -1769 9481
rect -1735 9447 -1701 9481
rect -1667 9447 -1633 9481
rect -1599 9447 -1565 9481
rect -1531 9447 -1497 9481
rect -1463 9447 -1429 9481
rect -1395 9447 -1361 9481
rect -1327 9447 -1293 9481
rect -1259 9447 -1225 9481
rect -1191 9447 -1157 9481
rect -1123 9447 -1089 9481
rect -1055 9447 -1021 9481
rect -987 9447 -953 9481
rect -919 9447 -885 9481
rect -851 9447 -817 9481
rect -783 9447 -749 9481
rect -715 9447 -681 9481
rect -647 9447 -613 9481
rect -579 9447 -545 9481
rect -511 9447 -477 9481
rect -443 9447 -409 9481
rect -375 9447 -341 9481
rect -307 9447 -273 9481
rect -2959 9378 -2925 9412
rect -2891 9378 -2857 9412
rect -2823 9378 -2789 9412
rect -2755 9378 -2721 9412
rect -2687 9378 -2653 9412
rect -2619 9378 -2585 9412
rect -2551 9378 -2517 9412
rect -2483 9378 -2449 9412
rect -2415 9378 -2381 9412
rect -2347 9378 -2313 9412
rect -2279 9378 -2245 9412
rect -2211 9378 -2177 9412
rect -2143 9378 -2109 9412
rect -2075 9378 -2041 9412
rect -2007 9378 -1973 9412
rect -1939 9378 -1905 9412
rect -1871 9378 -1837 9412
rect -1803 9378 -1769 9412
rect -1735 9378 -1701 9412
rect -1667 9378 -1633 9412
rect -1599 9378 -1565 9412
rect -1531 9378 -1497 9412
rect -1463 9378 -1429 9412
rect -1395 9378 -1361 9412
rect -1327 9378 -1293 9412
rect -1259 9378 -1225 9412
rect -1191 9378 -1157 9412
rect -1123 9378 -1089 9412
rect -1055 9378 -1021 9412
rect -987 9378 -953 9412
rect -919 9378 -885 9412
rect -851 9378 -817 9412
rect -783 9378 -749 9412
rect -715 9378 -681 9412
rect -647 9378 -613 9412
rect -579 9378 -545 9412
rect -511 9378 -477 9412
rect -443 9378 -409 9412
rect -375 9378 -341 9412
rect -307 9378 -273 9412
rect -2959 9309 -2925 9343
rect -2891 9309 -2857 9343
rect -2823 9309 -2789 9343
rect -2755 9309 -2721 9343
rect -2687 9309 -2653 9343
rect -2619 9309 -2585 9343
rect -2551 9309 -2517 9343
rect -2483 9309 -2449 9343
rect -2415 9309 -2381 9343
rect -2347 9309 -2313 9343
rect -2279 9309 -2245 9343
rect -2211 9309 -2177 9343
rect -2143 9309 -2109 9343
rect -2075 9309 -2041 9343
rect -2007 9309 -1973 9343
rect -1939 9309 -1905 9343
rect -1871 9309 -1837 9343
rect -1803 9309 -1769 9343
rect -1735 9309 -1701 9343
rect -1667 9309 -1633 9343
rect -1599 9309 -1565 9343
rect -1531 9309 -1497 9343
rect -1463 9309 -1429 9343
rect -1395 9309 -1361 9343
rect -1327 9309 -1293 9343
rect -1259 9309 -1225 9343
rect -1191 9309 -1157 9343
rect -1123 9309 -1089 9343
rect -1055 9309 -1021 9343
rect -987 9309 -953 9343
rect -919 9309 -885 9343
rect -851 9309 -817 9343
rect -783 9309 -749 9343
rect -715 9309 -681 9343
rect -647 9309 -613 9343
rect -579 9309 -545 9343
rect -511 9309 -477 9343
rect -443 9309 -409 9343
rect -375 9309 -341 9343
rect -307 9309 -273 9343
rect -2959 9240 -2925 9274
rect -2891 9240 -2857 9274
rect -2823 9240 -2789 9274
rect -2755 9240 -2721 9274
rect -2687 9240 -2653 9274
rect -2619 9240 -2585 9274
rect -2551 9240 -2517 9274
rect -2483 9240 -2449 9274
rect -2415 9240 -2381 9274
rect -2347 9240 -2313 9274
rect -2279 9240 -2245 9274
rect -2211 9240 -2177 9274
rect -2143 9240 -2109 9274
rect -2075 9240 -2041 9274
rect -2007 9240 -1973 9274
rect -1939 9240 -1905 9274
rect -1871 9240 -1837 9274
rect -1803 9240 -1769 9274
rect -1735 9240 -1701 9274
rect -1667 9240 -1633 9274
rect -1599 9240 -1565 9274
rect -1531 9240 -1497 9274
rect -1463 9240 -1429 9274
rect -1395 9240 -1361 9274
rect -1327 9240 -1293 9274
rect -1259 9240 -1225 9274
rect -1191 9240 -1157 9274
rect -1123 9240 -1089 9274
rect -1055 9240 -1021 9274
rect -987 9240 -953 9274
rect -919 9240 -885 9274
rect -851 9240 -817 9274
rect -783 9240 -749 9274
rect -715 9240 -681 9274
rect -647 9240 -613 9274
rect -579 9240 -545 9274
rect -511 9240 -477 9274
rect -443 9240 -409 9274
rect -375 9240 -341 9274
rect -307 9240 -273 9274
rect -2959 9171 -2925 9205
rect -2891 9171 -2857 9205
rect -2823 9171 -2789 9205
rect -2755 9171 -2721 9205
rect -2687 9171 -2653 9205
rect -2619 9171 -2585 9205
rect -2551 9171 -2517 9205
rect -2483 9171 -2449 9205
rect -2415 9171 -2381 9205
rect -2347 9171 -2313 9205
rect -2279 9171 -2245 9205
rect -2211 9171 -2177 9205
rect -2143 9171 -2109 9205
rect -2075 9171 -2041 9205
rect -2007 9171 -1973 9205
rect -1939 9171 -1905 9205
rect -1871 9171 -1837 9205
rect -1803 9171 -1769 9205
rect -1735 9171 -1701 9205
rect -1667 9171 -1633 9205
rect -1599 9171 -1565 9205
rect -1531 9171 -1497 9205
rect -1463 9171 -1429 9205
rect -1395 9171 -1361 9205
rect -1327 9171 -1293 9205
rect -1259 9171 -1225 9205
rect -1191 9171 -1157 9205
rect -1123 9171 -1089 9205
rect -1055 9171 -1021 9205
rect -987 9171 -953 9205
rect -919 9171 -885 9205
rect -851 9171 -817 9205
rect -783 9171 -749 9205
rect -715 9171 -681 9205
rect -647 9171 -613 9205
rect -579 9171 -545 9205
rect -511 9171 -477 9205
rect -443 9171 -409 9205
rect -375 9171 -341 9205
rect -307 9171 -273 9205
rect -2959 9102 -2925 9136
rect -2891 9102 -2857 9136
rect -2823 9102 -2789 9136
rect -2755 9102 -2721 9136
rect -2687 9102 -2653 9136
rect -2619 9102 -2585 9136
rect -2551 9102 -2517 9136
rect -2483 9102 -2449 9136
rect -2415 9102 -2381 9136
rect -2347 9102 -2313 9136
rect -2279 9102 -2245 9136
rect -2211 9102 -2177 9136
rect -2143 9102 -2109 9136
rect -2075 9102 -2041 9136
rect -2007 9102 -1973 9136
rect -1939 9102 -1905 9136
rect -1871 9102 -1837 9136
rect -1803 9102 -1769 9136
rect -1735 9102 -1701 9136
rect -1667 9102 -1633 9136
rect -1599 9102 -1565 9136
rect -1531 9102 -1497 9136
rect -1463 9102 -1429 9136
rect -1395 9102 -1361 9136
rect -1327 9102 -1293 9136
rect -1259 9102 -1225 9136
rect -1191 9102 -1157 9136
rect -1123 9102 -1089 9136
rect -1055 9102 -1021 9136
rect -987 9102 -953 9136
rect -919 9102 -885 9136
rect -851 9102 -817 9136
rect -783 9102 -749 9136
rect -715 9102 -681 9136
rect -647 9102 -613 9136
rect -579 9102 -545 9136
rect -511 9102 -477 9136
rect -443 9102 -409 9136
rect -375 9102 -341 9136
rect -307 9102 -273 9136
rect -2959 9033 -2925 9067
rect -2891 9033 -2857 9067
rect -2823 9033 -2789 9067
rect -2755 9033 -2721 9067
rect -2687 9033 -2653 9067
rect -2619 9033 -2585 9067
rect -2551 9033 -2517 9067
rect -2483 9033 -2449 9067
rect -2415 9033 -2381 9067
rect -2347 9033 -2313 9067
rect -2279 9033 -2245 9067
rect -2211 9033 -2177 9067
rect -2143 9033 -2109 9067
rect -2075 9033 -2041 9067
rect -2007 9033 -1973 9067
rect -1939 9033 -1905 9067
rect -1871 9033 -1837 9067
rect -1803 9033 -1769 9067
rect -1735 9033 -1701 9067
rect -1667 9033 -1633 9067
rect -1599 9033 -1565 9067
rect -1531 9033 -1497 9067
rect -1463 9033 -1429 9067
rect -1395 9033 -1361 9067
rect -1327 9033 -1293 9067
rect -1259 9033 -1225 9067
rect -1191 9033 -1157 9067
rect -1123 9033 -1089 9067
rect -1055 9033 -1021 9067
rect -987 9033 -953 9067
rect -919 9033 -885 9067
rect -851 9033 -817 9067
rect -783 9033 -749 9067
rect -715 9033 -681 9067
rect -647 9033 -613 9067
rect -579 9033 -545 9067
rect -511 9033 -477 9067
rect -443 9033 -409 9067
rect -375 9033 -341 9067
rect -307 9033 -273 9067
rect -2959 8964 -2925 8998
rect -2891 8964 -2857 8998
rect -2823 8964 -2789 8998
rect -2755 8964 -2721 8998
rect -2687 8964 -2653 8998
rect -2619 8964 -2585 8998
rect -2551 8964 -2517 8998
rect -2483 8964 -2449 8998
rect -2415 8964 -2381 8998
rect -2347 8964 -2313 8998
rect -2279 8964 -2245 8998
rect -2211 8964 -2177 8998
rect -2143 8964 -2109 8998
rect -2075 8964 -2041 8998
rect -2007 8964 -1973 8998
rect -1939 8964 -1905 8998
rect -1871 8964 -1837 8998
rect -1803 8964 -1769 8998
rect -1735 8964 -1701 8998
rect -1667 8964 -1633 8998
rect -1599 8964 -1565 8998
rect -1531 8964 -1497 8998
rect -1463 8964 -1429 8998
rect -1395 8964 -1361 8998
rect -1327 8964 -1293 8998
rect -1259 8964 -1225 8998
rect -1191 8964 -1157 8998
rect -1123 8964 -1089 8998
rect -1055 8964 -1021 8998
rect -987 8964 -953 8998
rect -919 8964 -885 8998
rect -851 8964 -817 8998
rect -783 8964 -749 8998
rect -715 8964 -681 8998
rect -647 8964 -613 8998
rect -579 8964 -545 8998
rect -511 8964 -477 8998
rect -443 8964 -409 8998
rect -375 8964 -341 8998
rect -307 8964 -273 8998
rect -2959 8895 -2925 8929
rect -2891 8895 -2857 8929
rect -2823 8895 -2789 8929
rect -2755 8895 -2721 8929
rect -2687 8895 -2653 8929
rect -2619 8895 -2585 8929
rect -2551 8895 -2517 8929
rect -2483 8895 -2449 8929
rect -2415 8895 -2381 8929
rect -2347 8895 -2313 8929
rect -2279 8895 -2245 8929
rect -2211 8895 -2177 8929
rect -2143 8895 -2109 8929
rect -2075 8895 -2041 8929
rect -2007 8895 -1973 8929
rect -1939 8895 -1905 8929
rect -1871 8895 -1837 8929
rect -1803 8895 -1769 8929
rect -1735 8895 -1701 8929
rect -1667 8895 -1633 8929
rect -1599 8895 -1565 8929
rect -1531 8895 -1497 8929
rect -1463 8895 -1429 8929
rect -1395 8895 -1361 8929
rect -1327 8895 -1293 8929
rect -1259 8895 -1225 8929
rect -1191 8895 -1157 8929
rect -1123 8895 -1089 8929
rect -1055 8895 -1021 8929
rect -987 8895 -953 8929
rect -919 8895 -885 8929
rect -851 8895 -817 8929
rect -783 8895 -749 8929
rect -715 8895 -681 8929
rect -647 8895 -613 8929
rect -579 8895 -545 8929
rect -511 8895 -477 8929
rect -443 8895 -409 8929
rect -375 8895 -341 8929
rect -307 8895 -273 8929
rect -2959 8826 -2925 8860
rect -2891 8826 -2857 8860
rect -2823 8826 -2789 8860
rect -2755 8826 -2721 8860
rect -2687 8826 -2653 8860
rect -2619 8826 -2585 8860
rect -2551 8826 -2517 8860
rect -2483 8826 -2449 8860
rect -2415 8826 -2381 8860
rect -2347 8826 -2313 8860
rect -2279 8826 -2245 8860
rect -2211 8826 -2177 8860
rect -2143 8826 -2109 8860
rect -2075 8826 -2041 8860
rect -2007 8826 -1973 8860
rect -1939 8826 -1905 8860
rect -1871 8826 -1837 8860
rect -1803 8826 -1769 8860
rect -1735 8826 -1701 8860
rect -1667 8826 -1633 8860
rect -1599 8826 -1565 8860
rect -1531 8826 -1497 8860
rect -1463 8826 -1429 8860
rect -1395 8826 -1361 8860
rect -1327 8826 -1293 8860
rect -1259 8826 -1225 8860
rect -1191 8826 -1157 8860
rect -1123 8826 -1089 8860
rect -1055 8826 -1021 8860
rect -987 8826 -953 8860
rect -919 8826 -885 8860
rect -851 8826 -817 8860
rect -783 8826 -749 8860
rect -715 8826 -681 8860
rect -647 8826 -613 8860
rect -579 8826 -545 8860
rect -511 8826 -477 8860
rect -443 8826 -409 8860
rect -375 8826 -341 8860
rect -307 8826 -273 8860
rect -2959 8757 -2925 8791
rect -2891 8757 -2857 8791
rect -2823 8757 -2789 8791
rect -2755 8757 -2721 8791
rect -2687 8757 -2653 8791
rect -2619 8757 -2585 8791
rect -2551 8757 -2517 8791
rect -2483 8757 -2449 8791
rect -2415 8757 -2381 8791
rect -2347 8757 -2313 8791
rect -2279 8757 -2245 8791
rect -2211 8757 -2177 8791
rect -2143 8757 -2109 8791
rect -2075 8757 -2041 8791
rect -2007 8757 -1973 8791
rect -1939 8757 -1905 8791
rect -1871 8757 -1837 8791
rect -1803 8757 -1769 8791
rect -1735 8757 -1701 8791
rect -1667 8757 -1633 8791
rect -1599 8757 -1565 8791
rect -1531 8757 -1497 8791
rect -1463 8757 -1429 8791
rect -1395 8757 -1361 8791
rect -1327 8757 -1293 8791
rect -1259 8757 -1225 8791
rect -1191 8757 -1157 8791
rect -1123 8757 -1089 8791
rect -1055 8757 -1021 8791
rect -987 8757 -953 8791
rect -919 8757 -885 8791
rect -851 8757 -817 8791
rect -783 8757 -749 8791
rect -715 8757 -681 8791
rect -647 8757 -613 8791
rect -579 8757 -545 8791
rect -511 8757 -477 8791
rect -443 8757 -409 8791
rect -375 8757 -341 8791
rect -307 8757 -273 8791
rect -2959 8688 -2925 8722
rect -2891 8688 -2857 8722
rect -2823 8688 -2789 8722
rect -2755 8688 -2721 8722
rect -2687 8688 -2653 8722
rect -2619 8688 -2585 8722
rect -2551 8688 -2517 8722
rect -2483 8688 -2449 8722
rect -2415 8688 -2381 8722
rect -2347 8688 -2313 8722
rect -2279 8688 -2245 8722
rect -2211 8688 -2177 8722
rect -2143 8688 -2109 8722
rect -2075 8688 -2041 8722
rect -2007 8688 -1973 8722
rect -1939 8688 -1905 8722
rect -1871 8688 -1837 8722
rect -1803 8688 -1769 8722
rect -1735 8688 -1701 8722
rect -1667 8688 -1633 8722
rect -1599 8688 -1565 8722
rect -1531 8688 -1497 8722
rect -1463 8688 -1429 8722
rect -1395 8688 -1361 8722
rect -1327 8688 -1293 8722
rect -1259 8688 -1225 8722
rect -1191 8688 -1157 8722
rect -1123 8688 -1089 8722
rect -1055 8688 -1021 8722
rect -987 8688 -953 8722
rect -919 8688 -885 8722
rect -851 8688 -817 8722
rect -783 8688 -749 8722
rect -715 8688 -681 8722
rect -647 8688 -613 8722
rect -579 8688 -545 8722
rect -511 8688 -477 8722
rect -443 8688 -409 8722
rect -375 8688 -341 8722
rect -307 8688 -273 8722
rect -2959 8619 -2925 8653
rect -2891 8619 -2857 8653
rect -2823 8619 -2789 8653
rect -2755 8619 -2721 8653
rect -2687 8619 -2653 8653
rect -2619 8619 -2585 8653
rect -2551 8619 -2517 8653
rect -2483 8619 -2449 8653
rect -2415 8619 -2381 8653
rect -2347 8619 -2313 8653
rect -2279 8619 -2245 8653
rect -2211 8619 -2177 8653
rect -2143 8619 -2109 8653
rect -2075 8619 -2041 8653
rect -2007 8619 -1973 8653
rect -1939 8619 -1905 8653
rect -1871 8619 -1837 8653
rect -1803 8619 -1769 8653
rect -1735 8619 -1701 8653
rect -1667 8619 -1633 8653
rect -1599 8619 -1565 8653
rect -1531 8619 -1497 8653
rect -1463 8619 -1429 8653
rect -1395 8619 -1361 8653
rect -1327 8619 -1293 8653
rect -1259 8619 -1225 8653
rect -1191 8619 -1157 8653
rect -1123 8619 -1089 8653
rect -1055 8619 -1021 8653
rect -987 8619 -953 8653
rect -919 8619 -885 8653
rect -851 8619 -817 8653
rect -783 8619 -749 8653
rect -715 8619 -681 8653
rect -647 8619 -613 8653
rect -579 8619 -545 8653
rect -511 8619 -477 8653
rect -443 8619 -409 8653
rect -375 8619 -341 8653
rect -307 8619 -273 8653
rect -2959 8550 -2925 8584
rect -2891 8550 -2857 8584
rect -2823 8550 -2789 8584
rect -2755 8550 -2721 8584
rect -2687 8550 -2653 8584
rect -2619 8550 -2585 8584
rect -2551 8550 -2517 8584
rect -2483 8550 -2449 8584
rect -2415 8550 -2381 8584
rect -2347 8550 -2313 8584
rect -2279 8550 -2245 8584
rect -2211 8550 -2177 8584
rect -2143 8550 -2109 8584
rect -2075 8550 -2041 8584
rect -2007 8550 -1973 8584
rect -1939 8550 -1905 8584
rect -1871 8550 -1837 8584
rect -1803 8550 -1769 8584
rect -1735 8550 -1701 8584
rect -1667 8550 -1633 8584
rect -1599 8550 -1565 8584
rect -1531 8550 -1497 8584
rect -1463 8550 -1429 8584
rect -1395 8550 -1361 8584
rect -1327 8550 -1293 8584
rect -1259 8550 -1225 8584
rect -1191 8550 -1157 8584
rect -1123 8550 -1089 8584
rect -1055 8550 -1021 8584
rect -987 8550 -953 8584
rect -919 8550 -885 8584
rect -851 8550 -817 8584
rect -783 8550 -749 8584
rect -715 8550 -681 8584
rect -647 8550 -613 8584
rect -579 8550 -545 8584
rect -511 8550 -477 8584
rect -443 8550 -409 8584
rect -375 8550 -341 8584
rect -307 8550 -273 8584
rect -2959 8481 -2925 8515
rect -2891 8481 -2857 8515
rect -2823 8481 -2789 8515
rect -2755 8481 -2721 8515
rect -2687 8481 -2653 8515
rect -2619 8481 -2585 8515
rect -2551 8481 -2517 8515
rect -2483 8481 -2449 8515
rect -2415 8481 -2381 8515
rect -2347 8481 -2313 8515
rect -2279 8481 -2245 8515
rect -2211 8481 -2177 8515
rect -2143 8481 -2109 8515
rect -2075 8481 -2041 8515
rect -2007 8481 -1973 8515
rect -1939 8481 -1905 8515
rect -1871 8481 -1837 8515
rect -1803 8481 -1769 8515
rect -1735 8481 -1701 8515
rect -1667 8481 -1633 8515
rect -1599 8481 -1565 8515
rect -1531 8481 -1497 8515
rect -1463 8481 -1429 8515
rect -1395 8481 -1361 8515
rect -1327 8481 -1293 8515
rect -1259 8481 -1225 8515
rect -1191 8481 -1157 8515
rect -1123 8481 -1089 8515
rect -1055 8481 -1021 8515
rect -987 8481 -953 8515
rect -919 8481 -885 8515
rect -851 8481 -817 8515
rect -783 8481 -749 8515
rect -715 8481 -681 8515
rect -647 8481 -613 8515
rect -579 8481 -545 8515
rect -511 8481 -477 8515
rect -443 8481 -409 8515
rect -375 8481 -341 8515
rect -307 8481 -273 8515
rect -2959 8412 -2925 8446
rect -2891 8412 -2857 8446
rect -2823 8412 -2789 8446
rect -2755 8412 -2721 8446
rect -2687 8412 -2653 8446
rect -2619 8412 -2585 8446
rect -2551 8412 -2517 8446
rect -2483 8412 -2449 8446
rect -2415 8412 -2381 8446
rect -2347 8412 -2313 8446
rect -2279 8412 -2245 8446
rect -2211 8412 -2177 8446
rect -2143 8412 -2109 8446
rect -2075 8412 -2041 8446
rect -2007 8412 -1973 8446
rect -1939 8412 -1905 8446
rect -1871 8412 -1837 8446
rect -1803 8412 -1769 8446
rect -1735 8412 -1701 8446
rect -1667 8412 -1633 8446
rect -1599 8412 -1565 8446
rect -1531 8412 -1497 8446
rect -1463 8412 -1429 8446
rect -1395 8412 -1361 8446
rect -1327 8412 -1293 8446
rect -1259 8412 -1225 8446
rect -1191 8412 -1157 8446
rect -1123 8412 -1089 8446
rect -1055 8412 -1021 8446
rect -987 8412 -953 8446
rect -919 8412 -885 8446
rect -851 8412 -817 8446
rect -783 8412 -749 8446
rect -715 8412 -681 8446
rect -647 8412 -613 8446
rect -579 8412 -545 8446
rect -511 8412 -477 8446
rect -443 8412 -409 8446
rect -375 8412 -341 8446
rect -307 8412 -273 8446
rect -2959 8343 -2925 8377
rect -2891 8343 -2857 8377
rect -2823 8343 -2789 8377
rect -2755 8343 -2721 8377
rect -2687 8343 -2653 8377
rect -2619 8343 -2585 8377
rect -2551 8343 -2517 8377
rect -2483 8343 -2449 8377
rect -2415 8343 -2381 8377
rect -2347 8343 -2313 8377
rect -2279 8343 -2245 8377
rect -2211 8343 -2177 8377
rect -2143 8343 -2109 8377
rect -2075 8343 -2041 8377
rect -2007 8343 -1973 8377
rect -1939 8343 -1905 8377
rect -1871 8343 -1837 8377
rect -1803 8343 -1769 8377
rect -1735 8343 -1701 8377
rect -1667 8343 -1633 8377
rect -1599 8343 -1565 8377
rect -1531 8343 -1497 8377
rect -1463 8343 -1429 8377
rect -1395 8343 -1361 8377
rect -1327 8343 -1293 8377
rect -1259 8343 -1225 8377
rect -1191 8343 -1157 8377
rect -1123 8343 -1089 8377
rect -1055 8343 -1021 8377
rect -987 8343 -953 8377
rect -919 8343 -885 8377
rect -851 8343 -817 8377
rect -783 8343 -749 8377
rect -715 8343 -681 8377
rect -647 8343 -613 8377
rect -579 8343 -545 8377
rect -511 8343 -477 8377
rect -443 8343 -409 8377
rect -375 8343 -341 8377
rect -307 8343 -273 8377
rect -2959 8274 -2925 8308
rect -2891 8274 -2857 8308
rect -2823 8274 -2789 8308
rect -2755 8274 -2721 8308
rect -2687 8274 -2653 8308
rect -2619 8274 -2585 8308
rect -2551 8274 -2517 8308
rect -2483 8274 -2449 8308
rect -2415 8274 -2381 8308
rect -2347 8274 -2313 8308
rect -2279 8274 -2245 8308
rect -2211 8274 -2177 8308
rect -2143 8274 -2109 8308
rect -2075 8274 -2041 8308
rect -2007 8274 -1973 8308
rect -1939 8274 -1905 8308
rect -1871 8274 -1837 8308
rect -1803 8274 -1769 8308
rect -1735 8274 -1701 8308
rect -1667 8274 -1633 8308
rect -1599 8274 -1565 8308
rect -1531 8274 -1497 8308
rect -1463 8274 -1429 8308
rect -1395 8274 -1361 8308
rect -1327 8274 -1293 8308
rect -1259 8274 -1225 8308
rect -1191 8274 -1157 8308
rect -1123 8274 -1089 8308
rect -1055 8274 -1021 8308
rect -987 8274 -953 8308
rect -919 8274 -885 8308
rect -851 8274 -817 8308
rect -783 8274 -749 8308
rect -715 8274 -681 8308
rect -647 8274 -613 8308
rect -579 8274 -545 8308
rect -511 8274 -477 8308
rect -443 8274 -409 8308
rect -375 8274 -341 8308
rect -307 8274 -273 8308
rect -2959 8205 -2925 8239
rect -2891 8205 -2857 8239
rect -2823 8205 -2789 8239
rect -2755 8205 -2721 8239
rect -2687 8205 -2653 8239
rect -2619 8205 -2585 8239
rect -2551 8205 -2517 8239
rect -2483 8205 -2449 8239
rect -2415 8205 -2381 8239
rect -2347 8205 -2313 8239
rect -2279 8205 -2245 8239
rect -2211 8205 -2177 8239
rect -2143 8205 -2109 8239
rect -2075 8205 -2041 8239
rect -2007 8205 -1973 8239
rect -1939 8205 -1905 8239
rect -1871 8205 -1837 8239
rect -1803 8205 -1769 8239
rect -1735 8205 -1701 8239
rect -1667 8205 -1633 8239
rect -1599 8205 -1565 8239
rect -1531 8205 -1497 8239
rect -1463 8205 -1429 8239
rect -1395 8205 -1361 8239
rect -1327 8205 -1293 8239
rect -1259 8205 -1225 8239
rect -1191 8205 -1157 8239
rect -1123 8205 -1089 8239
rect -1055 8205 -1021 8239
rect -987 8205 -953 8239
rect -919 8205 -885 8239
rect -851 8205 -817 8239
rect -783 8205 -749 8239
rect -715 8205 -681 8239
rect -647 8205 -613 8239
rect -579 8205 -545 8239
rect -511 8205 -477 8239
rect -443 8205 -409 8239
rect -375 8205 -341 8239
rect -307 8205 -273 8239
rect -2959 8136 -2925 8170
rect -2891 8136 -2857 8170
rect -2823 8136 -2789 8170
rect -2755 8136 -2721 8170
rect -2687 8136 -2653 8170
rect -2619 8136 -2585 8170
rect -2551 8136 -2517 8170
rect -2483 8136 -2449 8170
rect -2415 8136 -2381 8170
rect -2347 8136 -2313 8170
rect -2279 8136 -2245 8170
rect -2211 8136 -2177 8170
rect -2143 8136 -2109 8170
rect -2075 8136 -2041 8170
rect -2007 8136 -1973 8170
rect -1939 8136 -1905 8170
rect -1871 8136 -1837 8170
rect -1803 8136 -1769 8170
rect -1735 8136 -1701 8170
rect -1667 8136 -1633 8170
rect -1599 8136 -1565 8170
rect -1531 8136 -1497 8170
rect -1463 8136 -1429 8170
rect -1395 8136 -1361 8170
rect -1327 8136 -1293 8170
rect -1259 8136 -1225 8170
rect -1191 8136 -1157 8170
rect -1123 8136 -1089 8170
rect -1055 8136 -1021 8170
rect -987 8136 -953 8170
rect -919 8136 -885 8170
rect -851 8136 -817 8170
rect -783 8136 -749 8170
rect -715 8136 -681 8170
rect -647 8136 -613 8170
rect -579 8136 -545 8170
rect -511 8136 -477 8170
rect -443 8136 -409 8170
rect -375 8136 -341 8170
rect -307 8136 -273 8170
rect -2959 8067 -2925 8101
rect -2891 8067 -2857 8101
rect -2823 8067 -2789 8101
rect -2755 8067 -2721 8101
rect -2687 8067 -2653 8101
rect -2619 8067 -2585 8101
rect -2551 8067 -2517 8101
rect -2483 8067 -2449 8101
rect -2415 8067 -2381 8101
rect -2347 8067 -2313 8101
rect -2279 8067 -2245 8101
rect -2211 8067 -2177 8101
rect -2143 8067 -2109 8101
rect -2075 8067 -2041 8101
rect -2007 8067 -1973 8101
rect -1939 8067 -1905 8101
rect -1871 8067 -1837 8101
rect -1803 8067 -1769 8101
rect -1735 8067 -1701 8101
rect -1667 8067 -1633 8101
rect -1599 8067 -1565 8101
rect -1531 8067 -1497 8101
rect -1463 8067 -1429 8101
rect -1395 8067 -1361 8101
rect -1327 8067 -1293 8101
rect -1259 8067 -1225 8101
rect -1191 8067 -1157 8101
rect -1123 8067 -1089 8101
rect -1055 8067 -1021 8101
rect -987 8067 -953 8101
rect -919 8067 -885 8101
rect -851 8067 -817 8101
rect -783 8067 -749 8101
rect -715 8067 -681 8101
rect -647 8067 -613 8101
rect -579 8067 -545 8101
rect -511 8067 -477 8101
rect -443 8067 -409 8101
rect -375 8067 -341 8101
rect -307 8067 -273 8101
rect -2959 7998 -2925 8032
rect -2891 7998 -2857 8032
rect -2823 7998 -2789 8032
rect -2755 7998 -2721 8032
rect -2687 7998 -2653 8032
rect -2619 7998 -2585 8032
rect -2551 7998 -2517 8032
rect -2483 7998 -2449 8032
rect -2415 7998 -2381 8032
rect -2347 7998 -2313 8032
rect -2279 7998 -2245 8032
rect -2211 7998 -2177 8032
rect -2143 7998 -2109 8032
rect -2075 7998 -2041 8032
rect -2007 7998 -1973 8032
rect -1939 7998 -1905 8032
rect -1871 7998 -1837 8032
rect -1803 7998 -1769 8032
rect -1735 7998 -1701 8032
rect -1667 7998 -1633 8032
rect -1599 7998 -1565 8032
rect -1531 7998 -1497 8032
rect -1463 7998 -1429 8032
rect -1395 7998 -1361 8032
rect -1327 7998 -1293 8032
rect -1259 7998 -1225 8032
rect -1191 7998 -1157 8032
rect -1123 7998 -1089 8032
rect -1055 7998 -1021 8032
rect -987 7998 -953 8032
rect -919 7998 -885 8032
rect -851 7998 -817 8032
rect -783 7998 -749 8032
rect -715 7998 -681 8032
rect -647 7998 -613 8032
rect -579 7998 -545 8032
rect -511 7998 -477 8032
rect -443 7998 -409 8032
rect -375 7998 -341 8032
rect -307 7998 -273 8032
rect -2959 7929 -2925 7963
rect -2891 7929 -2857 7963
rect -2823 7929 -2789 7963
rect -2755 7929 -2721 7963
rect -2687 7929 -2653 7963
rect -2619 7929 -2585 7963
rect -2551 7929 -2517 7963
rect -2483 7929 -2449 7963
rect -2415 7929 -2381 7963
rect -2347 7929 -2313 7963
rect -2279 7929 -2245 7963
rect -2211 7929 -2177 7963
rect -2143 7929 -2109 7963
rect -2075 7929 -2041 7963
rect -2007 7929 -1973 7963
rect -1939 7929 -1905 7963
rect -1871 7929 -1837 7963
rect -1803 7929 -1769 7963
rect -1735 7929 -1701 7963
rect -1667 7929 -1633 7963
rect -1599 7929 -1565 7963
rect -1531 7929 -1497 7963
rect -1463 7929 -1429 7963
rect -1395 7929 -1361 7963
rect -1327 7929 -1293 7963
rect -1259 7929 -1225 7963
rect -1191 7929 -1157 7963
rect -1123 7929 -1089 7963
rect -1055 7929 -1021 7963
rect -987 7929 -953 7963
rect -919 7929 -885 7963
rect -851 7929 -817 7963
rect -783 7929 -749 7963
rect -715 7929 -681 7963
rect -647 7929 -613 7963
rect -579 7929 -545 7963
rect -511 7929 -477 7963
rect -443 7929 -409 7963
rect -375 7929 -341 7963
rect -307 7929 -273 7963
rect -2959 7860 -2925 7894
rect -2891 7860 -2857 7894
rect -2823 7860 -2789 7894
rect -2755 7860 -2721 7894
rect -2687 7860 -2653 7894
rect -2619 7860 -2585 7894
rect -2551 7860 -2517 7894
rect -2483 7860 -2449 7894
rect -2415 7860 -2381 7894
rect -2347 7860 -2313 7894
rect -2279 7860 -2245 7894
rect -2211 7860 -2177 7894
rect -2143 7860 -2109 7894
rect -2075 7860 -2041 7894
rect -2007 7860 -1973 7894
rect -1939 7860 -1905 7894
rect -1871 7860 -1837 7894
rect -1803 7860 -1769 7894
rect -1735 7860 -1701 7894
rect -1667 7860 -1633 7894
rect -1599 7860 -1565 7894
rect -1531 7860 -1497 7894
rect -1463 7860 -1429 7894
rect -1395 7860 -1361 7894
rect -1327 7860 -1293 7894
rect -1259 7860 -1225 7894
rect -1191 7860 -1157 7894
rect -1123 7860 -1089 7894
rect -1055 7860 -1021 7894
rect -987 7860 -953 7894
rect -919 7860 -885 7894
rect -851 7860 -817 7894
rect -783 7860 -749 7894
rect -715 7860 -681 7894
rect -647 7860 -613 7894
rect -579 7860 -545 7894
rect -511 7860 -477 7894
rect -443 7860 -409 7894
rect -375 7860 -341 7894
rect -307 7860 -273 7894
rect -2959 7791 -2925 7825
rect -2891 7791 -2857 7825
rect -2823 7791 -2789 7825
rect -2755 7791 -2721 7825
rect -2687 7791 -2653 7825
rect -2619 7791 -2585 7825
rect -2551 7791 -2517 7825
rect -2483 7791 -2449 7825
rect -2415 7791 -2381 7825
rect -2347 7791 -2313 7825
rect -2279 7791 -2245 7825
rect -2211 7791 -2177 7825
rect -2143 7791 -2109 7825
rect -2075 7791 -2041 7825
rect -2007 7791 -1973 7825
rect -1939 7791 -1905 7825
rect -1871 7791 -1837 7825
rect -1803 7791 -1769 7825
rect -1735 7791 -1701 7825
rect -1667 7791 -1633 7825
rect -1599 7791 -1565 7825
rect -1531 7791 -1497 7825
rect -1463 7791 -1429 7825
rect -1395 7791 -1361 7825
rect -1327 7791 -1293 7825
rect -1259 7791 -1225 7825
rect -1191 7791 -1157 7825
rect -1123 7791 -1089 7825
rect -1055 7791 -1021 7825
rect -987 7791 -953 7825
rect -919 7791 -885 7825
rect -851 7791 -817 7825
rect -783 7791 -749 7825
rect -715 7791 -681 7825
rect -647 7791 -613 7825
rect -579 7791 -545 7825
rect -511 7791 -477 7825
rect -443 7791 -409 7825
rect -375 7791 -341 7825
rect -307 7791 -273 7825
rect -2959 7722 -2925 7756
rect -2891 7722 -2857 7756
rect -2823 7722 -2789 7756
rect -2755 7722 -2721 7756
rect -2687 7722 -2653 7756
rect -2619 7722 -2585 7756
rect -2551 7722 -2517 7756
rect -2483 7722 -2449 7756
rect -2415 7722 -2381 7756
rect -2347 7722 -2313 7756
rect -2279 7722 -2245 7756
rect -2211 7722 -2177 7756
rect -2143 7722 -2109 7756
rect -2075 7722 -2041 7756
rect -2007 7722 -1973 7756
rect -1939 7722 -1905 7756
rect -1871 7722 -1837 7756
rect -1803 7722 -1769 7756
rect -1735 7722 -1701 7756
rect -1667 7722 -1633 7756
rect -1599 7722 -1565 7756
rect -1531 7722 -1497 7756
rect -1463 7722 -1429 7756
rect -1395 7722 -1361 7756
rect -1327 7722 -1293 7756
rect -1259 7722 -1225 7756
rect -1191 7722 -1157 7756
rect -1123 7722 -1089 7756
rect -1055 7722 -1021 7756
rect -987 7722 -953 7756
rect -919 7722 -885 7756
rect -851 7722 -817 7756
rect -783 7722 -749 7756
rect -715 7722 -681 7756
rect -647 7722 -613 7756
rect -579 7722 -545 7756
rect -511 7722 -477 7756
rect -443 7722 -409 7756
rect -375 7722 -341 7756
rect -307 7722 -273 7756
rect -2959 7653 -2925 7687
rect -2891 7653 -2857 7687
rect -2823 7653 -2789 7687
rect -2755 7653 -2721 7687
rect -2687 7653 -2653 7687
rect -2619 7653 -2585 7687
rect -2551 7653 -2517 7687
rect -2483 7653 -2449 7687
rect -2415 7653 -2381 7687
rect -2347 7653 -2313 7687
rect -2279 7653 -2245 7687
rect -2211 7653 -2177 7687
rect -2143 7653 -2109 7687
rect -2075 7653 -2041 7687
rect -2007 7653 -1973 7687
rect -1939 7653 -1905 7687
rect -1871 7653 -1837 7687
rect -1803 7653 -1769 7687
rect -1735 7653 -1701 7687
rect -1667 7653 -1633 7687
rect -1599 7653 -1565 7687
rect -1531 7653 -1497 7687
rect -1463 7653 -1429 7687
rect -1395 7653 -1361 7687
rect -1327 7653 -1293 7687
rect -1259 7653 -1225 7687
rect -1191 7653 -1157 7687
rect -1123 7653 -1089 7687
rect -1055 7653 -1021 7687
rect -987 7653 -953 7687
rect -919 7653 -885 7687
rect -851 7653 -817 7687
rect -783 7653 -749 7687
rect -715 7653 -681 7687
rect -647 7653 -613 7687
rect -579 7653 -545 7687
rect -511 7653 -477 7687
rect -443 7653 -409 7687
rect -375 7653 -341 7687
rect -307 7653 -273 7687
rect -2959 7584 -2925 7618
rect -2891 7584 -2857 7618
rect -2823 7584 -2789 7618
rect -2755 7584 -2721 7618
rect -2687 7584 -2653 7618
rect -2619 7584 -2585 7618
rect -2551 7584 -2517 7618
rect -2483 7584 -2449 7618
rect -2415 7584 -2381 7618
rect -2347 7584 -2313 7618
rect -2279 7584 -2245 7618
rect -2211 7584 -2177 7618
rect -2143 7584 -2109 7618
rect -2075 7584 -2041 7618
rect -2007 7584 -1973 7618
rect -1939 7584 -1905 7618
rect -1871 7584 -1837 7618
rect -1803 7584 -1769 7618
rect -1735 7584 -1701 7618
rect -1667 7584 -1633 7618
rect -1599 7584 -1565 7618
rect -1531 7584 -1497 7618
rect -1463 7584 -1429 7618
rect -1395 7584 -1361 7618
rect -1327 7584 -1293 7618
rect -1259 7584 -1225 7618
rect -1191 7584 -1157 7618
rect -1123 7584 -1089 7618
rect -1055 7584 -1021 7618
rect -987 7584 -953 7618
rect -919 7584 -885 7618
rect -851 7584 -817 7618
rect -783 7584 -749 7618
rect -715 7584 -681 7618
rect -647 7584 -613 7618
rect -579 7584 -545 7618
rect -511 7584 -477 7618
rect -443 7584 -409 7618
rect -375 7584 -341 7618
rect -307 7584 -273 7618
rect -2959 7515 -2925 7549
rect -2891 7515 -2857 7549
rect -2823 7515 -2789 7549
rect -2755 7515 -2721 7549
rect -2687 7515 -2653 7549
rect -2619 7515 -2585 7549
rect -2551 7515 -2517 7549
rect -2483 7515 -2449 7549
rect -2415 7515 -2381 7549
rect -2347 7515 -2313 7549
rect -2279 7515 -2245 7549
rect -2211 7515 -2177 7549
rect -2143 7515 -2109 7549
rect -2075 7515 -2041 7549
rect -2007 7515 -1973 7549
rect -1939 7515 -1905 7549
rect -1871 7515 -1837 7549
rect -1803 7515 -1769 7549
rect -1735 7515 -1701 7549
rect -1667 7515 -1633 7549
rect -1599 7515 -1565 7549
rect -1531 7515 -1497 7549
rect -1463 7515 -1429 7549
rect -1395 7515 -1361 7549
rect -1327 7515 -1293 7549
rect -1259 7515 -1225 7549
rect -1191 7515 -1157 7549
rect -1123 7515 -1089 7549
rect -1055 7515 -1021 7549
rect -987 7515 -953 7549
rect -919 7515 -885 7549
rect -851 7515 -817 7549
rect -783 7515 -749 7549
rect -715 7515 -681 7549
rect -647 7515 -613 7549
rect -579 7515 -545 7549
rect -511 7515 -477 7549
rect -443 7515 -409 7549
rect -375 7515 -341 7549
rect -307 7515 -273 7549
rect -2959 7446 -2925 7480
rect -2891 7446 -2857 7480
rect -2823 7446 -2789 7480
rect -2755 7446 -2721 7480
rect -2687 7446 -2653 7480
rect -2619 7446 -2585 7480
rect -2551 7446 -2517 7480
rect -2483 7446 -2449 7480
rect -2415 7446 -2381 7480
rect -2347 7446 -2313 7480
rect -2279 7446 -2245 7480
rect -2211 7446 -2177 7480
rect -2143 7446 -2109 7480
rect -2075 7446 -2041 7480
rect -2007 7446 -1973 7480
rect -1939 7446 -1905 7480
rect -1871 7446 -1837 7480
rect -1803 7446 -1769 7480
rect -1735 7446 -1701 7480
rect -1667 7446 -1633 7480
rect -1599 7446 -1565 7480
rect -1531 7446 -1497 7480
rect -1463 7446 -1429 7480
rect -1395 7446 -1361 7480
rect -1327 7446 -1293 7480
rect -1259 7446 -1225 7480
rect -1191 7446 -1157 7480
rect -1123 7446 -1089 7480
rect -1055 7446 -1021 7480
rect -987 7446 -953 7480
rect -919 7446 -885 7480
rect -851 7446 -817 7480
rect -783 7446 -749 7480
rect -715 7446 -681 7480
rect -647 7446 -613 7480
rect -579 7446 -545 7480
rect -511 7446 -477 7480
rect -443 7446 -409 7480
rect -375 7446 -341 7480
rect -307 7446 -273 7480
<< mvnsubdiffcont >>
rect 15 50602 49 50636
rect 87 50598 121 50632
rect 159 50593 193 50627
rect 15 50534 49 50568
rect 87 50530 121 50564
rect 159 50525 193 50559
rect 15 50466 49 50500
rect 87 50462 121 50496
rect 159 50457 193 50491
rect 15 50398 49 50432
rect 87 50394 121 50428
rect 159 50389 193 50423
rect 15 50330 49 50364
rect 87 50326 121 50360
rect 159 50321 193 50355
rect 15 50262 49 50296
rect 87 50258 121 50292
rect 159 50253 193 50287
rect 15 50194 49 50228
rect 87 50190 121 50224
rect 159 50185 193 50219
rect 15 50126 49 50160
rect 87 50122 121 50156
rect 159 50117 193 50151
rect 15 50058 49 50092
rect 87 50054 121 50088
rect 159 50049 193 50083
rect 15 49990 49 50024
rect 87 49986 121 50020
rect 159 49981 193 50015
rect 15 49922 49 49956
rect 87 49918 121 49952
rect 159 49913 193 49947
rect 15 49854 49 49888
rect 87 49850 121 49884
rect 159 49845 193 49879
rect 15 49786 49 49820
rect 87 49782 121 49816
rect 159 49777 193 49811
rect 15 49718 49 49752
rect 87 49714 121 49748
rect 159 49709 193 49743
rect 15 49650 49 49684
rect 87 49646 121 49680
rect 159 49641 193 49675
rect 15 49582 49 49616
rect 87 49578 121 49612
rect 159 49573 193 49607
rect 15 49514 49 49548
rect 87 49510 121 49544
rect 159 49505 193 49539
rect 15 49446 49 49480
rect 87 49442 121 49476
rect 159 49437 193 49471
rect 15 49378 49 49412
rect 87 49374 121 49408
rect 159 49369 193 49403
rect 15 49310 49 49344
rect 87 49306 121 49340
rect 159 49301 193 49335
rect 15 49242 49 49276
rect 87 49238 121 49272
rect 159 49233 193 49267
rect 15 49174 49 49208
rect 87 49170 121 49204
rect 159 49165 193 49199
rect 15 49106 49 49140
rect 87 49102 121 49136
rect 159 49097 193 49131
rect 15 49038 49 49072
rect 87 49034 121 49068
rect 159 49029 193 49063
rect 15 48970 49 49004
rect 87 48966 121 49000
rect 159 48961 193 48995
rect 15 48902 49 48936
rect 87 48898 121 48932
rect 159 48893 193 48927
rect 15 48834 49 48868
rect 87 48830 121 48864
rect 159 48825 193 48859
rect 15 48766 49 48800
rect 87 48762 121 48796
rect 159 48757 193 48791
rect 15 48698 49 48732
rect 87 48694 121 48728
rect 159 48689 193 48723
rect 15 48630 49 48664
rect 87 48626 121 48660
rect 159 48621 193 48655
rect 15 48562 49 48596
rect 87 48558 121 48592
rect 159 48553 193 48587
rect 15 48494 49 48528
rect 87 48490 121 48524
rect 159 48485 193 48519
rect 15 48426 49 48460
rect 87 48422 121 48456
rect 159 48417 193 48451
rect 15 48358 49 48392
rect 87 48354 121 48388
rect 159 48349 193 48383
rect 15 48290 49 48324
rect 87 48286 121 48320
rect 159 48281 193 48315
rect 15 48222 49 48256
rect 87 48218 121 48252
rect 159 48213 193 48247
rect 15 48154 49 48188
rect 87 48150 121 48184
rect 159 48145 193 48179
rect 15 48086 49 48120
rect 87 48082 121 48116
rect 159 48077 193 48111
rect 15 48018 49 48052
rect 87 48014 121 48048
rect 159 48009 193 48043
rect 15 47950 49 47984
rect 87 47946 121 47980
rect 159 47941 193 47975
rect 15 47882 49 47916
rect 87 47878 121 47912
rect 159 47873 193 47907
rect 15 47814 49 47848
rect 87 47810 121 47844
rect 159 47805 193 47839
rect 15 47746 49 47780
rect 87 47742 121 47776
rect 159 47737 193 47771
rect 15 47678 49 47712
rect 87 47674 121 47708
rect 159 47669 193 47703
rect 15 47610 49 47644
rect 87 47606 121 47640
rect 159 47601 193 47635
rect 15 47542 49 47576
rect 87 47538 121 47572
rect 159 47533 193 47567
rect 15 47474 49 47508
rect 87 47470 121 47504
rect 159 47465 193 47499
rect 15 47406 49 47440
rect 87 47402 121 47436
rect 159 47397 193 47431
rect 15 47338 49 47372
rect 87 47334 121 47368
rect 159 47329 193 47363
rect 15 47270 49 47304
rect 87 47266 121 47300
rect 159 47261 193 47295
rect 15 47202 49 47236
rect 87 47198 121 47232
rect 159 47193 193 47227
rect 15 47134 49 47168
rect 87 47130 121 47164
rect 159 47125 193 47159
rect 15 47066 49 47100
rect 87 47062 121 47096
rect 159 47057 193 47091
rect 15 46998 49 47032
rect 87 46994 121 47028
rect 159 46989 193 47023
rect 15 46930 49 46964
rect 87 46926 121 46960
rect 159 46921 193 46955
rect 15 46862 49 46896
rect 87 46858 121 46892
rect 159 46853 193 46887
rect 15 46794 49 46828
rect 87 46790 121 46824
rect 159 46785 193 46819
rect 15 46726 49 46760
rect 87 46722 121 46756
rect 159 46717 193 46751
rect 15 46658 49 46692
rect 87 46654 121 46688
rect 159 46649 193 46683
rect 15 46590 49 46624
rect 87 46586 121 46620
rect 159 46581 193 46615
rect 15 46522 49 46556
rect 87 46518 121 46552
rect 159 46513 193 46547
rect 15 46454 49 46488
rect 87 46450 121 46484
rect 159 46445 193 46479
rect 15 46386 49 46420
rect 87 46382 121 46416
rect 159 46377 193 46411
rect 15 46318 49 46352
rect 87 46314 121 46348
rect 159 46309 193 46343
rect 15 46250 49 46284
rect 87 46246 121 46280
rect 159 46241 193 46275
rect 15 46182 49 46216
rect 87 46178 121 46212
rect 159 46173 193 46207
rect 15 46114 49 46148
rect 87 46110 121 46144
rect 159 46105 193 46139
rect 15 46046 49 46080
rect 87 46042 121 46076
rect 159 46037 193 46071
rect 15 45978 49 46012
rect 87 45974 121 46008
rect 159 45969 193 46003
rect 15 45910 49 45944
rect 87 45906 121 45940
rect 159 45901 193 45935
rect 15 45842 49 45876
rect 87 45838 121 45872
rect 159 45833 193 45867
rect 15 45774 49 45808
rect 87 45770 121 45804
rect 159 45765 193 45799
rect 15 45706 49 45740
rect 87 45702 121 45736
rect 159 45697 193 45731
rect 15 45638 49 45672
rect 87 45634 121 45668
rect 159 45629 193 45663
rect 15 45570 49 45604
rect 87 45566 121 45600
rect 159 45561 193 45595
rect 15 45502 49 45536
rect 87 45498 121 45532
rect 159 45493 193 45527
rect 15 45434 49 45468
rect 87 45430 121 45464
rect 159 45425 193 45459
rect 15 45366 49 45400
rect 87 45362 121 45396
rect 159 45357 193 45391
rect 15 45298 49 45332
rect 87 45294 121 45328
rect 159 45289 193 45323
rect 15 45230 49 45264
rect 87 45226 121 45260
rect 159 45221 193 45255
rect 15 45162 49 45196
rect 87 45158 121 45192
rect 159 45153 193 45187
rect 15 45094 49 45128
rect 87 45090 121 45124
rect 159 45085 193 45119
rect 15 45026 49 45060
rect 87 45022 121 45056
rect 159 45017 193 45051
rect 15 44958 49 44992
rect 87 44954 121 44988
rect 159 44949 193 44983
rect 15 44890 49 44924
rect 87 44886 121 44920
rect 159 44881 193 44915
rect 15 44822 49 44856
rect 87 44818 121 44852
rect 159 44813 193 44847
rect 15 44754 49 44788
rect 87 44750 121 44784
rect 159 44745 193 44779
rect 15 44686 49 44720
rect 87 44682 121 44716
rect 159 44677 193 44711
rect 15 44618 49 44652
rect 87 44614 121 44648
rect 159 44609 193 44643
rect 15 44550 49 44584
rect 87 44546 121 44580
rect 159 44541 193 44575
rect 15 44482 49 44516
rect 87 44478 121 44512
rect 159 44473 193 44507
rect 15 44414 49 44448
rect 87 44410 121 44444
rect 159 44405 193 44439
rect 15 44346 49 44380
rect 87 44342 121 44376
rect 159 44337 193 44371
rect 15 44278 49 44312
rect 87 44274 121 44308
rect 159 44269 193 44303
rect 15 44210 49 44244
rect 87 44206 121 44240
rect 159 44201 193 44235
rect 15 44142 49 44176
rect 87 44138 121 44172
rect 159 44133 193 44167
rect 15 44074 49 44108
rect 87 44070 121 44104
rect 159 44065 193 44099
rect 15 44006 49 44040
rect 87 44002 121 44036
rect 159 43997 193 44031
rect 15 43938 49 43972
rect 87 43934 121 43968
rect 159 43929 193 43963
rect 15 43870 49 43904
rect 87 43866 121 43900
rect 159 43861 193 43895
rect 15 43802 49 43836
rect 87 43798 121 43832
rect 159 43793 193 43827
rect 15 43734 49 43768
rect 87 43730 121 43764
rect 159 43725 193 43759
rect 15 43666 49 43700
rect 87 43662 121 43696
rect 159 43657 193 43691
rect 15 43598 49 43632
rect 87 43594 121 43628
rect 159 43589 193 43623
rect 15 43530 49 43564
rect 87 43526 121 43560
rect 159 43521 193 43555
rect 15 43462 49 43496
rect 87 43458 121 43492
rect 159 43453 193 43487
rect 15 43394 49 43428
rect 87 43390 121 43424
rect 159 43385 193 43419
rect 15 43326 49 43360
rect 87 43322 121 43356
rect 159 43317 193 43351
rect 15 43258 49 43292
rect 87 43254 121 43288
rect 159 43249 193 43283
rect 15 43190 49 43224
rect 87 43186 121 43220
rect 159 43181 193 43215
rect 15 43122 49 43156
rect 87 43118 121 43152
rect 159 43113 193 43147
rect 15 43054 49 43088
rect 87 43050 121 43084
rect 159 43045 193 43079
rect 15 42986 49 43020
rect 87 42982 121 43016
rect 159 42977 193 43011
rect 15 42918 49 42952
rect 87 42914 121 42948
rect 159 42909 193 42943
rect 15 42850 49 42884
rect 87 42846 121 42880
rect 159 42841 193 42875
rect 15 42782 49 42816
rect 87 42778 121 42812
rect 159 42773 193 42807
rect 15 42714 49 42748
rect 87 42710 121 42744
rect 159 42705 193 42739
rect 15 42646 49 42680
rect 87 42642 121 42676
rect 159 42637 193 42671
rect 15 42578 49 42612
rect 87 42574 121 42608
rect 159 42569 193 42603
rect 15 42510 49 42544
rect 87 42506 121 42540
rect 159 42501 193 42535
rect 15 42442 49 42476
rect 87 42438 121 42472
rect 159 42433 193 42467
rect 15 42374 49 42408
rect 87 42370 121 42404
rect 159 42365 193 42399
rect 15 42306 49 42340
rect 87 42302 121 42336
rect 159 42297 193 42331
rect 15 42238 49 42272
rect 87 42234 121 42268
rect 159 42229 193 42263
rect 15 42170 49 42204
rect 87 42166 121 42200
rect 159 42161 193 42195
rect 15 42102 49 42136
rect 87 42098 121 42132
rect 159 42093 193 42127
rect 15 42034 49 42068
rect 87 42030 121 42064
rect 159 42025 193 42059
rect 15 41966 49 42000
rect 87 41962 121 41996
rect 159 41957 193 41991
rect 15 41898 49 41932
rect 87 41894 121 41928
rect 159 41889 193 41923
rect 15 41830 49 41864
rect 87 41826 121 41860
rect 159 41821 193 41855
rect 15 41762 49 41796
rect 87 41758 121 41792
rect 159 41753 193 41787
rect 15 41694 49 41728
rect 87 41690 121 41724
rect 159 41685 193 41719
rect 15 41626 49 41660
rect 87 41622 121 41656
rect 159 41617 193 41651
rect 15 41558 49 41592
rect 87 41554 121 41588
rect 159 41549 193 41583
rect 15 41490 49 41524
rect 87 41486 121 41520
rect 159 41481 193 41515
rect 15 41422 49 41456
rect 87 41418 121 41452
rect 159 41413 193 41447
rect 15 41354 49 41388
rect 87 41350 121 41384
rect 159 41345 193 41379
rect 15 41286 49 41320
rect 87 41282 121 41316
rect 159 41277 193 41311
rect 15 41218 49 41252
rect 87 41214 121 41248
rect 159 41209 193 41243
rect 15 41150 49 41184
rect 87 41146 121 41180
rect 159 41141 193 41175
rect 15 41082 49 41116
rect 87 41078 121 41112
rect 159 41073 193 41107
rect 15 41014 49 41048
rect 87 41010 121 41044
rect 159 41005 193 41039
rect 15 40946 49 40980
rect 87 40942 121 40976
rect 159 40937 193 40971
rect 15 40878 49 40912
rect 87 40874 121 40908
rect 159 40869 193 40903
rect 15 40810 49 40844
rect 87 40806 121 40840
rect 159 40801 193 40835
rect 15 40742 49 40776
rect 87 40738 121 40772
rect 159 40733 193 40767
rect 15 40674 49 40708
rect 87 40670 121 40704
rect 159 40665 193 40699
rect 15 40606 49 40640
rect 87 40602 121 40636
rect 159 40597 193 40631
rect 15 40538 49 40572
rect 87 40534 121 40568
rect 159 40529 193 40563
rect 15 40470 49 40504
rect 87 40466 121 40500
rect 159 40461 193 40495
rect 15 40402 49 40436
rect 87 40398 121 40432
rect 159 40393 193 40427
rect 15 40334 49 40368
rect 87 40330 121 40364
rect 159 40325 193 40359
rect 15 40266 49 40300
rect 87 40262 121 40296
rect 159 40257 193 40291
rect 15 40198 49 40232
rect 87 40194 121 40228
rect 159 40189 193 40223
rect 15 40130 49 40164
rect 87 40126 121 40160
rect 159 40121 193 40155
rect 15 40062 49 40096
rect 87 40058 121 40092
rect 159 40053 193 40087
rect 15 39994 49 40028
rect 87 39990 121 40024
rect 159 39985 193 40019
rect 15 39926 49 39960
rect 87 39922 121 39956
rect 159 39917 193 39951
rect 15 39858 49 39892
rect 87 39854 121 39888
rect 159 39849 193 39883
rect 15 39790 49 39824
rect 87 39786 121 39820
rect 159 39781 193 39815
rect 15 39722 49 39756
rect 87 39718 121 39752
rect 159 39713 193 39747
rect 15 39654 49 39688
rect 87 39650 121 39684
rect 159 39645 193 39679
rect 15 39586 49 39620
rect 87 39582 121 39616
rect 159 39577 193 39611
rect 15 39518 49 39552
rect 87 39514 121 39548
rect 159 39509 193 39543
rect 15 39450 49 39484
rect 87 39446 121 39480
rect 159 39441 193 39475
rect 15 39382 49 39416
rect 87 39378 121 39412
rect 159 39373 193 39407
rect 15 39314 49 39348
rect 87 39310 121 39344
rect 159 39305 193 39339
rect 15 39246 49 39280
rect 87 39242 121 39276
rect 159 39237 193 39271
rect 15 39178 49 39212
rect 87 39174 121 39208
rect 159 39169 193 39203
rect 15 39110 49 39144
rect 87 39106 121 39140
rect 159 39101 193 39135
rect 15 39042 49 39076
rect 87 39038 121 39072
rect 159 39033 193 39067
rect 15 38974 49 39008
rect 87 38970 121 39004
rect 159 38965 193 38999
rect 15 38906 49 38940
rect 87 38902 121 38936
rect 159 38897 193 38931
rect 15 38838 49 38872
rect 87 38834 121 38868
rect 159 38829 193 38863
rect 15 38770 49 38804
rect 87 38766 121 38800
rect 159 38761 193 38795
rect 15 38702 49 38736
rect 87 38698 121 38732
rect 159 38693 193 38727
rect 15 38634 49 38668
rect 87 38630 121 38664
rect 159 38625 193 38659
rect 15 38566 49 38600
rect 87 38562 121 38596
rect 159 38557 193 38591
rect 15 38498 49 38532
rect 87 38494 121 38528
rect 159 38489 193 38523
rect 15 38430 49 38464
rect 87 38426 121 38460
rect 159 38421 193 38455
rect 15 38362 49 38396
rect 87 38358 121 38392
rect 159 38353 193 38387
rect 15 38294 49 38328
rect 87 38290 121 38324
rect 159 38285 193 38319
rect 15 38226 49 38260
rect 87 38222 121 38256
rect 159 38217 193 38251
rect 15 38158 49 38192
rect 87 38154 121 38188
rect 159 38149 193 38183
rect 15 38090 49 38124
rect 87 38086 121 38120
rect 159 38081 193 38115
rect 15 38022 49 38056
rect 87 38018 121 38052
rect 159 38013 193 38047
rect 15 37954 49 37988
rect 87 37950 121 37984
rect 159 37945 193 37979
rect 15 37886 49 37920
rect 87 37882 121 37916
rect 159 37877 193 37911
rect 15 37818 49 37852
rect 87 37814 121 37848
rect 159 37809 193 37843
rect 15 37750 49 37784
rect 87 37746 121 37780
rect 159 37741 193 37775
rect 15 37682 49 37716
rect 87 37678 121 37712
rect 159 37673 193 37707
rect 15 37614 49 37648
rect 87 37610 121 37644
rect 159 37605 193 37639
rect 15 37546 49 37580
rect 87 37542 121 37576
rect 159 37537 193 37571
rect 15 37478 49 37512
rect 87 37474 121 37508
rect 159 37469 193 37503
rect 15 37410 49 37444
rect 87 37406 121 37440
rect 159 37401 193 37435
rect 15 37342 49 37376
rect 87 37338 121 37372
rect 159 37333 193 37367
rect 15 37274 49 37308
rect 87 37270 121 37304
rect 159 37265 193 37299
rect 15 37206 49 37240
rect 87 37202 121 37236
rect 159 37197 193 37231
rect 15 37138 49 37172
rect 87 37134 121 37168
rect 159 37129 193 37163
rect 15 37070 49 37104
rect 87 37066 121 37100
rect 159 37061 193 37095
rect 15 37002 49 37036
rect 87 36998 121 37032
rect 159 36993 193 37027
rect 15 36934 49 36968
rect 87 36930 121 36964
rect 159 36925 193 36959
rect 15 36866 49 36900
rect 87 36862 121 36896
rect 159 36857 193 36891
rect 15 36798 49 36832
rect 87 36794 121 36828
rect 159 36789 193 36823
rect 15 36730 49 36764
rect 87 36726 121 36760
rect 159 36721 193 36755
rect 15 36662 49 36696
rect 87 36658 121 36692
rect 159 36653 193 36687
rect 15 36594 49 36628
rect 87 36590 121 36624
rect 159 36585 193 36619
rect 15 36526 49 36560
rect 87 36522 121 36556
rect 159 36517 193 36551
rect 15 36458 49 36492
rect 87 36454 121 36488
rect 159 36449 193 36483
rect 15 36390 49 36424
rect 87 36386 121 36420
rect 159 36381 193 36415
rect 15 36322 49 36356
rect 87 36318 121 36352
rect 159 36313 193 36347
rect 15 36254 49 36288
rect 87 36250 121 36284
rect 159 36245 193 36279
rect 15 36186 49 36220
rect 87 36182 121 36216
rect 159 36177 193 36211
rect 15 36118 49 36152
rect 87 36114 121 36148
rect 159 36109 193 36143
rect 15 36050 49 36084
rect 87 36046 121 36080
rect 159 36041 193 36075
rect 15 35982 49 36016
rect 87 35978 121 36012
rect 159 35973 193 36007
rect 15 35914 49 35948
rect 87 35910 121 35944
rect 159 35905 193 35939
rect 15 35846 49 35880
rect 87 35842 121 35876
rect 159 35837 193 35871
rect 15 35778 49 35812
rect 87 35774 121 35808
rect 159 35769 193 35803
rect 15 35710 49 35744
rect 87 35706 121 35740
rect 159 35701 193 35735
rect 15 35642 49 35676
rect 87 35638 121 35672
rect 159 35633 193 35667
rect 15 35574 49 35608
rect 87 35570 121 35604
rect 159 35565 193 35599
rect 15 35506 49 35540
rect 87 35502 121 35536
rect 159 35497 193 35531
rect 15 35438 49 35472
rect 87 35434 121 35468
rect 159 35429 193 35463
rect 15 35370 49 35404
rect 87 35366 121 35400
rect 159 35361 193 35395
rect 15 35302 49 35336
rect 87 35298 121 35332
rect 159 35293 193 35327
rect 15 35234 49 35268
rect 87 35230 121 35264
rect 159 35225 193 35259
rect 15 35166 49 35200
rect 87 35162 121 35196
rect 159 35157 193 35191
rect 15 35098 49 35132
rect 87 35094 121 35128
rect 159 35089 193 35123
rect 15 35030 49 35064
rect 87 35026 121 35060
rect 159 35021 193 35055
rect 15 34962 49 34996
rect 87 34958 121 34992
rect 159 34953 193 34987
rect 15 34894 49 34928
rect 87 34890 121 34924
rect 159 34885 193 34919
rect -2833 34826 -2799 34860
rect -2765 34826 -2731 34860
rect -2697 34826 -2663 34860
rect -2629 34826 -2595 34860
rect -2561 34826 -2527 34860
rect -2493 34826 -2459 34860
rect -2425 34826 -2391 34860
rect -2357 34826 -2323 34860
rect -2289 34826 -2255 34860
rect -2221 34826 -2187 34860
rect -2153 34826 -2119 34860
rect -2085 34826 -2051 34860
rect -2017 34826 -1983 34860
rect -1949 34826 -1915 34860
rect -1881 34826 -1847 34860
rect -1813 34826 -1779 34860
rect -1745 34826 -1711 34860
rect -1677 34826 -1643 34860
rect -1609 34826 -1575 34860
rect -1541 34826 -1507 34860
rect -1473 34826 -1439 34860
rect -1405 34826 -1371 34860
rect -1337 34826 -1303 34860
rect -1269 34826 -1235 34860
rect -1201 34826 -1167 34860
rect -1133 34826 -1099 34860
rect -1065 34826 -1031 34860
rect -997 34826 -963 34860
rect -929 34826 -895 34860
rect -861 34826 -827 34860
rect -793 34826 -759 34860
rect -725 34826 -691 34860
rect -657 34826 -623 34860
rect -589 34826 -555 34860
rect -521 34826 -487 34860
rect -453 34826 -419 34860
rect -385 34826 -351 34860
rect -317 34826 -283 34860
rect -249 34826 -215 34860
rect -181 34826 -147 34860
rect -113 34826 -79 34860
rect 15 34826 49 34860
rect 87 34822 121 34856
rect 159 34817 193 34851
rect -2833 34754 -2799 34788
rect -2765 34754 -2731 34788
rect -2697 34754 -2663 34788
rect -2629 34754 -2595 34788
rect -2561 34754 -2527 34788
rect -2493 34754 -2459 34788
rect -2425 34754 -2391 34788
rect -2357 34754 -2323 34788
rect -2289 34754 -2255 34788
rect -2221 34754 -2187 34788
rect -2153 34754 -2119 34788
rect -2085 34754 -2051 34788
rect -2017 34754 -1983 34788
rect -1949 34754 -1915 34788
rect -1881 34754 -1847 34788
rect -1813 34754 -1779 34788
rect -1745 34754 -1711 34788
rect -1677 34754 -1643 34788
rect -1609 34754 -1575 34788
rect -1541 34754 -1507 34788
rect -1473 34754 -1439 34788
rect -1405 34754 -1371 34788
rect -1337 34754 -1303 34788
rect -1269 34754 -1235 34788
rect -1201 34754 -1167 34788
rect -1133 34754 -1099 34788
rect -1065 34754 -1031 34788
rect -997 34754 -963 34788
rect -929 34754 -895 34788
rect -861 34754 -827 34788
rect -793 34754 -759 34788
rect -725 34754 -691 34788
rect -657 34754 -623 34788
rect -589 34754 -555 34788
rect -521 34754 -487 34788
rect -453 34754 -419 34788
rect -385 34754 -351 34788
rect -317 34754 -283 34788
rect -249 34754 -215 34788
rect -181 34754 -147 34788
rect -113 34754 -79 34788
rect -45 34754 -11 34788
rect 87 34754 121 34788
rect 159 34749 193 34783
rect -2833 34682 -2799 34716
rect -2765 34682 -2731 34716
rect -2697 34682 -2663 34716
rect -2629 34682 -2595 34716
rect -2561 34682 -2527 34716
rect -2493 34682 -2459 34716
rect -2425 34682 -2391 34716
rect -2357 34682 -2323 34716
rect -2289 34682 -2255 34716
rect -2221 34682 -2187 34716
rect -2153 34682 -2119 34716
rect -2085 34682 -2051 34716
rect -2017 34682 -1983 34716
rect -1949 34682 -1915 34716
rect -1881 34682 -1847 34716
rect -1813 34682 -1779 34716
rect -1745 34682 -1711 34716
rect -1677 34682 -1643 34716
rect -1609 34682 -1575 34716
rect -1541 34682 -1507 34716
rect -1473 34682 -1439 34716
rect -1405 34682 -1371 34716
rect -1337 34682 -1303 34716
rect -1269 34682 -1235 34716
rect -1201 34682 -1167 34716
rect -1133 34682 -1099 34716
rect -1065 34682 -1031 34716
rect -997 34682 -963 34716
rect -929 34682 -895 34716
rect -861 34682 -827 34716
rect -793 34682 -759 34716
rect -725 34682 -691 34716
rect -657 34682 -623 34716
rect -589 34682 -555 34716
rect -521 34682 -487 34716
rect -453 34682 -419 34716
rect -385 34682 -351 34716
rect -317 34682 -283 34716
rect -249 34682 -215 34716
rect -181 34682 -147 34716
rect -113 34682 -79 34716
rect -45 34682 -11 34716
rect 23 34682 57 34716
rect 91 34682 125 34716
<< locali >>
rect -2969 50624 -153 50648
rect -2969 37942 -2938 50624
rect -184 37942 -153 50624
rect -2969 37907 -2829 37942
rect -275 37907 -153 37942
rect -2969 37873 -2938 37907
rect -2904 37873 -2870 37907
rect -2836 37901 -2829 37907
rect -2836 37873 -2802 37901
rect -2768 37873 -2734 37901
rect -2700 37873 -2666 37901
rect -2632 37873 -2598 37901
rect -2564 37873 -2530 37901
rect -2496 37873 -2462 37901
rect -2428 37873 -2394 37901
rect -2360 37873 -2326 37901
rect -2292 37873 -2258 37901
rect -2224 37873 -2190 37901
rect -2156 37873 -2122 37901
rect -2088 37873 -2054 37901
rect -2020 37873 -1986 37901
rect -1952 37873 -1918 37901
rect -1884 37873 -1850 37901
rect -1816 37873 -1782 37901
rect -1748 37873 -1714 37901
rect -1680 37873 -1646 37901
rect -1612 37873 -1578 37901
rect -1544 37873 -1510 37901
rect -1476 37873 -1442 37901
rect -1408 37873 -1374 37901
rect -1340 37873 -1306 37901
rect -1272 37873 -1238 37901
rect -1204 37873 -1170 37901
rect -1136 37873 -1102 37901
rect -1068 37873 -1034 37901
rect -1000 37873 -966 37901
rect -932 37873 -898 37901
rect -864 37873 -830 37901
rect -796 37873 -762 37901
rect -728 37873 -694 37901
rect -660 37873 -626 37901
rect -592 37873 -558 37901
rect -524 37873 -490 37901
rect -456 37873 -422 37901
rect -388 37873 -354 37901
rect -320 37873 -286 37901
rect -252 37873 -218 37907
rect -184 37873 -153 37907
rect -2969 37862 -153 37873
rect -2969 37838 -2829 37862
rect -2795 37838 -2757 37862
rect -2723 37838 -2685 37862
rect -2651 37838 -2613 37862
rect -2579 37838 -2541 37862
rect -2507 37838 -2469 37862
rect -2435 37838 -2397 37862
rect -2363 37838 -2325 37862
rect -2291 37838 -2253 37862
rect -2219 37838 -2181 37862
rect -2147 37838 -2109 37862
rect -2075 37838 -2037 37862
rect -2003 37838 -1965 37862
rect -1931 37838 -1893 37862
rect -1859 37838 -1821 37862
rect -1787 37838 -1749 37862
rect -1715 37838 -1677 37862
rect -1643 37838 -1605 37862
rect -1571 37838 -1533 37862
rect -1499 37838 -1461 37862
rect -1427 37838 -1389 37862
rect -1355 37838 -1317 37862
rect -1283 37838 -1245 37862
rect -1211 37838 -1173 37862
rect -1139 37838 -1101 37862
rect -1067 37838 -1029 37862
rect -995 37838 -957 37862
rect -923 37838 -885 37862
rect -851 37838 -813 37862
rect -779 37838 -741 37862
rect -707 37838 -669 37862
rect -635 37838 -597 37862
rect -563 37838 -525 37862
rect -491 37838 -453 37862
rect -419 37838 -381 37862
rect -347 37838 -309 37862
rect -275 37838 -153 37862
rect -2969 37804 -2938 37838
rect -2904 37804 -2870 37838
rect -2836 37828 -2829 37838
rect -2768 37828 -2757 37838
rect -2700 37828 -2685 37838
rect -2632 37828 -2613 37838
rect -2564 37828 -2541 37838
rect -2496 37828 -2469 37838
rect -2428 37828 -2397 37838
rect -2836 37804 -2802 37828
rect -2768 37804 -2734 37828
rect -2700 37804 -2666 37828
rect -2632 37804 -2598 37828
rect -2564 37804 -2530 37828
rect -2496 37804 -2462 37828
rect -2428 37804 -2394 37828
rect -2360 37804 -2326 37838
rect -2291 37828 -2258 37838
rect -2219 37828 -2190 37838
rect -2147 37828 -2122 37838
rect -2075 37828 -2054 37838
rect -2003 37828 -1986 37838
rect -1931 37828 -1918 37838
rect -1859 37828 -1850 37838
rect -1787 37828 -1782 37838
rect -1715 37828 -1714 37838
rect -2292 37804 -2258 37828
rect -2224 37804 -2190 37828
rect -2156 37804 -2122 37828
rect -2088 37804 -2054 37828
rect -2020 37804 -1986 37828
rect -1952 37804 -1918 37828
rect -1884 37804 -1850 37828
rect -1816 37804 -1782 37828
rect -1748 37804 -1714 37828
rect -1680 37828 -1677 37838
rect -1612 37828 -1605 37838
rect -1544 37828 -1533 37838
rect -1476 37828 -1461 37838
rect -1408 37828 -1389 37838
rect -1340 37828 -1317 37838
rect -1272 37828 -1245 37838
rect -1204 37828 -1173 37838
rect -1680 37804 -1646 37828
rect -1612 37804 -1578 37828
rect -1544 37804 -1510 37828
rect -1476 37804 -1442 37828
rect -1408 37804 -1374 37828
rect -1340 37804 -1306 37828
rect -1272 37804 -1238 37828
rect -1204 37804 -1170 37828
rect -1136 37804 -1102 37838
rect -1067 37828 -1034 37838
rect -995 37828 -966 37838
rect -923 37828 -898 37838
rect -851 37828 -830 37838
rect -779 37828 -762 37838
rect -707 37828 -694 37838
rect -635 37828 -626 37838
rect -563 37828 -558 37838
rect -491 37828 -490 37838
rect -1068 37804 -1034 37828
rect -1000 37804 -966 37828
rect -932 37804 -898 37828
rect -864 37804 -830 37828
rect -796 37804 -762 37828
rect -728 37804 -694 37828
rect -660 37804 -626 37828
rect -592 37804 -558 37828
rect -524 37804 -490 37828
rect -456 37828 -453 37838
rect -388 37828 -381 37838
rect -320 37828 -309 37838
rect -456 37804 -422 37828
rect -388 37804 -354 37828
rect -320 37804 -286 37828
rect -252 37804 -218 37838
rect -184 37804 -153 37838
rect -2969 37789 -153 37804
rect -2969 37769 -2829 37789
rect -2795 37769 -2757 37789
rect -2723 37769 -2685 37789
rect -2651 37769 -2613 37789
rect -2579 37769 -2541 37789
rect -2507 37769 -2469 37789
rect -2435 37769 -2397 37789
rect -2363 37769 -2325 37789
rect -2291 37769 -2253 37789
rect -2219 37769 -2181 37789
rect -2147 37769 -2109 37789
rect -2075 37769 -2037 37789
rect -2003 37769 -1965 37789
rect -1931 37769 -1893 37789
rect -1859 37769 -1821 37789
rect -1787 37769 -1749 37789
rect -1715 37769 -1677 37789
rect -1643 37769 -1605 37789
rect -1571 37769 -1533 37789
rect -1499 37769 -1461 37789
rect -1427 37769 -1389 37789
rect -1355 37769 -1317 37789
rect -1283 37769 -1245 37789
rect -1211 37769 -1173 37789
rect -1139 37769 -1101 37789
rect -1067 37769 -1029 37789
rect -995 37769 -957 37789
rect -923 37769 -885 37789
rect -851 37769 -813 37789
rect -779 37769 -741 37789
rect -707 37769 -669 37789
rect -635 37769 -597 37789
rect -563 37769 -525 37789
rect -491 37769 -453 37789
rect -419 37769 -381 37789
rect -347 37769 -309 37789
rect -275 37769 -153 37789
rect -2969 37735 -2938 37769
rect -2904 37735 -2870 37769
rect -2836 37755 -2829 37769
rect -2768 37755 -2757 37769
rect -2700 37755 -2685 37769
rect -2632 37755 -2613 37769
rect -2564 37755 -2541 37769
rect -2496 37755 -2469 37769
rect -2428 37755 -2397 37769
rect -2836 37735 -2802 37755
rect -2768 37735 -2734 37755
rect -2700 37735 -2666 37755
rect -2632 37735 -2598 37755
rect -2564 37735 -2530 37755
rect -2496 37735 -2462 37755
rect -2428 37735 -2394 37755
rect -2360 37735 -2326 37769
rect -2291 37755 -2258 37769
rect -2219 37755 -2190 37769
rect -2147 37755 -2122 37769
rect -2075 37755 -2054 37769
rect -2003 37755 -1986 37769
rect -1931 37755 -1918 37769
rect -1859 37755 -1850 37769
rect -1787 37755 -1782 37769
rect -1715 37755 -1714 37769
rect -2292 37735 -2258 37755
rect -2224 37735 -2190 37755
rect -2156 37735 -2122 37755
rect -2088 37735 -2054 37755
rect -2020 37735 -1986 37755
rect -1952 37735 -1918 37755
rect -1884 37735 -1850 37755
rect -1816 37735 -1782 37755
rect -1748 37735 -1714 37755
rect -1680 37755 -1677 37769
rect -1612 37755 -1605 37769
rect -1544 37755 -1533 37769
rect -1476 37755 -1461 37769
rect -1408 37755 -1389 37769
rect -1340 37755 -1317 37769
rect -1272 37755 -1245 37769
rect -1204 37755 -1173 37769
rect -1680 37735 -1646 37755
rect -1612 37735 -1578 37755
rect -1544 37735 -1510 37755
rect -1476 37735 -1442 37755
rect -1408 37735 -1374 37755
rect -1340 37735 -1306 37755
rect -1272 37735 -1238 37755
rect -1204 37735 -1170 37755
rect -1136 37735 -1102 37769
rect -1067 37755 -1034 37769
rect -995 37755 -966 37769
rect -923 37755 -898 37769
rect -851 37755 -830 37769
rect -779 37755 -762 37769
rect -707 37755 -694 37769
rect -635 37755 -626 37769
rect -563 37755 -558 37769
rect -491 37755 -490 37769
rect -1068 37735 -1034 37755
rect -1000 37735 -966 37755
rect -932 37735 -898 37755
rect -864 37735 -830 37755
rect -796 37735 -762 37755
rect -728 37735 -694 37755
rect -660 37735 -626 37755
rect -592 37735 -558 37755
rect -524 37735 -490 37755
rect -456 37755 -453 37769
rect -388 37755 -381 37769
rect -320 37755 -309 37769
rect -456 37735 -422 37755
rect -388 37735 -354 37755
rect -320 37735 -286 37755
rect -252 37735 -218 37769
rect -184 37735 -153 37769
rect -2969 37716 -153 37735
rect -2969 37700 -2829 37716
rect -2795 37700 -2757 37716
rect -2723 37700 -2685 37716
rect -2651 37700 -2613 37716
rect -2579 37700 -2541 37716
rect -2507 37700 -2469 37716
rect -2435 37700 -2397 37716
rect -2363 37700 -2325 37716
rect -2291 37700 -2253 37716
rect -2219 37700 -2181 37716
rect -2147 37700 -2109 37716
rect -2075 37700 -2037 37716
rect -2003 37700 -1965 37716
rect -1931 37700 -1893 37716
rect -1859 37700 -1821 37716
rect -1787 37700 -1749 37716
rect -1715 37700 -1677 37716
rect -1643 37700 -1605 37716
rect -1571 37700 -1533 37716
rect -1499 37700 -1461 37716
rect -1427 37700 -1389 37716
rect -1355 37700 -1317 37716
rect -1283 37700 -1245 37716
rect -1211 37700 -1173 37716
rect -1139 37700 -1101 37716
rect -1067 37700 -1029 37716
rect -995 37700 -957 37716
rect -923 37700 -885 37716
rect -851 37700 -813 37716
rect -779 37700 -741 37716
rect -707 37700 -669 37716
rect -635 37700 -597 37716
rect -563 37700 -525 37716
rect -491 37700 -453 37716
rect -419 37700 -381 37716
rect -347 37700 -309 37716
rect -275 37700 -153 37716
rect -2969 37666 -2938 37700
rect -2904 37666 -2870 37700
rect -2836 37682 -2829 37700
rect -2768 37682 -2757 37700
rect -2700 37682 -2685 37700
rect -2632 37682 -2613 37700
rect -2564 37682 -2541 37700
rect -2496 37682 -2469 37700
rect -2428 37682 -2397 37700
rect -2836 37666 -2802 37682
rect -2768 37666 -2734 37682
rect -2700 37666 -2666 37682
rect -2632 37666 -2598 37682
rect -2564 37666 -2530 37682
rect -2496 37666 -2462 37682
rect -2428 37666 -2394 37682
rect -2360 37666 -2326 37700
rect -2291 37682 -2258 37700
rect -2219 37682 -2190 37700
rect -2147 37682 -2122 37700
rect -2075 37682 -2054 37700
rect -2003 37682 -1986 37700
rect -1931 37682 -1918 37700
rect -1859 37682 -1850 37700
rect -1787 37682 -1782 37700
rect -1715 37682 -1714 37700
rect -2292 37666 -2258 37682
rect -2224 37666 -2190 37682
rect -2156 37666 -2122 37682
rect -2088 37666 -2054 37682
rect -2020 37666 -1986 37682
rect -1952 37666 -1918 37682
rect -1884 37666 -1850 37682
rect -1816 37666 -1782 37682
rect -1748 37666 -1714 37682
rect -1680 37682 -1677 37700
rect -1612 37682 -1605 37700
rect -1544 37682 -1533 37700
rect -1476 37682 -1461 37700
rect -1408 37682 -1389 37700
rect -1340 37682 -1317 37700
rect -1272 37682 -1245 37700
rect -1204 37682 -1173 37700
rect -1680 37666 -1646 37682
rect -1612 37666 -1578 37682
rect -1544 37666 -1510 37682
rect -1476 37666 -1442 37682
rect -1408 37666 -1374 37682
rect -1340 37666 -1306 37682
rect -1272 37666 -1238 37682
rect -1204 37666 -1170 37682
rect -1136 37666 -1102 37700
rect -1067 37682 -1034 37700
rect -995 37682 -966 37700
rect -923 37682 -898 37700
rect -851 37682 -830 37700
rect -779 37682 -762 37700
rect -707 37682 -694 37700
rect -635 37682 -626 37700
rect -563 37682 -558 37700
rect -491 37682 -490 37700
rect -1068 37666 -1034 37682
rect -1000 37666 -966 37682
rect -932 37666 -898 37682
rect -864 37666 -830 37682
rect -796 37666 -762 37682
rect -728 37666 -694 37682
rect -660 37666 -626 37682
rect -592 37666 -558 37682
rect -524 37666 -490 37682
rect -456 37682 -453 37700
rect -388 37682 -381 37700
rect -320 37682 -309 37700
rect -456 37666 -422 37682
rect -388 37666 -354 37682
rect -320 37666 -286 37682
rect -252 37666 -218 37700
rect -184 37666 -153 37700
rect -2969 37643 -153 37666
rect -2969 37631 -2829 37643
rect -2795 37631 -2757 37643
rect -2723 37631 -2685 37643
rect -2651 37631 -2613 37643
rect -2579 37631 -2541 37643
rect -2507 37631 -2469 37643
rect -2435 37631 -2397 37643
rect -2363 37631 -2325 37643
rect -2291 37631 -2253 37643
rect -2219 37631 -2181 37643
rect -2147 37631 -2109 37643
rect -2075 37631 -2037 37643
rect -2003 37631 -1965 37643
rect -1931 37631 -1893 37643
rect -1859 37631 -1821 37643
rect -1787 37631 -1749 37643
rect -1715 37631 -1677 37643
rect -1643 37631 -1605 37643
rect -1571 37631 -1533 37643
rect -1499 37631 -1461 37643
rect -1427 37631 -1389 37643
rect -1355 37631 -1317 37643
rect -1283 37631 -1245 37643
rect -1211 37631 -1173 37643
rect -1139 37631 -1101 37643
rect -1067 37631 -1029 37643
rect -995 37631 -957 37643
rect -923 37631 -885 37643
rect -851 37631 -813 37643
rect -779 37631 -741 37643
rect -707 37631 -669 37643
rect -635 37631 -597 37643
rect -563 37631 -525 37643
rect -491 37631 -453 37643
rect -419 37631 -381 37643
rect -347 37631 -309 37643
rect -275 37631 -153 37643
rect -2969 37597 -2938 37631
rect -2904 37597 -2870 37631
rect -2836 37609 -2829 37631
rect -2768 37609 -2757 37631
rect -2700 37609 -2685 37631
rect -2632 37609 -2613 37631
rect -2564 37609 -2541 37631
rect -2496 37609 -2469 37631
rect -2428 37609 -2397 37631
rect -2836 37597 -2802 37609
rect -2768 37597 -2734 37609
rect -2700 37597 -2666 37609
rect -2632 37597 -2598 37609
rect -2564 37597 -2530 37609
rect -2496 37597 -2462 37609
rect -2428 37597 -2394 37609
rect -2360 37597 -2326 37631
rect -2291 37609 -2258 37631
rect -2219 37609 -2190 37631
rect -2147 37609 -2122 37631
rect -2075 37609 -2054 37631
rect -2003 37609 -1986 37631
rect -1931 37609 -1918 37631
rect -1859 37609 -1850 37631
rect -1787 37609 -1782 37631
rect -1715 37609 -1714 37631
rect -2292 37597 -2258 37609
rect -2224 37597 -2190 37609
rect -2156 37597 -2122 37609
rect -2088 37597 -2054 37609
rect -2020 37597 -1986 37609
rect -1952 37597 -1918 37609
rect -1884 37597 -1850 37609
rect -1816 37597 -1782 37609
rect -1748 37597 -1714 37609
rect -1680 37609 -1677 37631
rect -1612 37609 -1605 37631
rect -1544 37609 -1533 37631
rect -1476 37609 -1461 37631
rect -1408 37609 -1389 37631
rect -1340 37609 -1317 37631
rect -1272 37609 -1245 37631
rect -1204 37609 -1173 37631
rect -1680 37597 -1646 37609
rect -1612 37597 -1578 37609
rect -1544 37597 -1510 37609
rect -1476 37597 -1442 37609
rect -1408 37597 -1374 37609
rect -1340 37597 -1306 37609
rect -1272 37597 -1238 37609
rect -1204 37597 -1170 37609
rect -1136 37597 -1102 37631
rect -1067 37609 -1034 37631
rect -995 37609 -966 37631
rect -923 37609 -898 37631
rect -851 37609 -830 37631
rect -779 37609 -762 37631
rect -707 37609 -694 37631
rect -635 37609 -626 37631
rect -563 37609 -558 37631
rect -491 37609 -490 37631
rect -1068 37597 -1034 37609
rect -1000 37597 -966 37609
rect -932 37597 -898 37609
rect -864 37597 -830 37609
rect -796 37597 -762 37609
rect -728 37597 -694 37609
rect -660 37597 -626 37609
rect -592 37597 -558 37609
rect -524 37597 -490 37609
rect -456 37609 -453 37631
rect -388 37609 -381 37631
rect -320 37609 -309 37631
rect -456 37597 -422 37609
rect -388 37597 -354 37609
rect -320 37597 -286 37609
rect -252 37597 -218 37631
rect -184 37597 -153 37631
rect -2969 37570 -153 37597
rect -2969 37562 -2829 37570
rect -2795 37562 -2757 37570
rect -2723 37562 -2685 37570
rect -2651 37562 -2613 37570
rect -2579 37562 -2541 37570
rect -2507 37562 -2469 37570
rect -2435 37562 -2397 37570
rect -2363 37562 -2325 37570
rect -2291 37562 -2253 37570
rect -2219 37562 -2181 37570
rect -2147 37562 -2109 37570
rect -2075 37562 -2037 37570
rect -2003 37562 -1965 37570
rect -1931 37562 -1893 37570
rect -1859 37562 -1821 37570
rect -1787 37562 -1749 37570
rect -1715 37562 -1677 37570
rect -1643 37562 -1605 37570
rect -1571 37562 -1533 37570
rect -1499 37562 -1461 37570
rect -1427 37562 -1389 37570
rect -1355 37562 -1317 37570
rect -1283 37562 -1245 37570
rect -1211 37562 -1173 37570
rect -1139 37562 -1101 37570
rect -1067 37562 -1029 37570
rect -995 37562 -957 37570
rect -923 37562 -885 37570
rect -851 37562 -813 37570
rect -779 37562 -741 37570
rect -707 37562 -669 37570
rect -635 37562 -597 37570
rect -563 37562 -525 37570
rect -491 37562 -453 37570
rect -419 37562 -381 37570
rect -347 37562 -309 37570
rect -275 37562 -153 37570
rect -2969 37528 -2938 37562
rect -2904 37528 -2870 37562
rect -2836 37536 -2829 37562
rect -2768 37536 -2757 37562
rect -2700 37536 -2685 37562
rect -2632 37536 -2613 37562
rect -2564 37536 -2541 37562
rect -2496 37536 -2469 37562
rect -2428 37536 -2397 37562
rect -2836 37528 -2802 37536
rect -2768 37528 -2734 37536
rect -2700 37528 -2666 37536
rect -2632 37528 -2598 37536
rect -2564 37528 -2530 37536
rect -2496 37528 -2462 37536
rect -2428 37528 -2394 37536
rect -2360 37528 -2326 37562
rect -2291 37536 -2258 37562
rect -2219 37536 -2190 37562
rect -2147 37536 -2122 37562
rect -2075 37536 -2054 37562
rect -2003 37536 -1986 37562
rect -1931 37536 -1918 37562
rect -1859 37536 -1850 37562
rect -1787 37536 -1782 37562
rect -1715 37536 -1714 37562
rect -2292 37528 -2258 37536
rect -2224 37528 -2190 37536
rect -2156 37528 -2122 37536
rect -2088 37528 -2054 37536
rect -2020 37528 -1986 37536
rect -1952 37528 -1918 37536
rect -1884 37528 -1850 37536
rect -1816 37528 -1782 37536
rect -1748 37528 -1714 37536
rect -1680 37536 -1677 37562
rect -1612 37536 -1605 37562
rect -1544 37536 -1533 37562
rect -1476 37536 -1461 37562
rect -1408 37536 -1389 37562
rect -1340 37536 -1317 37562
rect -1272 37536 -1245 37562
rect -1204 37536 -1173 37562
rect -1680 37528 -1646 37536
rect -1612 37528 -1578 37536
rect -1544 37528 -1510 37536
rect -1476 37528 -1442 37536
rect -1408 37528 -1374 37536
rect -1340 37528 -1306 37536
rect -1272 37528 -1238 37536
rect -1204 37528 -1170 37536
rect -1136 37528 -1102 37562
rect -1067 37536 -1034 37562
rect -995 37536 -966 37562
rect -923 37536 -898 37562
rect -851 37536 -830 37562
rect -779 37536 -762 37562
rect -707 37536 -694 37562
rect -635 37536 -626 37562
rect -563 37536 -558 37562
rect -491 37536 -490 37562
rect -1068 37528 -1034 37536
rect -1000 37528 -966 37536
rect -932 37528 -898 37536
rect -864 37528 -830 37536
rect -796 37528 -762 37536
rect -728 37528 -694 37536
rect -660 37528 -626 37536
rect -592 37528 -558 37536
rect -524 37528 -490 37536
rect -456 37536 -453 37562
rect -388 37536 -381 37562
rect -320 37536 -309 37562
rect -456 37528 -422 37536
rect -388 37528 -354 37536
rect -320 37528 -286 37536
rect -252 37528 -218 37562
rect -184 37528 -153 37562
rect -2969 37497 -153 37528
rect -2969 37493 -2829 37497
rect -2795 37493 -2757 37497
rect -2723 37493 -2685 37497
rect -2651 37493 -2613 37497
rect -2579 37493 -2541 37497
rect -2507 37493 -2469 37497
rect -2435 37493 -2397 37497
rect -2363 37493 -2325 37497
rect -2291 37493 -2253 37497
rect -2219 37493 -2181 37497
rect -2147 37493 -2109 37497
rect -2075 37493 -2037 37497
rect -2003 37493 -1965 37497
rect -1931 37493 -1893 37497
rect -1859 37493 -1821 37497
rect -1787 37493 -1749 37497
rect -1715 37493 -1677 37497
rect -1643 37493 -1605 37497
rect -1571 37493 -1533 37497
rect -1499 37493 -1461 37497
rect -1427 37493 -1389 37497
rect -1355 37493 -1317 37497
rect -1283 37493 -1245 37497
rect -1211 37493 -1173 37497
rect -1139 37493 -1101 37497
rect -1067 37493 -1029 37497
rect -995 37493 -957 37497
rect -923 37493 -885 37497
rect -851 37493 -813 37497
rect -779 37493 -741 37497
rect -707 37493 -669 37497
rect -635 37493 -597 37497
rect -563 37493 -525 37497
rect -491 37493 -453 37497
rect -419 37493 -381 37497
rect -347 37493 -309 37497
rect -275 37493 -153 37497
rect -2969 37459 -2938 37493
rect -2904 37459 -2870 37493
rect -2836 37463 -2829 37493
rect -2768 37463 -2757 37493
rect -2700 37463 -2685 37493
rect -2632 37463 -2613 37493
rect -2564 37463 -2541 37493
rect -2496 37463 -2469 37493
rect -2428 37463 -2397 37493
rect -2836 37459 -2802 37463
rect -2768 37459 -2734 37463
rect -2700 37459 -2666 37463
rect -2632 37459 -2598 37463
rect -2564 37459 -2530 37463
rect -2496 37459 -2462 37463
rect -2428 37459 -2394 37463
rect -2360 37459 -2326 37493
rect -2291 37463 -2258 37493
rect -2219 37463 -2190 37493
rect -2147 37463 -2122 37493
rect -2075 37463 -2054 37493
rect -2003 37463 -1986 37493
rect -1931 37463 -1918 37493
rect -1859 37463 -1850 37493
rect -1787 37463 -1782 37493
rect -1715 37463 -1714 37493
rect -2292 37459 -2258 37463
rect -2224 37459 -2190 37463
rect -2156 37459 -2122 37463
rect -2088 37459 -2054 37463
rect -2020 37459 -1986 37463
rect -1952 37459 -1918 37463
rect -1884 37459 -1850 37463
rect -1816 37459 -1782 37463
rect -1748 37459 -1714 37463
rect -1680 37463 -1677 37493
rect -1612 37463 -1605 37493
rect -1544 37463 -1533 37493
rect -1476 37463 -1461 37493
rect -1408 37463 -1389 37493
rect -1340 37463 -1317 37493
rect -1272 37463 -1245 37493
rect -1204 37463 -1173 37493
rect -1680 37459 -1646 37463
rect -1612 37459 -1578 37463
rect -1544 37459 -1510 37463
rect -1476 37459 -1442 37463
rect -1408 37459 -1374 37463
rect -1340 37459 -1306 37463
rect -1272 37459 -1238 37463
rect -1204 37459 -1170 37463
rect -1136 37459 -1102 37493
rect -1067 37463 -1034 37493
rect -995 37463 -966 37493
rect -923 37463 -898 37493
rect -851 37463 -830 37493
rect -779 37463 -762 37493
rect -707 37463 -694 37493
rect -635 37463 -626 37493
rect -563 37463 -558 37493
rect -491 37463 -490 37493
rect -1068 37459 -1034 37463
rect -1000 37459 -966 37463
rect -932 37459 -898 37463
rect -864 37459 -830 37463
rect -796 37459 -762 37463
rect -728 37459 -694 37463
rect -660 37459 -626 37463
rect -592 37459 -558 37463
rect -524 37459 -490 37463
rect -456 37463 -453 37493
rect -388 37463 -381 37493
rect -320 37463 -309 37493
rect -456 37459 -422 37463
rect -388 37459 -354 37463
rect -320 37459 -286 37463
rect -252 37459 -218 37493
rect -184 37459 -153 37493
rect -2969 37424 -153 37459
rect -2969 37390 -2938 37424
rect -2904 37390 -2870 37424
rect -2836 37390 -2829 37424
rect -2768 37390 -2757 37424
rect -2700 37390 -2685 37424
rect -2632 37390 -2613 37424
rect -2564 37390 -2541 37424
rect -2496 37390 -2469 37424
rect -2428 37390 -2397 37424
rect -2360 37390 -2326 37424
rect -2291 37390 -2258 37424
rect -2219 37390 -2190 37424
rect -2147 37390 -2122 37424
rect -2075 37390 -2054 37424
rect -2003 37390 -1986 37424
rect -1931 37390 -1918 37424
rect -1859 37390 -1850 37424
rect -1787 37390 -1782 37424
rect -1715 37390 -1714 37424
rect -1680 37390 -1677 37424
rect -1612 37390 -1605 37424
rect -1544 37390 -1533 37424
rect -1476 37390 -1461 37424
rect -1408 37390 -1389 37424
rect -1340 37390 -1317 37424
rect -1272 37390 -1245 37424
rect -1204 37390 -1173 37424
rect -1136 37390 -1102 37424
rect -1067 37390 -1034 37424
rect -995 37390 -966 37424
rect -923 37390 -898 37424
rect -851 37390 -830 37424
rect -779 37390 -762 37424
rect -707 37390 -694 37424
rect -635 37390 -626 37424
rect -563 37390 -558 37424
rect -491 37390 -490 37424
rect -456 37390 -453 37424
rect -388 37390 -381 37424
rect -320 37390 -309 37424
rect -252 37390 -218 37424
rect -184 37390 -153 37424
rect -2969 37355 -153 37390
rect -2969 37321 -2938 37355
rect -2904 37321 -2870 37355
rect -2836 37351 -2802 37355
rect -2768 37351 -2734 37355
rect -2700 37351 -2666 37355
rect -2632 37351 -2598 37355
rect -2564 37351 -2530 37355
rect -2496 37351 -2462 37355
rect -2428 37351 -2394 37355
rect -2836 37321 -2829 37351
rect -2768 37321 -2757 37351
rect -2700 37321 -2685 37351
rect -2632 37321 -2613 37351
rect -2564 37321 -2541 37351
rect -2496 37321 -2469 37351
rect -2428 37321 -2397 37351
rect -2360 37321 -2326 37355
rect -2292 37351 -2258 37355
rect -2224 37351 -2190 37355
rect -2156 37351 -2122 37355
rect -2088 37351 -2054 37355
rect -2020 37351 -1986 37355
rect -1952 37351 -1918 37355
rect -1884 37351 -1850 37355
rect -1816 37351 -1782 37355
rect -1748 37351 -1714 37355
rect -2291 37321 -2258 37351
rect -2219 37321 -2190 37351
rect -2147 37321 -2122 37351
rect -2075 37321 -2054 37351
rect -2003 37321 -1986 37351
rect -1931 37321 -1918 37351
rect -1859 37321 -1850 37351
rect -1787 37321 -1782 37351
rect -1715 37321 -1714 37351
rect -1680 37351 -1646 37355
rect -1612 37351 -1578 37355
rect -1544 37351 -1510 37355
rect -1476 37351 -1442 37355
rect -1408 37351 -1374 37355
rect -1340 37351 -1306 37355
rect -1272 37351 -1238 37355
rect -1204 37351 -1170 37355
rect -1680 37321 -1677 37351
rect -1612 37321 -1605 37351
rect -1544 37321 -1533 37351
rect -1476 37321 -1461 37351
rect -1408 37321 -1389 37351
rect -1340 37321 -1317 37351
rect -1272 37321 -1245 37351
rect -1204 37321 -1173 37351
rect -1136 37321 -1102 37355
rect -1068 37351 -1034 37355
rect -1000 37351 -966 37355
rect -932 37351 -898 37355
rect -864 37351 -830 37355
rect -796 37351 -762 37355
rect -728 37351 -694 37355
rect -660 37351 -626 37355
rect -592 37351 -558 37355
rect -524 37351 -490 37355
rect -1067 37321 -1034 37351
rect -995 37321 -966 37351
rect -923 37321 -898 37351
rect -851 37321 -830 37351
rect -779 37321 -762 37351
rect -707 37321 -694 37351
rect -635 37321 -626 37351
rect -563 37321 -558 37351
rect -491 37321 -490 37351
rect -456 37351 -422 37355
rect -388 37351 -354 37355
rect -320 37351 -286 37355
rect -456 37321 -453 37351
rect -388 37321 -381 37351
rect -320 37321 -309 37351
rect -252 37321 -218 37355
rect -184 37321 -153 37355
rect -2969 37317 -2829 37321
rect -2795 37317 -2757 37321
rect -2723 37317 -2685 37321
rect -2651 37317 -2613 37321
rect -2579 37317 -2541 37321
rect -2507 37317 -2469 37321
rect -2435 37317 -2397 37321
rect -2363 37317 -2325 37321
rect -2291 37317 -2253 37321
rect -2219 37317 -2181 37321
rect -2147 37317 -2109 37321
rect -2075 37317 -2037 37321
rect -2003 37317 -1965 37321
rect -1931 37317 -1893 37321
rect -1859 37317 -1821 37321
rect -1787 37317 -1749 37321
rect -1715 37317 -1677 37321
rect -1643 37317 -1605 37321
rect -1571 37317 -1533 37321
rect -1499 37317 -1461 37321
rect -1427 37317 -1389 37321
rect -1355 37317 -1317 37321
rect -1283 37317 -1245 37321
rect -1211 37317 -1173 37321
rect -1139 37317 -1101 37321
rect -1067 37317 -1029 37321
rect -995 37317 -957 37321
rect -923 37317 -885 37321
rect -851 37317 -813 37321
rect -779 37317 -741 37321
rect -707 37317 -669 37321
rect -635 37317 -597 37321
rect -563 37317 -525 37321
rect -491 37317 -453 37321
rect -419 37317 -381 37321
rect -347 37317 -309 37321
rect -275 37317 -153 37321
rect -2969 37286 -153 37317
rect -2969 37252 -2938 37286
rect -2904 37252 -2870 37286
rect -2836 37278 -2802 37286
rect -2768 37278 -2734 37286
rect -2700 37278 -2666 37286
rect -2632 37278 -2598 37286
rect -2564 37278 -2530 37286
rect -2496 37278 -2462 37286
rect -2428 37278 -2394 37286
rect -2836 37252 -2829 37278
rect -2768 37252 -2757 37278
rect -2700 37252 -2685 37278
rect -2632 37252 -2613 37278
rect -2564 37252 -2541 37278
rect -2496 37252 -2469 37278
rect -2428 37252 -2397 37278
rect -2360 37252 -2326 37286
rect -2292 37278 -2258 37286
rect -2224 37278 -2190 37286
rect -2156 37278 -2122 37286
rect -2088 37278 -2054 37286
rect -2020 37278 -1986 37286
rect -1952 37278 -1918 37286
rect -1884 37278 -1850 37286
rect -1816 37278 -1782 37286
rect -1748 37278 -1714 37286
rect -2291 37252 -2258 37278
rect -2219 37252 -2190 37278
rect -2147 37252 -2122 37278
rect -2075 37252 -2054 37278
rect -2003 37252 -1986 37278
rect -1931 37252 -1918 37278
rect -1859 37252 -1850 37278
rect -1787 37252 -1782 37278
rect -1715 37252 -1714 37278
rect -1680 37278 -1646 37286
rect -1612 37278 -1578 37286
rect -1544 37278 -1510 37286
rect -1476 37278 -1442 37286
rect -1408 37278 -1374 37286
rect -1340 37278 -1306 37286
rect -1272 37278 -1238 37286
rect -1204 37278 -1170 37286
rect -1680 37252 -1677 37278
rect -1612 37252 -1605 37278
rect -1544 37252 -1533 37278
rect -1476 37252 -1461 37278
rect -1408 37252 -1389 37278
rect -1340 37252 -1317 37278
rect -1272 37252 -1245 37278
rect -1204 37252 -1173 37278
rect -1136 37252 -1102 37286
rect -1068 37278 -1034 37286
rect -1000 37278 -966 37286
rect -932 37278 -898 37286
rect -864 37278 -830 37286
rect -796 37278 -762 37286
rect -728 37278 -694 37286
rect -660 37278 -626 37286
rect -592 37278 -558 37286
rect -524 37278 -490 37286
rect -1067 37252 -1034 37278
rect -995 37252 -966 37278
rect -923 37252 -898 37278
rect -851 37252 -830 37278
rect -779 37252 -762 37278
rect -707 37252 -694 37278
rect -635 37252 -626 37278
rect -563 37252 -558 37278
rect -491 37252 -490 37278
rect -456 37278 -422 37286
rect -388 37278 -354 37286
rect -320 37278 -286 37286
rect -456 37252 -453 37278
rect -388 37252 -381 37278
rect -320 37252 -309 37278
rect -252 37252 -218 37286
rect -184 37252 -153 37286
rect -2969 37244 -2829 37252
rect -2795 37244 -2757 37252
rect -2723 37244 -2685 37252
rect -2651 37244 -2613 37252
rect -2579 37244 -2541 37252
rect -2507 37244 -2469 37252
rect -2435 37244 -2397 37252
rect -2363 37244 -2325 37252
rect -2291 37244 -2253 37252
rect -2219 37244 -2181 37252
rect -2147 37244 -2109 37252
rect -2075 37244 -2037 37252
rect -2003 37244 -1965 37252
rect -1931 37244 -1893 37252
rect -1859 37244 -1821 37252
rect -1787 37244 -1749 37252
rect -1715 37244 -1677 37252
rect -1643 37244 -1605 37252
rect -1571 37244 -1533 37252
rect -1499 37244 -1461 37252
rect -1427 37244 -1389 37252
rect -1355 37244 -1317 37252
rect -1283 37244 -1245 37252
rect -1211 37244 -1173 37252
rect -1139 37244 -1101 37252
rect -1067 37244 -1029 37252
rect -995 37244 -957 37252
rect -923 37244 -885 37252
rect -851 37244 -813 37252
rect -779 37244 -741 37252
rect -707 37244 -669 37252
rect -635 37244 -597 37252
rect -563 37244 -525 37252
rect -491 37244 -453 37252
rect -419 37244 -381 37252
rect -347 37244 -309 37252
rect -275 37244 -153 37252
rect -2969 37217 -153 37244
rect -2969 37183 -2938 37217
rect -2904 37183 -2870 37217
rect -2836 37205 -2802 37217
rect -2768 37205 -2734 37217
rect -2700 37205 -2666 37217
rect -2632 37205 -2598 37217
rect -2564 37205 -2530 37217
rect -2496 37205 -2462 37217
rect -2428 37205 -2394 37217
rect -2836 37183 -2829 37205
rect -2768 37183 -2757 37205
rect -2700 37183 -2685 37205
rect -2632 37183 -2613 37205
rect -2564 37183 -2541 37205
rect -2496 37183 -2469 37205
rect -2428 37183 -2397 37205
rect -2360 37183 -2326 37217
rect -2292 37205 -2258 37217
rect -2224 37205 -2190 37217
rect -2156 37205 -2122 37217
rect -2088 37205 -2054 37217
rect -2020 37205 -1986 37217
rect -1952 37205 -1918 37217
rect -1884 37205 -1850 37217
rect -1816 37205 -1782 37217
rect -1748 37205 -1714 37217
rect -2291 37183 -2258 37205
rect -2219 37183 -2190 37205
rect -2147 37183 -2122 37205
rect -2075 37183 -2054 37205
rect -2003 37183 -1986 37205
rect -1931 37183 -1918 37205
rect -1859 37183 -1850 37205
rect -1787 37183 -1782 37205
rect -1715 37183 -1714 37205
rect -1680 37205 -1646 37217
rect -1612 37205 -1578 37217
rect -1544 37205 -1510 37217
rect -1476 37205 -1442 37217
rect -1408 37205 -1374 37217
rect -1340 37205 -1306 37217
rect -1272 37205 -1238 37217
rect -1204 37205 -1170 37217
rect -1680 37183 -1677 37205
rect -1612 37183 -1605 37205
rect -1544 37183 -1533 37205
rect -1476 37183 -1461 37205
rect -1408 37183 -1389 37205
rect -1340 37183 -1317 37205
rect -1272 37183 -1245 37205
rect -1204 37183 -1173 37205
rect -1136 37183 -1102 37217
rect -1068 37205 -1034 37217
rect -1000 37205 -966 37217
rect -932 37205 -898 37217
rect -864 37205 -830 37217
rect -796 37205 -762 37217
rect -728 37205 -694 37217
rect -660 37205 -626 37217
rect -592 37205 -558 37217
rect -524 37205 -490 37217
rect -1067 37183 -1034 37205
rect -995 37183 -966 37205
rect -923 37183 -898 37205
rect -851 37183 -830 37205
rect -779 37183 -762 37205
rect -707 37183 -694 37205
rect -635 37183 -626 37205
rect -563 37183 -558 37205
rect -491 37183 -490 37205
rect -456 37205 -422 37217
rect -388 37205 -354 37217
rect -320 37205 -286 37217
rect -456 37183 -453 37205
rect -388 37183 -381 37205
rect -320 37183 -309 37205
rect -252 37183 -218 37217
rect -184 37183 -153 37217
rect -2969 37171 -2829 37183
rect -2795 37171 -2757 37183
rect -2723 37171 -2685 37183
rect -2651 37171 -2613 37183
rect -2579 37171 -2541 37183
rect -2507 37171 -2469 37183
rect -2435 37171 -2397 37183
rect -2363 37171 -2325 37183
rect -2291 37171 -2253 37183
rect -2219 37171 -2181 37183
rect -2147 37171 -2109 37183
rect -2075 37171 -2037 37183
rect -2003 37171 -1965 37183
rect -1931 37171 -1893 37183
rect -1859 37171 -1821 37183
rect -1787 37171 -1749 37183
rect -1715 37171 -1677 37183
rect -1643 37171 -1605 37183
rect -1571 37171 -1533 37183
rect -1499 37171 -1461 37183
rect -1427 37171 -1389 37183
rect -1355 37171 -1317 37183
rect -1283 37171 -1245 37183
rect -1211 37171 -1173 37183
rect -1139 37171 -1101 37183
rect -1067 37171 -1029 37183
rect -995 37171 -957 37183
rect -923 37171 -885 37183
rect -851 37171 -813 37183
rect -779 37171 -741 37183
rect -707 37171 -669 37183
rect -635 37171 -597 37183
rect -563 37171 -525 37183
rect -491 37171 -453 37183
rect -419 37171 -381 37183
rect -347 37171 -309 37183
rect -275 37171 -153 37183
rect -2969 37148 -153 37171
rect -2969 37114 -2938 37148
rect -2904 37114 -2870 37148
rect -2836 37132 -2802 37148
rect -2768 37132 -2734 37148
rect -2700 37132 -2666 37148
rect -2632 37132 -2598 37148
rect -2564 37132 -2530 37148
rect -2496 37132 -2462 37148
rect -2428 37132 -2394 37148
rect -2836 37114 -2829 37132
rect -2768 37114 -2757 37132
rect -2700 37114 -2685 37132
rect -2632 37114 -2613 37132
rect -2564 37114 -2541 37132
rect -2496 37114 -2469 37132
rect -2428 37114 -2397 37132
rect -2360 37114 -2326 37148
rect -2292 37132 -2258 37148
rect -2224 37132 -2190 37148
rect -2156 37132 -2122 37148
rect -2088 37132 -2054 37148
rect -2020 37132 -1986 37148
rect -1952 37132 -1918 37148
rect -1884 37132 -1850 37148
rect -1816 37132 -1782 37148
rect -1748 37132 -1714 37148
rect -2291 37114 -2258 37132
rect -2219 37114 -2190 37132
rect -2147 37114 -2122 37132
rect -2075 37114 -2054 37132
rect -2003 37114 -1986 37132
rect -1931 37114 -1918 37132
rect -1859 37114 -1850 37132
rect -1787 37114 -1782 37132
rect -1715 37114 -1714 37132
rect -1680 37132 -1646 37148
rect -1612 37132 -1578 37148
rect -1544 37132 -1510 37148
rect -1476 37132 -1442 37148
rect -1408 37132 -1374 37148
rect -1340 37132 -1306 37148
rect -1272 37132 -1238 37148
rect -1204 37132 -1170 37148
rect -1680 37114 -1677 37132
rect -1612 37114 -1605 37132
rect -1544 37114 -1533 37132
rect -1476 37114 -1461 37132
rect -1408 37114 -1389 37132
rect -1340 37114 -1317 37132
rect -1272 37114 -1245 37132
rect -1204 37114 -1173 37132
rect -1136 37114 -1102 37148
rect -1068 37132 -1034 37148
rect -1000 37132 -966 37148
rect -932 37132 -898 37148
rect -864 37132 -830 37148
rect -796 37132 -762 37148
rect -728 37132 -694 37148
rect -660 37132 -626 37148
rect -592 37132 -558 37148
rect -524 37132 -490 37148
rect -1067 37114 -1034 37132
rect -995 37114 -966 37132
rect -923 37114 -898 37132
rect -851 37114 -830 37132
rect -779 37114 -762 37132
rect -707 37114 -694 37132
rect -635 37114 -626 37132
rect -563 37114 -558 37132
rect -491 37114 -490 37132
rect -456 37132 -422 37148
rect -388 37132 -354 37148
rect -320 37132 -286 37148
rect -456 37114 -453 37132
rect -388 37114 -381 37132
rect -320 37114 -309 37132
rect -252 37114 -218 37148
rect -184 37114 -153 37148
rect -2969 37098 -2829 37114
rect -2795 37098 -2757 37114
rect -2723 37098 -2685 37114
rect -2651 37098 -2613 37114
rect -2579 37098 -2541 37114
rect -2507 37098 -2469 37114
rect -2435 37098 -2397 37114
rect -2363 37098 -2325 37114
rect -2291 37098 -2253 37114
rect -2219 37098 -2181 37114
rect -2147 37098 -2109 37114
rect -2075 37098 -2037 37114
rect -2003 37098 -1965 37114
rect -1931 37098 -1893 37114
rect -1859 37098 -1821 37114
rect -1787 37098 -1749 37114
rect -1715 37098 -1677 37114
rect -1643 37098 -1605 37114
rect -1571 37098 -1533 37114
rect -1499 37098 -1461 37114
rect -1427 37098 -1389 37114
rect -1355 37098 -1317 37114
rect -1283 37098 -1245 37114
rect -1211 37098 -1173 37114
rect -1139 37098 -1101 37114
rect -1067 37098 -1029 37114
rect -995 37098 -957 37114
rect -923 37098 -885 37114
rect -851 37098 -813 37114
rect -779 37098 -741 37114
rect -707 37098 -669 37114
rect -635 37098 -597 37114
rect -563 37098 -525 37114
rect -491 37098 -453 37114
rect -419 37098 -381 37114
rect -347 37098 -309 37114
rect -275 37098 -153 37114
rect -2969 37079 -153 37098
rect -2969 37045 -2938 37079
rect -2904 37045 -2870 37079
rect -2836 37059 -2802 37079
rect -2768 37059 -2734 37079
rect -2700 37059 -2666 37079
rect -2632 37059 -2598 37079
rect -2564 37059 -2530 37079
rect -2496 37059 -2462 37079
rect -2428 37059 -2394 37079
rect -2836 37045 -2829 37059
rect -2768 37045 -2757 37059
rect -2700 37045 -2685 37059
rect -2632 37045 -2613 37059
rect -2564 37045 -2541 37059
rect -2496 37045 -2469 37059
rect -2428 37045 -2397 37059
rect -2360 37045 -2326 37079
rect -2292 37059 -2258 37079
rect -2224 37059 -2190 37079
rect -2156 37059 -2122 37079
rect -2088 37059 -2054 37079
rect -2020 37059 -1986 37079
rect -1952 37059 -1918 37079
rect -1884 37059 -1850 37079
rect -1816 37059 -1782 37079
rect -1748 37059 -1714 37079
rect -2291 37045 -2258 37059
rect -2219 37045 -2190 37059
rect -2147 37045 -2122 37059
rect -2075 37045 -2054 37059
rect -2003 37045 -1986 37059
rect -1931 37045 -1918 37059
rect -1859 37045 -1850 37059
rect -1787 37045 -1782 37059
rect -1715 37045 -1714 37059
rect -1680 37059 -1646 37079
rect -1612 37059 -1578 37079
rect -1544 37059 -1510 37079
rect -1476 37059 -1442 37079
rect -1408 37059 -1374 37079
rect -1340 37059 -1306 37079
rect -1272 37059 -1238 37079
rect -1204 37059 -1170 37079
rect -1680 37045 -1677 37059
rect -1612 37045 -1605 37059
rect -1544 37045 -1533 37059
rect -1476 37045 -1461 37059
rect -1408 37045 -1389 37059
rect -1340 37045 -1317 37059
rect -1272 37045 -1245 37059
rect -1204 37045 -1173 37059
rect -1136 37045 -1102 37079
rect -1068 37059 -1034 37079
rect -1000 37059 -966 37079
rect -932 37059 -898 37079
rect -864 37059 -830 37079
rect -796 37059 -762 37079
rect -728 37059 -694 37079
rect -660 37059 -626 37079
rect -592 37059 -558 37079
rect -524 37059 -490 37079
rect -1067 37045 -1034 37059
rect -995 37045 -966 37059
rect -923 37045 -898 37059
rect -851 37045 -830 37059
rect -779 37045 -762 37059
rect -707 37045 -694 37059
rect -635 37045 -626 37059
rect -563 37045 -558 37059
rect -491 37045 -490 37059
rect -456 37059 -422 37079
rect -388 37059 -354 37079
rect -320 37059 -286 37079
rect -456 37045 -453 37059
rect -388 37045 -381 37059
rect -320 37045 -309 37059
rect -252 37045 -218 37079
rect -184 37045 -153 37079
rect -2969 37025 -2829 37045
rect -2795 37025 -2757 37045
rect -2723 37025 -2685 37045
rect -2651 37025 -2613 37045
rect -2579 37025 -2541 37045
rect -2507 37025 -2469 37045
rect -2435 37025 -2397 37045
rect -2363 37025 -2325 37045
rect -2291 37025 -2253 37045
rect -2219 37025 -2181 37045
rect -2147 37025 -2109 37045
rect -2075 37025 -2037 37045
rect -2003 37025 -1965 37045
rect -1931 37025 -1893 37045
rect -1859 37025 -1821 37045
rect -1787 37025 -1749 37045
rect -1715 37025 -1677 37045
rect -1643 37025 -1605 37045
rect -1571 37025 -1533 37045
rect -1499 37025 -1461 37045
rect -1427 37025 -1389 37045
rect -1355 37025 -1317 37045
rect -1283 37025 -1245 37045
rect -1211 37025 -1173 37045
rect -1139 37025 -1101 37045
rect -1067 37025 -1029 37045
rect -995 37025 -957 37045
rect -923 37025 -885 37045
rect -851 37025 -813 37045
rect -779 37025 -741 37045
rect -707 37025 -669 37045
rect -635 37025 -597 37045
rect -563 37025 -525 37045
rect -491 37025 -453 37045
rect -419 37025 -381 37045
rect -347 37025 -309 37045
rect -275 37025 -153 37045
rect -2969 37010 -153 37025
rect -2969 36976 -2938 37010
rect -2904 36976 -2870 37010
rect -2836 36986 -2802 37010
rect -2768 36986 -2734 37010
rect -2700 36986 -2666 37010
rect -2632 36986 -2598 37010
rect -2564 36986 -2530 37010
rect -2496 36986 -2462 37010
rect -2428 36986 -2394 37010
rect -2836 36976 -2829 36986
rect -2768 36976 -2757 36986
rect -2700 36976 -2685 36986
rect -2632 36976 -2613 36986
rect -2564 36976 -2541 36986
rect -2496 36976 -2469 36986
rect -2428 36976 -2397 36986
rect -2360 36976 -2326 37010
rect -2292 36986 -2258 37010
rect -2224 36986 -2190 37010
rect -2156 36986 -2122 37010
rect -2088 36986 -2054 37010
rect -2020 36986 -1986 37010
rect -1952 36986 -1918 37010
rect -1884 36986 -1850 37010
rect -1816 36986 -1782 37010
rect -1748 36986 -1714 37010
rect -2291 36976 -2258 36986
rect -2219 36976 -2190 36986
rect -2147 36976 -2122 36986
rect -2075 36976 -2054 36986
rect -2003 36976 -1986 36986
rect -1931 36976 -1918 36986
rect -1859 36976 -1850 36986
rect -1787 36976 -1782 36986
rect -1715 36976 -1714 36986
rect -1680 36986 -1646 37010
rect -1612 36986 -1578 37010
rect -1544 36986 -1510 37010
rect -1476 36986 -1442 37010
rect -1408 36986 -1374 37010
rect -1340 36986 -1306 37010
rect -1272 36986 -1238 37010
rect -1204 36986 -1170 37010
rect -1680 36976 -1677 36986
rect -1612 36976 -1605 36986
rect -1544 36976 -1533 36986
rect -1476 36976 -1461 36986
rect -1408 36976 -1389 36986
rect -1340 36976 -1317 36986
rect -1272 36976 -1245 36986
rect -1204 36976 -1173 36986
rect -1136 36976 -1102 37010
rect -1068 36986 -1034 37010
rect -1000 36986 -966 37010
rect -932 36986 -898 37010
rect -864 36986 -830 37010
rect -796 36986 -762 37010
rect -728 36986 -694 37010
rect -660 36986 -626 37010
rect -592 36986 -558 37010
rect -524 36986 -490 37010
rect -1067 36976 -1034 36986
rect -995 36976 -966 36986
rect -923 36976 -898 36986
rect -851 36976 -830 36986
rect -779 36976 -762 36986
rect -707 36976 -694 36986
rect -635 36976 -626 36986
rect -563 36976 -558 36986
rect -491 36976 -490 36986
rect -456 36986 -422 37010
rect -388 36986 -354 37010
rect -320 36986 -286 37010
rect -456 36976 -453 36986
rect -388 36976 -381 36986
rect -320 36976 -309 36986
rect -252 36976 -218 37010
rect -184 36976 -153 37010
rect -2969 36952 -2829 36976
rect -2795 36952 -2757 36976
rect -2723 36952 -2685 36976
rect -2651 36952 -2613 36976
rect -2579 36952 -2541 36976
rect -2507 36952 -2469 36976
rect -2435 36952 -2397 36976
rect -2363 36952 -2325 36976
rect -2291 36952 -2253 36976
rect -2219 36952 -2181 36976
rect -2147 36952 -2109 36976
rect -2075 36952 -2037 36976
rect -2003 36952 -1965 36976
rect -1931 36952 -1893 36976
rect -1859 36952 -1821 36976
rect -1787 36952 -1749 36976
rect -1715 36952 -1677 36976
rect -1643 36952 -1605 36976
rect -1571 36952 -1533 36976
rect -1499 36952 -1461 36976
rect -1427 36952 -1389 36976
rect -1355 36952 -1317 36976
rect -1283 36952 -1245 36976
rect -1211 36952 -1173 36976
rect -1139 36952 -1101 36976
rect -1067 36952 -1029 36976
rect -995 36952 -957 36976
rect -923 36952 -885 36976
rect -851 36952 -813 36976
rect -779 36952 -741 36976
rect -707 36952 -669 36976
rect -635 36952 -597 36976
rect -563 36952 -525 36976
rect -491 36952 -453 36976
rect -419 36952 -381 36976
rect -347 36952 -309 36976
rect -275 36952 -153 36976
rect -2969 36941 -153 36952
rect -2969 36907 -2938 36941
rect -2904 36907 -2870 36941
rect -2836 36913 -2802 36941
rect -2768 36913 -2734 36941
rect -2700 36913 -2666 36941
rect -2632 36913 -2598 36941
rect -2564 36913 -2530 36941
rect -2496 36913 -2462 36941
rect -2428 36913 -2394 36941
rect -2836 36907 -2829 36913
rect -2768 36907 -2757 36913
rect -2700 36907 -2685 36913
rect -2632 36907 -2613 36913
rect -2564 36907 -2541 36913
rect -2496 36907 -2469 36913
rect -2428 36907 -2397 36913
rect -2360 36907 -2326 36941
rect -2292 36913 -2258 36941
rect -2224 36913 -2190 36941
rect -2156 36913 -2122 36941
rect -2088 36913 -2054 36941
rect -2020 36913 -1986 36941
rect -1952 36913 -1918 36941
rect -1884 36913 -1850 36941
rect -1816 36913 -1782 36941
rect -1748 36913 -1714 36941
rect -2291 36907 -2258 36913
rect -2219 36907 -2190 36913
rect -2147 36907 -2122 36913
rect -2075 36907 -2054 36913
rect -2003 36907 -1986 36913
rect -1931 36907 -1918 36913
rect -1859 36907 -1850 36913
rect -1787 36907 -1782 36913
rect -1715 36907 -1714 36913
rect -1680 36913 -1646 36941
rect -1612 36913 -1578 36941
rect -1544 36913 -1510 36941
rect -1476 36913 -1442 36941
rect -1408 36913 -1374 36941
rect -1340 36913 -1306 36941
rect -1272 36913 -1238 36941
rect -1204 36913 -1170 36941
rect -1680 36907 -1677 36913
rect -1612 36907 -1605 36913
rect -1544 36907 -1533 36913
rect -1476 36907 -1461 36913
rect -1408 36907 -1389 36913
rect -1340 36907 -1317 36913
rect -1272 36907 -1245 36913
rect -1204 36907 -1173 36913
rect -1136 36907 -1102 36941
rect -1068 36913 -1034 36941
rect -1000 36913 -966 36941
rect -932 36913 -898 36941
rect -864 36913 -830 36941
rect -796 36913 -762 36941
rect -728 36913 -694 36941
rect -660 36913 -626 36941
rect -592 36913 -558 36941
rect -524 36913 -490 36941
rect -1067 36907 -1034 36913
rect -995 36907 -966 36913
rect -923 36907 -898 36913
rect -851 36907 -830 36913
rect -779 36907 -762 36913
rect -707 36907 -694 36913
rect -635 36907 -626 36913
rect -563 36907 -558 36913
rect -491 36907 -490 36913
rect -456 36913 -422 36941
rect -388 36913 -354 36941
rect -320 36913 -286 36941
rect -456 36907 -453 36913
rect -388 36907 -381 36913
rect -320 36907 -309 36913
rect -252 36907 -218 36941
rect -184 36907 -153 36941
rect -2969 36879 -2829 36907
rect -2795 36879 -2757 36907
rect -2723 36879 -2685 36907
rect -2651 36879 -2613 36907
rect -2579 36879 -2541 36907
rect -2507 36879 -2469 36907
rect -2435 36879 -2397 36907
rect -2363 36879 -2325 36907
rect -2291 36879 -2253 36907
rect -2219 36879 -2181 36907
rect -2147 36879 -2109 36907
rect -2075 36879 -2037 36907
rect -2003 36879 -1965 36907
rect -1931 36879 -1893 36907
rect -1859 36879 -1821 36907
rect -1787 36879 -1749 36907
rect -1715 36879 -1677 36907
rect -1643 36879 -1605 36907
rect -1571 36879 -1533 36907
rect -1499 36879 -1461 36907
rect -1427 36879 -1389 36907
rect -1355 36879 -1317 36907
rect -1283 36879 -1245 36907
rect -1211 36879 -1173 36907
rect -1139 36879 -1101 36907
rect -1067 36879 -1029 36907
rect -995 36879 -957 36907
rect -923 36879 -885 36907
rect -851 36879 -813 36907
rect -779 36879 -741 36907
rect -707 36879 -669 36907
rect -635 36879 -597 36907
rect -563 36879 -525 36907
rect -491 36879 -453 36907
rect -419 36879 -381 36907
rect -347 36879 -309 36907
rect -275 36879 -153 36907
rect -2969 36872 -153 36879
rect -2969 36838 -2938 36872
rect -2904 36838 -2870 36872
rect -2836 36840 -2802 36872
rect -2768 36840 -2734 36872
rect -2700 36840 -2666 36872
rect -2632 36840 -2598 36872
rect -2564 36840 -2530 36872
rect -2496 36840 -2462 36872
rect -2428 36840 -2394 36872
rect -2836 36838 -2829 36840
rect -2768 36838 -2757 36840
rect -2700 36838 -2685 36840
rect -2632 36838 -2613 36840
rect -2564 36838 -2541 36840
rect -2496 36838 -2469 36840
rect -2428 36838 -2397 36840
rect -2360 36838 -2326 36872
rect -2292 36840 -2258 36872
rect -2224 36840 -2190 36872
rect -2156 36840 -2122 36872
rect -2088 36840 -2054 36872
rect -2020 36840 -1986 36872
rect -1952 36840 -1918 36872
rect -1884 36840 -1850 36872
rect -1816 36840 -1782 36872
rect -1748 36840 -1714 36872
rect -2291 36838 -2258 36840
rect -2219 36838 -2190 36840
rect -2147 36838 -2122 36840
rect -2075 36838 -2054 36840
rect -2003 36838 -1986 36840
rect -1931 36838 -1918 36840
rect -1859 36838 -1850 36840
rect -1787 36838 -1782 36840
rect -1715 36838 -1714 36840
rect -1680 36840 -1646 36872
rect -1612 36840 -1578 36872
rect -1544 36840 -1510 36872
rect -1476 36840 -1442 36872
rect -1408 36840 -1374 36872
rect -1340 36840 -1306 36872
rect -1272 36840 -1238 36872
rect -1204 36840 -1170 36872
rect -1680 36838 -1677 36840
rect -1612 36838 -1605 36840
rect -1544 36838 -1533 36840
rect -1476 36838 -1461 36840
rect -1408 36838 -1389 36840
rect -1340 36838 -1317 36840
rect -1272 36838 -1245 36840
rect -1204 36838 -1173 36840
rect -1136 36838 -1102 36872
rect -1068 36840 -1034 36872
rect -1000 36840 -966 36872
rect -932 36840 -898 36872
rect -864 36840 -830 36872
rect -796 36840 -762 36872
rect -728 36840 -694 36872
rect -660 36840 -626 36872
rect -592 36840 -558 36872
rect -524 36840 -490 36872
rect -1067 36838 -1034 36840
rect -995 36838 -966 36840
rect -923 36838 -898 36840
rect -851 36838 -830 36840
rect -779 36838 -762 36840
rect -707 36838 -694 36840
rect -635 36838 -626 36840
rect -563 36838 -558 36840
rect -491 36838 -490 36840
rect -456 36840 -422 36872
rect -388 36840 -354 36872
rect -320 36840 -286 36872
rect -456 36838 -453 36840
rect -388 36838 -381 36840
rect -320 36838 -309 36840
rect -252 36838 -218 36872
rect -184 36838 -153 36872
rect -2969 36806 -2829 36838
rect -2795 36806 -2757 36838
rect -2723 36806 -2685 36838
rect -2651 36806 -2613 36838
rect -2579 36806 -2541 36838
rect -2507 36806 -2469 36838
rect -2435 36806 -2397 36838
rect -2363 36806 -2325 36838
rect -2291 36806 -2253 36838
rect -2219 36806 -2181 36838
rect -2147 36806 -2109 36838
rect -2075 36806 -2037 36838
rect -2003 36806 -1965 36838
rect -1931 36806 -1893 36838
rect -1859 36806 -1821 36838
rect -1787 36806 -1749 36838
rect -1715 36806 -1677 36838
rect -1643 36806 -1605 36838
rect -1571 36806 -1533 36838
rect -1499 36806 -1461 36838
rect -1427 36806 -1389 36838
rect -1355 36806 -1317 36838
rect -1283 36806 -1245 36838
rect -1211 36806 -1173 36838
rect -1139 36806 -1101 36838
rect -1067 36806 -1029 36838
rect -995 36806 -957 36838
rect -923 36806 -885 36838
rect -851 36806 -813 36838
rect -779 36806 -741 36838
rect -707 36806 -669 36838
rect -635 36806 -597 36838
rect -563 36806 -525 36838
rect -491 36806 -453 36838
rect -419 36806 -381 36838
rect -347 36806 -309 36838
rect -275 36806 -153 36838
rect -2969 36803 -153 36806
rect -2969 36769 -2938 36803
rect -2904 36769 -2870 36803
rect -2836 36769 -2802 36803
rect -2768 36769 -2734 36803
rect -2700 36769 -2666 36803
rect -2632 36769 -2598 36803
rect -2564 36769 -2530 36803
rect -2496 36769 -2462 36803
rect -2428 36769 -2394 36803
rect -2360 36769 -2326 36803
rect -2292 36769 -2258 36803
rect -2224 36769 -2190 36803
rect -2156 36769 -2122 36803
rect -2088 36769 -2054 36803
rect -2020 36769 -1986 36803
rect -1952 36769 -1918 36803
rect -1884 36769 -1850 36803
rect -1816 36769 -1782 36803
rect -1748 36769 -1714 36803
rect -1680 36769 -1646 36803
rect -1612 36769 -1578 36803
rect -1544 36769 -1510 36803
rect -1476 36769 -1442 36803
rect -1408 36769 -1374 36803
rect -1340 36769 -1306 36803
rect -1272 36769 -1238 36803
rect -1204 36769 -1170 36803
rect -1136 36769 -1102 36803
rect -1068 36769 -1034 36803
rect -1000 36769 -966 36803
rect -932 36769 -898 36803
rect -864 36769 -830 36803
rect -796 36769 -762 36803
rect -728 36769 -694 36803
rect -660 36769 -626 36803
rect -592 36769 -558 36803
rect -524 36769 -490 36803
rect -456 36769 -422 36803
rect -388 36769 -354 36803
rect -320 36769 -286 36803
rect -252 36769 -218 36803
rect -184 36769 -153 36803
rect -2969 36767 -153 36769
rect -2969 36734 -2829 36767
rect -2795 36734 -2757 36767
rect -2723 36734 -2685 36767
rect -2651 36734 -2613 36767
rect -2579 36734 -2541 36767
rect -2507 36734 -2469 36767
rect -2435 36734 -2397 36767
rect -2363 36734 -2325 36767
rect -2291 36734 -2253 36767
rect -2219 36734 -2181 36767
rect -2147 36734 -2109 36767
rect -2075 36734 -2037 36767
rect -2003 36734 -1965 36767
rect -1931 36734 -1893 36767
rect -1859 36734 -1821 36767
rect -1787 36734 -1749 36767
rect -1715 36734 -1677 36767
rect -1643 36734 -1605 36767
rect -1571 36734 -1533 36767
rect -1499 36734 -1461 36767
rect -1427 36734 -1389 36767
rect -1355 36734 -1317 36767
rect -1283 36734 -1245 36767
rect -1211 36734 -1173 36767
rect -1139 36734 -1101 36767
rect -1067 36734 -1029 36767
rect -995 36734 -957 36767
rect -923 36734 -885 36767
rect -851 36734 -813 36767
rect -779 36734 -741 36767
rect -707 36734 -669 36767
rect -635 36734 -597 36767
rect -563 36734 -525 36767
rect -491 36734 -453 36767
rect -419 36734 -381 36767
rect -347 36734 -309 36767
rect -275 36734 -153 36767
rect -2969 36700 -2938 36734
rect -2904 36700 -2870 36734
rect -2836 36733 -2829 36734
rect -2768 36733 -2757 36734
rect -2700 36733 -2685 36734
rect -2632 36733 -2613 36734
rect -2564 36733 -2541 36734
rect -2496 36733 -2469 36734
rect -2428 36733 -2397 36734
rect -2836 36700 -2802 36733
rect -2768 36700 -2734 36733
rect -2700 36700 -2666 36733
rect -2632 36700 -2598 36733
rect -2564 36700 -2530 36733
rect -2496 36700 -2462 36733
rect -2428 36700 -2394 36733
rect -2360 36700 -2326 36734
rect -2291 36733 -2258 36734
rect -2219 36733 -2190 36734
rect -2147 36733 -2122 36734
rect -2075 36733 -2054 36734
rect -2003 36733 -1986 36734
rect -1931 36733 -1918 36734
rect -1859 36733 -1850 36734
rect -1787 36733 -1782 36734
rect -1715 36733 -1714 36734
rect -2292 36700 -2258 36733
rect -2224 36700 -2190 36733
rect -2156 36700 -2122 36733
rect -2088 36700 -2054 36733
rect -2020 36700 -1986 36733
rect -1952 36700 -1918 36733
rect -1884 36700 -1850 36733
rect -1816 36700 -1782 36733
rect -1748 36700 -1714 36733
rect -1680 36733 -1677 36734
rect -1612 36733 -1605 36734
rect -1544 36733 -1533 36734
rect -1476 36733 -1461 36734
rect -1408 36733 -1389 36734
rect -1340 36733 -1317 36734
rect -1272 36733 -1245 36734
rect -1204 36733 -1173 36734
rect -1680 36700 -1646 36733
rect -1612 36700 -1578 36733
rect -1544 36700 -1510 36733
rect -1476 36700 -1442 36733
rect -1408 36700 -1374 36733
rect -1340 36700 -1306 36733
rect -1272 36700 -1238 36733
rect -1204 36700 -1170 36733
rect -1136 36700 -1102 36734
rect -1067 36733 -1034 36734
rect -995 36733 -966 36734
rect -923 36733 -898 36734
rect -851 36733 -830 36734
rect -779 36733 -762 36734
rect -707 36733 -694 36734
rect -635 36733 -626 36734
rect -563 36733 -558 36734
rect -491 36733 -490 36734
rect -1068 36700 -1034 36733
rect -1000 36700 -966 36733
rect -932 36700 -898 36733
rect -864 36700 -830 36733
rect -796 36700 -762 36733
rect -728 36700 -694 36733
rect -660 36700 -626 36733
rect -592 36700 -558 36733
rect -524 36700 -490 36733
rect -456 36733 -453 36734
rect -388 36733 -381 36734
rect -320 36733 -309 36734
rect -456 36700 -422 36733
rect -388 36700 -354 36733
rect -320 36700 -286 36733
rect -252 36700 -218 36734
rect -184 36700 -153 36734
rect -2969 36694 -153 36700
rect -2969 36665 -2829 36694
rect -2795 36665 -2757 36694
rect -2723 36665 -2685 36694
rect -2651 36665 -2613 36694
rect -2579 36665 -2541 36694
rect -2507 36665 -2469 36694
rect -2435 36665 -2397 36694
rect -2363 36665 -2325 36694
rect -2291 36665 -2253 36694
rect -2219 36665 -2181 36694
rect -2147 36665 -2109 36694
rect -2075 36665 -2037 36694
rect -2003 36665 -1965 36694
rect -1931 36665 -1893 36694
rect -1859 36665 -1821 36694
rect -1787 36665 -1749 36694
rect -1715 36665 -1677 36694
rect -1643 36665 -1605 36694
rect -1571 36665 -1533 36694
rect -1499 36665 -1461 36694
rect -1427 36665 -1389 36694
rect -1355 36665 -1317 36694
rect -1283 36665 -1245 36694
rect -1211 36665 -1173 36694
rect -1139 36665 -1101 36694
rect -1067 36665 -1029 36694
rect -995 36665 -957 36694
rect -923 36665 -885 36694
rect -851 36665 -813 36694
rect -779 36665 -741 36694
rect -707 36665 -669 36694
rect -635 36665 -597 36694
rect -563 36665 -525 36694
rect -491 36665 -453 36694
rect -419 36665 -381 36694
rect -347 36665 -309 36694
rect -275 36665 -153 36694
rect -2969 36631 -2938 36665
rect -2904 36631 -2870 36665
rect -2836 36660 -2829 36665
rect -2768 36660 -2757 36665
rect -2700 36660 -2685 36665
rect -2632 36660 -2613 36665
rect -2564 36660 -2541 36665
rect -2496 36660 -2469 36665
rect -2428 36660 -2397 36665
rect -2836 36631 -2802 36660
rect -2768 36631 -2734 36660
rect -2700 36631 -2666 36660
rect -2632 36631 -2598 36660
rect -2564 36631 -2530 36660
rect -2496 36631 -2462 36660
rect -2428 36631 -2394 36660
rect -2360 36631 -2326 36665
rect -2291 36660 -2258 36665
rect -2219 36660 -2190 36665
rect -2147 36660 -2122 36665
rect -2075 36660 -2054 36665
rect -2003 36660 -1986 36665
rect -1931 36660 -1918 36665
rect -1859 36660 -1850 36665
rect -1787 36660 -1782 36665
rect -1715 36660 -1714 36665
rect -2292 36631 -2258 36660
rect -2224 36631 -2190 36660
rect -2156 36631 -2122 36660
rect -2088 36631 -2054 36660
rect -2020 36631 -1986 36660
rect -1952 36631 -1918 36660
rect -1884 36631 -1850 36660
rect -1816 36631 -1782 36660
rect -1748 36631 -1714 36660
rect -1680 36660 -1677 36665
rect -1612 36660 -1605 36665
rect -1544 36660 -1533 36665
rect -1476 36660 -1461 36665
rect -1408 36660 -1389 36665
rect -1340 36660 -1317 36665
rect -1272 36660 -1245 36665
rect -1204 36660 -1173 36665
rect -1680 36631 -1646 36660
rect -1612 36631 -1578 36660
rect -1544 36631 -1510 36660
rect -1476 36631 -1442 36660
rect -1408 36631 -1374 36660
rect -1340 36631 -1306 36660
rect -1272 36631 -1238 36660
rect -1204 36631 -1170 36660
rect -1136 36631 -1102 36665
rect -1067 36660 -1034 36665
rect -995 36660 -966 36665
rect -923 36660 -898 36665
rect -851 36660 -830 36665
rect -779 36660 -762 36665
rect -707 36660 -694 36665
rect -635 36660 -626 36665
rect -563 36660 -558 36665
rect -491 36660 -490 36665
rect -1068 36631 -1034 36660
rect -1000 36631 -966 36660
rect -932 36631 -898 36660
rect -864 36631 -830 36660
rect -796 36631 -762 36660
rect -728 36631 -694 36660
rect -660 36631 -626 36660
rect -592 36631 -558 36660
rect -524 36631 -490 36660
rect -456 36660 -453 36665
rect -388 36660 -381 36665
rect -320 36660 -309 36665
rect -456 36631 -422 36660
rect -388 36631 -354 36660
rect -320 36631 -286 36660
rect -252 36631 -218 36665
rect -184 36631 -153 36665
rect -2969 36621 -153 36631
rect -2969 36596 -2829 36621
rect -2795 36596 -2757 36621
rect -2723 36596 -2685 36621
rect -2651 36596 -2613 36621
rect -2579 36596 -2541 36621
rect -2507 36596 -2469 36621
rect -2435 36596 -2397 36621
rect -2363 36596 -2325 36621
rect -2291 36596 -2253 36621
rect -2219 36596 -2181 36621
rect -2147 36596 -2109 36621
rect -2075 36596 -2037 36621
rect -2003 36596 -1965 36621
rect -1931 36596 -1893 36621
rect -1859 36596 -1821 36621
rect -1787 36596 -1749 36621
rect -1715 36596 -1677 36621
rect -1643 36596 -1605 36621
rect -1571 36596 -1533 36621
rect -1499 36596 -1461 36621
rect -1427 36596 -1389 36621
rect -1355 36596 -1317 36621
rect -1283 36596 -1245 36621
rect -1211 36596 -1173 36621
rect -1139 36596 -1101 36621
rect -1067 36596 -1029 36621
rect -995 36596 -957 36621
rect -923 36596 -885 36621
rect -851 36596 -813 36621
rect -779 36596 -741 36621
rect -707 36596 -669 36621
rect -635 36596 -597 36621
rect -563 36596 -525 36621
rect -491 36596 -453 36621
rect -419 36596 -381 36621
rect -347 36596 -309 36621
rect -275 36596 -153 36621
rect -2969 36562 -2938 36596
rect -2904 36562 -2870 36596
rect -2836 36587 -2829 36596
rect -2768 36587 -2757 36596
rect -2700 36587 -2685 36596
rect -2632 36587 -2613 36596
rect -2564 36587 -2541 36596
rect -2496 36587 -2469 36596
rect -2428 36587 -2397 36596
rect -2836 36562 -2802 36587
rect -2768 36562 -2734 36587
rect -2700 36562 -2666 36587
rect -2632 36562 -2598 36587
rect -2564 36562 -2530 36587
rect -2496 36562 -2462 36587
rect -2428 36562 -2394 36587
rect -2360 36562 -2326 36596
rect -2291 36587 -2258 36596
rect -2219 36587 -2190 36596
rect -2147 36587 -2122 36596
rect -2075 36587 -2054 36596
rect -2003 36587 -1986 36596
rect -1931 36587 -1918 36596
rect -1859 36587 -1850 36596
rect -1787 36587 -1782 36596
rect -1715 36587 -1714 36596
rect -2292 36562 -2258 36587
rect -2224 36562 -2190 36587
rect -2156 36562 -2122 36587
rect -2088 36562 -2054 36587
rect -2020 36562 -1986 36587
rect -1952 36562 -1918 36587
rect -1884 36562 -1850 36587
rect -1816 36562 -1782 36587
rect -1748 36562 -1714 36587
rect -1680 36587 -1677 36596
rect -1612 36587 -1605 36596
rect -1544 36587 -1533 36596
rect -1476 36587 -1461 36596
rect -1408 36587 -1389 36596
rect -1340 36587 -1317 36596
rect -1272 36587 -1245 36596
rect -1204 36587 -1173 36596
rect -1680 36562 -1646 36587
rect -1612 36562 -1578 36587
rect -1544 36562 -1510 36587
rect -1476 36562 -1442 36587
rect -1408 36562 -1374 36587
rect -1340 36562 -1306 36587
rect -1272 36562 -1238 36587
rect -1204 36562 -1170 36587
rect -1136 36562 -1102 36596
rect -1067 36587 -1034 36596
rect -995 36587 -966 36596
rect -923 36587 -898 36596
rect -851 36587 -830 36596
rect -779 36587 -762 36596
rect -707 36587 -694 36596
rect -635 36587 -626 36596
rect -563 36587 -558 36596
rect -491 36587 -490 36596
rect -1068 36562 -1034 36587
rect -1000 36562 -966 36587
rect -932 36562 -898 36587
rect -864 36562 -830 36587
rect -796 36562 -762 36587
rect -728 36562 -694 36587
rect -660 36562 -626 36587
rect -592 36562 -558 36587
rect -524 36562 -490 36587
rect -456 36587 -453 36596
rect -388 36587 -381 36596
rect -320 36587 -309 36596
rect -456 36562 -422 36587
rect -388 36562 -354 36587
rect -320 36562 -286 36587
rect -252 36562 -218 36596
rect -184 36562 -153 36596
rect -2969 36548 -153 36562
rect -2969 36527 -2829 36548
rect -2795 36527 -2757 36548
rect -2723 36527 -2685 36548
rect -2651 36527 -2613 36548
rect -2579 36527 -2541 36548
rect -2507 36527 -2469 36548
rect -2435 36527 -2397 36548
rect -2363 36527 -2325 36548
rect -2291 36527 -2253 36548
rect -2219 36527 -2181 36548
rect -2147 36527 -2109 36548
rect -2075 36527 -2037 36548
rect -2003 36527 -1965 36548
rect -1931 36527 -1893 36548
rect -1859 36527 -1821 36548
rect -1787 36527 -1749 36548
rect -1715 36527 -1677 36548
rect -1643 36527 -1605 36548
rect -1571 36527 -1533 36548
rect -1499 36527 -1461 36548
rect -1427 36527 -1389 36548
rect -1355 36527 -1317 36548
rect -1283 36527 -1245 36548
rect -1211 36527 -1173 36548
rect -1139 36527 -1101 36548
rect -1067 36527 -1029 36548
rect -995 36527 -957 36548
rect -923 36527 -885 36548
rect -851 36527 -813 36548
rect -779 36527 -741 36548
rect -707 36527 -669 36548
rect -635 36527 -597 36548
rect -563 36527 -525 36548
rect -491 36527 -453 36548
rect -419 36527 -381 36548
rect -347 36527 -309 36548
rect -275 36527 -153 36548
rect -2969 36493 -2938 36527
rect -2904 36493 -2870 36527
rect -2836 36514 -2829 36527
rect -2768 36514 -2757 36527
rect -2700 36514 -2685 36527
rect -2632 36514 -2613 36527
rect -2564 36514 -2541 36527
rect -2496 36514 -2469 36527
rect -2428 36514 -2397 36527
rect -2836 36493 -2802 36514
rect -2768 36493 -2734 36514
rect -2700 36493 -2666 36514
rect -2632 36493 -2598 36514
rect -2564 36493 -2530 36514
rect -2496 36493 -2462 36514
rect -2428 36493 -2394 36514
rect -2360 36493 -2326 36527
rect -2291 36514 -2258 36527
rect -2219 36514 -2190 36527
rect -2147 36514 -2122 36527
rect -2075 36514 -2054 36527
rect -2003 36514 -1986 36527
rect -1931 36514 -1918 36527
rect -1859 36514 -1850 36527
rect -1787 36514 -1782 36527
rect -1715 36514 -1714 36527
rect -2292 36493 -2258 36514
rect -2224 36493 -2190 36514
rect -2156 36493 -2122 36514
rect -2088 36493 -2054 36514
rect -2020 36493 -1986 36514
rect -1952 36493 -1918 36514
rect -1884 36493 -1850 36514
rect -1816 36493 -1782 36514
rect -1748 36493 -1714 36514
rect -1680 36514 -1677 36527
rect -1612 36514 -1605 36527
rect -1544 36514 -1533 36527
rect -1476 36514 -1461 36527
rect -1408 36514 -1389 36527
rect -1340 36514 -1317 36527
rect -1272 36514 -1245 36527
rect -1204 36514 -1173 36527
rect -1680 36493 -1646 36514
rect -1612 36493 -1578 36514
rect -1544 36493 -1510 36514
rect -1476 36493 -1442 36514
rect -1408 36493 -1374 36514
rect -1340 36493 -1306 36514
rect -1272 36493 -1238 36514
rect -1204 36493 -1170 36514
rect -1136 36493 -1102 36527
rect -1067 36514 -1034 36527
rect -995 36514 -966 36527
rect -923 36514 -898 36527
rect -851 36514 -830 36527
rect -779 36514 -762 36527
rect -707 36514 -694 36527
rect -635 36514 -626 36527
rect -563 36514 -558 36527
rect -491 36514 -490 36527
rect -1068 36493 -1034 36514
rect -1000 36493 -966 36514
rect -932 36493 -898 36514
rect -864 36493 -830 36514
rect -796 36493 -762 36514
rect -728 36493 -694 36514
rect -660 36493 -626 36514
rect -592 36493 -558 36514
rect -524 36493 -490 36514
rect -456 36514 -453 36527
rect -388 36514 -381 36527
rect -320 36514 -309 36527
rect -456 36493 -422 36514
rect -388 36493 -354 36514
rect -320 36493 -286 36514
rect -252 36493 -218 36527
rect -184 36493 -153 36527
rect -2969 36475 -153 36493
rect -2969 36458 -2829 36475
rect -2795 36458 -2757 36475
rect -2723 36458 -2685 36475
rect -2651 36458 -2613 36475
rect -2579 36458 -2541 36475
rect -2507 36458 -2469 36475
rect -2435 36458 -2397 36475
rect -2363 36458 -2325 36475
rect -2291 36458 -2253 36475
rect -2219 36458 -2181 36475
rect -2147 36458 -2109 36475
rect -2075 36458 -2037 36475
rect -2003 36458 -1965 36475
rect -1931 36458 -1893 36475
rect -1859 36458 -1821 36475
rect -1787 36458 -1749 36475
rect -1715 36458 -1677 36475
rect -1643 36458 -1605 36475
rect -1571 36458 -1533 36475
rect -1499 36458 -1461 36475
rect -1427 36458 -1389 36475
rect -1355 36458 -1317 36475
rect -1283 36458 -1245 36475
rect -1211 36458 -1173 36475
rect -1139 36458 -1101 36475
rect -1067 36458 -1029 36475
rect -995 36458 -957 36475
rect -923 36458 -885 36475
rect -851 36458 -813 36475
rect -779 36458 -741 36475
rect -707 36458 -669 36475
rect -635 36458 -597 36475
rect -563 36458 -525 36475
rect -491 36458 -453 36475
rect -419 36458 -381 36475
rect -347 36458 -309 36475
rect -275 36458 -153 36475
rect -2969 36424 -2938 36458
rect -2904 36424 -2870 36458
rect -2836 36441 -2829 36458
rect -2768 36441 -2757 36458
rect -2700 36441 -2685 36458
rect -2632 36441 -2613 36458
rect -2564 36441 -2541 36458
rect -2496 36441 -2469 36458
rect -2428 36441 -2397 36458
rect -2836 36424 -2802 36441
rect -2768 36424 -2734 36441
rect -2700 36424 -2666 36441
rect -2632 36424 -2598 36441
rect -2564 36424 -2530 36441
rect -2496 36424 -2462 36441
rect -2428 36424 -2394 36441
rect -2360 36424 -2326 36458
rect -2291 36441 -2258 36458
rect -2219 36441 -2190 36458
rect -2147 36441 -2122 36458
rect -2075 36441 -2054 36458
rect -2003 36441 -1986 36458
rect -1931 36441 -1918 36458
rect -1859 36441 -1850 36458
rect -1787 36441 -1782 36458
rect -1715 36441 -1714 36458
rect -2292 36424 -2258 36441
rect -2224 36424 -2190 36441
rect -2156 36424 -2122 36441
rect -2088 36424 -2054 36441
rect -2020 36424 -1986 36441
rect -1952 36424 -1918 36441
rect -1884 36424 -1850 36441
rect -1816 36424 -1782 36441
rect -1748 36424 -1714 36441
rect -1680 36441 -1677 36458
rect -1612 36441 -1605 36458
rect -1544 36441 -1533 36458
rect -1476 36441 -1461 36458
rect -1408 36441 -1389 36458
rect -1340 36441 -1317 36458
rect -1272 36441 -1245 36458
rect -1204 36441 -1173 36458
rect -1680 36424 -1646 36441
rect -1612 36424 -1578 36441
rect -1544 36424 -1510 36441
rect -1476 36424 -1442 36441
rect -1408 36424 -1374 36441
rect -1340 36424 -1306 36441
rect -1272 36424 -1238 36441
rect -1204 36424 -1170 36441
rect -1136 36424 -1102 36458
rect -1067 36441 -1034 36458
rect -995 36441 -966 36458
rect -923 36441 -898 36458
rect -851 36441 -830 36458
rect -779 36441 -762 36458
rect -707 36441 -694 36458
rect -635 36441 -626 36458
rect -563 36441 -558 36458
rect -491 36441 -490 36458
rect -1068 36424 -1034 36441
rect -1000 36424 -966 36441
rect -932 36424 -898 36441
rect -864 36424 -830 36441
rect -796 36424 -762 36441
rect -728 36424 -694 36441
rect -660 36424 -626 36441
rect -592 36424 -558 36441
rect -524 36424 -490 36441
rect -456 36441 -453 36458
rect -388 36441 -381 36458
rect -320 36441 -309 36458
rect -456 36424 -422 36441
rect -388 36424 -354 36441
rect -320 36424 -286 36441
rect -252 36424 -218 36458
rect -184 36424 -153 36458
rect -2969 36402 -153 36424
rect -2969 36389 -2829 36402
rect -2795 36389 -2757 36402
rect -2723 36389 -2685 36402
rect -2651 36389 -2613 36402
rect -2579 36389 -2541 36402
rect -2507 36389 -2469 36402
rect -2435 36389 -2397 36402
rect -2363 36389 -2325 36402
rect -2291 36389 -2253 36402
rect -2219 36389 -2181 36402
rect -2147 36389 -2109 36402
rect -2075 36389 -2037 36402
rect -2003 36389 -1965 36402
rect -1931 36389 -1893 36402
rect -1859 36389 -1821 36402
rect -1787 36389 -1749 36402
rect -1715 36389 -1677 36402
rect -1643 36389 -1605 36402
rect -1571 36389 -1533 36402
rect -1499 36389 -1461 36402
rect -1427 36389 -1389 36402
rect -1355 36389 -1317 36402
rect -1283 36389 -1245 36402
rect -1211 36389 -1173 36402
rect -1139 36389 -1101 36402
rect -1067 36389 -1029 36402
rect -995 36389 -957 36402
rect -923 36389 -885 36402
rect -851 36389 -813 36402
rect -779 36389 -741 36402
rect -707 36389 -669 36402
rect -635 36389 -597 36402
rect -563 36389 -525 36402
rect -491 36389 -453 36402
rect -419 36389 -381 36402
rect -347 36389 -309 36402
rect -275 36389 -153 36402
rect -2969 36355 -2938 36389
rect -2904 36355 -2870 36389
rect -2836 36368 -2829 36389
rect -2768 36368 -2757 36389
rect -2700 36368 -2685 36389
rect -2632 36368 -2613 36389
rect -2564 36368 -2541 36389
rect -2496 36368 -2469 36389
rect -2428 36368 -2397 36389
rect -2836 36355 -2802 36368
rect -2768 36355 -2734 36368
rect -2700 36355 -2666 36368
rect -2632 36355 -2598 36368
rect -2564 36355 -2530 36368
rect -2496 36355 -2462 36368
rect -2428 36355 -2394 36368
rect -2360 36355 -2326 36389
rect -2291 36368 -2258 36389
rect -2219 36368 -2190 36389
rect -2147 36368 -2122 36389
rect -2075 36368 -2054 36389
rect -2003 36368 -1986 36389
rect -1931 36368 -1918 36389
rect -1859 36368 -1850 36389
rect -1787 36368 -1782 36389
rect -1715 36368 -1714 36389
rect -2292 36355 -2258 36368
rect -2224 36355 -2190 36368
rect -2156 36355 -2122 36368
rect -2088 36355 -2054 36368
rect -2020 36355 -1986 36368
rect -1952 36355 -1918 36368
rect -1884 36355 -1850 36368
rect -1816 36355 -1782 36368
rect -1748 36355 -1714 36368
rect -1680 36368 -1677 36389
rect -1612 36368 -1605 36389
rect -1544 36368 -1533 36389
rect -1476 36368 -1461 36389
rect -1408 36368 -1389 36389
rect -1340 36368 -1317 36389
rect -1272 36368 -1245 36389
rect -1204 36368 -1173 36389
rect -1680 36355 -1646 36368
rect -1612 36355 -1578 36368
rect -1544 36355 -1510 36368
rect -1476 36355 -1442 36368
rect -1408 36355 -1374 36368
rect -1340 36355 -1306 36368
rect -1272 36355 -1238 36368
rect -1204 36355 -1170 36368
rect -1136 36355 -1102 36389
rect -1067 36368 -1034 36389
rect -995 36368 -966 36389
rect -923 36368 -898 36389
rect -851 36368 -830 36389
rect -779 36368 -762 36389
rect -707 36368 -694 36389
rect -635 36368 -626 36389
rect -563 36368 -558 36389
rect -491 36368 -490 36389
rect -1068 36355 -1034 36368
rect -1000 36355 -966 36368
rect -932 36355 -898 36368
rect -864 36355 -830 36368
rect -796 36355 -762 36368
rect -728 36355 -694 36368
rect -660 36355 -626 36368
rect -592 36355 -558 36368
rect -524 36355 -490 36368
rect -456 36368 -453 36389
rect -388 36368 -381 36389
rect -320 36368 -309 36389
rect -456 36355 -422 36368
rect -388 36355 -354 36368
rect -320 36355 -286 36368
rect -252 36355 -218 36389
rect -184 36355 -153 36389
rect -2969 36329 -153 36355
rect -2969 36320 -2829 36329
rect -2795 36320 -2757 36329
rect -2723 36320 -2685 36329
rect -2651 36320 -2613 36329
rect -2579 36320 -2541 36329
rect -2507 36320 -2469 36329
rect -2435 36320 -2397 36329
rect -2363 36320 -2325 36329
rect -2291 36320 -2253 36329
rect -2219 36320 -2181 36329
rect -2147 36320 -2109 36329
rect -2075 36320 -2037 36329
rect -2003 36320 -1965 36329
rect -1931 36320 -1893 36329
rect -1859 36320 -1821 36329
rect -1787 36320 -1749 36329
rect -1715 36320 -1677 36329
rect -1643 36320 -1605 36329
rect -1571 36320 -1533 36329
rect -1499 36320 -1461 36329
rect -1427 36320 -1389 36329
rect -1355 36320 -1317 36329
rect -1283 36320 -1245 36329
rect -1211 36320 -1173 36329
rect -1139 36320 -1101 36329
rect -1067 36320 -1029 36329
rect -995 36320 -957 36329
rect -923 36320 -885 36329
rect -851 36320 -813 36329
rect -779 36320 -741 36329
rect -707 36320 -669 36329
rect -635 36320 -597 36329
rect -563 36320 -525 36329
rect -491 36320 -453 36329
rect -419 36320 -381 36329
rect -347 36320 -309 36329
rect -275 36320 -153 36329
rect -2969 36286 -2938 36320
rect -2904 36286 -2870 36320
rect -2836 36295 -2829 36320
rect -2768 36295 -2757 36320
rect -2700 36295 -2685 36320
rect -2632 36295 -2613 36320
rect -2564 36295 -2541 36320
rect -2496 36295 -2469 36320
rect -2428 36295 -2397 36320
rect -2836 36286 -2802 36295
rect -2768 36286 -2734 36295
rect -2700 36286 -2666 36295
rect -2632 36286 -2598 36295
rect -2564 36286 -2530 36295
rect -2496 36286 -2462 36295
rect -2428 36286 -2394 36295
rect -2360 36286 -2326 36320
rect -2291 36295 -2258 36320
rect -2219 36295 -2190 36320
rect -2147 36295 -2122 36320
rect -2075 36295 -2054 36320
rect -2003 36295 -1986 36320
rect -1931 36295 -1918 36320
rect -1859 36295 -1850 36320
rect -1787 36295 -1782 36320
rect -1715 36295 -1714 36320
rect -2292 36286 -2258 36295
rect -2224 36286 -2190 36295
rect -2156 36286 -2122 36295
rect -2088 36286 -2054 36295
rect -2020 36286 -1986 36295
rect -1952 36286 -1918 36295
rect -1884 36286 -1850 36295
rect -1816 36286 -1782 36295
rect -1748 36286 -1714 36295
rect -1680 36295 -1677 36320
rect -1612 36295 -1605 36320
rect -1544 36295 -1533 36320
rect -1476 36295 -1461 36320
rect -1408 36295 -1389 36320
rect -1340 36295 -1317 36320
rect -1272 36295 -1245 36320
rect -1204 36295 -1173 36320
rect -1680 36286 -1646 36295
rect -1612 36286 -1578 36295
rect -1544 36286 -1510 36295
rect -1476 36286 -1442 36295
rect -1408 36286 -1374 36295
rect -1340 36286 -1306 36295
rect -1272 36286 -1238 36295
rect -1204 36286 -1170 36295
rect -1136 36286 -1102 36320
rect -1067 36295 -1034 36320
rect -995 36295 -966 36320
rect -923 36295 -898 36320
rect -851 36295 -830 36320
rect -779 36295 -762 36320
rect -707 36295 -694 36320
rect -635 36295 -626 36320
rect -563 36295 -558 36320
rect -491 36295 -490 36320
rect -1068 36286 -1034 36295
rect -1000 36286 -966 36295
rect -932 36286 -898 36295
rect -864 36286 -830 36295
rect -796 36286 -762 36295
rect -728 36286 -694 36295
rect -660 36286 -626 36295
rect -592 36286 -558 36295
rect -524 36286 -490 36295
rect -456 36295 -453 36320
rect -388 36295 -381 36320
rect -320 36295 -309 36320
rect -456 36286 -422 36295
rect -388 36286 -354 36295
rect -320 36286 -286 36295
rect -252 36286 -218 36320
rect -184 36286 -153 36320
rect -2969 36256 -153 36286
rect -2969 36251 -2829 36256
rect -2795 36251 -2757 36256
rect -2723 36251 -2685 36256
rect -2651 36251 -2613 36256
rect -2579 36251 -2541 36256
rect -2507 36251 -2469 36256
rect -2435 36251 -2397 36256
rect -2363 36251 -2325 36256
rect -2291 36251 -2253 36256
rect -2219 36251 -2181 36256
rect -2147 36251 -2109 36256
rect -2075 36251 -2037 36256
rect -2003 36251 -1965 36256
rect -1931 36251 -1893 36256
rect -1859 36251 -1821 36256
rect -1787 36251 -1749 36256
rect -1715 36251 -1677 36256
rect -1643 36251 -1605 36256
rect -1571 36251 -1533 36256
rect -1499 36251 -1461 36256
rect -1427 36251 -1389 36256
rect -1355 36251 -1317 36256
rect -1283 36251 -1245 36256
rect -1211 36251 -1173 36256
rect -1139 36251 -1101 36256
rect -1067 36251 -1029 36256
rect -995 36251 -957 36256
rect -923 36251 -885 36256
rect -851 36251 -813 36256
rect -779 36251 -741 36256
rect -707 36251 -669 36256
rect -635 36251 -597 36256
rect -563 36251 -525 36256
rect -491 36251 -453 36256
rect -419 36251 -381 36256
rect -347 36251 -309 36256
rect -275 36251 -153 36256
rect -2969 36217 -2938 36251
rect -2904 36217 -2870 36251
rect -2836 36222 -2829 36251
rect -2768 36222 -2757 36251
rect -2700 36222 -2685 36251
rect -2632 36222 -2613 36251
rect -2564 36222 -2541 36251
rect -2496 36222 -2469 36251
rect -2428 36222 -2397 36251
rect -2836 36217 -2802 36222
rect -2768 36217 -2734 36222
rect -2700 36217 -2666 36222
rect -2632 36217 -2598 36222
rect -2564 36217 -2530 36222
rect -2496 36217 -2462 36222
rect -2428 36217 -2394 36222
rect -2360 36217 -2326 36251
rect -2291 36222 -2258 36251
rect -2219 36222 -2190 36251
rect -2147 36222 -2122 36251
rect -2075 36222 -2054 36251
rect -2003 36222 -1986 36251
rect -1931 36222 -1918 36251
rect -1859 36222 -1850 36251
rect -1787 36222 -1782 36251
rect -1715 36222 -1714 36251
rect -2292 36217 -2258 36222
rect -2224 36217 -2190 36222
rect -2156 36217 -2122 36222
rect -2088 36217 -2054 36222
rect -2020 36217 -1986 36222
rect -1952 36217 -1918 36222
rect -1884 36217 -1850 36222
rect -1816 36217 -1782 36222
rect -1748 36217 -1714 36222
rect -1680 36222 -1677 36251
rect -1612 36222 -1605 36251
rect -1544 36222 -1533 36251
rect -1476 36222 -1461 36251
rect -1408 36222 -1389 36251
rect -1340 36222 -1317 36251
rect -1272 36222 -1245 36251
rect -1204 36222 -1173 36251
rect -1680 36217 -1646 36222
rect -1612 36217 -1578 36222
rect -1544 36217 -1510 36222
rect -1476 36217 -1442 36222
rect -1408 36217 -1374 36222
rect -1340 36217 -1306 36222
rect -1272 36217 -1238 36222
rect -1204 36217 -1170 36222
rect -1136 36217 -1102 36251
rect -1067 36222 -1034 36251
rect -995 36222 -966 36251
rect -923 36222 -898 36251
rect -851 36222 -830 36251
rect -779 36222 -762 36251
rect -707 36222 -694 36251
rect -635 36222 -626 36251
rect -563 36222 -558 36251
rect -491 36222 -490 36251
rect -1068 36217 -1034 36222
rect -1000 36217 -966 36222
rect -932 36217 -898 36222
rect -864 36217 -830 36222
rect -796 36217 -762 36222
rect -728 36217 -694 36222
rect -660 36217 -626 36222
rect -592 36217 -558 36222
rect -524 36217 -490 36222
rect -456 36222 -453 36251
rect -388 36222 -381 36251
rect -320 36222 -309 36251
rect -456 36217 -422 36222
rect -388 36217 -354 36222
rect -320 36217 -286 36222
rect -252 36217 -218 36251
rect -184 36217 -153 36251
rect -2969 36183 -153 36217
rect -2969 36182 -2829 36183
rect -2795 36182 -2757 36183
rect -2723 36182 -2685 36183
rect -2651 36182 -2613 36183
rect -2579 36182 -2541 36183
rect -2507 36182 -2469 36183
rect -2435 36182 -2397 36183
rect -2363 36182 -2325 36183
rect -2291 36182 -2253 36183
rect -2219 36182 -2181 36183
rect -2147 36182 -2109 36183
rect -2075 36182 -2037 36183
rect -2003 36182 -1965 36183
rect -1931 36182 -1893 36183
rect -1859 36182 -1821 36183
rect -1787 36182 -1749 36183
rect -1715 36182 -1677 36183
rect -1643 36182 -1605 36183
rect -1571 36182 -1533 36183
rect -1499 36182 -1461 36183
rect -1427 36182 -1389 36183
rect -1355 36182 -1317 36183
rect -1283 36182 -1245 36183
rect -1211 36182 -1173 36183
rect -1139 36182 -1101 36183
rect -1067 36182 -1029 36183
rect -995 36182 -957 36183
rect -923 36182 -885 36183
rect -851 36182 -813 36183
rect -779 36182 -741 36183
rect -707 36182 -669 36183
rect -635 36182 -597 36183
rect -563 36182 -525 36183
rect -491 36182 -453 36183
rect -419 36182 -381 36183
rect -347 36182 -309 36183
rect -275 36182 -153 36183
rect -2969 36148 -2938 36182
rect -2904 36148 -2870 36182
rect -2836 36149 -2829 36182
rect -2768 36149 -2757 36182
rect -2700 36149 -2685 36182
rect -2632 36149 -2613 36182
rect -2564 36149 -2541 36182
rect -2496 36149 -2469 36182
rect -2428 36149 -2397 36182
rect -2836 36148 -2802 36149
rect -2768 36148 -2734 36149
rect -2700 36148 -2666 36149
rect -2632 36148 -2598 36149
rect -2564 36148 -2530 36149
rect -2496 36148 -2462 36149
rect -2428 36148 -2394 36149
rect -2360 36148 -2326 36182
rect -2291 36149 -2258 36182
rect -2219 36149 -2190 36182
rect -2147 36149 -2122 36182
rect -2075 36149 -2054 36182
rect -2003 36149 -1986 36182
rect -1931 36149 -1918 36182
rect -1859 36149 -1850 36182
rect -1787 36149 -1782 36182
rect -1715 36149 -1714 36182
rect -2292 36148 -2258 36149
rect -2224 36148 -2190 36149
rect -2156 36148 -2122 36149
rect -2088 36148 -2054 36149
rect -2020 36148 -1986 36149
rect -1952 36148 -1918 36149
rect -1884 36148 -1850 36149
rect -1816 36148 -1782 36149
rect -1748 36148 -1714 36149
rect -1680 36149 -1677 36182
rect -1612 36149 -1605 36182
rect -1544 36149 -1533 36182
rect -1476 36149 -1461 36182
rect -1408 36149 -1389 36182
rect -1340 36149 -1317 36182
rect -1272 36149 -1245 36182
rect -1204 36149 -1173 36182
rect -1680 36148 -1646 36149
rect -1612 36148 -1578 36149
rect -1544 36148 -1510 36149
rect -1476 36148 -1442 36149
rect -1408 36148 -1374 36149
rect -1340 36148 -1306 36149
rect -1272 36148 -1238 36149
rect -1204 36148 -1170 36149
rect -1136 36148 -1102 36182
rect -1067 36149 -1034 36182
rect -995 36149 -966 36182
rect -923 36149 -898 36182
rect -851 36149 -830 36182
rect -779 36149 -762 36182
rect -707 36149 -694 36182
rect -635 36149 -626 36182
rect -563 36149 -558 36182
rect -491 36149 -490 36182
rect -1068 36148 -1034 36149
rect -1000 36148 -966 36149
rect -932 36148 -898 36149
rect -864 36148 -830 36149
rect -796 36148 -762 36149
rect -728 36148 -694 36149
rect -660 36148 -626 36149
rect -592 36148 -558 36149
rect -524 36148 -490 36149
rect -456 36149 -453 36182
rect -388 36149 -381 36182
rect -320 36149 -309 36182
rect -456 36148 -422 36149
rect -388 36148 -354 36149
rect -320 36148 -286 36149
rect -252 36148 -218 36182
rect -184 36148 -153 36182
rect -2969 36113 -153 36148
rect -2969 36079 -2938 36113
rect -2904 36079 -2870 36113
rect -2836 36110 -2802 36113
rect -2768 36110 -2734 36113
rect -2700 36110 -2666 36113
rect -2632 36110 -2598 36113
rect -2564 36110 -2530 36113
rect -2496 36110 -2462 36113
rect -2428 36110 -2394 36113
rect -2836 36079 -2829 36110
rect -2768 36079 -2757 36110
rect -2700 36079 -2685 36110
rect -2632 36079 -2613 36110
rect -2564 36079 -2541 36110
rect -2496 36079 -2469 36110
rect -2428 36079 -2397 36110
rect -2360 36079 -2326 36113
rect -2292 36110 -2258 36113
rect -2224 36110 -2190 36113
rect -2156 36110 -2122 36113
rect -2088 36110 -2054 36113
rect -2020 36110 -1986 36113
rect -1952 36110 -1918 36113
rect -1884 36110 -1850 36113
rect -1816 36110 -1782 36113
rect -1748 36110 -1714 36113
rect -2291 36079 -2258 36110
rect -2219 36079 -2190 36110
rect -2147 36079 -2122 36110
rect -2075 36079 -2054 36110
rect -2003 36079 -1986 36110
rect -1931 36079 -1918 36110
rect -1859 36079 -1850 36110
rect -1787 36079 -1782 36110
rect -1715 36079 -1714 36110
rect -1680 36110 -1646 36113
rect -1612 36110 -1578 36113
rect -1544 36110 -1510 36113
rect -1476 36110 -1442 36113
rect -1408 36110 -1374 36113
rect -1340 36110 -1306 36113
rect -1272 36110 -1238 36113
rect -1204 36110 -1170 36113
rect -1680 36079 -1677 36110
rect -1612 36079 -1605 36110
rect -1544 36079 -1533 36110
rect -1476 36079 -1461 36110
rect -1408 36079 -1389 36110
rect -1340 36079 -1317 36110
rect -1272 36079 -1245 36110
rect -1204 36079 -1173 36110
rect -1136 36079 -1102 36113
rect -1068 36110 -1034 36113
rect -1000 36110 -966 36113
rect -932 36110 -898 36113
rect -864 36110 -830 36113
rect -796 36110 -762 36113
rect -728 36110 -694 36113
rect -660 36110 -626 36113
rect -592 36110 -558 36113
rect -524 36110 -490 36113
rect -1067 36079 -1034 36110
rect -995 36079 -966 36110
rect -923 36079 -898 36110
rect -851 36079 -830 36110
rect -779 36079 -762 36110
rect -707 36079 -694 36110
rect -635 36079 -626 36110
rect -563 36079 -558 36110
rect -491 36079 -490 36110
rect -456 36110 -422 36113
rect -388 36110 -354 36113
rect -320 36110 -286 36113
rect -456 36079 -453 36110
rect -388 36079 -381 36110
rect -320 36079 -309 36110
rect -252 36079 -218 36113
rect -184 36079 -153 36113
rect -2969 36076 -2829 36079
rect -2795 36076 -2757 36079
rect -2723 36076 -2685 36079
rect -2651 36076 -2613 36079
rect -2579 36076 -2541 36079
rect -2507 36076 -2469 36079
rect -2435 36076 -2397 36079
rect -2363 36076 -2325 36079
rect -2291 36076 -2253 36079
rect -2219 36076 -2181 36079
rect -2147 36076 -2109 36079
rect -2075 36076 -2037 36079
rect -2003 36076 -1965 36079
rect -1931 36076 -1893 36079
rect -1859 36076 -1821 36079
rect -1787 36076 -1749 36079
rect -1715 36076 -1677 36079
rect -1643 36076 -1605 36079
rect -1571 36076 -1533 36079
rect -1499 36076 -1461 36079
rect -1427 36076 -1389 36079
rect -1355 36076 -1317 36079
rect -1283 36076 -1245 36079
rect -1211 36076 -1173 36079
rect -1139 36076 -1101 36079
rect -1067 36076 -1029 36079
rect -995 36076 -957 36079
rect -923 36076 -885 36079
rect -851 36076 -813 36079
rect -779 36076 -741 36079
rect -707 36076 -669 36079
rect -635 36076 -597 36079
rect -563 36076 -525 36079
rect -491 36076 -453 36079
rect -419 36076 -381 36079
rect -347 36076 -309 36079
rect -275 36076 -153 36079
rect -2969 36044 -153 36076
rect -2969 36010 -2938 36044
rect -2904 36010 -2870 36044
rect -2836 36037 -2802 36044
rect -2768 36037 -2734 36044
rect -2700 36037 -2666 36044
rect -2632 36037 -2598 36044
rect -2564 36037 -2530 36044
rect -2496 36037 -2462 36044
rect -2428 36037 -2394 36044
rect -2836 36010 -2829 36037
rect -2768 36010 -2757 36037
rect -2700 36010 -2685 36037
rect -2632 36010 -2613 36037
rect -2564 36010 -2541 36037
rect -2496 36010 -2469 36037
rect -2428 36010 -2397 36037
rect -2360 36010 -2326 36044
rect -2292 36037 -2258 36044
rect -2224 36037 -2190 36044
rect -2156 36037 -2122 36044
rect -2088 36037 -2054 36044
rect -2020 36037 -1986 36044
rect -1952 36037 -1918 36044
rect -1884 36037 -1850 36044
rect -1816 36037 -1782 36044
rect -1748 36037 -1714 36044
rect -2291 36010 -2258 36037
rect -2219 36010 -2190 36037
rect -2147 36010 -2122 36037
rect -2075 36010 -2054 36037
rect -2003 36010 -1986 36037
rect -1931 36010 -1918 36037
rect -1859 36010 -1850 36037
rect -1787 36010 -1782 36037
rect -1715 36010 -1714 36037
rect -1680 36037 -1646 36044
rect -1612 36037 -1578 36044
rect -1544 36037 -1510 36044
rect -1476 36037 -1442 36044
rect -1408 36037 -1374 36044
rect -1340 36037 -1306 36044
rect -1272 36037 -1238 36044
rect -1204 36037 -1170 36044
rect -1680 36010 -1677 36037
rect -1612 36010 -1605 36037
rect -1544 36010 -1533 36037
rect -1476 36010 -1461 36037
rect -1408 36010 -1389 36037
rect -1340 36010 -1317 36037
rect -1272 36010 -1245 36037
rect -1204 36010 -1173 36037
rect -1136 36010 -1102 36044
rect -1068 36037 -1034 36044
rect -1000 36037 -966 36044
rect -932 36037 -898 36044
rect -864 36037 -830 36044
rect -796 36037 -762 36044
rect -728 36037 -694 36044
rect -660 36037 -626 36044
rect -592 36037 -558 36044
rect -524 36037 -490 36044
rect -1067 36010 -1034 36037
rect -995 36010 -966 36037
rect -923 36010 -898 36037
rect -851 36010 -830 36037
rect -779 36010 -762 36037
rect -707 36010 -694 36037
rect -635 36010 -626 36037
rect -563 36010 -558 36037
rect -491 36010 -490 36037
rect -456 36037 -422 36044
rect -388 36037 -354 36044
rect -320 36037 -286 36044
rect -456 36010 -453 36037
rect -388 36010 -381 36037
rect -320 36010 -309 36037
rect -252 36010 -218 36044
rect -184 36010 -153 36044
rect -2969 36003 -2829 36010
rect -2795 36003 -2757 36010
rect -2723 36003 -2685 36010
rect -2651 36003 -2613 36010
rect -2579 36003 -2541 36010
rect -2507 36003 -2469 36010
rect -2435 36003 -2397 36010
rect -2363 36003 -2325 36010
rect -2291 36003 -2253 36010
rect -2219 36003 -2181 36010
rect -2147 36003 -2109 36010
rect -2075 36003 -2037 36010
rect -2003 36003 -1965 36010
rect -1931 36003 -1893 36010
rect -1859 36003 -1821 36010
rect -1787 36003 -1749 36010
rect -1715 36003 -1677 36010
rect -1643 36003 -1605 36010
rect -1571 36003 -1533 36010
rect -1499 36003 -1461 36010
rect -1427 36003 -1389 36010
rect -1355 36003 -1317 36010
rect -1283 36003 -1245 36010
rect -1211 36003 -1173 36010
rect -1139 36003 -1101 36010
rect -1067 36003 -1029 36010
rect -995 36003 -957 36010
rect -923 36003 -885 36010
rect -851 36003 -813 36010
rect -779 36003 -741 36010
rect -707 36003 -669 36010
rect -635 36003 -597 36010
rect -563 36003 -525 36010
rect -491 36003 -453 36010
rect -419 36003 -381 36010
rect -347 36003 -309 36010
rect -275 36003 -153 36010
rect -2969 35975 -153 36003
rect -2969 35941 -2938 35975
rect -2904 35941 -2870 35975
rect -2836 35964 -2802 35975
rect -2768 35964 -2734 35975
rect -2700 35964 -2666 35975
rect -2632 35964 -2598 35975
rect -2564 35964 -2530 35975
rect -2496 35964 -2462 35975
rect -2428 35964 -2394 35975
rect -2836 35941 -2829 35964
rect -2768 35941 -2757 35964
rect -2700 35941 -2685 35964
rect -2632 35941 -2613 35964
rect -2564 35941 -2541 35964
rect -2496 35941 -2469 35964
rect -2428 35941 -2397 35964
rect -2360 35941 -2326 35975
rect -2292 35964 -2258 35975
rect -2224 35964 -2190 35975
rect -2156 35964 -2122 35975
rect -2088 35964 -2054 35975
rect -2020 35964 -1986 35975
rect -1952 35964 -1918 35975
rect -1884 35964 -1850 35975
rect -1816 35964 -1782 35975
rect -1748 35964 -1714 35975
rect -2291 35941 -2258 35964
rect -2219 35941 -2190 35964
rect -2147 35941 -2122 35964
rect -2075 35941 -2054 35964
rect -2003 35941 -1986 35964
rect -1931 35941 -1918 35964
rect -1859 35941 -1850 35964
rect -1787 35941 -1782 35964
rect -1715 35941 -1714 35964
rect -1680 35964 -1646 35975
rect -1612 35964 -1578 35975
rect -1544 35964 -1510 35975
rect -1476 35964 -1442 35975
rect -1408 35964 -1374 35975
rect -1340 35964 -1306 35975
rect -1272 35964 -1238 35975
rect -1204 35964 -1170 35975
rect -1680 35941 -1677 35964
rect -1612 35941 -1605 35964
rect -1544 35941 -1533 35964
rect -1476 35941 -1461 35964
rect -1408 35941 -1389 35964
rect -1340 35941 -1317 35964
rect -1272 35941 -1245 35964
rect -1204 35941 -1173 35964
rect -1136 35941 -1102 35975
rect -1068 35964 -1034 35975
rect -1000 35964 -966 35975
rect -932 35964 -898 35975
rect -864 35964 -830 35975
rect -796 35964 -762 35975
rect -728 35964 -694 35975
rect -660 35964 -626 35975
rect -592 35964 -558 35975
rect -524 35964 -490 35975
rect -1067 35941 -1034 35964
rect -995 35941 -966 35964
rect -923 35941 -898 35964
rect -851 35941 -830 35964
rect -779 35941 -762 35964
rect -707 35941 -694 35964
rect -635 35941 -626 35964
rect -563 35941 -558 35964
rect -491 35941 -490 35964
rect -456 35964 -422 35975
rect -388 35964 -354 35975
rect -320 35964 -286 35975
rect -456 35941 -453 35964
rect -388 35941 -381 35964
rect -320 35941 -309 35964
rect -252 35941 -218 35975
rect -184 35941 -153 35975
rect -2969 35930 -2829 35941
rect -2795 35930 -2757 35941
rect -2723 35930 -2685 35941
rect -2651 35930 -2613 35941
rect -2579 35930 -2541 35941
rect -2507 35930 -2469 35941
rect -2435 35930 -2397 35941
rect -2363 35930 -2325 35941
rect -2291 35930 -2253 35941
rect -2219 35930 -2181 35941
rect -2147 35930 -2109 35941
rect -2075 35930 -2037 35941
rect -2003 35930 -1965 35941
rect -1931 35930 -1893 35941
rect -1859 35930 -1821 35941
rect -1787 35930 -1749 35941
rect -1715 35930 -1677 35941
rect -1643 35930 -1605 35941
rect -1571 35930 -1533 35941
rect -1499 35930 -1461 35941
rect -1427 35930 -1389 35941
rect -1355 35930 -1317 35941
rect -1283 35930 -1245 35941
rect -1211 35930 -1173 35941
rect -1139 35930 -1101 35941
rect -1067 35930 -1029 35941
rect -995 35930 -957 35941
rect -923 35930 -885 35941
rect -851 35930 -813 35941
rect -779 35930 -741 35941
rect -707 35930 -669 35941
rect -635 35930 -597 35941
rect -563 35930 -525 35941
rect -491 35930 -453 35941
rect -419 35930 -381 35941
rect -347 35930 -309 35941
rect -275 35930 -153 35941
rect -2969 35906 -153 35930
rect -2969 35872 -2938 35906
rect -2904 35872 -2870 35906
rect -2836 35891 -2802 35906
rect -2768 35891 -2734 35906
rect -2700 35891 -2666 35906
rect -2632 35891 -2598 35906
rect -2564 35891 -2530 35906
rect -2496 35891 -2462 35906
rect -2428 35891 -2394 35906
rect -2836 35872 -2829 35891
rect -2768 35872 -2757 35891
rect -2700 35872 -2685 35891
rect -2632 35872 -2613 35891
rect -2564 35872 -2541 35891
rect -2496 35872 -2469 35891
rect -2428 35872 -2397 35891
rect -2360 35872 -2326 35906
rect -2292 35891 -2258 35906
rect -2224 35891 -2190 35906
rect -2156 35891 -2122 35906
rect -2088 35891 -2054 35906
rect -2020 35891 -1986 35906
rect -1952 35891 -1918 35906
rect -1884 35891 -1850 35906
rect -1816 35891 -1782 35906
rect -1748 35891 -1714 35906
rect -2291 35872 -2258 35891
rect -2219 35872 -2190 35891
rect -2147 35872 -2122 35891
rect -2075 35872 -2054 35891
rect -2003 35872 -1986 35891
rect -1931 35872 -1918 35891
rect -1859 35872 -1850 35891
rect -1787 35872 -1782 35891
rect -1715 35872 -1714 35891
rect -1680 35891 -1646 35906
rect -1612 35891 -1578 35906
rect -1544 35891 -1510 35906
rect -1476 35891 -1442 35906
rect -1408 35891 -1374 35906
rect -1340 35891 -1306 35906
rect -1272 35891 -1238 35906
rect -1204 35891 -1170 35906
rect -1680 35872 -1677 35891
rect -1612 35872 -1605 35891
rect -1544 35872 -1533 35891
rect -1476 35872 -1461 35891
rect -1408 35872 -1389 35891
rect -1340 35872 -1317 35891
rect -1272 35872 -1245 35891
rect -1204 35872 -1173 35891
rect -1136 35872 -1102 35906
rect -1068 35891 -1034 35906
rect -1000 35891 -966 35906
rect -932 35891 -898 35906
rect -864 35891 -830 35906
rect -796 35891 -762 35906
rect -728 35891 -694 35906
rect -660 35891 -626 35906
rect -592 35891 -558 35906
rect -524 35891 -490 35906
rect -1067 35872 -1034 35891
rect -995 35872 -966 35891
rect -923 35872 -898 35891
rect -851 35872 -830 35891
rect -779 35872 -762 35891
rect -707 35872 -694 35891
rect -635 35872 -626 35891
rect -563 35872 -558 35891
rect -491 35872 -490 35891
rect -456 35891 -422 35906
rect -388 35891 -354 35906
rect -320 35891 -286 35906
rect -456 35872 -453 35891
rect -388 35872 -381 35891
rect -320 35872 -309 35891
rect -252 35872 -218 35906
rect -184 35872 -153 35906
rect -2969 35857 -2829 35872
rect -2795 35857 -2757 35872
rect -2723 35857 -2685 35872
rect -2651 35857 -2613 35872
rect -2579 35857 -2541 35872
rect -2507 35857 -2469 35872
rect -2435 35857 -2397 35872
rect -2363 35857 -2325 35872
rect -2291 35857 -2253 35872
rect -2219 35857 -2181 35872
rect -2147 35857 -2109 35872
rect -2075 35857 -2037 35872
rect -2003 35857 -1965 35872
rect -1931 35857 -1893 35872
rect -1859 35857 -1821 35872
rect -1787 35857 -1749 35872
rect -1715 35857 -1677 35872
rect -1643 35857 -1605 35872
rect -1571 35857 -1533 35872
rect -1499 35857 -1461 35872
rect -1427 35857 -1389 35872
rect -1355 35857 -1317 35872
rect -1283 35857 -1245 35872
rect -1211 35857 -1173 35872
rect -1139 35857 -1101 35872
rect -1067 35857 -1029 35872
rect -995 35857 -957 35872
rect -923 35857 -885 35872
rect -851 35857 -813 35872
rect -779 35857 -741 35872
rect -707 35857 -669 35872
rect -635 35857 -597 35872
rect -563 35857 -525 35872
rect -491 35857 -453 35872
rect -419 35857 -381 35872
rect -347 35857 -309 35872
rect -275 35857 -153 35872
rect -2969 35837 -153 35857
rect -2969 35803 -2938 35837
rect -2904 35803 -2870 35837
rect -2836 35818 -2802 35837
rect -2768 35818 -2734 35837
rect -2700 35818 -2666 35837
rect -2632 35818 -2598 35837
rect -2564 35818 -2530 35837
rect -2496 35818 -2462 35837
rect -2428 35818 -2394 35837
rect -2836 35803 -2829 35818
rect -2768 35803 -2757 35818
rect -2700 35803 -2685 35818
rect -2632 35803 -2613 35818
rect -2564 35803 -2541 35818
rect -2496 35803 -2469 35818
rect -2428 35803 -2397 35818
rect -2360 35803 -2326 35837
rect -2292 35818 -2258 35837
rect -2224 35818 -2190 35837
rect -2156 35818 -2122 35837
rect -2088 35818 -2054 35837
rect -2020 35818 -1986 35837
rect -1952 35818 -1918 35837
rect -1884 35818 -1850 35837
rect -1816 35818 -1782 35837
rect -1748 35818 -1714 35837
rect -2291 35803 -2258 35818
rect -2219 35803 -2190 35818
rect -2147 35803 -2122 35818
rect -2075 35803 -2054 35818
rect -2003 35803 -1986 35818
rect -1931 35803 -1918 35818
rect -1859 35803 -1850 35818
rect -1787 35803 -1782 35818
rect -1715 35803 -1714 35818
rect -1680 35818 -1646 35837
rect -1612 35818 -1578 35837
rect -1544 35818 -1510 35837
rect -1476 35818 -1442 35837
rect -1408 35818 -1374 35837
rect -1340 35818 -1306 35837
rect -1272 35818 -1238 35837
rect -1204 35818 -1170 35837
rect -1680 35803 -1677 35818
rect -1612 35803 -1605 35818
rect -1544 35803 -1533 35818
rect -1476 35803 -1461 35818
rect -1408 35803 -1389 35818
rect -1340 35803 -1317 35818
rect -1272 35803 -1245 35818
rect -1204 35803 -1173 35818
rect -1136 35803 -1102 35837
rect -1068 35818 -1034 35837
rect -1000 35818 -966 35837
rect -932 35818 -898 35837
rect -864 35818 -830 35837
rect -796 35818 -762 35837
rect -728 35818 -694 35837
rect -660 35818 -626 35837
rect -592 35818 -558 35837
rect -524 35818 -490 35837
rect -1067 35803 -1034 35818
rect -995 35803 -966 35818
rect -923 35803 -898 35818
rect -851 35803 -830 35818
rect -779 35803 -762 35818
rect -707 35803 -694 35818
rect -635 35803 -626 35818
rect -563 35803 -558 35818
rect -491 35803 -490 35818
rect -456 35818 -422 35837
rect -388 35818 -354 35837
rect -320 35818 -286 35837
rect -456 35803 -453 35818
rect -388 35803 -381 35818
rect -320 35803 -309 35818
rect -252 35803 -218 35837
rect -184 35803 -153 35837
rect -2969 35784 -2829 35803
rect -2795 35784 -2757 35803
rect -2723 35784 -2685 35803
rect -2651 35784 -2613 35803
rect -2579 35784 -2541 35803
rect -2507 35784 -2469 35803
rect -2435 35784 -2397 35803
rect -2363 35784 -2325 35803
rect -2291 35784 -2253 35803
rect -2219 35784 -2181 35803
rect -2147 35784 -2109 35803
rect -2075 35784 -2037 35803
rect -2003 35784 -1965 35803
rect -1931 35784 -1893 35803
rect -1859 35784 -1821 35803
rect -1787 35784 -1749 35803
rect -1715 35784 -1677 35803
rect -1643 35784 -1605 35803
rect -1571 35784 -1533 35803
rect -1499 35784 -1461 35803
rect -1427 35784 -1389 35803
rect -1355 35784 -1317 35803
rect -1283 35784 -1245 35803
rect -1211 35784 -1173 35803
rect -1139 35784 -1101 35803
rect -1067 35784 -1029 35803
rect -995 35784 -957 35803
rect -923 35784 -885 35803
rect -851 35784 -813 35803
rect -779 35784 -741 35803
rect -707 35784 -669 35803
rect -635 35784 -597 35803
rect -563 35784 -525 35803
rect -491 35784 -453 35803
rect -419 35784 -381 35803
rect -347 35784 -309 35803
rect -275 35784 -153 35803
rect -2969 35768 -153 35784
rect -2969 35734 -2938 35768
rect -2904 35734 -2870 35768
rect -2836 35745 -2802 35768
rect -2768 35745 -2734 35768
rect -2700 35745 -2666 35768
rect -2632 35745 -2598 35768
rect -2564 35745 -2530 35768
rect -2496 35745 -2462 35768
rect -2428 35745 -2394 35768
rect -2836 35734 -2829 35745
rect -2768 35734 -2757 35745
rect -2700 35734 -2685 35745
rect -2632 35734 -2613 35745
rect -2564 35734 -2541 35745
rect -2496 35734 -2469 35745
rect -2428 35734 -2397 35745
rect -2360 35734 -2326 35768
rect -2292 35745 -2258 35768
rect -2224 35745 -2190 35768
rect -2156 35745 -2122 35768
rect -2088 35745 -2054 35768
rect -2020 35745 -1986 35768
rect -1952 35745 -1918 35768
rect -1884 35745 -1850 35768
rect -1816 35745 -1782 35768
rect -1748 35745 -1714 35768
rect -2291 35734 -2258 35745
rect -2219 35734 -2190 35745
rect -2147 35734 -2122 35745
rect -2075 35734 -2054 35745
rect -2003 35734 -1986 35745
rect -1931 35734 -1918 35745
rect -1859 35734 -1850 35745
rect -1787 35734 -1782 35745
rect -1715 35734 -1714 35745
rect -1680 35745 -1646 35768
rect -1612 35745 -1578 35768
rect -1544 35745 -1510 35768
rect -1476 35745 -1442 35768
rect -1408 35745 -1374 35768
rect -1340 35745 -1306 35768
rect -1272 35745 -1238 35768
rect -1204 35745 -1170 35768
rect -1680 35734 -1677 35745
rect -1612 35734 -1605 35745
rect -1544 35734 -1533 35745
rect -1476 35734 -1461 35745
rect -1408 35734 -1389 35745
rect -1340 35734 -1317 35745
rect -1272 35734 -1245 35745
rect -1204 35734 -1173 35745
rect -1136 35734 -1102 35768
rect -1068 35745 -1034 35768
rect -1000 35745 -966 35768
rect -932 35745 -898 35768
rect -864 35745 -830 35768
rect -796 35745 -762 35768
rect -728 35745 -694 35768
rect -660 35745 -626 35768
rect -592 35745 -558 35768
rect -524 35745 -490 35768
rect -1067 35734 -1034 35745
rect -995 35734 -966 35745
rect -923 35734 -898 35745
rect -851 35734 -830 35745
rect -779 35734 -762 35745
rect -707 35734 -694 35745
rect -635 35734 -626 35745
rect -563 35734 -558 35745
rect -491 35734 -490 35745
rect -456 35745 -422 35768
rect -388 35745 -354 35768
rect -320 35745 -286 35768
rect -456 35734 -453 35745
rect -388 35734 -381 35745
rect -320 35734 -309 35745
rect -252 35734 -218 35768
rect -184 35734 -153 35768
rect -2969 35711 -2829 35734
rect -2795 35711 -2757 35734
rect -2723 35711 -2685 35734
rect -2651 35711 -2613 35734
rect -2579 35711 -2541 35734
rect -2507 35711 -2469 35734
rect -2435 35711 -2397 35734
rect -2363 35711 -2325 35734
rect -2291 35711 -2253 35734
rect -2219 35711 -2181 35734
rect -2147 35711 -2109 35734
rect -2075 35711 -2037 35734
rect -2003 35711 -1965 35734
rect -1931 35711 -1893 35734
rect -1859 35711 -1821 35734
rect -1787 35711 -1749 35734
rect -1715 35711 -1677 35734
rect -1643 35711 -1605 35734
rect -1571 35711 -1533 35734
rect -1499 35711 -1461 35734
rect -1427 35711 -1389 35734
rect -1355 35711 -1317 35734
rect -1283 35711 -1245 35734
rect -1211 35711 -1173 35734
rect -1139 35711 -1101 35734
rect -1067 35711 -1029 35734
rect -995 35711 -957 35734
rect -923 35711 -885 35734
rect -851 35711 -813 35734
rect -779 35711 -741 35734
rect -707 35711 -669 35734
rect -635 35711 -597 35734
rect -563 35711 -525 35734
rect -491 35711 -453 35734
rect -419 35711 -381 35734
rect -347 35711 -309 35734
rect -275 35711 -153 35734
rect -2969 35699 -153 35711
rect -2969 35665 -2938 35699
rect -2904 35665 -2870 35699
rect -2836 35672 -2802 35699
rect -2768 35672 -2734 35699
rect -2700 35672 -2666 35699
rect -2632 35672 -2598 35699
rect -2564 35672 -2530 35699
rect -2496 35672 -2462 35699
rect -2428 35672 -2394 35699
rect -2836 35665 -2829 35672
rect -2768 35665 -2757 35672
rect -2700 35665 -2685 35672
rect -2632 35665 -2613 35672
rect -2564 35665 -2541 35672
rect -2496 35665 -2469 35672
rect -2428 35665 -2397 35672
rect -2360 35665 -2326 35699
rect -2292 35672 -2258 35699
rect -2224 35672 -2190 35699
rect -2156 35672 -2122 35699
rect -2088 35672 -2054 35699
rect -2020 35672 -1986 35699
rect -1952 35672 -1918 35699
rect -1884 35672 -1850 35699
rect -1816 35672 -1782 35699
rect -1748 35672 -1714 35699
rect -2291 35665 -2258 35672
rect -2219 35665 -2190 35672
rect -2147 35665 -2122 35672
rect -2075 35665 -2054 35672
rect -2003 35665 -1986 35672
rect -1931 35665 -1918 35672
rect -1859 35665 -1850 35672
rect -1787 35665 -1782 35672
rect -1715 35665 -1714 35672
rect -1680 35672 -1646 35699
rect -1612 35672 -1578 35699
rect -1544 35672 -1510 35699
rect -1476 35672 -1442 35699
rect -1408 35672 -1374 35699
rect -1340 35672 -1306 35699
rect -1272 35672 -1238 35699
rect -1204 35672 -1170 35699
rect -1680 35665 -1677 35672
rect -1612 35665 -1605 35672
rect -1544 35665 -1533 35672
rect -1476 35665 -1461 35672
rect -1408 35665 -1389 35672
rect -1340 35665 -1317 35672
rect -1272 35665 -1245 35672
rect -1204 35665 -1173 35672
rect -1136 35665 -1102 35699
rect -1068 35672 -1034 35699
rect -1000 35672 -966 35699
rect -932 35672 -898 35699
rect -864 35672 -830 35699
rect -796 35672 -762 35699
rect -728 35672 -694 35699
rect -660 35672 -626 35699
rect -592 35672 -558 35699
rect -524 35672 -490 35699
rect -1067 35665 -1034 35672
rect -995 35665 -966 35672
rect -923 35665 -898 35672
rect -851 35665 -830 35672
rect -779 35665 -762 35672
rect -707 35665 -694 35672
rect -635 35665 -626 35672
rect -563 35665 -558 35672
rect -491 35665 -490 35672
rect -456 35672 -422 35699
rect -388 35672 -354 35699
rect -320 35672 -286 35699
rect -456 35665 -453 35672
rect -388 35665 -381 35672
rect -320 35665 -309 35672
rect -252 35665 -218 35699
rect -184 35665 -153 35699
rect -2969 35638 -2829 35665
rect -2795 35638 -2757 35665
rect -2723 35638 -2685 35665
rect -2651 35638 -2613 35665
rect -2579 35638 -2541 35665
rect -2507 35638 -2469 35665
rect -2435 35638 -2397 35665
rect -2363 35638 -2325 35665
rect -2291 35638 -2253 35665
rect -2219 35638 -2181 35665
rect -2147 35638 -2109 35665
rect -2075 35638 -2037 35665
rect -2003 35638 -1965 35665
rect -1931 35638 -1893 35665
rect -1859 35638 -1821 35665
rect -1787 35638 -1749 35665
rect -1715 35638 -1677 35665
rect -1643 35638 -1605 35665
rect -1571 35638 -1533 35665
rect -1499 35638 -1461 35665
rect -1427 35638 -1389 35665
rect -1355 35638 -1317 35665
rect -1283 35638 -1245 35665
rect -1211 35638 -1173 35665
rect -1139 35638 -1101 35665
rect -1067 35638 -1029 35665
rect -995 35638 -957 35665
rect -923 35638 -885 35665
rect -851 35638 -813 35665
rect -779 35638 -741 35665
rect -707 35638 -669 35665
rect -635 35638 -597 35665
rect -563 35638 -525 35665
rect -491 35638 -453 35665
rect -419 35638 -381 35665
rect -347 35638 -309 35665
rect -275 35638 -153 35665
rect -2969 35630 -153 35638
rect -2969 35596 -2938 35630
rect -2904 35596 -2870 35630
rect -2836 35599 -2802 35630
rect -2768 35599 -2734 35630
rect -2700 35599 -2666 35630
rect -2632 35599 -2598 35630
rect -2564 35599 -2530 35630
rect -2496 35599 -2462 35630
rect -2428 35599 -2394 35630
rect -2836 35596 -2829 35599
rect -2768 35596 -2757 35599
rect -2700 35596 -2685 35599
rect -2632 35596 -2613 35599
rect -2564 35596 -2541 35599
rect -2496 35596 -2469 35599
rect -2428 35596 -2397 35599
rect -2360 35596 -2326 35630
rect -2292 35599 -2258 35630
rect -2224 35599 -2190 35630
rect -2156 35599 -2122 35630
rect -2088 35599 -2054 35630
rect -2020 35599 -1986 35630
rect -1952 35599 -1918 35630
rect -1884 35599 -1850 35630
rect -1816 35599 -1782 35630
rect -1748 35599 -1714 35630
rect -2291 35596 -2258 35599
rect -2219 35596 -2190 35599
rect -2147 35596 -2122 35599
rect -2075 35596 -2054 35599
rect -2003 35596 -1986 35599
rect -1931 35596 -1918 35599
rect -1859 35596 -1850 35599
rect -1787 35596 -1782 35599
rect -1715 35596 -1714 35599
rect -1680 35599 -1646 35630
rect -1612 35599 -1578 35630
rect -1544 35599 -1510 35630
rect -1476 35599 -1442 35630
rect -1408 35599 -1374 35630
rect -1340 35599 -1306 35630
rect -1272 35599 -1238 35630
rect -1204 35599 -1170 35630
rect -1680 35596 -1677 35599
rect -1612 35596 -1605 35599
rect -1544 35596 -1533 35599
rect -1476 35596 -1461 35599
rect -1408 35596 -1389 35599
rect -1340 35596 -1317 35599
rect -1272 35596 -1245 35599
rect -1204 35596 -1173 35599
rect -1136 35596 -1102 35630
rect -1068 35599 -1034 35630
rect -1000 35599 -966 35630
rect -932 35599 -898 35630
rect -864 35599 -830 35630
rect -796 35599 -762 35630
rect -728 35599 -694 35630
rect -660 35599 -626 35630
rect -592 35599 -558 35630
rect -524 35599 -490 35630
rect -1067 35596 -1034 35599
rect -995 35596 -966 35599
rect -923 35596 -898 35599
rect -851 35596 -830 35599
rect -779 35596 -762 35599
rect -707 35596 -694 35599
rect -635 35596 -626 35599
rect -563 35596 -558 35599
rect -491 35596 -490 35599
rect -456 35599 -422 35630
rect -388 35599 -354 35630
rect -320 35599 -286 35630
rect -456 35596 -453 35599
rect -388 35596 -381 35599
rect -320 35596 -309 35599
rect -252 35596 -218 35630
rect -184 35596 -153 35630
rect -2969 35565 -2829 35596
rect -2795 35565 -2757 35596
rect -2723 35565 -2685 35596
rect -2651 35565 -2613 35596
rect -2579 35565 -2541 35596
rect -2507 35565 -2469 35596
rect -2435 35565 -2397 35596
rect -2363 35565 -2325 35596
rect -2291 35565 -2253 35596
rect -2219 35565 -2181 35596
rect -2147 35565 -2109 35596
rect -2075 35565 -2037 35596
rect -2003 35565 -1965 35596
rect -1931 35565 -1893 35596
rect -1859 35565 -1821 35596
rect -1787 35565 -1749 35596
rect -1715 35565 -1677 35596
rect -1643 35565 -1605 35596
rect -1571 35565 -1533 35596
rect -1499 35565 -1461 35596
rect -1427 35565 -1389 35596
rect -1355 35565 -1317 35596
rect -1283 35565 -1245 35596
rect -1211 35565 -1173 35596
rect -1139 35565 -1101 35596
rect -1067 35565 -1029 35596
rect -995 35565 -957 35596
rect -923 35565 -885 35596
rect -851 35565 -813 35596
rect -779 35565 -741 35596
rect -707 35565 -669 35596
rect -635 35565 -597 35596
rect -563 35565 -525 35596
rect -491 35565 -453 35596
rect -419 35565 -381 35596
rect -347 35565 -309 35596
rect -275 35565 -153 35596
rect -2969 35561 -153 35565
rect -2969 35527 -2938 35561
rect -2904 35527 -2870 35561
rect -2836 35527 -2802 35561
rect -2768 35527 -2734 35561
rect -2700 35527 -2666 35561
rect -2632 35527 -2598 35561
rect -2564 35527 -2530 35561
rect -2496 35527 -2462 35561
rect -2428 35527 -2394 35561
rect -2360 35527 -2326 35561
rect -2292 35527 -2258 35561
rect -2224 35527 -2190 35561
rect -2156 35527 -2122 35561
rect -2088 35527 -2054 35561
rect -2020 35527 -1986 35561
rect -1952 35527 -1918 35561
rect -1884 35527 -1850 35561
rect -1816 35527 -1782 35561
rect -1748 35527 -1714 35561
rect -1680 35527 -1646 35561
rect -1612 35527 -1578 35561
rect -1544 35527 -1510 35561
rect -1476 35527 -1442 35561
rect -1408 35527 -1374 35561
rect -1340 35527 -1306 35561
rect -1272 35527 -1238 35561
rect -1204 35527 -1170 35561
rect -1136 35527 -1102 35561
rect -1068 35527 -1034 35561
rect -1000 35527 -966 35561
rect -932 35527 -898 35561
rect -864 35527 -830 35561
rect -796 35527 -762 35561
rect -728 35527 -694 35561
rect -660 35527 -626 35561
rect -592 35527 -558 35561
rect -524 35527 -490 35561
rect -456 35527 -422 35561
rect -388 35527 -354 35561
rect -320 35527 -286 35561
rect -252 35527 -218 35561
rect -184 35527 -153 35561
rect -2969 35526 -153 35527
rect -2969 35492 -2829 35526
rect -2795 35492 -2757 35526
rect -2723 35492 -2685 35526
rect -2651 35492 -2613 35526
rect -2579 35492 -2541 35526
rect -2507 35492 -2469 35526
rect -2435 35492 -2397 35526
rect -2363 35492 -2325 35526
rect -2291 35492 -2253 35526
rect -2219 35492 -2181 35526
rect -2147 35492 -2109 35526
rect -2075 35492 -2037 35526
rect -2003 35492 -1965 35526
rect -1931 35492 -1893 35526
rect -1859 35492 -1821 35526
rect -1787 35492 -1749 35526
rect -1715 35492 -1677 35526
rect -1643 35492 -1605 35526
rect -1571 35492 -1533 35526
rect -1499 35492 -1461 35526
rect -1427 35492 -1389 35526
rect -1355 35492 -1317 35526
rect -1283 35492 -1245 35526
rect -1211 35492 -1173 35526
rect -1139 35492 -1101 35526
rect -1067 35492 -1029 35526
rect -995 35492 -957 35526
rect -923 35492 -885 35526
rect -851 35492 -813 35526
rect -779 35492 -741 35526
rect -707 35492 -669 35526
rect -635 35492 -597 35526
rect -563 35492 -525 35526
rect -491 35492 -453 35526
rect -419 35492 -381 35526
rect -347 35492 -309 35526
rect -275 35492 -153 35526
rect -2969 35458 -2938 35492
rect -2904 35458 -2870 35492
rect -2836 35458 -2802 35492
rect -2768 35458 -2734 35492
rect -2700 35458 -2666 35492
rect -2632 35458 -2598 35492
rect -2564 35458 -2530 35492
rect -2496 35458 -2462 35492
rect -2428 35458 -2394 35492
rect -2360 35458 -2326 35492
rect -2292 35458 -2258 35492
rect -2224 35458 -2190 35492
rect -2156 35458 -2122 35492
rect -2088 35458 -2054 35492
rect -2020 35458 -1986 35492
rect -1952 35458 -1918 35492
rect -1884 35458 -1850 35492
rect -1816 35458 -1782 35492
rect -1748 35458 -1714 35492
rect -1680 35458 -1646 35492
rect -1612 35458 -1578 35492
rect -1544 35458 -1510 35492
rect -1476 35458 -1442 35492
rect -1408 35458 -1374 35492
rect -1340 35458 -1306 35492
rect -1272 35458 -1238 35492
rect -1204 35458 -1170 35492
rect -1136 35458 -1102 35492
rect -1068 35458 -1034 35492
rect -1000 35458 -966 35492
rect -932 35458 -898 35492
rect -864 35458 -830 35492
rect -796 35458 -762 35492
rect -728 35458 -694 35492
rect -660 35458 -626 35492
rect -592 35458 -558 35492
rect -524 35458 -490 35492
rect -456 35458 -422 35492
rect -388 35458 -354 35492
rect -320 35458 -286 35492
rect -252 35458 -218 35492
rect -184 35458 -153 35492
rect -2969 35453 -153 35458
rect -2969 35423 -2829 35453
rect -2795 35423 -2757 35453
rect -2723 35423 -2685 35453
rect -2651 35423 -2613 35453
rect -2579 35423 -2541 35453
rect -2507 35423 -2469 35453
rect -2435 35423 -2397 35453
rect -2363 35423 -2325 35453
rect -2291 35423 -2253 35453
rect -2219 35423 -2181 35453
rect -2147 35423 -2109 35453
rect -2075 35423 -2037 35453
rect -2003 35423 -1965 35453
rect -1931 35423 -1893 35453
rect -1859 35423 -1821 35453
rect -1787 35423 -1749 35453
rect -1715 35423 -1677 35453
rect -1643 35423 -1605 35453
rect -1571 35423 -1533 35453
rect -1499 35423 -1461 35453
rect -1427 35423 -1389 35453
rect -1355 35423 -1317 35453
rect -1283 35423 -1245 35453
rect -1211 35423 -1173 35453
rect -1139 35423 -1101 35453
rect -1067 35423 -1029 35453
rect -995 35423 -957 35453
rect -923 35423 -885 35453
rect -851 35423 -813 35453
rect -779 35423 -741 35453
rect -707 35423 -669 35453
rect -635 35423 -597 35453
rect -563 35423 -525 35453
rect -491 35423 -453 35453
rect -419 35423 -381 35453
rect -347 35423 -309 35453
rect -275 35423 -153 35453
rect -2969 35389 -2938 35423
rect -2904 35389 -2870 35423
rect -2836 35419 -2829 35423
rect -2768 35419 -2757 35423
rect -2700 35419 -2685 35423
rect -2632 35419 -2613 35423
rect -2564 35419 -2541 35423
rect -2496 35419 -2469 35423
rect -2428 35419 -2397 35423
rect -2836 35389 -2802 35419
rect -2768 35389 -2734 35419
rect -2700 35389 -2666 35419
rect -2632 35389 -2598 35419
rect -2564 35389 -2530 35419
rect -2496 35389 -2462 35419
rect -2428 35389 -2394 35419
rect -2360 35389 -2326 35423
rect -2291 35419 -2258 35423
rect -2219 35419 -2190 35423
rect -2147 35419 -2122 35423
rect -2075 35419 -2054 35423
rect -2003 35419 -1986 35423
rect -1931 35419 -1918 35423
rect -1859 35419 -1850 35423
rect -1787 35419 -1782 35423
rect -1715 35419 -1714 35423
rect -2292 35389 -2258 35419
rect -2224 35389 -2190 35419
rect -2156 35389 -2122 35419
rect -2088 35389 -2054 35419
rect -2020 35389 -1986 35419
rect -1952 35389 -1918 35419
rect -1884 35389 -1850 35419
rect -1816 35389 -1782 35419
rect -1748 35389 -1714 35419
rect -1680 35419 -1677 35423
rect -1612 35419 -1605 35423
rect -1544 35419 -1533 35423
rect -1476 35419 -1461 35423
rect -1408 35419 -1389 35423
rect -1340 35419 -1317 35423
rect -1272 35419 -1245 35423
rect -1204 35419 -1173 35423
rect -1680 35389 -1646 35419
rect -1612 35389 -1578 35419
rect -1544 35389 -1510 35419
rect -1476 35389 -1442 35419
rect -1408 35389 -1374 35419
rect -1340 35389 -1306 35419
rect -1272 35389 -1238 35419
rect -1204 35389 -1170 35419
rect -1136 35389 -1102 35423
rect -1067 35419 -1034 35423
rect -995 35419 -966 35423
rect -923 35419 -898 35423
rect -851 35419 -830 35423
rect -779 35419 -762 35423
rect -707 35419 -694 35423
rect -635 35419 -626 35423
rect -563 35419 -558 35423
rect -491 35419 -490 35423
rect -1068 35389 -1034 35419
rect -1000 35389 -966 35419
rect -932 35389 -898 35419
rect -864 35389 -830 35419
rect -796 35389 -762 35419
rect -728 35389 -694 35419
rect -660 35389 -626 35419
rect -592 35389 -558 35419
rect -524 35389 -490 35419
rect -456 35419 -453 35423
rect -388 35419 -381 35423
rect -320 35419 -309 35423
rect -456 35389 -422 35419
rect -388 35389 -354 35419
rect -320 35389 -286 35419
rect -252 35389 -218 35423
rect -184 35389 -153 35423
rect -2969 35380 -153 35389
rect -2969 35354 -2829 35380
rect -2795 35354 -2757 35380
rect -2723 35354 -2685 35380
rect -2651 35354 -2613 35380
rect -2579 35354 -2541 35380
rect -2507 35354 -2469 35380
rect -2435 35354 -2397 35380
rect -2363 35354 -2325 35380
rect -2291 35354 -2253 35380
rect -2219 35354 -2181 35380
rect -2147 35354 -2109 35380
rect -2075 35354 -2037 35380
rect -2003 35354 -1965 35380
rect -1931 35354 -1893 35380
rect -1859 35354 -1821 35380
rect -1787 35354 -1749 35380
rect -1715 35354 -1677 35380
rect -1643 35354 -1605 35380
rect -1571 35354 -1533 35380
rect -1499 35354 -1461 35380
rect -1427 35354 -1389 35380
rect -1355 35354 -1317 35380
rect -1283 35354 -1245 35380
rect -1211 35354 -1173 35380
rect -1139 35354 -1101 35380
rect -1067 35354 -1029 35380
rect -995 35354 -957 35380
rect -923 35354 -885 35380
rect -851 35354 -813 35380
rect -779 35354 -741 35380
rect -707 35354 -669 35380
rect -635 35354 -597 35380
rect -563 35354 -525 35380
rect -491 35354 -453 35380
rect -419 35354 -381 35380
rect -347 35354 -309 35380
rect -275 35354 -153 35380
rect -2969 35320 -2938 35354
rect -2904 35320 -2870 35354
rect -2836 35346 -2829 35354
rect -2768 35346 -2757 35354
rect -2700 35346 -2685 35354
rect -2632 35346 -2613 35354
rect -2564 35346 -2541 35354
rect -2496 35346 -2469 35354
rect -2428 35346 -2397 35354
rect -2836 35320 -2802 35346
rect -2768 35320 -2734 35346
rect -2700 35320 -2666 35346
rect -2632 35320 -2598 35346
rect -2564 35320 -2530 35346
rect -2496 35320 -2462 35346
rect -2428 35320 -2394 35346
rect -2360 35320 -2326 35354
rect -2291 35346 -2258 35354
rect -2219 35346 -2190 35354
rect -2147 35346 -2122 35354
rect -2075 35346 -2054 35354
rect -2003 35346 -1986 35354
rect -1931 35346 -1918 35354
rect -1859 35346 -1850 35354
rect -1787 35346 -1782 35354
rect -1715 35346 -1714 35354
rect -2292 35320 -2258 35346
rect -2224 35320 -2190 35346
rect -2156 35320 -2122 35346
rect -2088 35320 -2054 35346
rect -2020 35320 -1986 35346
rect -1952 35320 -1918 35346
rect -1884 35320 -1850 35346
rect -1816 35320 -1782 35346
rect -1748 35320 -1714 35346
rect -1680 35346 -1677 35354
rect -1612 35346 -1605 35354
rect -1544 35346 -1533 35354
rect -1476 35346 -1461 35354
rect -1408 35346 -1389 35354
rect -1340 35346 -1317 35354
rect -1272 35346 -1245 35354
rect -1204 35346 -1173 35354
rect -1680 35320 -1646 35346
rect -1612 35320 -1578 35346
rect -1544 35320 -1510 35346
rect -1476 35320 -1442 35346
rect -1408 35320 -1374 35346
rect -1340 35320 -1306 35346
rect -1272 35320 -1238 35346
rect -1204 35320 -1170 35346
rect -1136 35320 -1102 35354
rect -1067 35346 -1034 35354
rect -995 35346 -966 35354
rect -923 35346 -898 35354
rect -851 35346 -830 35354
rect -779 35346 -762 35354
rect -707 35346 -694 35354
rect -635 35346 -626 35354
rect -563 35346 -558 35354
rect -491 35346 -490 35354
rect -1068 35320 -1034 35346
rect -1000 35320 -966 35346
rect -932 35320 -898 35346
rect -864 35320 -830 35346
rect -796 35320 -762 35346
rect -728 35320 -694 35346
rect -660 35320 -626 35346
rect -592 35320 -558 35346
rect -524 35320 -490 35346
rect -456 35346 -453 35354
rect -388 35346 -381 35354
rect -320 35346 -309 35354
rect -456 35320 -422 35346
rect -388 35320 -354 35346
rect -320 35320 -286 35346
rect -252 35320 -218 35354
rect -184 35320 -153 35354
rect -2969 35307 -153 35320
rect -2969 35285 -2829 35307
rect -2795 35285 -2757 35307
rect -2723 35285 -2685 35307
rect -2651 35285 -2613 35307
rect -2579 35285 -2541 35307
rect -2507 35285 -2469 35307
rect -2435 35285 -2397 35307
rect -2363 35285 -2325 35307
rect -2291 35285 -2253 35307
rect -2219 35285 -2181 35307
rect -2147 35285 -2109 35307
rect -2075 35285 -2037 35307
rect -2003 35285 -1965 35307
rect -1931 35285 -1893 35307
rect -1859 35285 -1821 35307
rect -1787 35285 -1749 35307
rect -1715 35285 -1677 35307
rect -1643 35285 -1605 35307
rect -1571 35285 -1533 35307
rect -1499 35285 -1461 35307
rect -1427 35285 -1389 35307
rect -1355 35285 -1317 35307
rect -1283 35285 -1245 35307
rect -1211 35285 -1173 35307
rect -1139 35285 -1101 35307
rect -1067 35285 -1029 35307
rect -995 35285 -957 35307
rect -923 35285 -885 35307
rect -851 35285 -813 35307
rect -779 35285 -741 35307
rect -707 35285 -669 35307
rect -635 35285 -597 35307
rect -563 35285 -525 35307
rect -491 35285 -453 35307
rect -419 35285 -381 35307
rect -347 35285 -309 35307
rect -275 35285 -153 35307
rect -2969 35251 -2938 35285
rect -2904 35251 -2870 35285
rect -2836 35273 -2829 35285
rect -2768 35273 -2757 35285
rect -2700 35273 -2685 35285
rect -2632 35273 -2613 35285
rect -2564 35273 -2541 35285
rect -2496 35273 -2469 35285
rect -2428 35273 -2397 35285
rect -2836 35251 -2802 35273
rect -2768 35251 -2734 35273
rect -2700 35251 -2666 35273
rect -2632 35251 -2598 35273
rect -2564 35251 -2530 35273
rect -2496 35251 -2462 35273
rect -2428 35251 -2394 35273
rect -2360 35251 -2326 35285
rect -2291 35273 -2258 35285
rect -2219 35273 -2190 35285
rect -2147 35273 -2122 35285
rect -2075 35273 -2054 35285
rect -2003 35273 -1986 35285
rect -1931 35273 -1918 35285
rect -1859 35273 -1850 35285
rect -1787 35273 -1782 35285
rect -1715 35273 -1714 35285
rect -2292 35251 -2258 35273
rect -2224 35251 -2190 35273
rect -2156 35251 -2122 35273
rect -2088 35251 -2054 35273
rect -2020 35251 -1986 35273
rect -1952 35251 -1918 35273
rect -1884 35251 -1850 35273
rect -1816 35251 -1782 35273
rect -1748 35251 -1714 35273
rect -1680 35273 -1677 35285
rect -1612 35273 -1605 35285
rect -1544 35273 -1533 35285
rect -1476 35273 -1461 35285
rect -1408 35273 -1389 35285
rect -1340 35273 -1317 35285
rect -1272 35273 -1245 35285
rect -1204 35273 -1173 35285
rect -1680 35251 -1646 35273
rect -1612 35251 -1578 35273
rect -1544 35251 -1510 35273
rect -1476 35251 -1442 35273
rect -1408 35251 -1374 35273
rect -1340 35251 -1306 35273
rect -1272 35251 -1238 35273
rect -1204 35251 -1170 35273
rect -1136 35251 -1102 35285
rect -1067 35273 -1034 35285
rect -995 35273 -966 35285
rect -923 35273 -898 35285
rect -851 35273 -830 35285
rect -779 35273 -762 35285
rect -707 35273 -694 35285
rect -635 35273 -626 35285
rect -563 35273 -558 35285
rect -491 35273 -490 35285
rect -1068 35251 -1034 35273
rect -1000 35251 -966 35273
rect -932 35251 -898 35273
rect -864 35251 -830 35273
rect -796 35251 -762 35273
rect -728 35251 -694 35273
rect -660 35251 -626 35273
rect -592 35251 -558 35273
rect -524 35251 -490 35273
rect -456 35273 -453 35285
rect -388 35273 -381 35285
rect -320 35273 -309 35285
rect -456 35251 -422 35273
rect -388 35251 -354 35273
rect -320 35251 -286 35273
rect -252 35251 -218 35285
rect -184 35251 -153 35285
rect -2969 35234 -153 35251
rect -2969 35216 -2829 35234
rect -2795 35216 -2757 35234
rect -2723 35216 -2685 35234
rect -2651 35216 -2613 35234
rect -2579 35216 -2541 35234
rect -2507 35216 -2469 35234
rect -2435 35216 -2397 35234
rect -2363 35216 -2325 35234
rect -2291 35216 -2253 35234
rect -2219 35216 -2181 35234
rect -2147 35216 -2109 35234
rect -2075 35216 -2037 35234
rect -2003 35216 -1965 35234
rect -1931 35216 -1893 35234
rect -1859 35216 -1821 35234
rect -1787 35216 -1749 35234
rect -1715 35216 -1677 35234
rect -1643 35216 -1605 35234
rect -1571 35216 -1533 35234
rect -1499 35216 -1461 35234
rect -1427 35216 -1389 35234
rect -1355 35216 -1317 35234
rect -1283 35216 -1245 35234
rect -1211 35216 -1173 35234
rect -1139 35216 -1101 35234
rect -1067 35216 -1029 35234
rect -995 35216 -957 35234
rect -923 35216 -885 35234
rect -851 35216 -813 35234
rect -779 35216 -741 35234
rect -707 35216 -669 35234
rect -635 35216 -597 35234
rect -563 35216 -525 35234
rect -491 35216 -453 35234
rect -419 35216 -381 35234
rect -347 35216 -309 35234
rect -275 35216 -153 35234
rect -2969 35182 -2938 35216
rect -2904 35182 -2870 35216
rect -2836 35200 -2829 35216
rect -2768 35200 -2757 35216
rect -2700 35200 -2685 35216
rect -2632 35200 -2613 35216
rect -2564 35200 -2541 35216
rect -2496 35200 -2469 35216
rect -2428 35200 -2397 35216
rect -2836 35182 -2802 35200
rect -2768 35182 -2734 35200
rect -2700 35182 -2666 35200
rect -2632 35182 -2598 35200
rect -2564 35182 -2530 35200
rect -2496 35182 -2462 35200
rect -2428 35182 -2394 35200
rect -2360 35182 -2326 35216
rect -2291 35200 -2258 35216
rect -2219 35200 -2190 35216
rect -2147 35200 -2122 35216
rect -2075 35200 -2054 35216
rect -2003 35200 -1986 35216
rect -1931 35200 -1918 35216
rect -1859 35200 -1850 35216
rect -1787 35200 -1782 35216
rect -1715 35200 -1714 35216
rect -2292 35182 -2258 35200
rect -2224 35182 -2190 35200
rect -2156 35182 -2122 35200
rect -2088 35182 -2054 35200
rect -2020 35182 -1986 35200
rect -1952 35182 -1918 35200
rect -1884 35182 -1850 35200
rect -1816 35182 -1782 35200
rect -1748 35182 -1714 35200
rect -1680 35200 -1677 35216
rect -1612 35200 -1605 35216
rect -1544 35200 -1533 35216
rect -1476 35200 -1461 35216
rect -1408 35200 -1389 35216
rect -1340 35200 -1317 35216
rect -1272 35200 -1245 35216
rect -1204 35200 -1173 35216
rect -1680 35182 -1646 35200
rect -1612 35182 -1578 35200
rect -1544 35182 -1510 35200
rect -1476 35182 -1442 35200
rect -1408 35182 -1374 35200
rect -1340 35182 -1306 35200
rect -1272 35182 -1238 35200
rect -1204 35182 -1170 35200
rect -1136 35182 -1102 35216
rect -1067 35200 -1034 35216
rect -995 35200 -966 35216
rect -923 35200 -898 35216
rect -851 35200 -830 35216
rect -779 35200 -762 35216
rect -707 35200 -694 35216
rect -635 35200 -626 35216
rect -563 35200 -558 35216
rect -491 35200 -490 35216
rect -1068 35182 -1034 35200
rect -1000 35182 -966 35200
rect -932 35182 -898 35200
rect -864 35182 -830 35200
rect -796 35182 -762 35200
rect -728 35182 -694 35200
rect -660 35182 -626 35200
rect -592 35182 -558 35200
rect -524 35182 -490 35200
rect -456 35200 -453 35216
rect -388 35200 -381 35216
rect -320 35200 -309 35216
rect -456 35182 -422 35200
rect -388 35182 -354 35200
rect -320 35182 -286 35200
rect -252 35182 -218 35216
rect -184 35182 -153 35216
rect -2969 35161 -153 35182
rect -2969 35147 -2829 35161
rect -2795 35147 -2757 35161
rect -2723 35147 -2685 35161
rect -2651 35147 -2613 35161
rect -2579 35147 -2541 35161
rect -2507 35147 -2469 35161
rect -2435 35147 -2397 35161
rect -2363 35147 -2325 35161
rect -2291 35147 -2253 35161
rect -2219 35147 -2181 35161
rect -2147 35147 -2109 35161
rect -2075 35147 -2037 35161
rect -2003 35147 -1965 35161
rect -1931 35147 -1893 35161
rect -1859 35147 -1821 35161
rect -1787 35147 -1749 35161
rect -1715 35147 -1677 35161
rect -1643 35147 -1605 35161
rect -1571 35147 -1533 35161
rect -1499 35147 -1461 35161
rect -1427 35147 -1389 35161
rect -1355 35147 -1317 35161
rect -1283 35147 -1245 35161
rect -1211 35147 -1173 35161
rect -1139 35147 -1101 35161
rect -1067 35147 -1029 35161
rect -995 35147 -957 35161
rect -923 35147 -885 35161
rect -851 35147 -813 35161
rect -779 35147 -741 35161
rect -707 35147 -669 35161
rect -635 35147 -597 35161
rect -563 35147 -525 35161
rect -491 35147 -453 35161
rect -419 35147 -381 35161
rect -347 35147 -309 35161
rect -275 35147 -153 35161
rect -2969 35113 -2938 35147
rect -2904 35113 -2870 35147
rect -2836 35127 -2829 35147
rect -2768 35127 -2757 35147
rect -2700 35127 -2685 35147
rect -2632 35127 -2613 35147
rect -2564 35127 -2541 35147
rect -2496 35127 -2469 35147
rect -2428 35127 -2397 35147
rect -2836 35113 -2802 35127
rect -2768 35113 -2734 35127
rect -2700 35113 -2666 35127
rect -2632 35113 -2598 35127
rect -2564 35113 -2530 35127
rect -2496 35113 -2462 35127
rect -2428 35113 -2394 35127
rect -2360 35113 -2326 35147
rect -2291 35127 -2258 35147
rect -2219 35127 -2190 35147
rect -2147 35127 -2122 35147
rect -2075 35127 -2054 35147
rect -2003 35127 -1986 35147
rect -1931 35127 -1918 35147
rect -1859 35127 -1850 35147
rect -1787 35127 -1782 35147
rect -1715 35127 -1714 35147
rect -2292 35113 -2258 35127
rect -2224 35113 -2190 35127
rect -2156 35113 -2122 35127
rect -2088 35113 -2054 35127
rect -2020 35113 -1986 35127
rect -1952 35113 -1918 35127
rect -1884 35113 -1850 35127
rect -1816 35113 -1782 35127
rect -1748 35113 -1714 35127
rect -1680 35127 -1677 35147
rect -1612 35127 -1605 35147
rect -1544 35127 -1533 35147
rect -1476 35127 -1461 35147
rect -1408 35127 -1389 35147
rect -1340 35127 -1317 35147
rect -1272 35127 -1245 35147
rect -1204 35127 -1173 35147
rect -1680 35113 -1646 35127
rect -1612 35113 -1578 35127
rect -1544 35113 -1510 35127
rect -1476 35113 -1442 35127
rect -1408 35113 -1374 35127
rect -1340 35113 -1306 35127
rect -1272 35113 -1238 35127
rect -1204 35113 -1170 35127
rect -1136 35113 -1102 35147
rect -1067 35127 -1034 35147
rect -995 35127 -966 35147
rect -923 35127 -898 35147
rect -851 35127 -830 35147
rect -779 35127 -762 35147
rect -707 35127 -694 35147
rect -635 35127 -626 35147
rect -563 35127 -558 35147
rect -491 35127 -490 35147
rect -1068 35113 -1034 35127
rect -1000 35113 -966 35127
rect -932 35113 -898 35127
rect -864 35113 -830 35127
rect -796 35113 -762 35127
rect -728 35113 -694 35127
rect -660 35113 -626 35127
rect -592 35113 -558 35127
rect -524 35113 -490 35127
rect -456 35127 -453 35147
rect -388 35127 -381 35147
rect -320 35127 -309 35147
rect -456 35113 -422 35127
rect -388 35113 -354 35127
rect -320 35113 -286 35127
rect -252 35113 -218 35147
rect -184 35113 -153 35147
rect -2969 35078 -153 35113
rect -2969 35044 -2938 35078
rect -2904 35044 -2870 35078
rect -2836 35044 -2802 35078
rect -2768 35044 -2734 35078
rect -2700 35044 -2666 35078
rect -2632 35044 -2598 35078
rect -2564 35044 -2530 35078
rect -2496 35044 -2462 35078
rect -2428 35044 -2394 35078
rect -2360 35044 -2326 35078
rect -2292 35044 -2258 35078
rect -2224 35044 -2190 35078
rect -2156 35044 -2122 35078
rect -2088 35044 -2054 35078
rect -2020 35044 -1986 35078
rect -1952 35044 -1918 35078
rect -1884 35044 -1850 35078
rect -1816 35044 -1782 35078
rect -1748 35044 -1714 35078
rect -1680 35044 -1646 35078
rect -1612 35044 -1578 35078
rect -1544 35044 -1510 35078
rect -1476 35044 -1442 35078
rect -1408 35044 -1374 35078
rect -1340 35044 -1306 35078
rect -1272 35044 -1238 35078
rect -1204 35044 -1170 35078
rect -1136 35044 -1102 35078
rect -1068 35044 -1034 35078
rect -1000 35044 -966 35078
rect -932 35044 -898 35078
rect -864 35044 -830 35078
rect -796 35044 -762 35078
rect -728 35044 -694 35078
rect -660 35044 -626 35078
rect -592 35044 -558 35078
rect -524 35044 -490 35078
rect -456 35044 -422 35078
rect -388 35044 -354 35078
rect -320 35044 -286 35078
rect -252 35044 -218 35078
rect -184 35044 -153 35078
rect -2969 35020 -153 35044
rect 14 50636 228 50677
rect 14 50602 15 50636
rect 49 50632 228 50636
rect 49 50602 87 50632
rect 14 50598 87 50602
rect 121 50627 228 50632
rect 121 50598 159 50627
rect 14 50593 159 50598
rect 193 50593 228 50627
rect 14 50568 228 50593
rect 14 50534 15 50568
rect 49 50564 228 50568
rect 49 50534 87 50564
rect 14 50530 87 50534
rect 121 50559 228 50564
rect 121 50530 159 50559
rect 14 50525 159 50530
rect 193 50525 228 50559
rect 14 50500 228 50525
rect 14 50466 15 50500
rect 49 50496 228 50500
rect 49 50466 87 50496
rect 14 50462 87 50466
rect 121 50491 228 50496
rect 121 50462 159 50491
rect 14 50457 159 50462
rect 193 50457 228 50491
rect 14 50432 228 50457
rect 14 50398 15 50432
rect 49 50428 228 50432
rect 49 50398 87 50428
rect 14 50394 87 50398
rect 121 50423 228 50428
rect 121 50394 159 50423
rect 14 50389 159 50394
rect 193 50389 228 50423
rect 14 50364 228 50389
rect 14 50330 15 50364
rect 49 50360 228 50364
rect 49 50330 87 50360
rect 14 50326 87 50330
rect 121 50355 228 50360
rect 121 50326 159 50355
rect 14 50321 159 50326
rect 193 50321 228 50355
rect 14 50296 228 50321
rect 14 50262 15 50296
rect 49 50292 228 50296
rect 49 50262 87 50292
rect 14 50258 87 50262
rect 121 50287 228 50292
rect 121 50258 159 50287
rect 14 50253 159 50258
rect 193 50253 228 50287
rect 14 50228 228 50253
rect 14 50194 15 50228
rect 49 50224 228 50228
rect 49 50194 87 50224
rect 14 50190 87 50194
rect 121 50219 228 50224
rect 121 50190 159 50219
rect 14 50185 159 50190
rect 193 50185 228 50219
rect 14 50160 228 50185
rect 14 50126 15 50160
rect 49 50156 228 50160
rect 49 50126 87 50156
rect 14 50122 87 50126
rect 121 50151 228 50156
rect 121 50122 159 50151
rect 14 50117 159 50122
rect 193 50117 228 50151
rect 14 50092 228 50117
rect 14 50058 15 50092
rect 49 50088 228 50092
rect 49 50058 87 50088
rect 14 50054 87 50058
rect 121 50083 228 50088
rect 121 50054 159 50083
rect 14 50049 159 50054
rect 193 50049 228 50083
rect 14 50024 228 50049
rect 14 49990 15 50024
rect 49 50020 228 50024
rect 49 49990 87 50020
rect 14 49986 87 49990
rect 121 50015 228 50020
rect 121 49986 159 50015
rect 14 49981 159 49986
rect 193 49981 228 50015
rect 14 49956 228 49981
rect 14 49922 15 49956
rect 49 49952 228 49956
rect 49 49922 87 49952
rect 14 49918 87 49922
rect 121 49947 228 49952
rect 121 49918 159 49947
rect 14 49913 159 49918
rect 193 49913 228 49947
rect 14 49888 228 49913
rect 14 49854 15 49888
rect 49 49884 228 49888
rect 49 49854 87 49884
rect 14 49850 87 49854
rect 121 49879 228 49884
rect 121 49850 159 49879
rect 14 49845 159 49850
rect 193 49845 228 49879
rect 14 49820 228 49845
rect 14 49786 15 49820
rect 49 49816 228 49820
rect 49 49786 87 49816
rect 14 49782 87 49786
rect 121 49811 228 49816
rect 121 49782 159 49811
rect 14 49777 159 49782
rect 193 49777 228 49811
rect 14 49752 228 49777
rect 14 49718 15 49752
rect 49 49748 228 49752
rect 49 49718 87 49748
rect 14 49714 87 49718
rect 121 49743 228 49748
rect 121 49714 159 49743
rect 14 49709 159 49714
rect 193 49709 228 49743
rect 14 49684 228 49709
rect 14 49650 15 49684
rect 49 49680 228 49684
rect 49 49650 87 49680
rect 14 49646 87 49650
rect 121 49675 228 49680
rect 121 49646 159 49675
rect 14 49641 159 49646
rect 193 49641 228 49675
rect 14 49616 228 49641
rect 14 49582 15 49616
rect 49 49612 228 49616
rect 49 49582 87 49612
rect 14 49578 87 49582
rect 121 49607 228 49612
rect 121 49578 159 49607
rect 14 49573 159 49578
rect 193 49573 228 49607
rect 14 49548 228 49573
rect 14 49514 15 49548
rect 49 49544 228 49548
rect 49 49514 87 49544
rect 14 49510 87 49514
rect 121 49539 228 49544
rect 121 49510 159 49539
rect 14 49505 159 49510
rect 193 49505 228 49539
rect 14 49480 228 49505
rect 14 49446 15 49480
rect 49 49476 228 49480
rect 49 49446 87 49476
rect 14 49442 87 49446
rect 121 49471 228 49476
rect 121 49442 159 49471
rect 14 49437 159 49442
rect 193 49437 228 49471
rect 14 49412 228 49437
rect 14 49378 15 49412
rect 49 49408 228 49412
rect 49 49378 87 49408
rect 14 49374 87 49378
rect 121 49403 228 49408
rect 121 49374 159 49403
rect 14 49369 159 49374
rect 193 49369 228 49403
rect 14 49344 228 49369
rect 14 49310 15 49344
rect 49 49340 228 49344
rect 49 49310 87 49340
rect 14 49306 87 49310
rect 121 49335 228 49340
rect 121 49306 159 49335
rect 14 49301 159 49306
rect 193 49301 228 49335
rect 14 49276 228 49301
rect 14 49242 15 49276
rect 49 49272 228 49276
rect 49 49242 87 49272
rect 14 49238 87 49242
rect 121 49267 228 49272
rect 121 49238 159 49267
rect 14 49233 159 49238
rect 193 49233 228 49267
rect 14 49208 228 49233
rect 14 49174 15 49208
rect 49 49204 228 49208
rect 49 49174 87 49204
rect 14 49170 87 49174
rect 121 49199 228 49204
rect 121 49170 159 49199
rect 14 49165 159 49170
rect 193 49165 228 49199
rect 14 49140 228 49165
rect 14 49106 15 49140
rect 49 49136 228 49140
rect 49 49106 87 49136
rect 14 49102 87 49106
rect 121 49131 228 49136
rect 121 49102 159 49131
rect 14 49097 159 49102
rect 193 49097 228 49131
rect 14 49072 228 49097
rect 14 49038 15 49072
rect 49 49068 228 49072
rect 49 49038 87 49068
rect 14 49034 87 49038
rect 121 49063 228 49068
rect 121 49034 159 49063
rect 14 49029 159 49034
rect 193 49029 228 49063
rect 14 49004 228 49029
rect 14 48970 15 49004
rect 49 49000 228 49004
rect 49 48970 87 49000
rect 14 48966 87 48970
rect 121 48995 228 49000
rect 121 48966 159 48995
rect 14 48961 159 48966
rect 193 48961 228 48995
rect 14 48936 228 48961
rect 14 48902 15 48936
rect 49 48932 228 48936
rect 49 48902 87 48932
rect 14 48898 87 48902
rect 121 48927 228 48932
rect 121 48898 159 48927
rect 14 48893 159 48898
rect 193 48893 228 48927
rect 14 48868 228 48893
rect 14 48834 15 48868
rect 49 48864 228 48868
rect 49 48834 87 48864
rect 14 48830 87 48834
rect 121 48859 228 48864
rect 121 48830 159 48859
rect 14 48825 159 48830
rect 193 48825 228 48859
rect 14 48800 228 48825
rect 14 48766 15 48800
rect 49 48796 228 48800
rect 49 48766 87 48796
rect 14 48762 87 48766
rect 121 48791 228 48796
rect 121 48762 159 48791
rect 14 48757 159 48762
rect 193 48757 228 48791
rect 14 48732 228 48757
rect 14 48698 15 48732
rect 49 48728 228 48732
rect 49 48698 87 48728
rect 14 48694 87 48698
rect 121 48723 228 48728
rect 121 48694 159 48723
rect 14 48689 159 48694
rect 193 48689 228 48723
rect 14 48664 228 48689
rect 14 48630 15 48664
rect 49 48660 228 48664
rect 49 48630 87 48660
rect 14 48626 87 48630
rect 121 48655 228 48660
rect 121 48626 159 48655
rect 14 48621 159 48626
rect 193 48621 228 48655
rect 14 48596 228 48621
rect 14 48562 15 48596
rect 49 48592 228 48596
rect 49 48562 87 48592
rect 14 48558 87 48562
rect 121 48587 228 48592
rect 121 48558 159 48587
rect 14 48553 159 48558
rect 193 48553 228 48587
rect 14 48528 228 48553
rect 14 48494 15 48528
rect 49 48524 228 48528
rect 49 48494 87 48524
rect 14 48490 87 48494
rect 121 48519 228 48524
rect 121 48490 159 48519
rect 14 48485 159 48490
rect 193 48485 228 48519
rect 14 48460 228 48485
rect 14 48426 15 48460
rect 49 48456 228 48460
rect 49 48426 87 48456
rect 14 48422 87 48426
rect 121 48451 228 48456
rect 121 48422 159 48451
rect 14 48417 159 48422
rect 193 48417 228 48451
rect 14 48392 228 48417
rect 14 48358 15 48392
rect 49 48388 228 48392
rect 49 48358 87 48388
rect 14 48354 87 48358
rect 121 48383 228 48388
rect 121 48354 159 48383
rect 14 48349 159 48354
rect 193 48349 228 48383
rect 14 48324 228 48349
rect 14 48290 15 48324
rect 49 48320 228 48324
rect 49 48290 87 48320
rect 14 48286 87 48290
rect 121 48315 228 48320
rect 121 48286 159 48315
rect 14 48281 159 48286
rect 193 48281 228 48315
rect 14 48256 228 48281
rect 14 48222 15 48256
rect 49 48252 228 48256
rect 49 48222 87 48252
rect 14 48218 87 48222
rect 121 48247 228 48252
rect 121 48218 159 48247
rect 14 48213 159 48218
rect 193 48213 228 48247
rect 14 48188 228 48213
rect 14 48154 15 48188
rect 49 48184 228 48188
rect 49 48154 87 48184
rect 14 48150 87 48154
rect 121 48179 228 48184
rect 121 48150 159 48179
rect 14 48145 159 48150
rect 193 48145 228 48179
rect 14 48120 228 48145
rect 14 48086 15 48120
rect 49 48116 228 48120
rect 49 48086 87 48116
rect 14 48082 87 48086
rect 121 48111 228 48116
rect 121 48082 159 48111
rect 14 48077 159 48082
rect 193 48077 228 48111
rect 14 48052 228 48077
rect 14 48018 15 48052
rect 49 48048 228 48052
rect 49 48018 87 48048
rect 14 48014 87 48018
rect 121 48043 228 48048
rect 121 48014 159 48043
rect 14 48009 159 48014
rect 193 48009 228 48043
rect 14 47984 228 48009
rect 14 47950 15 47984
rect 49 47980 228 47984
rect 49 47950 87 47980
rect 14 47946 87 47950
rect 121 47975 228 47980
rect 121 47946 159 47975
rect 14 47941 159 47946
rect 193 47941 228 47975
rect 14 47916 228 47941
rect 14 47882 15 47916
rect 49 47912 228 47916
rect 49 47882 87 47912
rect 14 47878 87 47882
rect 121 47907 228 47912
rect 121 47878 159 47907
rect 14 47873 159 47878
rect 193 47873 228 47907
rect 14 47848 228 47873
rect 14 47814 15 47848
rect 49 47844 228 47848
rect 49 47814 87 47844
rect 14 47810 87 47814
rect 121 47839 228 47844
rect 121 47810 159 47839
rect 14 47805 159 47810
rect 193 47805 228 47839
rect 14 47780 228 47805
rect 14 47746 15 47780
rect 49 47776 228 47780
rect 49 47746 87 47776
rect 14 47742 87 47746
rect 121 47771 228 47776
rect 121 47742 159 47771
rect 14 47737 159 47742
rect 193 47737 228 47771
rect 14 47712 228 47737
rect 14 47678 15 47712
rect 49 47708 228 47712
rect 49 47678 87 47708
rect 14 47674 87 47678
rect 121 47703 228 47708
rect 121 47674 159 47703
rect 14 47669 159 47674
rect 193 47669 228 47703
rect 14 47644 228 47669
rect 14 47610 15 47644
rect 49 47640 228 47644
rect 49 47610 87 47640
rect 14 47606 87 47610
rect 121 47635 228 47640
rect 121 47606 159 47635
rect 14 47601 159 47606
rect 193 47601 228 47635
rect 14 47576 228 47601
rect 14 47542 15 47576
rect 49 47572 228 47576
rect 49 47542 87 47572
rect 14 47538 87 47542
rect 121 47567 228 47572
rect 121 47538 159 47567
rect 14 47533 159 47538
rect 193 47533 228 47567
rect 14 47508 228 47533
rect 14 47474 15 47508
rect 49 47504 228 47508
rect 49 47474 87 47504
rect 14 47470 87 47474
rect 121 47499 228 47504
rect 121 47470 159 47499
rect 14 47465 159 47470
rect 193 47465 228 47499
rect 14 47440 228 47465
rect 14 47406 15 47440
rect 49 47436 228 47440
rect 49 47406 87 47436
rect 14 47402 87 47406
rect 121 47431 228 47436
rect 121 47402 159 47431
rect 14 47397 159 47402
rect 193 47397 228 47431
rect 14 47372 228 47397
rect 14 47338 15 47372
rect 49 47368 228 47372
rect 49 47338 87 47368
rect 14 47334 87 47338
rect 121 47363 228 47368
rect 121 47334 159 47363
rect 14 47329 159 47334
rect 193 47329 228 47363
rect 14 47304 228 47329
rect 14 47270 15 47304
rect 49 47300 228 47304
rect 49 47270 87 47300
rect 14 47266 87 47270
rect 121 47295 228 47300
rect 121 47266 159 47295
rect 14 47261 159 47266
rect 193 47261 228 47295
rect 14 47236 228 47261
rect 14 47202 15 47236
rect 49 47232 228 47236
rect 49 47202 87 47232
rect 14 47198 87 47202
rect 121 47227 228 47232
rect 121 47198 159 47227
rect 14 47193 159 47198
rect 193 47193 228 47227
rect 14 47168 228 47193
rect 14 47134 15 47168
rect 49 47164 228 47168
rect 49 47134 87 47164
rect 14 47130 87 47134
rect 121 47159 228 47164
rect 121 47130 159 47159
rect 14 47125 159 47130
rect 193 47125 228 47159
rect 14 47100 228 47125
rect 14 47066 15 47100
rect 49 47096 228 47100
rect 49 47066 87 47096
rect 14 47062 87 47066
rect 121 47091 228 47096
rect 121 47062 159 47091
rect 14 47057 159 47062
rect 193 47057 228 47091
rect 14 47032 228 47057
rect 14 46998 15 47032
rect 49 47028 228 47032
rect 49 46998 87 47028
rect 14 46994 87 46998
rect 121 47023 228 47028
rect 121 46994 159 47023
rect 14 46989 159 46994
rect 193 46989 228 47023
rect 14 46964 228 46989
rect 14 46930 15 46964
rect 49 46960 228 46964
rect 49 46930 87 46960
rect 14 46926 87 46930
rect 121 46955 228 46960
rect 121 46926 159 46955
rect 14 46921 159 46926
rect 193 46921 228 46955
rect 14 46896 228 46921
rect 14 46862 15 46896
rect 49 46892 228 46896
rect 49 46862 87 46892
rect 14 46858 87 46862
rect 121 46887 228 46892
rect 121 46858 159 46887
rect 14 46853 159 46858
rect 193 46853 228 46887
rect 14 46828 228 46853
rect 14 46794 15 46828
rect 49 46824 228 46828
rect 49 46794 87 46824
rect 14 46790 87 46794
rect 121 46819 228 46824
rect 121 46790 159 46819
rect 14 46785 159 46790
rect 193 46785 228 46819
rect 14 46760 228 46785
rect 14 46726 15 46760
rect 49 46756 228 46760
rect 49 46726 87 46756
rect 14 46722 87 46726
rect 121 46751 228 46756
rect 121 46722 159 46751
rect 14 46717 159 46722
rect 193 46717 228 46751
rect 14 46692 228 46717
rect 14 46658 15 46692
rect 49 46688 228 46692
rect 49 46658 87 46688
rect 14 46654 87 46658
rect 121 46683 228 46688
rect 121 46654 159 46683
rect 14 46649 159 46654
rect 193 46649 228 46683
rect 14 46624 228 46649
rect 14 46590 15 46624
rect 49 46620 228 46624
rect 49 46590 87 46620
rect 14 46586 87 46590
rect 121 46615 228 46620
rect 121 46586 159 46615
rect 14 46581 159 46586
rect 193 46581 228 46615
rect 14 46556 228 46581
rect 14 46522 15 46556
rect 49 46552 228 46556
rect 49 46522 87 46552
rect 14 46518 87 46522
rect 121 46547 228 46552
rect 121 46518 159 46547
rect 14 46513 159 46518
rect 193 46513 228 46547
rect 14 46488 228 46513
rect 14 46454 15 46488
rect 49 46484 228 46488
rect 49 46454 87 46484
rect 14 46450 87 46454
rect 121 46479 228 46484
rect 121 46450 159 46479
rect 14 46445 159 46450
rect 193 46445 228 46479
rect 14 46420 228 46445
rect 14 46386 15 46420
rect 49 46416 228 46420
rect 49 46386 87 46416
rect 14 46382 87 46386
rect 121 46411 228 46416
rect 121 46382 159 46411
rect 14 46377 159 46382
rect 193 46377 228 46411
rect 14 46352 228 46377
rect 14 46318 15 46352
rect 49 46348 228 46352
rect 49 46318 87 46348
rect 14 46314 87 46318
rect 121 46343 228 46348
rect 121 46314 159 46343
rect 14 46309 159 46314
rect 193 46309 228 46343
rect 14 46284 228 46309
rect 14 46250 15 46284
rect 49 46280 228 46284
rect 49 46250 87 46280
rect 14 46246 87 46250
rect 121 46275 228 46280
rect 121 46246 159 46275
rect 14 46241 159 46246
rect 193 46241 228 46275
rect 14 46216 228 46241
rect 14 46182 15 46216
rect 49 46212 228 46216
rect 49 46182 87 46212
rect 14 46178 87 46182
rect 121 46207 228 46212
rect 121 46178 159 46207
rect 14 46173 159 46178
rect 193 46173 228 46207
rect 14 46148 228 46173
rect 14 46114 15 46148
rect 49 46144 228 46148
rect 49 46114 87 46144
rect 14 46110 87 46114
rect 121 46139 228 46144
rect 121 46110 159 46139
rect 14 46105 159 46110
rect 193 46105 228 46139
rect 14 46080 228 46105
rect 14 46046 15 46080
rect 49 46076 228 46080
rect 49 46046 87 46076
rect 14 46042 87 46046
rect 121 46071 228 46076
rect 121 46042 159 46071
rect 14 46037 159 46042
rect 193 46037 228 46071
rect 14 46012 228 46037
rect 14 45978 15 46012
rect 49 46008 228 46012
rect 49 45978 87 46008
rect 14 45974 87 45978
rect 121 46003 228 46008
rect 121 45974 159 46003
rect 14 45969 159 45974
rect 193 45969 228 46003
rect 14 45944 228 45969
rect 14 45910 15 45944
rect 49 45940 228 45944
rect 49 45910 87 45940
rect 14 45906 87 45910
rect 121 45935 228 45940
rect 121 45906 159 45935
rect 14 45901 159 45906
rect 193 45901 228 45935
rect 14 45876 228 45901
rect 14 45842 15 45876
rect 49 45872 228 45876
rect 49 45842 87 45872
rect 14 45838 87 45842
rect 121 45867 228 45872
rect 121 45838 159 45867
rect 14 45833 159 45838
rect 193 45833 228 45867
rect 14 45808 228 45833
rect 14 45774 15 45808
rect 49 45804 228 45808
rect 49 45774 87 45804
rect 14 45770 87 45774
rect 121 45799 228 45804
rect 121 45770 159 45799
rect 14 45765 159 45770
rect 193 45765 228 45799
rect 14 45740 228 45765
rect 14 45706 15 45740
rect 49 45736 228 45740
rect 49 45706 87 45736
rect 14 45702 87 45706
rect 121 45731 228 45736
rect 121 45702 159 45731
rect 14 45697 159 45702
rect 193 45697 228 45731
rect 14 45672 228 45697
rect 14 45638 15 45672
rect 49 45668 228 45672
rect 49 45638 87 45668
rect 14 45634 87 45638
rect 121 45663 228 45668
rect 121 45634 159 45663
rect 14 45629 159 45634
rect 193 45629 228 45663
rect 14 45604 228 45629
rect 14 45570 15 45604
rect 49 45600 228 45604
rect 49 45570 87 45600
rect 14 45566 87 45570
rect 121 45595 228 45600
rect 121 45566 159 45595
rect 14 45561 159 45566
rect 193 45561 228 45595
rect 14 45536 228 45561
rect 14 45502 15 45536
rect 49 45532 228 45536
rect 49 45502 87 45532
rect 14 45498 87 45502
rect 121 45527 228 45532
rect 121 45498 159 45527
rect 14 45493 159 45498
rect 193 45493 228 45527
rect 14 45468 228 45493
rect 14 45434 15 45468
rect 49 45464 228 45468
rect 49 45434 87 45464
rect 14 45430 87 45434
rect 121 45459 228 45464
rect 121 45430 159 45459
rect 14 45425 159 45430
rect 193 45425 228 45459
rect 14 45400 228 45425
rect 14 45366 15 45400
rect 49 45396 228 45400
rect 49 45366 87 45396
rect 14 45362 87 45366
rect 121 45391 228 45396
rect 121 45362 159 45391
rect 14 45357 159 45362
rect 193 45357 228 45391
rect 14 45332 228 45357
rect 14 45298 15 45332
rect 49 45328 228 45332
rect 49 45298 87 45328
rect 14 45294 87 45298
rect 121 45323 228 45328
rect 121 45294 159 45323
rect 14 45289 159 45294
rect 193 45289 228 45323
rect 14 45264 228 45289
rect 14 45230 15 45264
rect 49 45260 228 45264
rect 49 45230 87 45260
rect 14 45226 87 45230
rect 121 45255 228 45260
rect 121 45226 159 45255
rect 14 45221 159 45226
rect 193 45221 228 45255
rect 14 45196 228 45221
rect 14 45162 15 45196
rect 49 45192 228 45196
rect 49 45162 87 45192
rect 14 45158 87 45162
rect 121 45187 228 45192
rect 121 45158 159 45187
rect 14 45153 159 45158
rect 193 45153 228 45187
rect 14 45128 228 45153
rect 14 45094 15 45128
rect 49 45124 228 45128
rect 49 45094 87 45124
rect 14 45090 87 45094
rect 121 45119 228 45124
rect 121 45090 159 45119
rect 14 45085 159 45090
rect 193 45085 228 45119
rect 14 45060 228 45085
rect 14 45026 15 45060
rect 49 45056 228 45060
rect 49 45026 87 45056
rect 14 45022 87 45026
rect 121 45051 228 45056
rect 121 45022 159 45051
rect 14 45017 159 45022
rect 193 45017 228 45051
rect 14 44992 228 45017
rect 14 44958 15 44992
rect 49 44988 228 44992
rect 49 44958 87 44988
rect 14 44954 87 44958
rect 121 44983 228 44988
rect 121 44954 159 44983
rect 14 44949 159 44954
rect 193 44949 228 44983
rect 14 44924 228 44949
rect 14 44890 15 44924
rect 49 44920 228 44924
rect 49 44890 87 44920
rect 14 44886 87 44890
rect 121 44915 228 44920
rect 121 44886 159 44915
rect 14 44881 159 44886
rect 193 44881 228 44915
rect 14 44856 228 44881
rect 14 44822 15 44856
rect 49 44852 228 44856
rect 49 44822 87 44852
rect 14 44818 87 44822
rect 121 44847 228 44852
rect 121 44818 159 44847
rect 14 44813 159 44818
rect 193 44813 228 44847
rect 14 44788 228 44813
rect 14 44754 15 44788
rect 49 44784 228 44788
rect 49 44754 87 44784
rect 14 44750 87 44754
rect 121 44779 228 44784
rect 121 44750 159 44779
rect 14 44745 159 44750
rect 193 44745 228 44779
rect 14 44720 228 44745
rect 14 44686 15 44720
rect 49 44716 228 44720
rect 49 44686 87 44716
rect 14 44682 87 44686
rect 121 44711 228 44716
rect 121 44682 159 44711
rect 14 44677 159 44682
rect 193 44677 228 44711
rect 14 44652 228 44677
rect 14 44618 15 44652
rect 49 44648 228 44652
rect 49 44618 87 44648
rect 14 44614 87 44618
rect 121 44643 228 44648
rect 121 44614 159 44643
rect 14 44609 159 44614
rect 193 44609 228 44643
rect 14 44584 228 44609
rect 14 44550 15 44584
rect 49 44580 228 44584
rect 49 44550 87 44580
rect 14 44546 87 44550
rect 121 44575 228 44580
rect 121 44546 159 44575
rect 14 44541 159 44546
rect 193 44541 228 44575
rect 14 44516 228 44541
rect 14 44482 15 44516
rect 49 44512 228 44516
rect 49 44482 87 44512
rect 14 44478 87 44482
rect 121 44507 228 44512
rect 121 44478 159 44507
rect 14 44473 159 44478
rect 193 44473 228 44507
rect 14 44448 228 44473
rect 14 44414 15 44448
rect 49 44444 228 44448
rect 49 44414 87 44444
rect 14 44410 87 44414
rect 121 44439 228 44444
rect 121 44410 159 44439
rect 14 44405 159 44410
rect 193 44405 228 44439
rect 14 44380 228 44405
rect 14 44346 15 44380
rect 49 44376 228 44380
rect 49 44346 87 44376
rect 14 44342 87 44346
rect 121 44371 228 44376
rect 121 44342 159 44371
rect 14 44337 159 44342
rect 193 44337 228 44371
rect 14 44312 228 44337
rect 14 44278 15 44312
rect 49 44308 228 44312
rect 49 44278 87 44308
rect 14 44274 87 44278
rect 121 44303 228 44308
rect 121 44274 159 44303
rect 14 44269 159 44274
rect 193 44269 228 44303
rect 14 44244 228 44269
rect 14 44210 15 44244
rect 49 44240 228 44244
rect 49 44210 87 44240
rect 14 44206 87 44210
rect 121 44235 228 44240
rect 121 44206 159 44235
rect 14 44201 159 44206
rect 193 44201 228 44235
rect 14 44176 228 44201
rect 14 44142 15 44176
rect 49 44172 228 44176
rect 49 44142 87 44172
rect 14 44138 87 44142
rect 121 44167 228 44172
rect 121 44138 159 44167
rect 14 44133 159 44138
rect 193 44133 228 44167
rect 14 44108 228 44133
rect 14 44074 15 44108
rect 49 44104 228 44108
rect 49 44074 87 44104
rect 14 44070 87 44074
rect 121 44099 228 44104
rect 121 44070 159 44099
rect 14 44065 159 44070
rect 193 44065 228 44099
rect 14 44040 228 44065
rect 14 44006 15 44040
rect 49 44036 228 44040
rect 49 44006 87 44036
rect 14 44002 87 44006
rect 121 44031 228 44036
rect 121 44002 159 44031
rect 14 43997 159 44002
rect 193 43997 228 44031
rect 14 43972 228 43997
rect 14 43938 15 43972
rect 49 43968 228 43972
rect 49 43938 87 43968
rect 14 43934 87 43938
rect 121 43963 228 43968
rect 121 43934 159 43963
rect 14 43929 159 43934
rect 193 43929 228 43963
rect 14 43904 228 43929
rect 14 43870 15 43904
rect 49 43900 228 43904
rect 49 43870 87 43900
rect 14 43866 87 43870
rect 121 43895 228 43900
rect 121 43866 159 43895
rect 14 43861 159 43866
rect 193 43861 228 43895
rect 14 43836 228 43861
rect 14 43802 15 43836
rect 49 43832 228 43836
rect 49 43802 87 43832
rect 14 43798 87 43802
rect 121 43827 228 43832
rect 121 43798 159 43827
rect 14 43793 159 43798
rect 193 43793 228 43827
rect 14 43768 228 43793
rect 14 43734 15 43768
rect 49 43764 228 43768
rect 49 43734 87 43764
rect 14 43730 87 43734
rect 121 43759 228 43764
rect 121 43730 159 43759
rect 14 43725 159 43730
rect 193 43725 228 43759
rect 14 43700 228 43725
rect 14 43666 15 43700
rect 49 43696 228 43700
rect 49 43666 87 43696
rect 14 43662 87 43666
rect 121 43691 228 43696
rect 121 43662 159 43691
rect 14 43657 159 43662
rect 193 43657 228 43691
rect 14 43632 228 43657
rect 14 43598 15 43632
rect 49 43628 228 43632
rect 49 43598 87 43628
rect 14 43594 87 43598
rect 121 43623 228 43628
rect 121 43594 159 43623
rect 14 43589 159 43594
rect 193 43589 228 43623
rect 14 43564 228 43589
rect 14 43530 15 43564
rect 49 43560 228 43564
rect 49 43530 87 43560
rect 14 43526 87 43530
rect 121 43555 228 43560
rect 121 43526 159 43555
rect 14 43521 159 43526
rect 193 43521 228 43555
rect 14 43496 228 43521
rect 14 43462 15 43496
rect 49 43492 228 43496
rect 49 43462 87 43492
rect 14 43458 87 43462
rect 121 43487 228 43492
rect 121 43458 159 43487
rect 14 43453 159 43458
rect 193 43453 228 43487
rect 14 43428 228 43453
rect 14 43394 15 43428
rect 49 43424 228 43428
rect 49 43394 87 43424
rect 14 43390 87 43394
rect 121 43419 228 43424
rect 121 43390 159 43419
rect 14 43385 159 43390
rect 193 43385 228 43419
rect 14 43360 228 43385
rect 14 43326 15 43360
rect 49 43356 228 43360
rect 49 43326 87 43356
rect 14 43322 87 43326
rect 121 43351 228 43356
rect 121 43322 159 43351
rect 14 43317 159 43322
rect 193 43317 228 43351
rect 14 43292 228 43317
rect 14 43258 15 43292
rect 49 43288 228 43292
rect 49 43258 87 43288
rect 14 43254 87 43258
rect 121 43283 228 43288
rect 121 43254 159 43283
rect 14 43249 159 43254
rect 193 43249 228 43283
rect 14 43224 228 43249
rect 14 43190 15 43224
rect 49 43220 228 43224
rect 49 43190 87 43220
rect 14 43186 87 43190
rect 121 43215 228 43220
rect 121 43186 159 43215
rect 14 43181 159 43186
rect 193 43181 228 43215
rect 14 43156 228 43181
rect 14 43122 15 43156
rect 49 43152 228 43156
rect 49 43122 87 43152
rect 14 43118 87 43122
rect 121 43147 228 43152
rect 121 43118 159 43147
rect 14 43113 159 43118
rect 193 43113 228 43147
rect 14 43088 228 43113
rect 14 43054 15 43088
rect 49 43084 228 43088
rect 49 43054 87 43084
rect 14 43050 87 43054
rect 121 43079 228 43084
rect 121 43050 159 43079
rect 14 43045 159 43050
rect 193 43045 228 43079
rect 14 43020 228 43045
rect 14 42986 15 43020
rect 49 43016 228 43020
rect 49 42986 87 43016
rect 14 42982 87 42986
rect 121 43011 228 43016
rect 121 42982 159 43011
rect 14 42977 159 42982
rect 193 42977 228 43011
rect 14 42952 228 42977
rect 14 42918 15 42952
rect 49 42948 228 42952
rect 49 42918 87 42948
rect 14 42914 87 42918
rect 121 42943 228 42948
rect 121 42914 159 42943
rect 14 42909 159 42914
rect 193 42909 228 42943
rect 14 42884 228 42909
rect 14 42850 15 42884
rect 49 42880 228 42884
rect 49 42850 87 42880
rect 14 42846 87 42850
rect 121 42875 228 42880
rect 121 42846 159 42875
rect 14 42841 159 42846
rect 193 42841 228 42875
rect 14 42816 228 42841
rect 14 42782 15 42816
rect 49 42812 228 42816
rect 49 42782 87 42812
rect 14 42778 87 42782
rect 121 42807 228 42812
rect 121 42778 159 42807
rect 14 42773 159 42778
rect 193 42773 228 42807
rect 14 42748 228 42773
rect 14 42714 15 42748
rect 49 42744 228 42748
rect 49 42714 87 42744
rect 14 42710 87 42714
rect 121 42739 228 42744
rect 121 42710 159 42739
rect 14 42705 159 42710
rect 193 42705 228 42739
rect 14 42680 228 42705
rect 14 42646 15 42680
rect 49 42676 228 42680
rect 49 42646 87 42676
rect 14 42642 87 42646
rect 121 42671 228 42676
rect 121 42642 159 42671
rect 14 42637 159 42642
rect 193 42637 228 42671
rect 14 42612 228 42637
rect 14 42578 15 42612
rect 49 42608 228 42612
rect 49 42578 87 42608
rect 14 42574 87 42578
rect 121 42603 228 42608
rect 121 42574 159 42603
rect 14 42569 159 42574
rect 193 42569 228 42603
rect 14 42544 228 42569
rect 14 42510 15 42544
rect 49 42540 228 42544
rect 49 42510 87 42540
rect 14 42506 87 42510
rect 121 42535 228 42540
rect 121 42506 159 42535
rect 14 42501 159 42506
rect 193 42501 228 42535
rect 14 42476 228 42501
rect 14 42442 15 42476
rect 49 42472 228 42476
rect 49 42442 87 42472
rect 14 42438 87 42442
rect 121 42467 228 42472
rect 121 42438 159 42467
rect 14 42433 159 42438
rect 193 42433 228 42467
rect 14 42408 228 42433
rect 14 42374 15 42408
rect 49 42404 228 42408
rect 49 42374 87 42404
rect 14 42370 87 42374
rect 121 42399 228 42404
rect 121 42370 159 42399
rect 14 42365 159 42370
rect 193 42365 228 42399
rect 14 42340 228 42365
rect 14 42306 15 42340
rect 49 42336 228 42340
rect 49 42306 87 42336
rect 14 42302 87 42306
rect 121 42331 228 42336
rect 121 42302 159 42331
rect 14 42297 159 42302
rect 193 42297 228 42331
rect 14 42272 228 42297
rect 14 42238 15 42272
rect 49 42268 228 42272
rect 49 42238 87 42268
rect 14 42234 87 42238
rect 121 42263 228 42268
rect 121 42234 159 42263
rect 14 42229 159 42234
rect 193 42229 228 42263
rect 14 42204 228 42229
rect 14 42170 15 42204
rect 49 42200 228 42204
rect 49 42170 87 42200
rect 14 42166 87 42170
rect 121 42195 228 42200
rect 121 42166 159 42195
rect 14 42161 159 42166
rect 193 42161 228 42195
rect 14 42136 228 42161
rect 14 42102 15 42136
rect 49 42132 228 42136
rect 49 42102 87 42132
rect 14 42098 87 42102
rect 121 42127 228 42132
rect 121 42098 159 42127
rect 14 42093 159 42098
rect 193 42093 228 42127
rect 14 42068 228 42093
rect 14 42034 15 42068
rect 49 42064 228 42068
rect 49 42034 87 42064
rect 14 42030 87 42034
rect 121 42059 228 42064
rect 121 42030 159 42059
rect 14 42025 159 42030
rect 193 42025 228 42059
rect 14 42000 228 42025
rect 14 41966 15 42000
rect 49 41996 228 42000
rect 49 41966 87 41996
rect 14 41962 87 41966
rect 121 41991 228 41996
rect 121 41962 159 41991
rect 14 41957 159 41962
rect 193 41957 228 41991
rect 14 41932 228 41957
rect 14 41898 15 41932
rect 49 41928 228 41932
rect 49 41898 87 41928
rect 14 41894 87 41898
rect 121 41923 228 41928
rect 121 41894 159 41923
rect 14 41889 159 41894
rect 193 41889 228 41923
rect 14 41864 228 41889
rect 14 41830 15 41864
rect 49 41860 228 41864
rect 49 41830 87 41860
rect 14 41826 87 41830
rect 121 41855 228 41860
rect 121 41826 159 41855
rect 14 41821 159 41826
rect 193 41821 228 41855
rect 14 41796 228 41821
rect 14 41762 15 41796
rect 49 41792 228 41796
rect 49 41762 87 41792
rect 14 41758 87 41762
rect 121 41787 228 41792
rect 121 41758 159 41787
rect 14 41753 159 41758
rect 193 41753 228 41787
rect 14 41728 228 41753
rect 14 41694 15 41728
rect 49 41724 228 41728
rect 49 41694 87 41724
rect 14 41690 87 41694
rect 121 41719 228 41724
rect 121 41690 159 41719
rect 14 41685 159 41690
rect 193 41685 228 41719
rect 14 41660 228 41685
rect 14 41626 15 41660
rect 49 41656 228 41660
rect 49 41626 87 41656
rect 14 41622 87 41626
rect 121 41651 228 41656
rect 121 41622 159 41651
rect 14 41617 159 41622
rect 193 41617 228 41651
rect 14 41592 228 41617
rect 14 41558 15 41592
rect 49 41588 228 41592
rect 49 41558 87 41588
rect 14 41554 87 41558
rect 121 41583 228 41588
rect 121 41554 159 41583
rect 14 41549 159 41554
rect 193 41549 228 41583
rect 14 41524 228 41549
rect 14 41490 15 41524
rect 49 41520 228 41524
rect 49 41490 87 41520
rect 14 41486 87 41490
rect 121 41515 228 41520
rect 121 41486 159 41515
rect 14 41481 159 41486
rect 193 41481 228 41515
rect 14 41456 228 41481
rect 14 41422 15 41456
rect 49 41452 228 41456
rect 49 41422 87 41452
rect 14 41418 87 41422
rect 121 41447 228 41452
rect 121 41418 159 41447
rect 14 41413 159 41418
rect 193 41413 228 41447
rect 14 41388 228 41413
rect 14 41354 15 41388
rect 49 41384 228 41388
rect 49 41354 87 41384
rect 14 41350 87 41354
rect 121 41379 228 41384
rect 121 41350 159 41379
rect 14 41345 159 41350
rect 193 41345 228 41379
rect 14 41320 228 41345
rect 14 41286 15 41320
rect 49 41316 228 41320
rect 49 41286 87 41316
rect 14 41282 87 41286
rect 121 41311 228 41316
rect 121 41282 159 41311
rect 14 41277 159 41282
rect 193 41277 228 41311
rect 14 41252 228 41277
rect 14 41218 15 41252
rect 49 41248 228 41252
rect 49 41218 87 41248
rect 14 41214 87 41218
rect 121 41243 228 41248
rect 121 41214 159 41243
rect 14 41209 159 41214
rect 193 41209 228 41243
rect 14 41184 228 41209
rect 14 41150 15 41184
rect 49 41180 228 41184
rect 49 41150 87 41180
rect 14 41146 87 41150
rect 121 41175 228 41180
rect 121 41146 159 41175
rect 14 41141 159 41146
rect 193 41141 228 41175
rect 14 41116 228 41141
rect 14 41082 15 41116
rect 49 41112 228 41116
rect 49 41082 87 41112
rect 14 41078 87 41082
rect 121 41107 228 41112
rect 121 41078 159 41107
rect 14 41073 159 41078
rect 193 41073 228 41107
rect 14 41048 228 41073
rect 14 41014 15 41048
rect 49 41044 228 41048
rect 49 41014 87 41044
rect 14 41010 87 41014
rect 121 41039 228 41044
rect 121 41010 159 41039
rect 14 41005 159 41010
rect 193 41005 228 41039
rect 14 40980 228 41005
rect 14 40946 15 40980
rect 49 40976 228 40980
rect 49 40946 87 40976
rect 14 40942 87 40946
rect 121 40971 228 40976
rect 121 40942 159 40971
rect 14 40937 159 40942
rect 193 40937 228 40971
rect 14 40912 228 40937
rect 14 40878 15 40912
rect 49 40908 228 40912
rect 49 40878 87 40908
rect 14 40874 87 40878
rect 121 40903 228 40908
rect 121 40874 159 40903
rect 14 40869 159 40874
rect 193 40869 228 40903
rect 14 40844 228 40869
rect 14 40810 15 40844
rect 49 40840 228 40844
rect 49 40810 87 40840
rect 14 40806 87 40810
rect 121 40835 228 40840
rect 121 40806 159 40835
rect 14 40801 159 40806
rect 193 40801 228 40835
rect 14 40776 228 40801
rect 14 40742 15 40776
rect 49 40772 228 40776
rect 49 40742 87 40772
rect 14 40738 87 40742
rect 121 40767 228 40772
rect 121 40738 159 40767
rect 14 40733 159 40738
rect 193 40733 228 40767
rect 14 40708 228 40733
rect 14 40674 15 40708
rect 49 40704 228 40708
rect 49 40674 87 40704
rect 14 40670 87 40674
rect 121 40699 228 40704
rect 121 40670 159 40699
rect 14 40665 159 40670
rect 193 40665 228 40699
rect 14 40640 228 40665
rect 14 40606 15 40640
rect 49 40636 228 40640
rect 49 40606 87 40636
rect 14 40602 87 40606
rect 121 40631 228 40636
rect 121 40602 159 40631
rect 14 40597 159 40602
rect 193 40597 228 40631
rect 14 40572 228 40597
rect 14 40538 15 40572
rect 49 40568 228 40572
rect 49 40538 87 40568
rect 14 40534 87 40538
rect 121 40563 228 40568
rect 121 40534 159 40563
rect 14 40529 159 40534
rect 193 40529 228 40563
rect 14 40504 228 40529
rect 14 40470 15 40504
rect 49 40500 228 40504
rect 49 40470 87 40500
rect 14 40466 87 40470
rect 121 40495 228 40500
rect 121 40466 159 40495
rect 14 40461 159 40466
rect 193 40461 228 40495
rect 14 40436 228 40461
rect 14 40402 15 40436
rect 49 40432 228 40436
rect 49 40402 87 40432
rect 14 40398 87 40402
rect 121 40427 228 40432
rect 121 40398 159 40427
rect 14 40393 159 40398
rect 193 40393 228 40427
rect 14 40368 228 40393
rect 14 40334 15 40368
rect 49 40364 228 40368
rect 49 40334 87 40364
rect 14 40330 87 40334
rect 121 40359 228 40364
rect 121 40330 159 40359
rect 14 40325 159 40330
rect 193 40325 228 40359
rect 14 40300 228 40325
rect 14 40266 15 40300
rect 49 40296 228 40300
rect 49 40266 87 40296
rect 14 40262 87 40266
rect 121 40291 228 40296
rect 121 40262 159 40291
rect 14 40257 159 40262
rect 193 40257 228 40291
rect 14 40232 228 40257
rect 14 40198 15 40232
rect 49 40228 228 40232
rect 49 40198 87 40228
rect 14 40194 87 40198
rect 121 40223 228 40228
rect 121 40194 159 40223
rect 14 40189 159 40194
rect 193 40189 228 40223
rect 14 40164 228 40189
rect 14 40130 15 40164
rect 49 40160 228 40164
rect 49 40130 87 40160
rect 14 40126 87 40130
rect 121 40155 228 40160
rect 121 40126 159 40155
rect 14 40121 159 40126
rect 193 40121 228 40155
rect 14 40096 228 40121
rect 14 40062 15 40096
rect 49 40092 228 40096
rect 49 40062 87 40092
rect 14 40058 87 40062
rect 121 40087 228 40092
rect 121 40058 159 40087
rect 14 40053 159 40058
rect 193 40053 228 40087
rect 14 40028 228 40053
rect 14 39994 15 40028
rect 49 40024 228 40028
rect 49 39994 87 40024
rect 14 39990 87 39994
rect 121 40019 228 40024
rect 121 39990 159 40019
rect 14 39985 159 39990
rect 193 39985 228 40019
rect 14 39960 228 39985
rect 14 39926 15 39960
rect 49 39956 228 39960
rect 49 39926 87 39956
rect 14 39922 87 39926
rect 121 39951 228 39956
rect 121 39922 159 39951
rect 14 39917 159 39922
rect 193 39917 228 39951
rect 14 39892 228 39917
rect 14 39858 15 39892
rect 49 39888 228 39892
rect 49 39858 87 39888
rect 14 39854 87 39858
rect 121 39883 228 39888
rect 121 39854 159 39883
rect 14 39849 159 39854
rect 193 39849 228 39883
rect 14 39824 228 39849
rect 14 39790 15 39824
rect 49 39820 228 39824
rect 49 39790 87 39820
rect 14 39786 87 39790
rect 121 39815 228 39820
rect 121 39786 159 39815
rect 14 39781 159 39786
rect 193 39781 228 39815
rect 14 39756 228 39781
rect 14 39722 15 39756
rect 49 39752 228 39756
rect 49 39722 87 39752
rect 14 39718 87 39722
rect 121 39747 228 39752
rect 121 39718 159 39747
rect 14 39713 159 39718
rect 193 39713 228 39747
rect 14 39688 228 39713
rect 14 39654 15 39688
rect 49 39684 228 39688
rect 49 39654 87 39684
rect 14 39650 87 39654
rect 121 39679 228 39684
rect 121 39650 159 39679
rect 14 39645 159 39650
rect 193 39645 228 39679
rect 14 39620 228 39645
rect 14 39586 15 39620
rect 49 39616 228 39620
rect 49 39586 87 39616
rect 14 39582 87 39586
rect 121 39611 228 39616
rect 121 39582 159 39611
rect 14 39577 159 39582
rect 193 39577 228 39611
rect 14 39552 228 39577
rect 14 39518 15 39552
rect 49 39548 228 39552
rect 49 39518 87 39548
rect 14 39514 87 39518
rect 121 39543 228 39548
rect 121 39514 159 39543
rect 14 39509 159 39514
rect 193 39509 228 39543
rect 14 39484 228 39509
rect 14 39450 15 39484
rect 49 39480 228 39484
rect 49 39450 87 39480
rect 14 39446 87 39450
rect 121 39475 228 39480
rect 121 39446 159 39475
rect 14 39441 159 39446
rect 193 39441 228 39475
rect 14 39416 228 39441
rect 14 39382 15 39416
rect 49 39412 228 39416
rect 49 39382 87 39412
rect 14 39378 87 39382
rect 121 39407 228 39412
rect 121 39378 159 39407
rect 14 39373 159 39378
rect 193 39373 228 39407
rect 14 39348 228 39373
rect 14 39314 15 39348
rect 49 39344 228 39348
rect 49 39314 87 39344
rect 14 39310 87 39314
rect 121 39339 228 39344
rect 121 39310 159 39339
rect 14 39305 159 39310
rect 193 39305 228 39339
rect 14 39280 228 39305
rect 14 39246 15 39280
rect 49 39276 228 39280
rect 49 39246 87 39276
rect 14 39242 87 39246
rect 121 39271 228 39276
rect 121 39242 159 39271
rect 14 39237 159 39242
rect 193 39237 228 39271
rect 14 39212 228 39237
rect 14 39178 15 39212
rect 49 39208 228 39212
rect 49 39178 87 39208
rect 14 39174 87 39178
rect 121 39203 228 39208
rect 121 39174 159 39203
rect 14 39169 159 39174
rect 193 39169 228 39203
rect 14 39144 228 39169
rect 14 39110 15 39144
rect 49 39140 228 39144
rect 49 39110 87 39140
rect 14 39106 87 39110
rect 121 39135 228 39140
rect 121 39106 159 39135
rect 14 39101 159 39106
rect 193 39101 228 39135
rect 14 39076 228 39101
rect 14 39042 15 39076
rect 49 39072 228 39076
rect 49 39042 87 39072
rect 14 39038 87 39042
rect 121 39067 228 39072
rect 121 39038 159 39067
rect 14 39033 159 39038
rect 193 39033 228 39067
rect 14 39008 228 39033
rect 14 38974 15 39008
rect 49 39004 228 39008
rect 49 38974 87 39004
rect 14 38970 87 38974
rect 121 38999 228 39004
rect 121 38970 159 38999
rect 14 38965 159 38970
rect 193 38965 228 38999
rect 14 38940 228 38965
rect 14 38906 15 38940
rect 49 38936 228 38940
rect 49 38906 87 38936
rect 14 38902 87 38906
rect 121 38931 228 38936
rect 121 38902 159 38931
rect 14 38897 159 38902
rect 193 38897 228 38931
rect 14 38872 228 38897
rect 14 38838 15 38872
rect 49 38868 228 38872
rect 49 38838 87 38868
rect 14 38834 87 38838
rect 121 38863 228 38868
rect 121 38834 159 38863
rect 14 38829 159 38834
rect 193 38861 228 38863
rect 193 38829 194 38861
rect 14 38804 194 38829
rect 14 38770 15 38804
rect 49 38800 194 38804
rect 49 38770 87 38800
rect 14 38766 87 38770
rect 121 38795 194 38800
rect 121 38766 159 38795
rect 14 38761 159 38766
rect 193 38761 194 38795
rect 14 38736 194 38761
rect 14 38702 15 38736
rect 49 38732 194 38736
rect 49 38702 87 38732
rect 14 38698 87 38702
rect 121 38727 194 38732
rect 121 38698 159 38727
rect 14 38693 159 38698
rect 193 38693 194 38727
rect 14 38668 194 38693
rect 14 38634 15 38668
rect 49 38664 194 38668
rect 49 38634 87 38664
rect 14 38630 87 38634
rect 121 38659 194 38664
rect 121 38630 159 38659
rect 14 38625 159 38630
rect 193 38625 194 38659
rect 14 38600 194 38625
rect 14 38566 15 38600
rect 49 38596 194 38600
rect 49 38566 87 38596
rect 14 38562 87 38566
rect 121 38591 194 38596
rect 121 38562 159 38591
rect 14 38557 159 38562
rect 193 38557 194 38591
rect 14 38532 194 38557
rect 14 38498 15 38532
rect 49 38528 194 38532
rect 49 38498 87 38528
rect 14 38494 87 38498
rect 121 38523 194 38528
rect 121 38494 159 38523
rect 14 38489 159 38494
rect 193 38489 194 38523
rect 14 38464 194 38489
rect 14 38430 15 38464
rect 49 38460 194 38464
rect 49 38430 87 38460
rect 14 38426 87 38430
rect 121 38455 194 38460
rect 121 38426 159 38455
rect 14 38421 159 38426
rect 193 38421 194 38455
rect 14 38396 194 38421
rect 14 38362 15 38396
rect 49 38392 194 38396
rect 49 38362 87 38392
rect 14 38358 87 38362
rect 121 38387 194 38392
rect 121 38358 159 38387
rect 14 38353 159 38358
rect 193 38353 194 38387
rect 14 38328 194 38353
rect 14 38294 15 38328
rect 49 38324 194 38328
rect 49 38294 87 38324
rect 14 38290 87 38294
rect 121 38319 194 38324
rect 121 38290 159 38319
rect 14 38285 159 38290
rect 193 38285 194 38319
rect 14 38260 194 38285
rect 14 38226 15 38260
rect 49 38256 194 38260
rect 49 38226 87 38256
rect 14 38222 87 38226
rect 121 38251 194 38256
rect 121 38222 159 38251
rect 14 38217 159 38222
rect 193 38217 194 38251
rect 14 38192 194 38217
rect 14 38158 15 38192
rect 49 38188 194 38192
rect 49 38158 87 38188
rect 14 38154 87 38158
rect 121 38183 194 38188
rect 121 38154 159 38183
rect 14 38149 159 38154
rect 193 38149 194 38183
rect 14 38124 194 38149
rect 14 38090 15 38124
rect 49 38120 194 38124
rect 49 38090 87 38120
rect 14 38086 87 38090
rect 121 38115 194 38120
rect 121 38086 159 38115
rect 14 38081 159 38086
rect 193 38081 194 38115
rect 14 38056 194 38081
rect 14 38022 15 38056
rect 49 38052 194 38056
rect 49 38022 87 38052
rect 14 38018 87 38022
rect 121 38047 194 38052
rect 121 38018 159 38047
rect 14 38013 159 38018
rect 193 38013 194 38047
rect 14 37988 194 38013
rect 14 37954 15 37988
rect 49 37984 194 37988
rect 49 37954 87 37984
rect 14 37950 87 37954
rect 121 37979 194 37984
rect 121 37950 159 37979
rect 14 37945 159 37950
rect 193 37945 194 37979
rect 14 37920 194 37945
rect 14 37886 15 37920
rect 49 37916 194 37920
rect 49 37886 87 37916
rect 14 37882 87 37886
rect 121 37911 194 37916
rect 121 37882 159 37911
rect 14 37877 159 37882
rect 193 37877 194 37911
rect 14 37852 194 37877
rect 14 37818 15 37852
rect 49 37848 194 37852
rect 49 37818 87 37848
rect 14 37814 87 37818
rect 121 37843 194 37848
rect 121 37814 159 37843
rect 14 37809 159 37814
rect 193 37809 194 37843
rect 14 37784 194 37809
rect 14 37750 15 37784
rect 49 37780 194 37784
rect 49 37750 87 37780
rect 14 37746 87 37750
rect 121 37775 194 37780
rect 121 37746 159 37775
rect 14 37741 159 37746
rect 193 37741 194 37775
rect 14 37716 194 37741
rect 14 37682 15 37716
rect 49 37712 194 37716
rect 49 37682 87 37712
rect 14 37678 87 37682
rect 121 37707 194 37712
rect 121 37678 159 37707
rect 14 37673 159 37678
rect 193 37673 194 37707
rect 14 37648 194 37673
rect 14 37614 15 37648
rect 49 37644 194 37648
rect 49 37614 87 37644
rect 14 37610 87 37614
rect 121 37639 194 37644
rect 121 37610 159 37639
rect 14 37605 159 37610
rect 193 37605 194 37639
rect 14 37580 194 37605
rect 14 37546 15 37580
rect 49 37576 194 37580
rect 49 37546 87 37576
rect 14 37542 87 37546
rect 121 37571 194 37576
rect 121 37542 159 37571
rect 14 37537 159 37542
rect 193 37537 194 37571
rect 14 37512 194 37537
rect 14 37478 15 37512
rect 49 37508 194 37512
rect 49 37478 87 37508
rect 14 37474 87 37478
rect 121 37503 194 37508
rect 121 37474 159 37503
rect 14 37469 159 37474
rect 193 37469 194 37503
rect 14 37444 194 37469
rect 14 37410 15 37444
rect 49 37440 194 37444
rect 49 37410 87 37440
rect 14 37406 87 37410
rect 121 37435 194 37440
rect 121 37406 159 37435
rect 14 37401 159 37406
rect 193 37401 194 37435
rect 14 37376 194 37401
rect 14 37342 15 37376
rect 49 37372 194 37376
rect 49 37342 87 37372
rect 14 37338 87 37342
rect 121 37367 194 37372
rect 121 37338 159 37367
rect 14 37333 159 37338
rect 193 37333 194 37367
rect 14 37308 194 37333
rect 14 37274 15 37308
rect 49 37304 194 37308
rect 49 37274 87 37304
rect 14 37270 87 37274
rect 121 37299 194 37304
rect 121 37270 159 37299
rect 14 37265 159 37270
rect 193 37265 194 37299
rect 14 37240 194 37265
rect 14 37206 15 37240
rect 49 37236 194 37240
rect 49 37206 87 37236
rect 14 37202 87 37206
rect 121 37231 194 37236
rect 121 37202 159 37231
rect 14 37197 159 37202
rect 193 37197 194 37231
rect 14 37172 194 37197
rect 14 37138 15 37172
rect 49 37168 194 37172
rect 49 37138 87 37168
rect 14 37134 87 37138
rect 121 37163 194 37168
rect 121 37134 159 37163
rect 14 37129 159 37134
rect 193 37129 194 37163
rect 14 37104 194 37129
rect 14 37070 15 37104
rect 49 37100 194 37104
rect 49 37070 87 37100
rect 14 37066 87 37070
rect 121 37095 194 37100
rect 121 37066 159 37095
rect 14 37061 159 37066
rect 193 37061 194 37095
rect 14 37036 194 37061
rect 14 37002 15 37036
rect 49 37032 194 37036
rect 49 37002 87 37032
rect 14 36998 87 37002
rect 121 37027 194 37032
rect 121 36998 159 37027
rect 14 36993 159 36998
rect 193 36993 194 37027
rect 14 36968 194 36993
rect 14 36934 15 36968
rect 49 36964 194 36968
rect 49 36934 87 36964
rect 14 36930 87 36934
rect 121 36959 194 36964
rect 121 36930 159 36959
rect 14 36925 159 36930
rect 193 36925 194 36959
rect 14 36900 194 36925
rect 14 36866 15 36900
rect 49 36896 194 36900
rect 49 36866 87 36896
rect 14 36862 87 36866
rect 121 36891 194 36896
rect 121 36862 159 36891
rect 14 36857 159 36862
rect 193 36857 194 36891
rect 14 36832 194 36857
rect 14 36798 15 36832
rect 49 36828 194 36832
rect 49 36798 87 36828
rect 14 36794 87 36798
rect 121 36823 194 36828
rect 121 36794 159 36823
rect 14 36789 159 36794
rect 193 36789 194 36823
rect 14 36764 194 36789
rect 14 36730 15 36764
rect 49 36760 194 36764
rect 49 36730 87 36760
rect 14 36726 87 36730
rect 121 36755 194 36760
rect 121 36726 159 36755
rect 14 36721 159 36726
rect 193 36721 194 36755
rect 14 36696 194 36721
rect 14 36662 15 36696
rect 49 36692 194 36696
rect 49 36662 87 36692
rect 14 36658 87 36662
rect 121 36687 194 36692
rect 121 36658 159 36687
rect 14 36653 159 36658
rect 193 36653 194 36687
rect 14 36628 194 36653
rect 14 36594 15 36628
rect 49 36624 194 36628
rect 49 36594 87 36624
rect 14 36590 87 36594
rect 121 36619 194 36624
rect 121 36590 159 36619
rect 14 36585 159 36590
rect 193 36585 194 36619
rect 14 36560 194 36585
rect 14 36526 15 36560
rect 49 36556 194 36560
rect 49 36526 87 36556
rect 14 36522 87 36526
rect 121 36551 194 36556
rect 121 36522 159 36551
rect 14 36517 159 36522
rect 193 36517 194 36551
rect 14 36492 194 36517
rect 14 36458 15 36492
rect 49 36488 194 36492
rect 49 36458 87 36488
rect 14 36454 87 36458
rect 121 36483 194 36488
rect 121 36454 159 36483
rect 14 36449 159 36454
rect 193 36449 194 36483
rect 14 36424 194 36449
rect 14 36390 15 36424
rect 49 36420 194 36424
rect 49 36390 87 36420
rect 14 36386 87 36390
rect 121 36415 194 36420
rect 121 36386 159 36415
rect 14 36381 159 36386
rect 193 36381 194 36415
rect 14 36356 194 36381
rect 14 36322 15 36356
rect 49 36352 194 36356
rect 49 36322 87 36352
rect 14 36318 87 36322
rect 121 36347 194 36352
rect 121 36318 159 36347
rect 14 36313 159 36318
rect 193 36313 194 36347
rect 14 36288 194 36313
rect 14 36254 15 36288
rect 49 36284 194 36288
rect 49 36254 87 36284
rect 14 36250 87 36254
rect 121 36279 194 36284
rect 121 36250 159 36279
rect 14 36245 159 36250
rect 193 36245 194 36279
rect 14 36220 194 36245
rect 14 36186 15 36220
rect 49 36216 194 36220
rect 49 36186 87 36216
rect 14 36182 87 36186
rect 121 36211 194 36216
rect 121 36182 159 36211
rect 14 36177 159 36182
rect 193 36177 194 36211
rect 14 36152 194 36177
rect 14 36118 15 36152
rect 49 36148 194 36152
rect 49 36118 87 36148
rect 14 36114 87 36118
rect 121 36143 194 36148
rect 121 36114 159 36143
rect 14 36109 159 36114
rect 193 36109 194 36143
rect 14 36084 194 36109
rect 14 36050 15 36084
rect 49 36080 194 36084
rect 49 36050 87 36080
rect 14 36046 87 36050
rect 121 36075 194 36080
rect 121 36046 159 36075
rect 14 36041 159 36046
rect 193 36041 194 36075
rect 14 36016 194 36041
rect 14 35982 15 36016
rect 49 36012 194 36016
rect 49 35982 87 36012
rect 14 35978 87 35982
rect 121 36007 194 36012
rect 121 35978 159 36007
rect 14 35973 159 35978
rect 193 35973 194 36007
rect 14 35948 194 35973
rect 14 35914 15 35948
rect 49 35944 194 35948
rect 49 35914 87 35944
rect 14 35910 87 35914
rect 121 35939 194 35944
rect 121 35910 159 35939
rect 14 35905 159 35910
rect 193 35905 194 35939
rect 14 35880 194 35905
rect 14 35846 15 35880
rect 49 35876 194 35880
rect 49 35846 87 35876
rect 14 35842 87 35846
rect 121 35871 194 35876
rect 121 35842 159 35871
rect 14 35837 159 35842
rect 193 35837 194 35871
rect 14 35812 194 35837
rect 14 35778 15 35812
rect 49 35808 194 35812
rect 49 35778 87 35808
rect 14 35774 87 35778
rect 121 35803 194 35808
rect 121 35774 159 35803
rect 14 35769 159 35774
rect 193 35769 194 35803
rect 14 35744 194 35769
rect 14 35710 15 35744
rect 49 35740 194 35744
rect 49 35710 87 35740
rect 14 35706 87 35710
rect 121 35735 194 35740
rect 121 35706 159 35735
rect 14 35701 159 35706
rect 193 35701 194 35735
rect 14 35676 194 35701
rect 14 35642 15 35676
rect 49 35672 194 35676
rect 49 35642 87 35672
rect 14 35638 87 35642
rect 121 35667 194 35672
rect 121 35638 159 35667
rect 14 35633 159 35638
rect 193 35633 194 35667
rect 14 35608 194 35633
rect 14 35574 15 35608
rect 49 35604 194 35608
rect 49 35574 87 35604
rect 14 35570 87 35574
rect 121 35599 194 35604
rect 121 35570 159 35599
rect 14 35565 159 35570
rect 193 35565 194 35599
rect 14 35540 194 35565
rect 14 35506 15 35540
rect 49 35536 194 35540
rect 49 35506 87 35536
rect 14 35502 87 35506
rect 121 35531 194 35536
rect 121 35502 159 35531
rect 14 35497 159 35502
rect 193 35497 194 35531
rect 14 35472 194 35497
rect 14 35438 15 35472
rect 49 35468 194 35472
rect 49 35438 87 35468
rect 14 35434 87 35438
rect 121 35463 194 35468
rect 121 35434 159 35463
rect 14 35429 159 35434
rect 193 35429 194 35463
rect 14 35404 194 35429
rect 14 35370 15 35404
rect 49 35400 194 35404
rect 49 35370 87 35400
rect 14 35366 87 35370
rect 121 35395 194 35400
rect 121 35366 159 35395
rect 14 35361 159 35366
rect 193 35361 194 35395
rect 14 35336 194 35361
rect 14 35302 15 35336
rect 49 35332 194 35336
rect 49 35302 87 35332
rect 14 35298 87 35302
rect 121 35327 194 35332
rect 121 35298 159 35327
rect 14 35293 159 35298
rect 193 35293 194 35327
rect 14 35268 194 35293
rect 14 35234 15 35268
rect 49 35264 194 35268
rect 49 35234 87 35264
rect 14 35230 87 35234
rect 121 35259 194 35264
rect 121 35230 159 35259
rect 14 35225 159 35230
rect 193 35225 194 35259
rect 14 35200 194 35225
rect 14 35166 15 35200
rect 49 35196 194 35200
rect 49 35166 87 35196
rect 14 35162 87 35166
rect 121 35191 194 35196
rect 121 35162 159 35191
rect 14 35157 159 35162
rect 193 35157 194 35191
rect 14 35132 194 35157
rect 14 35098 15 35132
rect 49 35128 194 35132
rect 49 35098 87 35128
rect 14 35094 87 35098
rect 121 35123 194 35128
rect 121 35094 159 35123
rect 14 35089 159 35094
rect 193 35089 194 35123
rect 14 35064 194 35089
rect 14 35030 15 35064
rect 49 35060 194 35064
rect 49 35030 87 35060
rect 14 35026 87 35030
rect 121 35055 194 35060
rect 121 35026 159 35055
rect 14 35021 159 35026
rect 193 35021 194 35055
rect 14 34996 194 35021
rect 14 34962 15 34996
rect 49 34992 194 34996
rect 49 34962 87 34992
rect 14 34958 87 34962
rect 121 34987 194 34992
rect 121 34958 159 34987
rect 14 34953 159 34958
rect 193 34953 194 34987
rect 14 34928 194 34953
rect 14 34894 15 34928
rect 49 34924 194 34928
rect 49 34894 87 34924
rect 14 34890 87 34894
rect 121 34919 194 34924
rect 121 34890 159 34919
rect 14 34885 159 34890
rect 193 34885 194 34919
rect 14 34861 194 34885
rect -2867 34860 194 34861
rect -2867 34826 -2833 34860
rect -2799 34826 -2765 34860
rect -2731 34826 -2697 34860
rect -2663 34826 -2629 34860
rect -2595 34826 -2561 34860
rect -2527 34826 -2493 34860
rect -2459 34826 -2425 34860
rect -2391 34826 -2357 34860
rect -2323 34826 -2289 34860
rect -2255 34826 -2221 34860
rect -2187 34826 -2153 34860
rect -2119 34826 -2085 34860
rect -2051 34826 -2017 34860
rect -1983 34826 -1949 34860
rect -1915 34826 -1881 34860
rect -1847 34826 -1813 34860
rect -1779 34826 -1745 34860
rect -1711 34826 -1677 34860
rect -1643 34826 -1609 34860
rect -1575 34826 -1541 34860
rect -1507 34826 -1473 34860
rect -1439 34826 -1405 34860
rect -1371 34826 -1337 34860
rect -1303 34826 -1269 34860
rect -1235 34826 -1201 34860
rect -1167 34826 -1133 34860
rect -1099 34826 -1065 34860
rect -1031 34826 -997 34860
rect -963 34826 -929 34860
rect -895 34826 -861 34860
rect -827 34826 -793 34860
rect -759 34826 -725 34860
rect -691 34826 -657 34860
rect -623 34826 -589 34860
rect -555 34826 -521 34860
rect -487 34826 -453 34860
rect -419 34826 -385 34860
rect -351 34826 -317 34860
rect -283 34826 -249 34860
rect -215 34826 -181 34860
rect -147 34826 -113 34860
rect -79 34826 15 34860
rect 49 34856 194 34860
rect 49 34826 87 34856
rect -2867 34822 87 34826
rect 121 34851 194 34856
rect 121 34822 159 34851
rect -2867 34817 159 34822
rect 193 34817 194 34851
rect -2867 34788 194 34817
rect -2867 34754 -2833 34788
rect -2799 34754 -2765 34788
rect -2731 34754 -2697 34788
rect -2663 34754 -2629 34788
rect -2595 34754 -2561 34788
rect -2527 34754 -2493 34788
rect -2459 34754 -2425 34788
rect -2391 34754 -2357 34788
rect -2323 34754 -2289 34788
rect -2255 34754 -2221 34788
rect -2187 34754 -2153 34788
rect -2119 34754 -2085 34788
rect -2051 34754 -2017 34788
rect -1983 34754 -1949 34788
rect -1915 34754 -1881 34788
rect -1847 34754 -1813 34788
rect -1779 34754 -1745 34788
rect -1711 34754 -1677 34788
rect -1643 34754 -1609 34788
rect -1575 34754 -1541 34788
rect -1507 34754 -1473 34788
rect -1439 34754 -1405 34788
rect -1371 34754 -1337 34788
rect -1303 34754 -1269 34788
rect -1235 34754 -1201 34788
rect -1167 34754 -1133 34788
rect -1099 34754 -1065 34788
rect -1031 34754 -997 34788
rect -963 34754 -929 34788
rect -895 34754 -861 34788
rect -827 34754 -793 34788
rect -759 34754 -725 34788
rect -691 34754 -657 34788
rect -623 34754 -589 34788
rect -555 34754 -521 34788
rect -487 34754 -453 34788
rect -419 34754 -385 34788
rect -351 34754 -317 34788
rect -283 34754 -249 34788
rect -215 34754 -181 34788
rect -147 34754 -113 34788
rect -79 34754 -45 34788
rect -11 34754 87 34788
rect 121 34783 194 34788
rect 121 34754 159 34783
rect -2867 34749 159 34754
rect 193 34749 194 34783
rect -2867 34716 194 34749
rect -2867 34682 -2833 34716
rect -2799 34682 -2765 34716
rect -2731 34682 -2697 34716
rect -2663 34682 -2629 34716
rect -2595 34682 -2561 34716
rect -2527 34682 -2493 34716
rect -2459 34682 -2425 34716
rect -2391 34682 -2357 34716
rect -2323 34682 -2289 34716
rect -2255 34682 -2221 34716
rect -2187 34682 -2153 34716
rect -2119 34682 -2085 34716
rect -2051 34682 -2017 34716
rect -1983 34682 -1949 34716
rect -1915 34682 -1881 34716
rect -1847 34682 -1813 34716
rect -1779 34682 -1745 34716
rect -1711 34682 -1677 34716
rect -1643 34682 -1609 34716
rect -1575 34682 -1541 34716
rect -1507 34682 -1473 34716
rect -1439 34682 -1405 34716
rect -1371 34682 -1337 34716
rect -1303 34682 -1269 34716
rect -1235 34682 -1201 34716
rect -1167 34682 -1133 34716
rect -1099 34682 -1065 34716
rect -1031 34682 -997 34716
rect -963 34682 -929 34716
rect -895 34682 -861 34716
rect -827 34682 -793 34716
rect -759 34682 -725 34716
rect -691 34682 -657 34716
rect -623 34682 -589 34716
rect -555 34682 -521 34716
rect -487 34682 -453 34716
rect -419 34682 -385 34716
rect -351 34682 -317 34716
rect -283 34682 -249 34716
rect -215 34682 -181 34716
rect -147 34682 -113 34716
rect -79 34682 -45 34716
rect -11 34682 23 34716
rect 57 34682 91 34716
rect 125 34682 194 34716
rect -2867 34647 194 34682
rect -2856 19197 337 20380
rect -2969 18004 -17 19031
rect -2969 17940 2600 18004
rect -2969 17927 -17 17940
rect -2969 17925 -2959 17927
rect -2966 10413 -2959 17925
rect -273 17726 -17 17927
rect -273 10413 -266 17726
rect 10639 15870 10772 16576
rect 11631 15870 11774 16570
rect 10639 15836 10732 15870
rect 10766 15836 10772 15870
rect 10639 15773 10772 15836
rect 10639 15739 10732 15773
rect 10766 15739 10772 15773
rect 10639 15155 10772 15739
rect 10989 15751 11023 15836
rect 11341 15751 11375 15836
rect 11631 15836 11637 15870
rect 11671 15836 11774 15870
rect 11631 15751 11774 15836
rect 11631 15717 11637 15751
rect 11671 15717 11774 15751
rect 11631 15177 11774 15717
rect 10639 15121 10732 15155
rect 10766 15121 10772 15155
rect 10639 15102 10772 15121
rect 10659 15058 10772 15102
rect 10659 15024 10732 15058
rect 10766 15024 10772 15058
rect 10989 15058 11023 15143
rect 11341 15058 11375 15143
rect 11631 15143 11637 15177
rect 11671 15143 11723 15177
rect 11757 15143 11774 15177
rect 11631 15058 11774 15143
rect 11631 15024 11637 15058
rect 11671 15024 11723 15058
rect 11757 15024 11774 15058
rect 642 14245 819 14723
rect 5537 14461 5669 14727
rect 7137 14473 7269 14722
rect 10659 14510 10772 15024
rect 11631 14509 11774 15024
rect 5537 14248 5721 14461
rect 5537 14245 5735 14248
rect 642 14233 783 14245
rect 85 14199 124 14233
rect 158 14199 197 14233
rect 231 14199 270 14233
rect 304 14199 343 14233
rect 377 14199 416 14233
rect 450 14199 489 14233
rect 523 14199 563 14233
rect 597 14199 637 14233
rect 671 14199 711 14233
rect 745 14211 783 14233
rect 817 14211 822 14245
rect 745 14199 822 14211
rect 51 14168 822 14199
rect 51 14161 783 14168
rect 85 14127 124 14161
rect 158 14127 197 14161
rect 231 14127 270 14161
rect 304 14127 343 14161
rect 377 14127 416 14161
rect 450 14127 489 14161
rect 523 14127 563 14161
rect 597 14127 637 14161
rect 671 14127 711 14161
rect 745 14134 783 14161
rect 817 14134 822 14168
rect 1026 14211 1031 14245
rect 1065 14211 1070 14245
rect 1026 14171 1070 14211
rect 1026 14137 1031 14171
rect 1065 14137 1070 14171
rect 5537 14211 5588 14245
rect 5622 14211 5701 14245
rect 5537 14208 5735 14211
rect 745 14127 822 14134
rect 51 14091 822 14127
rect 51 14089 783 14091
rect 85 14055 124 14089
rect 158 14055 197 14089
rect 231 14055 270 14089
rect 304 14055 343 14089
rect 377 14055 416 14089
rect 450 14055 489 14089
rect 523 14055 563 14089
rect 597 14055 637 14089
rect 671 14055 711 14089
rect 745 14057 783 14089
rect 817 14057 822 14091
rect 745 14055 819 14057
rect 642 13723 819 14055
rect 5537 13727 5669 14208
rect 6259 14205 6293 14259
rect 6571 14205 6605 14259
rect 6883 14205 6917 14259
rect 7107 14206 7269 14473
rect 18281 14481 29669 14484
rect 18281 14447 18349 14481
rect 18383 14447 18418 14481
rect 18452 14447 18487 14481
rect 18521 14447 18556 14481
rect 18590 14447 18625 14481
rect 18659 14447 18694 14481
rect 18728 14447 18763 14481
rect 18797 14447 18832 14481
rect 18866 14447 18901 14481
rect 18935 14447 18970 14481
rect 19004 14447 19039 14481
rect 19073 14447 19108 14481
rect 19142 14447 19177 14481
rect 19211 14447 19246 14481
rect 19280 14447 19315 14481
rect 19349 14447 19384 14481
rect 19418 14447 19453 14481
rect 19487 14447 19522 14481
rect 19556 14447 19591 14481
rect 19625 14447 19660 14481
rect 19694 14447 19729 14481
rect 19763 14447 19798 14481
rect 19832 14447 19867 14481
rect 19901 14447 19936 14481
rect 19970 14447 20005 14481
rect 20039 14447 20074 14481
rect 20108 14447 20143 14481
rect 20177 14447 20212 14481
rect 20246 14447 20281 14481
rect 20315 14447 20350 14481
rect 20384 14447 20419 14481
rect 20453 14447 20488 14481
rect 20522 14447 20557 14481
rect 20591 14447 20626 14481
rect 20660 14447 20695 14481
rect 20729 14447 20764 14481
rect 20798 14447 20833 14481
rect 20867 14447 20902 14481
rect 20936 14447 20971 14481
rect 21005 14447 21040 14481
rect 21074 14447 21109 14481
rect 21143 14447 21178 14481
rect 21212 14447 21247 14481
rect 21281 14447 21315 14481
rect 21349 14447 21383 14481
rect 21417 14447 21451 14481
rect 21485 14447 21519 14481
rect 21553 14447 21587 14481
rect 21621 14447 21655 14481
rect 21689 14447 21723 14481
rect 21757 14447 21791 14481
rect 21825 14447 21859 14481
rect 21893 14447 21927 14481
rect 21961 14447 21995 14481
rect 22029 14447 22063 14481
rect 22097 14447 22131 14481
rect 22165 14447 22199 14481
rect 22233 14447 22267 14481
rect 22301 14447 22335 14481
rect 22369 14447 22403 14481
rect 22437 14447 22471 14481
rect 22505 14447 22539 14481
rect 22573 14447 22607 14481
rect 22641 14447 22675 14481
rect 22709 14447 22743 14481
rect 22777 14447 22811 14481
rect 22845 14447 22879 14481
rect 22913 14447 22947 14481
rect 22981 14447 23015 14481
rect 23049 14447 23083 14481
rect 23117 14447 23151 14481
rect 23185 14447 23219 14481
rect 23253 14447 23287 14481
rect 23321 14447 23355 14481
rect 23389 14447 23423 14481
rect 23457 14447 23491 14481
rect 23525 14447 23559 14481
rect 23593 14447 23627 14481
rect 23661 14447 23695 14481
rect 23729 14447 23763 14481
rect 23797 14447 23831 14481
rect 23865 14447 23899 14481
rect 23933 14447 23967 14481
rect 24001 14447 24035 14481
rect 24069 14447 24103 14481
rect 24137 14447 24171 14481
rect 24205 14447 24239 14481
rect 24273 14447 24307 14481
rect 24341 14447 24375 14481
rect 24409 14447 24443 14481
rect 24477 14447 24511 14481
rect 24545 14447 24579 14481
rect 24613 14447 24647 14481
rect 24681 14447 24715 14481
rect 24749 14447 24783 14481
rect 24817 14447 24851 14481
rect 24885 14447 24919 14481
rect 24953 14447 24987 14481
rect 25021 14447 25055 14481
rect 25089 14447 25123 14481
rect 25157 14447 25191 14481
rect 25225 14447 25259 14481
rect 25293 14447 25327 14481
rect 25361 14447 25395 14481
rect 25429 14447 25463 14481
rect 25497 14447 25531 14481
rect 25565 14447 25599 14481
rect 25633 14447 25667 14481
rect 25701 14447 25735 14481
rect 25769 14447 25803 14481
rect 25837 14447 25871 14481
rect 25905 14447 25939 14481
rect 25973 14447 26007 14481
rect 26041 14447 26075 14481
rect 26109 14447 26143 14481
rect 26177 14447 26211 14481
rect 26245 14447 26279 14481
rect 26313 14447 26347 14481
rect 26381 14447 26415 14481
rect 26449 14447 26483 14481
rect 26517 14447 26551 14481
rect 26585 14447 26619 14481
rect 26653 14447 26687 14481
rect 26721 14447 26755 14481
rect 26789 14447 26823 14481
rect 26857 14447 26891 14481
rect 26925 14447 26959 14481
rect 26993 14447 27027 14481
rect 27061 14447 27095 14481
rect 27129 14447 27163 14481
rect 27197 14447 27231 14481
rect 27265 14447 27299 14481
rect 27333 14447 27367 14481
rect 27401 14447 27435 14481
rect 27469 14447 27503 14481
rect 27537 14447 27571 14481
rect 27605 14447 27639 14481
rect 27673 14447 27707 14481
rect 27741 14447 27775 14481
rect 27809 14447 27843 14481
rect 27877 14447 27911 14481
rect 27945 14447 27979 14481
rect 28013 14447 28047 14481
rect 28081 14447 28115 14481
rect 28149 14447 28183 14481
rect 28217 14447 28251 14481
rect 28285 14447 28319 14481
rect 28353 14447 28387 14481
rect 28421 14447 28455 14481
rect 28489 14447 28523 14481
rect 28557 14447 28591 14481
rect 28625 14447 28659 14481
rect 28693 14447 28727 14481
rect 28761 14447 28795 14481
rect 28829 14447 28863 14481
rect 28897 14447 28931 14481
rect 28965 14447 28999 14481
rect 29033 14447 29067 14481
rect 29101 14447 29135 14481
rect 29169 14447 29203 14481
rect 29237 14447 29271 14481
rect 29305 14447 29339 14481
rect 29373 14447 29407 14481
rect 29441 14447 29475 14481
rect 29509 14447 29543 14481
rect 29577 14447 29611 14481
rect 29645 14447 29669 14481
rect 18281 14415 29669 14447
rect 18281 14381 18284 14415
rect 18318 14409 29669 14415
rect 18318 14381 18356 14409
rect 18390 14398 18425 14409
rect 18459 14398 18494 14409
rect 18528 14398 18563 14409
rect 18597 14398 18632 14409
rect 18666 14398 18701 14409
rect 18735 14398 18770 14409
rect 18804 14398 18839 14409
rect 18873 14398 18908 14409
rect 18281 14375 18356 14381
rect 18393 14375 18425 14398
rect 18466 14375 18494 14398
rect 18539 14375 18563 14398
rect 18612 14375 18632 14398
rect 18685 14375 18701 14398
rect 18758 14375 18770 14398
rect 18831 14375 18839 14398
rect 18904 14375 18908 14398
rect 18942 14398 18977 14409
rect 18942 14375 18943 14398
rect 18281 14364 18359 14375
rect 18393 14364 18432 14375
rect 18466 14364 18505 14375
rect 18539 14364 18578 14375
rect 18612 14364 18651 14375
rect 18685 14364 18724 14375
rect 18758 14364 18797 14375
rect 18831 14364 18870 14375
rect 18904 14364 18943 14375
rect 19011 14398 19046 14409
rect 19080 14398 19115 14409
rect 19149 14398 19184 14409
rect 19218 14398 19253 14409
rect 19287 14398 19322 14409
rect 19356 14398 19391 14409
rect 19425 14398 19460 14409
rect 19494 14398 19529 14409
rect 19011 14375 19016 14398
rect 19080 14375 19089 14398
rect 19149 14375 19162 14398
rect 19218 14375 19235 14398
rect 19287 14375 19308 14398
rect 19356 14375 19381 14398
rect 19425 14375 19454 14398
rect 19494 14375 19527 14398
rect 19563 14375 19598 14409
rect 19632 14398 19667 14409
rect 19701 14398 19736 14409
rect 19770 14398 19805 14409
rect 19839 14398 19874 14409
rect 19908 14398 19943 14409
rect 19977 14398 20012 14409
rect 20046 14398 20081 14409
rect 20115 14398 20150 14409
rect 19634 14375 19667 14398
rect 19707 14375 19736 14398
rect 19780 14375 19805 14398
rect 19853 14375 19874 14398
rect 19926 14375 19943 14398
rect 19999 14375 20012 14398
rect 20072 14375 20081 14398
rect 20145 14375 20150 14398
rect 20184 14398 20219 14409
rect 18977 14364 19016 14375
rect 19050 14364 19089 14375
rect 19123 14364 19162 14375
rect 19196 14364 19235 14375
rect 19269 14364 19308 14375
rect 19342 14364 19381 14375
rect 19415 14364 19454 14375
rect 19488 14364 19527 14375
rect 19561 14364 19600 14375
rect 19634 14364 19673 14375
rect 19707 14364 19746 14375
rect 19780 14364 19819 14375
rect 19853 14364 19892 14375
rect 19926 14364 19965 14375
rect 19999 14364 20038 14375
rect 20072 14364 20111 14375
rect 20145 14364 20184 14375
rect 20218 14375 20219 14398
rect 20253 14398 20288 14409
rect 20322 14398 20357 14409
rect 20391 14398 20426 14409
rect 20460 14398 20495 14409
rect 20529 14398 20564 14409
rect 20598 14398 20633 14409
rect 20667 14398 20702 14409
rect 20736 14398 20771 14409
rect 20253 14375 20257 14398
rect 20322 14375 20330 14398
rect 20391 14375 20403 14398
rect 20460 14375 20476 14398
rect 20529 14375 20549 14398
rect 20598 14375 20622 14398
rect 20667 14375 20695 14398
rect 20736 14375 20768 14398
rect 20805 14375 20839 14409
rect 20873 14398 20907 14409
rect 20941 14398 20975 14409
rect 21009 14398 21043 14409
rect 21077 14398 21111 14409
rect 21145 14398 21179 14409
rect 21213 14398 21247 14409
rect 21281 14398 21315 14409
rect 20875 14375 20907 14398
rect 20948 14375 20975 14398
rect 21021 14375 21043 14398
rect 21094 14375 21111 14398
rect 21167 14375 21179 14398
rect 21240 14375 21247 14398
rect 21313 14375 21315 14398
rect 21349 14398 21383 14409
rect 21417 14398 21451 14409
rect 21485 14398 21519 14409
rect 21553 14398 21587 14409
rect 21621 14398 21655 14409
rect 21689 14398 21723 14409
rect 21757 14398 21791 14409
rect 21349 14375 21352 14398
rect 21417 14375 21425 14398
rect 21485 14375 21498 14398
rect 21553 14375 21571 14398
rect 21621 14375 21644 14398
rect 21689 14375 21717 14398
rect 21757 14375 21790 14398
rect 21825 14375 21859 14409
rect 21893 14398 21927 14409
rect 21961 14398 21995 14409
rect 22029 14398 22063 14409
rect 22097 14398 22131 14409
rect 22165 14398 22199 14409
rect 22233 14398 22267 14409
rect 21897 14375 21927 14398
rect 21970 14375 21995 14398
rect 22043 14375 22063 14398
rect 22116 14375 22131 14398
rect 22189 14375 22199 14398
rect 22262 14375 22267 14398
rect 22301 14398 22335 14409
rect 20218 14364 20257 14375
rect 20291 14364 20330 14375
rect 20364 14364 20403 14375
rect 20437 14364 20476 14375
rect 20510 14364 20549 14375
rect 20583 14364 20622 14375
rect 20656 14364 20695 14375
rect 20729 14364 20768 14375
rect 20802 14364 20841 14375
rect 20875 14364 20914 14375
rect 20948 14364 20987 14375
rect 21021 14364 21060 14375
rect 21094 14364 21133 14375
rect 21167 14364 21206 14375
rect 21240 14364 21279 14375
rect 21313 14364 21352 14375
rect 21386 14364 21425 14375
rect 21459 14364 21498 14375
rect 21532 14364 21571 14375
rect 21605 14364 21644 14375
rect 21678 14364 21717 14375
rect 21751 14364 21790 14375
rect 21824 14364 21863 14375
rect 21897 14364 21936 14375
rect 21970 14364 22009 14375
rect 22043 14364 22082 14375
rect 22116 14364 22155 14375
rect 22189 14364 22228 14375
rect 22262 14364 22301 14375
rect 22369 14398 22403 14409
rect 22437 14398 22471 14409
rect 22505 14398 22539 14409
rect 22573 14398 22607 14409
rect 22641 14398 22675 14409
rect 22709 14398 22743 14409
rect 22777 14398 22811 14409
rect 22845 14398 22879 14409
rect 22369 14375 22373 14398
rect 22437 14375 22445 14398
rect 22505 14375 22517 14398
rect 22573 14375 22589 14398
rect 22641 14375 22661 14398
rect 22709 14375 22733 14398
rect 22777 14375 22805 14398
rect 22845 14375 22877 14398
rect 22913 14375 22947 14409
rect 22981 14398 23015 14409
rect 23049 14398 23083 14409
rect 23117 14398 23151 14409
rect 22983 14375 23015 14398
rect 23055 14375 23083 14398
rect 23127 14375 23151 14398
rect 23185 14375 23219 14409
rect 23253 14375 23287 14409
rect 23321 14375 23355 14409
rect 23389 14375 23423 14409
rect 23457 14398 23491 14409
rect 23525 14398 23559 14409
rect 23593 14398 23627 14409
rect 23661 14398 23695 14409
rect 23729 14398 23763 14409
rect 23797 14398 23831 14409
rect 23462 14375 23491 14398
rect 23535 14375 23559 14398
rect 23608 14375 23627 14398
rect 23681 14375 23695 14398
rect 23754 14375 23763 14398
rect 23827 14375 23831 14398
rect 23865 14398 23899 14409
rect 22335 14364 22373 14375
rect 22407 14364 22445 14375
rect 22479 14364 22517 14375
rect 22551 14364 22589 14375
rect 22623 14364 22661 14375
rect 22695 14364 22733 14375
rect 22767 14364 22805 14375
rect 22839 14364 22877 14375
rect 22911 14364 22949 14375
rect 22983 14364 23021 14375
rect 23055 14364 23093 14375
rect 23127 14364 23355 14375
rect 23389 14364 23428 14375
rect 23462 14364 23501 14375
rect 23535 14364 23574 14375
rect 23608 14364 23647 14375
rect 23681 14364 23720 14375
rect 23754 14364 23793 14375
rect 23827 14364 23865 14375
rect 23933 14398 23967 14409
rect 24001 14398 24035 14409
rect 24069 14398 24103 14409
rect 24137 14398 24171 14409
rect 24205 14398 24239 14409
rect 24273 14398 24307 14409
rect 24341 14398 24375 14409
rect 24409 14398 24443 14409
rect 23933 14375 23937 14398
rect 24001 14375 24009 14398
rect 24069 14375 24081 14398
rect 24137 14375 24153 14398
rect 24205 14375 24225 14398
rect 24273 14375 24297 14398
rect 24341 14375 24369 14398
rect 24409 14375 24441 14398
rect 24477 14375 24511 14409
rect 24545 14398 24579 14409
rect 24613 14398 24647 14409
rect 24681 14398 24715 14409
rect 24749 14398 24783 14409
rect 24817 14398 24851 14409
rect 24885 14398 24919 14409
rect 24953 14398 24987 14409
rect 25021 14398 25055 14409
rect 24547 14375 24579 14398
rect 24619 14375 24647 14398
rect 24691 14375 24715 14398
rect 24763 14375 24783 14398
rect 24835 14375 24851 14398
rect 24907 14375 24919 14398
rect 24979 14375 24987 14398
rect 25051 14375 25055 14398
rect 25089 14398 25123 14409
rect 23899 14364 23937 14375
rect 23971 14364 24009 14375
rect 24043 14364 24081 14375
rect 24115 14364 24153 14375
rect 24187 14364 24225 14375
rect 24259 14364 24297 14375
rect 24331 14364 24369 14375
rect 24403 14364 24441 14375
rect 24475 14364 24513 14375
rect 24547 14364 24585 14375
rect 24619 14364 24657 14375
rect 24691 14364 24729 14375
rect 24763 14364 24801 14375
rect 24835 14364 24873 14375
rect 24907 14364 24945 14375
rect 24979 14364 25017 14375
rect 25051 14364 25089 14375
rect 25157 14398 25191 14409
rect 25225 14398 25259 14409
rect 25293 14398 25327 14409
rect 25361 14398 25395 14409
rect 25429 14398 25463 14409
rect 25497 14398 25531 14409
rect 25565 14398 25599 14409
rect 25633 14398 25667 14409
rect 25157 14375 25161 14398
rect 25225 14375 25233 14398
rect 25293 14375 25305 14398
rect 25361 14375 25377 14398
rect 25429 14375 25449 14398
rect 25497 14375 25521 14398
rect 25565 14375 25593 14398
rect 25633 14375 25665 14398
rect 25701 14375 25735 14409
rect 25769 14398 25803 14409
rect 25837 14398 25871 14409
rect 25905 14398 25939 14409
rect 25973 14398 26007 14409
rect 26041 14398 26075 14409
rect 26109 14398 26143 14409
rect 26177 14398 26211 14409
rect 26245 14398 26279 14409
rect 25771 14375 25803 14398
rect 25843 14375 25871 14398
rect 25915 14375 25939 14398
rect 25987 14375 26007 14398
rect 26059 14375 26075 14398
rect 26131 14375 26143 14398
rect 26203 14375 26211 14398
rect 26275 14375 26279 14398
rect 26313 14398 26347 14409
rect 25123 14364 25161 14375
rect 25195 14364 25233 14375
rect 25267 14364 25305 14375
rect 25339 14364 25377 14375
rect 25411 14364 25449 14375
rect 25483 14364 25521 14375
rect 25555 14364 25593 14375
rect 25627 14364 25665 14375
rect 25699 14364 25737 14375
rect 25771 14364 25809 14375
rect 25843 14364 25881 14375
rect 25915 14364 25953 14375
rect 25987 14364 26025 14375
rect 26059 14364 26097 14375
rect 26131 14364 26169 14375
rect 26203 14364 26241 14375
rect 26275 14364 26313 14375
rect 26381 14398 26415 14409
rect 26449 14398 26483 14409
rect 26517 14398 26551 14409
rect 26585 14398 26619 14409
rect 26653 14398 26687 14409
rect 26721 14398 26755 14409
rect 26789 14398 26823 14409
rect 26857 14398 26891 14409
rect 26381 14375 26385 14398
rect 26449 14375 26457 14398
rect 26517 14375 26529 14398
rect 26585 14375 26601 14398
rect 26653 14375 26673 14398
rect 26721 14375 26745 14398
rect 26789 14375 26817 14398
rect 26857 14375 26889 14398
rect 26925 14375 26959 14409
rect 26993 14398 27027 14409
rect 27061 14398 27095 14409
rect 27129 14398 27163 14409
rect 27197 14398 27231 14409
rect 27265 14398 27299 14409
rect 27333 14398 27367 14409
rect 27401 14398 27435 14409
rect 27469 14398 27503 14409
rect 26995 14375 27027 14398
rect 27067 14375 27095 14398
rect 27139 14375 27163 14398
rect 27211 14375 27231 14398
rect 27283 14375 27299 14398
rect 27355 14375 27367 14398
rect 27427 14375 27435 14398
rect 27499 14375 27503 14398
rect 27537 14398 27571 14409
rect 26347 14364 26385 14375
rect 26419 14364 26457 14375
rect 26491 14364 26529 14375
rect 26563 14364 26601 14375
rect 26635 14364 26673 14375
rect 26707 14364 26745 14375
rect 26779 14364 26817 14375
rect 26851 14364 26889 14375
rect 26923 14364 26961 14375
rect 26995 14364 27033 14375
rect 27067 14364 27105 14375
rect 27139 14364 27177 14375
rect 27211 14364 27249 14375
rect 27283 14364 27321 14375
rect 27355 14364 27393 14375
rect 27427 14364 27465 14375
rect 27499 14364 27537 14375
rect 27605 14398 27639 14409
rect 27673 14398 27707 14409
rect 27741 14398 27775 14409
rect 27809 14398 27843 14409
rect 27877 14398 27911 14409
rect 27945 14398 27979 14409
rect 28013 14398 28047 14409
rect 28081 14398 28115 14409
rect 27605 14375 27609 14398
rect 27673 14375 27681 14398
rect 27741 14375 27753 14398
rect 27809 14375 27825 14398
rect 27877 14375 27897 14398
rect 27945 14375 27969 14398
rect 28013 14375 28041 14398
rect 28081 14375 28113 14398
rect 28149 14375 28183 14409
rect 28217 14398 28251 14409
rect 28285 14398 28319 14409
rect 28353 14398 28387 14409
rect 28421 14398 28455 14409
rect 28489 14398 28523 14409
rect 28557 14398 28591 14409
rect 28625 14398 28659 14409
rect 28693 14398 28727 14409
rect 28219 14375 28251 14398
rect 28291 14375 28319 14398
rect 28363 14375 28387 14398
rect 28435 14375 28455 14398
rect 28507 14375 28523 14398
rect 28579 14375 28591 14398
rect 28651 14375 28659 14398
rect 28723 14375 28727 14398
rect 28761 14398 28795 14409
rect 27571 14364 27609 14375
rect 27643 14364 27681 14375
rect 27715 14364 27753 14375
rect 27787 14364 27825 14375
rect 27859 14364 27897 14375
rect 27931 14364 27969 14375
rect 28003 14364 28041 14375
rect 28075 14364 28113 14375
rect 28147 14364 28185 14375
rect 28219 14364 28257 14375
rect 28291 14364 28329 14375
rect 28363 14364 28401 14375
rect 28435 14364 28473 14375
rect 28507 14364 28545 14375
rect 28579 14364 28617 14375
rect 28651 14364 28689 14375
rect 28723 14364 28761 14375
rect 28829 14398 28863 14409
rect 28897 14398 28931 14409
rect 28965 14398 28999 14409
rect 29033 14398 29067 14409
rect 29101 14398 29135 14409
rect 29169 14398 29203 14409
rect 29237 14398 29271 14409
rect 29305 14398 29339 14409
rect 28829 14375 28833 14398
rect 28897 14375 28905 14398
rect 28965 14375 28977 14398
rect 29033 14375 29049 14398
rect 29101 14375 29121 14398
rect 29169 14375 29193 14398
rect 29237 14375 29265 14398
rect 29305 14375 29337 14398
rect 29373 14375 29407 14409
rect 29441 14398 29475 14409
rect 29509 14398 29543 14409
rect 29577 14398 29611 14409
rect 29645 14398 29669 14409
rect 29443 14375 29475 14398
rect 29515 14375 29543 14398
rect 29587 14375 29611 14398
rect 28795 14364 28833 14375
rect 28867 14364 28905 14375
rect 28939 14364 28977 14375
rect 29011 14364 29049 14375
rect 29083 14364 29121 14375
rect 29155 14364 29193 14375
rect 29227 14364 29265 14375
rect 29299 14364 29337 14375
rect 29371 14364 29409 14375
rect 29443 14364 29481 14375
rect 29515 14364 29553 14375
rect 29587 14364 29625 14375
rect 29659 14364 29669 14398
rect 18281 14345 29669 14364
rect 18281 14311 18284 14345
rect 18318 14340 29669 14345
rect 18318 14311 18356 14340
rect 18281 14306 18356 14311
rect 18390 14337 29669 14340
rect 18390 14306 18428 14337
rect 18281 14303 18428 14306
rect 18462 14303 18497 14337
rect 18531 14303 18566 14337
rect 18600 14303 18635 14337
rect 18669 14303 18704 14337
rect 18738 14303 18773 14337
rect 18807 14303 18842 14337
rect 18876 14303 18911 14337
rect 18945 14303 18980 14337
rect 19014 14303 19049 14337
rect 19083 14303 19118 14337
rect 19152 14303 19187 14337
rect 19221 14303 19256 14337
rect 19290 14303 19325 14337
rect 19359 14303 19394 14337
rect 19428 14303 19463 14337
rect 19497 14303 19532 14337
rect 19566 14303 19601 14337
rect 19635 14303 19670 14337
rect 19704 14303 19739 14337
rect 19773 14303 19808 14337
rect 19842 14303 19877 14337
rect 19911 14303 19946 14337
rect 19980 14303 20015 14337
rect 20049 14303 20084 14337
rect 20118 14303 20153 14337
rect 20187 14303 20222 14337
rect 20256 14303 20291 14337
rect 20325 14303 20360 14337
rect 20394 14303 20429 14337
rect 20463 14303 20498 14337
rect 20532 14303 20567 14337
rect 20601 14303 20635 14337
rect 20669 14303 20703 14337
rect 20737 14303 20771 14337
rect 20805 14303 20839 14337
rect 20873 14303 20907 14337
rect 20941 14303 20975 14337
rect 21009 14303 21043 14337
rect 21077 14303 21111 14337
rect 21145 14303 21179 14337
rect 21213 14303 21247 14337
rect 21281 14303 21315 14337
rect 21349 14303 21383 14337
rect 21417 14303 21451 14337
rect 21485 14303 21519 14337
rect 21553 14303 21587 14337
rect 21621 14303 21655 14337
rect 21689 14303 21723 14337
rect 21757 14303 21791 14337
rect 21825 14303 21859 14337
rect 21893 14303 21927 14337
rect 21961 14303 21995 14337
rect 22029 14303 22063 14337
rect 22097 14303 22131 14337
rect 22165 14303 22199 14337
rect 22233 14303 22267 14337
rect 22301 14303 22335 14337
rect 22369 14303 22403 14337
rect 22437 14303 22471 14337
rect 22505 14303 22539 14337
rect 22573 14303 22607 14337
rect 22641 14303 22675 14337
rect 22709 14303 22743 14337
rect 22777 14303 22811 14337
rect 22845 14303 22879 14337
rect 22913 14303 22947 14337
rect 22981 14303 23015 14337
rect 23049 14303 23083 14337
rect 23117 14303 23151 14337
rect 23185 14303 23219 14337
rect 23253 14303 23287 14337
rect 23321 14303 23355 14337
rect 23389 14303 23423 14337
rect 23457 14303 23491 14337
rect 23525 14303 23559 14337
rect 23593 14303 23627 14337
rect 23661 14303 23695 14337
rect 23729 14303 23763 14337
rect 23797 14303 23831 14337
rect 23865 14303 23899 14337
rect 23933 14303 23967 14337
rect 24001 14303 24035 14337
rect 24069 14303 24103 14337
rect 24137 14303 24171 14337
rect 24205 14303 24239 14337
rect 24273 14303 24307 14337
rect 24341 14303 24375 14337
rect 24409 14303 24443 14337
rect 24477 14303 24511 14337
rect 24545 14303 24579 14337
rect 24613 14303 24647 14337
rect 24681 14303 24715 14337
rect 24749 14303 24783 14337
rect 24817 14303 24851 14337
rect 24885 14303 24919 14337
rect 24953 14303 24987 14337
rect 25021 14303 25055 14337
rect 25089 14303 25123 14337
rect 25157 14303 25191 14337
rect 25225 14303 25259 14337
rect 25293 14303 25327 14337
rect 25361 14303 25395 14337
rect 25429 14303 25463 14337
rect 25497 14303 25531 14337
rect 25565 14303 25599 14337
rect 25633 14303 25667 14337
rect 25701 14303 25735 14337
rect 25769 14303 25803 14337
rect 25837 14303 25871 14337
rect 25905 14303 25939 14337
rect 25973 14303 26007 14337
rect 26041 14303 26075 14337
rect 26109 14303 26143 14337
rect 26177 14303 26211 14337
rect 26245 14303 26279 14337
rect 26313 14303 26347 14337
rect 26381 14303 26415 14337
rect 26449 14303 26483 14337
rect 26517 14303 26551 14337
rect 26585 14303 26619 14337
rect 26653 14303 26687 14337
rect 26721 14303 26755 14337
rect 26789 14303 26823 14337
rect 26857 14303 26891 14337
rect 26925 14303 26959 14337
rect 26993 14303 27027 14337
rect 27061 14303 27095 14337
rect 27129 14303 27163 14337
rect 27197 14303 27231 14337
rect 27265 14303 27299 14337
rect 27333 14303 27367 14337
rect 27401 14303 27435 14337
rect 27469 14303 27503 14337
rect 27537 14303 27571 14337
rect 27605 14303 27639 14337
rect 27673 14303 27707 14337
rect 27741 14303 27775 14337
rect 27809 14303 27843 14337
rect 27877 14303 27911 14337
rect 27945 14303 27979 14337
rect 28013 14303 28047 14337
rect 28081 14303 28115 14337
rect 28149 14303 28183 14337
rect 28217 14303 28251 14337
rect 28285 14303 28319 14337
rect 28353 14303 28387 14337
rect 28421 14303 28455 14337
rect 28489 14303 28523 14337
rect 28557 14303 28591 14337
rect 28625 14303 28659 14337
rect 28693 14303 28727 14337
rect 28761 14303 28795 14337
rect 28829 14303 28863 14337
rect 28897 14303 28931 14337
rect 28965 14303 28999 14337
rect 29033 14303 29067 14337
rect 29101 14303 29135 14337
rect 29169 14303 29203 14337
rect 29237 14303 29271 14337
rect 29305 14303 29339 14337
rect 29373 14303 29407 14337
rect 29441 14303 29475 14337
rect 29509 14303 29543 14337
rect 29577 14303 29611 14337
rect 29645 14303 29669 14337
rect 18281 14275 29669 14303
rect 18281 14241 18284 14275
rect 18318 14271 29669 14275
rect 18318 14241 18356 14271
rect 18281 14237 18356 14241
rect 18390 14268 29669 14271
rect 18390 14237 18428 14268
rect 18281 14234 18428 14237
rect 18462 14265 29669 14268
rect 18462 14234 18500 14265
rect 18281 14231 18500 14234
rect 18534 14231 18569 14265
rect 18603 14231 18638 14265
rect 18672 14231 18707 14265
rect 18741 14231 18776 14265
rect 18810 14231 18845 14265
rect 18879 14231 18914 14265
rect 18948 14231 18983 14265
rect 19017 14231 19052 14265
rect 19086 14231 19121 14265
rect 19155 14231 19190 14265
rect 19224 14231 19259 14265
rect 19293 14231 19328 14265
rect 19362 14231 19397 14265
rect 19431 14231 19466 14265
rect 19500 14231 19535 14265
rect 19569 14231 19604 14265
rect 19638 14231 19673 14265
rect 19707 14231 19742 14265
rect 19776 14231 19811 14265
rect 19845 14231 19880 14265
rect 19914 14231 19949 14265
rect 19983 14231 20018 14265
rect 20052 14231 20087 14265
rect 20121 14231 20156 14265
rect 20190 14231 20225 14265
rect 20259 14231 20294 14265
rect 20328 14231 20363 14265
rect 20397 14231 20431 14265
rect 20465 14231 20499 14265
rect 20533 14231 20567 14265
rect 20601 14231 20635 14265
rect 20669 14231 20703 14265
rect 20737 14231 20771 14265
rect 20805 14231 20839 14265
rect 20873 14231 20907 14265
rect 20941 14231 20975 14265
rect 21009 14231 21043 14265
rect 21077 14231 21111 14265
rect 21145 14231 21179 14265
rect 21213 14231 21247 14265
rect 21281 14231 21315 14265
rect 21349 14231 21383 14265
rect 21417 14231 21451 14265
rect 21485 14231 21519 14265
rect 21553 14231 21587 14265
rect 21621 14231 21655 14265
rect 21689 14231 21723 14265
rect 21757 14231 21791 14265
rect 21825 14231 21859 14265
rect 21893 14231 21927 14265
rect 21961 14231 21995 14265
rect 22029 14231 22063 14265
rect 22097 14231 22131 14265
rect 22165 14231 22199 14265
rect 22233 14231 22267 14265
rect 22301 14231 22335 14265
rect 22369 14231 22403 14265
rect 22437 14231 22471 14265
rect 22505 14231 22539 14265
rect 22573 14231 22607 14265
rect 22641 14231 22675 14265
rect 22709 14231 22743 14265
rect 22777 14231 22811 14265
rect 22845 14231 22879 14265
rect 22913 14231 22947 14265
rect 22981 14231 23015 14265
rect 23049 14231 23083 14265
rect 23117 14231 23151 14265
rect 23185 14231 23219 14265
rect 23253 14231 23287 14265
rect 23321 14231 23355 14265
rect 23389 14231 23423 14265
rect 23457 14231 23491 14265
rect 23525 14231 23559 14265
rect 23593 14231 23627 14265
rect 23661 14231 23695 14265
rect 23729 14231 23763 14265
rect 23797 14231 23831 14265
rect 23865 14231 23899 14265
rect 23933 14231 23967 14265
rect 24001 14231 24035 14265
rect 24069 14231 24103 14265
rect 24137 14231 24171 14265
rect 24205 14231 24239 14265
rect 24273 14231 24307 14265
rect 24341 14231 24375 14265
rect 24409 14231 24443 14265
rect 24477 14231 24511 14265
rect 24545 14231 24579 14265
rect 24613 14231 24647 14265
rect 24681 14231 24715 14265
rect 24749 14231 24783 14265
rect 24817 14231 24851 14265
rect 24885 14231 24919 14265
rect 24953 14231 24987 14265
rect 25021 14231 25055 14265
rect 25089 14231 25123 14265
rect 25157 14231 25191 14265
rect 25225 14231 25259 14265
rect 25293 14231 25327 14265
rect 25361 14231 25395 14265
rect 25429 14231 25463 14265
rect 25497 14231 25531 14265
rect 25565 14231 25599 14265
rect 25633 14231 25667 14265
rect 25701 14231 25735 14265
rect 25769 14231 25803 14265
rect 25837 14231 25871 14265
rect 25905 14231 25939 14265
rect 25973 14231 26007 14265
rect 26041 14231 26075 14265
rect 26109 14231 26143 14265
rect 26177 14231 26211 14265
rect 26245 14231 26279 14265
rect 26313 14231 26347 14265
rect 26381 14231 26415 14265
rect 26449 14231 26483 14265
rect 26517 14231 26551 14265
rect 26585 14231 26619 14265
rect 26653 14231 26687 14265
rect 26721 14231 26755 14265
rect 26789 14231 26823 14265
rect 26857 14231 26891 14265
rect 26925 14231 26959 14265
rect 26993 14231 27027 14265
rect 27061 14231 27095 14265
rect 27129 14231 27163 14265
rect 27197 14231 27231 14265
rect 27265 14231 27299 14265
rect 27333 14231 27367 14265
rect 27401 14231 27435 14265
rect 27469 14231 27503 14265
rect 27537 14231 27571 14265
rect 27605 14231 27639 14265
rect 27673 14231 27707 14265
rect 27741 14231 27775 14265
rect 27809 14231 27843 14265
rect 27877 14231 27911 14265
rect 27945 14231 27979 14265
rect 28013 14231 28047 14265
rect 28081 14231 28115 14265
rect 28149 14231 28183 14265
rect 28217 14231 28251 14265
rect 28285 14231 28319 14265
rect 28353 14231 28387 14265
rect 28421 14231 28455 14265
rect 28489 14231 28523 14265
rect 28557 14231 28591 14265
rect 28625 14231 28659 14265
rect 28693 14231 28727 14265
rect 28761 14231 28795 14265
rect 28829 14231 28863 14265
rect 28897 14231 28931 14265
rect 28965 14231 28999 14265
rect 29033 14231 29067 14265
rect 29101 14231 29135 14265
rect 29169 14231 29203 14265
rect 29237 14231 29271 14265
rect 29305 14231 29339 14265
rect 29373 14231 29407 14265
rect 29441 14231 29475 14265
rect 29509 14231 29543 14265
rect 29577 14231 29611 14265
rect 29645 14231 29669 14265
rect 18281 14208 29669 14231
rect 7107 14172 7129 14206
rect 7163 14172 7269 14206
rect 7137 13785 7269 14172
rect 15831 14205 29669 14208
rect 15831 14171 15855 14205
rect 15889 14171 15925 14205
rect 15959 14171 15995 14205
rect 16029 14171 16065 14205
rect 16099 14171 16135 14205
rect 16169 14171 16205 14205
rect 16239 14171 16275 14205
rect 16309 14171 16345 14205
rect 16379 14171 16415 14205
rect 16449 14171 16485 14205
rect 16519 14171 16555 14205
rect 16589 14171 16625 14205
rect 16659 14171 16695 14205
rect 16729 14171 16765 14205
rect 16799 14171 16835 14205
rect 16869 14171 16904 14205
rect 16938 14171 16973 14205
rect 17007 14171 17042 14205
rect 17076 14171 17111 14205
rect 17145 14171 17180 14205
rect 17214 14171 17249 14205
rect 17283 14171 17318 14205
rect 17352 14171 17387 14205
rect 17421 14171 17456 14205
rect 17490 14171 17525 14205
rect 17559 14171 17594 14205
rect 17628 14171 17663 14205
rect 17697 14171 17732 14205
rect 17766 14171 17801 14205
rect 17835 14171 17870 14205
rect 17904 14171 17939 14205
rect 17973 14171 18008 14205
rect 18042 14171 18077 14205
rect 18111 14171 18146 14205
rect 18180 14171 18215 14205
rect 18249 14171 18284 14205
rect 18318 14202 29669 14205
rect 18318 14171 18356 14202
rect 15831 14168 18356 14171
rect 18390 14199 29669 14202
rect 18390 14168 18428 14199
rect 15831 14165 18428 14168
rect 18462 14196 29669 14199
rect 18462 14165 18500 14196
rect 15831 14162 18500 14165
rect 18534 14193 29669 14196
rect 18534 14162 18572 14193
rect 15831 14159 18572 14162
rect 18606 14159 18641 14193
rect 18675 14159 18710 14193
rect 18744 14159 18779 14193
rect 18813 14159 18848 14193
rect 18882 14159 18917 14193
rect 18951 14159 18986 14193
rect 19020 14159 19055 14193
rect 19089 14159 19124 14193
rect 19158 14159 19193 14193
rect 19227 14159 19262 14193
rect 19296 14159 19331 14193
rect 19365 14159 19400 14193
rect 19434 14159 19469 14193
rect 19503 14159 19538 14193
rect 19572 14159 19607 14193
rect 19641 14159 19676 14193
rect 19710 14159 19745 14193
rect 19779 14159 19814 14193
rect 19848 14159 19883 14193
rect 19917 14159 19952 14193
rect 19986 14159 20021 14193
rect 20055 14159 20090 14193
rect 20124 14159 20159 14193
rect 20193 14159 20227 14193
rect 20261 14159 20295 14193
rect 20329 14159 20363 14193
rect 20397 14159 20431 14193
rect 20465 14159 20499 14193
rect 20533 14159 20567 14193
rect 20601 14159 20635 14193
rect 20669 14159 20703 14193
rect 20737 14159 20771 14193
rect 20805 14159 20839 14193
rect 20873 14159 20907 14193
rect 20941 14159 20975 14193
rect 21009 14159 21043 14193
rect 21077 14159 21111 14193
rect 21145 14159 21179 14193
rect 21213 14159 21247 14193
rect 21281 14159 21315 14193
rect 21349 14159 21383 14193
rect 21417 14159 21451 14193
rect 21485 14159 21519 14193
rect 21553 14159 21587 14193
rect 21621 14159 21655 14193
rect 21689 14159 21723 14193
rect 21757 14159 21791 14193
rect 21825 14159 21859 14193
rect 21893 14159 21927 14193
rect 21961 14159 21995 14193
rect 22029 14159 22063 14193
rect 22097 14159 22131 14193
rect 22165 14159 22199 14193
rect 22233 14159 22267 14193
rect 22301 14159 22335 14193
rect 22369 14159 22403 14193
rect 22437 14159 22471 14193
rect 22505 14159 22539 14193
rect 22573 14159 22607 14193
rect 22641 14159 22675 14193
rect 22709 14159 22743 14193
rect 22777 14159 22811 14193
rect 22845 14159 22879 14193
rect 22913 14159 22947 14193
rect 22981 14159 23015 14193
rect 23049 14159 23083 14193
rect 23117 14159 23151 14193
rect 23185 14159 23219 14193
rect 23253 14159 23287 14193
rect 23321 14159 23355 14193
rect 23389 14159 23423 14193
rect 23457 14159 23491 14193
rect 23525 14159 23559 14193
rect 23593 14159 23627 14193
rect 23661 14159 23695 14193
rect 23729 14159 23763 14193
rect 23797 14159 23831 14193
rect 23865 14159 23899 14193
rect 23933 14159 23967 14193
rect 24001 14159 24035 14193
rect 24069 14159 24103 14193
rect 24137 14159 24171 14193
rect 24205 14159 24239 14193
rect 24273 14159 24307 14193
rect 24341 14159 24375 14193
rect 24409 14159 24443 14193
rect 24477 14159 24511 14193
rect 24545 14159 24579 14193
rect 24613 14159 24647 14193
rect 24681 14159 24715 14193
rect 24749 14159 24783 14193
rect 24817 14159 24851 14193
rect 24885 14159 24919 14193
rect 24953 14159 24987 14193
rect 25021 14159 25055 14193
rect 25089 14159 25123 14193
rect 25157 14159 25191 14193
rect 25225 14159 25259 14193
rect 25293 14159 25327 14193
rect 25361 14159 25395 14193
rect 25429 14159 25463 14193
rect 25497 14159 25531 14193
rect 25565 14159 25599 14193
rect 25633 14159 25667 14193
rect 25701 14159 25735 14193
rect 25769 14159 25803 14193
rect 25837 14159 25871 14193
rect 25905 14159 25939 14193
rect 25973 14159 26007 14193
rect 26041 14159 26075 14193
rect 26109 14159 26143 14193
rect 26177 14159 26211 14193
rect 26245 14159 26279 14193
rect 26313 14159 26347 14193
rect 26381 14159 26415 14193
rect 26449 14159 26483 14193
rect 26517 14159 26551 14193
rect 26585 14159 26619 14193
rect 26653 14159 26687 14193
rect 26721 14159 26755 14193
rect 26789 14159 26823 14193
rect 26857 14159 26891 14193
rect 26925 14159 26959 14193
rect 26993 14159 27027 14193
rect 27061 14159 27095 14193
rect 27129 14159 27163 14193
rect 27197 14159 27231 14193
rect 27265 14159 27299 14193
rect 27333 14159 27367 14193
rect 27401 14159 27435 14193
rect 27469 14159 27503 14193
rect 27537 14159 27571 14193
rect 27605 14159 27639 14193
rect 27673 14159 27707 14193
rect 27741 14159 27775 14193
rect 27809 14159 27843 14193
rect 27877 14159 27911 14193
rect 27945 14159 27979 14193
rect 28013 14159 28047 14193
rect 28081 14159 28115 14193
rect 28149 14159 28183 14193
rect 28217 14159 28251 14193
rect 28285 14159 28319 14193
rect 28353 14159 28387 14193
rect 28421 14159 28455 14193
rect 28489 14159 28523 14193
rect 28557 14159 28591 14193
rect 28625 14159 28659 14193
rect 28693 14159 28727 14193
rect 28761 14159 28795 14193
rect 28829 14159 28863 14193
rect 28897 14159 28931 14193
rect 28965 14159 28999 14193
rect 29033 14159 29067 14193
rect 29101 14159 29135 14193
rect 29169 14159 29203 14193
rect 29237 14159 29271 14193
rect 29305 14159 29339 14193
rect 29373 14159 29407 14193
rect 29441 14159 29475 14193
rect 29509 14159 29543 14193
rect 29577 14159 29611 14193
rect 29645 14159 29669 14193
rect 15831 14133 29669 14159
rect 15831 14099 15855 14133
rect 15889 14099 15925 14133
rect 15959 14099 15995 14133
rect 16029 14099 16065 14133
rect 16099 14099 16135 14133
rect 16169 14099 16205 14133
rect 16239 14099 16275 14133
rect 16309 14099 16345 14133
rect 16379 14099 16415 14133
rect 16449 14099 16485 14133
rect 16519 14099 16555 14133
rect 16589 14099 16625 14133
rect 16659 14099 16695 14133
rect 16729 14099 16765 14133
rect 16799 14099 16835 14133
rect 16869 14099 16905 14133
rect 16939 14099 16975 14133
rect 17009 14099 17045 14133
rect 17079 14099 17114 14133
rect 17148 14099 17183 14133
rect 17217 14099 17252 14133
rect 17286 14099 17321 14133
rect 17355 14099 17390 14133
rect 17424 14099 17459 14133
rect 17493 14099 17528 14133
rect 17562 14099 17597 14133
rect 17631 14099 17666 14133
rect 17700 14099 17735 14133
rect 17769 14099 17804 14133
rect 17838 14099 17873 14133
rect 17907 14099 17942 14133
rect 17976 14099 18011 14133
rect 18045 14099 18080 14133
rect 18114 14099 18149 14133
rect 18183 14099 18218 14133
rect 18252 14099 18287 14133
rect 18321 14099 18356 14133
rect 18390 14130 29669 14133
rect 18390 14099 18428 14130
rect 15831 14096 18428 14099
rect 18462 14127 29669 14130
rect 18462 14096 18500 14127
rect 15831 14093 18500 14096
rect 18534 14124 29669 14127
rect 18534 14093 18572 14124
rect 15831 14090 18572 14093
rect 18606 14121 29669 14124
rect 18606 14090 18644 14121
rect 15831 14087 18644 14090
rect 18678 14087 18713 14121
rect 18747 14087 18782 14121
rect 18816 14087 18851 14121
rect 18885 14087 18920 14121
rect 18954 14087 18989 14121
rect 19023 14087 19058 14121
rect 19092 14087 19127 14121
rect 19161 14087 19196 14121
rect 19230 14087 19265 14121
rect 19299 14087 19334 14121
rect 19368 14087 19403 14121
rect 19437 14087 19472 14121
rect 19506 14087 19541 14121
rect 19575 14087 19610 14121
rect 19644 14087 19679 14121
rect 19713 14087 19748 14121
rect 19782 14087 19817 14121
rect 19851 14087 19886 14121
rect 19920 14087 19955 14121
rect 19989 14087 20023 14121
rect 20057 14087 20091 14121
rect 20125 14087 20159 14121
rect 20193 14087 20227 14121
rect 20261 14087 20295 14121
rect 20329 14087 20363 14121
rect 20397 14087 20431 14121
rect 20465 14087 20499 14121
rect 20533 14087 20567 14121
rect 20601 14087 20635 14121
rect 20669 14087 20703 14121
rect 20737 14087 20771 14121
rect 20805 14087 20839 14121
rect 20873 14087 20907 14121
rect 20941 14087 20975 14121
rect 21009 14087 21043 14121
rect 21077 14087 21111 14121
rect 21145 14087 21179 14121
rect 21213 14087 21247 14121
rect 21281 14087 21315 14121
rect 21349 14087 21383 14121
rect 21417 14087 21451 14121
rect 21485 14087 21519 14121
rect 21553 14087 21587 14121
rect 21621 14087 21655 14121
rect 21689 14087 21723 14121
rect 21757 14087 21791 14121
rect 21825 14087 21859 14121
rect 21893 14087 21927 14121
rect 21961 14087 21995 14121
rect 22029 14087 22063 14121
rect 22097 14087 22131 14121
rect 22165 14087 22199 14121
rect 22233 14087 22267 14121
rect 22301 14087 22335 14121
rect 22369 14087 22403 14121
rect 22437 14087 22471 14121
rect 22505 14087 22539 14121
rect 22573 14087 22607 14121
rect 22641 14087 22675 14121
rect 22709 14087 22743 14121
rect 22777 14087 22811 14121
rect 22845 14087 22879 14121
rect 22913 14087 22947 14121
rect 22981 14087 23015 14121
rect 23049 14087 23083 14121
rect 23117 14087 23151 14121
rect 23185 14087 23219 14121
rect 23253 14087 23287 14121
rect 23321 14087 23355 14121
rect 23389 14087 23423 14121
rect 23457 14087 23491 14121
rect 23525 14087 23559 14121
rect 23593 14087 23627 14121
rect 23661 14087 23695 14121
rect 23729 14087 23763 14121
rect 23797 14087 23831 14121
rect 23865 14087 23899 14121
rect 23933 14087 23967 14121
rect 24001 14087 24035 14121
rect 24069 14087 24103 14121
rect 24137 14087 24171 14121
rect 24205 14087 24239 14121
rect 24273 14087 24307 14121
rect 24341 14087 24375 14121
rect 24409 14087 24443 14121
rect 24477 14087 24511 14121
rect 24545 14087 24579 14121
rect 24613 14087 24647 14121
rect 24681 14087 24715 14121
rect 24749 14087 24783 14121
rect 24817 14087 24851 14121
rect 24885 14087 24919 14121
rect 24953 14087 24987 14121
rect 25021 14087 25055 14121
rect 25089 14087 25123 14121
rect 25157 14087 25191 14121
rect 25225 14087 25259 14121
rect 25293 14087 25327 14121
rect 25361 14087 25395 14121
rect 25429 14087 25463 14121
rect 25497 14087 25531 14121
rect 25565 14087 25599 14121
rect 25633 14087 25667 14121
rect 25701 14087 25735 14121
rect 25769 14087 25803 14121
rect 25837 14087 25871 14121
rect 25905 14087 25939 14121
rect 25973 14087 26007 14121
rect 26041 14087 26075 14121
rect 26109 14087 26143 14121
rect 26177 14087 26211 14121
rect 26245 14087 26279 14121
rect 26313 14087 26347 14121
rect 26381 14087 26415 14121
rect 26449 14087 26483 14121
rect 26517 14087 26551 14121
rect 26585 14087 26619 14121
rect 26653 14087 26687 14121
rect 26721 14087 26755 14121
rect 26789 14087 26823 14121
rect 26857 14087 26891 14121
rect 26925 14087 26959 14121
rect 26993 14087 27027 14121
rect 27061 14087 27095 14121
rect 27129 14087 27163 14121
rect 27197 14087 27231 14121
rect 27265 14087 27299 14121
rect 27333 14087 27367 14121
rect 27401 14087 27435 14121
rect 27469 14087 27503 14121
rect 27537 14087 27571 14121
rect 27605 14087 27639 14121
rect 27673 14087 27707 14121
rect 27741 14087 27775 14121
rect 27809 14087 27843 14121
rect 27877 14087 27911 14121
rect 27945 14087 27979 14121
rect 28013 14087 28047 14121
rect 28081 14087 28115 14121
rect 28149 14087 28183 14121
rect 28217 14087 28251 14121
rect 28285 14087 28319 14121
rect 28353 14087 28387 14121
rect 28421 14087 28455 14121
rect 28489 14087 28523 14121
rect 28557 14087 28591 14121
rect 28625 14087 28659 14121
rect 28693 14087 28727 14121
rect 28761 14087 28795 14121
rect 28829 14087 28863 14121
rect 28897 14087 28931 14121
rect 28965 14087 28999 14121
rect 29033 14087 29067 14121
rect 29101 14087 29135 14121
rect 29169 14087 29203 14121
rect 29237 14087 29271 14121
rect 29305 14087 29339 14121
rect 29373 14087 29407 14121
rect 29441 14087 29475 14121
rect 29509 14087 29543 14121
rect 29577 14087 29611 14121
rect 29645 14087 29669 14121
rect 15831 14084 29669 14087
rect 15831 14061 18681 14084
rect 15831 14027 15855 14061
rect 15889 14027 15925 14061
rect 15959 14027 15995 14061
rect 16029 14027 16065 14061
rect 16099 14027 16135 14061
rect 16169 14027 16205 14061
rect 16239 14027 16275 14061
rect 16309 14027 16345 14061
rect 16379 14027 16415 14061
rect 16449 14027 16485 14061
rect 16519 14027 16555 14061
rect 16589 14027 16625 14061
rect 16659 14027 16695 14061
rect 16729 14027 16765 14061
rect 16799 14027 16835 14061
rect 16869 14027 16905 14061
rect 16939 14027 16975 14061
rect 17009 14027 17045 14061
rect 17079 14027 17115 14061
rect 17149 14027 17185 14061
rect 17219 14027 17255 14061
rect 17289 14027 17324 14061
rect 17358 14027 17393 14061
rect 17427 14027 17462 14061
rect 17496 14027 17531 14061
rect 17565 14027 17600 14061
rect 17634 14027 17669 14061
rect 17703 14027 17738 14061
rect 17772 14027 17807 14061
rect 17841 14027 17876 14061
rect 17910 14027 17945 14061
rect 17979 14027 18014 14061
rect 18048 14027 18083 14061
rect 18117 14027 18152 14061
rect 18186 14027 18221 14061
rect 18255 14027 18290 14061
rect 18324 14027 18359 14061
rect 18393 14027 18428 14061
rect 18462 14058 18681 14061
rect 18462 14027 18500 14058
rect 15831 14024 18500 14027
rect 18534 14055 18681 14058
rect 18534 14024 18572 14055
rect 15831 14021 18572 14024
rect 18606 14051 18681 14055
rect 18606 14021 18644 14051
rect 15831 14017 18644 14021
rect 18678 14017 18681 14051
rect 15831 13989 18681 14017
rect 15831 13955 15855 13989
rect 15889 13955 15925 13989
rect 15959 13955 15995 13989
rect 16029 13955 16065 13989
rect 16099 13955 16135 13989
rect 16169 13955 16205 13989
rect 16239 13955 16275 13989
rect 16309 13955 16345 13989
rect 16379 13955 16415 13989
rect 16449 13955 16485 13989
rect 16519 13955 16555 13989
rect 16589 13955 16625 13989
rect 16659 13955 16695 13989
rect 16729 13955 16765 13989
rect 16799 13955 16835 13989
rect 16869 13955 16905 13989
rect 16939 13955 16975 13989
rect 17009 13955 17045 13989
rect 17079 13955 17115 13989
rect 17149 13955 17185 13989
rect 17219 13955 17255 13989
rect 17289 13955 17325 13989
rect 17359 13955 17395 13989
rect 17429 13955 17465 13989
rect 17499 13955 17534 13989
rect 17568 13955 17603 13989
rect 17637 13955 17672 13989
rect 17706 13955 17741 13989
rect 17775 13955 17810 13989
rect 17844 13955 17879 13989
rect 17913 13955 17948 13989
rect 17982 13955 18017 13989
rect 18051 13955 18086 13989
rect 18120 13955 18155 13989
rect 18189 13955 18224 13989
rect 18258 13955 18293 13989
rect 18327 13955 18362 13989
rect 18396 13955 18431 13989
rect 18465 13955 18500 13989
rect 18534 13986 18681 13989
rect 18534 13955 18572 13986
rect 15831 13952 18572 13955
rect 18606 13981 18681 13986
rect 18606 13952 18644 13981
rect 15831 13947 18644 13952
rect 18678 13947 18681 13981
rect 15831 13917 18681 13947
rect 15831 13883 15855 13917
rect 15889 13883 15925 13917
rect 15959 13883 15995 13917
rect 16029 13883 16065 13917
rect 16099 13883 16135 13917
rect 16169 13883 16205 13917
rect 16239 13883 16275 13917
rect 16309 13883 16345 13917
rect 16379 13883 16415 13917
rect 16449 13883 16485 13917
rect 16519 13883 16555 13917
rect 16589 13883 16625 13917
rect 16659 13883 16695 13917
rect 16729 13883 16765 13917
rect 16799 13883 16835 13917
rect 16869 13883 16905 13917
rect 16939 13883 16975 13917
rect 17009 13883 17045 13917
rect 17079 13883 17115 13917
rect 17149 13883 17185 13917
rect 17219 13883 17255 13917
rect 17289 13883 17325 13917
rect 17359 13883 17395 13917
rect 17429 13883 17465 13917
rect 17499 13883 17535 13917
rect 17569 13883 17605 13917
rect 17639 13883 17675 13917
rect 17709 13883 17744 13917
rect 17778 13883 17813 13917
rect 17847 13883 17882 13917
rect 17916 13883 17951 13917
rect 17985 13883 18020 13917
rect 18054 13883 18089 13917
rect 18123 13883 18158 13917
rect 18192 13883 18227 13917
rect 18261 13883 18296 13917
rect 18330 13883 18365 13917
rect 18399 13883 18434 13917
rect 18468 13883 18503 13917
rect 18537 13883 18572 13917
rect 18606 13910 18681 13917
rect 18606 13883 18644 13910
rect 15831 13876 18644 13883
rect 18678 13876 18681 13910
rect 15831 13845 18681 13876
rect 15831 13811 15855 13845
rect 15889 13811 15924 13845
rect 15958 13811 15993 13845
rect 16027 13811 16062 13845
rect 16096 13811 16131 13845
rect 16165 13811 16199 13845
rect 16233 13811 16267 13845
rect 16301 13811 16335 13845
rect 16369 13811 16403 13845
rect 16437 13811 16471 13845
rect 16505 13811 16539 13845
rect 16573 13811 16607 13845
rect 16641 13811 16675 13845
rect 16709 13811 16743 13845
rect 16777 13811 16811 13845
rect 16845 13811 16879 13845
rect 16913 13811 16947 13845
rect 16981 13811 17015 13845
rect 17049 13811 17083 13845
rect 17117 13811 17151 13845
rect 17185 13811 17219 13845
rect 17253 13811 17287 13845
rect 17321 13811 17355 13845
rect 17389 13811 17423 13845
rect 17457 13811 17491 13845
rect 17525 13811 17559 13845
rect 17593 13811 17627 13845
rect 17661 13811 17695 13845
rect 17729 13811 17763 13845
rect 17797 13811 17831 13845
rect 17865 13811 17899 13845
rect 17933 13811 17967 13845
rect 18001 13811 18035 13845
rect 18069 13811 18103 13845
rect 18137 13811 18171 13845
rect 18205 13811 18239 13845
rect 18273 13811 18307 13845
rect 18341 13811 18375 13845
rect 18409 13811 18443 13845
rect 18477 13811 18511 13845
rect 18545 13811 18579 13845
rect 18613 13811 18681 13845
rect 15831 13808 18681 13811
rect 15225 12121 15968 12238
rect 13224 12087 13279 12121
rect 13313 12087 13347 12121
rect 13381 12087 13415 12121
rect 13449 12087 13483 12121
rect 13517 12087 13551 12121
rect 13585 12087 13619 12121
rect 13653 12087 13687 12121
rect 13721 12087 13755 12121
rect 13789 12087 13823 12121
rect 13857 12087 13891 12121
rect 13925 12087 13959 12121
rect 13993 12087 14027 12121
rect 14061 12087 14095 12121
rect 14129 12087 14163 12121
rect 14197 12087 14231 12121
rect 14265 12087 14299 12121
rect 14333 12087 14367 12121
rect 14401 12087 14435 12121
rect 14469 12087 14503 12121
rect 14537 12087 14571 12121
rect 14605 12087 14639 12121
rect 14673 12087 14707 12121
rect 14741 12087 14775 12121
rect 14809 12087 14843 12121
rect 14877 12087 14911 12121
rect 14945 12087 14979 12121
rect 15013 12087 15047 12121
rect 15081 12087 15115 12121
rect 15149 12087 15183 12121
rect 15217 12087 15251 12121
rect 15285 12087 15319 12121
rect 15353 12087 15387 12121
rect 15421 12087 15455 12121
rect 15489 12087 15523 12121
rect 15557 12087 15591 12121
rect 15625 12087 15659 12121
rect 15693 12087 15727 12121
rect 15761 12087 15795 12121
rect 15829 12087 15968 12121
rect 13224 12052 15968 12087
rect 13224 12018 13279 12052
rect 13313 12018 13347 12052
rect 13381 12018 13415 12052
rect 13449 12018 13483 12052
rect 13517 12018 13551 12052
rect 13585 12018 13619 12052
rect 13653 12018 13687 12052
rect 13721 12018 13755 12052
rect 13789 12018 13823 12052
rect 13857 12018 13891 12052
rect 13925 12018 13959 12052
rect 13993 12018 14027 12052
rect 14061 12018 14095 12052
rect 14129 12018 14163 12052
rect 14197 12018 14231 12052
rect 14265 12018 14299 12052
rect 14333 12018 14367 12052
rect 14401 12018 14435 12052
rect 14469 12018 14503 12052
rect 14537 12018 14571 12052
rect 14605 12018 14639 12052
rect 14673 12018 14707 12052
rect 14741 12018 14775 12052
rect 14809 12018 14843 12052
rect 14877 12018 14911 12052
rect 14945 12018 14979 12052
rect 15013 12018 15047 12052
rect 15081 12018 15115 12052
rect 15149 12018 15183 12052
rect 15217 12018 15251 12052
rect 15285 12018 15319 12052
rect 15353 12018 15387 12052
rect 15421 12018 15455 12052
rect 15489 12018 15523 12052
rect 15557 12018 15591 12052
rect 15625 12018 15659 12052
rect 15693 12018 15727 12052
rect 15761 12018 15795 12052
rect 15829 12043 15968 12052
rect 15829 12018 15884 12043
rect 13224 11983 15884 12018
rect 13224 11949 13279 11983
rect 13313 11949 13347 11983
rect 13381 11949 13415 11983
rect 13449 11949 13483 11983
rect 13517 11949 13551 11983
rect 13585 11949 13619 11983
rect 13653 11949 13687 11983
rect 13721 11949 13755 11983
rect 13789 11949 13823 11983
rect 13857 11949 13891 11983
rect 13925 11949 13959 11983
rect 13993 11949 14027 11983
rect 14061 11949 14095 11983
rect 14129 11949 14163 11983
rect 14197 11949 14231 11983
rect 14265 11949 14299 11983
rect 14333 11949 14367 11983
rect 14401 11949 14435 11983
rect 14469 11949 14503 11983
rect 14537 11949 14571 11983
rect 14605 11949 14639 11983
rect 14673 11949 14707 11983
rect 14741 11949 14775 11983
rect 14809 11949 14843 11983
rect 14877 11949 14911 11983
rect 14945 11949 14979 11983
rect 15013 11949 15047 11983
rect 15081 11949 15115 11983
rect 15149 11949 15183 11983
rect 15217 11949 15251 11983
rect 15285 11949 15319 11983
rect 15353 11949 15387 11983
rect 15421 11949 15455 11983
rect 15489 11949 15523 11983
rect 15557 11949 15591 11983
rect 15625 11949 15659 11983
rect 15693 11949 15727 11983
rect 15761 11949 15795 11983
rect 15829 11949 15884 11983
rect -2966 10378 -266 10413
rect -2966 10344 -2959 10378
rect -2925 10344 -2891 10378
rect -2857 10344 -2823 10378
rect -2789 10344 -2755 10378
rect -2721 10344 -2687 10378
rect -2653 10344 -2619 10378
rect -2585 10344 -2551 10378
rect -2517 10344 -2483 10378
rect -2449 10344 -2415 10378
rect -2381 10344 -2347 10378
rect -2313 10344 -2279 10378
rect -2245 10344 -2211 10378
rect -2177 10344 -2143 10378
rect -2109 10344 -2075 10378
rect -2041 10344 -2007 10378
rect -1973 10344 -1939 10378
rect -1905 10344 -1871 10378
rect -1837 10344 -1803 10378
rect -1769 10344 -1735 10378
rect -1701 10344 -1667 10378
rect -1633 10344 -1599 10378
rect -1565 10344 -1531 10378
rect -1497 10344 -1463 10378
rect -1429 10344 -1395 10378
rect -1361 10344 -1327 10378
rect -1293 10344 -1259 10378
rect -1225 10344 -1191 10378
rect -1157 10344 -1123 10378
rect -1089 10344 -1055 10378
rect -1021 10344 -987 10378
rect -953 10344 -919 10378
rect -885 10344 -851 10378
rect -817 10344 -783 10378
rect -749 10344 -715 10378
rect -681 10344 -647 10378
rect -613 10344 -579 10378
rect -545 10344 -511 10378
rect -477 10344 -443 10378
rect -409 10344 -375 10378
rect -341 10344 -307 10378
rect -273 10344 -266 10378
rect -2966 10309 -266 10344
rect -2966 10275 -2959 10309
rect -2925 10275 -2891 10309
rect -2857 10275 -2823 10309
rect -2789 10275 -2755 10309
rect -2721 10275 -2687 10309
rect -2653 10275 -2619 10309
rect -2585 10275 -2551 10309
rect -2517 10275 -2483 10309
rect -2449 10275 -2415 10309
rect -2381 10275 -2347 10309
rect -2313 10275 -2279 10309
rect -2245 10275 -2211 10309
rect -2177 10275 -2143 10309
rect -2109 10275 -2075 10309
rect -2041 10275 -2007 10309
rect -1973 10275 -1939 10309
rect -1905 10275 -1871 10309
rect -1837 10275 -1803 10309
rect -1769 10275 -1735 10309
rect -1701 10275 -1667 10309
rect -1633 10275 -1599 10309
rect -1565 10275 -1531 10309
rect -1497 10275 -1463 10309
rect -1429 10275 -1395 10309
rect -1361 10275 -1327 10309
rect -1293 10275 -1259 10309
rect -1225 10275 -1191 10309
rect -1157 10275 -1123 10309
rect -1089 10275 -1055 10309
rect -1021 10275 -987 10309
rect -953 10275 -919 10309
rect -885 10275 -851 10309
rect -817 10275 -783 10309
rect -749 10275 -715 10309
rect -681 10275 -647 10309
rect -613 10275 -579 10309
rect -545 10275 -511 10309
rect -477 10275 -443 10309
rect -409 10275 -375 10309
rect -341 10275 -307 10309
rect -273 10275 -266 10309
rect -2966 10240 -266 10275
rect -2966 10206 -2959 10240
rect -2925 10206 -2891 10240
rect -2857 10206 -2823 10240
rect -2789 10206 -2755 10240
rect -2721 10206 -2687 10240
rect -2653 10206 -2619 10240
rect -2585 10206 -2551 10240
rect -2517 10206 -2483 10240
rect -2449 10206 -2415 10240
rect -2381 10206 -2347 10240
rect -2313 10206 -2279 10240
rect -2245 10206 -2211 10240
rect -2177 10206 -2143 10240
rect -2109 10206 -2075 10240
rect -2041 10206 -2007 10240
rect -1973 10206 -1939 10240
rect -1905 10206 -1871 10240
rect -1837 10206 -1803 10240
rect -1769 10206 -1735 10240
rect -1701 10206 -1667 10240
rect -1633 10206 -1599 10240
rect -1565 10206 -1531 10240
rect -1497 10206 -1463 10240
rect -1429 10206 -1395 10240
rect -1361 10206 -1327 10240
rect -1293 10206 -1259 10240
rect -1225 10206 -1191 10240
rect -1157 10206 -1123 10240
rect -1089 10206 -1055 10240
rect -1021 10206 -987 10240
rect -953 10206 -919 10240
rect -885 10206 -851 10240
rect -817 10206 -783 10240
rect -749 10206 -715 10240
rect -681 10206 -647 10240
rect -613 10206 -579 10240
rect -545 10206 -511 10240
rect -477 10206 -443 10240
rect -409 10206 -375 10240
rect -341 10206 -307 10240
rect -273 10206 -266 10240
rect -2966 10171 -266 10206
rect -2966 10137 -2959 10171
rect -2925 10137 -2891 10171
rect -2857 10137 -2823 10171
rect -2789 10137 -2755 10171
rect -2721 10137 -2687 10171
rect -2653 10137 -2619 10171
rect -2585 10137 -2551 10171
rect -2517 10137 -2483 10171
rect -2449 10137 -2415 10171
rect -2381 10137 -2347 10171
rect -2313 10137 -2279 10171
rect -2245 10137 -2211 10171
rect -2177 10137 -2143 10171
rect -2109 10137 -2075 10171
rect -2041 10137 -2007 10171
rect -1973 10137 -1939 10171
rect -1905 10137 -1871 10171
rect -1837 10137 -1803 10171
rect -1769 10137 -1735 10171
rect -1701 10137 -1667 10171
rect -1633 10137 -1599 10171
rect -1565 10137 -1531 10171
rect -1497 10137 -1463 10171
rect -1429 10137 -1395 10171
rect -1361 10137 -1327 10171
rect -1293 10137 -1259 10171
rect -1225 10137 -1191 10171
rect -1157 10137 -1123 10171
rect -1089 10137 -1055 10171
rect -1021 10137 -987 10171
rect -953 10137 -919 10171
rect -885 10137 -851 10171
rect -817 10137 -783 10171
rect -749 10137 -715 10171
rect -681 10137 -647 10171
rect -613 10137 -579 10171
rect -545 10137 -511 10171
rect -477 10137 -443 10171
rect -409 10137 -375 10171
rect -341 10137 -307 10171
rect -273 10137 -266 10171
rect -2966 10102 -266 10137
rect -2966 10068 -2959 10102
rect -2925 10068 -2891 10102
rect -2857 10068 -2823 10102
rect -2789 10068 -2755 10102
rect -2721 10068 -2687 10102
rect -2653 10068 -2619 10102
rect -2585 10068 -2551 10102
rect -2517 10068 -2483 10102
rect -2449 10068 -2415 10102
rect -2381 10068 -2347 10102
rect -2313 10068 -2279 10102
rect -2245 10068 -2211 10102
rect -2177 10068 -2143 10102
rect -2109 10068 -2075 10102
rect -2041 10068 -2007 10102
rect -1973 10068 -1939 10102
rect -1905 10068 -1871 10102
rect -1837 10068 -1803 10102
rect -1769 10068 -1735 10102
rect -1701 10068 -1667 10102
rect -1633 10068 -1599 10102
rect -1565 10068 -1531 10102
rect -1497 10068 -1463 10102
rect -1429 10068 -1395 10102
rect -1361 10068 -1327 10102
rect -1293 10068 -1259 10102
rect -1225 10068 -1191 10102
rect -1157 10068 -1123 10102
rect -1089 10068 -1055 10102
rect -1021 10068 -987 10102
rect -953 10068 -919 10102
rect -885 10068 -851 10102
rect -817 10068 -783 10102
rect -749 10068 -715 10102
rect -681 10068 -647 10102
rect -613 10068 -579 10102
rect -545 10068 -511 10102
rect -477 10068 -443 10102
rect -409 10068 -375 10102
rect -341 10068 -307 10102
rect -273 10068 -266 10102
rect -2966 10033 -266 10068
rect 4421 11910 6239 11934
rect 4421 11332 4429 11910
rect 6231 11332 6239 11910
rect 4421 11297 6239 11332
rect 4421 11263 4429 11297
rect 4463 11263 4497 11297
rect 4531 11263 4565 11297
rect 4599 11263 4633 11297
rect 4667 11263 4701 11297
rect 4735 11263 4769 11297
rect 4803 11263 4837 11297
rect 4871 11263 4905 11297
rect 4939 11263 4973 11297
rect 5007 11263 5041 11297
rect 5075 11263 5109 11297
rect 5143 11263 5177 11297
rect 5211 11263 5245 11297
rect 5279 11263 5313 11297
rect 5347 11263 5381 11297
rect 5415 11263 5449 11297
rect 5483 11263 5517 11297
rect 5551 11263 5585 11297
rect 5619 11263 5653 11297
rect 5687 11263 5721 11297
rect 5755 11263 5789 11297
rect 5823 11263 5857 11297
rect 5891 11263 5925 11297
rect 5959 11263 5993 11297
rect 6027 11263 6061 11297
rect 6095 11263 6129 11297
rect 6163 11263 6197 11297
rect 6231 11263 6239 11297
rect 13224 11914 15884 11949
rect 13224 11880 13279 11914
rect 13313 11880 13347 11914
rect 13381 11880 13415 11914
rect 13449 11880 13483 11914
rect 13517 11880 13551 11914
rect 13585 11880 13619 11914
rect 13653 11880 13687 11914
rect 13721 11880 13755 11914
rect 13789 11880 13823 11914
rect 13857 11880 13891 11914
rect 13925 11880 13959 11914
rect 13993 11880 14027 11914
rect 14061 11880 14095 11914
rect 14129 11880 14163 11914
rect 14197 11880 14231 11914
rect 14265 11880 14299 11914
rect 14333 11880 14367 11914
rect 14401 11880 14435 11914
rect 14469 11880 14503 11914
rect 14537 11880 14571 11914
rect 14605 11880 14639 11914
rect 14673 11880 14707 11914
rect 14741 11880 14775 11914
rect 14809 11880 14843 11914
rect 14877 11880 14911 11914
rect 14945 11880 14979 11914
rect 15013 11880 15047 11914
rect 15081 11880 15115 11914
rect 15149 11880 15183 11914
rect 15217 11880 15251 11914
rect 15285 11880 15319 11914
rect 15353 11880 15387 11914
rect 15421 11880 15455 11914
rect 15489 11880 15523 11914
rect 15557 11880 15591 11914
rect 15625 11880 15659 11914
rect 15693 11880 15727 11914
rect 15761 11880 15795 11914
rect 15829 11880 15884 11914
rect 13224 11845 15884 11880
rect 13224 11811 13279 11845
rect 13313 11811 13347 11845
rect 13381 11811 13415 11845
rect 13449 11811 13483 11845
rect 13517 11811 13551 11845
rect 13585 11811 13619 11845
rect 13653 11811 13687 11845
rect 13721 11811 13755 11845
rect 13789 11811 13823 11845
rect 13857 11811 13891 11845
rect 13925 11811 13959 11845
rect 13993 11811 14027 11845
rect 14061 11811 14095 11845
rect 14129 11811 14163 11845
rect 14197 11811 14231 11845
rect 14265 11811 14299 11845
rect 14333 11811 14367 11845
rect 14401 11811 14435 11845
rect 14469 11811 14503 11845
rect 14537 11811 14571 11845
rect 14605 11811 14639 11845
rect 14673 11811 14707 11845
rect 14741 11811 14775 11845
rect 14809 11811 14843 11845
rect 14877 11811 14911 11845
rect 14945 11811 14979 11845
rect 15013 11811 15047 11845
rect 15081 11811 15115 11845
rect 15149 11811 15183 11845
rect 15217 11811 15251 11845
rect 15285 11811 15319 11845
rect 15353 11811 15387 11845
rect 15421 11811 15455 11845
rect 15489 11811 15523 11845
rect 15557 11811 15591 11845
rect 15625 11811 15659 11845
rect 15693 11811 15727 11845
rect 15761 11811 15795 11845
rect 15829 11811 15884 11845
rect 13224 11776 15884 11811
rect 13224 11742 13279 11776
rect 13313 11742 13347 11776
rect 13381 11742 13415 11776
rect 13449 11742 13483 11776
rect 13517 11742 13551 11776
rect 13585 11742 13619 11776
rect 13653 11742 13687 11776
rect 13721 11742 13755 11776
rect 13789 11742 13823 11776
rect 13857 11742 13891 11776
rect 13925 11742 13959 11776
rect 13993 11742 14027 11776
rect 14061 11742 14095 11776
rect 14129 11742 14163 11776
rect 14197 11742 14231 11776
rect 14265 11742 14299 11776
rect 14333 11742 14367 11776
rect 14401 11742 14435 11776
rect 14469 11742 14503 11776
rect 14537 11742 14571 11776
rect 14605 11742 14639 11776
rect 14673 11742 14707 11776
rect 14741 11742 14775 11776
rect 14809 11742 14843 11776
rect 14877 11742 14911 11776
rect 14945 11742 14979 11776
rect 15013 11742 15047 11776
rect 15081 11742 15115 11776
rect 15149 11742 15183 11776
rect 15217 11742 15251 11776
rect 15285 11742 15319 11776
rect 15353 11742 15387 11776
rect 15421 11742 15455 11776
rect 15489 11742 15523 11776
rect 15557 11742 15591 11776
rect 15625 11742 15659 11776
rect 15693 11742 15727 11776
rect 15761 11742 15795 11776
rect 15829 11742 15884 11776
rect 13224 11707 15884 11742
rect 13224 11673 13279 11707
rect 13313 11673 13347 11707
rect 13381 11673 13415 11707
rect 13449 11673 13483 11707
rect 13517 11673 13551 11707
rect 13585 11673 13619 11707
rect 13653 11673 13687 11707
rect 13721 11673 13755 11707
rect 13789 11673 13823 11707
rect 13857 11673 13891 11707
rect 13925 11673 13959 11707
rect 13993 11673 14027 11707
rect 14061 11673 14095 11707
rect 14129 11673 14163 11707
rect 14197 11673 14231 11707
rect 14265 11673 14299 11707
rect 14333 11673 14367 11707
rect 14401 11673 14435 11707
rect 14469 11673 14503 11707
rect 14537 11673 14571 11707
rect 14605 11673 14639 11707
rect 14673 11673 14707 11707
rect 14741 11673 14775 11707
rect 14809 11673 14843 11707
rect 14877 11673 14911 11707
rect 14945 11673 14979 11707
rect 15013 11673 15047 11707
rect 15081 11673 15115 11707
rect 15149 11673 15183 11707
rect 15217 11673 15251 11707
rect 15285 11673 15319 11707
rect 15353 11673 15387 11707
rect 15421 11673 15455 11707
rect 15489 11673 15523 11707
rect 15557 11673 15591 11707
rect 15625 11673 15659 11707
rect 15693 11673 15727 11707
rect 15761 11673 15795 11707
rect 15829 11673 15884 11707
rect 13224 11638 15884 11673
rect 13224 11604 13279 11638
rect 13313 11604 13347 11638
rect 13381 11604 13415 11638
rect 13449 11604 13483 11638
rect 13517 11604 13551 11638
rect 13585 11604 13619 11638
rect 13653 11604 13687 11638
rect 13721 11604 13755 11638
rect 13789 11604 13823 11638
rect 13857 11604 13891 11638
rect 13925 11604 13959 11638
rect 13993 11604 14027 11638
rect 14061 11604 14095 11638
rect 14129 11604 14163 11638
rect 14197 11604 14231 11638
rect 14265 11604 14299 11638
rect 14333 11604 14367 11638
rect 14401 11604 14435 11638
rect 14469 11604 14503 11638
rect 14537 11604 14571 11638
rect 14605 11604 14639 11638
rect 14673 11604 14707 11638
rect 14741 11604 14775 11638
rect 14809 11604 14843 11638
rect 14877 11604 14911 11638
rect 14945 11604 14979 11638
rect 15013 11604 15047 11638
rect 15081 11604 15115 11638
rect 15149 11604 15183 11638
rect 15217 11604 15251 11638
rect 15285 11604 15319 11638
rect 15353 11604 15387 11638
rect 15421 11604 15455 11638
rect 15489 11604 15523 11638
rect 15557 11604 15591 11638
rect 15625 11604 15659 11638
rect 15693 11604 15727 11638
rect 15761 11604 15795 11638
rect 15829 11604 15884 11638
rect 13224 11569 15884 11604
rect 13224 11535 13279 11569
rect 13313 11535 13347 11569
rect 13381 11535 13415 11569
rect 13449 11535 13483 11569
rect 13517 11535 13551 11569
rect 13585 11535 13619 11569
rect 13653 11535 13687 11569
rect 13721 11535 13755 11569
rect 13789 11535 13823 11569
rect 13857 11535 13891 11569
rect 13925 11535 13959 11569
rect 13993 11535 14027 11569
rect 14061 11535 14095 11569
rect 14129 11535 14163 11569
rect 14197 11535 14231 11569
rect 14265 11535 14299 11569
rect 14333 11535 14367 11569
rect 14401 11535 14435 11569
rect 14469 11535 14503 11569
rect 14537 11535 14571 11569
rect 14605 11535 14639 11569
rect 14673 11535 14707 11569
rect 14741 11535 14775 11569
rect 14809 11535 14843 11569
rect 14877 11535 14911 11569
rect 14945 11535 14979 11569
rect 15013 11535 15047 11569
rect 15081 11535 15115 11569
rect 15149 11535 15183 11569
rect 15217 11535 15251 11569
rect 15285 11535 15319 11569
rect 15353 11535 15387 11569
rect 15421 11535 15455 11569
rect 15489 11535 15523 11569
rect 15557 11535 15591 11569
rect 15625 11535 15659 11569
rect 15693 11535 15727 11569
rect 15761 11535 15795 11569
rect 15829 11535 15884 11569
rect 13224 11499 15884 11535
rect 13224 11465 13279 11499
rect 13313 11465 13347 11499
rect 13381 11465 13415 11499
rect 13449 11465 13483 11499
rect 13517 11465 13551 11499
rect 13585 11465 13619 11499
rect 13653 11465 13687 11499
rect 13721 11465 13755 11499
rect 13789 11465 13823 11499
rect 13857 11465 13891 11499
rect 13925 11465 13959 11499
rect 13993 11465 14027 11499
rect 14061 11465 14095 11499
rect 14129 11465 14163 11499
rect 14197 11465 14231 11499
rect 14265 11465 14299 11499
rect 14333 11465 14367 11499
rect 14401 11465 14435 11499
rect 14469 11465 14503 11499
rect 14537 11465 14571 11499
rect 14605 11465 14639 11499
rect 14673 11465 14707 11499
rect 14741 11465 14775 11499
rect 14809 11465 14843 11499
rect 14877 11465 14911 11499
rect 14945 11465 14979 11499
rect 15013 11465 15047 11499
rect 15081 11465 15115 11499
rect 15149 11465 15183 11499
rect 15217 11465 15251 11499
rect 15285 11465 15319 11499
rect 15353 11465 15387 11499
rect 15421 11465 15455 11499
rect 15489 11465 15523 11499
rect 15557 11465 15591 11499
rect 15625 11465 15659 11499
rect 15693 11465 15727 11499
rect 15761 11465 15795 11499
rect 15829 11465 15884 11499
rect 13224 11429 15884 11465
rect 13224 11395 13279 11429
rect 13313 11395 13347 11429
rect 13381 11395 13415 11429
rect 13449 11395 13483 11429
rect 13517 11395 13551 11429
rect 13585 11395 13619 11429
rect 13653 11395 13687 11429
rect 13721 11395 13755 11429
rect 13789 11395 13823 11429
rect 13857 11395 13891 11429
rect 13925 11395 13959 11429
rect 13993 11395 14027 11429
rect 14061 11395 14095 11429
rect 14129 11395 14163 11429
rect 14197 11395 14231 11429
rect 14265 11395 14299 11429
rect 14333 11395 14367 11429
rect 14401 11395 14435 11429
rect 14469 11395 14503 11429
rect 14537 11395 14571 11429
rect 14605 11395 14639 11429
rect 14673 11395 14707 11429
rect 14741 11395 14775 11429
rect 14809 11395 14843 11429
rect 14877 11395 14911 11429
rect 14945 11395 14979 11429
rect 15013 11395 15047 11429
rect 15081 11395 15115 11429
rect 15149 11395 15183 11429
rect 15217 11395 15251 11429
rect 15285 11395 15319 11429
rect 15353 11395 15387 11429
rect 15421 11395 15455 11429
rect 15489 11395 15523 11429
rect 15557 11395 15591 11429
rect 15625 11395 15659 11429
rect 15693 11395 15727 11429
rect 15761 11395 15795 11429
rect 15829 11395 15884 11429
rect 13224 11359 15884 11395
rect 13224 11325 13279 11359
rect 13313 11325 13347 11359
rect 13381 11325 13415 11359
rect 13449 11325 13483 11359
rect 13517 11325 13551 11359
rect 13585 11325 13619 11359
rect 13653 11325 13687 11359
rect 13721 11325 13755 11359
rect 13789 11325 13823 11359
rect 13857 11325 13891 11359
rect 13925 11325 13959 11359
rect 13993 11325 14027 11359
rect 14061 11325 14095 11359
rect 14129 11325 14163 11359
rect 14197 11325 14231 11359
rect 14265 11325 14299 11359
rect 14333 11325 14367 11359
rect 14401 11325 14435 11359
rect 14469 11325 14503 11359
rect 14537 11325 14571 11359
rect 14605 11325 14639 11359
rect 14673 11325 14707 11359
rect 14741 11325 14775 11359
rect 14809 11325 14843 11359
rect 14877 11325 14911 11359
rect 14945 11325 14979 11359
rect 15013 11325 15047 11359
rect 15081 11325 15115 11359
rect 15149 11325 15183 11359
rect 15217 11325 15251 11359
rect 15285 11325 15319 11359
rect 15353 11325 15387 11359
rect 15421 11325 15455 11359
rect 15489 11325 15523 11359
rect 15557 11325 15591 11359
rect 15625 11325 15659 11359
rect 15693 11325 15727 11359
rect 15761 11325 15795 11359
rect 15829 11325 15884 11359
rect 13224 11289 15884 11325
rect 13224 11265 13279 11289
rect 13313 11265 13347 11289
rect 13381 11265 13415 11289
rect 4421 11228 6239 11263
rect 13118 11231 13157 11265
rect 13191 11231 13230 11265
rect 13264 11255 13279 11265
rect 13337 11255 13347 11265
rect 13410 11255 13415 11265
rect 13449 11265 13483 11289
rect 13264 11231 13303 11255
rect 13337 11231 13376 11255
rect 13410 11231 13449 11255
rect 13517 11265 13551 11289
rect 13585 11265 13619 11289
rect 13653 11265 13687 11289
rect 13721 11265 13755 11289
rect 13789 11265 13823 11289
rect 13857 11265 13891 11289
rect 13517 11255 13522 11265
rect 13585 11255 13595 11265
rect 13653 11255 13668 11265
rect 13721 11255 13741 11265
rect 13789 11255 13814 11265
rect 13857 11255 13887 11265
rect 13925 11255 13959 11289
rect 13993 11265 14027 11289
rect 14061 11265 14095 11289
rect 14129 11265 14163 11289
rect 14197 11265 14231 11289
rect 14265 11265 14299 11289
rect 14333 11265 14367 11289
rect 14401 11265 14435 11289
rect 13994 11255 14027 11265
rect 14067 11255 14095 11265
rect 14140 11255 14163 11265
rect 14213 11255 14231 11265
rect 14286 11255 14299 11265
rect 14359 11255 14367 11265
rect 14432 11255 14435 11265
rect 14469 11265 14503 11289
rect 14537 11265 14571 11289
rect 14605 11265 14639 11289
rect 14673 11265 14707 11289
rect 14741 11265 14775 11289
rect 14809 11265 14843 11289
rect 14877 11265 14911 11289
rect 14469 11255 14471 11265
rect 14537 11255 14544 11265
rect 14605 11255 14617 11265
rect 14673 11255 14690 11265
rect 14741 11255 14763 11265
rect 14809 11255 14836 11265
rect 14877 11255 14909 11265
rect 14945 11255 14979 11289
rect 15013 11265 15047 11289
rect 15081 11265 15115 11289
rect 15149 11265 15183 11289
rect 15217 11265 15251 11289
rect 15285 11265 15319 11289
rect 15353 11265 15387 11289
rect 15421 11265 15455 11289
rect 15016 11255 15047 11265
rect 15089 11255 15115 11265
rect 15162 11255 15183 11265
rect 15235 11255 15251 11265
rect 15307 11255 15319 11265
rect 15379 11255 15387 11265
rect 15451 11255 15455 11265
rect 15489 11265 15523 11289
rect 13483 11231 13522 11255
rect 13556 11231 13595 11255
rect 13629 11231 13668 11255
rect 13702 11231 13741 11255
rect 13775 11231 13814 11255
rect 13848 11231 13887 11255
rect 13921 11231 13960 11255
rect 13994 11231 14033 11255
rect 14067 11231 14106 11255
rect 14140 11231 14179 11255
rect 14213 11231 14252 11255
rect 14286 11231 14325 11255
rect 14359 11231 14398 11255
rect 14432 11231 14471 11255
rect 14505 11231 14544 11255
rect 14578 11231 14617 11255
rect 14651 11231 14690 11255
rect 14724 11231 14763 11255
rect 14797 11231 14836 11255
rect 14870 11231 14909 11255
rect 14943 11231 14982 11255
rect 15016 11231 15055 11255
rect 15089 11231 15128 11255
rect 15162 11231 15201 11255
rect 15235 11231 15273 11255
rect 15307 11231 15345 11255
rect 15379 11231 15417 11255
rect 15451 11231 15489 11255
rect 15557 11265 15591 11289
rect 15625 11265 15659 11289
rect 15693 11265 15727 11289
rect 15761 11265 15795 11289
rect 15829 11265 15884 11289
rect 15557 11255 15561 11265
rect 15625 11255 15633 11265
rect 15693 11255 15705 11265
rect 15761 11255 15777 11265
rect 15829 11255 15849 11265
rect 15523 11231 15561 11255
rect 15595 11231 15633 11255
rect 15667 11231 15705 11255
rect 15739 11231 15777 11255
rect 15811 11231 15849 11255
rect 15883 11231 15921 11265
rect 4421 11194 4429 11228
rect 4463 11194 4497 11228
rect 4531 11194 4565 11228
rect 4599 11194 4633 11228
rect 4667 11194 4701 11228
rect 4735 11194 4769 11228
rect 4803 11194 4837 11228
rect 4871 11194 4905 11228
rect 4939 11194 4973 11228
rect 5007 11194 5041 11228
rect 5075 11194 5109 11228
rect 5143 11194 5177 11228
rect 5211 11194 5245 11228
rect 5279 11194 5313 11228
rect 5347 11194 5381 11228
rect 5415 11194 5449 11228
rect 5483 11194 5517 11228
rect 5551 11194 5585 11228
rect 5619 11194 5653 11228
rect 5687 11194 5721 11228
rect 5755 11194 5789 11228
rect 5823 11194 5857 11228
rect 5891 11194 5925 11228
rect 5959 11194 5993 11228
rect 6027 11194 6061 11228
rect 6095 11194 6129 11228
rect 6163 11194 6197 11228
rect 6231 11194 6239 11228
rect 4421 11159 6239 11194
rect 4421 11125 4429 11159
rect 4463 11125 4497 11159
rect 4531 11125 4565 11159
rect 4599 11125 4633 11159
rect 4667 11125 4701 11159
rect 4735 11125 4769 11159
rect 4803 11125 4837 11159
rect 4871 11125 4905 11159
rect 4939 11125 4973 11159
rect 5007 11125 5041 11159
rect 5075 11125 5109 11159
rect 5143 11125 5177 11159
rect 5211 11125 5245 11159
rect 5279 11125 5313 11159
rect 5347 11125 5381 11159
rect 5415 11125 5449 11159
rect 5483 11125 5517 11159
rect 5551 11125 5585 11159
rect 5619 11125 5653 11159
rect 5687 11125 5721 11159
rect 5755 11125 5789 11159
rect 5823 11125 5857 11159
rect 5891 11125 5925 11159
rect 5959 11125 5993 11159
rect 6027 11125 6061 11159
rect 6095 11125 6129 11159
rect 6163 11125 6197 11159
rect 6231 11125 6239 11159
rect 4421 11090 6239 11125
rect 4421 11056 4429 11090
rect 4463 11056 4497 11090
rect 4531 11056 4565 11090
rect 4599 11056 4633 11090
rect 4667 11056 4701 11090
rect 4735 11056 4769 11090
rect 4803 11056 4837 11090
rect 4871 11056 4905 11090
rect 4939 11056 4973 11090
rect 5007 11056 5041 11090
rect 5075 11056 5109 11090
rect 5143 11056 5177 11090
rect 5211 11056 5245 11090
rect 5279 11056 5313 11090
rect 5347 11056 5381 11090
rect 5415 11056 5449 11090
rect 5483 11056 5517 11090
rect 5551 11056 5585 11090
rect 5619 11056 5653 11090
rect 5687 11056 5721 11090
rect 5755 11056 5789 11090
rect 5823 11056 5857 11090
rect 5891 11056 5925 11090
rect 5959 11056 5993 11090
rect 6027 11056 6061 11090
rect 6095 11056 6129 11090
rect 6163 11056 6197 11090
rect 6231 11056 6239 11090
rect 4421 11021 6239 11056
rect 4421 10987 4429 11021
rect 4463 10987 4497 11021
rect 4531 10987 4565 11021
rect 4599 10987 4633 11021
rect 4667 10987 4701 11021
rect 4735 10987 4769 11021
rect 4803 10987 4837 11021
rect 4871 10987 4905 11021
rect 4939 10987 4973 11021
rect 5007 10987 5041 11021
rect 5075 10987 5109 11021
rect 5143 10987 5177 11021
rect 5211 10987 5245 11021
rect 5279 10987 5313 11021
rect 5347 10987 5381 11021
rect 5415 10987 5449 11021
rect 5483 10987 5517 11021
rect 5551 10987 5585 11021
rect 5619 10987 5653 11021
rect 5687 10987 5721 11021
rect 5755 10987 5789 11021
rect 5823 10987 5857 11021
rect 5891 10987 5925 11021
rect 5959 10987 5993 11021
rect 6027 10987 6061 11021
rect 6095 10987 6129 11021
rect 6163 10987 6197 11021
rect 6231 10987 6239 11021
rect 4421 10952 6239 10987
rect 4421 10918 4429 10952
rect 4463 10937 4497 10952
rect 4531 10937 4565 10952
rect 4599 10937 4633 10952
rect 4667 10937 4701 10952
rect 4735 10937 4769 10952
rect 4467 10918 4497 10937
rect 4541 10918 4565 10937
rect 4615 10918 4633 10937
rect 4689 10918 4701 10937
rect 4763 10918 4769 10937
rect 4803 10937 4837 10952
rect 4421 10903 4433 10918
rect 4467 10903 4507 10918
rect 4541 10903 4581 10918
rect 4615 10903 4655 10918
rect 4689 10903 4729 10918
rect 4763 10903 4803 10918
rect 4871 10937 4905 10952
rect 4939 10937 4973 10952
rect 5007 10937 5041 10952
rect 5075 10937 5109 10952
rect 5143 10937 5177 10952
rect 5211 10937 5245 10952
rect 4871 10918 4876 10937
rect 4939 10918 4949 10937
rect 5007 10918 5022 10937
rect 5075 10918 5095 10937
rect 5143 10918 5168 10937
rect 5211 10918 5241 10937
rect 5279 10918 5313 10952
rect 5347 10937 5381 10952
rect 5415 10937 5449 10952
rect 5483 10937 5517 10952
rect 5551 10937 5585 10952
rect 5619 10937 5653 10952
rect 5687 10937 5721 10952
rect 5755 10937 5789 10952
rect 5348 10918 5381 10937
rect 5421 10918 5449 10937
rect 5494 10918 5517 10937
rect 5567 10918 5585 10937
rect 5640 10918 5653 10937
rect 5713 10918 5721 10937
rect 5786 10918 5789 10937
rect 5823 10937 5857 10952
rect 5891 10937 5925 10952
rect 5959 10937 5993 10952
rect 6027 10937 6061 10952
rect 6095 10937 6129 10952
rect 6163 10937 6197 10952
rect 5823 10918 5825 10937
rect 5891 10918 5898 10937
rect 5959 10918 5971 10937
rect 6027 10918 6044 10937
rect 6095 10918 6117 10937
rect 6163 10918 6190 10937
rect 6231 10918 6239 10952
rect 4837 10903 4876 10918
rect 4910 10903 4949 10918
rect 4983 10903 5022 10918
rect 5056 10903 5095 10918
rect 5129 10903 5168 10918
rect 5202 10903 5241 10918
rect 5275 10903 5314 10918
rect 5348 10903 5387 10918
rect 5421 10903 5460 10918
rect 5494 10903 5533 10918
rect 5567 10903 5606 10918
rect 5640 10903 5679 10918
rect 5713 10903 5752 10918
rect 5786 10903 5825 10918
rect 5859 10903 5898 10918
rect 5932 10903 5971 10918
rect 6005 10903 6044 10918
rect 6078 10903 6117 10918
rect 6151 10903 6190 10918
rect 6224 10903 6239 10918
rect 4421 10883 6239 10903
rect 4421 10849 4429 10883
rect 4463 10861 4497 10883
rect 4531 10861 4565 10883
rect 4599 10861 4633 10883
rect 4667 10861 4701 10883
rect 4735 10861 4769 10883
rect 4467 10849 4497 10861
rect 4541 10849 4565 10861
rect 4615 10849 4633 10861
rect 4689 10849 4701 10861
rect 4763 10849 4769 10861
rect 4803 10861 4837 10883
rect 4421 10827 4433 10849
rect 4467 10827 4507 10849
rect 4541 10827 4581 10849
rect 4615 10827 4655 10849
rect 4689 10827 4729 10849
rect 4763 10827 4803 10849
rect 4871 10861 4905 10883
rect 4939 10861 4973 10883
rect 5007 10861 5041 10883
rect 5075 10861 5109 10883
rect 5143 10861 5177 10883
rect 5211 10861 5245 10883
rect 4871 10849 4876 10861
rect 4939 10849 4949 10861
rect 5007 10849 5022 10861
rect 5075 10849 5095 10861
rect 5143 10849 5168 10861
rect 5211 10849 5241 10861
rect 5279 10849 5313 10883
rect 5347 10861 5381 10883
rect 5415 10861 5449 10883
rect 5483 10861 5517 10883
rect 5551 10861 5585 10883
rect 5619 10861 5653 10883
rect 5687 10861 5721 10883
rect 5755 10861 5789 10883
rect 5348 10849 5381 10861
rect 5421 10849 5449 10861
rect 5494 10849 5517 10861
rect 5567 10849 5585 10861
rect 5640 10849 5653 10861
rect 5713 10849 5721 10861
rect 5786 10849 5789 10861
rect 5823 10861 5857 10883
rect 5891 10861 5925 10883
rect 5959 10861 5993 10883
rect 6027 10861 6061 10883
rect 6095 10861 6129 10883
rect 6163 10861 6197 10883
rect 5823 10849 5825 10861
rect 5891 10849 5898 10861
rect 5959 10849 5971 10861
rect 6027 10849 6044 10861
rect 6095 10849 6117 10861
rect 6163 10849 6190 10861
rect 6231 10849 6239 10883
rect 13224 11219 15884 11231
rect 13224 11185 13279 11219
rect 13313 11185 13347 11219
rect 13381 11185 13415 11219
rect 13449 11185 13483 11219
rect 13517 11185 13551 11219
rect 13585 11185 13619 11219
rect 13653 11185 13687 11219
rect 13721 11185 13755 11219
rect 13789 11185 13823 11219
rect 13857 11185 13891 11219
rect 13925 11185 13959 11219
rect 13993 11185 14027 11219
rect 14061 11185 14095 11219
rect 14129 11185 14163 11219
rect 14197 11185 14231 11219
rect 14265 11185 14299 11219
rect 14333 11185 14367 11219
rect 14401 11185 14435 11219
rect 14469 11185 14503 11219
rect 14537 11185 14571 11219
rect 14605 11185 14639 11219
rect 14673 11185 14707 11219
rect 14741 11185 14775 11219
rect 14809 11185 14843 11219
rect 14877 11185 14911 11219
rect 14945 11185 14979 11219
rect 15013 11185 15047 11219
rect 15081 11185 15115 11219
rect 15149 11185 15183 11219
rect 15217 11185 15251 11219
rect 15285 11185 15319 11219
rect 15353 11185 15387 11219
rect 15421 11185 15455 11219
rect 15489 11185 15523 11219
rect 15557 11185 15591 11219
rect 15625 11185 15659 11219
rect 15693 11185 15727 11219
rect 15761 11185 15795 11219
rect 15829 11185 15884 11219
rect 13224 11149 15884 11185
rect 13224 11115 13279 11149
rect 13313 11115 13347 11149
rect 13381 11115 13415 11149
rect 13449 11115 13483 11149
rect 13517 11115 13551 11149
rect 13585 11115 13619 11149
rect 13653 11115 13687 11149
rect 13721 11115 13755 11149
rect 13789 11115 13823 11149
rect 13857 11115 13891 11149
rect 13925 11115 13959 11149
rect 13993 11115 14027 11149
rect 14061 11115 14095 11149
rect 14129 11115 14163 11149
rect 14197 11115 14231 11149
rect 14265 11115 14299 11149
rect 14333 11115 14367 11149
rect 14401 11115 14435 11149
rect 14469 11115 14503 11149
rect 14537 11115 14571 11149
rect 14605 11115 14639 11149
rect 14673 11115 14707 11149
rect 14741 11115 14775 11149
rect 14809 11115 14843 11149
rect 14877 11115 14911 11149
rect 14945 11115 14979 11149
rect 15013 11115 15047 11149
rect 15081 11115 15115 11149
rect 15149 11115 15183 11149
rect 15217 11115 15251 11149
rect 15285 11115 15319 11149
rect 15353 11115 15387 11149
rect 15421 11115 15455 11149
rect 15489 11115 15523 11149
rect 15557 11115 15591 11149
rect 15625 11115 15659 11149
rect 15693 11115 15727 11149
rect 15761 11115 15795 11149
rect 15829 11115 15884 11149
rect 13224 11079 15884 11115
rect 13224 11045 13279 11079
rect 13313 11045 13347 11079
rect 13381 11045 13415 11079
rect 13449 11045 13483 11079
rect 13517 11045 13551 11079
rect 13585 11045 13619 11079
rect 13653 11045 13687 11079
rect 13721 11045 13755 11079
rect 13789 11045 13823 11079
rect 13857 11045 13891 11079
rect 13925 11045 13959 11079
rect 13993 11045 14027 11079
rect 14061 11045 14095 11079
rect 14129 11045 14163 11079
rect 14197 11045 14231 11079
rect 14265 11045 14299 11079
rect 14333 11045 14367 11079
rect 14401 11045 14435 11079
rect 14469 11045 14503 11079
rect 14537 11045 14571 11079
rect 14605 11045 14639 11079
rect 14673 11045 14707 11079
rect 14741 11045 14775 11079
rect 14809 11045 14843 11079
rect 14877 11045 14911 11079
rect 14945 11045 14979 11079
rect 15013 11045 15047 11079
rect 15081 11045 15115 11079
rect 15149 11045 15183 11079
rect 15217 11045 15251 11079
rect 15285 11045 15319 11079
rect 15353 11045 15387 11079
rect 15421 11045 15455 11079
rect 15489 11045 15523 11079
rect 15557 11045 15591 11079
rect 15625 11045 15659 11079
rect 15693 11045 15727 11079
rect 15761 11045 15795 11079
rect 15829 11045 15884 11079
rect 13224 11009 15884 11045
rect 13224 10975 13279 11009
rect 13313 10975 13347 11009
rect 13381 10975 13415 11009
rect 13449 10975 13483 11009
rect 13517 10975 13551 11009
rect 13585 10975 13619 11009
rect 13653 10975 13687 11009
rect 13721 10975 13755 11009
rect 13789 10975 13823 11009
rect 13857 10975 13891 11009
rect 13925 10975 13959 11009
rect 13993 10975 14027 11009
rect 14061 10975 14095 11009
rect 14129 10975 14163 11009
rect 14197 10975 14231 11009
rect 14265 10975 14299 11009
rect 14333 10975 14367 11009
rect 14401 10975 14435 11009
rect 14469 10975 14503 11009
rect 14537 10975 14571 11009
rect 14605 10975 14639 11009
rect 14673 10975 14707 11009
rect 14741 10975 14775 11009
rect 14809 10975 14843 11009
rect 14877 10975 14911 11009
rect 14945 10975 14979 11009
rect 15013 10975 15047 11009
rect 15081 10975 15115 11009
rect 15149 10975 15183 11009
rect 15217 10975 15251 11009
rect 15285 10975 15319 11009
rect 15353 10975 15387 11009
rect 15421 10975 15455 11009
rect 15489 10975 15523 11009
rect 15557 10975 15591 11009
rect 15625 10975 15659 11009
rect 15693 10975 15727 11009
rect 15761 10975 15795 11009
rect 15829 10975 15884 11009
rect 13224 10939 15884 10975
rect 13224 10905 13279 10939
rect 13313 10905 13347 10939
rect 13381 10934 13415 10939
rect 13449 10934 13483 10939
rect 13517 10934 13551 10939
rect 13398 10905 13415 10934
rect 13472 10905 13483 10934
rect 13546 10905 13551 10934
rect 13585 10934 13619 10939
rect 13224 10900 13364 10905
rect 13398 10900 13438 10905
rect 13472 10900 13512 10905
rect 13546 10900 13585 10905
rect 13653 10934 13687 10939
rect 13721 10934 13755 10939
rect 13789 10934 13823 10939
rect 13857 10934 13891 10939
rect 13925 10934 13959 10939
rect 13993 10934 14027 10939
rect 13653 10905 13658 10934
rect 13721 10905 13731 10934
rect 13789 10905 13804 10934
rect 13857 10905 13877 10934
rect 13925 10905 13950 10934
rect 13993 10905 14023 10934
rect 14061 10905 14095 10939
rect 14129 10934 14163 10939
rect 14197 10934 14231 10939
rect 14265 10934 14299 10939
rect 14333 10934 14367 10939
rect 14401 10934 14435 10939
rect 14469 10934 14503 10939
rect 14537 10934 14571 10939
rect 14130 10905 14163 10934
rect 14203 10905 14231 10934
rect 14276 10905 14299 10934
rect 14349 10905 14367 10934
rect 14422 10905 14435 10934
rect 14495 10905 14503 10934
rect 14568 10905 14571 10934
rect 14605 10934 14639 10939
rect 14673 10934 14707 10939
rect 14741 10934 14775 10939
rect 14809 10934 14843 10939
rect 14877 10934 14911 10939
rect 14945 10934 14979 10939
rect 15013 10934 15047 10939
rect 14605 10905 14607 10934
rect 14673 10905 14680 10934
rect 14741 10905 14753 10934
rect 14809 10905 14826 10934
rect 14877 10905 14899 10934
rect 14945 10905 14972 10934
rect 15013 10905 15045 10934
rect 15081 10905 15115 10939
rect 15149 10934 15183 10939
rect 15217 10934 15251 10939
rect 15285 10934 15319 10939
rect 15353 10934 15387 10939
rect 15421 10934 15455 10939
rect 15489 10934 15523 10939
rect 15557 10934 15591 10939
rect 15152 10905 15183 10934
rect 15225 10905 15251 10934
rect 15298 10905 15319 10934
rect 15371 10905 15387 10934
rect 15444 10905 15455 10934
rect 15517 10905 15523 10934
rect 15590 10905 15591 10934
rect 15625 10934 15659 10939
rect 15693 10934 15727 10939
rect 15761 10934 15795 10939
rect 15829 10934 15884 10939
rect 15625 10905 15629 10934
rect 15693 10905 15702 10934
rect 15761 10905 15775 10934
rect 15829 10905 15848 10934
rect 13619 10900 13658 10905
rect 13692 10900 13731 10905
rect 13765 10900 13804 10905
rect 13838 10900 13877 10905
rect 13911 10900 13950 10905
rect 13984 10900 14023 10905
rect 14057 10900 14096 10905
rect 14130 10900 14169 10905
rect 14203 10900 14242 10905
rect 14276 10900 14315 10905
rect 14349 10900 14388 10905
rect 14422 10900 14461 10905
rect 14495 10900 14534 10905
rect 14568 10900 14607 10905
rect 14641 10900 14680 10905
rect 14714 10900 14753 10905
rect 14787 10900 14826 10905
rect 14860 10900 14899 10905
rect 14933 10900 14972 10905
rect 15006 10900 15045 10905
rect 15079 10900 15118 10905
rect 15152 10900 15191 10905
rect 15225 10900 15264 10905
rect 15298 10900 15337 10905
rect 15371 10900 15410 10905
rect 15444 10900 15483 10905
rect 15517 10900 15556 10905
rect 15590 10900 15629 10905
rect 15663 10900 15702 10905
rect 15736 10900 15775 10905
rect 15809 10900 15848 10905
rect 15882 10900 15884 10934
rect 4837 10827 4876 10849
rect 4910 10827 4949 10849
rect 4983 10827 5022 10849
rect 5056 10827 5095 10849
rect 5129 10827 5168 10849
rect 5202 10827 5241 10849
rect 5275 10827 5314 10849
rect 5348 10827 5387 10849
rect 5421 10827 5460 10849
rect 5494 10827 5533 10849
rect 5567 10827 5606 10849
rect 5640 10827 5679 10849
rect 5713 10827 5752 10849
rect 5786 10827 5825 10849
rect 5859 10827 5898 10849
rect 5932 10827 5971 10849
rect 6005 10827 6044 10849
rect 6078 10827 6117 10849
rect 6151 10827 6190 10849
rect 6224 10827 6239 10849
rect 4421 10814 6239 10827
rect 4421 10780 4429 10814
rect 4463 10785 4497 10814
rect 4531 10785 4565 10814
rect 4599 10785 4633 10814
rect 4667 10785 4701 10814
rect 4735 10785 4769 10814
rect 4467 10780 4497 10785
rect 4541 10780 4565 10785
rect 4615 10780 4633 10785
rect 4689 10780 4701 10785
rect 4763 10780 4769 10785
rect 4803 10785 4837 10814
rect 4421 10751 4433 10780
rect 4467 10751 4507 10780
rect 4541 10751 4581 10780
rect 4615 10751 4655 10780
rect 4689 10751 4729 10780
rect 4763 10751 4803 10780
rect 4871 10785 4905 10814
rect 4939 10785 4973 10814
rect 5007 10785 5041 10814
rect 5075 10785 5109 10814
rect 5143 10785 5177 10814
rect 5211 10785 5245 10814
rect 4871 10780 4876 10785
rect 4939 10780 4949 10785
rect 5007 10780 5022 10785
rect 5075 10780 5095 10785
rect 5143 10780 5168 10785
rect 5211 10780 5241 10785
rect 5279 10780 5313 10814
rect 5347 10785 5381 10814
rect 5415 10785 5449 10814
rect 5483 10785 5517 10814
rect 5551 10785 5585 10814
rect 5619 10785 5653 10814
rect 5687 10785 5721 10814
rect 5755 10785 5789 10814
rect 5348 10780 5381 10785
rect 5421 10780 5449 10785
rect 5494 10780 5517 10785
rect 5567 10780 5585 10785
rect 5640 10780 5653 10785
rect 5713 10780 5721 10785
rect 5786 10780 5789 10785
rect 5823 10785 5857 10814
rect 5891 10785 5925 10814
rect 5959 10785 5993 10814
rect 6027 10785 6061 10814
rect 6095 10785 6129 10814
rect 6163 10785 6197 10814
rect 5823 10780 5825 10785
rect 5891 10780 5898 10785
rect 5959 10780 5971 10785
rect 6027 10780 6044 10785
rect 6095 10780 6117 10785
rect 6163 10780 6190 10785
rect 6231 10780 6239 10814
rect 4837 10751 4876 10780
rect 4910 10751 4949 10780
rect 4983 10751 5022 10780
rect 5056 10751 5095 10780
rect 5129 10751 5168 10780
rect 5202 10751 5241 10780
rect 5275 10751 5314 10780
rect 5348 10751 5387 10780
rect 5421 10751 5460 10780
rect 5494 10751 5533 10780
rect 5567 10751 5606 10780
rect 5640 10751 5679 10780
rect 5713 10751 5752 10780
rect 5786 10751 5825 10780
rect 5859 10751 5898 10780
rect 5932 10751 5971 10780
rect 6005 10751 6044 10780
rect 6078 10751 6117 10780
rect 6151 10751 6190 10780
rect 6224 10751 6239 10780
rect 4421 10745 6239 10751
rect 4421 10711 4429 10745
rect 4463 10711 4497 10745
rect 4531 10711 4565 10745
rect 4599 10711 4633 10745
rect 4667 10711 4701 10745
rect 4735 10711 4769 10745
rect 4803 10711 4837 10745
rect 4871 10711 4905 10745
rect 4939 10711 4973 10745
rect 5007 10711 5041 10745
rect 5075 10711 5109 10745
rect 5143 10711 5177 10745
rect 5211 10711 5245 10745
rect 5279 10711 5313 10745
rect 5347 10711 5381 10745
rect 5415 10711 5449 10745
rect 5483 10711 5517 10745
rect 5551 10711 5585 10745
rect 5619 10711 5653 10745
rect 5687 10711 5721 10745
rect 5755 10711 5789 10745
rect 5823 10711 5857 10745
rect 5891 10711 5925 10745
rect 5959 10711 5993 10745
rect 6027 10711 6061 10745
rect 6095 10711 6129 10745
rect 6163 10711 6197 10745
rect 6231 10711 6239 10745
rect 4421 10676 6239 10711
rect 12508 10684 12844 10877
rect 13224 10869 15884 10900
rect 13224 10835 13279 10869
rect 13313 10835 13347 10869
rect 13381 10860 13415 10869
rect 13449 10860 13483 10869
rect 13517 10860 13551 10869
rect 13398 10835 13415 10860
rect 13472 10835 13483 10860
rect 13546 10835 13551 10860
rect 13585 10860 13619 10869
rect 13224 10826 13364 10835
rect 13398 10826 13438 10835
rect 13472 10826 13512 10835
rect 13546 10826 13585 10835
rect 13653 10860 13687 10869
rect 13721 10860 13755 10869
rect 13789 10860 13823 10869
rect 13857 10860 13891 10869
rect 13925 10860 13959 10869
rect 13993 10860 14027 10869
rect 13653 10835 13658 10860
rect 13721 10835 13731 10860
rect 13789 10835 13804 10860
rect 13857 10835 13877 10860
rect 13925 10835 13950 10860
rect 13993 10835 14023 10860
rect 14061 10835 14095 10869
rect 14129 10860 14163 10869
rect 14197 10860 14231 10869
rect 14265 10860 14299 10869
rect 14333 10860 14367 10869
rect 14401 10860 14435 10869
rect 14469 10860 14503 10869
rect 14537 10860 14571 10869
rect 14130 10835 14163 10860
rect 14203 10835 14231 10860
rect 14276 10835 14299 10860
rect 14349 10835 14367 10860
rect 14422 10835 14435 10860
rect 14495 10835 14503 10860
rect 14568 10835 14571 10860
rect 14605 10860 14639 10869
rect 14673 10860 14707 10869
rect 14741 10860 14775 10869
rect 14809 10860 14843 10869
rect 14877 10860 14911 10869
rect 14945 10860 14979 10869
rect 15013 10860 15047 10869
rect 14605 10835 14607 10860
rect 14673 10835 14680 10860
rect 14741 10835 14753 10860
rect 14809 10835 14826 10860
rect 14877 10835 14899 10860
rect 14945 10835 14972 10860
rect 15013 10835 15045 10860
rect 15081 10835 15115 10869
rect 15149 10860 15183 10869
rect 15217 10860 15251 10869
rect 15285 10860 15319 10869
rect 15353 10860 15387 10869
rect 15421 10860 15455 10869
rect 15489 10860 15523 10869
rect 15557 10860 15591 10869
rect 15152 10835 15183 10860
rect 15225 10835 15251 10860
rect 15298 10835 15319 10860
rect 15371 10835 15387 10860
rect 15444 10835 15455 10860
rect 15517 10835 15523 10860
rect 15590 10835 15591 10860
rect 15625 10860 15659 10869
rect 15693 10860 15727 10869
rect 15761 10860 15795 10869
rect 15829 10860 15884 10869
rect 15625 10835 15629 10860
rect 15693 10835 15702 10860
rect 15761 10835 15775 10860
rect 15829 10835 15848 10860
rect 13619 10826 13658 10835
rect 13692 10826 13731 10835
rect 13765 10826 13804 10835
rect 13838 10826 13877 10835
rect 13911 10826 13950 10835
rect 13984 10826 14023 10835
rect 14057 10826 14096 10835
rect 14130 10826 14169 10835
rect 14203 10826 14242 10835
rect 14276 10826 14315 10835
rect 14349 10826 14388 10835
rect 14422 10826 14461 10835
rect 14495 10826 14534 10835
rect 14568 10826 14607 10835
rect 14641 10826 14680 10835
rect 14714 10826 14753 10835
rect 14787 10826 14826 10835
rect 14860 10826 14899 10835
rect 14933 10826 14972 10835
rect 15006 10826 15045 10835
rect 15079 10826 15118 10835
rect 15152 10826 15191 10835
rect 15225 10826 15264 10835
rect 15298 10826 15337 10835
rect 15371 10826 15410 10835
rect 15444 10826 15483 10835
rect 15517 10826 15556 10835
rect 15590 10826 15629 10835
rect 15663 10826 15702 10835
rect 15736 10826 15775 10835
rect 15809 10826 15848 10835
rect 15882 10826 15884 10860
rect 13224 10799 15884 10826
rect 13224 10765 13279 10799
rect 13313 10765 13347 10799
rect 13381 10786 13415 10799
rect 13449 10786 13483 10799
rect 13517 10786 13551 10799
rect 13398 10765 13415 10786
rect 13472 10765 13483 10786
rect 13546 10765 13551 10786
rect 13585 10786 13619 10799
rect 13224 10752 13364 10765
rect 13398 10752 13438 10765
rect 13472 10752 13512 10765
rect 13546 10752 13585 10765
rect 13653 10786 13687 10799
rect 13721 10786 13755 10799
rect 13789 10786 13823 10799
rect 13857 10786 13891 10799
rect 13925 10786 13959 10799
rect 13993 10786 14027 10799
rect 13653 10765 13658 10786
rect 13721 10765 13731 10786
rect 13789 10765 13804 10786
rect 13857 10765 13877 10786
rect 13925 10765 13950 10786
rect 13993 10765 14023 10786
rect 14061 10765 14095 10799
rect 14129 10786 14163 10799
rect 14197 10786 14231 10799
rect 14265 10786 14299 10799
rect 14333 10786 14367 10799
rect 14401 10786 14435 10799
rect 14469 10786 14503 10799
rect 14537 10786 14571 10799
rect 14130 10765 14163 10786
rect 14203 10765 14231 10786
rect 14276 10765 14299 10786
rect 14349 10765 14367 10786
rect 14422 10765 14435 10786
rect 14495 10765 14503 10786
rect 14568 10765 14571 10786
rect 14605 10786 14639 10799
rect 14673 10786 14707 10799
rect 14741 10786 14775 10799
rect 14809 10786 14843 10799
rect 14877 10786 14911 10799
rect 14945 10786 14979 10799
rect 15013 10786 15047 10799
rect 14605 10765 14607 10786
rect 14673 10765 14680 10786
rect 14741 10765 14753 10786
rect 14809 10765 14826 10786
rect 14877 10765 14899 10786
rect 14945 10765 14972 10786
rect 15013 10765 15045 10786
rect 15081 10765 15115 10799
rect 15149 10786 15183 10799
rect 15217 10786 15251 10799
rect 15285 10786 15319 10799
rect 15353 10786 15387 10799
rect 15421 10786 15455 10799
rect 15489 10786 15523 10799
rect 15557 10786 15591 10799
rect 15152 10765 15183 10786
rect 15225 10765 15251 10786
rect 15298 10765 15319 10786
rect 15371 10765 15387 10786
rect 15444 10765 15455 10786
rect 15517 10765 15523 10786
rect 15590 10765 15591 10786
rect 15625 10786 15659 10799
rect 15693 10786 15727 10799
rect 15761 10786 15795 10799
rect 15829 10786 15884 10799
rect 15625 10765 15629 10786
rect 15693 10765 15702 10786
rect 15761 10765 15775 10786
rect 15829 10765 15848 10786
rect 13619 10752 13658 10765
rect 13692 10752 13731 10765
rect 13765 10752 13804 10765
rect 13838 10752 13877 10765
rect 13911 10752 13950 10765
rect 13984 10752 14023 10765
rect 14057 10752 14096 10765
rect 14130 10752 14169 10765
rect 14203 10752 14242 10765
rect 14276 10752 14315 10765
rect 14349 10752 14388 10765
rect 14422 10752 14461 10765
rect 14495 10752 14534 10765
rect 14568 10752 14607 10765
rect 14641 10752 14680 10765
rect 14714 10752 14753 10765
rect 14787 10752 14826 10765
rect 14860 10752 14899 10765
rect 14933 10752 14972 10765
rect 15006 10752 15045 10765
rect 15079 10752 15118 10765
rect 15152 10752 15191 10765
rect 15225 10752 15264 10765
rect 15298 10752 15337 10765
rect 15371 10752 15410 10765
rect 15444 10752 15483 10765
rect 15517 10752 15556 10765
rect 15590 10752 15629 10765
rect 15663 10752 15702 10765
rect 15736 10752 15775 10765
rect 15809 10752 15848 10765
rect 15882 10752 15884 10786
rect 13224 10729 15884 10752
rect 13224 10695 13279 10729
rect 13313 10695 13347 10729
rect 13381 10695 13415 10729
rect 13449 10695 13483 10729
rect 13517 10695 13551 10729
rect 13585 10695 13619 10729
rect 13653 10695 13687 10729
rect 13721 10695 13755 10729
rect 13789 10695 13823 10729
rect 13857 10695 13891 10729
rect 13925 10695 13959 10729
rect 13993 10695 14027 10729
rect 14061 10695 14095 10729
rect 14129 10695 14163 10729
rect 14197 10695 14231 10729
rect 14265 10695 14299 10729
rect 14333 10695 14367 10729
rect 14401 10695 14435 10729
rect 14469 10695 14503 10729
rect 14537 10695 14571 10729
rect 14605 10695 14639 10729
rect 14673 10695 14707 10729
rect 14741 10695 14775 10729
rect 14809 10695 14843 10729
rect 14877 10695 14911 10729
rect 14945 10695 14979 10729
rect 15013 10695 15047 10729
rect 15081 10695 15115 10729
rect 15149 10695 15183 10729
rect 15217 10695 15251 10729
rect 15285 10695 15319 10729
rect 15353 10695 15387 10729
rect 15421 10695 15455 10729
rect 15489 10695 15523 10729
rect 15557 10695 15591 10729
rect 15625 10695 15659 10729
rect 15693 10695 15727 10729
rect 15761 10695 15795 10729
rect 15829 10695 15884 10729
rect 4421 10642 4429 10676
rect 4463 10642 4497 10676
rect 4531 10642 4565 10676
rect 4599 10642 4633 10676
rect 4667 10642 4701 10676
rect 4735 10642 4769 10676
rect 4803 10642 4837 10676
rect 4871 10642 4905 10676
rect 4939 10642 4973 10676
rect 5007 10642 5041 10676
rect 5075 10642 5109 10676
rect 5143 10642 5177 10676
rect 5211 10642 5245 10676
rect 5279 10642 5313 10676
rect 5347 10642 5381 10676
rect 5415 10642 5449 10676
rect 5483 10642 5517 10676
rect 5551 10642 5585 10676
rect 5619 10642 5653 10676
rect 5687 10642 5721 10676
rect 5755 10642 5789 10676
rect 5823 10642 5857 10676
rect 5891 10642 5925 10676
rect 5959 10642 5993 10676
rect 6027 10642 6061 10676
rect 6095 10642 6129 10676
rect 6163 10642 6197 10676
rect 6231 10642 6239 10676
rect 4421 10607 6239 10642
rect 4421 10573 4429 10607
rect 4463 10573 4497 10607
rect 4531 10573 4565 10607
rect 4599 10573 4633 10607
rect 4667 10573 4701 10607
rect 4735 10573 4769 10607
rect 4803 10573 4837 10607
rect 4871 10573 4905 10607
rect 4939 10573 4973 10607
rect 5007 10573 5041 10607
rect 5075 10573 5109 10607
rect 5143 10573 5177 10607
rect 5211 10573 5245 10607
rect 5279 10573 5313 10607
rect 5347 10573 5381 10607
rect 5415 10573 5449 10607
rect 5483 10573 5517 10607
rect 5551 10573 5585 10607
rect 5619 10573 5653 10607
rect 5687 10573 5721 10607
rect 5755 10573 5789 10607
rect 5823 10573 5857 10607
rect 5891 10573 5925 10607
rect 5959 10573 5993 10607
rect 6027 10573 6061 10607
rect 6095 10573 6129 10607
rect 6163 10573 6197 10607
rect 6231 10573 6239 10607
rect 4421 10538 6239 10573
rect 13224 10659 15884 10695
rect 13224 10625 13279 10659
rect 13313 10625 13347 10659
rect 13381 10625 13415 10659
rect 13449 10625 13483 10659
rect 13517 10625 13551 10659
rect 13585 10625 13619 10659
rect 13653 10625 13687 10659
rect 13721 10625 13755 10659
rect 13789 10625 13823 10659
rect 13857 10625 13891 10659
rect 13925 10625 13959 10659
rect 13993 10625 14027 10659
rect 14061 10625 14095 10659
rect 14129 10625 14163 10659
rect 14197 10625 14231 10659
rect 14265 10625 14299 10659
rect 14333 10625 14367 10659
rect 14401 10625 14435 10659
rect 14469 10625 14503 10659
rect 14537 10625 14571 10659
rect 14605 10625 14639 10659
rect 14673 10625 14707 10659
rect 14741 10625 14775 10659
rect 14809 10625 14843 10659
rect 14877 10625 14911 10659
rect 14945 10625 14979 10659
rect 15013 10625 15047 10659
rect 15081 10625 15115 10659
rect 15149 10625 15183 10659
rect 15217 10625 15251 10659
rect 15285 10625 15319 10659
rect 15353 10625 15387 10659
rect 15421 10625 15455 10659
rect 15489 10625 15523 10659
rect 15557 10625 15591 10659
rect 15625 10625 15659 10659
rect 15693 10625 15727 10659
rect 15761 10625 15795 10659
rect 15829 10625 15884 10659
rect 13224 10589 15884 10625
rect 13224 10555 13279 10589
rect 13313 10555 13347 10589
rect 13381 10555 13415 10589
rect 13449 10555 13483 10589
rect 13517 10555 13551 10589
rect 13585 10555 13619 10589
rect 13653 10555 13687 10589
rect 13721 10555 13755 10589
rect 13789 10555 13823 10589
rect 13857 10555 13891 10589
rect 13925 10555 13959 10589
rect 13993 10555 14027 10589
rect 14061 10555 14095 10589
rect 14129 10555 14163 10589
rect 14197 10555 14231 10589
rect 14265 10555 14299 10589
rect 14333 10555 14367 10589
rect 14401 10555 14435 10589
rect 14469 10555 14503 10589
rect 14537 10555 14571 10589
rect 14605 10555 14639 10589
rect 14673 10555 14707 10589
rect 14741 10555 14775 10589
rect 14809 10555 14843 10589
rect 14877 10555 14911 10589
rect 14945 10555 14979 10589
rect 15013 10555 15047 10589
rect 15081 10555 15115 10589
rect 15149 10555 15183 10589
rect 15217 10555 15251 10589
rect 15285 10555 15319 10589
rect 15353 10555 15387 10589
rect 15421 10555 15455 10589
rect 15489 10555 15523 10589
rect 15557 10555 15591 10589
rect 15625 10555 15659 10589
rect 15693 10555 15727 10589
rect 15761 10555 15795 10589
rect 15829 10555 15884 10589
rect 13224 10542 15884 10555
rect 4421 10504 4429 10538
rect 4463 10504 4497 10538
rect 4531 10504 4565 10538
rect 4599 10504 4633 10538
rect 4667 10504 4701 10538
rect 4735 10504 4769 10538
rect 4803 10504 4837 10538
rect 4871 10504 4905 10538
rect 4939 10504 4973 10538
rect 5007 10504 5041 10538
rect 5075 10504 5109 10538
rect 5143 10504 5177 10538
rect 5211 10504 5245 10538
rect 5279 10504 5313 10538
rect 5347 10504 5381 10538
rect 5415 10504 5449 10538
rect 5483 10504 5517 10538
rect 5551 10504 5585 10538
rect 5619 10504 5653 10538
rect 5687 10504 5721 10538
rect 5755 10504 5789 10538
rect 5823 10504 5857 10538
rect 5891 10504 5925 10538
rect 5959 10504 5993 10538
rect 6027 10504 6061 10538
rect 6095 10504 6129 10538
rect 6163 10504 6197 10538
rect 6231 10504 6239 10538
rect 13150 10508 13190 10542
rect 13224 10508 13264 10542
rect 13298 10519 13338 10542
rect 13372 10519 13412 10542
rect 13446 10519 13486 10542
rect 13520 10519 13560 10542
rect 13594 10519 13634 10542
rect 13668 10519 13708 10542
rect 13742 10519 13782 10542
rect 13816 10519 13856 10542
rect 13890 10519 13930 10542
rect 13964 10519 14004 10542
rect 14038 10519 14078 10542
rect 14112 10519 14152 10542
rect 14186 10519 14226 10542
rect 14260 10519 14300 10542
rect 14334 10519 14374 10542
rect 14408 10519 14448 10542
rect 14482 10519 14522 10542
rect 14556 10519 14596 10542
rect 14630 10519 14670 10542
rect 14704 10519 14744 10542
rect 14778 10519 14818 10542
rect 14852 10519 14892 10542
rect 14926 10519 14966 10542
rect 15000 10519 15040 10542
rect 15074 10519 15114 10542
rect 15148 10519 15188 10542
rect 15222 10519 15261 10542
rect 15295 10519 15334 10542
rect 15368 10519 15407 10542
rect 15441 10519 15480 10542
rect 15514 10519 15553 10542
rect 15587 10519 15626 10542
rect 15660 10519 15699 10542
rect 15733 10519 15884 10542
rect 13313 10508 13338 10519
rect 13381 10508 13412 10519
rect 4421 10469 6239 10504
rect 4421 10435 4429 10469
rect 4463 10435 4497 10469
rect 4531 10435 4565 10469
rect 4599 10435 4633 10469
rect 4667 10435 4701 10469
rect 4735 10435 4769 10469
rect 4803 10435 4837 10469
rect 4871 10435 4905 10469
rect 4939 10435 4973 10469
rect 5007 10435 5041 10469
rect 5075 10435 5109 10469
rect 5143 10435 5177 10469
rect 5211 10435 5245 10469
rect 5279 10435 5313 10469
rect 5347 10435 5381 10469
rect 5415 10435 5449 10469
rect 5483 10435 5517 10469
rect 5551 10435 5585 10469
rect 5619 10435 5653 10469
rect 5687 10435 5721 10469
rect 5755 10435 5789 10469
rect 5823 10435 5857 10469
rect 5891 10435 5925 10469
rect 5959 10435 5993 10469
rect 6027 10435 6061 10469
rect 6095 10435 6129 10469
rect 6163 10435 6197 10469
rect 6231 10435 6239 10469
rect 4421 10400 6239 10435
rect 4421 10366 4429 10400
rect 4463 10366 4497 10400
rect 4531 10366 4565 10400
rect 4599 10366 4633 10400
rect 4667 10366 4701 10400
rect 4735 10366 4769 10400
rect 4803 10366 4837 10400
rect 4871 10366 4905 10400
rect 4939 10366 4973 10400
rect 5007 10366 5041 10400
rect 5075 10366 5109 10400
rect 5143 10366 5177 10400
rect 5211 10366 5245 10400
rect 5279 10366 5313 10400
rect 5347 10366 5381 10400
rect 5415 10366 5449 10400
rect 5483 10366 5517 10400
rect 5551 10366 5585 10400
rect 5619 10366 5653 10400
rect 5687 10366 5721 10400
rect 5755 10366 5789 10400
rect 5823 10366 5857 10400
rect 5891 10366 5925 10400
rect 5959 10366 5993 10400
rect 6027 10366 6061 10400
rect 6095 10366 6129 10400
rect 6163 10366 6197 10400
rect 6231 10366 6239 10400
rect 4421 10331 6239 10366
rect 4421 10297 4429 10331
rect 4463 10297 4497 10331
rect 4531 10297 4565 10331
rect 4599 10297 4633 10331
rect 4667 10297 4701 10331
rect 4735 10297 4769 10331
rect 4803 10297 4837 10331
rect 4871 10297 4905 10331
rect 4939 10297 4973 10331
rect 5007 10297 5041 10331
rect 5075 10297 5109 10331
rect 5143 10297 5177 10331
rect 5211 10297 5245 10331
rect 5279 10297 5313 10331
rect 5347 10297 5381 10331
rect 5415 10297 5449 10331
rect 5483 10297 5517 10331
rect 5551 10297 5585 10331
rect 5619 10297 5653 10331
rect 5687 10297 5721 10331
rect 5755 10297 5789 10331
rect 5823 10297 5857 10331
rect 5891 10297 5925 10331
rect 5959 10297 5993 10331
rect 6027 10297 6061 10331
rect 6095 10297 6129 10331
rect 6163 10297 6197 10331
rect 6231 10297 6239 10331
rect 13224 10485 13279 10508
rect 13313 10485 13347 10508
rect 13381 10485 13415 10508
rect 13449 10485 13483 10519
rect 13520 10508 13551 10519
rect 13594 10508 13619 10519
rect 13668 10508 13687 10519
rect 13742 10508 13755 10519
rect 13816 10508 13823 10519
rect 13890 10508 13891 10519
rect 13517 10485 13551 10508
rect 13585 10485 13619 10508
rect 13653 10485 13687 10508
rect 13721 10485 13755 10508
rect 13789 10485 13823 10508
rect 13857 10485 13891 10508
rect 13925 10508 13930 10519
rect 13993 10508 14004 10519
rect 14061 10508 14078 10519
rect 14129 10508 14152 10519
rect 14197 10508 14226 10519
rect 13925 10485 13959 10508
rect 13993 10485 14027 10508
rect 14061 10485 14095 10508
rect 14129 10485 14163 10508
rect 14197 10485 14231 10508
rect 14265 10485 14299 10519
rect 14334 10508 14367 10519
rect 14408 10508 14435 10519
rect 14482 10508 14503 10519
rect 14556 10508 14571 10519
rect 14630 10508 14639 10519
rect 14704 10508 14707 10519
rect 14333 10485 14367 10508
rect 14401 10485 14435 10508
rect 14469 10485 14503 10508
rect 14537 10485 14571 10508
rect 14605 10485 14639 10508
rect 14673 10485 14707 10508
rect 14741 10508 14744 10519
rect 14809 10508 14818 10519
rect 14877 10508 14892 10519
rect 14945 10508 14966 10519
rect 15013 10508 15040 10519
rect 15081 10508 15114 10519
rect 14741 10485 14775 10508
rect 14809 10485 14843 10508
rect 14877 10485 14911 10508
rect 14945 10485 14979 10508
rect 15013 10485 15047 10508
rect 15081 10485 15115 10508
rect 15149 10485 15183 10519
rect 15222 10508 15251 10519
rect 15295 10508 15319 10519
rect 15368 10508 15387 10519
rect 15441 10508 15455 10519
rect 15514 10508 15523 10519
rect 15587 10508 15591 10519
rect 15217 10485 15251 10508
rect 15285 10485 15319 10508
rect 15353 10485 15387 10508
rect 15421 10485 15455 10508
rect 15489 10485 15523 10508
rect 15557 10485 15591 10508
rect 15625 10508 15626 10519
rect 15693 10508 15699 10519
rect 15625 10485 15659 10508
rect 15693 10485 15727 10508
rect 15761 10485 15795 10519
rect 15829 10485 15884 10519
rect 13224 10449 15884 10485
rect 13224 10415 13279 10449
rect 13313 10415 13347 10449
rect 13381 10415 13415 10449
rect 13449 10415 13483 10449
rect 13517 10415 13551 10449
rect 13585 10415 13619 10449
rect 13653 10415 13687 10449
rect 13721 10415 13755 10449
rect 13789 10415 13823 10449
rect 13857 10415 13891 10449
rect 13925 10415 13959 10449
rect 13993 10415 14027 10449
rect 14061 10415 14095 10449
rect 14129 10415 14163 10449
rect 14197 10415 14231 10449
rect 14265 10415 14299 10449
rect 14333 10415 14367 10449
rect 14401 10415 14435 10449
rect 14469 10415 14503 10449
rect 14537 10415 14571 10449
rect 14605 10415 14639 10449
rect 14673 10415 14707 10449
rect 14741 10415 14775 10449
rect 14809 10415 14843 10449
rect 14877 10415 14911 10449
rect 14945 10415 14979 10449
rect 15013 10415 15047 10449
rect 15081 10415 15115 10449
rect 15149 10415 15183 10449
rect 15217 10415 15251 10449
rect 15285 10415 15319 10449
rect 15353 10415 15387 10449
rect 15421 10415 15455 10449
rect 15489 10415 15523 10449
rect 15557 10415 15591 10449
rect 15625 10415 15659 10449
rect 15693 10415 15727 10449
rect 15761 10415 15795 10449
rect 15829 10415 15884 10449
rect 13224 10379 15884 10415
rect 13224 10345 13279 10379
rect 13313 10345 13347 10379
rect 13381 10345 13415 10379
rect 13449 10345 13483 10379
rect 13517 10345 13551 10379
rect 13585 10345 13619 10379
rect 13653 10345 13687 10379
rect 13721 10345 13755 10379
rect 13789 10345 13823 10379
rect 13857 10345 13891 10379
rect 13925 10345 13959 10379
rect 13993 10345 14027 10379
rect 14061 10345 14095 10379
rect 14129 10345 14163 10379
rect 14197 10345 14231 10379
rect 14265 10345 14299 10379
rect 14333 10345 14367 10379
rect 14401 10345 14435 10379
rect 14469 10345 14503 10379
rect 14537 10345 14571 10379
rect 14605 10345 14639 10379
rect 14673 10345 14707 10379
rect 14741 10345 14775 10379
rect 14809 10345 14843 10379
rect 14877 10345 14911 10379
rect 14945 10345 14979 10379
rect 15013 10345 15047 10379
rect 15081 10345 15115 10379
rect 15149 10345 15183 10379
rect 15217 10345 15251 10379
rect 15285 10345 15319 10379
rect 15353 10345 15387 10379
rect 15421 10345 15455 10379
rect 15489 10345 15523 10379
rect 15557 10345 15591 10379
rect 15625 10345 15659 10379
rect 15693 10345 15727 10379
rect 15761 10345 15795 10379
rect 15829 10345 15884 10379
rect 13224 10311 15884 10345
rect 4421 10262 6239 10297
rect 4421 10228 4429 10262
rect 4463 10228 4497 10262
rect 4531 10228 4565 10262
rect 4599 10228 4633 10262
rect 4667 10228 4701 10262
rect 4735 10228 4769 10262
rect 4803 10228 4837 10262
rect 4871 10228 4905 10262
rect 4939 10228 4973 10262
rect 5007 10228 5041 10262
rect 5075 10228 5109 10262
rect 5143 10228 5177 10262
rect 5211 10228 5245 10262
rect 5279 10228 5313 10262
rect 5347 10228 5381 10262
rect 5415 10228 5449 10262
rect 5483 10228 5517 10262
rect 5551 10228 5585 10262
rect 5619 10228 5653 10262
rect 5687 10228 5721 10262
rect 5755 10228 5789 10262
rect 5823 10228 5857 10262
rect 5891 10228 5925 10262
rect 5959 10228 5993 10262
rect 6027 10228 6061 10262
rect 6095 10228 6129 10262
rect 6163 10228 6197 10262
rect 6231 10228 6239 10262
rect 4421 10193 6239 10228
rect 4421 10159 4429 10193
rect 4463 10159 4497 10193
rect 4531 10159 4565 10193
rect 4599 10159 4633 10193
rect 4667 10159 4701 10193
rect 4735 10159 4769 10193
rect 4803 10159 4837 10193
rect 4871 10159 4905 10193
rect 4939 10159 4973 10193
rect 5007 10159 5041 10193
rect 5075 10159 5109 10193
rect 5143 10159 5177 10193
rect 5211 10159 5245 10193
rect 5279 10159 5313 10193
rect 5347 10159 5381 10193
rect 5415 10159 5449 10193
rect 5483 10159 5517 10193
rect 5551 10159 5585 10193
rect 5619 10159 5653 10193
rect 5687 10159 5721 10193
rect 5755 10159 5789 10193
rect 5823 10159 5857 10193
rect 5891 10159 5925 10193
rect 5959 10159 5993 10193
rect 6027 10159 6061 10193
rect 6095 10159 6129 10193
rect 6163 10159 6197 10193
rect 6231 10159 6239 10193
rect 4421 10124 6239 10159
rect 4421 10090 4429 10124
rect 4463 10090 4497 10124
rect 4531 10090 4565 10124
rect 4599 10090 4633 10124
rect 4667 10090 4701 10124
rect 4735 10090 4769 10124
rect 4803 10090 4837 10124
rect 4871 10090 4905 10124
rect 4939 10090 4973 10124
rect 5007 10090 5041 10124
rect 5075 10090 5109 10124
rect 5143 10090 5177 10124
rect 5211 10090 5245 10124
rect 5279 10090 5313 10124
rect 5347 10090 5381 10124
rect 5415 10090 5449 10124
rect 5483 10090 5517 10124
rect 5551 10090 5585 10124
rect 5619 10090 5653 10124
rect 5687 10090 5721 10124
rect 5755 10090 5789 10124
rect 5823 10090 5857 10124
rect 5891 10090 5925 10124
rect 5959 10090 5993 10124
rect 6027 10090 6061 10124
rect 6095 10090 6129 10124
rect 6163 10090 6197 10124
rect 6231 10090 6239 10124
rect 4421 10066 6239 10090
rect 12479 10309 15884 10311
rect 12479 10275 13279 10309
rect 13313 10275 13347 10309
rect 13381 10275 13415 10309
rect 13449 10275 13483 10309
rect 13517 10275 13551 10309
rect 13585 10275 13619 10309
rect 13653 10275 13687 10309
rect 13721 10275 13755 10309
rect 13789 10275 13823 10309
rect 13857 10275 13891 10309
rect 13925 10275 13959 10309
rect 13993 10275 14027 10309
rect 14061 10275 14095 10309
rect 14129 10275 14163 10309
rect 14197 10275 14231 10309
rect 14265 10275 14299 10309
rect 14333 10275 14367 10309
rect 14401 10275 14435 10309
rect 14469 10275 14503 10309
rect 14537 10275 14571 10309
rect 14605 10275 14639 10309
rect 14673 10275 14707 10309
rect 14741 10275 14775 10309
rect 14809 10275 14843 10309
rect 14877 10275 14911 10309
rect 14945 10275 14979 10309
rect 15013 10275 15047 10309
rect 15081 10275 15115 10309
rect 15149 10275 15183 10309
rect 15217 10275 15251 10309
rect 15285 10275 15319 10309
rect 15353 10275 15387 10309
rect 15421 10275 15455 10309
rect 15489 10275 15523 10309
rect 15557 10275 15591 10309
rect 15625 10275 15659 10309
rect 15693 10275 15727 10309
rect 15761 10275 15795 10309
rect 15829 10275 15884 10309
rect 12479 10239 15884 10275
rect 12479 10205 13279 10239
rect 13313 10205 13347 10239
rect 13381 10205 13415 10239
rect 13449 10205 13483 10239
rect 13517 10205 13551 10239
rect 13585 10205 13619 10239
rect 13653 10205 13687 10239
rect 13721 10205 13755 10239
rect 13789 10205 13823 10239
rect 13857 10205 13891 10239
rect 13925 10205 13959 10239
rect 13993 10205 14027 10239
rect 14061 10205 14095 10239
rect 14129 10205 14163 10239
rect 14197 10205 14231 10239
rect 14265 10205 14299 10239
rect 14333 10205 14367 10239
rect 14401 10205 14435 10239
rect 14469 10205 14503 10239
rect 14537 10205 14571 10239
rect 14605 10205 14639 10239
rect 14673 10205 14707 10239
rect 14741 10205 14775 10239
rect 14809 10205 14843 10239
rect 14877 10205 14911 10239
rect 14945 10205 14979 10239
rect 15013 10205 15047 10239
rect 15081 10205 15115 10239
rect 15149 10205 15183 10239
rect 15217 10205 15251 10239
rect 15285 10205 15319 10239
rect 15353 10205 15387 10239
rect 15421 10205 15455 10239
rect 15489 10205 15523 10239
rect 15557 10205 15591 10239
rect 15625 10205 15659 10239
rect 15693 10205 15727 10239
rect 15761 10205 15795 10239
rect 15829 10205 15884 10239
rect 12479 10169 15884 10205
rect 12479 10162 13279 10169
rect 12479 10128 12504 10162
rect 12538 10128 12599 10162
rect 12633 10128 12694 10162
rect 12728 10128 12788 10162
rect 12822 10128 12882 10162
rect 12916 10128 12976 10162
rect 13010 10135 13279 10162
rect 13313 10135 13347 10169
rect 13381 10135 13415 10169
rect 13449 10135 13483 10169
rect 13517 10135 13551 10169
rect 13585 10135 13619 10169
rect 13653 10135 13687 10169
rect 13721 10135 13755 10169
rect 13789 10135 13823 10169
rect 13857 10135 13891 10169
rect 13925 10135 13959 10169
rect 13993 10135 14027 10169
rect 14061 10135 14095 10169
rect 14129 10135 14163 10169
rect 14197 10135 14231 10169
rect 14265 10135 14299 10169
rect 14333 10135 14367 10169
rect 14401 10135 14435 10169
rect 14469 10135 14503 10169
rect 14537 10135 14571 10169
rect 14605 10135 14639 10169
rect 14673 10135 14707 10169
rect 14741 10135 14775 10169
rect 14809 10135 14843 10169
rect 14877 10135 14911 10169
rect 14945 10135 14979 10169
rect 15013 10135 15047 10169
rect 15081 10135 15115 10169
rect 15149 10135 15183 10169
rect 15217 10135 15251 10169
rect 15285 10135 15319 10169
rect 15353 10135 15387 10169
rect 15421 10135 15455 10169
rect 15489 10135 15523 10169
rect 15557 10135 15591 10169
rect 15625 10135 15659 10169
rect 15693 10135 15727 10169
rect 15761 10135 15795 10169
rect 15829 10135 15884 10169
rect 13010 10128 15884 10135
rect 12479 10099 15884 10128
rect 12479 10094 13279 10099
rect 12479 10081 12504 10094
rect -2966 9999 -2959 10033
rect -2925 9999 -2891 10033
rect -2857 9999 -2823 10033
rect -2789 9999 -2755 10033
rect -2721 9999 -2687 10033
rect -2653 9999 -2619 10033
rect -2585 9999 -2551 10033
rect -2517 9999 -2483 10033
rect -2449 9999 -2415 10033
rect -2381 9999 -2347 10033
rect -2313 9999 -2279 10033
rect -2245 9999 -2211 10033
rect -2177 9999 -2143 10033
rect -2109 9999 -2075 10033
rect -2041 9999 -2007 10033
rect -1973 9999 -1939 10033
rect -1905 9999 -1871 10033
rect -1837 9999 -1803 10033
rect -1769 9999 -1735 10033
rect -1701 9999 -1667 10033
rect -1633 9999 -1599 10033
rect -1565 9999 -1531 10033
rect -1497 9999 -1463 10033
rect -1429 9999 -1395 10033
rect -1361 9999 -1327 10033
rect -1293 9999 -1259 10033
rect -1225 9999 -1191 10033
rect -1157 9999 -1123 10033
rect -1089 9999 -1055 10033
rect -1021 9999 -987 10033
rect -953 9999 -919 10033
rect -885 9999 -851 10033
rect -817 9999 -783 10033
rect -749 9999 -715 10033
rect -681 9999 -647 10033
rect -613 9999 -579 10033
rect -545 9999 -511 10033
rect -477 9999 -443 10033
rect -409 9999 -375 10033
rect -341 9999 -307 10033
rect -273 9999 -266 10033
rect -2966 9964 -266 9999
rect 12416 10060 12504 10081
rect 12538 10060 12599 10094
rect 12633 10060 12694 10094
rect 12728 10060 12788 10094
rect 12822 10060 12882 10094
rect 12916 10060 12976 10094
rect 13010 10065 13279 10094
rect 13313 10065 13347 10099
rect 13381 10065 13415 10099
rect 13449 10065 13483 10099
rect 13517 10065 13551 10099
rect 13585 10065 13619 10099
rect 13653 10065 13687 10099
rect 13721 10065 13755 10099
rect 13789 10065 13823 10099
rect 13857 10065 13891 10099
rect 13925 10065 13959 10099
rect 13993 10065 14027 10099
rect 14061 10065 14095 10099
rect 14129 10065 14163 10099
rect 14197 10065 14231 10099
rect 14265 10065 14299 10099
rect 14333 10065 14367 10099
rect 14401 10065 14435 10099
rect 14469 10065 14503 10099
rect 14537 10065 14571 10099
rect 14605 10065 14639 10099
rect 14673 10065 14707 10099
rect 14741 10065 14775 10099
rect 14809 10065 14843 10099
rect 14877 10065 14911 10099
rect 14945 10065 14979 10099
rect 15013 10065 15047 10099
rect 15081 10065 15115 10099
rect 15149 10065 15183 10099
rect 15217 10065 15251 10099
rect 15285 10065 15319 10099
rect 15353 10065 15387 10099
rect 15421 10065 15455 10099
rect 15489 10065 15523 10099
rect 15557 10065 15591 10099
rect 15625 10065 15659 10099
rect 15693 10065 15727 10099
rect 15761 10065 15795 10099
rect 15829 10065 15884 10099
rect 13010 10060 15884 10065
rect 12416 10056 15884 10060
rect 12416 10026 13077 10056
rect 12416 9992 12504 10026
rect 12538 9992 12599 10026
rect 12633 9992 12694 10026
rect 12728 9992 12788 10026
rect 12822 9992 12882 10026
rect 12916 9992 12976 10026
rect 13010 10022 13077 10026
rect 13111 10022 13160 10056
rect 13194 10029 15884 10056
rect 13194 10022 13279 10029
rect 13010 9995 13279 10022
rect 13313 9995 13347 10029
rect 13381 9995 13415 10029
rect 13449 9995 13483 10029
rect 13517 9995 13551 10029
rect 13585 9995 13619 10029
rect 13653 9995 13687 10029
rect 13721 9995 13755 10029
rect 13789 9995 13823 10029
rect 13857 9995 13891 10029
rect 13925 9995 13959 10029
rect 13993 9995 14027 10029
rect 14061 9995 14095 10029
rect 14129 9995 14163 10029
rect 14197 9995 14231 10029
rect 14265 9995 14299 10029
rect 14333 9995 14367 10029
rect 14401 9995 14435 10029
rect 14469 9995 14503 10029
rect 14537 9995 14571 10029
rect 14605 9995 14639 10029
rect 14673 9995 14707 10029
rect 14741 9995 14775 10029
rect 14809 9995 14843 10029
rect 14877 9995 14911 10029
rect 14945 9995 14979 10029
rect 15013 9995 15047 10029
rect 15081 9995 15115 10029
rect 15149 9995 15183 10029
rect 15217 9995 15251 10029
rect 15285 9995 15319 10029
rect 15353 9995 15387 10029
rect 15421 9995 15455 10029
rect 15489 9995 15523 10029
rect 15557 9995 15591 10029
rect 15625 9995 15659 10029
rect 15693 9995 15727 10029
rect 15761 9995 15795 10029
rect 15829 9995 15884 10029
rect 13010 9992 15194 9995
rect -2966 9930 -2959 9964
rect -2925 9930 -2891 9964
rect -2857 9930 -2823 9964
rect -2789 9930 -2755 9964
rect -2721 9930 -2687 9964
rect -2653 9930 -2619 9964
rect -2585 9930 -2551 9964
rect -2517 9930 -2483 9964
rect -2449 9930 -2415 9964
rect -2381 9930 -2347 9964
rect -2313 9930 -2279 9964
rect -2245 9930 -2211 9964
rect -2177 9930 -2143 9964
rect -2109 9930 -2075 9964
rect -2041 9930 -2007 9964
rect -1973 9930 -1939 9964
rect -1905 9930 -1871 9964
rect -1837 9930 -1803 9964
rect -1769 9930 -1735 9964
rect -1701 9930 -1667 9964
rect -1633 9930 -1599 9964
rect -1565 9930 -1531 9964
rect -1497 9930 -1463 9964
rect -1429 9930 -1395 9964
rect -1361 9930 -1327 9964
rect -1293 9930 -1259 9964
rect -1225 9930 -1191 9964
rect -1157 9930 -1123 9964
rect -1089 9930 -1055 9964
rect -1021 9930 -987 9964
rect -953 9930 -919 9964
rect -885 9930 -851 9964
rect -817 9930 -783 9964
rect -749 9930 -715 9964
rect -681 9930 -647 9964
rect -613 9930 -579 9964
rect -545 9930 -511 9964
rect -477 9930 -443 9964
rect -409 9930 -375 9964
rect -341 9930 -307 9964
rect -273 9930 -266 9964
rect -2966 9895 -266 9930
rect 7505 9925 7555 9980
rect 12416 9958 15194 9992
rect 12416 9952 13587 9958
rect 12416 9947 12553 9952
rect -2966 9861 -2959 9895
rect -2925 9861 -2891 9895
rect -2857 9861 -2823 9895
rect -2789 9861 -2755 9895
rect -2721 9861 -2687 9895
rect -2653 9861 -2619 9895
rect -2585 9861 -2551 9895
rect -2517 9861 -2483 9895
rect -2449 9861 -2415 9895
rect -2381 9861 -2347 9895
rect -2313 9861 -2279 9895
rect -2245 9861 -2211 9895
rect -2177 9861 -2143 9895
rect -2109 9861 -2075 9895
rect -2041 9861 -2007 9895
rect -1973 9861 -1939 9895
rect -1905 9861 -1871 9895
rect -1837 9861 -1803 9895
rect -1769 9861 -1735 9895
rect -1701 9861 -1667 9895
rect -1633 9861 -1599 9895
rect -1565 9861 -1531 9895
rect -1497 9861 -1463 9895
rect -1429 9861 -1395 9895
rect -1361 9861 -1327 9895
rect -1293 9861 -1259 9895
rect -1225 9861 -1191 9895
rect -1157 9861 -1123 9895
rect -1089 9861 -1055 9895
rect -1021 9861 -987 9895
rect -953 9861 -919 9895
rect -885 9861 -851 9895
rect -817 9861 -783 9895
rect -749 9861 -715 9895
rect -681 9861 -647 9895
rect -613 9861 -579 9895
rect -545 9861 -511 9895
rect -477 9861 -443 9895
rect -409 9861 -375 9895
rect -341 9861 -307 9895
rect -273 9861 -266 9895
rect -2966 9826 -266 9861
rect 11650 9850 11696 9864
rect -2966 9792 -2959 9826
rect -2925 9792 -2891 9826
rect -2857 9792 -2823 9826
rect -2789 9792 -2755 9826
rect -2721 9792 -2687 9826
rect -2653 9792 -2619 9826
rect -2585 9792 -2551 9826
rect -2517 9792 -2483 9826
rect -2449 9792 -2415 9826
rect -2381 9792 -2347 9826
rect -2313 9792 -2279 9826
rect -2245 9792 -2211 9826
rect -2177 9792 -2143 9826
rect -2109 9792 -2075 9826
rect -2041 9792 -2007 9826
rect -1973 9792 -1939 9826
rect -1905 9792 -1871 9826
rect -1837 9792 -1803 9826
rect -1769 9792 -1735 9826
rect -1701 9792 -1667 9826
rect -1633 9792 -1599 9826
rect -1565 9792 -1531 9826
rect -1497 9792 -1463 9826
rect -1429 9792 -1395 9826
rect -1361 9792 -1327 9826
rect -1293 9792 -1259 9826
rect -1225 9792 -1191 9826
rect -1157 9792 -1123 9826
rect -1089 9792 -1055 9826
rect -1021 9792 -987 9826
rect -953 9792 -919 9826
rect -885 9792 -851 9826
rect -817 9792 -783 9826
rect -749 9792 -715 9826
rect -681 9792 -647 9826
rect -613 9792 -579 9826
rect -545 9792 -511 9826
rect -477 9792 -443 9826
rect -409 9792 -375 9826
rect -341 9792 -307 9826
rect -273 9792 -266 9826
rect -2966 9757 -266 9792
rect -2966 9723 -2959 9757
rect -2925 9723 -2891 9757
rect -2857 9723 -2823 9757
rect -2789 9723 -2755 9757
rect -2721 9723 -2687 9757
rect -2653 9723 -2619 9757
rect -2585 9723 -2551 9757
rect -2517 9723 -2483 9757
rect -2449 9723 -2415 9757
rect -2381 9723 -2347 9757
rect -2313 9723 -2279 9757
rect -2245 9723 -2211 9757
rect -2177 9723 -2143 9757
rect -2109 9723 -2075 9757
rect -2041 9723 -2007 9757
rect -1973 9723 -1939 9757
rect -1905 9723 -1871 9757
rect -1837 9723 -1803 9757
rect -1769 9723 -1735 9757
rect -1701 9723 -1667 9757
rect -1633 9723 -1599 9757
rect -1565 9723 -1531 9757
rect -1497 9723 -1463 9757
rect -1429 9723 -1395 9757
rect -1361 9723 -1327 9757
rect -1293 9723 -1259 9757
rect -1225 9723 -1191 9757
rect -1157 9723 -1123 9757
rect -1089 9723 -1055 9757
rect -1021 9723 -987 9757
rect -953 9723 -919 9757
rect -885 9723 -851 9757
rect -817 9723 -783 9757
rect -749 9723 -715 9757
rect -681 9723 -647 9757
rect -613 9723 -579 9757
rect -545 9723 -511 9757
rect -477 9723 -443 9757
rect -409 9723 -375 9757
rect -341 9723 -307 9757
rect -273 9723 -266 9757
rect -2966 9688 -266 9723
rect -2966 9654 -2959 9688
rect -2925 9654 -2891 9688
rect -2857 9654 -2823 9688
rect -2789 9654 -2755 9688
rect -2721 9654 -2687 9688
rect -2653 9654 -2619 9688
rect -2585 9654 -2551 9688
rect -2517 9654 -2483 9688
rect -2449 9654 -2415 9688
rect -2381 9654 -2347 9688
rect -2313 9654 -2279 9688
rect -2245 9654 -2211 9688
rect -2177 9654 -2143 9688
rect -2109 9654 -2075 9688
rect -2041 9654 -2007 9688
rect -1973 9654 -1939 9688
rect -1905 9654 -1871 9688
rect -1837 9654 -1803 9688
rect -1769 9654 -1735 9688
rect -1701 9654 -1667 9688
rect -1633 9654 -1599 9688
rect -1565 9654 -1531 9688
rect -1497 9654 -1463 9688
rect -1429 9654 -1395 9688
rect -1361 9654 -1327 9688
rect -1293 9654 -1259 9688
rect -1225 9654 -1191 9688
rect -1157 9654 -1123 9688
rect -1089 9654 -1055 9688
rect -1021 9654 -987 9688
rect -953 9654 -919 9688
rect -885 9654 -851 9688
rect -817 9654 -783 9688
rect -749 9654 -715 9688
rect -681 9654 -647 9688
rect -613 9654 -579 9688
rect -545 9654 -511 9688
rect -477 9654 -443 9688
rect -409 9654 -375 9688
rect -341 9654 -307 9688
rect -273 9654 -266 9688
rect -2966 9619 -266 9654
rect -2966 9585 -2959 9619
rect -2925 9585 -2891 9619
rect -2857 9585 -2823 9619
rect -2789 9585 -2755 9619
rect -2721 9585 -2687 9619
rect -2653 9585 -2619 9619
rect -2585 9585 -2551 9619
rect -2517 9585 -2483 9619
rect -2449 9585 -2415 9619
rect -2381 9585 -2347 9619
rect -2313 9585 -2279 9619
rect -2245 9585 -2211 9619
rect -2177 9585 -2143 9619
rect -2109 9585 -2075 9619
rect -2041 9585 -2007 9619
rect -1973 9585 -1939 9619
rect -1905 9585 -1871 9619
rect -1837 9585 -1803 9619
rect -1769 9585 -1735 9619
rect -1701 9585 -1667 9619
rect -1633 9585 -1599 9619
rect -1565 9585 -1531 9619
rect -1497 9585 -1463 9619
rect -1429 9585 -1395 9619
rect -1361 9585 -1327 9619
rect -1293 9585 -1259 9619
rect -1225 9585 -1191 9619
rect -1157 9585 -1123 9619
rect -1089 9585 -1055 9619
rect -1021 9585 -987 9619
rect -953 9585 -919 9619
rect -885 9585 -851 9619
rect -817 9585 -783 9619
rect -749 9585 -715 9619
rect -681 9585 -647 9619
rect -613 9585 -579 9619
rect -545 9585 -511 9619
rect -477 9585 -443 9619
rect -409 9585 -375 9619
rect -341 9585 -307 9619
rect -273 9585 -266 9619
rect -2966 9550 -266 9585
rect -2966 9516 -2959 9550
rect -2925 9516 -2891 9550
rect -2857 9516 -2823 9550
rect -2789 9516 -2755 9550
rect -2721 9516 -2687 9550
rect -2653 9516 -2619 9550
rect -2585 9516 -2551 9550
rect -2517 9516 -2483 9550
rect -2449 9516 -2415 9550
rect -2381 9516 -2347 9550
rect -2313 9516 -2279 9550
rect -2245 9516 -2211 9550
rect -2177 9516 -2143 9550
rect -2109 9516 -2075 9550
rect -2041 9516 -2007 9550
rect -1973 9516 -1939 9550
rect -1905 9516 -1871 9550
rect -1837 9516 -1803 9550
rect -1769 9516 -1735 9550
rect -1701 9516 -1667 9550
rect -1633 9516 -1599 9550
rect -1565 9516 -1531 9550
rect -1497 9516 -1463 9550
rect -1429 9516 -1395 9550
rect -1361 9516 -1327 9550
rect -1293 9516 -1259 9550
rect -1225 9516 -1191 9550
rect -1157 9516 -1123 9550
rect -1089 9516 -1055 9550
rect -1021 9516 -987 9550
rect -953 9516 -919 9550
rect -885 9516 -851 9550
rect -817 9516 -783 9550
rect -749 9516 -715 9550
rect -681 9516 -647 9550
rect -613 9516 -579 9550
rect -545 9516 -511 9550
rect -477 9516 -443 9550
rect -409 9516 -375 9550
rect -341 9516 -307 9550
rect -273 9516 -266 9550
rect -2966 9481 -266 9516
rect -2966 9447 -2959 9481
rect -2925 9447 -2891 9481
rect -2857 9447 -2823 9481
rect -2789 9447 -2755 9481
rect -2721 9447 -2687 9481
rect -2653 9447 -2619 9481
rect -2585 9447 -2551 9481
rect -2517 9447 -2483 9481
rect -2449 9447 -2415 9481
rect -2381 9447 -2347 9481
rect -2313 9447 -2279 9481
rect -2245 9447 -2211 9481
rect -2177 9447 -2143 9481
rect -2109 9447 -2075 9481
rect -2041 9447 -2007 9481
rect -1973 9447 -1939 9481
rect -1905 9447 -1871 9481
rect -1837 9447 -1803 9481
rect -1769 9447 -1735 9481
rect -1701 9447 -1667 9481
rect -1633 9447 -1599 9481
rect -1565 9447 -1531 9481
rect -1497 9447 -1463 9481
rect -1429 9447 -1395 9481
rect -1361 9447 -1327 9481
rect -1293 9447 -1259 9481
rect -1225 9447 -1191 9481
rect -1157 9447 -1123 9481
rect -1089 9447 -1055 9481
rect -1021 9447 -987 9481
rect -953 9447 -919 9481
rect -885 9447 -851 9481
rect -817 9447 -783 9481
rect -749 9447 -715 9481
rect -681 9447 -647 9481
rect -613 9447 -579 9481
rect -545 9447 -511 9481
rect -477 9447 -443 9481
rect -409 9447 -375 9481
rect -341 9447 -307 9481
rect -273 9447 -266 9481
rect -2966 9412 -266 9447
rect -2966 9378 -2959 9412
rect -2925 9378 -2891 9412
rect -2857 9378 -2823 9412
rect -2789 9378 -2755 9412
rect -2721 9378 -2687 9412
rect -2653 9378 -2619 9412
rect -2585 9378 -2551 9412
rect -2517 9378 -2483 9412
rect -2449 9378 -2415 9412
rect -2381 9378 -2347 9412
rect -2313 9378 -2279 9412
rect -2245 9378 -2211 9412
rect -2177 9378 -2143 9412
rect -2109 9378 -2075 9412
rect -2041 9378 -2007 9412
rect -1973 9378 -1939 9412
rect -1905 9378 -1871 9412
rect -1837 9378 -1803 9412
rect -1769 9378 -1735 9412
rect -1701 9378 -1667 9412
rect -1633 9378 -1599 9412
rect -1565 9378 -1531 9412
rect -1497 9378 -1463 9412
rect -1429 9378 -1395 9412
rect -1361 9378 -1327 9412
rect -1293 9378 -1259 9412
rect -1225 9378 -1191 9412
rect -1157 9378 -1123 9412
rect -1089 9378 -1055 9412
rect -1021 9378 -987 9412
rect -953 9378 -919 9412
rect -885 9378 -851 9412
rect -817 9378 -783 9412
rect -749 9378 -715 9412
rect -681 9378 -647 9412
rect -613 9378 -579 9412
rect -545 9378 -511 9412
rect -477 9378 -443 9412
rect -409 9378 -375 9412
rect -341 9378 -307 9412
rect -273 9378 -266 9412
rect -2966 9343 -266 9378
rect -2966 9309 -2959 9343
rect -2925 9309 -2891 9343
rect -2857 9309 -2823 9343
rect -2789 9309 -2755 9343
rect -2721 9309 -2687 9343
rect -2653 9309 -2619 9343
rect -2585 9309 -2551 9343
rect -2517 9309 -2483 9343
rect -2449 9309 -2415 9343
rect -2381 9309 -2347 9343
rect -2313 9309 -2279 9343
rect -2245 9309 -2211 9343
rect -2177 9309 -2143 9343
rect -2109 9309 -2075 9343
rect -2041 9309 -2007 9343
rect -1973 9309 -1939 9343
rect -1905 9309 -1871 9343
rect -1837 9309 -1803 9343
rect -1769 9309 -1735 9343
rect -1701 9309 -1667 9343
rect -1633 9309 -1599 9343
rect -1565 9309 -1531 9343
rect -1497 9309 -1463 9343
rect -1429 9309 -1395 9343
rect -1361 9309 -1327 9343
rect -1293 9309 -1259 9343
rect -1225 9309 -1191 9343
rect -1157 9309 -1123 9343
rect -1089 9309 -1055 9343
rect -1021 9309 -987 9343
rect -953 9309 -919 9343
rect -885 9309 -851 9343
rect -817 9309 -783 9343
rect -749 9309 -715 9343
rect -681 9309 -647 9343
rect -613 9309 -579 9343
rect -545 9309 -511 9343
rect -477 9309 -443 9343
rect -409 9309 -375 9343
rect -341 9309 -307 9343
rect -273 9309 -266 9343
rect -2966 9274 -266 9309
rect -2966 9240 -2959 9274
rect -2925 9240 -2891 9274
rect -2857 9240 -2823 9274
rect -2789 9240 -2755 9274
rect -2721 9240 -2687 9274
rect -2653 9240 -2619 9274
rect -2585 9240 -2551 9274
rect -2517 9240 -2483 9274
rect -2449 9240 -2415 9274
rect -2381 9240 -2347 9274
rect -2313 9240 -2279 9274
rect -2245 9240 -2211 9274
rect -2177 9240 -2143 9274
rect -2109 9240 -2075 9274
rect -2041 9240 -2007 9274
rect -1973 9240 -1939 9274
rect -1905 9240 -1871 9274
rect -1837 9240 -1803 9274
rect -1769 9240 -1735 9274
rect -1701 9240 -1667 9274
rect -1633 9240 -1599 9274
rect -1565 9240 -1531 9274
rect -1497 9240 -1463 9274
rect -1429 9240 -1395 9274
rect -1361 9240 -1327 9274
rect -1293 9240 -1259 9274
rect -1225 9240 -1191 9274
rect -1157 9240 -1123 9274
rect -1089 9240 -1055 9274
rect -1021 9240 -987 9274
rect -953 9240 -919 9274
rect -885 9240 -851 9274
rect -817 9240 -783 9274
rect -749 9240 -715 9274
rect -681 9240 -647 9274
rect -613 9240 -579 9274
rect -545 9240 -511 9274
rect -477 9240 -443 9274
rect -409 9240 -375 9274
rect -341 9240 -307 9274
rect -273 9240 -266 9274
rect -2966 9205 -266 9240
rect -2966 9171 -2959 9205
rect -2925 9171 -2891 9205
rect -2857 9171 -2823 9205
rect -2789 9171 -2755 9205
rect -2721 9171 -2687 9205
rect -2653 9171 -2619 9205
rect -2585 9171 -2551 9205
rect -2517 9171 -2483 9205
rect -2449 9171 -2415 9205
rect -2381 9171 -2347 9205
rect -2313 9171 -2279 9205
rect -2245 9171 -2211 9205
rect -2177 9171 -2143 9205
rect -2109 9171 -2075 9205
rect -2041 9171 -2007 9205
rect -1973 9171 -1939 9205
rect -1905 9171 -1871 9205
rect -1837 9171 -1803 9205
rect -1769 9171 -1735 9205
rect -1701 9171 -1667 9205
rect -1633 9171 -1599 9205
rect -1565 9171 -1531 9205
rect -1497 9171 -1463 9205
rect -1429 9171 -1395 9205
rect -1361 9171 -1327 9205
rect -1293 9171 -1259 9205
rect -1225 9171 -1191 9205
rect -1157 9171 -1123 9205
rect -1089 9171 -1055 9205
rect -1021 9171 -987 9205
rect -953 9171 -919 9205
rect -885 9171 -851 9205
rect -817 9171 -783 9205
rect -749 9171 -715 9205
rect -681 9171 -647 9205
rect -613 9171 -579 9205
rect -545 9171 -511 9205
rect -477 9171 -443 9205
rect -409 9171 -375 9205
rect -341 9171 -307 9205
rect -273 9171 -266 9205
rect -2966 9136 -266 9171
rect -2966 9102 -2959 9136
rect -2925 9102 -2891 9136
rect -2857 9102 -2823 9136
rect -2789 9102 -2755 9136
rect -2721 9102 -2687 9136
rect -2653 9102 -2619 9136
rect -2585 9102 -2551 9136
rect -2517 9102 -2483 9136
rect -2449 9102 -2415 9136
rect -2381 9102 -2347 9136
rect -2313 9102 -2279 9136
rect -2245 9102 -2211 9136
rect -2177 9102 -2143 9136
rect -2109 9102 -2075 9136
rect -2041 9102 -2007 9136
rect -1973 9102 -1939 9136
rect -1905 9102 -1871 9136
rect -1837 9102 -1803 9136
rect -1769 9102 -1735 9136
rect -1701 9102 -1667 9136
rect -1633 9102 -1599 9136
rect -1565 9102 -1531 9136
rect -1497 9102 -1463 9136
rect -1429 9102 -1395 9136
rect -1361 9102 -1327 9136
rect -1293 9102 -1259 9136
rect -1225 9102 -1191 9136
rect -1157 9102 -1123 9136
rect -1089 9102 -1055 9136
rect -1021 9102 -987 9136
rect -953 9102 -919 9136
rect -885 9102 -851 9136
rect -817 9102 -783 9136
rect -749 9102 -715 9136
rect -681 9102 -647 9136
rect -613 9102 -579 9136
rect -545 9102 -511 9136
rect -477 9102 -443 9136
rect -409 9102 -375 9136
rect -341 9102 -307 9136
rect -273 9102 -266 9136
rect -2966 9067 -266 9102
rect -2966 9033 -2959 9067
rect -2925 9033 -2891 9067
rect -2857 9033 -2823 9067
rect -2789 9033 -2755 9067
rect -2721 9033 -2687 9067
rect -2653 9033 -2619 9067
rect -2585 9033 -2551 9067
rect -2517 9033 -2483 9067
rect -2449 9033 -2415 9067
rect -2381 9033 -2347 9067
rect -2313 9033 -2279 9067
rect -2245 9033 -2211 9067
rect -2177 9033 -2143 9067
rect -2109 9033 -2075 9067
rect -2041 9033 -2007 9067
rect -1973 9033 -1939 9067
rect -1905 9033 -1871 9067
rect -1837 9033 -1803 9067
rect -1769 9033 -1735 9067
rect -1701 9033 -1667 9067
rect -1633 9033 -1599 9067
rect -1565 9033 -1531 9067
rect -1497 9033 -1463 9067
rect -1429 9033 -1395 9067
rect -1361 9033 -1327 9067
rect -1293 9033 -1259 9067
rect -1225 9033 -1191 9067
rect -1157 9033 -1123 9067
rect -1089 9033 -1055 9067
rect -1021 9033 -987 9067
rect -953 9033 -919 9067
rect -885 9033 -851 9067
rect -817 9033 -783 9067
rect -749 9033 -715 9067
rect -681 9033 -647 9067
rect -613 9033 -579 9067
rect -545 9033 -511 9067
rect -477 9033 -443 9067
rect -409 9033 -375 9067
rect -341 9033 -307 9067
rect -273 9033 -266 9067
rect -2966 8998 -266 9033
rect -2966 8964 -2959 8998
rect -2925 8964 -2891 8998
rect -2857 8964 -2823 8998
rect -2789 8964 -2755 8998
rect -2721 8964 -2687 8998
rect -2653 8964 -2619 8998
rect -2585 8964 -2551 8998
rect -2517 8964 -2483 8998
rect -2449 8964 -2415 8998
rect -2381 8964 -2347 8998
rect -2313 8964 -2279 8998
rect -2245 8964 -2211 8998
rect -2177 8964 -2143 8998
rect -2109 8964 -2075 8998
rect -2041 8964 -2007 8998
rect -1973 8964 -1939 8998
rect -1905 8964 -1871 8998
rect -1837 8964 -1803 8998
rect -1769 8964 -1735 8998
rect -1701 8964 -1667 8998
rect -1633 8964 -1599 8998
rect -1565 8964 -1531 8998
rect -1497 8964 -1463 8998
rect -1429 8964 -1395 8998
rect -1361 8964 -1327 8998
rect -1293 8964 -1259 8998
rect -1225 8964 -1191 8998
rect -1157 8964 -1123 8998
rect -1089 8964 -1055 8998
rect -1021 8964 -987 8998
rect -953 8964 -919 8998
rect -885 8964 -851 8998
rect -817 8964 -783 8998
rect -749 8964 -715 8998
rect -681 8964 -647 8998
rect -613 8964 -579 8998
rect -545 8964 -511 8998
rect -477 8964 -443 8998
rect -409 8964 -375 8998
rect -341 8964 -307 8998
rect -273 8964 -266 8998
rect -2966 8929 -266 8964
rect -2966 8895 -2959 8929
rect -2925 8895 -2891 8929
rect -2857 8895 -2823 8929
rect -2789 8895 -2755 8929
rect -2721 8895 -2687 8929
rect -2653 8895 -2619 8929
rect -2585 8895 -2551 8929
rect -2517 8895 -2483 8929
rect -2449 8895 -2415 8929
rect -2381 8895 -2347 8929
rect -2313 8895 -2279 8929
rect -2245 8895 -2211 8929
rect -2177 8895 -2143 8929
rect -2109 8895 -2075 8929
rect -2041 8895 -2007 8929
rect -1973 8895 -1939 8929
rect -1905 8895 -1871 8929
rect -1837 8895 -1803 8929
rect -1769 8895 -1735 8929
rect -1701 8895 -1667 8929
rect -1633 8895 -1599 8929
rect -1565 8895 -1531 8929
rect -1497 8895 -1463 8929
rect -1429 8895 -1395 8929
rect -1361 8895 -1327 8929
rect -1293 8895 -1259 8929
rect -1225 8895 -1191 8929
rect -1157 8895 -1123 8929
rect -1089 8895 -1055 8929
rect -1021 8895 -987 8929
rect -953 8895 -919 8929
rect -885 8895 -851 8929
rect -817 8895 -783 8929
rect -749 8895 -715 8929
rect -681 8895 -647 8929
rect -613 8895 -579 8929
rect -545 8895 -511 8929
rect -477 8895 -443 8929
rect -409 8895 -375 8929
rect -341 8895 -307 8929
rect -273 8895 -266 8929
rect -2966 8860 -266 8895
rect -2966 8826 -2959 8860
rect -2925 8826 -2891 8860
rect -2857 8826 -2823 8860
rect -2789 8826 -2755 8860
rect -2721 8826 -2687 8860
rect -2653 8826 -2619 8860
rect -2585 8826 -2551 8860
rect -2517 8826 -2483 8860
rect -2449 8826 -2415 8860
rect -2381 8826 -2347 8860
rect -2313 8826 -2279 8860
rect -2245 8826 -2211 8860
rect -2177 8826 -2143 8860
rect -2109 8826 -2075 8860
rect -2041 8826 -2007 8860
rect -1973 8826 -1939 8860
rect -1905 8826 -1871 8860
rect -1837 8826 -1803 8860
rect -1769 8826 -1735 8860
rect -1701 8826 -1667 8860
rect -1633 8826 -1599 8860
rect -1565 8826 -1531 8860
rect -1497 8826 -1463 8860
rect -1429 8826 -1395 8860
rect -1361 8826 -1327 8860
rect -1293 8826 -1259 8860
rect -1225 8826 -1191 8860
rect -1157 8826 -1123 8860
rect -1089 8826 -1055 8860
rect -1021 8826 -987 8860
rect -953 8826 -919 8860
rect -885 8826 -851 8860
rect -817 8826 -783 8860
rect -749 8826 -715 8860
rect -681 8826 -647 8860
rect -613 8826 -579 8860
rect -545 8826 -511 8860
rect -477 8826 -443 8860
rect -409 8826 -375 8860
rect -341 8826 -307 8860
rect -273 8826 -266 8860
rect -2966 8791 -266 8826
rect -2966 8757 -2959 8791
rect -2925 8757 -2891 8791
rect -2857 8757 -2823 8791
rect -2789 8757 -2755 8791
rect -2721 8757 -2687 8791
rect -2653 8757 -2619 8791
rect -2585 8757 -2551 8791
rect -2517 8757 -2483 8791
rect -2449 8757 -2415 8791
rect -2381 8757 -2347 8791
rect -2313 8757 -2279 8791
rect -2245 8757 -2211 8791
rect -2177 8757 -2143 8791
rect -2109 8757 -2075 8791
rect -2041 8757 -2007 8791
rect -1973 8757 -1939 8791
rect -1905 8757 -1871 8791
rect -1837 8757 -1803 8791
rect -1769 8757 -1735 8791
rect -1701 8757 -1667 8791
rect -1633 8757 -1599 8791
rect -1565 8757 -1531 8791
rect -1497 8757 -1463 8791
rect -1429 8757 -1395 8791
rect -1361 8757 -1327 8791
rect -1293 8757 -1259 8791
rect -1225 8757 -1191 8791
rect -1157 8757 -1123 8791
rect -1089 8757 -1055 8791
rect -1021 8757 -987 8791
rect -953 8757 -919 8791
rect -885 8757 -851 8791
rect -817 8757 -783 8791
rect -749 8757 -715 8791
rect -681 8757 -647 8791
rect -613 8757 -579 8791
rect -545 8757 -511 8791
rect -477 8757 -443 8791
rect -409 8757 -375 8791
rect -341 8757 -307 8791
rect -273 8757 -266 8791
rect -2966 8722 -266 8757
rect -2966 8688 -2959 8722
rect -2925 8688 -2891 8722
rect -2857 8688 -2823 8722
rect -2789 8688 -2755 8722
rect -2721 8688 -2687 8722
rect -2653 8688 -2619 8722
rect -2585 8688 -2551 8722
rect -2517 8688 -2483 8722
rect -2449 8688 -2415 8722
rect -2381 8688 -2347 8722
rect -2313 8688 -2279 8722
rect -2245 8688 -2211 8722
rect -2177 8688 -2143 8722
rect -2109 8688 -2075 8722
rect -2041 8688 -2007 8722
rect -1973 8688 -1939 8722
rect -1905 8688 -1871 8722
rect -1837 8688 -1803 8722
rect -1769 8688 -1735 8722
rect -1701 8688 -1667 8722
rect -1633 8688 -1599 8722
rect -1565 8688 -1531 8722
rect -1497 8688 -1463 8722
rect -1429 8688 -1395 8722
rect -1361 8688 -1327 8722
rect -1293 8688 -1259 8722
rect -1225 8688 -1191 8722
rect -1157 8688 -1123 8722
rect -1089 8688 -1055 8722
rect -1021 8688 -987 8722
rect -953 8688 -919 8722
rect -885 8688 -851 8722
rect -817 8688 -783 8722
rect -749 8688 -715 8722
rect -681 8688 -647 8722
rect -613 8688 -579 8722
rect -545 8688 -511 8722
rect -477 8688 -443 8722
rect -409 8688 -375 8722
rect -341 8688 -307 8722
rect -273 8688 -266 8722
rect -2966 8653 -266 8688
rect -2966 8619 -2959 8653
rect -2925 8619 -2891 8653
rect -2857 8619 -2823 8653
rect -2789 8619 -2755 8653
rect -2721 8619 -2687 8653
rect -2653 8619 -2619 8653
rect -2585 8619 -2551 8653
rect -2517 8619 -2483 8653
rect -2449 8619 -2415 8653
rect -2381 8619 -2347 8653
rect -2313 8619 -2279 8653
rect -2245 8619 -2211 8653
rect -2177 8619 -2143 8653
rect -2109 8619 -2075 8653
rect -2041 8619 -2007 8653
rect -1973 8619 -1939 8653
rect -1905 8619 -1871 8653
rect -1837 8619 -1803 8653
rect -1769 8619 -1735 8653
rect -1701 8619 -1667 8653
rect -1633 8619 -1599 8653
rect -1565 8619 -1531 8653
rect -1497 8619 -1463 8653
rect -1429 8619 -1395 8653
rect -1361 8619 -1327 8653
rect -1293 8619 -1259 8653
rect -1225 8619 -1191 8653
rect -1157 8619 -1123 8653
rect -1089 8619 -1055 8653
rect -1021 8619 -987 8653
rect -953 8619 -919 8653
rect -885 8619 -851 8653
rect -817 8619 -783 8653
rect -749 8619 -715 8653
rect -681 8619 -647 8653
rect -613 8619 -579 8653
rect -545 8619 -511 8653
rect -477 8619 -443 8653
rect -409 8619 -375 8653
rect -341 8619 -307 8653
rect -273 8619 -266 8653
rect -2966 8584 -266 8619
rect -2966 8550 -2959 8584
rect -2925 8550 -2891 8584
rect -2857 8550 -2823 8584
rect -2789 8550 -2755 8584
rect -2721 8550 -2687 8584
rect -2653 8550 -2619 8584
rect -2585 8550 -2551 8584
rect -2517 8550 -2483 8584
rect -2449 8550 -2415 8584
rect -2381 8550 -2347 8584
rect -2313 8550 -2279 8584
rect -2245 8550 -2211 8584
rect -2177 8550 -2143 8584
rect -2109 8550 -2075 8584
rect -2041 8550 -2007 8584
rect -1973 8550 -1939 8584
rect -1905 8550 -1871 8584
rect -1837 8550 -1803 8584
rect -1769 8550 -1735 8584
rect -1701 8550 -1667 8584
rect -1633 8550 -1599 8584
rect -1565 8550 -1531 8584
rect -1497 8550 -1463 8584
rect -1429 8550 -1395 8584
rect -1361 8550 -1327 8584
rect -1293 8550 -1259 8584
rect -1225 8550 -1191 8584
rect -1157 8550 -1123 8584
rect -1089 8550 -1055 8584
rect -1021 8550 -987 8584
rect -953 8550 -919 8584
rect -885 8550 -851 8584
rect -817 8550 -783 8584
rect -749 8550 -715 8584
rect -681 8550 -647 8584
rect -613 8550 -579 8584
rect -545 8550 -511 8584
rect -477 8550 -443 8584
rect -409 8550 -375 8584
rect -341 8550 -307 8584
rect -273 8550 -266 8584
rect -2966 8515 -266 8550
rect -2966 8481 -2959 8515
rect -2925 8481 -2891 8515
rect -2857 8481 -2823 8515
rect -2789 8481 -2755 8515
rect -2721 8481 -2687 8515
rect -2653 8481 -2619 8515
rect -2585 8481 -2551 8515
rect -2517 8481 -2483 8515
rect -2449 8481 -2415 8515
rect -2381 8481 -2347 8515
rect -2313 8481 -2279 8515
rect -2245 8481 -2211 8515
rect -2177 8481 -2143 8515
rect -2109 8481 -2075 8515
rect -2041 8481 -2007 8515
rect -1973 8481 -1939 8515
rect -1905 8481 -1871 8515
rect -1837 8481 -1803 8515
rect -1769 8481 -1735 8515
rect -1701 8481 -1667 8515
rect -1633 8481 -1599 8515
rect -1565 8481 -1531 8515
rect -1497 8481 -1463 8515
rect -1429 8481 -1395 8515
rect -1361 8481 -1327 8515
rect -1293 8481 -1259 8515
rect -1225 8481 -1191 8515
rect -1157 8481 -1123 8515
rect -1089 8481 -1055 8515
rect -1021 8481 -987 8515
rect -953 8481 -919 8515
rect -885 8481 -851 8515
rect -817 8481 -783 8515
rect -749 8481 -715 8515
rect -681 8481 -647 8515
rect -613 8481 -579 8515
rect -545 8481 -511 8515
rect -477 8481 -443 8515
rect -409 8481 -375 8515
rect -341 8481 -307 8515
rect -273 8481 -266 8515
rect -2966 8446 -266 8481
rect -2966 8412 -2959 8446
rect -2925 8412 -2891 8446
rect -2857 8412 -2823 8446
rect -2789 8412 -2755 8446
rect -2721 8412 -2687 8446
rect -2653 8412 -2619 8446
rect -2585 8412 -2551 8446
rect -2517 8412 -2483 8446
rect -2449 8412 -2415 8446
rect -2381 8412 -2347 8446
rect -2313 8412 -2279 8446
rect -2245 8412 -2211 8446
rect -2177 8412 -2143 8446
rect -2109 8412 -2075 8446
rect -2041 8412 -2007 8446
rect -1973 8412 -1939 8446
rect -1905 8412 -1871 8446
rect -1837 8412 -1803 8446
rect -1769 8412 -1735 8446
rect -1701 8412 -1667 8446
rect -1633 8412 -1599 8446
rect -1565 8412 -1531 8446
rect -1497 8412 -1463 8446
rect -1429 8412 -1395 8446
rect -1361 8412 -1327 8446
rect -1293 8412 -1259 8446
rect -1225 8412 -1191 8446
rect -1157 8412 -1123 8446
rect -1089 8412 -1055 8446
rect -1021 8412 -987 8446
rect -953 8412 -919 8446
rect -885 8412 -851 8446
rect -817 8412 -783 8446
rect -749 8412 -715 8446
rect -681 8412 -647 8446
rect -613 8412 -579 8446
rect -545 8412 -511 8446
rect -477 8412 -443 8446
rect -409 8412 -375 8446
rect -341 8412 -307 8446
rect -273 8412 -266 8446
rect -2966 8377 -266 8412
rect -2966 8343 -2959 8377
rect -2925 8343 -2891 8377
rect -2857 8343 -2823 8377
rect -2789 8343 -2755 8377
rect -2721 8343 -2687 8377
rect -2653 8343 -2619 8377
rect -2585 8343 -2551 8377
rect -2517 8343 -2483 8377
rect -2449 8343 -2415 8377
rect -2381 8343 -2347 8377
rect -2313 8343 -2279 8377
rect -2245 8343 -2211 8377
rect -2177 8343 -2143 8377
rect -2109 8343 -2075 8377
rect -2041 8343 -2007 8377
rect -1973 8343 -1939 8377
rect -1905 8343 -1871 8377
rect -1837 8343 -1803 8377
rect -1769 8343 -1735 8377
rect -1701 8343 -1667 8377
rect -1633 8343 -1599 8377
rect -1565 8343 -1531 8377
rect -1497 8343 -1463 8377
rect -1429 8343 -1395 8377
rect -1361 8343 -1327 8377
rect -1293 8343 -1259 8377
rect -1225 8343 -1191 8377
rect -1157 8343 -1123 8377
rect -1089 8343 -1055 8377
rect -1021 8343 -987 8377
rect -953 8343 -919 8377
rect -885 8343 -851 8377
rect -817 8343 -783 8377
rect -749 8343 -715 8377
rect -681 8343 -647 8377
rect -613 8343 -579 8377
rect -545 8343 -511 8377
rect -477 8343 -443 8377
rect -409 8343 -375 8377
rect -341 8343 -307 8377
rect -273 8343 -266 8377
rect 32028 8355 32061 8542
rect 32028 8348 32085 8355
rect -2966 8308 -266 8343
rect -2966 8274 -2959 8308
rect -2925 8274 -2891 8308
rect -2857 8274 -2823 8308
rect -2789 8274 -2755 8308
rect -2721 8274 -2687 8308
rect -2653 8274 -2619 8308
rect -2585 8274 -2551 8308
rect -2517 8274 -2483 8308
rect -2449 8274 -2415 8308
rect -2381 8274 -2347 8308
rect -2313 8274 -2279 8308
rect -2245 8274 -2211 8308
rect -2177 8274 -2143 8308
rect -2109 8274 -2075 8308
rect -2041 8274 -2007 8308
rect -1973 8274 -1939 8308
rect -1905 8274 -1871 8308
rect -1837 8274 -1803 8308
rect -1769 8274 -1735 8308
rect -1701 8274 -1667 8308
rect -1633 8274 -1599 8308
rect -1565 8274 -1531 8308
rect -1497 8274 -1463 8308
rect -1429 8274 -1395 8308
rect -1361 8274 -1327 8308
rect -1293 8274 -1259 8308
rect -1225 8274 -1191 8308
rect -1157 8274 -1123 8308
rect -1089 8274 -1055 8308
rect -1021 8274 -987 8308
rect -953 8274 -919 8308
rect -885 8274 -851 8308
rect -817 8274 -783 8308
rect -749 8274 -715 8308
rect -681 8274 -647 8308
rect -613 8274 -579 8308
rect -545 8274 -511 8308
rect -477 8274 -443 8308
rect -409 8274 -375 8308
rect -341 8274 -307 8308
rect -273 8274 -266 8308
rect -2966 8239 -266 8274
rect -2966 8205 -2959 8239
rect -2925 8205 -2891 8239
rect -2857 8205 -2823 8239
rect -2789 8205 -2755 8239
rect -2721 8205 -2687 8239
rect -2653 8205 -2619 8239
rect -2585 8205 -2551 8239
rect -2517 8205 -2483 8239
rect -2449 8205 -2415 8239
rect -2381 8205 -2347 8239
rect -2313 8205 -2279 8239
rect -2245 8205 -2211 8239
rect -2177 8205 -2143 8239
rect -2109 8205 -2075 8239
rect -2041 8205 -2007 8239
rect -1973 8205 -1939 8239
rect -1905 8205 -1871 8239
rect -1837 8205 -1803 8239
rect -1769 8205 -1735 8239
rect -1701 8205 -1667 8239
rect -1633 8205 -1599 8239
rect -1565 8205 -1531 8239
rect -1497 8205 -1463 8239
rect -1429 8205 -1395 8239
rect -1361 8205 -1327 8239
rect -1293 8205 -1259 8239
rect -1225 8205 -1191 8239
rect -1157 8205 -1123 8239
rect -1089 8205 -1055 8239
rect -1021 8205 -987 8239
rect -953 8205 -919 8239
rect -885 8205 -851 8239
rect -817 8205 -783 8239
rect -749 8205 -715 8239
rect -681 8205 -647 8239
rect -613 8205 -579 8239
rect -545 8205 -511 8239
rect -477 8205 -443 8239
rect -409 8205 -375 8239
rect -341 8205 -307 8239
rect -273 8205 -266 8239
rect -2966 8170 -266 8205
rect -2966 8136 -2959 8170
rect -2925 8136 -2891 8170
rect -2857 8136 -2823 8170
rect -2789 8136 -2755 8170
rect -2721 8136 -2687 8170
rect -2653 8136 -2619 8170
rect -2585 8136 -2551 8170
rect -2517 8136 -2483 8170
rect -2449 8136 -2415 8170
rect -2381 8136 -2347 8170
rect -2313 8136 -2279 8170
rect -2245 8136 -2211 8170
rect -2177 8136 -2143 8170
rect -2109 8136 -2075 8170
rect -2041 8136 -2007 8170
rect -1973 8136 -1939 8170
rect -1905 8136 -1871 8170
rect -1837 8136 -1803 8170
rect -1769 8136 -1735 8170
rect -1701 8136 -1667 8170
rect -1633 8136 -1599 8170
rect -1565 8136 -1531 8170
rect -1497 8136 -1463 8170
rect -1429 8136 -1395 8170
rect -1361 8136 -1327 8170
rect -1293 8136 -1259 8170
rect -1225 8136 -1191 8170
rect -1157 8136 -1123 8170
rect -1089 8136 -1055 8170
rect -1021 8136 -987 8170
rect -953 8136 -919 8170
rect -885 8136 -851 8170
rect -817 8136 -783 8170
rect -749 8136 -715 8170
rect -681 8136 -647 8170
rect -613 8136 -579 8170
rect -545 8136 -511 8170
rect -477 8136 -443 8170
rect -409 8136 -375 8170
rect -341 8136 -307 8170
rect -273 8136 -266 8170
rect -2966 8101 -266 8136
rect -2966 8067 -2959 8101
rect -2925 8067 -2891 8101
rect -2857 8067 -2823 8101
rect -2789 8067 -2755 8101
rect -2721 8067 -2687 8101
rect -2653 8067 -2619 8101
rect -2585 8067 -2551 8101
rect -2517 8067 -2483 8101
rect -2449 8067 -2415 8101
rect -2381 8067 -2347 8101
rect -2313 8067 -2279 8101
rect -2245 8067 -2211 8101
rect -2177 8067 -2143 8101
rect -2109 8067 -2075 8101
rect -2041 8067 -2007 8101
rect -1973 8067 -1939 8101
rect -1905 8067 -1871 8101
rect -1837 8067 -1803 8101
rect -1769 8067 -1735 8101
rect -1701 8067 -1667 8101
rect -1633 8067 -1599 8101
rect -1565 8067 -1531 8101
rect -1497 8067 -1463 8101
rect -1429 8067 -1395 8101
rect -1361 8067 -1327 8101
rect -1293 8067 -1259 8101
rect -1225 8067 -1191 8101
rect -1157 8067 -1123 8101
rect -1089 8067 -1055 8101
rect -1021 8067 -987 8101
rect -953 8067 -919 8101
rect -885 8067 -851 8101
rect -817 8067 -783 8101
rect -749 8067 -715 8101
rect -681 8067 -647 8101
rect -613 8067 -579 8101
rect -545 8067 -511 8101
rect -477 8067 -443 8101
rect -409 8067 -375 8101
rect -341 8067 -307 8101
rect -273 8067 -266 8101
rect -2966 8032 -266 8067
rect -2966 7998 -2959 8032
rect -2925 7998 -2891 8032
rect -2857 7998 -2823 8032
rect -2789 7998 -2755 8032
rect -2721 7998 -2687 8032
rect -2653 7998 -2619 8032
rect -2585 7998 -2551 8032
rect -2517 7998 -2483 8032
rect -2449 7998 -2415 8032
rect -2381 7998 -2347 8032
rect -2313 7998 -2279 8032
rect -2245 7998 -2211 8032
rect -2177 7998 -2143 8032
rect -2109 7998 -2075 8032
rect -2041 7998 -2007 8032
rect -1973 7998 -1939 8032
rect -1905 7998 -1871 8032
rect -1837 7998 -1803 8032
rect -1769 7998 -1735 8032
rect -1701 7998 -1667 8032
rect -1633 7998 -1599 8032
rect -1565 7998 -1531 8032
rect -1497 7998 -1463 8032
rect -1429 7998 -1395 8032
rect -1361 7998 -1327 8032
rect -1293 7998 -1259 8032
rect -1225 7998 -1191 8032
rect -1157 7998 -1123 8032
rect -1089 7998 -1055 8032
rect -1021 7998 -987 8032
rect -953 7998 -919 8032
rect -885 7998 -851 8032
rect -817 7998 -783 8032
rect -749 7998 -715 8032
rect -681 7998 -647 8032
rect -613 7998 -579 8032
rect -545 7998 -511 8032
rect -477 7998 -443 8032
rect -409 7998 -375 8032
rect -341 7998 -307 8032
rect -273 7998 -266 8032
rect -2966 7963 -266 7998
rect -2966 7929 -2959 7963
rect -2925 7929 -2891 7963
rect -2857 7929 -2823 7963
rect -2789 7929 -2755 7963
rect -2721 7929 -2687 7963
rect -2653 7929 -2619 7963
rect -2585 7929 -2551 7963
rect -2517 7929 -2483 7963
rect -2449 7929 -2415 7963
rect -2381 7929 -2347 7963
rect -2313 7929 -2279 7963
rect -2245 7929 -2211 7963
rect -2177 7929 -2143 7963
rect -2109 7929 -2075 7963
rect -2041 7929 -2007 7963
rect -1973 7929 -1939 7963
rect -1905 7929 -1871 7963
rect -1837 7929 -1803 7963
rect -1769 7929 -1735 7963
rect -1701 7929 -1667 7963
rect -1633 7929 -1599 7963
rect -1565 7929 -1531 7963
rect -1497 7929 -1463 7963
rect -1429 7929 -1395 7963
rect -1361 7929 -1327 7963
rect -1293 7929 -1259 7963
rect -1225 7929 -1191 7963
rect -1157 7929 -1123 7963
rect -1089 7929 -1055 7963
rect -1021 7929 -987 7963
rect -953 7929 -919 7963
rect -885 7929 -851 7963
rect -817 7929 -783 7963
rect -749 7929 -715 7963
rect -681 7929 -647 7963
rect -613 7929 -579 7963
rect -545 7929 -511 7963
rect -477 7929 -443 7963
rect -409 7929 -375 7963
rect -341 7929 -307 7963
rect -273 7929 -266 7963
rect -2966 7894 -266 7929
rect -2966 7860 -2959 7894
rect -2925 7860 -2891 7894
rect -2857 7860 -2823 7894
rect -2789 7860 -2755 7894
rect -2721 7860 -2687 7894
rect -2653 7860 -2619 7894
rect -2585 7860 -2551 7894
rect -2517 7860 -2483 7894
rect -2449 7860 -2415 7894
rect -2381 7860 -2347 7894
rect -2313 7860 -2279 7894
rect -2245 7860 -2211 7894
rect -2177 7860 -2143 7894
rect -2109 7860 -2075 7894
rect -2041 7860 -2007 7894
rect -1973 7860 -1939 7894
rect -1905 7860 -1871 7894
rect -1837 7860 -1803 7894
rect -1769 7860 -1735 7894
rect -1701 7860 -1667 7894
rect -1633 7860 -1599 7894
rect -1565 7860 -1531 7894
rect -1497 7860 -1463 7894
rect -1429 7860 -1395 7894
rect -1361 7860 -1327 7894
rect -1293 7860 -1259 7894
rect -1225 7860 -1191 7894
rect -1157 7860 -1123 7894
rect -1089 7860 -1055 7894
rect -1021 7860 -987 7894
rect -953 7860 -919 7894
rect -885 7860 -851 7894
rect -817 7860 -783 7894
rect -749 7860 -715 7894
rect -681 7860 -647 7894
rect -613 7860 -579 7894
rect -545 7860 -511 7894
rect -477 7860 -443 7894
rect -409 7860 -375 7894
rect -341 7860 -307 7894
rect -273 7860 -266 7894
rect -2966 7825 -266 7860
rect -2966 7791 -2959 7825
rect -2925 7791 -2891 7825
rect -2857 7791 -2823 7825
rect -2789 7791 -2755 7825
rect -2721 7791 -2687 7825
rect -2653 7791 -2619 7825
rect -2585 7791 -2551 7825
rect -2517 7791 -2483 7825
rect -2449 7791 -2415 7825
rect -2381 7791 -2347 7825
rect -2313 7791 -2279 7825
rect -2245 7791 -2211 7825
rect -2177 7791 -2143 7825
rect -2109 7791 -2075 7825
rect -2041 7791 -2007 7825
rect -1973 7791 -1939 7825
rect -1905 7791 -1871 7825
rect -1837 7791 -1803 7825
rect -1769 7791 -1735 7825
rect -1701 7791 -1667 7825
rect -1633 7791 -1599 7825
rect -1565 7791 -1531 7825
rect -1497 7791 -1463 7825
rect -1429 7791 -1395 7825
rect -1361 7791 -1327 7825
rect -1293 7791 -1259 7825
rect -1225 7791 -1191 7825
rect -1157 7791 -1123 7825
rect -1089 7791 -1055 7825
rect -1021 7791 -987 7825
rect -953 7791 -919 7825
rect -885 7791 -851 7825
rect -817 7791 -783 7825
rect -749 7791 -715 7825
rect -681 7791 -647 7825
rect -613 7791 -579 7825
rect -545 7791 -511 7825
rect -477 7791 -443 7825
rect -409 7791 -375 7825
rect -341 7791 -307 7825
rect -273 7791 -266 7825
rect -2966 7756 -266 7791
rect -2966 7722 -2959 7756
rect -2925 7722 -2891 7756
rect -2857 7722 -2823 7756
rect -2789 7722 -2755 7756
rect -2721 7722 -2687 7756
rect -2653 7722 -2619 7756
rect -2585 7722 -2551 7756
rect -2517 7722 -2483 7756
rect -2449 7722 -2415 7756
rect -2381 7722 -2347 7756
rect -2313 7722 -2279 7756
rect -2245 7722 -2211 7756
rect -2177 7722 -2143 7756
rect -2109 7722 -2075 7756
rect -2041 7722 -2007 7756
rect -1973 7722 -1939 7756
rect -1905 7722 -1871 7756
rect -1837 7722 -1803 7756
rect -1769 7722 -1735 7756
rect -1701 7722 -1667 7756
rect -1633 7722 -1599 7756
rect -1565 7722 -1531 7756
rect -1497 7722 -1463 7756
rect -1429 7722 -1395 7756
rect -1361 7722 -1327 7756
rect -1293 7722 -1259 7756
rect -1225 7722 -1191 7756
rect -1157 7722 -1123 7756
rect -1089 7722 -1055 7756
rect -1021 7722 -987 7756
rect -953 7722 -919 7756
rect -885 7722 -851 7756
rect -817 7722 -783 7756
rect -749 7722 -715 7756
rect -681 7722 -647 7756
rect -613 7722 -579 7756
rect -545 7722 -511 7756
rect -477 7722 -443 7756
rect -409 7722 -375 7756
rect -341 7722 -307 7756
rect -273 7722 -266 7756
rect -2966 7687 -266 7722
rect -2966 7653 -2959 7687
rect -2925 7653 -2891 7687
rect -2857 7653 -2823 7687
rect -2789 7653 -2755 7687
rect -2721 7653 -2687 7687
rect -2653 7653 -2619 7687
rect -2585 7653 -2551 7687
rect -2517 7653 -2483 7687
rect -2449 7653 -2415 7687
rect -2381 7653 -2347 7687
rect -2313 7653 -2279 7687
rect -2245 7653 -2211 7687
rect -2177 7653 -2143 7687
rect -2109 7653 -2075 7687
rect -2041 7653 -2007 7687
rect -1973 7653 -1939 7687
rect -1905 7653 -1871 7687
rect -1837 7653 -1803 7687
rect -1769 7653 -1735 7687
rect -1701 7653 -1667 7687
rect -1633 7653 -1599 7687
rect -1565 7653 -1531 7687
rect -1497 7653 -1463 7687
rect -1429 7653 -1395 7687
rect -1361 7653 -1327 7687
rect -1293 7653 -1259 7687
rect -1225 7653 -1191 7687
rect -1157 7653 -1123 7687
rect -1089 7653 -1055 7687
rect -1021 7653 -987 7687
rect -953 7653 -919 7687
rect -885 7653 -851 7687
rect -817 7653 -783 7687
rect -749 7653 -715 7687
rect -681 7653 -647 7687
rect -613 7653 -579 7687
rect -545 7653 -511 7687
rect -477 7653 -443 7687
rect -409 7653 -375 7687
rect -341 7653 -307 7687
rect -273 7653 -266 7687
rect -2966 7618 -266 7653
rect -2966 7584 -2959 7618
rect -2925 7584 -2891 7618
rect -2857 7584 -2823 7618
rect -2789 7584 -2755 7618
rect -2721 7584 -2687 7618
rect -2653 7584 -2619 7618
rect -2585 7584 -2551 7618
rect -2517 7584 -2483 7618
rect -2449 7584 -2415 7618
rect -2381 7584 -2347 7618
rect -2313 7584 -2279 7618
rect -2245 7584 -2211 7618
rect -2177 7584 -2143 7618
rect -2109 7584 -2075 7618
rect -2041 7584 -2007 7618
rect -1973 7584 -1939 7618
rect -1905 7584 -1871 7618
rect -1837 7584 -1803 7618
rect -1769 7584 -1735 7618
rect -1701 7584 -1667 7618
rect -1633 7584 -1599 7618
rect -1565 7584 -1531 7618
rect -1497 7584 -1463 7618
rect -1429 7584 -1395 7618
rect -1361 7584 -1327 7618
rect -1293 7584 -1259 7618
rect -1225 7584 -1191 7618
rect -1157 7584 -1123 7618
rect -1089 7584 -1055 7618
rect -1021 7584 -987 7618
rect -953 7584 -919 7618
rect -885 7584 -851 7618
rect -817 7584 -783 7618
rect -749 7584 -715 7618
rect -681 7584 -647 7618
rect -613 7584 -579 7618
rect -545 7584 -511 7618
rect -477 7584 -443 7618
rect -409 7584 -375 7618
rect -341 7584 -307 7618
rect -273 7584 -266 7618
rect -2966 7549 -266 7584
rect -2966 7515 -2959 7549
rect -2925 7515 -2891 7549
rect -2857 7515 -2823 7549
rect -2789 7515 -2755 7549
rect -2721 7515 -2687 7549
rect -2653 7515 -2619 7549
rect -2585 7515 -2551 7549
rect -2517 7515 -2483 7549
rect -2449 7515 -2415 7549
rect -2381 7515 -2347 7549
rect -2313 7515 -2279 7549
rect -2245 7515 -2211 7549
rect -2177 7515 -2143 7549
rect -2109 7515 -2075 7549
rect -2041 7515 -2007 7549
rect -1973 7515 -1939 7549
rect -1905 7515 -1871 7549
rect -1837 7515 -1803 7549
rect -1769 7515 -1735 7549
rect -1701 7515 -1667 7549
rect -1633 7515 -1599 7549
rect -1565 7515 -1531 7549
rect -1497 7515 -1463 7549
rect -1429 7515 -1395 7549
rect -1361 7515 -1327 7549
rect -1293 7515 -1259 7549
rect -1225 7515 -1191 7549
rect -1157 7515 -1123 7549
rect -1089 7515 -1055 7549
rect -1021 7515 -987 7549
rect -953 7515 -919 7549
rect -885 7515 -851 7549
rect -817 7515 -783 7549
rect -749 7515 -715 7549
rect -681 7515 -647 7549
rect -613 7515 -579 7549
rect -545 7515 -511 7549
rect -477 7515 -443 7549
rect -409 7515 -375 7549
rect -341 7515 -307 7549
rect -273 7515 -266 7549
rect -2966 7480 -266 7515
rect -2966 7446 -2959 7480
rect -2925 7446 -2891 7480
rect -2857 7446 -2823 7480
rect -2789 7446 -2755 7480
rect -2721 7446 -2687 7480
rect -2653 7446 -2619 7480
rect -2585 7446 -2551 7480
rect -2517 7446 -2483 7480
rect -2449 7446 -2415 7480
rect -2381 7446 -2347 7480
rect -2313 7446 -2279 7480
rect -2245 7446 -2211 7480
rect -2177 7446 -2143 7480
rect -2109 7446 -2075 7480
rect -2041 7446 -2007 7480
rect -1973 7446 -1939 7480
rect -1905 7446 -1871 7480
rect -1837 7446 -1803 7480
rect -1769 7446 -1735 7480
rect -1701 7446 -1667 7480
rect -1633 7446 -1599 7480
rect -1565 7446 -1531 7480
rect -1497 7446 -1463 7480
rect -1429 7446 -1395 7480
rect -1361 7446 -1327 7480
rect -1293 7446 -1259 7480
rect -1225 7446 -1191 7480
rect -1157 7446 -1123 7480
rect -1089 7446 -1055 7480
rect -1021 7446 -987 7480
rect -953 7446 -919 7480
rect -885 7446 -851 7480
rect -817 7446 -783 7480
rect -749 7446 -715 7480
rect -681 7446 -647 7480
rect -613 7446 -579 7480
rect -545 7446 -511 7480
rect -477 7446 -443 7480
rect -409 7446 -375 7480
rect -341 7446 -307 7480
rect -273 7446 -266 7480
rect -2966 7422 -266 7446
rect 6294 4588 6334 4617
rect 6243 3827 6319 4230
rect 6243 3771 6641 3827
rect 6243 3732 6319 3771
<< viali >>
rect -2829 37942 -275 50607
rect -2829 37907 -275 37942
rect -2829 37901 -2802 37907
rect -2802 37901 -2768 37907
rect -2768 37901 -2734 37907
rect -2734 37901 -2700 37907
rect -2700 37901 -2666 37907
rect -2666 37901 -2632 37907
rect -2632 37901 -2598 37907
rect -2598 37901 -2564 37907
rect -2564 37901 -2530 37907
rect -2530 37901 -2496 37907
rect -2496 37901 -2462 37907
rect -2462 37901 -2428 37907
rect -2428 37901 -2394 37907
rect -2394 37901 -2360 37907
rect -2360 37901 -2326 37907
rect -2326 37901 -2292 37907
rect -2292 37901 -2258 37907
rect -2258 37901 -2224 37907
rect -2224 37901 -2190 37907
rect -2190 37901 -2156 37907
rect -2156 37901 -2122 37907
rect -2122 37901 -2088 37907
rect -2088 37901 -2054 37907
rect -2054 37901 -2020 37907
rect -2020 37901 -1986 37907
rect -1986 37901 -1952 37907
rect -1952 37901 -1918 37907
rect -1918 37901 -1884 37907
rect -1884 37901 -1850 37907
rect -1850 37901 -1816 37907
rect -1816 37901 -1782 37907
rect -1782 37901 -1748 37907
rect -1748 37901 -1714 37907
rect -1714 37901 -1680 37907
rect -1680 37901 -1646 37907
rect -1646 37901 -1612 37907
rect -1612 37901 -1578 37907
rect -1578 37901 -1544 37907
rect -1544 37901 -1510 37907
rect -1510 37901 -1476 37907
rect -1476 37901 -1442 37907
rect -1442 37901 -1408 37907
rect -1408 37901 -1374 37907
rect -1374 37901 -1340 37907
rect -1340 37901 -1306 37907
rect -1306 37901 -1272 37907
rect -1272 37901 -1238 37907
rect -1238 37901 -1204 37907
rect -1204 37901 -1170 37907
rect -1170 37901 -1136 37907
rect -1136 37901 -1102 37907
rect -1102 37901 -1068 37907
rect -1068 37901 -1034 37907
rect -1034 37901 -1000 37907
rect -1000 37901 -966 37907
rect -966 37901 -932 37907
rect -932 37901 -898 37907
rect -898 37901 -864 37907
rect -864 37901 -830 37907
rect -830 37901 -796 37907
rect -796 37901 -762 37907
rect -762 37901 -728 37907
rect -728 37901 -694 37907
rect -694 37901 -660 37907
rect -660 37901 -626 37907
rect -626 37901 -592 37907
rect -592 37901 -558 37907
rect -558 37901 -524 37907
rect -524 37901 -490 37907
rect -490 37901 -456 37907
rect -456 37901 -422 37907
rect -422 37901 -388 37907
rect -388 37901 -354 37907
rect -354 37901 -320 37907
rect -320 37901 -286 37907
rect -286 37901 -275 37907
rect -2829 37838 -2795 37862
rect -2757 37838 -2723 37862
rect -2685 37838 -2651 37862
rect -2613 37838 -2579 37862
rect -2541 37838 -2507 37862
rect -2469 37838 -2435 37862
rect -2397 37838 -2363 37862
rect -2325 37838 -2291 37862
rect -2253 37838 -2219 37862
rect -2181 37838 -2147 37862
rect -2109 37838 -2075 37862
rect -2037 37838 -2003 37862
rect -1965 37838 -1931 37862
rect -1893 37838 -1859 37862
rect -1821 37838 -1787 37862
rect -1749 37838 -1715 37862
rect -1677 37838 -1643 37862
rect -1605 37838 -1571 37862
rect -1533 37838 -1499 37862
rect -1461 37838 -1427 37862
rect -1389 37838 -1355 37862
rect -1317 37838 -1283 37862
rect -1245 37838 -1211 37862
rect -1173 37838 -1139 37862
rect -1101 37838 -1067 37862
rect -1029 37838 -995 37862
rect -957 37838 -923 37862
rect -885 37838 -851 37862
rect -813 37838 -779 37862
rect -741 37838 -707 37862
rect -669 37838 -635 37862
rect -597 37838 -563 37862
rect -525 37838 -491 37862
rect -453 37838 -419 37862
rect -381 37838 -347 37862
rect -309 37838 -275 37862
rect -2829 37828 -2802 37838
rect -2802 37828 -2795 37838
rect -2757 37828 -2734 37838
rect -2734 37828 -2723 37838
rect -2685 37828 -2666 37838
rect -2666 37828 -2651 37838
rect -2613 37828 -2598 37838
rect -2598 37828 -2579 37838
rect -2541 37828 -2530 37838
rect -2530 37828 -2507 37838
rect -2469 37828 -2462 37838
rect -2462 37828 -2435 37838
rect -2397 37828 -2394 37838
rect -2394 37828 -2363 37838
rect -2325 37828 -2292 37838
rect -2292 37828 -2291 37838
rect -2253 37828 -2224 37838
rect -2224 37828 -2219 37838
rect -2181 37828 -2156 37838
rect -2156 37828 -2147 37838
rect -2109 37828 -2088 37838
rect -2088 37828 -2075 37838
rect -2037 37828 -2020 37838
rect -2020 37828 -2003 37838
rect -1965 37828 -1952 37838
rect -1952 37828 -1931 37838
rect -1893 37828 -1884 37838
rect -1884 37828 -1859 37838
rect -1821 37828 -1816 37838
rect -1816 37828 -1787 37838
rect -1749 37828 -1748 37838
rect -1748 37828 -1715 37838
rect -1677 37828 -1646 37838
rect -1646 37828 -1643 37838
rect -1605 37828 -1578 37838
rect -1578 37828 -1571 37838
rect -1533 37828 -1510 37838
rect -1510 37828 -1499 37838
rect -1461 37828 -1442 37838
rect -1442 37828 -1427 37838
rect -1389 37828 -1374 37838
rect -1374 37828 -1355 37838
rect -1317 37828 -1306 37838
rect -1306 37828 -1283 37838
rect -1245 37828 -1238 37838
rect -1238 37828 -1211 37838
rect -1173 37828 -1170 37838
rect -1170 37828 -1139 37838
rect -1101 37828 -1068 37838
rect -1068 37828 -1067 37838
rect -1029 37828 -1000 37838
rect -1000 37828 -995 37838
rect -957 37828 -932 37838
rect -932 37828 -923 37838
rect -885 37828 -864 37838
rect -864 37828 -851 37838
rect -813 37828 -796 37838
rect -796 37828 -779 37838
rect -741 37828 -728 37838
rect -728 37828 -707 37838
rect -669 37828 -660 37838
rect -660 37828 -635 37838
rect -597 37828 -592 37838
rect -592 37828 -563 37838
rect -525 37828 -524 37838
rect -524 37828 -491 37838
rect -453 37828 -422 37838
rect -422 37828 -419 37838
rect -381 37828 -354 37838
rect -354 37828 -347 37838
rect -309 37828 -286 37838
rect -286 37828 -275 37838
rect -2829 37769 -2795 37789
rect -2757 37769 -2723 37789
rect -2685 37769 -2651 37789
rect -2613 37769 -2579 37789
rect -2541 37769 -2507 37789
rect -2469 37769 -2435 37789
rect -2397 37769 -2363 37789
rect -2325 37769 -2291 37789
rect -2253 37769 -2219 37789
rect -2181 37769 -2147 37789
rect -2109 37769 -2075 37789
rect -2037 37769 -2003 37789
rect -1965 37769 -1931 37789
rect -1893 37769 -1859 37789
rect -1821 37769 -1787 37789
rect -1749 37769 -1715 37789
rect -1677 37769 -1643 37789
rect -1605 37769 -1571 37789
rect -1533 37769 -1499 37789
rect -1461 37769 -1427 37789
rect -1389 37769 -1355 37789
rect -1317 37769 -1283 37789
rect -1245 37769 -1211 37789
rect -1173 37769 -1139 37789
rect -1101 37769 -1067 37789
rect -1029 37769 -995 37789
rect -957 37769 -923 37789
rect -885 37769 -851 37789
rect -813 37769 -779 37789
rect -741 37769 -707 37789
rect -669 37769 -635 37789
rect -597 37769 -563 37789
rect -525 37769 -491 37789
rect -453 37769 -419 37789
rect -381 37769 -347 37789
rect -309 37769 -275 37789
rect -2829 37755 -2802 37769
rect -2802 37755 -2795 37769
rect -2757 37755 -2734 37769
rect -2734 37755 -2723 37769
rect -2685 37755 -2666 37769
rect -2666 37755 -2651 37769
rect -2613 37755 -2598 37769
rect -2598 37755 -2579 37769
rect -2541 37755 -2530 37769
rect -2530 37755 -2507 37769
rect -2469 37755 -2462 37769
rect -2462 37755 -2435 37769
rect -2397 37755 -2394 37769
rect -2394 37755 -2363 37769
rect -2325 37755 -2292 37769
rect -2292 37755 -2291 37769
rect -2253 37755 -2224 37769
rect -2224 37755 -2219 37769
rect -2181 37755 -2156 37769
rect -2156 37755 -2147 37769
rect -2109 37755 -2088 37769
rect -2088 37755 -2075 37769
rect -2037 37755 -2020 37769
rect -2020 37755 -2003 37769
rect -1965 37755 -1952 37769
rect -1952 37755 -1931 37769
rect -1893 37755 -1884 37769
rect -1884 37755 -1859 37769
rect -1821 37755 -1816 37769
rect -1816 37755 -1787 37769
rect -1749 37755 -1748 37769
rect -1748 37755 -1715 37769
rect -1677 37755 -1646 37769
rect -1646 37755 -1643 37769
rect -1605 37755 -1578 37769
rect -1578 37755 -1571 37769
rect -1533 37755 -1510 37769
rect -1510 37755 -1499 37769
rect -1461 37755 -1442 37769
rect -1442 37755 -1427 37769
rect -1389 37755 -1374 37769
rect -1374 37755 -1355 37769
rect -1317 37755 -1306 37769
rect -1306 37755 -1283 37769
rect -1245 37755 -1238 37769
rect -1238 37755 -1211 37769
rect -1173 37755 -1170 37769
rect -1170 37755 -1139 37769
rect -1101 37755 -1068 37769
rect -1068 37755 -1067 37769
rect -1029 37755 -1000 37769
rect -1000 37755 -995 37769
rect -957 37755 -932 37769
rect -932 37755 -923 37769
rect -885 37755 -864 37769
rect -864 37755 -851 37769
rect -813 37755 -796 37769
rect -796 37755 -779 37769
rect -741 37755 -728 37769
rect -728 37755 -707 37769
rect -669 37755 -660 37769
rect -660 37755 -635 37769
rect -597 37755 -592 37769
rect -592 37755 -563 37769
rect -525 37755 -524 37769
rect -524 37755 -491 37769
rect -453 37755 -422 37769
rect -422 37755 -419 37769
rect -381 37755 -354 37769
rect -354 37755 -347 37769
rect -309 37755 -286 37769
rect -286 37755 -275 37769
rect -2829 37700 -2795 37716
rect -2757 37700 -2723 37716
rect -2685 37700 -2651 37716
rect -2613 37700 -2579 37716
rect -2541 37700 -2507 37716
rect -2469 37700 -2435 37716
rect -2397 37700 -2363 37716
rect -2325 37700 -2291 37716
rect -2253 37700 -2219 37716
rect -2181 37700 -2147 37716
rect -2109 37700 -2075 37716
rect -2037 37700 -2003 37716
rect -1965 37700 -1931 37716
rect -1893 37700 -1859 37716
rect -1821 37700 -1787 37716
rect -1749 37700 -1715 37716
rect -1677 37700 -1643 37716
rect -1605 37700 -1571 37716
rect -1533 37700 -1499 37716
rect -1461 37700 -1427 37716
rect -1389 37700 -1355 37716
rect -1317 37700 -1283 37716
rect -1245 37700 -1211 37716
rect -1173 37700 -1139 37716
rect -1101 37700 -1067 37716
rect -1029 37700 -995 37716
rect -957 37700 -923 37716
rect -885 37700 -851 37716
rect -813 37700 -779 37716
rect -741 37700 -707 37716
rect -669 37700 -635 37716
rect -597 37700 -563 37716
rect -525 37700 -491 37716
rect -453 37700 -419 37716
rect -381 37700 -347 37716
rect -309 37700 -275 37716
rect -2829 37682 -2802 37700
rect -2802 37682 -2795 37700
rect -2757 37682 -2734 37700
rect -2734 37682 -2723 37700
rect -2685 37682 -2666 37700
rect -2666 37682 -2651 37700
rect -2613 37682 -2598 37700
rect -2598 37682 -2579 37700
rect -2541 37682 -2530 37700
rect -2530 37682 -2507 37700
rect -2469 37682 -2462 37700
rect -2462 37682 -2435 37700
rect -2397 37682 -2394 37700
rect -2394 37682 -2363 37700
rect -2325 37682 -2292 37700
rect -2292 37682 -2291 37700
rect -2253 37682 -2224 37700
rect -2224 37682 -2219 37700
rect -2181 37682 -2156 37700
rect -2156 37682 -2147 37700
rect -2109 37682 -2088 37700
rect -2088 37682 -2075 37700
rect -2037 37682 -2020 37700
rect -2020 37682 -2003 37700
rect -1965 37682 -1952 37700
rect -1952 37682 -1931 37700
rect -1893 37682 -1884 37700
rect -1884 37682 -1859 37700
rect -1821 37682 -1816 37700
rect -1816 37682 -1787 37700
rect -1749 37682 -1748 37700
rect -1748 37682 -1715 37700
rect -1677 37682 -1646 37700
rect -1646 37682 -1643 37700
rect -1605 37682 -1578 37700
rect -1578 37682 -1571 37700
rect -1533 37682 -1510 37700
rect -1510 37682 -1499 37700
rect -1461 37682 -1442 37700
rect -1442 37682 -1427 37700
rect -1389 37682 -1374 37700
rect -1374 37682 -1355 37700
rect -1317 37682 -1306 37700
rect -1306 37682 -1283 37700
rect -1245 37682 -1238 37700
rect -1238 37682 -1211 37700
rect -1173 37682 -1170 37700
rect -1170 37682 -1139 37700
rect -1101 37682 -1068 37700
rect -1068 37682 -1067 37700
rect -1029 37682 -1000 37700
rect -1000 37682 -995 37700
rect -957 37682 -932 37700
rect -932 37682 -923 37700
rect -885 37682 -864 37700
rect -864 37682 -851 37700
rect -813 37682 -796 37700
rect -796 37682 -779 37700
rect -741 37682 -728 37700
rect -728 37682 -707 37700
rect -669 37682 -660 37700
rect -660 37682 -635 37700
rect -597 37682 -592 37700
rect -592 37682 -563 37700
rect -525 37682 -524 37700
rect -524 37682 -491 37700
rect -453 37682 -422 37700
rect -422 37682 -419 37700
rect -381 37682 -354 37700
rect -354 37682 -347 37700
rect -309 37682 -286 37700
rect -286 37682 -275 37700
rect -2829 37631 -2795 37643
rect -2757 37631 -2723 37643
rect -2685 37631 -2651 37643
rect -2613 37631 -2579 37643
rect -2541 37631 -2507 37643
rect -2469 37631 -2435 37643
rect -2397 37631 -2363 37643
rect -2325 37631 -2291 37643
rect -2253 37631 -2219 37643
rect -2181 37631 -2147 37643
rect -2109 37631 -2075 37643
rect -2037 37631 -2003 37643
rect -1965 37631 -1931 37643
rect -1893 37631 -1859 37643
rect -1821 37631 -1787 37643
rect -1749 37631 -1715 37643
rect -1677 37631 -1643 37643
rect -1605 37631 -1571 37643
rect -1533 37631 -1499 37643
rect -1461 37631 -1427 37643
rect -1389 37631 -1355 37643
rect -1317 37631 -1283 37643
rect -1245 37631 -1211 37643
rect -1173 37631 -1139 37643
rect -1101 37631 -1067 37643
rect -1029 37631 -995 37643
rect -957 37631 -923 37643
rect -885 37631 -851 37643
rect -813 37631 -779 37643
rect -741 37631 -707 37643
rect -669 37631 -635 37643
rect -597 37631 -563 37643
rect -525 37631 -491 37643
rect -453 37631 -419 37643
rect -381 37631 -347 37643
rect -309 37631 -275 37643
rect -2829 37609 -2802 37631
rect -2802 37609 -2795 37631
rect -2757 37609 -2734 37631
rect -2734 37609 -2723 37631
rect -2685 37609 -2666 37631
rect -2666 37609 -2651 37631
rect -2613 37609 -2598 37631
rect -2598 37609 -2579 37631
rect -2541 37609 -2530 37631
rect -2530 37609 -2507 37631
rect -2469 37609 -2462 37631
rect -2462 37609 -2435 37631
rect -2397 37609 -2394 37631
rect -2394 37609 -2363 37631
rect -2325 37609 -2292 37631
rect -2292 37609 -2291 37631
rect -2253 37609 -2224 37631
rect -2224 37609 -2219 37631
rect -2181 37609 -2156 37631
rect -2156 37609 -2147 37631
rect -2109 37609 -2088 37631
rect -2088 37609 -2075 37631
rect -2037 37609 -2020 37631
rect -2020 37609 -2003 37631
rect -1965 37609 -1952 37631
rect -1952 37609 -1931 37631
rect -1893 37609 -1884 37631
rect -1884 37609 -1859 37631
rect -1821 37609 -1816 37631
rect -1816 37609 -1787 37631
rect -1749 37609 -1748 37631
rect -1748 37609 -1715 37631
rect -1677 37609 -1646 37631
rect -1646 37609 -1643 37631
rect -1605 37609 -1578 37631
rect -1578 37609 -1571 37631
rect -1533 37609 -1510 37631
rect -1510 37609 -1499 37631
rect -1461 37609 -1442 37631
rect -1442 37609 -1427 37631
rect -1389 37609 -1374 37631
rect -1374 37609 -1355 37631
rect -1317 37609 -1306 37631
rect -1306 37609 -1283 37631
rect -1245 37609 -1238 37631
rect -1238 37609 -1211 37631
rect -1173 37609 -1170 37631
rect -1170 37609 -1139 37631
rect -1101 37609 -1068 37631
rect -1068 37609 -1067 37631
rect -1029 37609 -1000 37631
rect -1000 37609 -995 37631
rect -957 37609 -932 37631
rect -932 37609 -923 37631
rect -885 37609 -864 37631
rect -864 37609 -851 37631
rect -813 37609 -796 37631
rect -796 37609 -779 37631
rect -741 37609 -728 37631
rect -728 37609 -707 37631
rect -669 37609 -660 37631
rect -660 37609 -635 37631
rect -597 37609 -592 37631
rect -592 37609 -563 37631
rect -525 37609 -524 37631
rect -524 37609 -491 37631
rect -453 37609 -422 37631
rect -422 37609 -419 37631
rect -381 37609 -354 37631
rect -354 37609 -347 37631
rect -309 37609 -286 37631
rect -286 37609 -275 37631
rect -2829 37562 -2795 37570
rect -2757 37562 -2723 37570
rect -2685 37562 -2651 37570
rect -2613 37562 -2579 37570
rect -2541 37562 -2507 37570
rect -2469 37562 -2435 37570
rect -2397 37562 -2363 37570
rect -2325 37562 -2291 37570
rect -2253 37562 -2219 37570
rect -2181 37562 -2147 37570
rect -2109 37562 -2075 37570
rect -2037 37562 -2003 37570
rect -1965 37562 -1931 37570
rect -1893 37562 -1859 37570
rect -1821 37562 -1787 37570
rect -1749 37562 -1715 37570
rect -1677 37562 -1643 37570
rect -1605 37562 -1571 37570
rect -1533 37562 -1499 37570
rect -1461 37562 -1427 37570
rect -1389 37562 -1355 37570
rect -1317 37562 -1283 37570
rect -1245 37562 -1211 37570
rect -1173 37562 -1139 37570
rect -1101 37562 -1067 37570
rect -1029 37562 -995 37570
rect -957 37562 -923 37570
rect -885 37562 -851 37570
rect -813 37562 -779 37570
rect -741 37562 -707 37570
rect -669 37562 -635 37570
rect -597 37562 -563 37570
rect -525 37562 -491 37570
rect -453 37562 -419 37570
rect -381 37562 -347 37570
rect -309 37562 -275 37570
rect -2829 37536 -2802 37562
rect -2802 37536 -2795 37562
rect -2757 37536 -2734 37562
rect -2734 37536 -2723 37562
rect -2685 37536 -2666 37562
rect -2666 37536 -2651 37562
rect -2613 37536 -2598 37562
rect -2598 37536 -2579 37562
rect -2541 37536 -2530 37562
rect -2530 37536 -2507 37562
rect -2469 37536 -2462 37562
rect -2462 37536 -2435 37562
rect -2397 37536 -2394 37562
rect -2394 37536 -2363 37562
rect -2325 37536 -2292 37562
rect -2292 37536 -2291 37562
rect -2253 37536 -2224 37562
rect -2224 37536 -2219 37562
rect -2181 37536 -2156 37562
rect -2156 37536 -2147 37562
rect -2109 37536 -2088 37562
rect -2088 37536 -2075 37562
rect -2037 37536 -2020 37562
rect -2020 37536 -2003 37562
rect -1965 37536 -1952 37562
rect -1952 37536 -1931 37562
rect -1893 37536 -1884 37562
rect -1884 37536 -1859 37562
rect -1821 37536 -1816 37562
rect -1816 37536 -1787 37562
rect -1749 37536 -1748 37562
rect -1748 37536 -1715 37562
rect -1677 37536 -1646 37562
rect -1646 37536 -1643 37562
rect -1605 37536 -1578 37562
rect -1578 37536 -1571 37562
rect -1533 37536 -1510 37562
rect -1510 37536 -1499 37562
rect -1461 37536 -1442 37562
rect -1442 37536 -1427 37562
rect -1389 37536 -1374 37562
rect -1374 37536 -1355 37562
rect -1317 37536 -1306 37562
rect -1306 37536 -1283 37562
rect -1245 37536 -1238 37562
rect -1238 37536 -1211 37562
rect -1173 37536 -1170 37562
rect -1170 37536 -1139 37562
rect -1101 37536 -1068 37562
rect -1068 37536 -1067 37562
rect -1029 37536 -1000 37562
rect -1000 37536 -995 37562
rect -957 37536 -932 37562
rect -932 37536 -923 37562
rect -885 37536 -864 37562
rect -864 37536 -851 37562
rect -813 37536 -796 37562
rect -796 37536 -779 37562
rect -741 37536 -728 37562
rect -728 37536 -707 37562
rect -669 37536 -660 37562
rect -660 37536 -635 37562
rect -597 37536 -592 37562
rect -592 37536 -563 37562
rect -525 37536 -524 37562
rect -524 37536 -491 37562
rect -453 37536 -422 37562
rect -422 37536 -419 37562
rect -381 37536 -354 37562
rect -354 37536 -347 37562
rect -309 37536 -286 37562
rect -286 37536 -275 37562
rect -2829 37493 -2795 37497
rect -2757 37493 -2723 37497
rect -2685 37493 -2651 37497
rect -2613 37493 -2579 37497
rect -2541 37493 -2507 37497
rect -2469 37493 -2435 37497
rect -2397 37493 -2363 37497
rect -2325 37493 -2291 37497
rect -2253 37493 -2219 37497
rect -2181 37493 -2147 37497
rect -2109 37493 -2075 37497
rect -2037 37493 -2003 37497
rect -1965 37493 -1931 37497
rect -1893 37493 -1859 37497
rect -1821 37493 -1787 37497
rect -1749 37493 -1715 37497
rect -1677 37493 -1643 37497
rect -1605 37493 -1571 37497
rect -1533 37493 -1499 37497
rect -1461 37493 -1427 37497
rect -1389 37493 -1355 37497
rect -1317 37493 -1283 37497
rect -1245 37493 -1211 37497
rect -1173 37493 -1139 37497
rect -1101 37493 -1067 37497
rect -1029 37493 -995 37497
rect -957 37493 -923 37497
rect -885 37493 -851 37497
rect -813 37493 -779 37497
rect -741 37493 -707 37497
rect -669 37493 -635 37497
rect -597 37493 -563 37497
rect -525 37493 -491 37497
rect -453 37493 -419 37497
rect -381 37493 -347 37497
rect -309 37493 -275 37497
rect -2829 37463 -2802 37493
rect -2802 37463 -2795 37493
rect -2757 37463 -2734 37493
rect -2734 37463 -2723 37493
rect -2685 37463 -2666 37493
rect -2666 37463 -2651 37493
rect -2613 37463 -2598 37493
rect -2598 37463 -2579 37493
rect -2541 37463 -2530 37493
rect -2530 37463 -2507 37493
rect -2469 37463 -2462 37493
rect -2462 37463 -2435 37493
rect -2397 37463 -2394 37493
rect -2394 37463 -2363 37493
rect -2325 37463 -2292 37493
rect -2292 37463 -2291 37493
rect -2253 37463 -2224 37493
rect -2224 37463 -2219 37493
rect -2181 37463 -2156 37493
rect -2156 37463 -2147 37493
rect -2109 37463 -2088 37493
rect -2088 37463 -2075 37493
rect -2037 37463 -2020 37493
rect -2020 37463 -2003 37493
rect -1965 37463 -1952 37493
rect -1952 37463 -1931 37493
rect -1893 37463 -1884 37493
rect -1884 37463 -1859 37493
rect -1821 37463 -1816 37493
rect -1816 37463 -1787 37493
rect -1749 37463 -1748 37493
rect -1748 37463 -1715 37493
rect -1677 37463 -1646 37493
rect -1646 37463 -1643 37493
rect -1605 37463 -1578 37493
rect -1578 37463 -1571 37493
rect -1533 37463 -1510 37493
rect -1510 37463 -1499 37493
rect -1461 37463 -1442 37493
rect -1442 37463 -1427 37493
rect -1389 37463 -1374 37493
rect -1374 37463 -1355 37493
rect -1317 37463 -1306 37493
rect -1306 37463 -1283 37493
rect -1245 37463 -1238 37493
rect -1238 37463 -1211 37493
rect -1173 37463 -1170 37493
rect -1170 37463 -1139 37493
rect -1101 37463 -1068 37493
rect -1068 37463 -1067 37493
rect -1029 37463 -1000 37493
rect -1000 37463 -995 37493
rect -957 37463 -932 37493
rect -932 37463 -923 37493
rect -885 37463 -864 37493
rect -864 37463 -851 37493
rect -813 37463 -796 37493
rect -796 37463 -779 37493
rect -741 37463 -728 37493
rect -728 37463 -707 37493
rect -669 37463 -660 37493
rect -660 37463 -635 37493
rect -597 37463 -592 37493
rect -592 37463 -563 37493
rect -525 37463 -524 37493
rect -524 37463 -491 37493
rect -453 37463 -422 37493
rect -422 37463 -419 37493
rect -381 37463 -354 37493
rect -354 37463 -347 37493
rect -309 37463 -286 37493
rect -286 37463 -275 37493
rect -2829 37390 -2802 37424
rect -2802 37390 -2795 37424
rect -2757 37390 -2734 37424
rect -2734 37390 -2723 37424
rect -2685 37390 -2666 37424
rect -2666 37390 -2651 37424
rect -2613 37390 -2598 37424
rect -2598 37390 -2579 37424
rect -2541 37390 -2530 37424
rect -2530 37390 -2507 37424
rect -2469 37390 -2462 37424
rect -2462 37390 -2435 37424
rect -2397 37390 -2394 37424
rect -2394 37390 -2363 37424
rect -2325 37390 -2292 37424
rect -2292 37390 -2291 37424
rect -2253 37390 -2224 37424
rect -2224 37390 -2219 37424
rect -2181 37390 -2156 37424
rect -2156 37390 -2147 37424
rect -2109 37390 -2088 37424
rect -2088 37390 -2075 37424
rect -2037 37390 -2020 37424
rect -2020 37390 -2003 37424
rect -1965 37390 -1952 37424
rect -1952 37390 -1931 37424
rect -1893 37390 -1884 37424
rect -1884 37390 -1859 37424
rect -1821 37390 -1816 37424
rect -1816 37390 -1787 37424
rect -1749 37390 -1748 37424
rect -1748 37390 -1715 37424
rect -1677 37390 -1646 37424
rect -1646 37390 -1643 37424
rect -1605 37390 -1578 37424
rect -1578 37390 -1571 37424
rect -1533 37390 -1510 37424
rect -1510 37390 -1499 37424
rect -1461 37390 -1442 37424
rect -1442 37390 -1427 37424
rect -1389 37390 -1374 37424
rect -1374 37390 -1355 37424
rect -1317 37390 -1306 37424
rect -1306 37390 -1283 37424
rect -1245 37390 -1238 37424
rect -1238 37390 -1211 37424
rect -1173 37390 -1170 37424
rect -1170 37390 -1139 37424
rect -1101 37390 -1068 37424
rect -1068 37390 -1067 37424
rect -1029 37390 -1000 37424
rect -1000 37390 -995 37424
rect -957 37390 -932 37424
rect -932 37390 -923 37424
rect -885 37390 -864 37424
rect -864 37390 -851 37424
rect -813 37390 -796 37424
rect -796 37390 -779 37424
rect -741 37390 -728 37424
rect -728 37390 -707 37424
rect -669 37390 -660 37424
rect -660 37390 -635 37424
rect -597 37390 -592 37424
rect -592 37390 -563 37424
rect -525 37390 -524 37424
rect -524 37390 -491 37424
rect -453 37390 -422 37424
rect -422 37390 -419 37424
rect -381 37390 -354 37424
rect -354 37390 -347 37424
rect -309 37390 -286 37424
rect -286 37390 -275 37424
rect -2829 37321 -2802 37351
rect -2802 37321 -2795 37351
rect -2757 37321 -2734 37351
rect -2734 37321 -2723 37351
rect -2685 37321 -2666 37351
rect -2666 37321 -2651 37351
rect -2613 37321 -2598 37351
rect -2598 37321 -2579 37351
rect -2541 37321 -2530 37351
rect -2530 37321 -2507 37351
rect -2469 37321 -2462 37351
rect -2462 37321 -2435 37351
rect -2397 37321 -2394 37351
rect -2394 37321 -2363 37351
rect -2325 37321 -2292 37351
rect -2292 37321 -2291 37351
rect -2253 37321 -2224 37351
rect -2224 37321 -2219 37351
rect -2181 37321 -2156 37351
rect -2156 37321 -2147 37351
rect -2109 37321 -2088 37351
rect -2088 37321 -2075 37351
rect -2037 37321 -2020 37351
rect -2020 37321 -2003 37351
rect -1965 37321 -1952 37351
rect -1952 37321 -1931 37351
rect -1893 37321 -1884 37351
rect -1884 37321 -1859 37351
rect -1821 37321 -1816 37351
rect -1816 37321 -1787 37351
rect -1749 37321 -1748 37351
rect -1748 37321 -1715 37351
rect -1677 37321 -1646 37351
rect -1646 37321 -1643 37351
rect -1605 37321 -1578 37351
rect -1578 37321 -1571 37351
rect -1533 37321 -1510 37351
rect -1510 37321 -1499 37351
rect -1461 37321 -1442 37351
rect -1442 37321 -1427 37351
rect -1389 37321 -1374 37351
rect -1374 37321 -1355 37351
rect -1317 37321 -1306 37351
rect -1306 37321 -1283 37351
rect -1245 37321 -1238 37351
rect -1238 37321 -1211 37351
rect -1173 37321 -1170 37351
rect -1170 37321 -1139 37351
rect -1101 37321 -1068 37351
rect -1068 37321 -1067 37351
rect -1029 37321 -1000 37351
rect -1000 37321 -995 37351
rect -957 37321 -932 37351
rect -932 37321 -923 37351
rect -885 37321 -864 37351
rect -864 37321 -851 37351
rect -813 37321 -796 37351
rect -796 37321 -779 37351
rect -741 37321 -728 37351
rect -728 37321 -707 37351
rect -669 37321 -660 37351
rect -660 37321 -635 37351
rect -597 37321 -592 37351
rect -592 37321 -563 37351
rect -525 37321 -524 37351
rect -524 37321 -491 37351
rect -453 37321 -422 37351
rect -422 37321 -419 37351
rect -381 37321 -354 37351
rect -354 37321 -347 37351
rect -309 37321 -286 37351
rect -286 37321 -275 37351
rect -2829 37317 -2795 37321
rect -2757 37317 -2723 37321
rect -2685 37317 -2651 37321
rect -2613 37317 -2579 37321
rect -2541 37317 -2507 37321
rect -2469 37317 -2435 37321
rect -2397 37317 -2363 37321
rect -2325 37317 -2291 37321
rect -2253 37317 -2219 37321
rect -2181 37317 -2147 37321
rect -2109 37317 -2075 37321
rect -2037 37317 -2003 37321
rect -1965 37317 -1931 37321
rect -1893 37317 -1859 37321
rect -1821 37317 -1787 37321
rect -1749 37317 -1715 37321
rect -1677 37317 -1643 37321
rect -1605 37317 -1571 37321
rect -1533 37317 -1499 37321
rect -1461 37317 -1427 37321
rect -1389 37317 -1355 37321
rect -1317 37317 -1283 37321
rect -1245 37317 -1211 37321
rect -1173 37317 -1139 37321
rect -1101 37317 -1067 37321
rect -1029 37317 -995 37321
rect -957 37317 -923 37321
rect -885 37317 -851 37321
rect -813 37317 -779 37321
rect -741 37317 -707 37321
rect -669 37317 -635 37321
rect -597 37317 -563 37321
rect -525 37317 -491 37321
rect -453 37317 -419 37321
rect -381 37317 -347 37321
rect -309 37317 -275 37321
rect -2829 37252 -2802 37278
rect -2802 37252 -2795 37278
rect -2757 37252 -2734 37278
rect -2734 37252 -2723 37278
rect -2685 37252 -2666 37278
rect -2666 37252 -2651 37278
rect -2613 37252 -2598 37278
rect -2598 37252 -2579 37278
rect -2541 37252 -2530 37278
rect -2530 37252 -2507 37278
rect -2469 37252 -2462 37278
rect -2462 37252 -2435 37278
rect -2397 37252 -2394 37278
rect -2394 37252 -2363 37278
rect -2325 37252 -2292 37278
rect -2292 37252 -2291 37278
rect -2253 37252 -2224 37278
rect -2224 37252 -2219 37278
rect -2181 37252 -2156 37278
rect -2156 37252 -2147 37278
rect -2109 37252 -2088 37278
rect -2088 37252 -2075 37278
rect -2037 37252 -2020 37278
rect -2020 37252 -2003 37278
rect -1965 37252 -1952 37278
rect -1952 37252 -1931 37278
rect -1893 37252 -1884 37278
rect -1884 37252 -1859 37278
rect -1821 37252 -1816 37278
rect -1816 37252 -1787 37278
rect -1749 37252 -1748 37278
rect -1748 37252 -1715 37278
rect -1677 37252 -1646 37278
rect -1646 37252 -1643 37278
rect -1605 37252 -1578 37278
rect -1578 37252 -1571 37278
rect -1533 37252 -1510 37278
rect -1510 37252 -1499 37278
rect -1461 37252 -1442 37278
rect -1442 37252 -1427 37278
rect -1389 37252 -1374 37278
rect -1374 37252 -1355 37278
rect -1317 37252 -1306 37278
rect -1306 37252 -1283 37278
rect -1245 37252 -1238 37278
rect -1238 37252 -1211 37278
rect -1173 37252 -1170 37278
rect -1170 37252 -1139 37278
rect -1101 37252 -1068 37278
rect -1068 37252 -1067 37278
rect -1029 37252 -1000 37278
rect -1000 37252 -995 37278
rect -957 37252 -932 37278
rect -932 37252 -923 37278
rect -885 37252 -864 37278
rect -864 37252 -851 37278
rect -813 37252 -796 37278
rect -796 37252 -779 37278
rect -741 37252 -728 37278
rect -728 37252 -707 37278
rect -669 37252 -660 37278
rect -660 37252 -635 37278
rect -597 37252 -592 37278
rect -592 37252 -563 37278
rect -525 37252 -524 37278
rect -524 37252 -491 37278
rect -453 37252 -422 37278
rect -422 37252 -419 37278
rect -381 37252 -354 37278
rect -354 37252 -347 37278
rect -309 37252 -286 37278
rect -286 37252 -275 37278
rect -2829 37244 -2795 37252
rect -2757 37244 -2723 37252
rect -2685 37244 -2651 37252
rect -2613 37244 -2579 37252
rect -2541 37244 -2507 37252
rect -2469 37244 -2435 37252
rect -2397 37244 -2363 37252
rect -2325 37244 -2291 37252
rect -2253 37244 -2219 37252
rect -2181 37244 -2147 37252
rect -2109 37244 -2075 37252
rect -2037 37244 -2003 37252
rect -1965 37244 -1931 37252
rect -1893 37244 -1859 37252
rect -1821 37244 -1787 37252
rect -1749 37244 -1715 37252
rect -1677 37244 -1643 37252
rect -1605 37244 -1571 37252
rect -1533 37244 -1499 37252
rect -1461 37244 -1427 37252
rect -1389 37244 -1355 37252
rect -1317 37244 -1283 37252
rect -1245 37244 -1211 37252
rect -1173 37244 -1139 37252
rect -1101 37244 -1067 37252
rect -1029 37244 -995 37252
rect -957 37244 -923 37252
rect -885 37244 -851 37252
rect -813 37244 -779 37252
rect -741 37244 -707 37252
rect -669 37244 -635 37252
rect -597 37244 -563 37252
rect -525 37244 -491 37252
rect -453 37244 -419 37252
rect -381 37244 -347 37252
rect -309 37244 -275 37252
rect -2829 37183 -2802 37205
rect -2802 37183 -2795 37205
rect -2757 37183 -2734 37205
rect -2734 37183 -2723 37205
rect -2685 37183 -2666 37205
rect -2666 37183 -2651 37205
rect -2613 37183 -2598 37205
rect -2598 37183 -2579 37205
rect -2541 37183 -2530 37205
rect -2530 37183 -2507 37205
rect -2469 37183 -2462 37205
rect -2462 37183 -2435 37205
rect -2397 37183 -2394 37205
rect -2394 37183 -2363 37205
rect -2325 37183 -2292 37205
rect -2292 37183 -2291 37205
rect -2253 37183 -2224 37205
rect -2224 37183 -2219 37205
rect -2181 37183 -2156 37205
rect -2156 37183 -2147 37205
rect -2109 37183 -2088 37205
rect -2088 37183 -2075 37205
rect -2037 37183 -2020 37205
rect -2020 37183 -2003 37205
rect -1965 37183 -1952 37205
rect -1952 37183 -1931 37205
rect -1893 37183 -1884 37205
rect -1884 37183 -1859 37205
rect -1821 37183 -1816 37205
rect -1816 37183 -1787 37205
rect -1749 37183 -1748 37205
rect -1748 37183 -1715 37205
rect -1677 37183 -1646 37205
rect -1646 37183 -1643 37205
rect -1605 37183 -1578 37205
rect -1578 37183 -1571 37205
rect -1533 37183 -1510 37205
rect -1510 37183 -1499 37205
rect -1461 37183 -1442 37205
rect -1442 37183 -1427 37205
rect -1389 37183 -1374 37205
rect -1374 37183 -1355 37205
rect -1317 37183 -1306 37205
rect -1306 37183 -1283 37205
rect -1245 37183 -1238 37205
rect -1238 37183 -1211 37205
rect -1173 37183 -1170 37205
rect -1170 37183 -1139 37205
rect -1101 37183 -1068 37205
rect -1068 37183 -1067 37205
rect -1029 37183 -1000 37205
rect -1000 37183 -995 37205
rect -957 37183 -932 37205
rect -932 37183 -923 37205
rect -885 37183 -864 37205
rect -864 37183 -851 37205
rect -813 37183 -796 37205
rect -796 37183 -779 37205
rect -741 37183 -728 37205
rect -728 37183 -707 37205
rect -669 37183 -660 37205
rect -660 37183 -635 37205
rect -597 37183 -592 37205
rect -592 37183 -563 37205
rect -525 37183 -524 37205
rect -524 37183 -491 37205
rect -453 37183 -422 37205
rect -422 37183 -419 37205
rect -381 37183 -354 37205
rect -354 37183 -347 37205
rect -309 37183 -286 37205
rect -286 37183 -275 37205
rect -2829 37171 -2795 37183
rect -2757 37171 -2723 37183
rect -2685 37171 -2651 37183
rect -2613 37171 -2579 37183
rect -2541 37171 -2507 37183
rect -2469 37171 -2435 37183
rect -2397 37171 -2363 37183
rect -2325 37171 -2291 37183
rect -2253 37171 -2219 37183
rect -2181 37171 -2147 37183
rect -2109 37171 -2075 37183
rect -2037 37171 -2003 37183
rect -1965 37171 -1931 37183
rect -1893 37171 -1859 37183
rect -1821 37171 -1787 37183
rect -1749 37171 -1715 37183
rect -1677 37171 -1643 37183
rect -1605 37171 -1571 37183
rect -1533 37171 -1499 37183
rect -1461 37171 -1427 37183
rect -1389 37171 -1355 37183
rect -1317 37171 -1283 37183
rect -1245 37171 -1211 37183
rect -1173 37171 -1139 37183
rect -1101 37171 -1067 37183
rect -1029 37171 -995 37183
rect -957 37171 -923 37183
rect -885 37171 -851 37183
rect -813 37171 -779 37183
rect -741 37171 -707 37183
rect -669 37171 -635 37183
rect -597 37171 -563 37183
rect -525 37171 -491 37183
rect -453 37171 -419 37183
rect -381 37171 -347 37183
rect -309 37171 -275 37183
rect -2829 37114 -2802 37132
rect -2802 37114 -2795 37132
rect -2757 37114 -2734 37132
rect -2734 37114 -2723 37132
rect -2685 37114 -2666 37132
rect -2666 37114 -2651 37132
rect -2613 37114 -2598 37132
rect -2598 37114 -2579 37132
rect -2541 37114 -2530 37132
rect -2530 37114 -2507 37132
rect -2469 37114 -2462 37132
rect -2462 37114 -2435 37132
rect -2397 37114 -2394 37132
rect -2394 37114 -2363 37132
rect -2325 37114 -2292 37132
rect -2292 37114 -2291 37132
rect -2253 37114 -2224 37132
rect -2224 37114 -2219 37132
rect -2181 37114 -2156 37132
rect -2156 37114 -2147 37132
rect -2109 37114 -2088 37132
rect -2088 37114 -2075 37132
rect -2037 37114 -2020 37132
rect -2020 37114 -2003 37132
rect -1965 37114 -1952 37132
rect -1952 37114 -1931 37132
rect -1893 37114 -1884 37132
rect -1884 37114 -1859 37132
rect -1821 37114 -1816 37132
rect -1816 37114 -1787 37132
rect -1749 37114 -1748 37132
rect -1748 37114 -1715 37132
rect -1677 37114 -1646 37132
rect -1646 37114 -1643 37132
rect -1605 37114 -1578 37132
rect -1578 37114 -1571 37132
rect -1533 37114 -1510 37132
rect -1510 37114 -1499 37132
rect -1461 37114 -1442 37132
rect -1442 37114 -1427 37132
rect -1389 37114 -1374 37132
rect -1374 37114 -1355 37132
rect -1317 37114 -1306 37132
rect -1306 37114 -1283 37132
rect -1245 37114 -1238 37132
rect -1238 37114 -1211 37132
rect -1173 37114 -1170 37132
rect -1170 37114 -1139 37132
rect -1101 37114 -1068 37132
rect -1068 37114 -1067 37132
rect -1029 37114 -1000 37132
rect -1000 37114 -995 37132
rect -957 37114 -932 37132
rect -932 37114 -923 37132
rect -885 37114 -864 37132
rect -864 37114 -851 37132
rect -813 37114 -796 37132
rect -796 37114 -779 37132
rect -741 37114 -728 37132
rect -728 37114 -707 37132
rect -669 37114 -660 37132
rect -660 37114 -635 37132
rect -597 37114 -592 37132
rect -592 37114 -563 37132
rect -525 37114 -524 37132
rect -524 37114 -491 37132
rect -453 37114 -422 37132
rect -422 37114 -419 37132
rect -381 37114 -354 37132
rect -354 37114 -347 37132
rect -309 37114 -286 37132
rect -286 37114 -275 37132
rect -2829 37098 -2795 37114
rect -2757 37098 -2723 37114
rect -2685 37098 -2651 37114
rect -2613 37098 -2579 37114
rect -2541 37098 -2507 37114
rect -2469 37098 -2435 37114
rect -2397 37098 -2363 37114
rect -2325 37098 -2291 37114
rect -2253 37098 -2219 37114
rect -2181 37098 -2147 37114
rect -2109 37098 -2075 37114
rect -2037 37098 -2003 37114
rect -1965 37098 -1931 37114
rect -1893 37098 -1859 37114
rect -1821 37098 -1787 37114
rect -1749 37098 -1715 37114
rect -1677 37098 -1643 37114
rect -1605 37098 -1571 37114
rect -1533 37098 -1499 37114
rect -1461 37098 -1427 37114
rect -1389 37098 -1355 37114
rect -1317 37098 -1283 37114
rect -1245 37098 -1211 37114
rect -1173 37098 -1139 37114
rect -1101 37098 -1067 37114
rect -1029 37098 -995 37114
rect -957 37098 -923 37114
rect -885 37098 -851 37114
rect -813 37098 -779 37114
rect -741 37098 -707 37114
rect -669 37098 -635 37114
rect -597 37098 -563 37114
rect -525 37098 -491 37114
rect -453 37098 -419 37114
rect -381 37098 -347 37114
rect -309 37098 -275 37114
rect -2829 37045 -2802 37059
rect -2802 37045 -2795 37059
rect -2757 37045 -2734 37059
rect -2734 37045 -2723 37059
rect -2685 37045 -2666 37059
rect -2666 37045 -2651 37059
rect -2613 37045 -2598 37059
rect -2598 37045 -2579 37059
rect -2541 37045 -2530 37059
rect -2530 37045 -2507 37059
rect -2469 37045 -2462 37059
rect -2462 37045 -2435 37059
rect -2397 37045 -2394 37059
rect -2394 37045 -2363 37059
rect -2325 37045 -2292 37059
rect -2292 37045 -2291 37059
rect -2253 37045 -2224 37059
rect -2224 37045 -2219 37059
rect -2181 37045 -2156 37059
rect -2156 37045 -2147 37059
rect -2109 37045 -2088 37059
rect -2088 37045 -2075 37059
rect -2037 37045 -2020 37059
rect -2020 37045 -2003 37059
rect -1965 37045 -1952 37059
rect -1952 37045 -1931 37059
rect -1893 37045 -1884 37059
rect -1884 37045 -1859 37059
rect -1821 37045 -1816 37059
rect -1816 37045 -1787 37059
rect -1749 37045 -1748 37059
rect -1748 37045 -1715 37059
rect -1677 37045 -1646 37059
rect -1646 37045 -1643 37059
rect -1605 37045 -1578 37059
rect -1578 37045 -1571 37059
rect -1533 37045 -1510 37059
rect -1510 37045 -1499 37059
rect -1461 37045 -1442 37059
rect -1442 37045 -1427 37059
rect -1389 37045 -1374 37059
rect -1374 37045 -1355 37059
rect -1317 37045 -1306 37059
rect -1306 37045 -1283 37059
rect -1245 37045 -1238 37059
rect -1238 37045 -1211 37059
rect -1173 37045 -1170 37059
rect -1170 37045 -1139 37059
rect -1101 37045 -1068 37059
rect -1068 37045 -1067 37059
rect -1029 37045 -1000 37059
rect -1000 37045 -995 37059
rect -957 37045 -932 37059
rect -932 37045 -923 37059
rect -885 37045 -864 37059
rect -864 37045 -851 37059
rect -813 37045 -796 37059
rect -796 37045 -779 37059
rect -741 37045 -728 37059
rect -728 37045 -707 37059
rect -669 37045 -660 37059
rect -660 37045 -635 37059
rect -597 37045 -592 37059
rect -592 37045 -563 37059
rect -525 37045 -524 37059
rect -524 37045 -491 37059
rect -453 37045 -422 37059
rect -422 37045 -419 37059
rect -381 37045 -354 37059
rect -354 37045 -347 37059
rect -309 37045 -286 37059
rect -286 37045 -275 37059
rect -2829 37025 -2795 37045
rect -2757 37025 -2723 37045
rect -2685 37025 -2651 37045
rect -2613 37025 -2579 37045
rect -2541 37025 -2507 37045
rect -2469 37025 -2435 37045
rect -2397 37025 -2363 37045
rect -2325 37025 -2291 37045
rect -2253 37025 -2219 37045
rect -2181 37025 -2147 37045
rect -2109 37025 -2075 37045
rect -2037 37025 -2003 37045
rect -1965 37025 -1931 37045
rect -1893 37025 -1859 37045
rect -1821 37025 -1787 37045
rect -1749 37025 -1715 37045
rect -1677 37025 -1643 37045
rect -1605 37025 -1571 37045
rect -1533 37025 -1499 37045
rect -1461 37025 -1427 37045
rect -1389 37025 -1355 37045
rect -1317 37025 -1283 37045
rect -1245 37025 -1211 37045
rect -1173 37025 -1139 37045
rect -1101 37025 -1067 37045
rect -1029 37025 -995 37045
rect -957 37025 -923 37045
rect -885 37025 -851 37045
rect -813 37025 -779 37045
rect -741 37025 -707 37045
rect -669 37025 -635 37045
rect -597 37025 -563 37045
rect -525 37025 -491 37045
rect -453 37025 -419 37045
rect -381 37025 -347 37045
rect -309 37025 -275 37045
rect -2829 36976 -2802 36986
rect -2802 36976 -2795 36986
rect -2757 36976 -2734 36986
rect -2734 36976 -2723 36986
rect -2685 36976 -2666 36986
rect -2666 36976 -2651 36986
rect -2613 36976 -2598 36986
rect -2598 36976 -2579 36986
rect -2541 36976 -2530 36986
rect -2530 36976 -2507 36986
rect -2469 36976 -2462 36986
rect -2462 36976 -2435 36986
rect -2397 36976 -2394 36986
rect -2394 36976 -2363 36986
rect -2325 36976 -2292 36986
rect -2292 36976 -2291 36986
rect -2253 36976 -2224 36986
rect -2224 36976 -2219 36986
rect -2181 36976 -2156 36986
rect -2156 36976 -2147 36986
rect -2109 36976 -2088 36986
rect -2088 36976 -2075 36986
rect -2037 36976 -2020 36986
rect -2020 36976 -2003 36986
rect -1965 36976 -1952 36986
rect -1952 36976 -1931 36986
rect -1893 36976 -1884 36986
rect -1884 36976 -1859 36986
rect -1821 36976 -1816 36986
rect -1816 36976 -1787 36986
rect -1749 36976 -1748 36986
rect -1748 36976 -1715 36986
rect -1677 36976 -1646 36986
rect -1646 36976 -1643 36986
rect -1605 36976 -1578 36986
rect -1578 36976 -1571 36986
rect -1533 36976 -1510 36986
rect -1510 36976 -1499 36986
rect -1461 36976 -1442 36986
rect -1442 36976 -1427 36986
rect -1389 36976 -1374 36986
rect -1374 36976 -1355 36986
rect -1317 36976 -1306 36986
rect -1306 36976 -1283 36986
rect -1245 36976 -1238 36986
rect -1238 36976 -1211 36986
rect -1173 36976 -1170 36986
rect -1170 36976 -1139 36986
rect -1101 36976 -1068 36986
rect -1068 36976 -1067 36986
rect -1029 36976 -1000 36986
rect -1000 36976 -995 36986
rect -957 36976 -932 36986
rect -932 36976 -923 36986
rect -885 36976 -864 36986
rect -864 36976 -851 36986
rect -813 36976 -796 36986
rect -796 36976 -779 36986
rect -741 36976 -728 36986
rect -728 36976 -707 36986
rect -669 36976 -660 36986
rect -660 36976 -635 36986
rect -597 36976 -592 36986
rect -592 36976 -563 36986
rect -525 36976 -524 36986
rect -524 36976 -491 36986
rect -453 36976 -422 36986
rect -422 36976 -419 36986
rect -381 36976 -354 36986
rect -354 36976 -347 36986
rect -309 36976 -286 36986
rect -286 36976 -275 36986
rect -2829 36952 -2795 36976
rect -2757 36952 -2723 36976
rect -2685 36952 -2651 36976
rect -2613 36952 -2579 36976
rect -2541 36952 -2507 36976
rect -2469 36952 -2435 36976
rect -2397 36952 -2363 36976
rect -2325 36952 -2291 36976
rect -2253 36952 -2219 36976
rect -2181 36952 -2147 36976
rect -2109 36952 -2075 36976
rect -2037 36952 -2003 36976
rect -1965 36952 -1931 36976
rect -1893 36952 -1859 36976
rect -1821 36952 -1787 36976
rect -1749 36952 -1715 36976
rect -1677 36952 -1643 36976
rect -1605 36952 -1571 36976
rect -1533 36952 -1499 36976
rect -1461 36952 -1427 36976
rect -1389 36952 -1355 36976
rect -1317 36952 -1283 36976
rect -1245 36952 -1211 36976
rect -1173 36952 -1139 36976
rect -1101 36952 -1067 36976
rect -1029 36952 -995 36976
rect -957 36952 -923 36976
rect -885 36952 -851 36976
rect -813 36952 -779 36976
rect -741 36952 -707 36976
rect -669 36952 -635 36976
rect -597 36952 -563 36976
rect -525 36952 -491 36976
rect -453 36952 -419 36976
rect -381 36952 -347 36976
rect -309 36952 -275 36976
rect -2829 36907 -2802 36913
rect -2802 36907 -2795 36913
rect -2757 36907 -2734 36913
rect -2734 36907 -2723 36913
rect -2685 36907 -2666 36913
rect -2666 36907 -2651 36913
rect -2613 36907 -2598 36913
rect -2598 36907 -2579 36913
rect -2541 36907 -2530 36913
rect -2530 36907 -2507 36913
rect -2469 36907 -2462 36913
rect -2462 36907 -2435 36913
rect -2397 36907 -2394 36913
rect -2394 36907 -2363 36913
rect -2325 36907 -2292 36913
rect -2292 36907 -2291 36913
rect -2253 36907 -2224 36913
rect -2224 36907 -2219 36913
rect -2181 36907 -2156 36913
rect -2156 36907 -2147 36913
rect -2109 36907 -2088 36913
rect -2088 36907 -2075 36913
rect -2037 36907 -2020 36913
rect -2020 36907 -2003 36913
rect -1965 36907 -1952 36913
rect -1952 36907 -1931 36913
rect -1893 36907 -1884 36913
rect -1884 36907 -1859 36913
rect -1821 36907 -1816 36913
rect -1816 36907 -1787 36913
rect -1749 36907 -1748 36913
rect -1748 36907 -1715 36913
rect -1677 36907 -1646 36913
rect -1646 36907 -1643 36913
rect -1605 36907 -1578 36913
rect -1578 36907 -1571 36913
rect -1533 36907 -1510 36913
rect -1510 36907 -1499 36913
rect -1461 36907 -1442 36913
rect -1442 36907 -1427 36913
rect -1389 36907 -1374 36913
rect -1374 36907 -1355 36913
rect -1317 36907 -1306 36913
rect -1306 36907 -1283 36913
rect -1245 36907 -1238 36913
rect -1238 36907 -1211 36913
rect -1173 36907 -1170 36913
rect -1170 36907 -1139 36913
rect -1101 36907 -1068 36913
rect -1068 36907 -1067 36913
rect -1029 36907 -1000 36913
rect -1000 36907 -995 36913
rect -957 36907 -932 36913
rect -932 36907 -923 36913
rect -885 36907 -864 36913
rect -864 36907 -851 36913
rect -813 36907 -796 36913
rect -796 36907 -779 36913
rect -741 36907 -728 36913
rect -728 36907 -707 36913
rect -669 36907 -660 36913
rect -660 36907 -635 36913
rect -597 36907 -592 36913
rect -592 36907 -563 36913
rect -525 36907 -524 36913
rect -524 36907 -491 36913
rect -453 36907 -422 36913
rect -422 36907 -419 36913
rect -381 36907 -354 36913
rect -354 36907 -347 36913
rect -309 36907 -286 36913
rect -286 36907 -275 36913
rect -2829 36879 -2795 36907
rect -2757 36879 -2723 36907
rect -2685 36879 -2651 36907
rect -2613 36879 -2579 36907
rect -2541 36879 -2507 36907
rect -2469 36879 -2435 36907
rect -2397 36879 -2363 36907
rect -2325 36879 -2291 36907
rect -2253 36879 -2219 36907
rect -2181 36879 -2147 36907
rect -2109 36879 -2075 36907
rect -2037 36879 -2003 36907
rect -1965 36879 -1931 36907
rect -1893 36879 -1859 36907
rect -1821 36879 -1787 36907
rect -1749 36879 -1715 36907
rect -1677 36879 -1643 36907
rect -1605 36879 -1571 36907
rect -1533 36879 -1499 36907
rect -1461 36879 -1427 36907
rect -1389 36879 -1355 36907
rect -1317 36879 -1283 36907
rect -1245 36879 -1211 36907
rect -1173 36879 -1139 36907
rect -1101 36879 -1067 36907
rect -1029 36879 -995 36907
rect -957 36879 -923 36907
rect -885 36879 -851 36907
rect -813 36879 -779 36907
rect -741 36879 -707 36907
rect -669 36879 -635 36907
rect -597 36879 -563 36907
rect -525 36879 -491 36907
rect -453 36879 -419 36907
rect -381 36879 -347 36907
rect -309 36879 -275 36907
rect -2829 36838 -2802 36840
rect -2802 36838 -2795 36840
rect -2757 36838 -2734 36840
rect -2734 36838 -2723 36840
rect -2685 36838 -2666 36840
rect -2666 36838 -2651 36840
rect -2613 36838 -2598 36840
rect -2598 36838 -2579 36840
rect -2541 36838 -2530 36840
rect -2530 36838 -2507 36840
rect -2469 36838 -2462 36840
rect -2462 36838 -2435 36840
rect -2397 36838 -2394 36840
rect -2394 36838 -2363 36840
rect -2325 36838 -2292 36840
rect -2292 36838 -2291 36840
rect -2253 36838 -2224 36840
rect -2224 36838 -2219 36840
rect -2181 36838 -2156 36840
rect -2156 36838 -2147 36840
rect -2109 36838 -2088 36840
rect -2088 36838 -2075 36840
rect -2037 36838 -2020 36840
rect -2020 36838 -2003 36840
rect -1965 36838 -1952 36840
rect -1952 36838 -1931 36840
rect -1893 36838 -1884 36840
rect -1884 36838 -1859 36840
rect -1821 36838 -1816 36840
rect -1816 36838 -1787 36840
rect -1749 36838 -1748 36840
rect -1748 36838 -1715 36840
rect -1677 36838 -1646 36840
rect -1646 36838 -1643 36840
rect -1605 36838 -1578 36840
rect -1578 36838 -1571 36840
rect -1533 36838 -1510 36840
rect -1510 36838 -1499 36840
rect -1461 36838 -1442 36840
rect -1442 36838 -1427 36840
rect -1389 36838 -1374 36840
rect -1374 36838 -1355 36840
rect -1317 36838 -1306 36840
rect -1306 36838 -1283 36840
rect -1245 36838 -1238 36840
rect -1238 36838 -1211 36840
rect -1173 36838 -1170 36840
rect -1170 36838 -1139 36840
rect -1101 36838 -1068 36840
rect -1068 36838 -1067 36840
rect -1029 36838 -1000 36840
rect -1000 36838 -995 36840
rect -957 36838 -932 36840
rect -932 36838 -923 36840
rect -885 36838 -864 36840
rect -864 36838 -851 36840
rect -813 36838 -796 36840
rect -796 36838 -779 36840
rect -741 36838 -728 36840
rect -728 36838 -707 36840
rect -669 36838 -660 36840
rect -660 36838 -635 36840
rect -597 36838 -592 36840
rect -592 36838 -563 36840
rect -525 36838 -524 36840
rect -524 36838 -491 36840
rect -453 36838 -422 36840
rect -422 36838 -419 36840
rect -381 36838 -354 36840
rect -354 36838 -347 36840
rect -309 36838 -286 36840
rect -286 36838 -275 36840
rect -2829 36806 -2795 36838
rect -2757 36806 -2723 36838
rect -2685 36806 -2651 36838
rect -2613 36806 -2579 36838
rect -2541 36806 -2507 36838
rect -2469 36806 -2435 36838
rect -2397 36806 -2363 36838
rect -2325 36806 -2291 36838
rect -2253 36806 -2219 36838
rect -2181 36806 -2147 36838
rect -2109 36806 -2075 36838
rect -2037 36806 -2003 36838
rect -1965 36806 -1931 36838
rect -1893 36806 -1859 36838
rect -1821 36806 -1787 36838
rect -1749 36806 -1715 36838
rect -1677 36806 -1643 36838
rect -1605 36806 -1571 36838
rect -1533 36806 -1499 36838
rect -1461 36806 -1427 36838
rect -1389 36806 -1355 36838
rect -1317 36806 -1283 36838
rect -1245 36806 -1211 36838
rect -1173 36806 -1139 36838
rect -1101 36806 -1067 36838
rect -1029 36806 -995 36838
rect -957 36806 -923 36838
rect -885 36806 -851 36838
rect -813 36806 -779 36838
rect -741 36806 -707 36838
rect -669 36806 -635 36838
rect -597 36806 -563 36838
rect -525 36806 -491 36838
rect -453 36806 -419 36838
rect -381 36806 -347 36838
rect -309 36806 -275 36838
rect -2829 36734 -2795 36767
rect -2757 36734 -2723 36767
rect -2685 36734 -2651 36767
rect -2613 36734 -2579 36767
rect -2541 36734 -2507 36767
rect -2469 36734 -2435 36767
rect -2397 36734 -2363 36767
rect -2325 36734 -2291 36767
rect -2253 36734 -2219 36767
rect -2181 36734 -2147 36767
rect -2109 36734 -2075 36767
rect -2037 36734 -2003 36767
rect -1965 36734 -1931 36767
rect -1893 36734 -1859 36767
rect -1821 36734 -1787 36767
rect -1749 36734 -1715 36767
rect -1677 36734 -1643 36767
rect -1605 36734 -1571 36767
rect -1533 36734 -1499 36767
rect -1461 36734 -1427 36767
rect -1389 36734 -1355 36767
rect -1317 36734 -1283 36767
rect -1245 36734 -1211 36767
rect -1173 36734 -1139 36767
rect -1101 36734 -1067 36767
rect -1029 36734 -995 36767
rect -957 36734 -923 36767
rect -885 36734 -851 36767
rect -813 36734 -779 36767
rect -741 36734 -707 36767
rect -669 36734 -635 36767
rect -597 36734 -563 36767
rect -525 36734 -491 36767
rect -453 36734 -419 36767
rect -381 36734 -347 36767
rect -309 36734 -275 36767
rect -2829 36733 -2802 36734
rect -2802 36733 -2795 36734
rect -2757 36733 -2734 36734
rect -2734 36733 -2723 36734
rect -2685 36733 -2666 36734
rect -2666 36733 -2651 36734
rect -2613 36733 -2598 36734
rect -2598 36733 -2579 36734
rect -2541 36733 -2530 36734
rect -2530 36733 -2507 36734
rect -2469 36733 -2462 36734
rect -2462 36733 -2435 36734
rect -2397 36733 -2394 36734
rect -2394 36733 -2363 36734
rect -2325 36733 -2292 36734
rect -2292 36733 -2291 36734
rect -2253 36733 -2224 36734
rect -2224 36733 -2219 36734
rect -2181 36733 -2156 36734
rect -2156 36733 -2147 36734
rect -2109 36733 -2088 36734
rect -2088 36733 -2075 36734
rect -2037 36733 -2020 36734
rect -2020 36733 -2003 36734
rect -1965 36733 -1952 36734
rect -1952 36733 -1931 36734
rect -1893 36733 -1884 36734
rect -1884 36733 -1859 36734
rect -1821 36733 -1816 36734
rect -1816 36733 -1787 36734
rect -1749 36733 -1748 36734
rect -1748 36733 -1715 36734
rect -1677 36733 -1646 36734
rect -1646 36733 -1643 36734
rect -1605 36733 -1578 36734
rect -1578 36733 -1571 36734
rect -1533 36733 -1510 36734
rect -1510 36733 -1499 36734
rect -1461 36733 -1442 36734
rect -1442 36733 -1427 36734
rect -1389 36733 -1374 36734
rect -1374 36733 -1355 36734
rect -1317 36733 -1306 36734
rect -1306 36733 -1283 36734
rect -1245 36733 -1238 36734
rect -1238 36733 -1211 36734
rect -1173 36733 -1170 36734
rect -1170 36733 -1139 36734
rect -1101 36733 -1068 36734
rect -1068 36733 -1067 36734
rect -1029 36733 -1000 36734
rect -1000 36733 -995 36734
rect -957 36733 -932 36734
rect -932 36733 -923 36734
rect -885 36733 -864 36734
rect -864 36733 -851 36734
rect -813 36733 -796 36734
rect -796 36733 -779 36734
rect -741 36733 -728 36734
rect -728 36733 -707 36734
rect -669 36733 -660 36734
rect -660 36733 -635 36734
rect -597 36733 -592 36734
rect -592 36733 -563 36734
rect -525 36733 -524 36734
rect -524 36733 -491 36734
rect -453 36733 -422 36734
rect -422 36733 -419 36734
rect -381 36733 -354 36734
rect -354 36733 -347 36734
rect -309 36733 -286 36734
rect -286 36733 -275 36734
rect -2829 36665 -2795 36694
rect -2757 36665 -2723 36694
rect -2685 36665 -2651 36694
rect -2613 36665 -2579 36694
rect -2541 36665 -2507 36694
rect -2469 36665 -2435 36694
rect -2397 36665 -2363 36694
rect -2325 36665 -2291 36694
rect -2253 36665 -2219 36694
rect -2181 36665 -2147 36694
rect -2109 36665 -2075 36694
rect -2037 36665 -2003 36694
rect -1965 36665 -1931 36694
rect -1893 36665 -1859 36694
rect -1821 36665 -1787 36694
rect -1749 36665 -1715 36694
rect -1677 36665 -1643 36694
rect -1605 36665 -1571 36694
rect -1533 36665 -1499 36694
rect -1461 36665 -1427 36694
rect -1389 36665 -1355 36694
rect -1317 36665 -1283 36694
rect -1245 36665 -1211 36694
rect -1173 36665 -1139 36694
rect -1101 36665 -1067 36694
rect -1029 36665 -995 36694
rect -957 36665 -923 36694
rect -885 36665 -851 36694
rect -813 36665 -779 36694
rect -741 36665 -707 36694
rect -669 36665 -635 36694
rect -597 36665 -563 36694
rect -525 36665 -491 36694
rect -453 36665 -419 36694
rect -381 36665 -347 36694
rect -309 36665 -275 36694
rect -2829 36660 -2802 36665
rect -2802 36660 -2795 36665
rect -2757 36660 -2734 36665
rect -2734 36660 -2723 36665
rect -2685 36660 -2666 36665
rect -2666 36660 -2651 36665
rect -2613 36660 -2598 36665
rect -2598 36660 -2579 36665
rect -2541 36660 -2530 36665
rect -2530 36660 -2507 36665
rect -2469 36660 -2462 36665
rect -2462 36660 -2435 36665
rect -2397 36660 -2394 36665
rect -2394 36660 -2363 36665
rect -2325 36660 -2292 36665
rect -2292 36660 -2291 36665
rect -2253 36660 -2224 36665
rect -2224 36660 -2219 36665
rect -2181 36660 -2156 36665
rect -2156 36660 -2147 36665
rect -2109 36660 -2088 36665
rect -2088 36660 -2075 36665
rect -2037 36660 -2020 36665
rect -2020 36660 -2003 36665
rect -1965 36660 -1952 36665
rect -1952 36660 -1931 36665
rect -1893 36660 -1884 36665
rect -1884 36660 -1859 36665
rect -1821 36660 -1816 36665
rect -1816 36660 -1787 36665
rect -1749 36660 -1748 36665
rect -1748 36660 -1715 36665
rect -1677 36660 -1646 36665
rect -1646 36660 -1643 36665
rect -1605 36660 -1578 36665
rect -1578 36660 -1571 36665
rect -1533 36660 -1510 36665
rect -1510 36660 -1499 36665
rect -1461 36660 -1442 36665
rect -1442 36660 -1427 36665
rect -1389 36660 -1374 36665
rect -1374 36660 -1355 36665
rect -1317 36660 -1306 36665
rect -1306 36660 -1283 36665
rect -1245 36660 -1238 36665
rect -1238 36660 -1211 36665
rect -1173 36660 -1170 36665
rect -1170 36660 -1139 36665
rect -1101 36660 -1068 36665
rect -1068 36660 -1067 36665
rect -1029 36660 -1000 36665
rect -1000 36660 -995 36665
rect -957 36660 -932 36665
rect -932 36660 -923 36665
rect -885 36660 -864 36665
rect -864 36660 -851 36665
rect -813 36660 -796 36665
rect -796 36660 -779 36665
rect -741 36660 -728 36665
rect -728 36660 -707 36665
rect -669 36660 -660 36665
rect -660 36660 -635 36665
rect -597 36660 -592 36665
rect -592 36660 -563 36665
rect -525 36660 -524 36665
rect -524 36660 -491 36665
rect -453 36660 -422 36665
rect -422 36660 -419 36665
rect -381 36660 -354 36665
rect -354 36660 -347 36665
rect -309 36660 -286 36665
rect -286 36660 -275 36665
rect -2829 36596 -2795 36621
rect -2757 36596 -2723 36621
rect -2685 36596 -2651 36621
rect -2613 36596 -2579 36621
rect -2541 36596 -2507 36621
rect -2469 36596 -2435 36621
rect -2397 36596 -2363 36621
rect -2325 36596 -2291 36621
rect -2253 36596 -2219 36621
rect -2181 36596 -2147 36621
rect -2109 36596 -2075 36621
rect -2037 36596 -2003 36621
rect -1965 36596 -1931 36621
rect -1893 36596 -1859 36621
rect -1821 36596 -1787 36621
rect -1749 36596 -1715 36621
rect -1677 36596 -1643 36621
rect -1605 36596 -1571 36621
rect -1533 36596 -1499 36621
rect -1461 36596 -1427 36621
rect -1389 36596 -1355 36621
rect -1317 36596 -1283 36621
rect -1245 36596 -1211 36621
rect -1173 36596 -1139 36621
rect -1101 36596 -1067 36621
rect -1029 36596 -995 36621
rect -957 36596 -923 36621
rect -885 36596 -851 36621
rect -813 36596 -779 36621
rect -741 36596 -707 36621
rect -669 36596 -635 36621
rect -597 36596 -563 36621
rect -525 36596 -491 36621
rect -453 36596 -419 36621
rect -381 36596 -347 36621
rect -309 36596 -275 36621
rect -2829 36587 -2802 36596
rect -2802 36587 -2795 36596
rect -2757 36587 -2734 36596
rect -2734 36587 -2723 36596
rect -2685 36587 -2666 36596
rect -2666 36587 -2651 36596
rect -2613 36587 -2598 36596
rect -2598 36587 -2579 36596
rect -2541 36587 -2530 36596
rect -2530 36587 -2507 36596
rect -2469 36587 -2462 36596
rect -2462 36587 -2435 36596
rect -2397 36587 -2394 36596
rect -2394 36587 -2363 36596
rect -2325 36587 -2292 36596
rect -2292 36587 -2291 36596
rect -2253 36587 -2224 36596
rect -2224 36587 -2219 36596
rect -2181 36587 -2156 36596
rect -2156 36587 -2147 36596
rect -2109 36587 -2088 36596
rect -2088 36587 -2075 36596
rect -2037 36587 -2020 36596
rect -2020 36587 -2003 36596
rect -1965 36587 -1952 36596
rect -1952 36587 -1931 36596
rect -1893 36587 -1884 36596
rect -1884 36587 -1859 36596
rect -1821 36587 -1816 36596
rect -1816 36587 -1787 36596
rect -1749 36587 -1748 36596
rect -1748 36587 -1715 36596
rect -1677 36587 -1646 36596
rect -1646 36587 -1643 36596
rect -1605 36587 -1578 36596
rect -1578 36587 -1571 36596
rect -1533 36587 -1510 36596
rect -1510 36587 -1499 36596
rect -1461 36587 -1442 36596
rect -1442 36587 -1427 36596
rect -1389 36587 -1374 36596
rect -1374 36587 -1355 36596
rect -1317 36587 -1306 36596
rect -1306 36587 -1283 36596
rect -1245 36587 -1238 36596
rect -1238 36587 -1211 36596
rect -1173 36587 -1170 36596
rect -1170 36587 -1139 36596
rect -1101 36587 -1068 36596
rect -1068 36587 -1067 36596
rect -1029 36587 -1000 36596
rect -1000 36587 -995 36596
rect -957 36587 -932 36596
rect -932 36587 -923 36596
rect -885 36587 -864 36596
rect -864 36587 -851 36596
rect -813 36587 -796 36596
rect -796 36587 -779 36596
rect -741 36587 -728 36596
rect -728 36587 -707 36596
rect -669 36587 -660 36596
rect -660 36587 -635 36596
rect -597 36587 -592 36596
rect -592 36587 -563 36596
rect -525 36587 -524 36596
rect -524 36587 -491 36596
rect -453 36587 -422 36596
rect -422 36587 -419 36596
rect -381 36587 -354 36596
rect -354 36587 -347 36596
rect -309 36587 -286 36596
rect -286 36587 -275 36596
rect -2829 36527 -2795 36548
rect -2757 36527 -2723 36548
rect -2685 36527 -2651 36548
rect -2613 36527 -2579 36548
rect -2541 36527 -2507 36548
rect -2469 36527 -2435 36548
rect -2397 36527 -2363 36548
rect -2325 36527 -2291 36548
rect -2253 36527 -2219 36548
rect -2181 36527 -2147 36548
rect -2109 36527 -2075 36548
rect -2037 36527 -2003 36548
rect -1965 36527 -1931 36548
rect -1893 36527 -1859 36548
rect -1821 36527 -1787 36548
rect -1749 36527 -1715 36548
rect -1677 36527 -1643 36548
rect -1605 36527 -1571 36548
rect -1533 36527 -1499 36548
rect -1461 36527 -1427 36548
rect -1389 36527 -1355 36548
rect -1317 36527 -1283 36548
rect -1245 36527 -1211 36548
rect -1173 36527 -1139 36548
rect -1101 36527 -1067 36548
rect -1029 36527 -995 36548
rect -957 36527 -923 36548
rect -885 36527 -851 36548
rect -813 36527 -779 36548
rect -741 36527 -707 36548
rect -669 36527 -635 36548
rect -597 36527 -563 36548
rect -525 36527 -491 36548
rect -453 36527 -419 36548
rect -381 36527 -347 36548
rect -309 36527 -275 36548
rect -2829 36514 -2802 36527
rect -2802 36514 -2795 36527
rect -2757 36514 -2734 36527
rect -2734 36514 -2723 36527
rect -2685 36514 -2666 36527
rect -2666 36514 -2651 36527
rect -2613 36514 -2598 36527
rect -2598 36514 -2579 36527
rect -2541 36514 -2530 36527
rect -2530 36514 -2507 36527
rect -2469 36514 -2462 36527
rect -2462 36514 -2435 36527
rect -2397 36514 -2394 36527
rect -2394 36514 -2363 36527
rect -2325 36514 -2292 36527
rect -2292 36514 -2291 36527
rect -2253 36514 -2224 36527
rect -2224 36514 -2219 36527
rect -2181 36514 -2156 36527
rect -2156 36514 -2147 36527
rect -2109 36514 -2088 36527
rect -2088 36514 -2075 36527
rect -2037 36514 -2020 36527
rect -2020 36514 -2003 36527
rect -1965 36514 -1952 36527
rect -1952 36514 -1931 36527
rect -1893 36514 -1884 36527
rect -1884 36514 -1859 36527
rect -1821 36514 -1816 36527
rect -1816 36514 -1787 36527
rect -1749 36514 -1748 36527
rect -1748 36514 -1715 36527
rect -1677 36514 -1646 36527
rect -1646 36514 -1643 36527
rect -1605 36514 -1578 36527
rect -1578 36514 -1571 36527
rect -1533 36514 -1510 36527
rect -1510 36514 -1499 36527
rect -1461 36514 -1442 36527
rect -1442 36514 -1427 36527
rect -1389 36514 -1374 36527
rect -1374 36514 -1355 36527
rect -1317 36514 -1306 36527
rect -1306 36514 -1283 36527
rect -1245 36514 -1238 36527
rect -1238 36514 -1211 36527
rect -1173 36514 -1170 36527
rect -1170 36514 -1139 36527
rect -1101 36514 -1068 36527
rect -1068 36514 -1067 36527
rect -1029 36514 -1000 36527
rect -1000 36514 -995 36527
rect -957 36514 -932 36527
rect -932 36514 -923 36527
rect -885 36514 -864 36527
rect -864 36514 -851 36527
rect -813 36514 -796 36527
rect -796 36514 -779 36527
rect -741 36514 -728 36527
rect -728 36514 -707 36527
rect -669 36514 -660 36527
rect -660 36514 -635 36527
rect -597 36514 -592 36527
rect -592 36514 -563 36527
rect -525 36514 -524 36527
rect -524 36514 -491 36527
rect -453 36514 -422 36527
rect -422 36514 -419 36527
rect -381 36514 -354 36527
rect -354 36514 -347 36527
rect -309 36514 -286 36527
rect -286 36514 -275 36527
rect -2829 36458 -2795 36475
rect -2757 36458 -2723 36475
rect -2685 36458 -2651 36475
rect -2613 36458 -2579 36475
rect -2541 36458 -2507 36475
rect -2469 36458 -2435 36475
rect -2397 36458 -2363 36475
rect -2325 36458 -2291 36475
rect -2253 36458 -2219 36475
rect -2181 36458 -2147 36475
rect -2109 36458 -2075 36475
rect -2037 36458 -2003 36475
rect -1965 36458 -1931 36475
rect -1893 36458 -1859 36475
rect -1821 36458 -1787 36475
rect -1749 36458 -1715 36475
rect -1677 36458 -1643 36475
rect -1605 36458 -1571 36475
rect -1533 36458 -1499 36475
rect -1461 36458 -1427 36475
rect -1389 36458 -1355 36475
rect -1317 36458 -1283 36475
rect -1245 36458 -1211 36475
rect -1173 36458 -1139 36475
rect -1101 36458 -1067 36475
rect -1029 36458 -995 36475
rect -957 36458 -923 36475
rect -885 36458 -851 36475
rect -813 36458 -779 36475
rect -741 36458 -707 36475
rect -669 36458 -635 36475
rect -597 36458 -563 36475
rect -525 36458 -491 36475
rect -453 36458 -419 36475
rect -381 36458 -347 36475
rect -309 36458 -275 36475
rect -2829 36441 -2802 36458
rect -2802 36441 -2795 36458
rect -2757 36441 -2734 36458
rect -2734 36441 -2723 36458
rect -2685 36441 -2666 36458
rect -2666 36441 -2651 36458
rect -2613 36441 -2598 36458
rect -2598 36441 -2579 36458
rect -2541 36441 -2530 36458
rect -2530 36441 -2507 36458
rect -2469 36441 -2462 36458
rect -2462 36441 -2435 36458
rect -2397 36441 -2394 36458
rect -2394 36441 -2363 36458
rect -2325 36441 -2292 36458
rect -2292 36441 -2291 36458
rect -2253 36441 -2224 36458
rect -2224 36441 -2219 36458
rect -2181 36441 -2156 36458
rect -2156 36441 -2147 36458
rect -2109 36441 -2088 36458
rect -2088 36441 -2075 36458
rect -2037 36441 -2020 36458
rect -2020 36441 -2003 36458
rect -1965 36441 -1952 36458
rect -1952 36441 -1931 36458
rect -1893 36441 -1884 36458
rect -1884 36441 -1859 36458
rect -1821 36441 -1816 36458
rect -1816 36441 -1787 36458
rect -1749 36441 -1748 36458
rect -1748 36441 -1715 36458
rect -1677 36441 -1646 36458
rect -1646 36441 -1643 36458
rect -1605 36441 -1578 36458
rect -1578 36441 -1571 36458
rect -1533 36441 -1510 36458
rect -1510 36441 -1499 36458
rect -1461 36441 -1442 36458
rect -1442 36441 -1427 36458
rect -1389 36441 -1374 36458
rect -1374 36441 -1355 36458
rect -1317 36441 -1306 36458
rect -1306 36441 -1283 36458
rect -1245 36441 -1238 36458
rect -1238 36441 -1211 36458
rect -1173 36441 -1170 36458
rect -1170 36441 -1139 36458
rect -1101 36441 -1068 36458
rect -1068 36441 -1067 36458
rect -1029 36441 -1000 36458
rect -1000 36441 -995 36458
rect -957 36441 -932 36458
rect -932 36441 -923 36458
rect -885 36441 -864 36458
rect -864 36441 -851 36458
rect -813 36441 -796 36458
rect -796 36441 -779 36458
rect -741 36441 -728 36458
rect -728 36441 -707 36458
rect -669 36441 -660 36458
rect -660 36441 -635 36458
rect -597 36441 -592 36458
rect -592 36441 -563 36458
rect -525 36441 -524 36458
rect -524 36441 -491 36458
rect -453 36441 -422 36458
rect -422 36441 -419 36458
rect -381 36441 -354 36458
rect -354 36441 -347 36458
rect -309 36441 -286 36458
rect -286 36441 -275 36458
rect -2829 36389 -2795 36402
rect -2757 36389 -2723 36402
rect -2685 36389 -2651 36402
rect -2613 36389 -2579 36402
rect -2541 36389 -2507 36402
rect -2469 36389 -2435 36402
rect -2397 36389 -2363 36402
rect -2325 36389 -2291 36402
rect -2253 36389 -2219 36402
rect -2181 36389 -2147 36402
rect -2109 36389 -2075 36402
rect -2037 36389 -2003 36402
rect -1965 36389 -1931 36402
rect -1893 36389 -1859 36402
rect -1821 36389 -1787 36402
rect -1749 36389 -1715 36402
rect -1677 36389 -1643 36402
rect -1605 36389 -1571 36402
rect -1533 36389 -1499 36402
rect -1461 36389 -1427 36402
rect -1389 36389 -1355 36402
rect -1317 36389 -1283 36402
rect -1245 36389 -1211 36402
rect -1173 36389 -1139 36402
rect -1101 36389 -1067 36402
rect -1029 36389 -995 36402
rect -957 36389 -923 36402
rect -885 36389 -851 36402
rect -813 36389 -779 36402
rect -741 36389 -707 36402
rect -669 36389 -635 36402
rect -597 36389 -563 36402
rect -525 36389 -491 36402
rect -453 36389 -419 36402
rect -381 36389 -347 36402
rect -309 36389 -275 36402
rect -2829 36368 -2802 36389
rect -2802 36368 -2795 36389
rect -2757 36368 -2734 36389
rect -2734 36368 -2723 36389
rect -2685 36368 -2666 36389
rect -2666 36368 -2651 36389
rect -2613 36368 -2598 36389
rect -2598 36368 -2579 36389
rect -2541 36368 -2530 36389
rect -2530 36368 -2507 36389
rect -2469 36368 -2462 36389
rect -2462 36368 -2435 36389
rect -2397 36368 -2394 36389
rect -2394 36368 -2363 36389
rect -2325 36368 -2292 36389
rect -2292 36368 -2291 36389
rect -2253 36368 -2224 36389
rect -2224 36368 -2219 36389
rect -2181 36368 -2156 36389
rect -2156 36368 -2147 36389
rect -2109 36368 -2088 36389
rect -2088 36368 -2075 36389
rect -2037 36368 -2020 36389
rect -2020 36368 -2003 36389
rect -1965 36368 -1952 36389
rect -1952 36368 -1931 36389
rect -1893 36368 -1884 36389
rect -1884 36368 -1859 36389
rect -1821 36368 -1816 36389
rect -1816 36368 -1787 36389
rect -1749 36368 -1748 36389
rect -1748 36368 -1715 36389
rect -1677 36368 -1646 36389
rect -1646 36368 -1643 36389
rect -1605 36368 -1578 36389
rect -1578 36368 -1571 36389
rect -1533 36368 -1510 36389
rect -1510 36368 -1499 36389
rect -1461 36368 -1442 36389
rect -1442 36368 -1427 36389
rect -1389 36368 -1374 36389
rect -1374 36368 -1355 36389
rect -1317 36368 -1306 36389
rect -1306 36368 -1283 36389
rect -1245 36368 -1238 36389
rect -1238 36368 -1211 36389
rect -1173 36368 -1170 36389
rect -1170 36368 -1139 36389
rect -1101 36368 -1068 36389
rect -1068 36368 -1067 36389
rect -1029 36368 -1000 36389
rect -1000 36368 -995 36389
rect -957 36368 -932 36389
rect -932 36368 -923 36389
rect -885 36368 -864 36389
rect -864 36368 -851 36389
rect -813 36368 -796 36389
rect -796 36368 -779 36389
rect -741 36368 -728 36389
rect -728 36368 -707 36389
rect -669 36368 -660 36389
rect -660 36368 -635 36389
rect -597 36368 -592 36389
rect -592 36368 -563 36389
rect -525 36368 -524 36389
rect -524 36368 -491 36389
rect -453 36368 -422 36389
rect -422 36368 -419 36389
rect -381 36368 -354 36389
rect -354 36368 -347 36389
rect -309 36368 -286 36389
rect -286 36368 -275 36389
rect -2829 36320 -2795 36329
rect -2757 36320 -2723 36329
rect -2685 36320 -2651 36329
rect -2613 36320 -2579 36329
rect -2541 36320 -2507 36329
rect -2469 36320 -2435 36329
rect -2397 36320 -2363 36329
rect -2325 36320 -2291 36329
rect -2253 36320 -2219 36329
rect -2181 36320 -2147 36329
rect -2109 36320 -2075 36329
rect -2037 36320 -2003 36329
rect -1965 36320 -1931 36329
rect -1893 36320 -1859 36329
rect -1821 36320 -1787 36329
rect -1749 36320 -1715 36329
rect -1677 36320 -1643 36329
rect -1605 36320 -1571 36329
rect -1533 36320 -1499 36329
rect -1461 36320 -1427 36329
rect -1389 36320 -1355 36329
rect -1317 36320 -1283 36329
rect -1245 36320 -1211 36329
rect -1173 36320 -1139 36329
rect -1101 36320 -1067 36329
rect -1029 36320 -995 36329
rect -957 36320 -923 36329
rect -885 36320 -851 36329
rect -813 36320 -779 36329
rect -741 36320 -707 36329
rect -669 36320 -635 36329
rect -597 36320 -563 36329
rect -525 36320 -491 36329
rect -453 36320 -419 36329
rect -381 36320 -347 36329
rect -309 36320 -275 36329
rect -2829 36295 -2802 36320
rect -2802 36295 -2795 36320
rect -2757 36295 -2734 36320
rect -2734 36295 -2723 36320
rect -2685 36295 -2666 36320
rect -2666 36295 -2651 36320
rect -2613 36295 -2598 36320
rect -2598 36295 -2579 36320
rect -2541 36295 -2530 36320
rect -2530 36295 -2507 36320
rect -2469 36295 -2462 36320
rect -2462 36295 -2435 36320
rect -2397 36295 -2394 36320
rect -2394 36295 -2363 36320
rect -2325 36295 -2292 36320
rect -2292 36295 -2291 36320
rect -2253 36295 -2224 36320
rect -2224 36295 -2219 36320
rect -2181 36295 -2156 36320
rect -2156 36295 -2147 36320
rect -2109 36295 -2088 36320
rect -2088 36295 -2075 36320
rect -2037 36295 -2020 36320
rect -2020 36295 -2003 36320
rect -1965 36295 -1952 36320
rect -1952 36295 -1931 36320
rect -1893 36295 -1884 36320
rect -1884 36295 -1859 36320
rect -1821 36295 -1816 36320
rect -1816 36295 -1787 36320
rect -1749 36295 -1748 36320
rect -1748 36295 -1715 36320
rect -1677 36295 -1646 36320
rect -1646 36295 -1643 36320
rect -1605 36295 -1578 36320
rect -1578 36295 -1571 36320
rect -1533 36295 -1510 36320
rect -1510 36295 -1499 36320
rect -1461 36295 -1442 36320
rect -1442 36295 -1427 36320
rect -1389 36295 -1374 36320
rect -1374 36295 -1355 36320
rect -1317 36295 -1306 36320
rect -1306 36295 -1283 36320
rect -1245 36295 -1238 36320
rect -1238 36295 -1211 36320
rect -1173 36295 -1170 36320
rect -1170 36295 -1139 36320
rect -1101 36295 -1068 36320
rect -1068 36295 -1067 36320
rect -1029 36295 -1000 36320
rect -1000 36295 -995 36320
rect -957 36295 -932 36320
rect -932 36295 -923 36320
rect -885 36295 -864 36320
rect -864 36295 -851 36320
rect -813 36295 -796 36320
rect -796 36295 -779 36320
rect -741 36295 -728 36320
rect -728 36295 -707 36320
rect -669 36295 -660 36320
rect -660 36295 -635 36320
rect -597 36295 -592 36320
rect -592 36295 -563 36320
rect -525 36295 -524 36320
rect -524 36295 -491 36320
rect -453 36295 -422 36320
rect -422 36295 -419 36320
rect -381 36295 -354 36320
rect -354 36295 -347 36320
rect -309 36295 -286 36320
rect -286 36295 -275 36320
rect -2829 36251 -2795 36256
rect -2757 36251 -2723 36256
rect -2685 36251 -2651 36256
rect -2613 36251 -2579 36256
rect -2541 36251 -2507 36256
rect -2469 36251 -2435 36256
rect -2397 36251 -2363 36256
rect -2325 36251 -2291 36256
rect -2253 36251 -2219 36256
rect -2181 36251 -2147 36256
rect -2109 36251 -2075 36256
rect -2037 36251 -2003 36256
rect -1965 36251 -1931 36256
rect -1893 36251 -1859 36256
rect -1821 36251 -1787 36256
rect -1749 36251 -1715 36256
rect -1677 36251 -1643 36256
rect -1605 36251 -1571 36256
rect -1533 36251 -1499 36256
rect -1461 36251 -1427 36256
rect -1389 36251 -1355 36256
rect -1317 36251 -1283 36256
rect -1245 36251 -1211 36256
rect -1173 36251 -1139 36256
rect -1101 36251 -1067 36256
rect -1029 36251 -995 36256
rect -957 36251 -923 36256
rect -885 36251 -851 36256
rect -813 36251 -779 36256
rect -741 36251 -707 36256
rect -669 36251 -635 36256
rect -597 36251 -563 36256
rect -525 36251 -491 36256
rect -453 36251 -419 36256
rect -381 36251 -347 36256
rect -309 36251 -275 36256
rect -2829 36222 -2802 36251
rect -2802 36222 -2795 36251
rect -2757 36222 -2734 36251
rect -2734 36222 -2723 36251
rect -2685 36222 -2666 36251
rect -2666 36222 -2651 36251
rect -2613 36222 -2598 36251
rect -2598 36222 -2579 36251
rect -2541 36222 -2530 36251
rect -2530 36222 -2507 36251
rect -2469 36222 -2462 36251
rect -2462 36222 -2435 36251
rect -2397 36222 -2394 36251
rect -2394 36222 -2363 36251
rect -2325 36222 -2292 36251
rect -2292 36222 -2291 36251
rect -2253 36222 -2224 36251
rect -2224 36222 -2219 36251
rect -2181 36222 -2156 36251
rect -2156 36222 -2147 36251
rect -2109 36222 -2088 36251
rect -2088 36222 -2075 36251
rect -2037 36222 -2020 36251
rect -2020 36222 -2003 36251
rect -1965 36222 -1952 36251
rect -1952 36222 -1931 36251
rect -1893 36222 -1884 36251
rect -1884 36222 -1859 36251
rect -1821 36222 -1816 36251
rect -1816 36222 -1787 36251
rect -1749 36222 -1748 36251
rect -1748 36222 -1715 36251
rect -1677 36222 -1646 36251
rect -1646 36222 -1643 36251
rect -1605 36222 -1578 36251
rect -1578 36222 -1571 36251
rect -1533 36222 -1510 36251
rect -1510 36222 -1499 36251
rect -1461 36222 -1442 36251
rect -1442 36222 -1427 36251
rect -1389 36222 -1374 36251
rect -1374 36222 -1355 36251
rect -1317 36222 -1306 36251
rect -1306 36222 -1283 36251
rect -1245 36222 -1238 36251
rect -1238 36222 -1211 36251
rect -1173 36222 -1170 36251
rect -1170 36222 -1139 36251
rect -1101 36222 -1068 36251
rect -1068 36222 -1067 36251
rect -1029 36222 -1000 36251
rect -1000 36222 -995 36251
rect -957 36222 -932 36251
rect -932 36222 -923 36251
rect -885 36222 -864 36251
rect -864 36222 -851 36251
rect -813 36222 -796 36251
rect -796 36222 -779 36251
rect -741 36222 -728 36251
rect -728 36222 -707 36251
rect -669 36222 -660 36251
rect -660 36222 -635 36251
rect -597 36222 -592 36251
rect -592 36222 -563 36251
rect -525 36222 -524 36251
rect -524 36222 -491 36251
rect -453 36222 -422 36251
rect -422 36222 -419 36251
rect -381 36222 -354 36251
rect -354 36222 -347 36251
rect -309 36222 -286 36251
rect -286 36222 -275 36251
rect -2829 36182 -2795 36183
rect -2757 36182 -2723 36183
rect -2685 36182 -2651 36183
rect -2613 36182 -2579 36183
rect -2541 36182 -2507 36183
rect -2469 36182 -2435 36183
rect -2397 36182 -2363 36183
rect -2325 36182 -2291 36183
rect -2253 36182 -2219 36183
rect -2181 36182 -2147 36183
rect -2109 36182 -2075 36183
rect -2037 36182 -2003 36183
rect -1965 36182 -1931 36183
rect -1893 36182 -1859 36183
rect -1821 36182 -1787 36183
rect -1749 36182 -1715 36183
rect -1677 36182 -1643 36183
rect -1605 36182 -1571 36183
rect -1533 36182 -1499 36183
rect -1461 36182 -1427 36183
rect -1389 36182 -1355 36183
rect -1317 36182 -1283 36183
rect -1245 36182 -1211 36183
rect -1173 36182 -1139 36183
rect -1101 36182 -1067 36183
rect -1029 36182 -995 36183
rect -957 36182 -923 36183
rect -885 36182 -851 36183
rect -813 36182 -779 36183
rect -741 36182 -707 36183
rect -669 36182 -635 36183
rect -597 36182 -563 36183
rect -525 36182 -491 36183
rect -453 36182 -419 36183
rect -381 36182 -347 36183
rect -309 36182 -275 36183
rect -2829 36149 -2802 36182
rect -2802 36149 -2795 36182
rect -2757 36149 -2734 36182
rect -2734 36149 -2723 36182
rect -2685 36149 -2666 36182
rect -2666 36149 -2651 36182
rect -2613 36149 -2598 36182
rect -2598 36149 -2579 36182
rect -2541 36149 -2530 36182
rect -2530 36149 -2507 36182
rect -2469 36149 -2462 36182
rect -2462 36149 -2435 36182
rect -2397 36149 -2394 36182
rect -2394 36149 -2363 36182
rect -2325 36149 -2292 36182
rect -2292 36149 -2291 36182
rect -2253 36149 -2224 36182
rect -2224 36149 -2219 36182
rect -2181 36149 -2156 36182
rect -2156 36149 -2147 36182
rect -2109 36149 -2088 36182
rect -2088 36149 -2075 36182
rect -2037 36149 -2020 36182
rect -2020 36149 -2003 36182
rect -1965 36149 -1952 36182
rect -1952 36149 -1931 36182
rect -1893 36149 -1884 36182
rect -1884 36149 -1859 36182
rect -1821 36149 -1816 36182
rect -1816 36149 -1787 36182
rect -1749 36149 -1748 36182
rect -1748 36149 -1715 36182
rect -1677 36149 -1646 36182
rect -1646 36149 -1643 36182
rect -1605 36149 -1578 36182
rect -1578 36149 -1571 36182
rect -1533 36149 -1510 36182
rect -1510 36149 -1499 36182
rect -1461 36149 -1442 36182
rect -1442 36149 -1427 36182
rect -1389 36149 -1374 36182
rect -1374 36149 -1355 36182
rect -1317 36149 -1306 36182
rect -1306 36149 -1283 36182
rect -1245 36149 -1238 36182
rect -1238 36149 -1211 36182
rect -1173 36149 -1170 36182
rect -1170 36149 -1139 36182
rect -1101 36149 -1068 36182
rect -1068 36149 -1067 36182
rect -1029 36149 -1000 36182
rect -1000 36149 -995 36182
rect -957 36149 -932 36182
rect -932 36149 -923 36182
rect -885 36149 -864 36182
rect -864 36149 -851 36182
rect -813 36149 -796 36182
rect -796 36149 -779 36182
rect -741 36149 -728 36182
rect -728 36149 -707 36182
rect -669 36149 -660 36182
rect -660 36149 -635 36182
rect -597 36149 -592 36182
rect -592 36149 -563 36182
rect -525 36149 -524 36182
rect -524 36149 -491 36182
rect -453 36149 -422 36182
rect -422 36149 -419 36182
rect -381 36149 -354 36182
rect -354 36149 -347 36182
rect -309 36149 -286 36182
rect -286 36149 -275 36182
rect -2829 36079 -2802 36110
rect -2802 36079 -2795 36110
rect -2757 36079 -2734 36110
rect -2734 36079 -2723 36110
rect -2685 36079 -2666 36110
rect -2666 36079 -2651 36110
rect -2613 36079 -2598 36110
rect -2598 36079 -2579 36110
rect -2541 36079 -2530 36110
rect -2530 36079 -2507 36110
rect -2469 36079 -2462 36110
rect -2462 36079 -2435 36110
rect -2397 36079 -2394 36110
rect -2394 36079 -2363 36110
rect -2325 36079 -2292 36110
rect -2292 36079 -2291 36110
rect -2253 36079 -2224 36110
rect -2224 36079 -2219 36110
rect -2181 36079 -2156 36110
rect -2156 36079 -2147 36110
rect -2109 36079 -2088 36110
rect -2088 36079 -2075 36110
rect -2037 36079 -2020 36110
rect -2020 36079 -2003 36110
rect -1965 36079 -1952 36110
rect -1952 36079 -1931 36110
rect -1893 36079 -1884 36110
rect -1884 36079 -1859 36110
rect -1821 36079 -1816 36110
rect -1816 36079 -1787 36110
rect -1749 36079 -1748 36110
rect -1748 36079 -1715 36110
rect -1677 36079 -1646 36110
rect -1646 36079 -1643 36110
rect -1605 36079 -1578 36110
rect -1578 36079 -1571 36110
rect -1533 36079 -1510 36110
rect -1510 36079 -1499 36110
rect -1461 36079 -1442 36110
rect -1442 36079 -1427 36110
rect -1389 36079 -1374 36110
rect -1374 36079 -1355 36110
rect -1317 36079 -1306 36110
rect -1306 36079 -1283 36110
rect -1245 36079 -1238 36110
rect -1238 36079 -1211 36110
rect -1173 36079 -1170 36110
rect -1170 36079 -1139 36110
rect -1101 36079 -1068 36110
rect -1068 36079 -1067 36110
rect -1029 36079 -1000 36110
rect -1000 36079 -995 36110
rect -957 36079 -932 36110
rect -932 36079 -923 36110
rect -885 36079 -864 36110
rect -864 36079 -851 36110
rect -813 36079 -796 36110
rect -796 36079 -779 36110
rect -741 36079 -728 36110
rect -728 36079 -707 36110
rect -669 36079 -660 36110
rect -660 36079 -635 36110
rect -597 36079 -592 36110
rect -592 36079 -563 36110
rect -525 36079 -524 36110
rect -524 36079 -491 36110
rect -453 36079 -422 36110
rect -422 36079 -419 36110
rect -381 36079 -354 36110
rect -354 36079 -347 36110
rect -309 36079 -286 36110
rect -286 36079 -275 36110
rect -2829 36076 -2795 36079
rect -2757 36076 -2723 36079
rect -2685 36076 -2651 36079
rect -2613 36076 -2579 36079
rect -2541 36076 -2507 36079
rect -2469 36076 -2435 36079
rect -2397 36076 -2363 36079
rect -2325 36076 -2291 36079
rect -2253 36076 -2219 36079
rect -2181 36076 -2147 36079
rect -2109 36076 -2075 36079
rect -2037 36076 -2003 36079
rect -1965 36076 -1931 36079
rect -1893 36076 -1859 36079
rect -1821 36076 -1787 36079
rect -1749 36076 -1715 36079
rect -1677 36076 -1643 36079
rect -1605 36076 -1571 36079
rect -1533 36076 -1499 36079
rect -1461 36076 -1427 36079
rect -1389 36076 -1355 36079
rect -1317 36076 -1283 36079
rect -1245 36076 -1211 36079
rect -1173 36076 -1139 36079
rect -1101 36076 -1067 36079
rect -1029 36076 -995 36079
rect -957 36076 -923 36079
rect -885 36076 -851 36079
rect -813 36076 -779 36079
rect -741 36076 -707 36079
rect -669 36076 -635 36079
rect -597 36076 -563 36079
rect -525 36076 -491 36079
rect -453 36076 -419 36079
rect -381 36076 -347 36079
rect -309 36076 -275 36079
rect -2829 36010 -2802 36037
rect -2802 36010 -2795 36037
rect -2757 36010 -2734 36037
rect -2734 36010 -2723 36037
rect -2685 36010 -2666 36037
rect -2666 36010 -2651 36037
rect -2613 36010 -2598 36037
rect -2598 36010 -2579 36037
rect -2541 36010 -2530 36037
rect -2530 36010 -2507 36037
rect -2469 36010 -2462 36037
rect -2462 36010 -2435 36037
rect -2397 36010 -2394 36037
rect -2394 36010 -2363 36037
rect -2325 36010 -2292 36037
rect -2292 36010 -2291 36037
rect -2253 36010 -2224 36037
rect -2224 36010 -2219 36037
rect -2181 36010 -2156 36037
rect -2156 36010 -2147 36037
rect -2109 36010 -2088 36037
rect -2088 36010 -2075 36037
rect -2037 36010 -2020 36037
rect -2020 36010 -2003 36037
rect -1965 36010 -1952 36037
rect -1952 36010 -1931 36037
rect -1893 36010 -1884 36037
rect -1884 36010 -1859 36037
rect -1821 36010 -1816 36037
rect -1816 36010 -1787 36037
rect -1749 36010 -1748 36037
rect -1748 36010 -1715 36037
rect -1677 36010 -1646 36037
rect -1646 36010 -1643 36037
rect -1605 36010 -1578 36037
rect -1578 36010 -1571 36037
rect -1533 36010 -1510 36037
rect -1510 36010 -1499 36037
rect -1461 36010 -1442 36037
rect -1442 36010 -1427 36037
rect -1389 36010 -1374 36037
rect -1374 36010 -1355 36037
rect -1317 36010 -1306 36037
rect -1306 36010 -1283 36037
rect -1245 36010 -1238 36037
rect -1238 36010 -1211 36037
rect -1173 36010 -1170 36037
rect -1170 36010 -1139 36037
rect -1101 36010 -1068 36037
rect -1068 36010 -1067 36037
rect -1029 36010 -1000 36037
rect -1000 36010 -995 36037
rect -957 36010 -932 36037
rect -932 36010 -923 36037
rect -885 36010 -864 36037
rect -864 36010 -851 36037
rect -813 36010 -796 36037
rect -796 36010 -779 36037
rect -741 36010 -728 36037
rect -728 36010 -707 36037
rect -669 36010 -660 36037
rect -660 36010 -635 36037
rect -597 36010 -592 36037
rect -592 36010 -563 36037
rect -525 36010 -524 36037
rect -524 36010 -491 36037
rect -453 36010 -422 36037
rect -422 36010 -419 36037
rect -381 36010 -354 36037
rect -354 36010 -347 36037
rect -309 36010 -286 36037
rect -286 36010 -275 36037
rect -2829 36003 -2795 36010
rect -2757 36003 -2723 36010
rect -2685 36003 -2651 36010
rect -2613 36003 -2579 36010
rect -2541 36003 -2507 36010
rect -2469 36003 -2435 36010
rect -2397 36003 -2363 36010
rect -2325 36003 -2291 36010
rect -2253 36003 -2219 36010
rect -2181 36003 -2147 36010
rect -2109 36003 -2075 36010
rect -2037 36003 -2003 36010
rect -1965 36003 -1931 36010
rect -1893 36003 -1859 36010
rect -1821 36003 -1787 36010
rect -1749 36003 -1715 36010
rect -1677 36003 -1643 36010
rect -1605 36003 -1571 36010
rect -1533 36003 -1499 36010
rect -1461 36003 -1427 36010
rect -1389 36003 -1355 36010
rect -1317 36003 -1283 36010
rect -1245 36003 -1211 36010
rect -1173 36003 -1139 36010
rect -1101 36003 -1067 36010
rect -1029 36003 -995 36010
rect -957 36003 -923 36010
rect -885 36003 -851 36010
rect -813 36003 -779 36010
rect -741 36003 -707 36010
rect -669 36003 -635 36010
rect -597 36003 -563 36010
rect -525 36003 -491 36010
rect -453 36003 -419 36010
rect -381 36003 -347 36010
rect -309 36003 -275 36010
rect -2829 35941 -2802 35964
rect -2802 35941 -2795 35964
rect -2757 35941 -2734 35964
rect -2734 35941 -2723 35964
rect -2685 35941 -2666 35964
rect -2666 35941 -2651 35964
rect -2613 35941 -2598 35964
rect -2598 35941 -2579 35964
rect -2541 35941 -2530 35964
rect -2530 35941 -2507 35964
rect -2469 35941 -2462 35964
rect -2462 35941 -2435 35964
rect -2397 35941 -2394 35964
rect -2394 35941 -2363 35964
rect -2325 35941 -2292 35964
rect -2292 35941 -2291 35964
rect -2253 35941 -2224 35964
rect -2224 35941 -2219 35964
rect -2181 35941 -2156 35964
rect -2156 35941 -2147 35964
rect -2109 35941 -2088 35964
rect -2088 35941 -2075 35964
rect -2037 35941 -2020 35964
rect -2020 35941 -2003 35964
rect -1965 35941 -1952 35964
rect -1952 35941 -1931 35964
rect -1893 35941 -1884 35964
rect -1884 35941 -1859 35964
rect -1821 35941 -1816 35964
rect -1816 35941 -1787 35964
rect -1749 35941 -1748 35964
rect -1748 35941 -1715 35964
rect -1677 35941 -1646 35964
rect -1646 35941 -1643 35964
rect -1605 35941 -1578 35964
rect -1578 35941 -1571 35964
rect -1533 35941 -1510 35964
rect -1510 35941 -1499 35964
rect -1461 35941 -1442 35964
rect -1442 35941 -1427 35964
rect -1389 35941 -1374 35964
rect -1374 35941 -1355 35964
rect -1317 35941 -1306 35964
rect -1306 35941 -1283 35964
rect -1245 35941 -1238 35964
rect -1238 35941 -1211 35964
rect -1173 35941 -1170 35964
rect -1170 35941 -1139 35964
rect -1101 35941 -1068 35964
rect -1068 35941 -1067 35964
rect -1029 35941 -1000 35964
rect -1000 35941 -995 35964
rect -957 35941 -932 35964
rect -932 35941 -923 35964
rect -885 35941 -864 35964
rect -864 35941 -851 35964
rect -813 35941 -796 35964
rect -796 35941 -779 35964
rect -741 35941 -728 35964
rect -728 35941 -707 35964
rect -669 35941 -660 35964
rect -660 35941 -635 35964
rect -597 35941 -592 35964
rect -592 35941 -563 35964
rect -525 35941 -524 35964
rect -524 35941 -491 35964
rect -453 35941 -422 35964
rect -422 35941 -419 35964
rect -381 35941 -354 35964
rect -354 35941 -347 35964
rect -309 35941 -286 35964
rect -286 35941 -275 35964
rect -2829 35930 -2795 35941
rect -2757 35930 -2723 35941
rect -2685 35930 -2651 35941
rect -2613 35930 -2579 35941
rect -2541 35930 -2507 35941
rect -2469 35930 -2435 35941
rect -2397 35930 -2363 35941
rect -2325 35930 -2291 35941
rect -2253 35930 -2219 35941
rect -2181 35930 -2147 35941
rect -2109 35930 -2075 35941
rect -2037 35930 -2003 35941
rect -1965 35930 -1931 35941
rect -1893 35930 -1859 35941
rect -1821 35930 -1787 35941
rect -1749 35930 -1715 35941
rect -1677 35930 -1643 35941
rect -1605 35930 -1571 35941
rect -1533 35930 -1499 35941
rect -1461 35930 -1427 35941
rect -1389 35930 -1355 35941
rect -1317 35930 -1283 35941
rect -1245 35930 -1211 35941
rect -1173 35930 -1139 35941
rect -1101 35930 -1067 35941
rect -1029 35930 -995 35941
rect -957 35930 -923 35941
rect -885 35930 -851 35941
rect -813 35930 -779 35941
rect -741 35930 -707 35941
rect -669 35930 -635 35941
rect -597 35930 -563 35941
rect -525 35930 -491 35941
rect -453 35930 -419 35941
rect -381 35930 -347 35941
rect -309 35930 -275 35941
rect -2829 35872 -2802 35891
rect -2802 35872 -2795 35891
rect -2757 35872 -2734 35891
rect -2734 35872 -2723 35891
rect -2685 35872 -2666 35891
rect -2666 35872 -2651 35891
rect -2613 35872 -2598 35891
rect -2598 35872 -2579 35891
rect -2541 35872 -2530 35891
rect -2530 35872 -2507 35891
rect -2469 35872 -2462 35891
rect -2462 35872 -2435 35891
rect -2397 35872 -2394 35891
rect -2394 35872 -2363 35891
rect -2325 35872 -2292 35891
rect -2292 35872 -2291 35891
rect -2253 35872 -2224 35891
rect -2224 35872 -2219 35891
rect -2181 35872 -2156 35891
rect -2156 35872 -2147 35891
rect -2109 35872 -2088 35891
rect -2088 35872 -2075 35891
rect -2037 35872 -2020 35891
rect -2020 35872 -2003 35891
rect -1965 35872 -1952 35891
rect -1952 35872 -1931 35891
rect -1893 35872 -1884 35891
rect -1884 35872 -1859 35891
rect -1821 35872 -1816 35891
rect -1816 35872 -1787 35891
rect -1749 35872 -1748 35891
rect -1748 35872 -1715 35891
rect -1677 35872 -1646 35891
rect -1646 35872 -1643 35891
rect -1605 35872 -1578 35891
rect -1578 35872 -1571 35891
rect -1533 35872 -1510 35891
rect -1510 35872 -1499 35891
rect -1461 35872 -1442 35891
rect -1442 35872 -1427 35891
rect -1389 35872 -1374 35891
rect -1374 35872 -1355 35891
rect -1317 35872 -1306 35891
rect -1306 35872 -1283 35891
rect -1245 35872 -1238 35891
rect -1238 35872 -1211 35891
rect -1173 35872 -1170 35891
rect -1170 35872 -1139 35891
rect -1101 35872 -1068 35891
rect -1068 35872 -1067 35891
rect -1029 35872 -1000 35891
rect -1000 35872 -995 35891
rect -957 35872 -932 35891
rect -932 35872 -923 35891
rect -885 35872 -864 35891
rect -864 35872 -851 35891
rect -813 35872 -796 35891
rect -796 35872 -779 35891
rect -741 35872 -728 35891
rect -728 35872 -707 35891
rect -669 35872 -660 35891
rect -660 35872 -635 35891
rect -597 35872 -592 35891
rect -592 35872 -563 35891
rect -525 35872 -524 35891
rect -524 35872 -491 35891
rect -453 35872 -422 35891
rect -422 35872 -419 35891
rect -381 35872 -354 35891
rect -354 35872 -347 35891
rect -309 35872 -286 35891
rect -286 35872 -275 35891
rect -2829 35857 -2795 35872
rect -2757 35857 -2723 35872
rect -2685 35857 -2651 35872
rect -2613 35857 -2579 35872
rect -2541 35857 -2507 35872
rect -2469 35857 -2435 35872
rect -2397 35857 -2363 35872
rect -2325 35857 -2291 35872
rect -2253 35857 -2219 35872
rect -2181 35857 -2147 35872
rect -2109 35857 -2075 35872
rect -2037 35857 -2003 35872
rect -1965 35857 -1931 35872
rect -1893 35857 -1859 35872
rect -1821 35857 -1787 35872
rect -1749 35857 -1715 35872
rect -1677 35857 -1643 35872
rect -1605 35857 -1571 35872
rect -1533 35857 -1499 35872
rect -1461 35857 -1427 35872
rect -1389 35857 -1355 35872
rect -1317 35857 -1283 35872
rect -1245 35857 -1211 35872
rect -1173 35857 -1139 35872
rect -1101 35857 -1067 35872
rect -1029 35857 -995 35872
rect -957 35857 -923 35872
rect -885 35857 -851 35872
rect -813 35857 -779 35872
rect -741 35857 -707 35872
rect -669 35857 -635 35872
rect -597 35857 -563 35872
rect -525 35857 -491 35872
rect -453 35857 -419 35872
rect -381 35857 -347 35872
rect -309 35857 -275 35872
rect -2829 35803 -2802 35818
rect -2802 35803 -2795 35818
rect -2757 35803 -2734 35818
rect -2734 35803 -2723 35818
rect -2685 35803 -2666 35818
rect -2666 35803 -2651 35818
rect -2613 35803 -2598 35818
rect -2598 35803 -2579 35818
rect -2541 35803 -2530 35818
rect -2530 35803 -2507 35818
rect -2469 35803 -2462 35818
rect -2462 35803 -2435 35818
rect -2397 35803 -2394 35818
rect -2394 35803 -2363 35818
rect -2325 35803 -2292 35818
rect -2292 35803 -2291 35818
rect -2253 35803 -2224 35818
rect -2224 35803 -2219 35818
rect -2181 35803 -2156 35818
rect -2156 35803 -2147 35818
rect -2109 35803 -2088 35818
rect -2088 35803 -2075 35818
rect -2037 35803 -2020 35818
rect -2020 35803 -2003 35818
rect -1965 35803 -1952 35818
rect -1952 35803 -1931 35818
rect -1893 35803 -1884 35818
rect -1884 35803 -1859 35818
rect -1821 35803 -1816 35818
rect -1816 35803 -1787 35818
rect -1749 35803 -1748 35818
rect -1748 35803 -1715 35818
rect -1677 35803 -1646 35818
rect -1646 35803 -1643 35818
rect -1605 35803 -1578 35818
rect -1578 35803 -1571 35818
rect -1533 35803 -1510 35818
rect -1510 35803 -1499 35818
rect -1461 35803 -1442 35818
rect -1442 35803 -1427 35818
rect -1389 35803 -1374 35818
rect -1374 35803 -1355 35818
rect -1317 35803 -1306 35818
rect -1306 35803 -1283 35818
rect -1245 35803 -1238 35818
rect -1238 35803 -1211 35818
rect -1173 35803 -1170 35818
rect -1170 35803 -1139 35818
rect -1101 35803 -1068 35818
rect -1068 35803 -1067 35818
rect -1029 35803 -1000 35818
rect -1000 35803 -995 35818
rect -957 35803 -932 35818
rect -932 35803 -923 35818
rect -885 35803 -864 35818
rect -864 35803 -851 35818
rect -813 35803 -796 35818
rect -796 35803 -779 35818
rect -741 35803 -728 35818
rect -728 35803 -707 35818
rect -669 35803 -660 35818
rect -660 35803 -635 35818
rect -597 35803 -592 35818
rect -592 35803 -563 35818
rect -525 35803 -524 35818
rect -524 35803 -491 35818
rect -453 35803 -422 35818
rect -422 35803 -419 35818
rect -381 35803 -354 35818
rect -354 35803 -347 35818
rect -309 35803 -286 35818
rect -286 35803 -275 35818
rect -2829 35784 -2795 35803
rect -2757 35784 -2723 35803
rect -2685 35784 -2651 35803
rect -2613 35784 -2579 35803
rect -2541 35784 -2507 35803
rect -2469 35784 -2435 35803
rect -2397 35784 -2363 35803
rect -2325 35784 -2291 35803
rect -2253 35784 -2219 35803
rect -2181 35784 -2147 35803
rect -2109 35784 -2075 35803
rect -2037 35784 -2003 35803
rect -1965 35784 -1931 35803
rect -1893 35784 -1859 35803
rect -1821 35784 -1787 35803
rect -1749 35784 -1715 35803
rect -1677 35784 -1643 35803
rect -1605 35784 -1571 35803
rect -1533 35784 -1499 35803
rect -1461 35784 -1427 35803
rect -1389 35784 -1355 35803
rect -1317 35784 -1283 35803
rect -1245 35784 -1211 35803
rect -1173 35784 -1139 35803
rect -1101 35784 -1067 35803
rect -1029 35784 -995 35803
rect -957 35784 -923 35803
rect -885 35784 -851 35803
rect -813 35784 -779 35803
rect -741 35784 -707 35803
rect -669 35784 -635 35803
rect -597 35784 -563 35803
rect -525 35784 -491 35803
rect -453 35784 -419 35803
rect -381 35784 -347 35803
rect -309 35784 -275 35803
rect -2829 35734 -2802 35745
rect -2802 35734 -2795 35745
rect -2757 35734 -2734 35745
rect -2734 35734 -2723 35745
rect -2685 35734 -2666 35745
rect -2666 35734 -2651 35745
rect -2613 35734 -2598 35745
rect -2598 35734 -2579 35745
rect -2541 35734 -2530 35745
rect -2530 35734 -2507 35745
rect -2469 35734 -2462 35745
rect -2462 35734 -2435 35745
rect -2397 35734 -2394 35745
rect -2394 35734 -2363 35745
rect -2325 35734 -2292 35745
rect -2292 35734 -2291 35745
rect -2253 35734 -2224 35745
rect -2224 35734 -2219 35745
rect -2181 35734 -2156 35745
rect -2156 35734 -2147 35745
rect -2109 35734 -2088 35745
rect -2088 35734 -2075 35745
rect -2037 35734 -2020 35745
rect -2020 35734 -2003 35745
rect -1965 35734 -1952 35745
rect -1952 35734 -1931 35745
rect -1893 35734 -1884 35745
rect -1884 35734 -1859 35745
rect -1821 35734 -1816 35745
rect -1816 35734 -1787 35745
rect -1749 35734 -1748 35745
rect -1748 35734 -1715 35745
rect -1677 35734 -1646 35745
rect -1646 35734 -1643 35745
rect -1605 35734 -1578 35745
rect -1578 35734 -1571 35745
rect -1533 35734 -1510 35745
rect -1510 35734 -1499 35745
rect -1461 35734 -1442 35745
rect -1442 35734 -1427 35745
rect -1389 35734 -1374 35745
rect -1374 35734 -1355 35745
rect -1317 35734 -1306 35745
rect -1306 35734 -1283 35745
rect -1245 35734 -1238 35745
rect -1238 35734 -1211 35745
rect -1173 35734 -1170 35745
rect -1170 35734 -1139 35745
rect -1101 35734 -1068 35745
rect -1068 35734 -1067 35745
rect -1029 35734 -1000 35745
rect -1000 35734 -995 35745
rect -957 35734 -932 35745
rect -932 35734 -923 35745
rect -885 35734 -864 35745
rect -864 35734 -851 35745
rect -813 35734 -796 35745
rect -796 35734 -779 35745
rect -741 35734 -728 35745
rect -728 35734 -707 35745
rect -669 35734 -660 35745
rect -660 35734 -635 35745
rect -597 35734 -592 35745
rect -592 35734 -563 35745
rect -525 35734 -524 35745
rect -524 35734 -491 35745
rect -453 35734 -422 35745
rect -422 35734 -419 35745
rect -381 35734 -354 35745
rect -354 35734 -347 35745
rect -309 35734 -286 35745
rect -286 35734 -275 35745
rect -2829 35711 -2795 35734
rect -2757 35711 -2723 35734
rect -2685 35711 -2651 35734
rect -2613 35711 -2579 35734
rect -2541 35711 -2507 35734
rect -2469 35711 -2435 35734
rect -2397 35711 -2363 35734
rect -2325 35711 -2291 35734
rect -2253 35711 -2219 35734
rect -2181 35711 -2147 35734
rect -2109 35711 -2075 35734
rect -2037 35711 -2003 35734
rect -1965 35711 -1931 35734
rect -1893 35711 -1859 35734
rect -1821 35711 -1787 35734
rect -1749 35711 -1715 35734
rect -1677 35711 -1643 35734
rect -1605 35711 -1571 35734
rect -1533 35711 -1499 35734
rect -1461 35711 -1427 35734
rect -1389 35711 -1355 35734
rect -1317 35711 -1283 35734
rect -1245 35711 -1211 35734
rect -1173 35711 -1139 35734
rect -1101 35711 -1067 35734
rect -1029 35711 -995 35734
rect -957 35711 -923 35734
rect -885 35711 -851 35734
rect -813 35711 -779 35734
rect -741 35711 -707 35734
rect -669 35711 -635 35734
rect -597 35711 -563 35734
rect -525 35711 -491 35734
rect -453 35711 -419 35734
rect -381 35711 -347 35734
rect -309 35711 -275 35734
rect -2829 35665 -2802 35672
rect -2802 35665 -2795 35672
rect -2757 35665 -2734 35672
rect -2734 35665 -2723 35672
rect -2685 35665 -2666 35672
rect -2666 35665 -2651 35672
rect -2613 35665 -2598 35672
rect -2598 35665 -2579 35672
rect -2541 35665 -2530 35672
rect -2530 35665 -2507 35672
rect -2469 35665 -2462 35672
rect -2462 35665 -2435 35672
rect -2397 35665 -2394 35672
rect -2394 35665 -2363 35672
rect -2325 35665 -2292 35672
rect -2292 35665 -2291 35672
rect -2253 35665 -2224 35672
rect -2224 35665 -2219 35672
rect -2181 35665 -2156 35672
rect -2156 35665 -2147 35672
rect -2109 35665 -2088 35672
rect -2088 35665 -2075 35672
rect -2037 35665 -2020 35672
rect -2020 35665 -2003 35672
rect -1965 35665 -1952 35672
rect -1952 35665 -1931 35672
rect -1893 35665 -1884 35672
rect -1884 35665 -1859 35672
rect -1821 35665 -1816 35672
rect -1816 35665 -1787 35672
rect -1749 35665 -1748 35672
rect -1748 35665 -1715 35672
rect -1677 35665 -1646 35672
rect -1646 35665 -1643 35672
rect -1605 35665 -1578 35672
rect -1578 35665 -1571 35672
rect -1533 35665 -1510 35672
rect -1510 35665 -1499 35672
rect -1461 35665 -1442 35672
rect -1442 35665 -1427 35672
rect -1389 35665 -1374 35672
rect -1374 35665 -1355 35672
rect -1317 35665 -1306 35672
rect -1306 35665 -1283 35672
rect -1245 35665 -1238 35672
rect -1238 35665 -1211 35672
rect -1173 35665 -1170 35672
rect -1170 35665 -1139 35672
rect -1101 35665 -1068 35672
rect -1068 35665 -1067 35672
rect -1029 35665 -1000 35672
rect -1000 35665 -995 35672
rect -957 35665 -932 35672
rect -932 35665 -923 35672
rect -885 35665 -864 35672
rect -864 35665 -851 35672
rect -813 35665 -796 35672
rect -796 35665 -779 35672
rect -741 35665 -728 35672
rect -728 35665 -707 35672
rect -669 35665 -660 35672
rect -660 35665 -635 35672
rect -597 35665 -592 35672
rect -592 35665 -563 35672
rect -525 35665 -524 35672
rect -524 35665 -491 35672
rect -453 35665 -422 35672
rect -422 35665 -419 35672
rect -381 35665 -354 35672
rect -354 35665 -347 35672
rect -309 35665 -286 35672
rect -286 35665 -275 35672
rect -2829 35638 -2795 35665
rect -2757 35638 -2723 35665
rect -2685 35638 -2651 35665
rect -2613 35638 -2579 35665
rect -2541 35638 -2507 35665
rect -2469 35638 -2435 35665
rect -2397 35638 -2363 35665
rect -2325 35638 -2291 35665
rect -2253 35638 -2219 35665
rect -2181 35638 -2147 35665
rect -2109 35638 -2075 35665
rect -2037 35638 -2003 35665
rect -1965 35638 -1931 35665
rect -1893 35638 -1859 35665
rect -1821 35638 -1787 35665
rect -1749 35638 -1715 35665
rect -1677 35638 -1643 35665
rect -1605 35638 -1571 35665
rect -1533 35638 -1499 35665
rect -1461 35638 -1427 35665
rect -1389 35638 -1355 35665
rect -1317 35638 -1283 35665
rect -1245 35638 -1211 35665
rect -1173 35638 -1139 35665
rect -1101 35638 -1067 35665
rect -1029 35638 -995 35665
rect -957 35638 -923 35665
rect -885 35638 -851 35665
rect -813 35638 -779 35665
rect -741 35638 -707 35665
rect -669 35638 -635 35665
rect -597 35638 -563 35665
rect -525 35638 -491 35665
rect -453 35638 -419 35665
rect -381 35638 -347 35665
rect -309 35638 -275 35665
rect -2829 35596 -2802 35599
rect -2802 35596 -2795 35599
rect -2757 35596 -2734 35599
rect -2734 35596 -2723 35599
rect -2685 35596 -2666 35599
rect -2666 35596 -2651 35599
rect -2613 35596 -2598 35599
rect -2598 35596 -2579 35599
rect -2541 35596 -2530 35599
rect -2530 35596 -2507 35599
rect -2469 35596 -2462 35599
rect -2462 35596 -2435 35599
rect -2397 35596 -2394 35599
rect -2394 35596 -2363 35599
rect -2325 35596 -2292 35599
rect -2292 35596 -2291 35599
rect -2253 35596 -2224 35599
rect -2224 35596 -2219 35599
rect -2181 35596 -2156 35599
rect -2156 35596 -2147 35599
rect -2109 35596 -2088 35599
rect -2088 35596 -2075 35599
rect -2037 35596 -2020 35599
rect -2020 35596 -2003 35599
rect -1965 35596 -1952 35599
rect -1952 35596 -1931 35599
rect -1893 35596 -1884 35599
rect -1884 35596 -1859 35599
rect -1821 35596 -1816 35599
rect -1816 35596 -1787 35599
rect -1749 35596 -1748 35599
rect -1748 35596 -1715 35599
rect -1677 35596 -1646 35599
rect -1646 35596 -1643 35599
rect -1605 35596 -1578 35599
rect -1578 35596 -1571 35599
rect -1533 35596 -1510 35599
rect -1510 35596 -1499 35599
rect -1461 35596 -1442 35599
rect -1442 35596 -1427 35599
rect -1389 35596 -1374 35599
rect -1374 35596 -1355 35599
rect -1317 35596 -1306 35599
rect -1306 35596 -1283 35599
rect -1245 35596 -1238 35599
rect -1238 35596 -1211 35599
rect -1173 35596 -1170 35599
rect -1170 35596 -1139 35599
rect -1101 35596 -1068 35599
rect -1068 35596 -1067 35599
rect -1029 35596 -1000 35599
rect -1000 35596 -995 35599
rect -957 35596 -932 35599
rect -932 35596 -923 35599
rect -885 35596 -864 35599
rect -864 35596 -851 35599
rect -813 35596 -796 35599
rect -796 35596 -779 35599
rect -741 35596 -728 35599
rect -728 35596 -707 35599
rect -669 35596 -660 35599
rect -660 35596 -635 35599
rect -597 35596 -592 35599
rect -592 35596 -563 35599
rect -525 35596 -524 35599
rect -524 35596 -491 35599
rect -453 35596 -422 35599
rect -422 35596 -419 35599
rect -381 35596 -354 35599
rect -354 35596 -347 35599
rect -309 35596 -286 35599
rect -286 35596 -275 35599
rect -2829 35565 -2795 35596
rect -2757 35565 -2723 35596
rect -2685 35565 -2651 35596
rect -2613 35565 -2579 35596
rect -2541 35565 -2507 35596
rect -2469 35565 -2435 35596
rect -2397 35565 -2363 35596
rect -2325 35565 -2291 35596
rect -2253 35565 -2219 35596
rect -2181 35565 -2147 35596
rect -2109 35565 -2075 35596
rect -2037 35565 -2003 35596
rect -1965 35565 -1931 35596
rect -1893 35565 -1859 35596
rect -1821 35565 -1787 35596
rect -1749 35565 -1715 35596
rect -1677 35565 -1643 35596
rect -1605 35565 -1571 35596
rect -1533 35565 -1499 35596
rect -1461 35565 -1427 35596
rect -1389 35565 -1355 35596
rect -1317 35565 -1283 35596
rect -1245 35565 -1211 35596
rect -1173 35565 -1139 35596
rect -1101 35565 -1067 35596
rect -1029 35565 -995 35596
rect -957 35565 -923 35596
rect -885 35565 -851 35596
rect -813 35565 -779 35596
rect -741 35565 -707 35596
rect -669 35565 -635 35596
rect -597 35565 -563 35596
rect -525 35565 -491 35596
rect -453 35565 -419 35596
rect -381 35565 -347 35596
rect -309 35565 -275 35596
rect -2829 35492 -2795 35526
rect -2757 35492 -2723 35526
rect -2685 35492 -2651 35526
rect -2613 35492 -2579 35526
rect -2541 35492 -2507 35526
rect -2469 35492 -2435 35526
rect -2397 35492 -2363 35526
rect -2325 35492 -2291 35526
rect -2253 35492 -2219 35526
rect -2181 35492 -2147 35526
rect -2109 35492 -2075 35526
rect -2037 35492 -2003 35526
rect -1965 35492 -1931 35526
rect -1893 35492 -1859 35526
rect -1821 35492 -1787 35526
rect -1749 35492 -1715 35526
rect -1677 35492 -1643 35526
rect -1605 35492 -1571 35526
rect -1533 35492 -1499 35526
rect -1461 35492 -1427 35526
rect -1389 35492 -1355 35526
rect -1317 35492 -1283 35526
rect -1245 35492 -1211 35526
rect -1173 35492 -1139 35526
rect -1101 35492 -1067 35526
rect -1029 35492 -995 35526
rect -957 35492 -923 35526
rect -885 35492 -851 35526
rect -813 35492 -779 35526
rect -741 35492 -707 35526
rect -669 35492 -635 35526
rect -597 35492 -563 35526
rect -525 35492 -491 35526
rect -453 35492 -419 35526
rect -381 35492 -347 35526
rect -309 35492 -275 35526
rect -2829 35423 -2795 35453
rect -2757 35423 -2723 35453
rect -2685 35423 -2651 35453
rect -2613 35423 -2579 35453
rect -2541 35423 -2507 35453
rect -2469 35423 -2435 35453
rect -2397 35423 -2363 35453
rect -2325 35423 -2291 35453
rect -2253 35423 -2219 35453
rect -2181 35423 -2147 35453
rect -2109 35423 -2075 35453
rect -2037 35423 -2003 35453
rect -1965 35423 -1931 35453
rect -1893 35423 -1859 35453
rect -1821 35423 -1787 35453
rect -1749 35423 -1715 35453
rect -1677 35423 -1643 35453
rect -1605 35423 -1571 35453
rect -1533 35423 -1499 35453
rect -1461 35423 -1427 35453
rect -1389 35423 -1355 35453
rect -1317 35423 -1283 35453
rect -1245 35423 -1211 35453
rect -1173 35423 -1139 35453
rect -1101 35423 -1067 35453
rect -1029 35423 -995 35453
rect -957 35423 -923 35453
rect -885 35423 -851 35453
rect -813 35423 -779 35453
rect -741 35423 -707 35453
rect -669 35423 -635 35453
rect -597 35423 -563 35453
rect -525 35423 -491 35453
rect -453 35423 -419 35453
rect -381 35423 -347 35453
rect -309 35423 -275 35453
rect -2829 35419 -2802 35423
rect -2802 35419 -2795 35423
rect -2757 35419 -2734 35423
rect -2734 35419 -2723 35423
rect -2685 35419 -2666 35423
rect -2666 35419 -2651 35423
rect -2613 35419 -2598 35423
rect -2598 35419 -2579 35423
rect -2541 35419 -2530 35423
rect -2530 35419 -2507 35423
rect -2469 35419 -2462 35423
rect -2462 35419 -2435 35423
rect -2397 35419 -2394 35423
rect -2394 35419 -2363 35423
rect -2325 35419 -2292 35423
rect -2292 35419 -2291 35423
rect -2253 35419 -2224 35423
rect -2224 35419 -2219 35423
rect -2181 35419 -2156 35423
rect -2156 35419 -2147 35423
rect -2109 35419 -2088 35423
rect -2088 35419 -2075 35423
rect -2037 35419 -2020 35423
rect -2020 35419 -2003 35423
rect -1965 35419 -1952 35423
rect -1952 35419 -1931 35423
rect -1893 35419 -1884 35423
rect -1884 35419 -1859 35423
rect -1821 35419 -1816 35423
rect -1816 35419 -1787 35423
rect -1749 35419 -1748 35423
rect -1748 35419 -1715 35423
rect -1677 35419 -1646 35423
rect -1646 35419 -1643 35423
rect -1605 35419 -1578 35423
rect -1578 35419 -1571 35423
rect -1533 35419 -1510 35423
rect -1510 35419 -1499 35423
rect -1461 35419 -1442 35423
rect -1442 35419 -1427 35423
rect -1389 35419 -1374 35423
rect -1374 35419 -1355 35423
rect -1317 35419 -1306 35423
rect -1306 35419 -1283 35423
rect -1245 35419 -1238 35423
rect -1238 35419 -1211 35423
rect -1173 35419 -1170 35423
rect -1170 35419 -1139 35423
rect -1101 35419 -1068 35423
rect -1068 35419 -1067 35423
rect -1029 35419 -1000 35423
rect -1000 35419 -995 35423
rect -957 35419 -932 35423
rect -932 35419 -923 35423
rect -885 35419 -864 35423
rect -864 35419 -851 35423
rect -813 35419 -796 35423
rect -796 35419 -779 35423
rect -741 35419 -728 35423
rect -728 35419 -707 35423
rect -669 35419 -660 35423
rect -660 35419 -635 35423
rect -597 35419 -592 35423
rect -592 35419 -563 35423
rect -525 35419 -524 35423
rect -524 35419 -491 35423
rect -453 35419 -422 35423
rect -422 35419 -419 35423
rect -381 35419 -354 35423
rect -354 35419 -347 35423
rect -309 35419 -286 35423
rect -286 35419 -275 35423
rect -2829 35354 -2795 35380
rect -2757 35354 -2723 35380
rect -2685 35354 -2651 35380
rect -2613 35354 -2579 35380
rect -2541 35354 -2507 35380
rect -2469 35354 -2435 35380
rect -2397 35354 -2363 35380
rect -2325 35354 -2291 35380
rect -2253 35354 -2219 35380
rect -2181 35354 -2147 35380
rect -2109 35354 -2075 35380
rect -2037 35354 -2003 35380
rect -1965 35354 -1931 35380
rect -1893 35354 -1859 35380
rect -1821 35354 -1787 35380
rect -1749 35354 -1715 35380
rect -1677 35354 -1643 35380
rect -1605 35354 -1571 35380
rect -1533 35354 -1499 35380
rect -1461 35354 -1427 35380
rect -1389 35354 -1355 35380
rect -1317 35354 -1283 35380
rect -1245 35354 -1211 35380
rect -1173 35354 -1139 35380
rect -1101 35354 -1067 35380
rect -1029 35354 -995 35380
rect -957 35354 -923 35380
rect -885 35354 -851 35380
rect -813 35354 -779 35380
rect -741 35354 -707 35380
rect -669 35354 -635 35380
rect -597 35354 -563 35380
rect -525 35354 -491 35380
rect -453 35354 -419 35380
rect -381 35354 -347 35380
rect -309 35354 -275 35380
rect -2829 35346 -2802 35354
rect -2802 35346 -2795 35354
rect -2757 35346 -2734 35354
rect -2734 35346 -2723 35354
rect -2685 35346 -2666 35354
rect -2666 35346 -2651 35354
rect -2613 35346 -2598 35354
rect -2598 35346 -2579 35354
rect -2541 35346 -2530 35354
rect -2530 35346 -2507 35354
rect -2469 35346 -2462 35354
rect -2462 35346 -2435 35354
rect -2397 35346 -2394 35354
rect -2394 35346 -2363 35354
rect -2325 35346 -2292 35354
rect -2292 35346 -2291 35354
rect -2253 35346 -2224 35354
rect -2224 35346 -2219 35354
rect -2181 35346 -2156 35354
rect -2156 35346 -2147 35354
rect -2109 35346 -2088 35354
rect -2088 35346 -2075 35354
rect -2037 35346 -2020 35354
rect -2020 35346 -2003 35354
rect -1965 35346 -1952 35354
rect -1952 35346 -1931 35354
rect -1893 35346 -1884 35354
rect -1884 35346 -1859 35354
rect -1821 35346 -1816 35354
rect -1816 35346 -1787 35354
rect -1749 35346 -1748 35354
rect -1748 35346 -1715 35354
rect -1677 35346 -1646 35354
rect -1646 35346 -1643 35354
rect -1605 35346 -1578 35354
rect -1578 35346 -1571 35354
rect -1533 35346 -1510 35354
rect -1510 35346 -1499 35354
rect -1461 35346 -1442 35354
rect -1442 35346 -1427 35354
rect -1389 35346 -1374 35354
rect -1374 35346 -1355 35354
rect -1317 35346 -1306 35354
rect -1306 35346 -1283 35354
rect -1245 35346 -1238 35354
rect -1238 35346 -1211 35354
rect -1173 35346 -1170 35354
rect -1170 35346 -1139 35354
rect -1101 35346 -1068 35354
rect -1068 35346 -1067 35354
rect -1029 35346 -1000 35354
rect -1000 35346 -995 35354
rect -957 35346 -932 35354
rect -932 35346 -923 35354
rect -885 35346 -864 35354
rect -864 35346 -851 35354
rect -813 35346 -796 35354
rect -796 35346 -779 35354
rect -741 35346 -728 35354
rect -728 35346 -707 35354
rect -669 35346 -660 35354
rect -660 35346 -635 35354
rect -597 35346 -592 35354
rect -592 35346 -563 35354
rect -525 35346 -524 35354
rect -524 35346 -491 35354
rect -453 35346 -422 35354
rect -422 35346 -419 35354
rect -381 35346 -354 35354
rect -354 35346 -347 35354
rect -309 35346 -286 35354
rect -286 35346 -275 35354
rect -2829 35285 -2795 35307
rect -2757 35285 -2723 35307
rect -2685 35285 -2651 35307
rect -2613 35285 -2579 35307
rect -2541 35285 -2507 35307
rect -2469 35285 -2435 35307
rect -2397 35285 -2363 35307
rect -2325 35285 -2291 35307
rect -2253 35285 -2219 35307
rect -2181 35285 -2147 35307
rect -2109 35285 -2075 35307
rect -2037 35285 -2003 35307
rect -1965 35285 -1931 35307
rect -1893 35285 -1859 35307
rect -1821 35285 -1787 35307
rect -1749 35285 -1715 35307
rect -1677 35285 -1643 35307
rect -1605 35285 -1571 35307
rect -1533 35285 -1499 35307
rect -1461 35285 -1427 35307
rect -1389 35285 -1355 35307
rect -1317 35285 -1283 35307
rect -1245 35285 -1211 35307
rect -1173 35285 -1139 35307
rect -1101 35285 -1067 35307
rect -1029 35285 -995 35307
rect -957 35285 -923 35307
rect -885 35285 -851 35307
rect -813 35285 -779 35307
rect -741 35285 -707 35307
rect -669 35285 -635 35307
rect -597 35285 -563 35307
rect -525 35285 -491 35307
rect -453 35285 -419 35307
rect -381 35285 -347 35307
rect -309 35285 -275 35307
rect -2829 35273 -2802 35285
rect -2802 35273 -2795 35285
rect -2757 35273 -2734 35285
rect -2734 35273 -2723 35285
rect -2685 35273 -2666 35285
rect -2666 35273 -2651 35285
rect -2613 35273 -2598 35285
rect -2598 35273 -2579 35285
rect -2541 35273 -2530 35285
rect -2530 35273 -2507 35285
rect -2469 35273 -2462 35285
rect -2462 35273 -2435 35285
rect -2397 35273 -2394 35285
rect -2394 35273 -2363 35285
rect -2325 35273 -2292 35285
rect -2292 35273 -2291 35285
rect -2253 35273 -2224 35285
rect -2224 35273 -2219 35285
rect -2181 35273 -2156 35285
rect -2156 35273 -2147 35285
rect -2109 35273 -2088 35285
rect -2088 35273 -2075 35285
rect -2037 35273 -2020 35285
rect -2020 35273 -2003 35285
rect -1965 35273 -1952 35285
rect -1952 35273 -1931 35285
rect -1893 35273 -1884 35285
rect -1884 35273 -1859 35285
rect -1821 35273 -1816 35285
rect -1816 35273 -1787 35285
rect -1749 35273 -1748 35285
rect -1748 35273 -1715 35285
rect -1677 35273 -1646 35285
rect -1646 35273 -1643 35285
rect -1605 35273 -1578 35285
rect -1578 35273 -1571 35285
rect -1533 35273 -1510 35285
rect -1510 35273 -1499 35285
rect -1461 35273 -1442 35285
rect -1442 35273 -1427 35285
rect -1389 35273 -1374 35285
rect -1374 35273 -1355 35285
rect -1317 35273 -1306 35285
rect -1306 35273 -1283 35285
rect -1245 35273 -1238 35285
rect -1238 35273 -1211 35285
rect -1173 35273 -1170 35285
rect -1170 35273 -1139 35285
rect -1101 35273 -1068 35285
rect -1068 35273 -1067 35285
rect -1029 35273 -1000 35285
rect -1000 35273 -995 35285
rect -957 35273 -932 35285
rect -932 35273 -923 35285
rect -885 35273 -864 35285
rect -864 35273 -851 35285
rect -813 35273 -796 35285
rect -796 35273 -779 35285
rect -741 35273 -728 35285
rect -728 35273 -707 35285
rect -669 35273 -660 35285
rect -660 35273 -635 35285
rect -597 35273 -592 35285
rect -592 35273 -563 35285
rect -525 35273 -524 35285
rect -524 35273 -491 35285
rect -453 35273 -422 35285
rect -422 35273 -419 35285
rect -381 35273 -354 35285
rect -354 35273 -347 35285
rect -309 35273 -286 35285
rect -286 35273 -275 35285
rect -2829 35216 -2795 35234
rect -2757 35216 -2723 35234
rect -2685 35216 -2651 35234
rect -2613 35216 -2579 35234
rect -2541 35216 -2507 35234
rect -2469 35216 -2435 35234
rect -2397 35216 -2363 35234
rect -2325 35216 -2291 35234
rect -2253 35216 -2219 35234
rect -2181 35216 -2147 35234
rect -2109 35216 -2075 35234
rect -2037 35216 -2003 35234
rect -1965 35216 -1931 35234
rect -1893 35216 -1859 35234
rect -1821 35216 -1787 35234
rect -1749 35216 -1715 35234
rect -1677 35216 -1643 35234
rect -1605 35216 -1571 35234
rect -1533 35216 -1499 35234
rect -1461 35216 -1427 35234
rect -1389 35216 -1355 35234
rect -1317 35216 -1283 35234
rect -1245 35216 -1211 35234
rect -1173 35216 -1139 35234
rect -1101 35216 -1067 35234
rect -1029 35216 -995 35234
rect -957 35216 -923 35234
rect -885 35216 -851 35234
rect -813 35216 -779 35234
rect -741 35216 -707 35234
rect -669 35216 -635 35234
rect -597 35216 -563 35234
rect -525 35216 -491 35234
rect -453 35216 -419 35234
rect -381 35216 -347 35234
rect -309 35216 -275 35234
rect -2829 35200 -2802 35216
rect -2802 35200 -2795 35216
rect -2757 35200 -2734 35216
rect -2734 35200 -2723 35216
rect -2685 35200 -2666 35216
rect -2666 35200 -2651 35216
rect -2613 35200 -2598 35216
rect -2598 35200 -2579 35216
rect -2541 35200 -2530 35216
rect -2530 35200 -2507 35216
rect -2469 35200 -2462 35216
rect -2462 35200 -2435 35216
rect -2397 35200 -2394 35216
rect -2394 35200 -2363 35216
rect -2325 35200 -2292 35216
rect -2292 35200 -2291 35216
rect -2253 35200 -2224 35216
rect -2224 35200 -2219 35216
rect -2181 35200 -2156 35216
rect -2156 35200 -2147 35216
rect -2109 35200 -2088 35216
rect -2088 35200 -2075 35216
rect -2037 35200 -2020 35216
rect -2020 35200 -2003 35216
rect -1965 35200 -1952 35216
rect -1952 35200 -1931 35216
rect -1893 35200 -1884 35216
rect -1884 35200 -1859 35216
rect -1821 35200 -1816 35216
rect -1816 35200 -1787 35216
rect -1749 35200 -1748 35216
rect -1748 35200 -1715 35216
rect -1677 35200 -1646 35216
rect -1646 35200 -1643 35216
rect -1605 35200 -1578 35216
rect -1578 35200 -1571 35216
rect -1533 35200 -1510 35216
rect -1510 35200 -1499 35216
rect -1461 35200 -1442 35216
rect -1442 35200 -1427 35216
rect -1389 35200 -1374 35216
rect -1374 35200 -1355 35216
rect -1317 35200 -1306 35216
rect -1306 35200 -1283 35216
rect -1245 35200 -1238 35216
rect -1238 35200 -1211 35216
rect -1173 35200 -1170 35216
rect -1170 35200 -1139 35216
rect -1101 35200 -1068 35216
rect -1068 35200 -1067 35216
rect -1029 35200 -1000 35216
rect -1000 35200 -995 35216
rect -957 35200 -932 35216
rect -932 35200 -923 35216
rect -885 35200 -864 35216
rect -864 35200 -851 35216
rect -813 35200 -796 35216
rect -796 35200 -779 35216
rect -741 35200 -728 35216
rect -728 35200 -707 35216
rect -669 35200 -660 35216
rect -660 35200 -635 35216
rect -597 35200 -592 35216
rect -592 35200 -563 35216
rect -525 35200 -524 35216
rect -524 35200 -491 35216
rect -453 35200 -422 35216
rect -422 35200 -419 35216
rect -381 35200 -354 35216
rect -354 35200 -347 35216
rect -309 35200 -286 35216
rect -286 35200 -275 35216
rect -2829 35147 -2795 35161
rect -2757 35147 -2723 35161
rect -2685 35147 -2651 35161
rect -2613 35147 -2579 35161
rect -2541 35147 -2507 35161
rect -2469 35147 -2435 35161
rect -2397 35147 -2363 35161
rect -2325 35147 -2291 35161
rect -2253 35147 -2219 35161
rect -2181 35147 -2147 35161
rect -2109 35147 -2075 35161
rect -2037 35147 -2003 35161
rect -1965 35147 -1931 35161
rect -1893 35147 -1859 35161
rect -1821 35147 -1787 35161
rect -1749 35147 -1715 35161
rect -1677 35147 -1643 35161
rect -1605 35147 -1571 35161
rect -1533 35147 -1499 35161
rect -1461 35147 -1427 35161
rect -1389 35147 -1355 35161
rect -1317 35147 -1283 35161
rect -1245 35147 -1211 35161
rect -1173 35147 -1139 35161
rect -1101 35147 -1067 35161
rect -1029 35147 -995 35161
rect -957 35147 -923 35161
rect -885 35147 -851 35161
rect -813 35147 -779 35161
rect -741 35147 -707 35161
rect -669 35147 -635 35161
rect -597 35147 -563 35161
rect -525 35147 -491 35161
rect -453 35147 -419 35161
rect -381 35147 -347 35161
rect -309 35147 -275 35161
rect -2829 35127 -2802 35147
rect -2802 35127 -2795 35147
rect -2757 35127 -2734 35147
rect -2734 35127 -2723 35147
rect -2685 35127 -2666 35147
rect -2666 35127 -2651 35147
rect -2613 35127 -2598 35147
rect -2598 35127 -2579 35147
rect -2541 35127 -2530 35147
rect -2530 35127 -2507 35147
rect -2469 35127 -2462 35147
rect -2462 35127 -2435 35147
rect -2397 35127 -2394 35147
rect -2394 35127 -2363 35147
rect -2325 35127 -2292 35147
rect -2292 35127 -2291 35147
rect -2253 35127 -2224 35147
rect -2224 35127 -2219 35147
rect -2181 35127 -2156 35147
rect -2156 35127 -2147 35147
rect -2109 35127 -2088 35147
rect -2088 35127 -2075 35147
rect -2037 35127 -2020 35147
rect -2020 35127 -2003 35147
rect -1965 35127 -1952 35147
rect -1952 35127 -1931 35147
rect -1893 35127 -1884 35147
rect -1884 35127 -1859 35147
rect -1821 35127 -1816 35147
rect -1816 35127 -1787 35147
rect -1749 35127 -1748 35147
rect -1748 35127 -1715 35147
rect -1677 35127 -1646 35147
rect -1646 35127 -1643 35147
rect -1605 35127 -1578 35147
rect -1578 35127 -1571 35147
rect -1533 35127 -1510 35147
rect -1510 35127 -1499 35147
rect -1461 35127 -1442 35147
rect -1442 35127 -1427 35147
rect -1389 35127 -1374 35147
rect -1374 35127 -1355 35147
rect -1317 35127 -1306 35147
rect -1306 35127 -1283 35147
rect -1245 35127 -1238 35147
rect -1238 35127 -1211 35147
rect -1173 35127 -1170 35147
rect -1170 35127 -1139 35147
rect -1101 35127 -1068 35147
rect -1068 35127 -1067 35147
rect -1029 35127 -1000 35147
rect -1000 35127 -995 35147
rect -957 35127 -932 35147
rect -932 35127 -923 35147
rect -885 35127 -864 35147
rect -864 35127 -851 35147
rect -813 35127 -796 35147
rect -796 35127 -779 35147
rect -741 35127 -728 35147
rect -728 35127 -707 35147
rect -669 35127 -660 35147
rect -660 35127 -635 35147
rect -597 35127 -592 35147
rect -592 35127 -563 35147
rect -525 35127 -524 35147
rect -524 35127 -491 35147
rect -453 35127 -422 35147
rect -422 35127 -419 35147
rect -381 35127 -354 35147
rect -354 35127 -347 35147
rect -309 35127 -286 35147
rect -286 35127 -275 35147
rect 10732 15836 10766 15870
rect 10732 15739 10766 15773
rect 10989 15836 11023 15870
rect 10989 15717 11023 15751
rect 11341 15836 11375 15870
rect 11341 15717 11375 15751
rect 11637 15836 11671 15870
rect 11637 15717 11671 15751
rect 10732 15121 10766 15155
rect 10732 15024 10766 15058
rect 10989 15143 11023 15177
rect 10989 15024 11023 15058
rect 11341 15143 11375 15177
rect 11341 15024 11375 15058
rect 11637 15143 11671 15177
rect 11723 15143 11757 15177
rect 11637 15024 11671 15058
rect 11723 15024 11757 15058
rect 51 14199 85 14233
rect 124 14199 158 14233
rect 197 14199 231 14233
rect 270 14199 304 14233
rect 343 14199 377 14233
rect 416 14199 450 14233
rect 489 14199 523 14233
rect 563 14199 597 14233
rect 637 14199 671 14233
rect 711 14199 745 14233
rect 783 14211 817 14245
rect 51 14127 85 14161
rect 124 14127 158 14161
rect 197 14127 231 14161
rect 270 14127 304 14161
rect 343 14127 377 14161
rect 416 14127 450 14161
rect 489 14127 523 14161
rect 563 14127 597 14161
rect 637 14127 671 14161
rect 711 14127 745 14161
rect 783 14134 817 14168
rect 1031 14211 1065 14245
rect 1031 14137 1065 14171
rect 5588 14211 5622 14245
rect 5701 14211 5735 14245
rect 51 14055 85 14089
rect 124 14055 158 14089
rect 197 14055 231 14089
rect 270 14055 304 14089
rect 343 14055 377 14089
rect 416 14055 450 14089
rect 489 14055 523 14089
rect 563 14055 597 14089
rect 637 14055 671 14089
rect 711 14055 745 14089
rect 783 14057 817 14091
rect 6259 14171 6293 14205
rect 6571 14171 6605 14205
rect 6883 14171 6917 14205
rect 18359 14375 18390 14398
rect 18390 14375 18393 14398
rect 18432 14375 18459 14398
rect 18459 14375 18466 14398
rect 18505 14375 18528 14398
rect 18528 14375 18539 14398
rect 18578 14375 18597 14398
rect 18597 14375 18612 14398
rect 18651 14375 18666 14398
rect 18666 14375 18685 14398
rect 18724 14375 18735 14398
rect 18735 14375 18758 14398
rect 18797 14375 18804 14398
rect 18804 14375 18831 14398
rect 18870 14375 18873 14398
rect 18873 14375 18904 14398
rect 18359 14364 18393 14375
rect 18432 14364 18466 14375
rect 18505 14364 18539 14375
rect 18578 14364 18612 14375
rect 18651 14364 18685 14375
rect 18724 14364 18758 14375
rect 18797 14364 18831 14375
rect 18870 14364 18904 14375
rect 18943 14364 18977 14398
rect 19016 14375 19046 14398
rect 19046 14375 19050 14398
rect 19089 14375 19115 14398
rect 19115 14375 19123 14398
rect 19162 14375 19184 14398
rect 19184 14375 19196 14398
rect 19235 14375 19253 14398
rect 19253 14375 19269 14398
rect 19308 14375 19322 14398
rect 19322 14375 19342 14398
rect 19381 14375 19391 14398
rect 19391 14375 19415 14398
rect 19454 14375 19460 14398
rect 19460 14375 19488 14398
rect 19527 14375 19529 14398
rect 19529 14375 19561 14398
rect 19600 14375 19632 14398
rect 19632 14375 19634 14398
rect 19673 14375 19701 14398
rect 19701 14375 19707 14398
rect 19746 14375 19770 14398
rect 19770 14375 19780 14398
rect 19819 14375 19839 14398
rect 19839 14375 19853 14398
rect 19892 14375 19908 14398
rect 19908 14375 19926 14398
rect 19965 14375 19977 14398
rect 19977 14375 19999 14398
rect 20038 14375 20046 14398
rect 20046 14375 20072 14398
rect 20111 14375 20115 14398
rect 20115 14375 20145 14398
rect 19016 14364 19050 14375
rect 19089 14364 19123 14375
rect 19162 14364 19196 14375
rect 19235 14364 19269 14375
rect 19308 14364 19342 14375
rect 19381 14364 19415 14375
rect 19454 14364 19488 14375
rect 19527 14364 19561 14375
rect 19600 14364 19634 14375
rect 19673 14364 19707 14375
rect 19746 14364 19780 14375
rect 19819 14364 19853 14375
rect 19892 14364 19926 14375
rect 19965 14364 19999 14375
rect 20038 14364 20072 14375
rect 20111 14364 20145 14375
rect 20184 14364 20218 14398
rect 20257 14375 20288 14398
rect 20288 14375 20291 14398
rect 20330 14375 20357 14398
rect 20357 14375 20364 14398
rect 20403 14375 20426 14398
rect 20426 14375 20437 14398
rect 20476 14375 20495 14398
rect 20495 14375 20510 14398
rect 20549 14375 20564 14398
rect 20564 14375 20583 14398
rect 20622 14375 20633 14398
rect 20633 14375 20656 14398
rect 20695 14375 20702 14398
rect 20702 14375 20729 14398
rect 20768 14375 20771 14398
rect 20771 14375 20802 14398
rect 20841 14375 20873 14398
rect 20873 14375 20875 14398
rect 20914 14375 20941 14398
rect 20941 14375 20948 14398
rect 20987 14375 21009 14398
rect 21009 14375 21021 14398
rect 21060 14375 21077 14398
rect 21077 14375 21094 14398
rect 21133 14375 21145 14398
rect 21145 14375 21167 14398
rect 21206 14375 21213 14398
rect 21213 14375 21240 14398
rect 21279 14375 21281 14398
rect 21281 14375 21313 14398
rect 21352 14375 21383 14398
rect 21383 14375 21386 14398
rect 21425 14375 21451 14398
rect 21451 14375 21459 14398
rect 21498 14375 21519 14398
rect 21519 14375 21532 14398
rect 21571 14375 21587 14398
rect 21587 14375 21605 14398
rect 21644 14375 21655 14398
rect 21655 14375 21678 14398
rect 21717 14375 21723 14398
rect 21723 14375 21751 14398
rect 21790 14375 21791 14398
rect 21791 14375 21824 14398
rect 21863 14375 21893 14398
rect 21893 14375 21897 14398
rect 21936 14375 21961 14398
rect 21961 14375 21970 14398
rect 22009 14375 22029 14398
rect 22029 14375 22043 14398
rect 22082 14375 22097 14398
rect 22097 14375 22116 14398
rect 22155 14375 22165 14398
rect 22165 14375 22189 14398
rect 22228 14375 22233 14398
rect 22233 14375 22262 14398
rect 20257 14364 20291 14375
rect 20330 14364 20364 14375
rect 20403 14364 20437 14375
rect 20476 14364 20510 14375
rect 20549 14364 20583 14375
rect 20622 14364 20656 14375
rect 20695 14364 20729 14375
rect 20768 14364 20802 14375
rect 20841 14364 20875 14375
rect 20914 14364 20948 14375
rect 20987 14364 21021 14375
rect 21060 14364 21094 14375
rect 21133 14364 21167 14375
rect 21206 14364 21240 14375
rect 21279 14364 21313 14375
rect 21352 14364 21386 14375
rect 21425 14364 21459 14375
rect 21498 14364 21532 14375
rect 21571 14364 21605 14375
rect 21644 14364 21678 14375
rect 21717 14364 21751 14375
rect 21790 14364 21824 14375
rect 21863 14364 21897 14375
rect 21936 14364 21970 14375
rect 22009 14364 22043 14375
rect 22082 14364 22116 14375
rect 22155 14364 22189 14375
rect 22228 14364 22262 14375
rect 22301 14364 22335 14398
rect 22373 14375 22403 14398
rect 22403 14375 22407 14398
rect 22445 14375 22471 14398
rect 22471 14375 22479 14398
rect 22517 14375 22539 14398
rect 22539 14375 22551 14398
rect 22589 14375 22607 14398
rect 22607 14375 22623 14398
rect 22661 14375 22675 14398
rect 22675 14375 22695 14398
rect 22733 14375 22743 14398
rect 22743 14375 22767 14398
rect 22805 14375 22811 14398
rect 22811 14375 22839 14398
rect 22877 14375 22879 14398
rect 22879 14375 22911 14398
rect 22949 14375 22981 14398
rect 22981 14375 22983 14398
rect 23021 14375 23049 14398
rect 23049 14375 23055 14398
rect 23093 14375 23117 14398
rect 23117 14375 23127 14398
rect 23355 14375 23389 14398
rect 23428 14375 23457 14398
rect 23457 14375 23462 14398
rect 23501 14375 23525 14398
rect 23525 14375 23535 14398
rect 23574 14375 23593 14398
rect 23593 14375 23608 14398
rect 23647 14375 23661 14398
rect 23661 14375 23681 14398
rect 23720 14375 23729 14398
rect 23729 14375 23754 14398
rect 23793 14375 23797 14398
rect 23797 14375 23827 14398
rect 22373 14364 22407 14375
rect 22445 14364 22479 14375
rect 22517 14364 22551 14375
rect 22589 14364 22623 14375
rect 22661 14364 22695 14375
rect 22733 14364 22767 14375
rect 22805 14364 22839 14375
rect 22877 14364 22911 14375
rect 22949 14364 22983 14375
rect 23021 14364 23055 14375
rect 23093 14364 23127 14375
rect 23355 14364 23389 14375
rect 23428 14364 23462 14375
rect 23501 14364 23535 14375
rect 23574 14364 23608 14375
rect 23647 14364 23681 14375
rect 23720 14364 23754 14375
rect 23793 14364 23827 14375
rect 23865 14364 23899 14398
rect 23937 14375 23967 14398
rect 23967 14375 23971 14398
rect 24009 14375 24035 14398
rect 24035 14375 24043 14398
rect 24081 14375 24103 14398
rect 24103 14375 24115 14398
rect 24153 14375 24171 14398
rect 24171 14375 24187 14398
rect 24225 14375 24239 14398
rect 24239 14375 24259 14398
rect 24297 14375 24307 14398
rect 24307 14375 24331 14398
rect 24369 14375 24375 14398
rect 24375 14375 24403 14398
rect 24441 14375 24443 14398
rect 24443 14375 24475 14398
rect 24513 14375 24545 14398
rect 24545 14375 24547 14398
rect 24585 14375 24613 14398
rect 24613 14375 24619 14398
rect 24657 14375 24681 14398
rect 24681 14375 24691 14398
rect 24729 14375 24749 14398
rect 24749 14375 24763 14398
rect 24801 14375 24817 14398
rect 24817 14375 24835 14398
rect 24873 14375 24885 14398
rect 24885 14375 24907 14398
rect 24945 14375 24953 14398
rect 24953 14375 24979 14398
rect 25017 14375 25021 14398
rect 25021 14375 25051 14398
rect 23937 14364 23971 14375
rect 24009 14364 24043 14375
rect 24081 14364 24115 14375
rect 24153 14364 24187 14375
rect 24225 14364 24259 14375
rect 24297 14364 24331 14375
rect 24369 14364 24403 14375
rect 24441 14364 24475 14375
rect 24513 14364 24547 14375
rect 24585 14364 24619 14375
rect 24657 14364 24691 14375
rect 24729 14364 24763 14375
rect 24801 14364 24835 14375
rect 24873 14364 24907 14375
rect 24945 14364 24979 14375
rect 25017 14364 25051 14375
rect 25089 14364 25123 14398
rect 25161 14375 25191 14398
rect 25191 14375 25195 14398
rect 25233 14375 25259 14398
rect 25259 14375 25267 14398
rect 25305 14375 25327 14398
rect 25327 14375 25339 14398
rect 25377 14375 25395 14398
rect 25395 14375 25411 14398
rect 25449 14375 25463 14398
rect 25463 14375 25483 14398
rect 25521 14375 25531 14398
rect 25531 14375 25555 14398
rect 25593 14375 25599 14398
rect 25599 14375 25627 14398
rect 25665 14375 25667 14398
rect 25667 14375 25699 14398
rect 25737 14375 25769 14398
rect 25769 14375 25771 14398
rect 25809 14375 25837 14398
rect 25837 14375 25843 14398
rect 25881 14375 25905 14398
rect 25905 14375 25915 14398
rect 25953 14375 25973 14398
rect 25973 14375 25987 14398
rect 26025 14375 26041 14398
rect 26041 14375 26059 14398
rect 26097 14375 26109 14398
rect 26109 14375 26131 14398
rect 26169 14375 26177 14398
rect 26177 14375 26203 14398
rect 26241 14375 26245 14398
rect 26245 14375 26275 14398
rect 25161 14364 25195 14375
rect 25233 14364 25267 14375
rect 25305 14364 25339 14375
rect 25377 14364 25411 14375
rect 25449 14364 25483 14375
rect 25521 14364 25555 14375
rect 25593 14364 25627 14375
rect 25665 14364 25699 14375
rect 25737 14364 25771 14375
rect 25809 14364 25843 14375
rect 25881 14364 25915 14375
rect 25953 14364 25987 14375
rect 26025 14364 26059 14375
rect 26097 14364 26131 14375
rect 26169 14364 26203 14375
rect 26241 14364 26275 14375
rect 26313 14364 26347 14398
rect 26385 14375 26415 14398
rect 26415 14375 26419 14398
rect 26457 14375 26483 14398
rect 26483 14375 26491 14398
rect 26529 14375 26551 14398
rect 26551 14375 26563 14398
rect 26601 14375 26619 14398
rect 26619 14375 26635 14398
rect 26673 14375 26687 14398
rect 26687 14375 26707 14398
rect 26745 14375 26755 14398
rect 26755 14375 26779 14398
rect 26817 14375 26823 14398
rect 26823 14375 26851 14398
rect 26889 14375 26891 14398
rect 26891 14375 26923 14398
rect 26961 14375 26993 14398
rect 26993 14375 26995 14398
rect 27033 14375 27061 14398
rect 27061 14375 27067 14398
rect 27105 14375 27129 14398
rect 27129 14375 27139 14398
rect 27177 14375 27197 14398
rect 27197 14375 27211 14398
rect 27249 14375 27265 14398
rect 27265 14375 27283 14398
rect 27321 14375 27333 14398
rect 27333 14375 27355 14398
rect 27393 14375 27401 14398
rect 27401 14375 27427 14398
rect 27465 14375 27469 14398
rect 27469 14375 27499 14398
rect 26385 14364 26419 14375
rect 26457 14364 26491 14375
rect 26529 14364 26563 14375
rect 26601 14364 26635 14375
rect 26673 14364 26707 14375
rect 26745 14364 26779 14375
rect 26817 14364 26851 14375
rect 26889 14364 26923 14375
rect 26961 14364 26995 14375
rect 27033 14364 27067 14375
rect 27105 14364 27139 14375
rect 27177 14364 27211 14375
rect 27249 14364 27283 14375
rect 27321 14364 27355 14375
rect 27393 14364 27427 14375
rect 27465 14364 27499 14375
rect 27537 14364 27571 14398
rect 27609 14375 27639 14398
rect 27639 14375 27643 14398
rect 27681 14375 27707 14398
rect 27707 14375 27715 14398
rect 27753 14375 27775 14398
rect 27775 14375 27787 14398
rect 27825 14375 27843 14398
rect 27843 14375 27859 14398
rect 27897 14375 27911 14398
rect 27911 14375 27931 14398
rect 27969 14375 27979 14398
rect 27979 14375 28003 14398
rect 28041 14375 28047 14398
rect 28047 14375 28075 14398
rect 28113 14375 28115 14398
rect 28115 14375 28147 14398
rect 28185 14375 28217 14398
rect 28217 14375 28219 14398
rect 28257 14375 28285 14398
rect 28285 14375 28291 14398
rect 28329 14375 28353 14398
rect 28353 14375 28363 14398
rect 28401 14375 28421 14398
rect 28421 14375 28435 14398
rect 28473 14375 28489 14398
rect 28489 14375 28507 14398
rect 28545 14375 28557 14398
rect 28557 14375 28579 14398
rect 28617 14375 28625 14398
rect 28625 14375 28651 14398
rect 28689 14375 28693 14398
rect 28693 14375 28723 14398
rect 27609 14364 27643 14375
rect 27681 14364 27715 14375
rect 27753 14364 27787 14375
rect 27825 14364 27859 14375
rect 27897 14364 27931 14375
rect 27969 14364 28003 14375
rect 28041 14364 28075 14375
rect 28113 14364 28147 14375
rect 28185 14364 28219 14375
rect 28257 14364 28291 14375
rect 28329 14364 28363 14375
rect 28401 14364 28435 14375
rect 28473 14364 28507 14375
rect 28545 14364 28579 14375
rect 28617 14364 28651 14375
rect 28689 14364 28723 14375
rect 28761 14364 28795 14398
rect 28833 14375 28863 14398
rect 28863 14375 28867 14398
rect 28905 14375 28931 14398
rect 28931 14375 28939 14398
rect 28977 14375 28999 14398
rect 28999 14375 29011 14398
rect 29049 14375 29067 14398
rect 29067 14375 29083 14398
rect 29121 14375 29135 14398
rect 29135 14375 29155 14398
rect 29193 14375 29203 14398
rect 29203 14375 29227 14398
rect 29265 14375 29271 14398
rect 29271 14375 29299 14398
rect 29337 14375 29339 14398
rect 29339 14375 29371 14398
rect 29409 14375 29441 14398
rect 29441 14375 29443 14398
rect 29481 14375 29509 14398
rect 29509 14375 29515 14398
rect 29553 14375 29577 14398
rect 29577 14375 29587 14398
rect 29625 14375 29645 14398
rect 29645 14375 29659 14398
rect 28833 14364 28867 14375
rect 28905 14364 28939 14375
rect 28977 14364 29011 14375
rect 29049 14364 29083 14375
rect 29121 14364 29155 14375
rect 29193 14364 29227 14375
rect 29265 14364 29299 14375
rect 29337 14364 29371 14375
rect 29409 14364 29443 14375
rect 29481 14364 29515 14375
rect 29553 14364 29587 14375
rect 29625 14364 29659 14375
rect 7129 14172 7163 14206
rect 13084 11231 13118 11265
rect 13157 11231 13191 11265
rect 13230 11231 13264 11265
rect 13303 11255 13313 11265
rect 13313 11255 13337 11265
rect 13376 11255 13381 11265
rect 13381 11255 13410 11265
rect 13303 11231 13337 11255
rect 13376 11231 13410 11255
rect 13449 11231 13483 11265
rect 13522 11255 13551 11265
rect 13551 11255 13556 11265
rect 13595 11255 13619 11265
rect 13619 11255 13629 11265
rect 13668 11255 13687 11265
rect 13687 11255 13702 11265
rect 13741 11255 13755 11265
rect 13755 11255 13775 11265
rect 13814 11255 13823 11265
rect 13823 11255 13848 11265
rect 13887 11255 13891 11265
rect 13891 11255 13921 11265
rect 13960 11255 13993 11265
rect 13993 11255 13994 11265
rect 14033 11255 14061 11265
rect 14061 11255 14067 11265
rect 14106 11255 14129 11265
rect 14129 11255 14140 11265
rect 14179 11255 14197 11265
rect 14197 11255 14213 11265
rect 14252 11255 14265 11265
rect 14265 11255 14286 11265
rect 14325 11255 14333 11265
rect 14333 11255 14359 11265
rect 14398 11255 14401 11265
rect 14401 11255 14432 11265
rect 14471 11255 14503 11265
rect 14503 11255 14505 11265
rect 14544 11255 14571 11265
rect 14571 11255 14578 11265
rect 14617 11255 14639 11265
rect 14639 11255 14651 11265
rect 14690 11255 14707 11265
rect 14707 11255 14724 11265
rect 14763 11255 14775 11265
rect 14775 11255 14797 11265
rect 14836 11255 14843 11265
rect 14843 11255 14870 11265
rect 14909 11255 14911 11265
rect 14911 11255 14943 11265
rect 14982 11255 15013 11265
rect 15013 11255 15016 11265
rect 15055 11255 15081 11265
rect 15081 11255 15089 11265
rect 15128 11255 15149 11265
rect 15149 11255 15162 11265
rect 15201 11255 15217 11265
rect 15217 11255 15235 11265
rect 15273 11255 15285 11265
rect 15285 11255 15307 11265
rect 15345 11255 15353 11265
rect 15353 11255 15379 11265
rect 15417 11255 15421 11265
rect 15421 11255 15451 11265
rect 13522 11231 13556 11255
rect 13595 11231 13629 11255
rect 13668 11231 13702 11255
rect 13741 11231 13775 11255
rect 13814 11231 13848 11255
rect 13887 11231 13921 11255
rect 13960 11231 13994 11255
rect 14033 11231 14067 11255
rect 14106 11231 14140 11255
rect 14179 11231 14213 11255
rect 14252 11231 14286 11255
rect 14325 11231 14359 11255
rect 14398 11231 14432 11255
rect 14471 11231 14505 11255
rect 14544 11231 14578 11255
rect 14617 11231 14651 11255
rect 14690 11231 14724 11255
rect 14763 11231 14797 11255
rect 14836 11231 14870 11255
rect 14909 11231 14943 11255
rect 14982 11231 15016 11255
rect 15055 11231 15089 11255
rect 15128 11231 15162 11255
rect 15201 11231 15235 11255
rect 15273 11231 15307 11255
rect 15345 11231 15379 11255
rect 15417 11231 15451 11255
rect 15489 11231 15523 11265
rect 15561 11255 15591 11265
rect 15591 11255 15595 11265
rect 15633 11255 15659 11265
rect 15659 11255 15667 11265
rect 15705 11255 15727 11265
rect 15727 11255 15739 11265
rect 15777 11255 15795 11265
rect 15795 11255 15811 11265
rect 15561 11231 15595 11255
rect 15633 11231 15667 11255
rect 15705 11231 15739 11255
rect 15777 11231 15811 11255
rect 15849 11231 15883 11265
rect 15921 11231 15955 11265
rect 4433 10918 4463 10937
rect 4463 10918 4467 10937
rect 4507 10918 4531 10937
rect 4531 10918 4541 10937
rect 4581 10918 4599 10937
rect 4599 10918 4615 10937
rect 4655 10918 4667 10937
rect 4667 10918 4689 10937
rect 4729 10918 4735 10937
rect 4735 10918 4763 10937
rect 4433 10903 4467 10918
rect 4507 10903 4541 10918
rect 4581 10903 4615 10918
rect 4655 10903 4689 10918
rect 4729 10903 4763 10918
rect 4803 10903 4837 10937
rect 4876 10918 4905 10937
rect 4905 10918 4910 10937
rect 4949 10918 4973 10937
rect 4973 10918 4983 10937
rect 5022 10918 5041 10937
rect 5041 10918 5056 10937
rect 5095 10918 5109 10937
rect 5109 10918 5129 10937
rect 5168 10918 5177 10937
rect 5177 10918 5202 10937
rect 5241 10918 5245 10937
rect 5245 10918 5275 10937
rect 5314 10918 5347 10937
rect 5347 10918 5348 10937
rect 5387 10918 5415 10937
rect 5415 10918 5421 10937
rect 5460 10918 5483 10937
rect 5483 10918 5494 10937
rect 5533 10918 5551 10937
rect 5551 10918 5567 10937
rect 5606 10918 5619 10937
rect 5619 10918 5640 10937
rect 5679 10918 5687 10937
rect 5687 10918 5713 10937
rect 5752 10918 5755 10937
rect 5755 10918 5786 10937
rect 5825 10918 5857 10937
rect 5857 10918 5859 10937
rect 5898 10918 5925 10937
rect 5925 10918 5932 10937
rect 5971 10918 5993 10937
rect 5993 10918 6005 10937
rect 6044 10918 6061 10937
rect 6061 10918 6078 10937
rect 6117 10918 6129 10937
rect 6129 10918 6151 10937
rect 6190 10918 6197 10937
rect 6197 10918 6224 10937
rect 4876 10903 4910 10918
rect 4949 10903 4983 10918
rect 5022 10903 5056 10918
rect 5095 10903 5129 10918
rect 5168 10903 5202 10918
rect 5241 10903 5275 10918
rect 5314 10903 5348 10918
rect 5387 10903 5421 10918
rect 5460 10903 5494 10918
rect 5533 10903 5567 10918
rect 5606 10903 5640 10918
rect 5679 10903 5713 10918
rect 5752 10903 5786 10918
rect 5825 10903 5859 10918
rect 5898 10903 5932 10918
rect 5971 10903 6005 10918
rect 6044 10903 6078 10918
rect 6117 10903 6151 10918
rect 6190 10903 6224 10918
rect 4433 10849 4463 10861
rect 4463 10849 4467 10861
rect 4507 10849 4531 10861
rect 4531 10849 4541 10861
rect 4581 10849 4599 10861
rect 4599 10849 4615 10861
rect 4655 10849 4667 10861
rect 4667 10849 4689 10861
rect 4729 10849 4735 10861
rect 4735 10849 4763 10861
rect 4433 10827 4467 10849
rect 4507 10827 4541 10849
rect 4581 10827 4615 10849
rect 4655 10827 4689 10849
rect 4729 10827 4763 10849
rect 4803 10827 4837 10861
rect 4876 10849 4905 10861
rect 4905 10849 4910 10861
rect 4949 10849 4973 10861
rect 4973 10849 4983 10861
rect 5022 10849 5041 10861
rect 5041 10849 5056 10861
rect 5095 10849 5109 10861
rect 5109 10849 5129 10861
rect 5168 10849 5177 10861
rect 5177 10849 5202 10861
rect 5241 10849 5245 10861
rect 5245 10849 5275 10861
rect 5314 10849 5347 10861
rect 5347 10849 5348 10861
rect 5387 10849 5415 10861
rect 5415 10849 5421 10861
rect 5460 10849 5483 10861
rect 5483 10849 5494 10861
rect 5533 10849 5551 10861
rect 5551 10849 5567 10861
rect 5606 10849 5619 10861
rect 5619 10849 5640 10861
rect 5679 10849 5687 10861
rect 5687 10849 5713 10861
rect 5752 10849 5755 10861
rect 5755 10849 5786 10861
rect 5825 10849 5857 10861
rect 5857 10849 5859 10861
rect 5898 10849 5925 10861
rect 5925 10849 5932 10861
rect 5971 10849 5993 10861
rect 5993 10849 6005 10861
rect 6044 10849 6061 10861
rect 6061 10849 6078 10861
rect 6117 10849 6129 10861
rect 6129 10849 6151 10861
rect 6190 10849 6197 10861
rect 6197 10849 6224 10861
rect 13364 10905 13381 10934
rect 13381 10905 13398 10934
rect 13438 10905 13449 10934
rect 13449 10905 13472 10934
rect 13512 10905 13517 10934
rect 13517 10905 13546 10934
rect 13364 10900 13398 10905
rect 13438 10900 13472 10905
rect 13512 10900 13546 10905
rect 13585 10900 13619 10934
rect 13658 10905 13687 10934
rect 13687 10905 13692 10934
rect 13731 10905 13755 10934
rect 13755 10905 13765 10934
rect 13804 10905 13823 10934
rect 13823 10905 13838 10934
rect 13877 10905 13891 10934
rect 13891 10905 13911 10934
rect 13950 10905 13959 10934
rect 13959 10905 13984 10934
rect 14023 10905 14027 10934
rect 14027 10905 14057 10934
rect 14096 10905 14129 10934
rect 14129 10905 14130 10934
rect 14169 10905 14197 10934
rect 14197 10905 14203 10934
rect 14242 10905 14265 10934
rect 14265 10905 14276 10934
rect 14315 10905 14333 10934
rect 14333 10905 14349 10934
rect 14388 10905 14401 10934
rect 14401 10905 14422 10934
rect 14461 10905 14469 10934
rect 14469 10905 14495 10934
rect 14534 10905 14537 10934
rect 14537 10905 14568 10934
rect 14607 10905 14639 10934
rect 14639 10905 14641 10934
rect 14680 10905 14707 10934
rect 14707 10905 14714 10934
rect 14753 10905 14775 10934
rect 14775 10905 14787 10934
rect 14826 10905 14843 10934
rect 14843 10905 14860 10934
rect 14899 10905 14911 10934
rect 14911 10905 14933 10934
rect 14972 10905 14979 10934
rect 14979 10905 15006 10934
rect 15045 10905 15047 10934
rect 15047 10905 15079 10934
rect 15118 10905 15149 10934
rect 15149 10905 15152 10934
rect 15191 10905 15217 10934
rect 15217 10905 15225 10934
rect 15264 10905 15285 10934
rect 15285 10905 15298 10934
rect 15337 10905 15353 10934
rect 15353 10905 15371 10934
rect 15410 10905 15421 10934
rect 15421 10905 15444 10934
rect 15483 10905 15489 10934
rect 15489 10905 15517 10934
rect 15556 10905 15557 10934
rect 15557 10905 15590 10934
rect 15629 10905 15659 10934
rect 15659 10905 15663 10934
rect 15702 10905 15727 10934
rect 15727 10905 15736 10934
rect 15775 10905 15795 10934
rect 15795 10905 15809 10934
rect 13658 10900 13692 10905
rect 13731 10900 13765 10905
rect 13804 10900 13838 10905
rect 13877 10900 13911 10905
rect 13950 10900 13984 10905
rect 14023 10900 14057 10905
rect 14096 10900 14130 10905
rect 14169 10900 14203 10905
rect 14242 10900 14276 10905
rect 14315 10900 14349 10905
rect 14388 10900 14422 10905
rect 14461 10900 14495 10905
rect 14534 10900 14568 10905
rect 14607 10900 14641 10905
rect 14680 10900 14714 10905
rect 14753 10900 14787 10905
rect 14826 10900 14860 10905
rect 14899 10900 14933 10905
rect 14972 10900 15006 10905
rect 15045 10900 15079 10905
rect 15118 10900 15152 10905
rect 15191 10900 15225 10905
rect 15264 10900 15298 10905
rect 15337 10900 15371 10905
rect 15410 10900 15444 10905
rect 15483 10900 15517 10905
rect 15556 10900 15590 10905
rect 15629 10900 15663 10905
rect 15702 10900 15736 10905
rect 15775 10900 15809 10905
rect 15848 10900 15882 10934
rect 4876 10827 4910 10849
rect 4949 10827 4983 10849
rect 5022 10827 5056 10849
rect 5095 10827 5129 10849
rect 5168 10827 5202 10849
rect 5241 10827 5275 10849
rect 5314 10827 5348 10849
rect 5387 10827 5421 10849
rect 5460 10827 5494 10849
rect 5533 10827 5567 10849
rect 5606 10827 5640 10849
rect 5679 10827 5713 10849
rect 5752 10827 5786 10849
rect 5825 10827 5859 10849
rect 5898 10827 5932 10849
rect 5971 10827 6005 10849
rect 6044 10827 6078 10849
rect 6117 10827 6151 10849
rect 6190 10827 6224 10849
rect 4433 10780 4463 10785
rect 4463 10780 4467 10785
rect 4507 10780 4531 10785
rect 4531 10780 4541 10785
rect 4581 10780 4599 10785
rect 4599 10780 4615 10785
rect 4655 10780 4667 10785
rect 4667 10780 4689 10785
rect 4729 10780 4735 10785
rect 4735 10780 4763 10785
rect 4433 10751 4467 10780
rect 4507 10751 4541 10780
rect 4581 10751 4615 10780
rect 4655 10751 4689 10780
rect 4729 10751 4763 10780
rect 4803 10751 4837 10785
rect 4876 10780 4905 10785
rect 4905 10780 4910 10785
rect 4949 10780 4973 10785
rect 4973 10780 4983 10785
rect 5022 10780 5041 10785
rect 5041 10780 5056 10785
rect 5095 10780 5109 10785
rect 5109 10780 5129 10785
rect 5168 10780 5177 10785
rect 5177 10780 5202 10785
rect 5241 10780 5245 10785
rect 5245 10780 5275 10785
rect 5314 10780 5347 10785
rect 5347 10780 5348 10785
rect 5387 10780 5415 10785
rect 5415 10780 5421 10785
rect 5460 10780 5483 10785
rect 5483 10780 5494 10785
rect 5533 10780 5551 10785
rect 5551 10780 5567 10785
rect 5606 10780 5619 10785
rect 5619 10780 5640 10785
rect 5679 10780 5687 10785
rect 5687 10780 5713 10785
rect 5752 10780 5755 10785
rect 5755 10780 5786 10785
rect 5825 10780 5857 10785
rect 5857 10780 5859 10785
rect 5898 10780 5925 10785
rect 5925 10780 5932 10785
rect 5971 10780 5993 10785
rect 5993 10780 6005 10785
rect 6044 10780 6061 10785
rect 6061 10780 6078 10785
rect 6117 10780 6129 10785
rect 6129 10780 6151 10785
rect 6190 10780 6197 10785
rect 6197 10780 6224 10785
rect 4876 10751 4910 10780
rect 4949 10751 4983 10780
rect 5022 10751 5056 10780
rect 5095 10751 5129 10780
rect 5168 10751 5202 10780
rect 5241 10751 5275 10780
rect 5314 10751 5348 10780
rect 5387 10751 5421 10780
rect 5460 10751 5494 10780
rect 5533 10751 5567 10780
rect 5606 10751 5640 10780
rect 5679 10751 5713 10780
rect 5752 10751 5786 10780
rect 5825 10751 5859 10780
rect 5898 10751 5932 10780
rect 5971 10751 6005 10780
rect 6044 10751 6078 10780
rect 6117 10751 6151 10780
rect 6190 10751 6224 10780
rect 13364 10835 13381 10860
rect 13381 10835 13398 10860
rect 13438 10835 13449 10860
rect 13449 10835 13472 10860
rect 13512 10835 13517 10860
rect 13517 10835 13546 10860
rect 13364 10826 13398 10835
rect 13438 10826 13472 10835
rect 13512 10826 13546 10835
rect 13585 10826 13619 10860
rect 13658 10835 13687 10860
rect 13687 10835 13692 10860
rect 13731 10835 13755 10860
rect 13755 10835 13765 10860
rect 13804 10835 13823 10860
rect 13823 10835 13838 10860
rect 13877 10835 13891 10860
rect 13891 10835 13911 10860
rect 13950 10835 13959 10860
rect 13959 10835 13984 10860
rect 14023 10835 14027 10860
rect 14027 10835 14057 10860
rect 14096 10835 14129 10860
rect 14129 10835 14130 10860
rect 14169 10835 14197 10860
rect 14197 10835 14203 10860
rect 14242 10835 14265 10860
rect 14265 10835 14276 10860
rect 14315 10835 14333 10860
rect 14333 10835 14349 10860
rect 14388 10835 14401 10860
rect 14401 10835 14422 10860
rect 14461 10835 14469 10860
rect 14469 10835 14495 10860
rect 14534 10835 14537 10860
rect 14537 10835 14568 10860
rect 14607 10835 14639 10860
rect 14639 10835 14641 10860
rect 14680 10835 14707 10860
rect 14707 10835 14714 10860
rect 14753 10835 14775 10860
rect 14775 10835 14787 10860
rect 14826 10835 14843 10860
rect 14843 10835 14860 10860
rect 14899 10835 14911 10860
rect 14911 10835 14933 10860
rect 14972 10835 14979 10860
rect 14979 10835 15006 10860
rect 15045 10835 15047 10860
rect 15047 10835 15079 10860
rect 15118 10835 15149 10860
rect 15149 10835 15152 10860
rect 15191 10835 15217 10860
rect 15217 10835 15225 10860
rect 15264 10835 15285 10860
rect 15285 10835 15298 10860
rect 15337 10835 15353 10860
rect 15353 10835 15371 10860
rect 15410 10835 15421 10860
rect 15421 10835 15444 10860
rect 15483 10835 15489 10860
rect 15489 10835 15517 10860
rect 15556 10835 15557 10860
rect 15557 10835 15590 10860
rect 15629 10835 15659 10860
rect 15659 10835 15663 10860
rect 15702 10835 15727 10860
rect 15727 10835 15736 10860
rect 15775 10835 15795 10860
rect 15795 10835 15809 10860
rect 13658 10826 13692 10835
rect 13731 10826 13765 10835
rect 13804 10826 13838 10835
rect 13877 10826 13911 10835
rect 13950 10826 13984 10835
rect 14023 10826 14057 10835
rect 14096 10826 14130 10835
rect 14169 10826 14203 10835
rect 14242 10826 14276 10835
rect 14315 10826 14349 10835
rect 14388 10826 14422 10835
rect 14461 10826 14495 10835
rect 14534 10826 14568 10835
rect 14607 10826 14641 10835
rect 14680 10826 14714 10835
rect 14753 10826 14787 10835
rect 14826 10826 14860 10835
rect 14899 10826 14933 10835
rect 14972 10826 15006 10835
rect 15045 10826 15079 10835
rect 15118 10826 15152 10835
rect 15191 10826 15225 10835
rect 15264 10826 15298 10835
rect 15337 10826 15371 10835
rect 15410 10826 15444 10835
rect 15483 10826 15517 10835
rect 15556 10826 15590 10835
rect 15629 10826 15663 10835
rect 15702 10826 15736 10835
rect 15775 10826 15809 10835
rect 15848 10826 15882 10860
rect 13364 10765 13381 10786
rect 13381 10765 13398 10786
rect 13438 10765 13449 10786
rect 13449 10765 13472 10786
rect 13512 10765 13517 10786
rect 13517 10765 13546 10786
rect 13364 10752 13398 10765
rect 13438 10752 13472 10765
rect 13512 10752 13546 10765
rect 13585 10752 13619 10786
rect 13658 10765 13687 10786
rect 13687 10765 13692 10786
rect 13731 10765 13755 10786
rect 13755 10765 13765 10786
rect 13804 10765 13823 10786
rect 13823 10765 13838 10786
rect 13877 10765 13891 10786
rect 13891 10765 13911 10786
rect 13950 10765 13959 10786
rect 13959 10765 13984 10786
rect 14023 10765 14027 10786
rect 14027 10765 14057 10786
rect 14096 10765 14129 10786
rect 14129 10765 14130 10786
rect 14169 10765 14197 10786
rect 14197 10765 14203 10786
rect 14242 10765 14265 10786
rect 14265 10765 14276 10786
rect 14315 10765 14333 10786
rect 14333 10765 14349 10786
rect 14388 10765 14401 10786
rect 14401 10765 14422 10786
rect 14461 10765 14469 10786
rect 14469 10765 14495 10786
rect 14534 10765 14537 10786
rect 14537 10765 14568 10786
rect 14607 10765 14639 10786
rect 14639 10765 14641 10786
rect 14680 10765 14707 10786
rect 14707 10765 14714 10786
rect 14753 10765 14775 10786
rect 14775 10765 14787 10786
rect 14826 10765 14843 10786
rect 14843 10765 14860 10786
rect 14899 10765 14911 10786
rect 14911 10765 14933 10786
rect 14972 10765 14979 10786
rect 14979 10765 15006 10786
rect 15045 10765 15047 10786
rect 15047 10765 15079 10786
rect 15118 10765 15149 10786
rect 15149 10765 15152 10786
rect 15191 10765 15217 10786
rect 15217 10765 15225 10786
rect 15264 10765 15285 10786
rect 15285 10765 15298 10786
rect 15337 10765 15353 10786
rect 15353 10765 15371 10786
rect 15410 10765 15421 10786
rect 15421 10765 15444 10786
rect 15483 10765 15489 10786
rect 15489 10765 15517 10786
rect 15556 10765 15557 10786
rect 15557 10765 15590 10786
rect 15629 10765 15659 10786
rect 15659 10765 15663 10786
rect 15702 10765 15727 10786
rect 15727 10765 15736 10786
rect 15775 10765 15795 10786
rect 15795 10765 15809 10786
rect 13658 10752 13692 10765
rect 13731 10752 13765 10765
rect 13804 10752 13838 10765
rect 13877 10752 13911 10765
rect 13950 10752 13984 10765
rect 14023 10752 14057 10765
rect 14096 10752 14130 10765
rect 14169 10752 14203 10765
rect 14242 10752 14276 10765
rect 14315 10752 14349 10765
rect 14388 10752 14422 10765
rect 14461 10752 14495 10765
rect 14534 10752 14568 10765
rect 14607 10752 14641 10765
rect 14680 10752 14714 10765
rect 14753 10752 14787 10765
rect 14826 10752 14860 10765
rect 14899 10752 14933 10765
rect 14972 10752 15006 10765
rect 15045 10752 15079 10765
rect 15118 10752 15152 10765
rect 15191 10752 15225 10765
rect 15264 10752 15298 10765
rect 15337 10752 15371 10765
rect 15410 10752 15444 10765
rect 15483 10752 15517 10765
rect 15556 10752 15590 10765
rect 15629 10752 15663 10765
rect 15702 10752 15736 10765
rect 15775 10752 15809 10765
rect 15848 10752 15882 10786
rect 13116 10508 13150 10542
rect 13190 10508 13224 10542
rect 13264 10519 13298 10542
rect 13338 10519 13372 10542
rect 13412 10519 13446 10542
rect 13486 10519 13520 10542
rect 13560 10519 13594 10542
rect 13634 10519 13668 10542
rect 13708 10519 13742 10542
rect 13782 10519 13816 10542
rect 13856 10519 13890 10542
rect 13930 10519 13964 10542
rect 14004 10519 14038 10542
rect 14078 10519 14112 10542
rect 14152 10519 14186 10542
rect 14226 10519 14260 10542
rect 14300 10519 14334 10542
rect 14374 10519 14408 10542
rect 14448 10519 14482 10542
rect 14522 10519 14556 10542
rect 14596 10519 14630 10542
rect 14670 10519 14704 10542
rect 14744 10519 14778 10542
rect 14818 10519 14852 10542
rect 14892 10519 14926 10542
rect 14966 10519 15000 10542
rect 15040 10519 15074 10542
rect 15114 10519 15148 10542
rect 15188 10519 15222 10542
rect 15261 10519 15295 10542
rect 15334 10519 15368 10542
rect 15407 10519 15441 10542
rect 15480 10519 15514 10542
rect 15553 10519 15587 10542
rect 15626 10519 15660 10542
rect 15699 10519 15733 10542
rect 13264 10508 13279 10519
rect 13279 10508 13298 10519
rect 13338 10508 13347 10519
rect 13347 10508 13372 10519
rect 13412 10508 13415 10519
rect 13415 10508 13446 10519
rect 13486 10508 13517 10519
rect 13517 10508 13520 10519
rect 13560 10508 13585 10519
rect 13585 10508 13594 10519
rect 13634 10508 13653 10519
rect 13653 10508 13668 10519
rect 13708 10508 13721 10519
rect 13721 10508 13742 10519
rect 13782 10508 13789 10519
rect 13789 10508 13816 10519
rect 13856 10508 13857 10519
rect 13857 10508 13890 10519
rect 13930 10508 13959 10519
rect 13959 10508 13964 10519
rect 14004 10508 14027 10519
rect 14027 10508 14038 10519
rect 14078 10508 14095 10519
rect 14095 10508 14112 10519
rect 14152 10508 14163 10519
rect 14163 10508 14186 10519
rect 14226 10508 14231 10519
rect 14231 10508 14260 10519
rect 14300 10508 14333 10519
rect 14333 10508 14334 10519
rect 14374 10508 14401 10519
rect 14401 10508 14408 10519
rect 14448 10508 14469 10519
rect 14469 10508 14482 10519
rect 14522 10508 14537 10519
rect 14537 10508 14556 10519
rect 14596 10508 14605 10519
rect 14605 10508 14630 10519
rect 14670 10508 14673 10519
rect 14673 10508 14704 10519
rect 14744 10508 14775 10519
rect 14775 10508 14778 10519
rect 14818 10508 14843 10519
rect 14843 10508 14852 10519
rect 14892 10508 14911 10519
rect 14911 10508 14926 10519
rect 14966 10508 14979 10519
rect 14979 10508 15000 10519
rect 15040 10508 15047 10519
rect 15047 10508 15074 10519
rect 15114 10508 15115 10519
rect 15115 10508 15148 10519
rect 15188 10508 15217 10519
rect 15217 10508 15222 10519
rect 15261 10508 15285 10519
rect 15285 10508 15295 10519
rect 15334 10508 15353 10519
rect 15353 10508 15368 10519
rect 15407 10508 15421 10519
rect 15421 10508 15441 10519
rect 15480 10508 15489 10519
rect 15489 10508 15514 10519
rect 15553 10508 15557 10519
rect 15557 10508 15587 10519
rect 15626 10508 15659 10519
rect 15659 10508 15660 10519
rect 15699 10508 15727 10519
rect 15727 10508 15733 10519
<< metal1 >>
rect -2842 50607 -262 50619
rect -2842 37901 -2829 50607
rect -275 37901 -262 50607
rect 645 43689 1083 43695
rect 645 43637 646 43689
rect 698 43637 710 43689
rect 762 43637 774 43689
rect 826 43637 838 43689
rect 890 43637 902 43689
rect 954 43637 966 43689
rect 1018 43637 1030 43689
rect 1082 43637 1083 43689
rect 645 43623 1083 43637
rect 645 43571 646 43623
rect 698 43571 710 43623
rect 762 43571 774 43623
rect 826 43571 838 43623
rect 890 43571 902 43623
rect 954 43571 966 43623
rect 1018 43571 1030 43623
rect 1082 43571 1083 43623
rect 645 43557 1083 43571
rect 645 43505 646 43557
rect 698 43505 710 43557
rect 762 43505 774 43557
rect 826 43505 838 43557
rect 890 43505 902 43557
rect 954 43505 966 43557
rect 1018 43505 1030 43557
rect 1082 43505 1083 43557
rect 645 43491 1083 43505
rect 645 43439 646 43491
rect 698 43439 710 43491
rect 762 43439 774 43491
rect 826 43439 838 43491
rect 890 43439 902 43491
rect 954 43439 966 43491
rect 1018 43439 1030 43491
rect 1082 43439 1083 43491
rect 645 43425 1083 43439
rect 645 43373 646 43425
rect 698 43373 710 43425
rect 762 43373 774 43425
rect 826 43373 838 43425
rect 890 43373 902 43425
rect 954 43373 966 43425
rect 1018 43373 1030 43425
rect 1082 43373 1083 43425
rect 645 43359 1083 43373
rect 645 43307 646 43359
rect 698 43307 710 43359
rect 762 43307 774 43359
rect 826 43307 838 43359
rect 890 43307 902 43359
rect 954 43307 966 43359
rect 1018 43307 1030 43359
rect 1082 43307 1083 43359
rect 645 43293 1083 43307
rect 645 43241 646 43293
rect 698 43241 710 43293
rect 762 43241 774 43293
rect 826 43241 838 43293
rect 890 43241 902 43293
rect 954 43241 966 43293
rect 1018 43241 1030 43293
rect 1082 43241 1083 43293
rect 645 43226 1083 43241
rect 645 43174 646 43226
rect 698 43174 710 43226
rect 762 43174 774 43226
rect 826 43174 838 43226
rect 890 43174 902 43226
rect 954 43174 966 43226
rect 1018 43174 1030 43226
rect 1082 43174 1083 43226
rect 645 43168 1083 43174
tri 24138 40260 24144 40266 se
rect 24144 40260 24149 40266
rect 31407 40072 31413 40188
rect 31529 40136 32301 40188
rect 31529 40072 31535 40136
tri 31535 40072 31599 40136 nw
rect 31593 39827 31599 39943
rect 31715 39897 32301 39943
rect 31715 39827 31721 39897
tri 31721 39827 31791 39897 nw
rect -2842 37862 -262 37901
rect -2842 37828 -2829 37862
rect -2795 37828 -2757 37862
rect -2723 37828 -2685 37862
rect -2651 37828 -2613 37862
rect -2579 37828 -2541 37862
rect -2507 37828 -2469 37862
rect -2435 37828 -2397 37862
rect -2363 37828 -2325 37862
rect -2291 37828 -2253 37862
rect -2219 37828 -2181 37862
rect -2147 37828 -2109 37862
rect -2075 37828 -2037 37862
rect -2003 37828 -1965 37862
rect -1931 37828 -1893 37862
rect -1859 37828 -1821 37862
rect -1787 37828 -1749 37862
rect -1715 37828 -1677 37862
rect -1643 37828 -1605 37862
rect -1571 37828 -1533 37862
rect -1499 37828 -1461 37862
rect -1427 37828 -1389 37862
rect -1355 37828 -1317 37862
rect -1283 37828 -1245 37862
rect -1211 37828 -1173 37862
rect -1139 37828 -1101 37862
rect -1067 37828 -1029 37862
rect -995 37828 -957 37862
rect -923 37828 -885 37862
rect -851 37828 -813 37862
rect -779 37828 -741 37862
rect -707 37828 -669 37862
rect -635 37828 -597 37862
rect -563 37828 -525 37862
rect -491 37828 -453 37862
rect -419 37828 -381 37862
rect -347 37828 -309 37862
rect -275 37828 -262 37862
rect -2842 37789 -262 37828
rect -2842 37755 -2829 37789
rect -2795 37755 -2757 37789
rect -2723 37755 -2685 37789
rect -2651 37755 -2613 37789
rect -2579 37755 -2541 37789
rect -2507 37755 -2469 37789
rect -2435 37755 -2397 37789
rect -2363 37755 -2325 37789
rect -2291 37755 -2253 37789
rect -2219 37755 -2181 37789
rect -2147 37755 -2109 37789
rect -2075 37755 -2037 37789
rect -2003 37755 -1965 37789
rect -1931 37755 -1893 37789
rect -1859 37755 -1821 37789
rect -1787 37755 -1749 37789
rect -1715 37755 -1677 37789
rect -1643 37755 -1605 37789
rect -1571 37755 -1533 37789
rect -1499 37755 -1461 37789
rect -1427 37755 -1389 37789
rect -1355 37755 -1317 37789
rect -1283 37755 -1245 37789
rect -1211 37755 -1173 37789
rect -1139 37755 -1101 37789
rect -1067 37755 -1029 37789
rect -995 37755 -957 37789
rect -923 37755 -885 37789
rect -851 37755 -813 37789
rect -779 37755 -741 37789
rect -707 37755 -669 37789
rect -635 37755 -597 37789
rect -563 37755 -525 37789
rect -491 37755 -453 37789
rect -419 37755 -381 37789
rect -347 37755 -309 37789
rect -275 37755 -262 37789
rect -2842 37716 -262 37755
rect -2842 37682 -2829 37716
rect -2795 37682 -2757 37716
rect -2723 37682 -2685 37716
rect -2651 37682 -2613 37716
rect -2579 37682 -2541 37716
rect -2507 37682 -2469 37716
rect -2435 37682 -2397 37716
rect -2363 37682 -2325 37716
rect -2291 37682 -2253 37716
rect -2219 37682 -2181 37716
rect -2147 37682 -2109 37716
rect -2075 37682 -2037 37716
rect -2003 37682 -1965 37716
rect -1931 37682 -1893 37716
rect -1859 37682 -1821 37716
rect -1787 37682 -1749 37716
rect -1715 37682 -1677 37716
rect -1643 37682 -1605 37716
rect -1571 37682 -1533 37716
rect -1499 37682 -1461 37716
rect -1427 37682 -1389 37716
rect -1355 37682 -1317 37716
rect -1283 37682 -1245 37716
rect -1211 37682 -1173 37716
rect -1139 37682 -1101 37716
rect -1067 37682 -1029 37716
rect -995 37682 -957 37716
rect -923 37682 -885 37716
rect -851 37682 -813 37716
rect -779 37682 -741 37716
rect -707 37682 -669 37716
rect -635 37682 -597 37716
rect -563 37682 -525 37716
rect -491 37682 -453 37716
rect -419 37682 -381 37716
rect -347 37682 -309 37716
rect -275 37682 -262 37716
rect -2842 37643 -262 37682
rect -2842 37609 -2829 37643
rect -2795 37609 -2757 37643
rect -2723 37609 -2685 37643
rect -2651 37609 -2613 37643
rect -2579 37609 -2541 37643
rect -2507 37609 -2469 37643
rect -2435 37609 -2397 37643
rect -2363 37609 -2325 37643
rect -2291 37609 -2253 37643
rect -2219 37609 -2181 37643
rect -2147 37609 -2109 37643
rect -2075 37609 -2037 37643
rect -2003 37609 -1965 37643
rect -1931 37609 -1893 37643
rect -1859 37609 -1821 37643
rect -1787 37609 -1749 37643
rect -1715 37609 -1677 37643
rect -1643 37609 -1605 37643
rect -1571 37609 -1533 37643
rect -1499 37609 -1461 37643
rect -1427 37609 -1389 37643
rect -1355 37609 -1317 37643
rect -1283 37609 -1245 37643
rect -1211 37609 -1173 37643
rect -1139 37609 -1101 37643
rect -1067 37609 -1029 37643
rect -995 37609 -957 37643
rect -923 37609 -885 37643
rect -851 37609 -813 37643
rect -779 37609 -741 37643
rect -707 37609 -669 37643
rect -635 37609 -597 37643
rect -563 37609 -525 37643
rect -491 37609 -453 37643
rect -419 37609 -381 37643
rect -347 37609 -309 37643
rect -275 37609 -262 37643
rect -2842 37570 -262 37609
rect -2842 37536 -2829 37570
rect -2795 37536 -2757 37570
rect -2723 37536 -2685 37570
rect -2651 37536 -2613 37570
rect -2579 37536 -2541 37570
rect -2507 37536 -2469 37570
rect -2435 37536 -2397 37570
rect -2363 37536 -2325 37570
rect -2291 37536 -2253 37570
rect -2219 37536 -2181 37570
rect -2147 37536 -2109 37570
rect -2075 37536 -2037 37570
rect -2003 37536 -1965 37570
rect -1931 37536 -1893 37570
rect -1859 37536 -1821 37570
rect -1787 37536 -1749 37570
rect -1715 37536 -1677 37570
rect -1643 37536 -1605 37570
rect -1571 37536 -1533 37570
rect -1499 37536 -1461 37570
rect -1427 37536 -1389 37570
rect -1355 37536 -1317 37570
rect -1283 37536 -1245 37570
rect -1211 37536 -1173 37570
rect -1139 37536 -1101 37570
rect -1067 37536 -1029 37570
rect -995 37536 -957 37570
rect -923 37536 -885 37570
rect -851 37536 -813 37570
rect -779 37536 -741 37570
rect -707 37536 -669 37570
rect -635 37536 -597 37570
rect -563 37536 -525 37570
rect -491 37536 -453 37570
rect -419 37536 -381 37570
rect -347 37536 -309 37570
rect -275 37536 -262 37570
rect -2842 37497 -262 37536
rect -2842 37463 -2829 37497
rect -2795 37463 -2757 37497
rect -2723 37463 -2685 37497
rect -2651 37463 -2613 37497
rect -2579 37463 -2541 37497
rect -2507 37463 -2469 37497
rect -2435 37463 -2397 37497
rect -2363 37463 -2325 37497
rect -2291 37463 -2253 37497
rect -2219 37463 -2181 37497
rect -2147 37463 -2109 37497
rect -2075 37463 -2037 37497
rect -2003 37463 -1965 37497
rect -1931 37463 -1893 37497
rect -1859 37463 -1821 37497
rect -1787 37463 -1749 37497
rect -1715 37463 -1677 37497
rect -1643 37463 -1605 37497
rect -1571 37463 -1533 37497
rect -1499 37463 -1461 37497
rect -1427 37463 -1389 37497
rect -1355 37463 -1317 37497
rect -1283 37463 -1245 37497
rect -1211 37463 -1173 37497
rect -1139 37463 -1101 37497
rect -1067 37463 -1029 37497
rect -995 37463 -957 37497
rect -923 37463 -885 37497
rect -851 37463 -813 37497
rect -779 37463 -741 37497
rect -707 37463 -669 37497
rect -635 37463 -597 37497
rect -563 37463 -525 37497
rect -491 37463 -453 37497
rect -419 37463 -381 37497
rect -347 37463 -309 37497
rect -275 37463 -262 37497
rect -2842 37424 -262 37463
rect -2842 37390 -2829 37424
rect -2795 37390 -2757 37424
rect -2723 37390 -2685 37424
rect -2651 37390 -2613 37424
rect -2579 37390 -2541 37424
rect -2507 37390 -2469 37424
rect -2435 37390 -2397 37424
rect -2363 37390 -2325 37424
rect -2291 37390 -2253 37424
rect -2219 37390 -2181 37424
rect -2147 37390 -2109 37424
rect -2075 37390 -2037 37424
rect -2003 37390 -1965 37424
rect -1931 37390 -1893 37424
rect -1859 37390 -1821 37424
rect -1787 37390 -1749 37424
rect -1715 37390 -1677 37424
rect -1643 37390 -1605 37424
rect -1571 37390 -1533 37424
rect -1499 37390 -1461 37424
rect -1427 37390 -1389 37424
rect -1355 37390 -1317 37424
rect -1283 37390 -1245 37424
rect -1211 37390 -1173 37424
rect -1139 37390 -1101 37424
rect -1067 37390 -1029 37424
rect -995 37390 -957 37424
rect -923 37390 -885 37424
rect -851 37390 -813 37424
rect -779 37390 -741 37424
rect -707 37390 -669 37424
rect -635 37390 -597 37424
rect -563 37390 -525 37424
rect -491 37390 -453 37424
rect -419 37390 -381 37424
rect -347 37390 -309 37424
rect -275 37390 -262 37424
rect -2842 37351 -262 37390
rect -2842 37317 -2829 37351
rect -2795 37317 -2757 37351
rect -2723 37317 -2685 37351
rect -2651 37317 -2613 37351
rect -2579 37317 -2541 37351
rect -2507 37317 -2469 37351
rect -2435 37317 -2397 37351
rect -2363 37317 -2325 37351
rect -2291 37317 -2253 37351
rect -2219 37317 -2181 37351
rect -2147 37317 -2109 37351
rect -2075 37317 -2037 37351
rect -2003 37317 -1965 37351
rect -1931 37317 -1893 37351
rect -1859 37317 -1821 37351
rect -1787 37317 -1749 37351
rect -1715 37317 -1677 37351
rect -1643 37317 -1605 37351
rect -1571 37317 -1533 37351
rect -1499 37317 -1461 37351
rect -1427 37317 -1389 37351
rect -1355 37317 -1317 37351
rect -1283 37317 -1245 37351
rect -1211 37317 -1173 37351
rect -1139 37317 -1101 37351
rect -1067 37317 -1029 37351
rect -995 37317 -957 37351
rect -923 37317 -885 37351
rect -851 37317 -813 37351
rect -779 37317 -741 37351
rect -707 37317 -669 37351
rect -635 37317 -597 37351
rect -563 37317 -525 37351
rect -491 37317 -453 37351
rect -419 37317 -381 37351
rect -347 37317 -309 37351
rect -275 37317 -262 37351
rect -2842 37278 -262 37317
rect -2842 37244 -2829 37278
rect -2795 37244 -2757 37278
rect -2723 37244 -2685 37278
rect -2651 37244 -2613 37278
rect -2579 37244 -2541 37278
rect -2507 37244 -2469 37278
rect -2435 37244 -2397 37278
rect -2363 37244 -2325 37278
rect -2291 37244 -2253 37278
rect -2219 37244 -2181 37278
rect -2147 37244 -2109 37278
rect -2075 37244 -2037 37278
rect -2003 37244 -1965 37278
rect -1931 37244 -1893 37278
rect -1859 37244 -1821 37278
rect -1787 37244 -1749 37278
rect -1715 37244 -1677 37278
rect -1643 37244 -1605 37278
rect -1571 37244 -1533 37278
rect -1499 37244 -1461 37278
rect -1427 37244 -1389 37278
rect -1355 37244 -1317 37278
rect -1283 37244 -1245 37278
rect -1211 37244 -1173 37278
rect -1139 37244 -1101 37278
rect -1067 37244 -1029 37278
rect -995 37244 -957 37278
rect -923 37244 -885 37278
rect -851 37244 -813 37278
rect -779 37244 -741 37278
rect -707 37244 -669 37278
rect -635 37244 -597 37278
rect -563 37244 -525 37278
rect -491 37244 -453 37278
rect -419 37244 -381 37278
rect -347 37244 -309 37278
rect -275 37244 -262 37278
rect -2842 37205 -262 37244
rect -2842 37171 -2829 37205
rect -2795 37171 -2757 37205
rect -2723 37171 -2685 37205
rect -2651 37171 -2613 37205
rect -2579 37171 -2541 37205
rect -2507 37171 -2469 37205
rect -2435 37171 -2397 37205
rect -2363 37171 -2325 37205
rect -2291 37171 -2253 37205
rect -2219 37171 -2181 37205
rect -2147 37171 -2109 37205
rect -2075 37171 -2037 37205
rect -2003 37171 -1965 37205
rect -1931 37171 -1893 37205
rect -1859 37171 -1821 37205
rect -1787 37171 -1749 37205
rect -1715 37171 -1677 37205
rect -1643 37171 -1605 37205
rect -1571 37171 -1533 37205
rect -1499 37171 -1461 37205
rect -1427 37171 -1389 37205
rect -1355 37171 -1317 37205
rect -1283 37171 -1245 37205
rect -1211 37171 -1173 37205
rect -1139 37171 -1101 37205
rect -1067 37171 -1029 37205
rect -995 37171 -957 37205
rect -923 37171 -885 37205
rect -851 37171 -813 37205
rect -779 37171 -741 37205
rect -707 37171 -669 37205
rect -635 37171 -597 37205
rect -563 37171 -525 37205
rect -491 37171 -453 37205
rect -419 37171 -381 37205
rect -347 37171 -309 37205
rect -275 37171 -262 37205
rect -2842 37132 -262 37171
rect -2842 37098 -2829 37132
rect -2795 37098 -2757 37132
rect -2723 37098 -2685 37132
rect -2651 37098 -2613 37132
rect -2579 37098 -2541 37132
rect -2507 37098 -2469 37132
rect -2435 37098 -2397 37132
rect -2363 37098 -2325 37132
rect -2291 37098 -2253 37132
rect -2219 37098 -2181 37132
rect -2147 37098 -2109 37132
rect -2075 37098 -2037 37132
rect -2003 37098 -1965 37132
rect -1931 37098 -1893 37132
rect -1859 37098 -1821 37132
rect -1787 37098 -1749 37132
rect -1715 37098 -1677 37132
rect -1643 37098 -1605 37132
rect -1571 37098 -1533 37132
rect -1499 37098 -1461 37132
rect -1427 37098 -1389 37132
rect -1355 37098 -1317 37132
rect -1283 37098 -1245 37132
rect -1211 37098 -1173 37132
rect -1139 37098 -1101 37132
rect -1067 37098 -1029 37132
rect -995 37098 -957 37132
rect -923 37098 -885 37132
rect -851 37098 -813 37132
rect -779 37098 -741 37132
rect -707 37098 -669 37132
rect -635 37098 -597 37132
rect -563 37098 -525 37132
rect -491 37098 -453 37132
rect -419 37098 -381 37132
rect -347 37098 -309 37132
rect -275 37098 -262 37132
rect -2842 37059 -262 37098
tri 24138 37090 24144 37096 se
rect 24144 37090 24149 37096
rect -2842 37025 -2829 37059
rect -2795 37025 -2757 37059
rect -2723 37025 -2685 37059
rect -2651 37025 -2613 37059
rect -2579 37025 -2541 37059
rect -2507 37025 -2469 37059
rect -2435 37025 -2397 37059
rect -2363 37025 -2325 37059
rect -2291 37025 -2253 37059
rect -2219 37025 -2181 37059
rect -2147 37025 -2109 37059
rect -2075 37025 -2037 37059
rect -2003 37025 -1965 37059
rect -1931 37025 -1893 37059
rect -1859 37025 -1821 37059
rect -1787 37025 -1749 37059
rect -1715 37025 -1677 37059
rect -1643 37025 -1605 37059
rect -1571 37025 -1533 37059
rect -1499 37025 -1461 37059
rect -1427 37025 -1389 37059
rect -1355 37025 -1317 37059
rect -1283 37025 -1245 37059
rect -1211 37025 -1173 37059
rect -1139 37025 -1101 37059
rect -1067 37025 -1029 37059
rect -995 37025 -957 37059
rect -923 37025 -885 37059
rect -851 37025 -813 37059
rect -779 37025 -741 37059
rect -707 37025 -669 37059
rect -635 37025 -597 37059
rect -563 37025 -525 37059
rect -491 37025 -453 37059
rect -419 37025 -381 37059
rect -347 37025 -309 37059
rect -275 37025 -262 37059
rect -2842 36986 -262 37025
rect -2842 36952 -2829 36986
rect -2795 36952 -2757 36986
rect -2723 36952 -2685 36986
rect -2651 36952 -2613 36986
rect -2579 36952 -2541 36986
rect -2507 36952 -2469 36986
rect -2435 36952 -2397 36986
rect -2363 36952 -2325 36986
rect -2291 36952 -2253 36986
rect -2219 36952 -2181 36986
rect -2147 36952 -2109 36986
rect -2075 36952 -2037 36986
rect -2003 36952 -1965 36986
rect -1931 36952 -1893 36986
rect -1859 36952 -1821 36986
rect -1787 36952 -1749 36986
rect -1715 36952 -1677 36986
rect -1643 36952 -1605 36986
rect -1571 36952 -1533 36986
rect -1499 36952 -1461 36986
rect -1427 36952 -1389 36986
rect -1355 36952 -1317 36986
rect -1283 36952 -1245 36986
rect -1211 36952 -1173 36986
rect -1139 36952 -1101 36986
rect -1067 36952 -1029 36986
rect -995 36952 -957 36986
rect -923 36952 -885 36986
rect -851 36952 -813 36986
rect -779 36952 -741 36986
rect -707 36952 -669 36986
rect -635 36952 -597 36986
rect -563 36952 -525 36986
rect -491 36952 -453 36986
rect -419 36952 -381 36986
rect -347 36952 -309 36986
rect -275 36952 -262 36986
rect -2842 36913 -262 36952
rect -2842 36879 -2829 36913
rect -2795 36879 -2757 36913
rect -2723 36879 -2685 36913
rect -2651 36879 -2613 36913
rect -2579 36879 -2541 36913
rect -2507 36879 -2469 36913
rect -2435 36879 -2397 36913
rect -2363 36879 -2325 36913
rect -2291 36879 -2253 36913
rect -2219 36879 -2181 36913
rect -2147 36879 -2109 36913
rect -2075 36879 -2037 36913
rect -2003 36879 -1965 36913
rect -1931 36879 -1893 36913
rect -1859 36879 -1821 36913
rect -1787 36879 -1749 36913
rect -1715 36879 -1677 36913
rect -1643 36879 -1605 36913
rect -1571 36879 -1533 36913
rect -1499 36879 -1461 36913
rect -1427 36879 -1389 36913
rect -1355 36879 -1317 36913
rect -1283 36879 -1245 36913
rect -1211 36879 -1173 36913
rect -1139 36879 -1101 36913
rect -1067 36879 -1029 36913
rect -995 36879 -957 36913
rect -923 36879 -885 36913
rect -851 36879 -813 36913
rect -779 36879 -741 36913
rect -707 36879 -669 36913
rect -635 36879 -597 36913
rect -563 36879 -525 36913
rect -491 36879 -453 36913
rect -419 36879 -381 36913
rect -347 36879 -309 36913
rect -275 36879 -262 36913
rect -2842 36840 -262 36879
rect -2842 36806 -2829 36840
rect -2795 36806 -2757 36840
rect -2723 36806 -2685 36840
rect -2651 36806 -2613 36840
rect -2579 36806 -2541 36840
rect -2507 36806 -2469 36840
rect -2435 36806 -2397 36840
rect -2363 36806 -2325 36840
rect -2291 36806 -2253 36840
rect -2219 36806 -2181 36840
rect -2147 36806 -2109 36840
rect -2075 36806 -2037 36840
rect -2003 36806 -1965 36840
rect -1931 36806 -1893 36840
rect -1859 36806 -1821 36840
rect -1787 36806 -1749 36840
rect -1715 36806 -1677 36840
rect -1643 36806 -1605 36840
rect -1571 36806 -1533 36840
rect -1499 36806 -1461 36840
rect -1427 36806 -1389 36840
rect -1355 36806 -1317 36840
rect -1283 36806 -1245 36840
rect -1211 36806 -1173 36840
rect -1139 36806 -1101 36840
rect -1067 36806 -1029 36840
rect -995 36806 -957 36840
rect -923 36806 -885 36840
rect -851 36806 -813 36840
rect -779 36806 -741 36840
rect -707 36806 -669 36840
rect -635 36806 -597 36840
rect -563 36806 -525 36840
rect -491 36806 -453 36840
rect -419 36806 -381 36840
rect -347 36806 -309 36840
rect -275 36806 -262 36840
rect -2842 36767 -262 36806
rect -2842 36733 -2829 36767
rect -2795 36733 -2757 36767
rect -2723 36733 -2685 36767
rect -2651 36733 -2613 36767
rect -2579 36733 -2541 36767
rect -2507 36733 -2469 36767
rect -2435 36733 -2397 36767
rect -2363 36733 -2325 36767
rect -2291 36733 -2253 36767
rect -2219 36733 -2181 36767
rect -2147 36733 -2109 36767
rect -2075 36733 -2037 36767
rect -2003 36733 -1965 36767
rect -1931 36733 -1893 36767
rect -1859 36733 -1821 36767
rect -1787 36733 -1749 36767
rect -1715 36733 -1677 36767
rect -1643 36733 -1605 36767
rect -1571 36733 -1533 36767
rect -1499 36733 -1461 36767
rect -1427 36733 -1389 36767
rect -1355 36733 -1317 36767
rect -1283 36733 -1245 36767
rect -1211 36733 -1173 36767
rect -1139 36733 -1101 36767
rect -1067 36733 -1029 36767
rect -995 36733 -957 36767
rect -923 36733 -885 36767
rect -851 36733 -813 36767
rect -779 36733 -741 36767
rect -707 36733 -669 36767
rect -635 36733 -597 36767
rect -563 36733 -525 36767
rect -491 36733 -453 36767
rect -419 36733 -381 36767
rect -347 36733 -309 36767
rect -275 36733 -262 36767
rect -2842 36694 -262 36733
rect -2842 36660 -2829 36694
rect -2795 36660 -2757 36694
rect -2723 36660 -2685 36694
rect -2651 36660 -2613 36694
rect -2579 36660 -2541 36694
rect -2507 36660 -2469 36694
rect -2435 36660 -2397 36694
rect -2363 36660 -2325 36694
rect -2291 36660 -2253 36694
rect -2219 36660 -2181 36694
rect -2147 36660 -2109 36694
rect -2075 36660 -2037 36694
rect -2003 36660 -1965 36694
rect -1931 36660 -1893 36694
rect -1859 36660 -1821 36694
rect -1787 36660 -1749 36694
rect -1715 36660 -1677 36694
rect -1643 36660 -1605 36694
rect -1571 36660 -1533 36694
rect -1499 36660 -1461 36694
rect -1427 36660 -1389 36694
rect -1355 36660 -1317 36694
rect -1283 36660 -1245 36694
rect -1211 36660 -1173 36694
rect -1139 36660 -1101 36694
rect -1067 36660 -1029 36694
rect -995 36660 -957 36694
rect -923 36660 -885 36694
rect -851 36660 -813 36694
rect -779 36660 -741 36694
rect -707 36660 -669 36694
rect -635 36660 -597 36694
rect -563 36660 -525 36694
rect -491 36660 -453 36694
rect -419 36660 -381 36694
rect -347 36660 -309 36694
rect -275 36660 -262 36694
rect -2842 36621 -262 36660
rect -2842 36587 -2829 36621
rect -2795 36587 -2757 36621
rect -2723 36587 -2685 36621
rect -2651 36587 -2613 36621
rect -2579 36587 -2541 36621
rect -2507 36587 -2469 36621
rect -2435 36587 -2397 36621
rect -2363 36587 -2325 36621
rect -2291 36587 -2253 36621
rect -2219 36587 -2181 36621
rect -2147 36587 -2109 36621
rect -2075 36587 -2037 36621
rect -2003 36587 -1965 36621
rect -1931 36587 -1893 36621
rect -1859 36587 -1821 36621
rect -1787 36587 -1749 36621
rect -1715 36587 -1677 36621
rect -1643 36587 -1605 36621
rect -1571 36587 -1533 36621
rect -1499 36587 -1461 36621
rect -1427 36587 -1389 36621
rect -1355 36587 -1317 36621
rect -1283 36587 -1245 36621
rect -1211 36587 -1173 36621
rect -1139 36587 -1101 36621
rect -1067 36587 -1029 36621
rect -995 36587 -957 36621
rect -923 36587 -885 36621
rect -851 36587 -813 36621
rect -779 36587 -741 36621
rect -707 36587 -669 36621
rect -635 36587 -597 36621
rect -563 36587 -525 36621
rect -491 36587 -453 36621
rect -419 36587 -381 36621
rect -347 36587 -309 36621
rect -275 36587 -262 36621
rect -2842 36548 -262 36587
rect -2842 36514 -2829 36548
rect -2795 36514 -2757 36548
rect -2723 36514 -2685 36548
rect -2651 36514 -2613 36548
rect -2579 36514 -2541 36548
rect -2507 36514 -2469 36548
rect -2435 36514 -2397 36548
rect -2363 36514 -2325 36548
rect -2291 36514 -2253 36548
rect -2219 36514 -2181 36548
rect -2147 36514 -2109 36548
rect -2075 36514 -2037 36548
rect -2003 36514 -1965 36548
rect -1931 36514 -1893 36548
rect -1859 36514 -1821 36548
rect -1787 36514 -1749 36548
rect -1715 36514 -1677 36548
rect -1643 36514 -1605 36548
rect -1571 36514 -1533 36548
rect -1499 36514 -1461 36548
rect -1427 36514 -1389 36548
rect -1355 36514 -1317 36548
rect -1283 36514 -1245 36548
rect -1211 36514 -1173 36548
rect -1139 36514 -1101 36548
rect -1067 36514 -1029 36548
rect -995 36514 -957 36548
rect -923 36514 -885 36548
rect -851 36514 -813 36548
rect -779 36514 -741 36548
rect -707 36514 -669 36548
rect -635 36514 -597 36548
rect -563 36514 -525 36548
rect -491 36514 -453 36548
rect -419 36514 -381 36548
rect -347 36514 -309 36548
rect -275 36514 -262 36548
rect -2842 36475 -262 36514
rect -2842 36441 -2829 36475
rect -2795 36441 -2757 36475
rect -2723 36441 -2685 36475
rect -2651 36441 -2613 36475
rect -2579 36441 -2541 36475
rect -2507 36441 -2469 36475
rect -2435 36441 -2397 36475
rect -2363 36441 -2325 36475
rect -2291 36441 -2253 36475
rect -2219 36441 -2181 36475
rect -2147 36441 -2109 36475
rect -2075 36441 -2037 36475
rect -2003 36441 -1965 36475
rect -1931 36441 -1893 36475
rect -1859 36441 -1821 36475
rect -1787 36441 -1749 36475
rect -1715 36441 -1677 36475
rect -1643 36441 -1605 36475
rect -1571 36441 -1533 36475
rect -1499 36441 -1461 36475
rect -1427 36441 -1389 36475
rect -1355 36441 -1317 36475
rect -1283 36441 -1245 36475
rect -1211 36441 -1173 36475
rect -1139 36441 -1101 36475
rect -1067 36441 -1029 36475
rect -995 36441 -957 36475
rect -923 36441 -885 36475
rect -851 36441 -813 36475
rect -779 36441 -741 36475
rect -707 36441 -669 36475
rect -635 36441 -597 36475
rect -563 36441 -525 36475
rect -491 36441 -453 36475
rect -419 36441 -381 36475
rect -347 36441 -309 36475
rect -275 36441 -262 36475
rect -2842 36402 -262 36441
rect -2842 36368 -2829 36402
rect -2795 36368 -2757 36402
rect -2723 36368 -2685 36402
rect -2651 36368 -2613 36402
rect -2579 36368 -2541 36402
rect -2507 36368 -2469 36402
rect -2435 36368 -2397 36402
rect -2363 36368 -2325 36402
rect -2291 36368 -2253 36402
rect -2219 36368 -2181 36402
rect -2147 36368 -2109 36402
rect -2075 36368 -2037 36402
rect -2003 36368 -1965 36402
rect -1931 36368 -1893 36402
rect -1859 36368 -1821 36402
rect -1787 36368 -1749 36402
rect -1715 36368 -1677 36402
rect -1643 36368 -1605 36402
rect -1571 36368 -1533 36402
rect -1499 36368 -1461 36402
rect -1427 36368 -1389 36402
rect -1355 36368 -1317 36402
rect -1283 36368 -1245 36402
rect -1211 36368 -1173 36402
rect -1139 36368 -1101 36402
rect -1067 36368 -1029 36402
rect -995 36368 -957 36402
rect -923 36368 -885 36402
rect -851 36368 -813 36402
rect -779 36368 -741 36402
rect -707 36368 -669 36402
rect -635 36368 -597 36402
rect -563 36368 -525 36402
rect -491 36368 -453 36402
rect -419 36368 -381 36402
rect -347 36368 -309 36402
rect -275 36368 -262 36402
rect -2842 36329 -262 36368
rect -2842 36295 -2829 36329
rect -2795 36295 -2757 36329
rect -2723 36295 -2685 36329
rect -2651 36295 -2613 36329
rect -2579 36295 -2541 36329
rect -2507 36295 -2469 36329
rect -2435 36295 -2397 36329
rect -2363 36295 -2325 36329
rect -2291 36295 -2253 36329
rect -2219 36295 -2181 36329
rect -2147 36295 -2109 36329
rect -2075 36295 -2037 36329
rect -2003 36295 -1965 36329
rect -1931 36295 -1893 36329
rect -1859 36295 -1821 36329
rect -1787 36295 -1749 36329
rect -1715 36295 -1677 36329
rect -1643 36295 -1605 36329
rect -1571 36295 -1533 36329
rect -1499 36295 -1461 36329
rect -1427 36295 -1389 36329
rect -1355 36295 -1317 36329
rect -1283 36295 -1245 36329
rect -1211 36295 -1173 36329
rect -1139 36295 -1101 36329
rect -1067 36295 -1029 36329
rect -995 36295 -957 36329
rect -923 36295 -885 36329
rect -851 36295 -813 36329
rect -779 36295 -741 36329
rect -707 36295 -669 36329
rect -635 36295 -597 36329
rect -563 36295 -525 36329
rect -491 36295 -453 36329
rect -419 36295 -381 36329
rect -347 36295 -309 36329
rect -275 36295 -262 36329
rect -2842 36256 -262 36295
rect -2842 36222 -2829 36256
rect -2795 36222 -2757 36256
rect -2723 36222 -2685 36256
rect -2651 36222 -2613 36256
rect -2579 36222 -2541 36256
rect -2507 36222 -2469 36256
rect -2435 36222 -2397 36256
rect -2363 36222 -2325 36256
rect -2291 36222 -2253 36256
rect -2219 36222 -2181 36256
rect -2147 36222 -2109 36256
rect -2075 36222 -2037 36256
rect -2003 36222 -1965 36256
rect -1931 36222 -1893 36256
rect -1859 36222 -1821 36256
rect -1787 36222 -1749 36256
rect -1715 36222 -1677 36256
rect -1643 36222 -1605 36256
rect -1571 36222 -1533 36256
rect -1499 36222 -1461 36256
rect -1427 36222 -1389 36256
rect -1355 36222 -1317 36256
rect -1283 36222 -1245 36256
rect -1211 36222 -1173 36256
rect -1139 36222 -1101 36256
rect -1067 36222 -1029 36256
rect -995 36222 -957 36256
rect -923 36222 -885 36256
rect -851 36222 -813 36256
rect -779 36222 -741 36256
rect -707 36222 -669 36256
rect -635 36222 -597 36256
rect -563 36222 -525 36256
rect -491 36222 -453 36256
rect -419 36222 -381 36256
rect -347 36222 -309 36256
rect -275 36222 -262 36256
rect -2842 36183 -262 36222
rect -2842 36149 -2829 36183
rect -2795 36149 -2757 36183
rect -2723 36149 -2685 36183
rect -2651 36149 -2613 36183
rect -2579 36149 -2541 36183
rect -2507 36149 -2469 36183
rect -2435 36149 -2397 36183
rect -2363 36149 -2325 36183
rect -2291 36149 -2253 36183
rect -2219 36149 -2181 36183
rect -2147 36149 -2109 36183
rect -2075 36149 -2037 36183
rect -2003 36149 -1965 36183
rect -1931 36149 -1893 36183
rect -1859 36149 -1821 36183
rect -1787 36149 -1749 36183
rect -1715 36149 -1677 36183
rect -1643 36149 -1605 36183
rect -1571 36149 -1533 36183
rect -1499 36149 -1461 36183
rect -1427 36149 -1389 36183
rect -1355 36149 -1317 36183
rect -1283 36149 -1245 36183
rect -1211 36149 -1173 36183
rect -1139 36149 -1101 36183
rect -1067 36149 -1029 36183
rect -995 36149 -957 36183
rect -923 36149 -885 36183
rect -851 36149 -813 36183
rect -779 36149 -741 36183
rect -707 36149 -669 36183
rect -635 36149 -597 36183
rect -563 36149 -525 36183
rect -491 36149 -453 36183
rect -419 36149 -381 36183
rect -347 36149 -309 36183
rect -275 36149 -262 36183
rect -2842 36110 -262 36149
rect -2842 36076 -2829 36110
rect -2795 36076 -2757 36110
rect -2723 36076 -2685 36110
rect -2651 36076 -2613 36110
rect -2579 36076 -2541 36110
rect -2507 36076 -2469 36110
rect -2435 36076 -2397 36110
rect -2363 36076 -2325 36110
rect -2291 36076 -2253 36110
rect -2219 36076 -2181 36110
rect -2147 36076 -2109 36110
rect -2075 36076 -2037 36110
rect -2003 36076 -1965 36110
rect -1931 36076 -1893 36110
rect -1859 36076 -1821 36110
rect -1787 36076 -1749 36110
rect -1715 36076 -1677 36110
rect -1643 36076 -1605 36110
rect -1571 36076 -1533 36110
rect -1499 36076 -1461 36110
rect -1427 36076 -1389 36110
rect -1355 36076 -1317 36110
rect -1283 36076 -1245 36110
rect -1211 36076 -1173 36110
rect -1139 36076 -1101 36110
rect -1067 36076 -1029 36110
rect -995 36076 -957 36110
rect -923 36076 -885 36110
rect -851 36076 -813 36110
rect -779 36076 -741 36110
rect -707 36076 -669 36110
rect -635 36076 -597 36110
rect -563 36076 -525 36110
rect -491 36076 -453 36110
rect -419 36076 -381 36110
rect -347 36076 -309 36110
rect -275 36076 -262 36110
rect -2842 36037 -262 36076
rect -2842 36003 -2829 36037
rect -2795 36003 -2757 36037
rect -2723 36003 -2685 36037
rect -2651 36003 -2613 36037
rect -2579 36003 -2541 36037
rect -2507 36003 -2469 36037
rect -2435 36003 -2397 36037
rect -2363 36003 -2325 36037
rect -2291 36003 -2253 36037
rect -2219 36003 -2181 36037
rect -2147 36003 -2109 36037
rect -2075 36003 -2037 36037
rect -2003 36003 -1965 36037
rect -1931 36003 -1893 36037
rect -1859 36003 -1821 36037
rect -1787 36003 -1749 36037
rect -1715 36003 -1677 36037
rect -1643 36003 -1605 36037
rect -1571 36003 -1533 36037
rect -1499 36003 -1461 36037
rect -1427 36003 -1389 36037
rect -1355 36003 -1317 36037
rect -1283 36003 -1245 36037
rect -1211 36003 -1173 36037
rect -1139 36003 -1101 36037
rect -1067 36003 -1029 36037
rect -995 36003 -957 36037
rect -923 36003 -885 36037
rect -851 36003 -813 36037
rect -779 36003 -741 36037
rect -707 36003 -669 36037
rect -635 36003 -597 36037
rect -563 36003 -525 36037
rect -491 36003 -453 36037
rect -419 36003 -381 36037
rect -347 36003 -309 36037
rect -275 36003 -262 36037
rect -2842 35964 -262 36003
rect -2842 35930 -2829 35964
rect -2795 35930 -2757 35964
rect -2723 35930 -2685 35964
rect -2651 35930 -2613 35964
rect -2579 35930 -2541 35964
rect -2507 35930 -2469 35964
rect -2435 35930 -2397 35964
rect -2363 35930 -2325 35964
rect -2291 35930 -2253 35964
rect -2219 35930 -2181 35964
rect -2147 35930 -2109 35964
rect -2075 35930 -2037 35964
rect -2003 35930 -1965 35964
rect -1931 35930 -1893 35964
rect -1859 35930 -1821 35964
rect -1787 35930 -1749 35964
rect -1715 35930 -1677 35964
rect -1643 35930 -1605 35964
rect -1571 35930 -1533 35964
rect -1499 35930 -1461 35964
rect -1427 35930 -1389 35964
rect -1355 35930 -1317 35964
rect -1283 35930 -1245 35964
rect -1211 35930 -1173 35964
rect -1139 35930 -1101 35964
rect -1067 35930 -1029 35964
rect -995 35930 -957 35964
rect -923 35930 -885 35964
rect -851 35930 -813 35964
rect -779 35930 -741 35964
rect -707 35930 -669 35964
rect -635 35930 -597 35964
rect -563 35930 -525 35964
rect -491 35930 -453 35964
rect -419 35930 -381 35964
rect -347 35930 -309 35964
rect -275 35930 -262 35964
rect -2842 35891 -262 35930
rect -2842 35857 -2829 35891
rect -2795 35857 -2757 35891
rect -2723 35857 -2685 35891
rect -2651 35857 -2613 35891
rect -2579 35857 -2541 35891
rect -2507 35857 -2469 35891
rect -2435 35857 -2397 35891
rect -2363 35857 -2325 35891
rect -2291 35857 -2253 35891
rect -2219 35857 -2181 35891
rect -2147 35857 -2109 35891
rect -2075 35857 -2037 35891
rect -2003 35857 -1965 35891
rect -1931 35857 -1893 35891
rect -1859 35857 -1821 35891
rect -1787 35857 -1749 35891
rect -1715 35857 -1677 35891
rect -1643 35857 -1605 35891
rect -1571 35857 -1533 35891
rect -1499 35857 -1461 35891
rect -1427 35857 -1389 35891
rect -1355 35857 -1317 35891
rect -1283 35857 -1245 35891
rect -1211 35857 -1173 35891
rect -1139 35857 -1101 35891
rect -1067 35857 -1029 35891
rect -995 35857 -957 35891
rect -923 35857 -885 35891
rect -851 35857 -813 35891
rect -779 35857 -741 35891
rect -707 35857 -669 35891
rect -635 35857 -597 35891
rect -563 35857 -525 35891
rect -491 35857 -453 35891
rect -419 35857 -381 35891
rect -347 35857 -309 35891
rect -275 35857 -262 35891
rect -2842 35818 -262 35857
rect -2842 35784 -2829 35818
rect -2795 35784 -2757 35818
rect -2723 35784 -2685 35818
rect -2651 35784 -2613 35818
rect -2579 35784 -2541 35818
rect -2507 35784 -2469 35818
rect -2435 35784 -2397 35818
rect -2363 35784 -2325 35818
rect -2291 35784 -2253 35818
rect -2219 35784 -2181 35818
rect -2147 35784 -2109 35818
rect -2075 35784 -2037 35818
rect -2003 35784 -1965 35818
rect -1931 35784 -1893 35818
rect -1859 35784 -1821 35818
rect -1787 35784 -1749 35818
rect -1715 35784 -1677 35818
rect -1643 35784 -1605 35818
rect -1571 35784 -1533 35818
rect -1499 35784 -1461 35818
rect -1427 35784 -1389 35818
rect -1355 35784 -1317 35818
rect -1283 35784 -1245 35818
rect -1211 35784 -1173 35818
rect -1139 35784 -1101 35818
rect -1067 35784 -1029 35818
rect -995 35784 -957 35818
rect -923 35784 -885 35818
rect -851 35784 -813 35818
rect -779 35784 -741 35818
rect -707 35784 -669 35818
rect -635 35784 -597 35818
rect -563 35784 -525 35818
rect -491 35784 -453 35818
rect -419 35784 -381 35818
rect -347 35784 -309 35818
rect -275 35784 -262 35818
rect -2842 35745 -262 35784
rect -2842 35711 -2829 35745
rect -2795 35711 -2757 35745
rect -2723 35711 -2685 35745
rect -2651 35711 -2613 35745
rect -2579 35711 -2541 35745
rect -2507 35711 -2469 35745
rect -2435 35711 -2397 35745
rect -2363 35711 -2325 35745
rect -2291 35711 -2253 35745
rect -2219 35711 -2181 35745
rect -2147 35711 -2109 35745
rect -2075 35711 -2037 35745
rect -2003 35711 -1965 35745
rect -1931 35711 -1893 35745
rect -1859 35711 -1821 35745
rect -1787 35711 -1749 35745
rect -1715 35711 -1677 35745
rect -1643 35711 -1605 35745
rect -1571 35711 -1533 35745
rect -1499 35711 -1461 35745
rect -1427 35711 -1389 35745
rect -1355 35711 -1317 35745
rect -1283 35711 -1245 35745
rect -1211 35711 -1173 35745
rect -1139 35711 -1101 35745
rect -1067 35711 -1029 35745
rect -995 35711 -957 35745
rect -923 35711 -885 35745
rect -851 35711 -813 35745
rect -779 35711 -741 35745
rect -707 35711 -669 35745
rect -635 35711 -597 35745
rect -563 35711 -525 35745
rect -491 35711 -453 35745
rect -419 35711 -381 35745
rect -347 35711 -309 35745
rect -275 35711 -262 35745
rect -2842 35672 -262 35711
rect -2842 35638 -2829 35672
rect -2795 35638 -2757 35672
rect -2723 35638 -2685 35672
rect -2651 35638 -2613 35672
rect -2579 35638 -2541 35672
rect -2507 35638 -2469 35672
rect -2435 35638 -2397 35672
rect -2363 35638 -2325 35672
rect -2291 35638 -2253 35672
rect -2219 35638 -2181 35672
rect -2147 35638 -2109 35672
rect -2075 35638 -2037 35672
rect -2003 35638 -1965 35672
rect -1931 35638 -1893 35672
rect -1859 35638 -1821 35672
rect -1787 35638 -1749 35672
rect -1715 35638 -1677 35672
rect -1643 35638 -1605 35672
rect -1571 35638 -1533 35672
rect -1499 35638 -1461 35672
rect -1427 35638 -1389 35672
rect -1355 35638 -1317 35672
rect -1283 35638 -1245 35672
rect -1211 35638 -1173 35672
rect -1139 35638 -1101 35672
rect -1067 35638 -1029 35672
rect -995 35638 -957 35672
rect -923 35638 -885 35672
rect -851 35638 -813 35672
rect -779 35638 -741 35672
rect -707 35638 -669 35672
rect -635 35638 -597 35672
rect -563 35638 -525 35672
rect -491 35638 -453 35672
rect -419 35638 -381 35672
rect -347 35638 -309 35672
rect -275 35638 -262 35672
rect -2842 35599 -262 35638
rect -2842 35565 -2829 35599
rect -2795 35565 -2757 35599
rect -2723 35565 -2685 35599
rect -2651 35565 -2613 35599
rect -2579 35565 -2541 35599
rect -2507 35565 -2469 35599
rect -2435 35565 -2397 35599
rect -2363 35565 -2325 35599
rect -2291 35565 -2253 35599
rect -2219 35565 -2181 35599
rect -2147 35565 -2109 35599
rect -2075 35565 -2037 35599
rect -2003 35565 -1965 35599
rect -1931 35565 -1893 35599
rect -1859 35565 -1821 35599
rect -1787 35565 -1749 35599
rect -1715 35565 -1677 35599
rect -1643 35565 -1605 35599
rect -1571 35565 -1533 35599
rect -1499 35565 -1461 35599
rect -1427 35565 -1389 35599
rect -1355 35565 -1317 35599
rect -1283 35565 -1245 35599
rect -1211 35565 -1173 35599
rect -1139 35565 -1101 35599
rect -1067 35565 -1029 35599
rect -995 35565 -957 35599
rect -923 35565 -885 35599
rect -851 35565 -813 35599
rect -779 35565 -741 35599
rect -707 35565 -669 35599
rect -635 35565 -597 35599
rect -563 35565 -525 35599
rect -491 35565 -453 35599
rect -419 35565 -381 35599
rect -347 35565 -309 35599
rect -275 35565 -262 35599
rect -2842 35526 -262 35565
rect -2842 35492 -2829 35526
rect -2795 35492 -2757 35526
rect -2723 35492 -2685 35526
rect -2651 35492 -2613 35526
rect -2579 35492 -2541 35526
rect -2507 35492 -2469 35526
rect -2435 35492 -2397 35526
rect -2363 35492 -2325 35526
rect -2291 35492 -2253 35526
rect -2219 35492 -2181 35526
rect -2147 35492 -2109 35526
rect -2075 35492 -2037 35526
rect -2003 35492 -1965 35526
rect -1931 35492 -1893 35526
rect -1859 35492 -1821 35526
rect -1787 35492 -1749 35526
rect -1715 35492 -1677 35526
rect -1643 35492 -1605 35526
rect -1571 35492 -1533 35526
rect -1499 35492 -1461 35526
rect -1427 35492 -1389 35526
rect -1355 35492 -1317 35526
rect -1283 35492 -1245 35526
rect -1211 35492 -1173 35526
rect -1139 35492 -1101 35526
rect -1067 35492 -1029 35526
rect -995 35492 -957 35526
rect -923 35492 -885 35526
rect -851 35492 -813 35526
rect -779 35492 -741 35526
rect -707 35492 -669 35526
rect -635 35492 -597 35526
rect -563 35492 -525 35526
rect -491 35492 -453 35526
rect -419 35492 -381 35526
rect -347 35492 -309 35526
rect -275 35492 -262 35526
rect -2842 35453 -262 35492
rect -2842 35419 -2829 35453
rect -2795 35419 -2757 35453
rect -2723 35419 -2685 35453
rect -2651 35419 -2613 35453
rect -2579 35419 -2541 35453
rect -2507 35419 -2469 35453
rect -2435 35419 -2397 35453
rect -2363 35419 -2325 35453
rect -2291 35419 -2253 35453
rect -2219 35419 -2181 35453
rect -2147 35419 -2109 35453
rect -2075 35419 -2037 35453
rect -2003 35419 -1965 35453
rect -1931 35419 -1893 35453
rect -1859 35419 -1821 35453
rect -1787 35419 -1749 35453
rect -1715 35419 -1677 35453
rect -1643 35419 -1605 35453
rect -1571 35419 -1533 35453
rect -1499 35419 -1461 35453
rect -1427 35419 -1389 35453
rect -1355 35419 -1317 35453
rect -1283 35419 -1245 35453
rect -1211 35419 -1173 35453
rect -1139 35419 -1101 35453
rect -1067 35419 -1029 35453
rect -995 35419 -957 35453
rect -923 35419 -885 35453
rect -851 35419 -813 35453
rect -779 35419 -741 35453
rect -707 35419 -669 35453
rect -635 35419 -597 35453
rect -563 35419 -525 35453
rect -491 35419 -453 35453
rect -419 35419 -381 35453
rect -347 35419 -309 35453
rect -275 35419 -262 35453
rect -2842 35380 -262 35419
rect -2842 35346 -2829 35380
rect -2795 35346 -2757 35380
rect -2723 35346 -2685 35380
rect -2651 35346 -2613 35380
rect -2579 35346 -2541 35380
rect -2507 35346 -2469 35380
rect -2435 35346 -2397 35380
rect -2363 35346 -2325 35380
rect -2291 35346 -2253 35380
rect -2219 35346 -2181 35380
rect -2147 35346 -2109 35380
rect -2075 35346 -2037 35380
rect -2003 35346 -1965 35380
rect -1931 35346 -1893 35380
rect -1859 35346 -1821 35380
rect -1787 35346 -1749 35380
rect -1715 35346 -1677 35380
rect -1643 35346 -1605 35380
rect -1571 35346 -1533 35380
rect -1499 35346 -1461 35380
rect -1427 35346 -1389 35380
rect -1355 35346 -1317 35380
rect -1283 35346 -1245 35380
rect -1211 35346 -1173 35380
rect -1139 35346 -1101 35380
rect -1067 35346 -1029 35380
rect -995 35346 -957 35380
rect -923 35346 -885 35380
rect -851 35346 -813 35380
rect -779 35346 -741 35380
rect -707 35346 -669 35380
rect -635 35346 -597 35380
rect -563 35346 -525 35380
rect -491 35346 -453 35380
rect -419 35346 -381 35380
rect -347 35346 -309 35380
rect -275 35346 -262 35380
rect -2842 35307 -262 35346
rect -2842 35273 -2829 35307
rect -2795 35273 -2757 35307
rect -2723 35273 -2685 35307
rect -2651 35273 -2613 35307
rect -2579 35273 -2541 35307
rect -2507 35273 -2469 35307
rect -2435 35273 -2397 35307
rect -2363 35273 -2325 35307
rect -2291 35273 -2253 35307
rect -2219 35273 -2181 35307
rect -2147 35273 -2109 35307
rect -2075 35273 -2037 35307
rect -2003 35273 -1965 35307
rect -1931 35273 -1893 35307
rect -1859 35273 -1821 35307
rect -1787 35273 -1749 35307
rect -1715 35273 -1677 35307
rect -1643 35273 -1605 35307
rect -1571 35273 -1533 35307
rect -1499 35273 -1461 35307
rect -1427 35273 -1389 35307
rect -1355 35273 -1317 35307
rect -1283 35273 -1245 35307
rect -1211 35273 -1173 35307
rect -1139 35273 -1101 35307
rect -1067 35273 -1029 35307
rect -995 35273 -957 35307
rect -923 35273 -885 35307
rect -851 35273 -813 35307
rect -779 35273 -741 35307
rect -707 35273 -669 35307
rect -635 35273 -597 35307
rect -563 35273 -525 35307
rect -491 35273 -453 35307
rect -419 35273 -381 35307
rect -347 35273 -309 35307
rect -275 35273 -262 35307
rect -2842 35234 -262 35273
rect -2842 35200 -2829 35234
rect -2795 35200 -2757 35234
rect -2723 35200 -2685 35234
rect -2651 35200 -2613 35234
rect -2579 35200 -2541 35234
rect -2507 35200 -2469 35234
rect -2435 35200 -2397 35234
rect -2363 35200 -2325 35234
rect -2291 35200 -2253 35234
rect -2219 35200 -2181 35234
rect -2147 35200 -2109 35234
rect -2075 35200 -2037 35234
rect -2003 35200 -1965 35234
rect -1931 35200 -1893 35234
rect -1859 35200 -1821 35234
rect -1787 35200 -1749 35234
rect -1715 35200 -1677 35234
rect -1643 35200 -1605 35234
rect -1571 35200 -1533 35234
rect -1499 35200 -1461 35234
rect -1427 35200 -1389 35234
rect -1355 35200 -1317 35234
rect -1283 35200 -1245 35234
rect -1211 35200 -1173 35234
rect -1139 35200 -1101 35234
rect -1067 35200 -1029 35234
rect -995 35200 -957 35234
rect -923 35200 -885 35234
rect -851 35200 -813 35234
rect -779 35200 -741 35234
rect -707 35200 -669 35234
rect -635 35200 -597 35234
rect -563 35200 -525 35234
rect -491 35200 -453 35234
rect -419 35200 -381 35234
rect -347 35200 -309 35234
rect -275 35200 -262 35234
rect -2842 35161 -262 35200
rect -2842 35127 -2829 35161
rect -2795 35127 -2757 35161
rect -2723 35127 -2685 35161
rect -2651 35127 -2613 35161
rect -2579 35127 -2541 35161
rect -2507 35127 -2469 35161
rect -2435 35127 -2397 35161
rect -2363 35127 -2325 35161
rect -2291 35127 -2253 35161
rect -2219 35127 -2181 35161
rect -2147 35127 -2109 35161
rect -2075 35127 -2037 35161
rect -2003 35127 -1965 35161
rect -1931 35127 -1893 35161
rect -1859 35127 -1821 35161
rect -1787 35127 -1749 35161
rect -1715 35127 -1677 35161
rect -1643 35127 -1605 35161
rect -1571 35127 -1533 35161
rect -1499 35127 -1461 35161
rect -1427 35127 -1389 35161
rect -1355 35127 -1317 35161
rect -1283 35127 -1245 35161
rect -1211 35127 -1173 35161
rect -1139 35127 -1101 35161
rect -1067 35127 -1029 35161
rect -995 35127 -957 35161
rect -923 35127 -885 35161
rect -851 35127 -813 35161
rect -779 35127 -741 35161
rect -707 35127 -669 35161
rect -635 35127 -597 35161
rect -563 35127 -525 35161
rect -491 35127 -453 35161
rect -419 35127 -381 35161
rect -347 35127 -309 35161
rect -275 35127 -262 35161
rect -2842 35115 -262 35127
tri 24138 34614 24144 34620 se
rect 24144 34614 24149 34620
tri 24138 30832 24144 30838 ne
rect 24144 30832 24149 30838
rect -1190 25161 -590 25167
rect -1190 25109 -1188 25161
rect -1136 25109 -1120 25161
rect -1068 25109 -1052 25161
rect -1000 25109 -984 25161
rect -932 25109 -916 25161
rect -864 25109 -848 25161
rect -796 25109 -780 25161
rect -728 25109 -712 25161
rect -660 25109 -644 25161
rect -592 25109 -590 25161
rect -1190 25097 -590 25109
rect -1190 25045 -1188 25097
rect -1136 25045 -1120 25097
rect -1068 25045 -1052 25097
rect -1000 25045 -984 25097
rect -932 25045 -916 25097
rect -864 25045 -848 25097
rect -796 25045 -780 25097
rect -728 25045 -712 25097
rect -660 25045 -644 25097
rect -592 25045 -590 25097
rect -1190 25033 -590 25045
rect -1190 24981 -1188 25033
rect -1136 24981 -1120 25033
rect -1068 24981 -1052 25033
rect -1000 24981 -984 25033
rect -932 24981 -916 25033
rect -864 24981 -848 25033
rect -796 24981 -780 25033
rect -728 24981 -712 25033
rect -660 24981 -644 25033
rect -592 24981 -590 25033
rect -1190 24969 -590 24981
rect -1190 24917 -1188 24969
rect -1136 24917 -1120 24969
rect -1068 24917 -1052 24969
rect -1000 24917 -984 24969
rect -932 24917 -916 24969
rect -864 24917 -848 24969
rect -796 24917 -780 24969
rect -728 24917 -712 24969
rect -660 24917 -644 24969
rect -592 24917 -590 24969
rect -1190 24905 -590 24917
rect -1190 24853 -1188 24905
rect -1136 24853 -1120 24905
rect -1068 24853 -1052 24905
rect -1000 24853 -984 24905
rect -932 24853 -916 24905
rect -864 24853 -848 24905
rect -796 24853 -780 24905
rect -728 24853 -712 24905
rect -660 24853 -644 24905
rect -592 24853 -590 24905
rect -1190 24841 -590 24853
rect -1190 24789 -1188 24841
rect -1136 24789 -1120 24841
rect -1068 24789 -1052 24841
rect -1000 24789 -984 24841
rect -932 24789 -916 24841
rect -864 24789 -848 24841
rect -796 24789 -780 24841
rect -728 24789 -712 24841
rect -660 24789 -644 24841
rect -592 24789 -590 24841
rect -1190 24777 -590 24789
rect -1190 24725 -1188 24777
rect -1136 24725 -1120 24777
rect -1068 24725 -1052 24777
rect -1000 24725 -984 24777
rect -932 24725 -916 24777
rect -864 24725 -848 24777
rect -796 24725 -780 24777
rect -728 24725 -712 24777
rect -660 24725 -644 24777
rect -592 24725 -590 24777
rect -1190 24713 -590 24725
rect -1190 24661 -1188 24713
rect -1136 24661 -1120 24713
rect -1068 24661 -1052 24713
rect -1000 24661 -984 24713
rect -932 24661 -916 24713
rect -864 24661 -848 24713
rect -796 24661 -780 24713
rect -728 24661 -712 24713
rect -660 24661 -644 24713
rect -592 24661 -590 24713
rect -1190 24649 -590 24661
rect -1190 24597 -1188 24649
rect -1136 24597 -1120 24649
rect -1068 24597 -1052 24649
rect -1000 24597 -984 24649
rect -932 24597 -916 24649
rect -864 24597 -848 24649
rect -796 24597 -780 24649
rect -728 24597 -712 24649
rect -660 24597 -644 24649
rect -592 24597 -590 24649
rect -1190 24585 -590 24597
rect -1190 24533 -1188 24585
rect -1136 24533 -1120 24585
rect -1068 24533 -1052 24585
rect -1000 24533 -984 24585
rect -932 24533 -916 24585
rect -864 24533 -848 24585
rect -796 24533 -780 24585
rect -728 24533 -712 24585
rect -660 24533 -644 24585
rect -592 24533 -590 24585
rect -1190 24521 -590 24533
rect -1190 24469 -1188 24521
rect -1136 24469 -1120 24521
rect -1068 24469 -1052 24521
rect -1000 24469 -984 24521
rect -932 24469 -916 24521
rect -864 24469 -848 24521
rect -796 24469 -780 24521
rect -728 24469 -712 24521
rect -660 24469 -644 24521
rect -592 24469 -590 24521
rect -1190 24457 -590 24469
rect -1190 24405 -1188 24457
rect -1136 24405 -1120 24457
rect -1068 24405 -1052 24457
rect -1000 24405 -984 24457
rect -932 24405 -916 24457
rect -864 24405 -848 24457
rect -796 24405 -780 24457
rect -728 24405 -712 24457
rect -660 24405 -644 24457
rect -592 24405 -590 24457
rect -1190 24393 -590 24405
rect -1190 24341 -1188 24393
rect -1136 24341 -1120 24393
rect -1068 24341 -1052 24393
rect -1000 24341 -984 24393
rect -932 24341 -916 24393
rect -864 24341 -848 24393
rect -796 24341 -780 24393
rect -728 24341 -712 24393
rect -660 24341 -644 24393
rect -592 24341 -590 24393
rect -1190 24329 -590 24341
rect -1190 24277 -1188 24329
rect -1136 24277 -1120 24329
rect -1068 24277 -1052 24329
rect -1000 24277 -984 24329
rect -932 24277 -916 24329
rect -864 24277 -848 24329
rect -796 24277 -780 24329
rect -728 24277 -712 24329
rect -660 24277 -644 24329
rect -592 24277 -590 24329
rect -1190 24265 -590 24277
rect -1190 24213 -1188 24265
rect -1136 24213 -1120 24265
rect -1068 24213 -1052 24265
rect -1000 24213 -984 24265
rect -932 24213 -916 24265
rect -864 24213 -848 24265
rect -796 24213 -780 24265
rect -728 24213 -712 24265
rect -660 24213 -644 24265
rect -592 24213 -590 24265
rect -1190 24201 -590 24213
rect -1190 24149 -1188 24201
rect -1136 24149 -1120 24201
rect -1068 24149 -1052 24201
rect -1000 24149 -984 24201
rect -932 24149 -916 24201
rect -864 24149 -848 24201
rect -796 24149 -780 24201
rect -728 24149 -712 24201
rect -660 24149 -644 24201
rect -592 24149 -590 24201
rect -1190 24137 -590 24149
rect -1190 24085 -1188 24137
rect -1136 24085 -1120 24137
rect -1068 24085 -1052 24137
rect -1000 24085 -984 24137
rect -932 24085 -916 24137
rect -864 24085 -848 24137
rect -796 24085 -780 24137
rect -728 24085 -712 24137
rect -660 24085 -644 24137
rect -592 24085 -590 24137
rect -1190 24073 -590 24085
rect -1190 24021 -1188 24073
rect -1136 24021 -1120 24073
rect -1068 24021 -1052 24073
rect -1000 24021 -984 24073
rect -932 24021 -916 24073
rect -864 24021 -848 24073
rect -796 24021 -780 24073
rect -728 24021 -712 24073
rect -660 24021 -644 24073
rect -592 24021 -590 24073
rect -1190 24009 -590 24021
rect -1190 23957 -1188 24009
rect -1136 23957 -1120 24009
rect -1068 23957 -1052 24009
rect -1000 23957 -984 24009
rect -932 23957 -916 24009
rect -864 23957 -848 24009
rect -796 23957 -780 24009
rect -728 23957 -712 24009
rect -660 23957 -644 24009
rect -592 23957 -590 24009
rect -1190 23945 -590 23957
rect -1190 23893 -1188 23945
rect -1136 23893 -1120 23945
rect -1068 23893 -1052 23945
rect -1000 23893 -984 23945
rect -932 23893 -916 23945
rect -864 23893 -848 23945
rect -796 23893 -780 23945
rect -728 23893 -712 23945
rect -660 23893 -644 23945
rect -592 23893 -590 23945
rect -1190 23880 -590 23893
rect -1190 23828 -1188 23880
rect -1136 23828 -1120 23880
rect -1068 23828 -1052 23880
rect -1000 23828 -984 23880
rect -932 23828 -916 23880
rect -864 23828 -848 23880
rect -796 23828 -780 23880
rect -728 23828 -712 23880
rect -660 23828 -644 23880
rect -592 23828 -590 23880
rect -1190 23815 -590 23828
rect -1190 23763 -1188 23815
rect -1136 23763 -1120 23815
rect -1068 23763 -1052 23815
rect -1000 23763 -984 23815
rect -932 23763 -916 23815
rect -864 23763 -848 23815
rect -796 23763 -780 23815
rect -728 23763 -712 23815
rect -660 23763 -644 23815
rect -592 23763 -590 23815
rect -1190 23750 -590 23763
rect -1190 23698 -1188 23750
rect -1136 23698 -1120 23750
rect -1068 23698 -1052 23750
rect -1000 23698 -984 23750
rect -932 23698 -916 23750
rect -864 23698 -848 23750
rect -796 23698 -780 23750
rect -728 23698 -712 23750
rect -660 23698 -644 23750
rect -592 23698 -590 23750
rect -1190 23685 -590 23698
rect -1190 23633 -1188 23685
rect -1136 23633 -1120 23685
rect -1068 23633 -1052 23685
rect -1000 23633 -984 23685
rect -932 23633 -916 23685
rect -864 23633 -848 23685
rect -796 23633 -780 23685
rect -728 23633 -712 23685
rect -660 23633 -644 23685
rect -592 23633 -590 23685
rect -1190 23620 -590 23633
rect -1190 23568 -1188 23620
rect -1136 23568 -1120 23620
rect -1068 23568 -1052 23620
rect -1000 23568 -984 23620
rect -932 23568 -916 23620
rect -864 23568 -848 23620
rect -796 23568 -780 23620
rect -728 23568 -712 23620
rect -660 23568 -644 23620
rect -592 23568 -590 23620
rect -1190 23555 -590 23568
rect -1190 23503 -1188 23555
rect -1136 23503 -1120 23555
rect -1068 23503 -1052 23555
rect -1000 23503 -984 23555
rect -932 23503 -916 23555
rect -864 23503 -848 23555
rect -796 23503 -780 23555
rect -728 23503 -712 23555
rect -660 23503 -644 23555
rect -592 23503 -590 23555
rect -1190 23490 -590 23503
rect -1190 23438 -1188 23490
rect -1136 23438 -1120 23490
rect -1068 23438 -1052 23490
rect -1000 23438 -984 23490
rect -932 23438 -916 23490
rect -864 23438 -848 23490
rect -796 23438 -780 23490
rect -728 23438 -712 23490
rect -660 23438 -644 23490
rect -592 23438 -590 23490
rect -1190 23425 -590 23438
rect -1190 23373 -1188 23425
rect -1136 23373 -1120 23425
rect -1068 23373 -1052 23425
rect -1000 23373 -984 23425
rect -932 23373 -916 23425
rect -864 23373 -848 23425
rect -796 23373 -780 23425
rect -728 23373 -712 23425
rect -660 23373 -644 23425
rect -592 23373 -590 23425
rect -1190 23360 -590 23373
rect -1190 23308 -1188 23360
rect -1136 23308 -1120 23360
rect -1068 23308 -1052 23360
rect -1000 23308 -984 23360
rect -932 23308 -916 23360
rect -864 23308 -848 23360
rect -796 23308 -780 23360
rect -728 23308 -712 23360
rect -660 23308 -644 23360
rect -592 23308 -590 23360
rect -1190 23295 -590 23308
rect -1190 23243 -1188 23295
rect -1136 23243 -1120 23295
rect -1068 23243 -1052 23295
rect -1000 23243 -984 23295
rect -932 23243 -916 23295
rect -864 23243 -848 23295
rect -796 23243 -780 23295
rect -728 23243 -712 23295
rect -660 23243 -644 23295
rect -592 23243 -590 23295
rect -1190 23230 -590 23243
rect -1190 23178 -1188 23230
rect -1136 23178 -1120 23230
rect -1068 23178 -1052 23230
rect -1000 23178 -984 23230
rect -932 23178 -916 23230
rect -864 23178 -848 23230
rect -796 23178 -780 23230
rect -728 23178 -712 23230
rect -660 23178 -644 23230
rect -592 23178 -590 23230
rect -1190 23165 -590 23178
rect -1190 23113 -1188 23165
rect -1136 23113 -1120 23165
rect -1068 23113 -1052 23165
rect -1000 23113 -984 23165
rect -932 23113 -916 23165
rect -864 23113 -848 23165
rect -796 23113 -780 23165
rect -728 23113 -712 23165
rect -660 23113 -644 23165
rect -592 23113 -590 23165
rect -1190 23100 -590 23113
rect -1190 23048 -1188 23100
rect -1136 23048 -1120 23100
rect -1068 23048 -1052 23100
rect -1000 23048 -984 23100
rect -932 23048 -916 23100
rect -864 23048 -848 23100
rect -796 23048 -780 23100
rect -728 23048 -712 23100
rect -660 23048 -644 23100
rect -592 23048 -590 23100
rect -1190 23035 -590 23048
rect -1190 22983 -1188 23035
rect -1136 22983 -1120 23035
rect -1068 22983 -1052 23035
rect -1000 22983 -984 23035
rect -932 22983 -916 23035
rect -864 22983 -848 23035
rect -796 22983 -780 23035
rect -728 22983 -712 23035
rect -660 22983 -644 23035
rect -592 22983 -590 23035
rect -1190 22970 -590 22983
rect -1190 22918 -1188 22970
rect -1136 22918 -1120 22970
rect -1068 22918 -1052 22970
rect -1000 22918 -984 22970
rect -932 22918 -916 22970
rect -864 22918 -848 22970
rect -796 22918 -780 22970
rect -728 22918 -712 22970
rect -660 22918 -644 22970
rect -592 22918 -590 22970
rect -1190 22905 -590 22918
rect -1190 22853 -1188 22905
rect -1136 22853 -1120 22905
rect -1068 22853 -1052 22905
rect -1000 22853 -984 22905
rect -932 22853 -916 22905
rect -864 22853 -848 22905
rect -796 22853 -780 22905
rect -728 22853 -712 22905
rect -660 22853 -644 22905
rect -592 22853 -590 22905
rect -1190 22840 -590 22853
rect -1190 22788 -1188 22840
rect -1136 22788 -1120 22840
rect -1068 22788 -1052 22840
rect -1000 22788 -984 22840
rect -932 22788 -916 22840
rect -864 22788 -848 22840
rect -796 22788 -780 22840
rect -728 22788 -712 22840
rect -660 22788 -644 22840
rect -592 22788 -590 22840
rect -1190 22782 -590 22788
tri 10553 15882 10567 15896 ne
rect 10567 15882 11814 15896
tri 11814 15882 11828 15896 nw
tri 10567 15870 10579 15882 ne
rect 10579 15870 11677 15882
tri 10579 15836 10613 15870 ne
rect 10613 15836 10732 15870
rect 10766 15836 10989 15870
rect 11023 15836 11341 15870
rect 11375 15836 11637 15870
rect 11671 15836 11677 15870
tri 10613 15773 10676 15836 ne
rect 10676 15773 11677 15836
tri 10676 15739 10710 15773 ne
rect 10710 15739 10732 15773
rect 10766 15751 11677 15773
rect 10766 15739 10989 15751
tri 10710 15727 10722 15739 ne
rect 10722 15727 10989 15739
tri 10722 15717 10732 15727 ne
rect 10732 15717 10989 15727
rect 11023 15717 11341 15751
rect 11375 15717 11637 15751
rect 11671 15717 11677 15751
tri 11677 15745 11814 15882 nw
tri 10732 15705 10744 15717 ne
rect 10744 15705 11677 15717
tri 10732 15177 10744 15189 se
rect 10744 15177 11763 15189
tri 10722 15167 10732 15177 se
rect 10732 15167 10989 15177
tri 10710 15155 10722 15167 se
rect 10722 15155 10989 15167
tri 10676 15121 10710 15155 se
rect 10710 15121 10732 15155
rect 10766 15143 10989 15155
rect 11023 15143 11341 15177
rect 11375 15143 11637 15177
rect 11671 15143 11723 15177
rect 11757 15167 11763 15177
tri 11763 15167 11784 15188 sw
rect 11757 15143 11784 15167
rect 10766 15121 11784 15143
tri 10613 15058 10676 15121 se
rect 10676 15058 11784 15121
tri 10579 15024 10613 15058 se
rect 10613 15024 10732 15058
rect 10766 15024 10989 15058
rect 11023 15024 11341 15058
rect 11375 15024 11637 15058
rect 11671 15024 11723 15058
rect 11757 15024 11784 15058
tri 10567 15012 10579 15024 se
rect 10579 15012 11784 15024
tri 11784 15012 11939 15167 sw
tri 10553 14998 10567 15012 se
rect 10567 14998 11939 15012
tri 11939 14998 11953 15012 sw
rect 18347 14398 23139 14407
rect 18347 14364 18359 14398
rect 18393 14364 18432 14398
rect 18466 14364 18505 14398
rect 18539 14364 18578 14398
rect 18612 14364 18651 14398
rect 18685 14364 18724 14398
rect 18758 14364 18797 14398
rect 18831 14364 18870 14398
rect 18904 14364 18943 14398
rect 18977 14364 19016 14398
rect 19050 14364 19089 14398
rect 19123 14364 19162 14398
rect 19196 14364 19235 14398
rect 19269 14364 19308 14398
rect 19342 14364 19381 14398
rect 19415 14364 19454 14398
rect 19488 14364 19527 14398
rect 19561 14364 19600 14398
rect 19634 14364 19673 14398
rect 19707 14364 19746 14398
rect 19780 14364 19819 14398
rect 19853 14364 19892 14398
rect 19926 14364 19965 14398
rect 19999 14364 20038 14398
rect 20072 14364 20111 14398
rect 20145 14364 20184 14398
rect 20218 14364 20257 14398
rect 20291 14364 20330 14398
rect 20364 14364 20403 14398
rect 20437 14364 20476 14398
rect 20510 14364 20549 14398
rect 20583 14364 20622 14398
rect 20656 14364 20695 14398
rect 20729 14364 20768 14398
rect 20802 14364 20841 14398
rect 20875 14364 20914 14398
rect 20948 14364 20987 14398
rect 21021 14364 21060 14398
rect 21094 14364 21133 14398
rect 21167 14364 21206 14398
rect 21240 14364 21279 14398
rect 21313 14364 21352 14398
rect 21386 14364 21425 14398
rect 21459 14364 21498 14398
rect 21532 14364 21571 14398
rect 21605 14364 21644 14398
rect 21678 14364 21717 14398
rect 21751 14364 21790 14398
rect 21824 14364 21863 14398
rect 21897 14364 21936 14398
rect 21970 14364 22009 14398
rect 22043 14364 22082 14398
rect 22116 14364 22155 14398
rect 22189 14364 22228 14398
rect 22262 14364 22301 14398
rect 22335 14364 22373 14398
rect 22407 14364 22445 14398
rect 22479 14364 22517 14398
rect 22551 14364 22589 14398
rect 22623 14364 22661 14398
rect 22695 14364 22733 14398
rect 22767 14364 22805 14398
rect 22839 14364 22877 14398
rect 22911 14364 22949 14398
rect 22983 14364 23021 14398
rect 23055 14364 23093 14398
rect 23127 14364 23139 14398
rect 18347 14355 23139 14364
rect 23343 14398 29671 14407
rect 23343 14364 23355 14398
rect 23389 14364 23428 14398
rect 23462 14364 23501 14398
rect 23535 14364 23574 14398
rect 23608 14364 23647 14398
rect 23681 14364 23720 14398
rect 23754 14364 23793 14398
rect 23827 14364 23865 14398
rect 23899 14364 23937 14398
rect 23971 14364 24009 14398
rect 24043 14364 24081 14398
rect 24115 14364 24153 14398
rect 24187 14364 24225 14398
rect 24259 14364 24297 14398
rect 24331 14364 24369 14398
rect 24403 14364 24441 14398
rect 24475 14364 24513 14398
rect 24547 14364 24585 14398
rect 24619 14364 24657 14398
rect 24691 14364 24729 14398
rect 24763 14364 24801 14398
rect 24835 14364 24873 14398
rect 24907 14364 24945 14398
rect 24979 14364 25017 14398
rect 25051 14364 25089 14398
rect 25123 14364 25161 14398
rect 25195 14364 25233 14398
rect 25267 14364 25305 14398
rect 25339 14364 25377 14398
rect 25411 14364 25449 14398
rect 25483 14364 25521 14398
rect 25555 14364 25593 14398
rect 25627 14364 25665 14398
rect 25699 14364 25737 14398
rect 25771 14364 25809 14398
rect 25843 14364 25881 14398
rect 25915 14364 25953 14398
rect 25987 14364 26025 14398
rect 26059 14364 26097 14398
rect 26131 14364 26169 14398
rect 26203 14364 26241 14398
rect 26275 14364 26313 14398
rect 26347 14364 26385 14398
rect 26419 14364 26457 14398
rect 26491 14364 26529 14398
rect 26563 14364 26601 14398
rect 26635 14364 26673 14398
rect 26707 14364 26745 14398
rect 26779 14364 26817 14398
rect 26851 14364 26889 14398
rect 26923 14364 26961 14398
rect 26995 14364 27033 14398
rect 27067 14364 27105 14398
rect 27139 14364 27177 14398
rect 27211 14364 27249 14398
rect 27283 14364 27321 14398
rect 27355 14364 27393 14398
rect 27427 14364 27465 14398
rect 27499 14364 27537 14398
rect 27571 14364 27609 14398
rect 27643 14364 27681 14398
rect 27715 14364 27753 14398
rect 27787 14364 27825 14398
rect 27859 14364 27897 14398
rect 27931 14364 27969 14398
rect 28003 14364 28041 14398
rect 28075 14364 28113 14398
rect 28147 14364 28185 14398
rect 28219 14364 28257 14398
rect 28291 14364 28329 14398
rect 28363 14364 28401 14398
rect 28435 14364 28473 14398
rect 28507 14364 28545 14398
rect 28579 14364 28617 14398
rect 28651 14364 28689 14398
rect 28723 14364 28761 14398
rect 28795 14364 28833 14398
rect 28867 14364 28905 14398
rect 28939 14364 28977 14398
rect 29011 14364 29049 14398
rect 29083 14364 29121 14398
rect 29155 14364 29193 14398
rect 29227 14364 29265 14398
rect 29299 14364 29337 14398
rect 29371 14364 29409 14398
rect 29443 14364 29481 14398
rect 29515 14364 29553 14398
rect 29587 14364 29625 14398
rect 29659 14364 29671 14398
rect 23343 14355 29671 14364
rect 5493 14285 7306 14331
tri 5493 14272 5506 14285 ne
rect 5506 14272 7306 14285
rect 38 14271 1222 14272
tri 1222 14271 1223 14272 nw
tri 5506 14271 5507 14272 ne
rect 5507 14271 7194 14272
rect 38 14257 1208 14271
tri 1208 14257 1222 14271 nw
tri 5507 14257 5521 14271 ne
rect 5521 14257 5800 14271
rect 38 14254 1205 14257
tri 1205 14254 1208 14257 nw
tri 5521 14254 5524 14257 ne
rect 5524 14254 5800 14257
tri 5800 14254 5817 14271 nw
tri 6017 14254 6034 14271 ne
rect 6034 14254 7194 14271
rect 38 14245 1196 14254
tri 1196 14245 1205 14254 nw
tri 5524 14245 5533 14254 ne
rect 5533 14245 5752 14254
rect 38 14233 783 14245
rect 38 14199 51 14233
rect 85 14199 124 14233
rect 158 14199 197 14233
rect 231 14199 270 14233
rect 304 14199 343 14233
rect 377 14199 416 14233
rect 450 14199 489 14233
rect 523 14199 563 14233
rect 597 14199 637 14233
rect 671 14199 711 14233
rect 745 14211 783 14233
rect 817 14211 1031 14245
rect 1065 14211 1162 14245
tri 1162 14211 1196 14245 nw
tri 5533 14211 5567 14245 ne
rect 5567 14211 5588 14245
rect 5622 14211 5701 14245
rect 5735 14211 5752 14245
rect 745 14206 1157 14211
tri 1157 14206 1162 14211 nw
tri 5567 14206 5572 14211 ne
rect 5572 14206 5752 14211
tri 5752 14206 5800 14254 nw
tri 6034 14206 6082 14254 ne
rect 6082 14206 7194 14254
rect 745 14205 1156 14206
tri 1156 14205 1157 14206 nw
tri 5572 14205 5573 14206 ne
rect 5573 14205 5751 14206
tri 5751 14205 5752 14206 nw
tri 6082 14205 6083 14206 ne
rect 6083 14205 7129 14206
rect 745 14202 1153 14205
tri 1153 14202 1156 14205 nw
tri 5573 14202 5576 14205 ne
rect 5576 14202 5748 14205
tri 5748 14202 5751 14205 nw
tri 6083 14202 6086 14205 ne
rect 6086 14202 6259 14205
rect 745 14199 1122 14202
rect 38 14171 1122 14199
tri 1122 14171 1153 14202 nw
tri 6086 14171 6117 14202 ne
rect 6117 14171 6259 14202
rect 6293 14171 6571 14205
rect 6605 14171 6883 14205
rect 6917 14172 7129 14205
rect 7163 14172 7194 14206
rect 6917 14171 7194 14172
rect 38 14168 1031 14171
rect 38 14161 783 14168
rect 38 14127 51 14161
rect 85 14127 124 14161
rect 158 14127 197 14161
rect 231 14127 270 14161
rect 304 14127 343 14161
rect 377 14127 416 14161
rect 450 14127 489 14161
rect 523 14127 563 14161
rect 597 14127 637 14161
rect 671 14127 711 14161
rect 745 14134 783 14161
rect 817 14137 1031 14168
rect 1065 14159 1110 14171
tri 1110 14159 1122 14171 nw
tri 6117 14159 6129 14171 ne
rect 6129 14160 7194 14171
tri 7194 14160 7306 14272 nw
rect 6129 14159 7193 14160
tri 7193 14159 7194 14160 nw
rect 1065 14158 1109 14159
tri 1109 14158 1110 14159 nw
tri 6129 14158 6130 14159 ne
rect 6130 14158 7192 14159
tri 7192 14158 7193 14159 nw
rect 1065 14137 1076 14158
rect 817 14134 1076 14137
rect 745 14127 1076 14134
rect 38 14125 1076 14127
tri 1076 14125 1109 14158 nw
rect 38 14091 996 14125
rect 38 14089 783 14091
rect 38 14055 51 14089
rect 85 14055 124 14089
rect 158 14055 197 14089
rect 231 14055 270 14089
rect 304 14055 343 14089
rect 377 14055 416 14089
rect 450 14055 489 14089
rect 523 14055 563 14089
rect 597 14055 637 14089
rect 671 14055 711 14089
rect 745 14057 783 14089
rect 817 14057 996 14091
rect 745 14055 996 14057
rect 38 14045 996 14055
tri 996 14045 1076 14125 nw
rect 31468 14066 31674 14072
rect 38 14044 995 14045
tri 995 14044 996 14045 nw
rect 31468 14014 31469 14066
rect 31521 14014 31545 14066
rect 31597 14014 31621 14066
rect 31673 14014 31674 14066
rect 31468 14002 31674 14014
rect 31468 13950 31469 14002
rect 31521 13950 31545 14002
rect 31597 13950 31621 14002
rect 31673 13950 31674 14002
rect 31468 13938 31674 13950
rect 31468 13886 31469 13938
rect 31521 13886 31545 13938
rect 31597 13886 31621 13938
rect 31673 13886 31674 13938
rect 31468 13874 31674 13886
rect 31468 13822 31469 13874
rect 31521 13822 31545 13874
rect 31597 13822 31621 13874
rect 31673 13822 31674 13874
rect 31468 13810 31674 13822
rect 31468 13758 31469 13810
rect 31521 13758 31545 13810
rect 31597 13758 31621 13810
rect 31673 13758 31674 13810
rect 31468 13745 31674 13758
rect 31468 13693 31469 13745
rect 31521 13693 31545 13745
rect 31597 13693 31621 13745
rect 31673 13693 31674 13745
rect 31468 13680 31674 13693
rect 31468 13628 31469 13680
rect 31521 13628 31545 13680
rect 31597 13628 31621 13680
rect 31673 13628 31674 13680
rect 31468 13615 31674 13628
rect 31468 13563 31469 13615
rect 31521 13563 31545 13615
rect 31597 13563 31621 13615
rect 31673 13563 31674 13615
rect 31468 13550 31674 13563
rect 31468 13498 31469 13550
rect 31521 13498 31545 13550
rect 31597 13498 31621 13550
rect 31673 13498 31674 13550
rect 31468 13485 31674 13498
rect 31468 13433 31469 13485
rect 31521 13433 31545 13485
rect 31597 13433 31621 13485
rect 31673 13433 31674 13485
rect 31468 13420 31674 13433
rect 31468 13368 31469 13420
rect 31521 13368 31545 13420
rect 31597 13368 31621 13420
rect 31673 13368 31674 13420
rect 31468 13355 31674 13368
rect 31468 13303 31469 13355
rect 31521 13303 31545 13355
rect 31597 13303 31621 13355
rect 31673 13303 31674 13355
rect 31468 13290 31674 13303
rect 31468 13238 31469 13290
rect 31521 13238 31545 13290
rect 31597 13238 31621 13290
rect 31673 13238 31674 13290
rect 31468 13225 31674 13238
rect 31468 13173 31469 13225
rect 31521 13173 31545 13225
rect 31597 13173 31621 13225
rect 31673 13173 31674 13225
rect 31468 13160 31674 13173
rect 31468 13108 31469 13160
rect 31521 13108 31545 13160
rect 31597 13108 31621 13160
rect 31673 13108 31674 13160
rect 31468 13095 31674 13108
rect 31468 13043 31469 13095
rect 31521 13043 31545 13095
rect 31597 13043 31621 13095
rect 31673 13043 31674 13095
rect 15143 13032 16541 13033
rect 15143 12980 15149 13032
rect 15201 12980 15213 13032
rect 15265 12980 15277 13032
rect 15329 12980 15341 13032
rect 15393 12980 15405 13032
rect 15457 12980 16541 13032
rect 15143 12962 16541 12980
rect 15143 12910 15149 12962
rect 15201 12910 15213 12962
rect 15265 12910 15277 12962
rect 15329 12910 15341 12962
rect 15393 12910 15405 12962
rect 15457 12910 16541 12962
rect 15143 12892 16541 12910
rect 15143 12840 15149 12892
rect 15201 12840 15213 12892
rect 15265 12840 15277 12892
rect 15329 12840 15341 12892
rect 15393 12840 15405 12892
rect 15457 12840 16541 12892
rect 15143 12822 16541 12840
rect 15143 12770 15149 12822
rect 15201 12770 15213 12822
rect 15265 12770 15277 12822
rect 15329 12770 15341 12822
rect 15393 12770 15405 12822
rect 15457 12770 16541 12822
rect 15143 12769 16541 12770
rect 31468 13030 31674 13043
rect 31468 12978 31469 13030
rect 31521 12978 31545 13030
rect 31597 12978 31621 13030
rect 31673 12978 31674 13030
rect 31468 12965 31674 12978
rect 31468 12913 31469 12965
rect 31521 12913 31545 12965
rect 31597 12913 31621 12965
rect 31673 12913 31674 12965
rect 31468 12900 31674 12913
rect 31468 12848 31469 12900
rect 31521 12848 31545 12900
rect 31597 12848 31621 12900
rect 31673 12848 31674 12900
rect 31468 12835 31674 12848
rect 31468 12783 31469 12835
rect 31521 12783 31545 12835
rect 31597 12783 31621 12835
rect 31673 12783 31674 12835
rect 31468 12770 31674 12783
rect 31468 12718 31469 12770
rect 31521 12718 31545 12770
rect 31597 12718 31621 12770
rect 31673 12718 31674 12770
rect 31468 12705 31674 12718
rect 31468 12653 31469 12705
rect 31521 12653 31545 12705
rect 31597 12653 31621 12705
rect 31673 12653 31674 12705
rect 31468 12640 31674 12653
rect 31468 12588 31469 12640
rect 31521 12588 31545 12640
rect 31597 12588 31621 12640
rect 31673 12588 31674 12640
rect 31468 12575 31674 12588
rect 31468 12523 31469 12575
rect 31521 12523 31545 12575
rect 31597 12523 31621 12575
rect 31673 12523 31674 12575
rect 31468 12510 31674 12523
rect 31468 12458 31469 12510
rect 31521 12458 31545 12510
rect 31597 12458 31621 12510
rect 31673 12458 31674 12510
rect 31468 12445 31674 12458
rect 31468 12393 31469 12445
rect 31521 12393 31545 12445
rect 31597 12393 31621 12445
rect 31673 12393 31674 12445
rect 31468 12380 31674 12393
rect 31468 12328 31469 12380
rect 31521 12328 31545 12380
rect 31597 12328 31621 12380
rect 31673 12328 31674 12380
rect 31468 12315 31674 12328
rect 31468 12263 31469 12315
rect 31521 12263 31545 12315
rect 31597 12263 31621 12315
rect 31673 12263 31674 12315
rect 31468 12250 31674 12263
rect 31468 12198 31469 12250
rect 31521 12198 31545 12250
rect 31597 12198 31621 12250
rect 31673 12198 31674 12250
rect 31468 12185 31674 12198
rect 31468 12133 31469 12185
rect 31521 12133 31545 12185
rect 31597 12133 31621 12185
rect 31673 12133 31674 12185
rect 31468 12120 31674 12133
rect 31468 12068 31469 12120
rect 31521 12068 31545 12120
rect 31597 12068 31621 12120
rect 31673 12068 31674 12120
rect 31468 12055 31674 12068
rect 17608 12039 17901 12041
rect 17608 12037 18413 12039
rect 17608 11985 17617 12037
rect 17669 11985 17685 12037
rect 17737 11985 17752 12037
rect 17804 11985 17819 12037
rect 17871 11985 17886 12037
rect 17938 11985 17953 12037
rect 18005 11985 18020 12037
rect 18072 11985 18087 12037
rect 18139 11985 18154 12037
rect 18206 11985 18221 12037
rect 18273 11985 18288 12037
rect 18340 11985 18355 12037
rect 18407 11985 18413 12037
rect 17608 11965 18413 11985
rect 17608 11913 17617 11965
rect 17669 11913 17685 11965
rect 17737 11913 17752 11965
rect 17804 11913 17819 11965
rect 17871 11913 17886 11965
rect 17938 11913 17953 11965
rect 18005 11913 18020 11965
rect 18072 11913 18087 11965
rect 18139 11913 18154 11965
rect 18206 11913 18221 11965
rect 18273 11913 18288 11965
rect 18340 11913 18355 11965
rect 18407 11913 18413 11965
rect 17608 11893 18413 11913
rect 17608 11841 17617 11893
rect 17669 11841 17685 11893
rect 17737 11841 17752 11893
rect 17804 11841 17819 11893
rect 17871 11841 17886 11893
rect 17938 11841 17953 11893
rect 18005 11841 18020 11893
rect 18072 11841 18087 11893
rect 18139 11841 18154 11893
rect 18206 11841 18221 11893
rect 18273 11841 18288 11893
rect 18340 11841 18355 11893
rect 18407 11841 18413 11893
rect 17608 11821 18413 11841
rect 17608 11769 17617 11821
rect 17669 11769 17685 11821
rect 17737 11769 17752 11821
rect 17804 11769 17819 11821
rect 17871 11769 17886 11821
rect 17938 11769 17953 11821
rect 18005 11769 18020 11821
rect 18072 11769 18087 11821
rect 18139 11769 18154 11821
rect 18206 11769 18221 11821
rect 18273 11769 18288 11821
rect 18340 11769 18355 11821
rect 18407 11769 18413 11821
rect 17608 11767 18413 11769
rect 31468 12003 31469 12055
rect 31521 12003 31545 12055
rect 31597 12003 31621 12055
rect 31673 12003 31674 12055
rect 31468 11990 31674 12003
rect 31468 11938 31469 11990
rect 31521 11938 31545 11990
rect 31597 11938 31621 11990
rect 31673 11938 31674 11990
rect 31468 11925 31674 11938
rect 31468 11873 31469 11925
rect 31521 11873 31545 11925
rect 31597 11873 31621 11925
rect 31673 11873 31674 11925
rect 31468 11860 31674 11873
rect 31468 11808 31469 11860
rect 31521 11808 31545 11860
rect 31597 11808 31621 11860
rect 31673 11808 31674 11860
rect 31468 11795 31674 11808
rect 17608 11765 17901 11767
rect 31468 11743 31469 11795
rect 31521 11743 31545 11795
rect 31597 11743 31621 11795
rect 31673 11743 31674 11795
rect 31468 11730 31674 11743
rect 4073 11653 4079 11705
rect 4131 11653 4143 11705
rect 4195 11653 5115 11705
rect 5167 11653 5179 11705
rect 5231 11653 5237 11705
rect 31468 11678 31469 11730
rect 31521 11678 31545 11730
rect 31597 11678 31621 11730
rect 31673 11678 31674 11730
rect 31468 11665 31674 11678
rect 31468 11613 31469 11665
rect 31521 11613 31545 11665
rect 31597 11613 31621 11665
rect 31673 11613 31674 11665
rect 31468 11600 31674 11613
rect 19533 11582 20334 11589
rect 19533 11530 19836 11582
rect 19888 11530 19908 11582
rect 19960 11530 19979 11582
rect 20031 11530 20050 11582
rect 20102 11530 20121 11582
rect 20173 11530 20192 11582
rect 20244 11530 20263 11582
rect 20315 11530 20334 11582
rect 19533 11514 20334 11530
rect 19533 11462 19836 11514
rect 19888 11462 19908 11514
rect 19960 11462 19979 11514
rect 20031 11462 20050 11514
rect 20102 11462 20121 11514
rect 20173 11462 20192 11514
rect 20244 11462 20263 11514
rect 20315 11462 20334 11514
rect 19533 11446 20334 11462
rect 19533 11394 19836 11446
rect 19888 11394 19908 11446
rect 19960 11394 19979 11446
rect 20031 11394 20050 11446
rect 20102 11394 20121 11446
rect 20173 11394 20192 11446
rect 20244 11394 20263 11446
rect 20315 11394 20334 11446
tri 15891 11274 15999 11382 se
rect 19533 11378 20334 11394
rect 19533 11326 19836 11378
rect 19888 11326 19908 11378
rect 19960 11326 19979 11378
rect 20031 11326 20050 11378
rect 20102 11326 20121 11378
rect 20173 11326 20192 11378
rect 20244 11326 20263 11378
rect 20315 11326 20334 11378
rect 19533 11313 20334 11326
rect 31468 11548 31469 11600
rect 31521 11548 31545 11600
rect 31597 11548 31621 11600
rect 31673 11548 31674 11600
rect 31468 11535 31674 11548
rect 31468 11483 31469 11535
rect 31521 11483 31545 11535
rect 31597 11483 31621 11535
rect 31673 11483 31674 11535
rect 31468 11470 31674 11483
rect 31468 11418 31469 11470
rect 31521 11418 31545 11470
rect 31597 11418 31621 11470
rect 31673 11418 31674 11470
rect 31468 11405 31674 11418
rect 31468 11353 31469 11405
rect 31521 11353 31545 11405
rect 31597 11353 31621 11405
rect 31673 11353 31674 11405
rect 31468 11340 31674 11353
tri 13881 11271 13884 11274 se
rect 13884 11271 13890 11274
rect 13072 11265 13890 11271
rect 13942 11265 13981 11274
rect 14033 11265 14071 11274
rect 14123 11271 14129 11274
tri 14129 11271 14132 11274 sw
tri 14415 11271 14418 11274 se
rect 14418 11271 14424 11274
rect 14123 11265 14424 11271
rect 14476 11265 14489 11274
rect 14541 11265 14553 11274
rect 13072 11231 13084 11265
rect 13118 11231 13157 11265
rect 13191 11231 13230 11265
rect 13264 11231 13303 11265
rect 13337 11231 13376 11265
rect 13410 11231 13449 11265
rect 13483 11231 13522 11265
rect 13556 11231 13595 11265
rect 13629 11231 13668 11265
rect 13702 11231 13741 11265
rect 13775 11231 13814 11265
rect 13848 11231 13887 11265
rect 13942 11231 13960 11265
rect 14067 11231 14071 11265
rect 14140 11231 14179 11265
rect 14213 11231 14252 11265
rect 14286 11231 14325 11265
rect 14359 11231 14398 11265
rect 14541 11231 14544 11265
rect 13072 11225 13890 11231
tri 13881 11222 13884 11225 ne
rect 13884 11222 13890 11225
rect 13942 11222 13981 11231
rect 14033 11222 14071 11231
rect 14123 11225 14424 11231
rect 14123 11222 14129 11225
tri 14129 11222 14132 11225 nw
tri 14415 11222 14418 11225 ne
rect 14418 11222 14424 11225
rect 14476 11222 14489 11231
rect 14541 11222 14553 11231
rect 14605 11222 14617 11274
rect 14669 11222 14681 11274
rect 14733 11271 14739 11274
tri 14739 11271 14742 11274 sw
tri 15888 11271 15891 11274 se
rect 15891 11271 15999 11274
rect 14733 11265 15999 11271
rect 14733 11231 14763 11265
rect 14797 11231 14836 11265
rect 14870 11231 14909 11265
rect 14943 11231 14982 11265
rect 15016 11231 15055 11265
rect 15089 11231 15128 11265
rect 15162 11231 15201 11265
rect 15235 11231 15273 11265
rect 15307 11231 15345 11265
rect 15379 11231 15417 11265
rect 15451 11231 15489 11265
rect 15523 11231 15561 11265
rect 15595 11231 15633 11265
rect 15667 11231 15705 11265
rect 15739 11231 15777 11265
rect 15811 11231 15849 11265
rect 15883 11231 15921 11265
rect 15955 11231 15999 11265
rect 14733 11225 15999 11231
rect 14733 11222 14739 11225
tri 14739 11222 14742 11225 nw
tri 15976 11222 15979 11225 ne
rect 15979 11222 15999 11225
tri 15979 11202 15999 11222 ne
rect 31468 11288 31469 11340
rect 31521 11288 31545 11340
rect 31597 11288 31621 11340
rect 31673 11288 31674 11340
rect 31468 11275 31674 11288
rect 31468 11223 31469 11275
rect 31521 11223 31545 11275
rect 31597 11223 31621 11275
rect 31673 11223 31674 11275
rect 31468 11210 31674 11223
rect 31468 11158 31469 11210
rect 31521 11158 31545 11210
rect 31597 11158 31621 11210
rect 31673 11158 31674 11210
rect 4084 11142 4202 11148
rect 4084 11090 4085 11142
rect 4137 11090 4149 11142
rect 4201 11090 4202 11142
rect 4084 11084 4202 11090
rect 31468 11145 31674 11158
rect 31468 11093 31469 11145
rect 31521 11093 31545 11145
rect 31597 11093 31621 11145
rect 31673 11093 31674 11145
rect 31468 11087 31674 11093
rect 4421 10937 6236 10944
rect 4421 10903 4433 10937
rect 4467 10903 4507 10937
rect 4541 10903 4581 10937
rect 4615 10903 4655 10937
rect 4689 10903 4729 10937
rect 4763 10903 4803 10937
rect 4837 10903 4876 10937
rect 4910 10903 4949 10937
rect 4983 10903 5022 10937
rect 5056 10903 5095 10937
rect 5129 10903 5168 10937
rect 5202 10903 5241 10937
rect 5275 10903 5314 10937
rect 5348 10903 5387 10937
rect 5421 10903 5460 10937
rect 5494 10903 5533 10937
rect 5567 10903 5606 10937
rect 5640 10903 5679 10937
rect 5713 10903 5752 10937
rect 5786 10903 5825 10937
rect 5859 10903 5898 10937
rect 5932 10903 5971 10937
rect 6005 10903 6044 10937
rect 6078 10903 6117 10937
rect 6151 10903 6190 10937
rect 6224 10903 6236 10937
rect 4421 10861 6236 10903
rect 4421 10827 4433 10861
rect 4467 10827 4507 10861
rect 4541 10827 4581 10861
rect 4615 10827 4655 10861
rect 4689 10827 4729 10861
rect 4763 10827 4803 10861
rect 4837 10827 4876 10861
rect 4910 10827 4949 10861
rect 4983 10827 5022 10861
rect 5056 10827 5095 10861
rect 5129 10827 5168 10861
rect 5202 10827 5241 10861
rect 5275 10827 5314 10861
rect 5348 10827 5387 10861
rect 5421 10827 5460 10861
rect 5494 10827 5533 10861
rect 5567 10827 5606 10861
rect 5640 10827 5679 10861
rect 5713 10827 5752 10861
rect 5786 10827 5825 10861
rect 5859 10827 5898 10861
rect 5932 10827 5971 10861
rect 6005 10827 6044 10861
rect 6078 10827 6117 10861
rect 6151 10827 6190 10861
rect 6224 10827 6236 10861
rect 4421 10785 6236 10827
rect 4421 10751 4433 10785
rect 4467 10751 4507 10785
rect 4541 10751 4581 10785
rect 4615 10751 4655 10785
rect 4689 10751 4729 10785
rect 4763 10751 4803 10785
rect 4837 10751 4876 10785
rect 4910 10751 4949 10785
rect 4983 10751 5022 10785
rect 5056 10751 5095 10785
rect 5129 10751 5168 10785
rect 5202 10751 5241 10785
rect 5275 10751 5314 10785
rect 5348 10751 5387 10785
rect 5421 10751 5460 10785
rect 5494 10751 5533 10785
rect 5567 10751 5606 10785
rect 5640 10751 5679 10785
rect 5713 10751 5752 10785
rect 5786 10751 5825 10785
rect 5859 10751 5898 10785
rect 5932 10751 5971 10785
rect 6005 10751 6044 10785
rect 6078 10751 6117 10785
rect 6151 10751 6190 10785
rect 6224 10751 6236 10785
rect 4421 10744 6236 10751
rect 13352 10934 15894 10940
rect 13352 10900 13364 10934
rect 13398 10900 13438 10934
rect 13472 10900 13512 10934
rect 13546 10900 13585 10934
rect 13619 10900 13658 10934
rect 13692 10900 13731 10934
rect 13765 10900 13804 10934
rect 13838 10900 13877 10934
rect 13911 10900 13950 10934
rect 13984 10900 14023 10934
rect 14057 10900 14096 10934
rect 14130 10900 14169 10934
rect 14203 10900 14242 10934
rect 14276 10900 14315 10934
rect 14349 10900 14388 10934
rect 14422 10900 14461 10934
rect 14495 10900 14534 10934
rect 14568 10900 14607 10934
rect 14641 10900 14680 10934
rect 14714 10900 14753 10934
rect 14787 10900 14826 10934
rect 14860 10900 14899 10934
rect 14933 10900 14972 10934
rect 15006 10900 15045 10934
rect 15079 10900 15118 10934
rect 15152 10900 15191 10934
rect 15225 10900 15264 10934
rect 15298 10900 15337 10934
rect 15371 10900 15410 10934
rect 15444 10900 15483 10934
rect 15517 10900 15556 10934
rect 15590 10900 15629 10934
rect 15663 10900 15702 10934
rect 15736 10900 15775 10934
rect 15809 10900 15848 10934
rect 15882 10900 15894 10934
rect 13352 10860 15894 10900
rect 13352 10826 13364 10860
rect 13398 10826 13438 10860
rect 13472 10826 13512 10860
rect 13546 10826 13585 10860
rect 13619 10826 13658 10860
rect 13692 10826 13731 10860
rect 13765 10826 13804 10860
rect 13838 10826 13877 10860
rect 13911 10826 13950 10860
rect 13984 10826 14023 10860
rect 14057 10826 14096 10860
rect 14130 10826 14169 10860
rect 14203 10826 14242 10860
rect 14276 10826 14315 10860
rect 14349 10826 14388 10860
rect 14422 10826 14461 10860
rect 14495 10826 14534 10860
rect 14568 10826 14607 10860
rect 14641 10826 14680 10860
rect 14714 10826 14753 10860
rect 14787 10826 14826 10860
rect 14860 10826 14899 10860
rect 14933 10826 14972 10860
rect 15006 10826 15045 10860
rect 15079 10826 15118 10860
rect 15152 10826 15191 10860
rect 15225 10826 15264 10860
rect 15298 10826 15337 10860
rect 15371 10826 15410 10860
rect 15444 10826 15483 10860
rect 15517 10826 15556 10860
rect 15590 10826 15629 10860
rect 15663 10826 15702 10860
rect 15736 10826 15775 10860
rect 15809 10826 15848 10860
rect 15882 10826 15894 10860
rect 13352 10786 15894 10826
rect 13352 10752 13364 10786
rect 13398 10752 13438 10786
rect 13472 10752 13512 10786
rect 13546 10752 13585 10786
rect 13619 10752 13658 10786
rect 13692 10752 13731 10786
rect 13765 10752 13804 10786
rect 13838 10752 13877 10786
rect 13911 10752 13950 10786
rect 13984 10752 14023 10786
rect 14057 10752 14096 10786
rect 14130 10752 14169 10786
rect 14203 10752 14242 10786
rect 14276 10752 14315 10786
rect 14349 10752 14388 10786
rect 14422 10752 14461 10786
rect 14495 10752 14534 10786
rect 14568 10752 14607 10786
rect 14641 10752 14680 10786
rect 14714 10752 14753 10786
rect 14787 10752 14826 10786
rect 14860 10752 14899 10786
rect 14933 10752 14972 10786
rect 15006 10752 15045 10786
rect 15079 10752 15118 10786
rect 15152 10752 15191 10786
rect 15225 10752 15264 10786
rect 15298 10752 15337 10786
rect 15371 10752 15410 10786
rect 15444 10752 15483 10786
rect 15517 10752 15556 10786
rect 15590 10752 15629 10786
rect 15663 10752 15702 10786
rect 15736 10752 15775 10786
rect 15809 10752 15848 10786
rect 15882 10752 15894 10786
rect 13352 10746 15894 10752
tri 13881 10548 13884 10551 se
rect 13884 10548 13890 10551
rect 13104 10542 13890 10548
rect 13942 10542 13981 10551
rect 14033 10542 14071 10551
rect 14123 10548 14129 10551
tri 14129 10548 14132 10551 sw
tri 14415 10548 14418 10551 se
rect 14418 10548 14424 10551
rect 14123 10542 14424 10548
rect 14476 10542 14489 10551
rect 14541 10542 14553 10551
rect 14605 10542 14617 10551
rect 14669 10542 14681 10551
rect 14733 10548 14739 10551
tri 14739 10548 14742 10551 sw
rect 14733 10542 15745 10548
rect 13104 10508 13116 10542
rect 13150 10508 13190 10542
rect 13224 10508 13264 10542
rect 13298 10508 13338 10542
rect 13372 10508 13412 10542
rect 13446 10508 13486 10542
rect 13520 10508 13560 10542
rect 13594 10508 13634 10542
rect 13668 10508 13708 10542
rect 13742 10508 13782 10542
rect 13816 10508 13856 10542
rect 13964 10508 13981 10542
rect 14038 10508 14071 10542
rect 14123 10508 14152 10542
rect 14186 10508 14226 10542
rect 14260 10508 14300 10542
rect 14334 10508 14374 10542
rect 14408 10508 14424 10542
rect 14482 10508 14489 10542
rect 14669 10508 14670 10542
rect 14733 10508 14744 10542
rect 14778 10508 14818 10542
rect 14852 10508 14892 10542
rect 14926 10508 14966 10542
rect 15000 10508 15040 10542
rect 15074 10508 15114 10542
rect 15148 10508 15188 10542
rect 15222 10508 15261 10542
rect 15295 10508 15334 10542
rect 15368 10508 15407 10542
rect 15441 10508 15480 10542
rect 15514 10508 15553 10542
rect 15587 10508 15626 10542
rect 15660 10508 15699 10542
rect 15733 10508 15745 10542
rect 13104 10502 13890 10508
tri 13881 10499 13884 10502 ne
rect 13884 10499 13890 10502
rect 13942 10499 13981 10508
rect 14033 10499 14071 10508
rect 14123 10502 14424 10508
rect 14123 10499 14129 10502
tri 14129 10499 14132 10502 nw
tri 14415 10499 14418 10502 ne
rect 14418 10499 14424 10502
rect 14476 10499 14489 10508
rect 14541 10499 14553 10508
rect 14605 10499 14617 10508
rect 14669 10499 14681 10508
rect 14733 10502 15745 10508
rect 14733 10499 14739 10502
tri 14739 10499 14742 10502 nw
rect 6019 9871 6025 9923
rect 6077 9871 6089 9923
rect 6141 9877 6891 9923
rect 6141 9871 6147 9877
tri 6147 9871 6153 9877 nw
rect 5623 9221 5675 9227
rect 6114 9195 6123 9247
rect 6175 9195 6187 9247
rect 6239 9227 6245 9247
tri 10045 9244 10048 9247 se
rect 10048 9244 10054 9247
tri 6245 9227 6262 9244 sw
tri 10028 9227 10045 9244 se
rect 10045 9227 10054 9244
rect 6239 9195 10054 9227
rect 10106 9195 10118 9247
rect 10170 9195 10176 9247
rect 10779 9204 10785 9256
rect 10837 9204 10849 9256
rect 10901 9204 10907 9256
rect 5623 9157 5675 9169
rect 5623 9099 5675 9105
rect 18531 8371 18537 8423
rect 18589 8371 18601 8423
rect 18653 8371 18665 8423
rect 18717 8371 18729 8423
rect 18781 8371 18793 8423
rect 18845 8371 18857 8423
rect 18909 8371 18915 8423
rect 5298 7488 5350 7497
tri 5350 7481 5366 7497 sw
rect 5350 7436 6123 7481
rect 5298 7429 6123 7436
rect 6175 7429 6187 7481
rect 6239 7429 6245 7481
rect 5298 7424 5350 7429
tri 5350 7395 5384 7429 nw
rect 5298 7366 5350 7372
rect 13259 7379 13375 7385
rect 13311 7327 13323 7379
rect 13259 7321 13375 7327
rect -593 7009 -587 7061
rect -535 7009 -505 7061
rect -453 7009 -423 7061
rect -371 7009 -341 7061
rect -289 7009 -259 7061
rect -207 7009 -201 7061
tri -600 7001 -593 7008 se
rect -593 6997 -201 7009
tri -201 7001 -198 7004 sw
rect -593 6945 -587 6997
rect -535 6945 -505 6997
rect -453 6945 -423 6997
rect -371 6945 -341 6997
rect -289 6945 -259 6997
rect -207 6945 -201 6997
rect 18300 6480 18341 6647
rect 18343 6480 18384 6647
rect 23952 6302 23958 6354
rect 24010 6302 24042 6354
rect 24094 6302 24126 6354
rect 24178 6302 24209 6354
rect 24261 6302 24267 6354
rect 23952 6288 24267 6302
rect 23952 6236 23958 6288
rect 24010 6236 24042 6288
rect 24094 6236 24126 6288
rect 24178 6236 24209 6288
rect 24261 6236 24267 6288
rect 23952 6222 24267 6236
rect 23952 6170 23958 6222
rect 24010 6170 24042 6222
rect 24094 6170 24126 6222
rect 24178 6170 24209 6222
rect 24261 6170 24267 6222
rect 8303 5997 8319 6049
rect 76 5764 2263 5770
rect 192 5763 2263 5764
rect 192 5648 2145 5763
rect 76 5647 2145 5648
rect 2261 5647 2263 5763
rect 32274 5699 32301 5751
rect 32729 5699 32781 5750
rect 76 5642 2263 5647
rect 2145 5641 2261 5642
rect -600 4816 -200 4846
rect -600 4764 -594 4816
rect -542 4764 -510 4816
rect -458 4764 -426 4816
rect -374 4764 -342 4816
rect -290 4764 -258 4816
rect -206 4764 -200 4816
rect -600 4734 -200 4764
tri 4803 3214 4847 3258 se
rect 4847 3252 4899 3258
rect 3582 3200 4847 3214
rect 3582 3188 4899 3200
rect 3582 3136 4847 3188
rect 3582 3130 4899 3136
tri 3582 3074 3638 3130 nw
rect 5964 2536 6126 2542
rect 5964 2484 5987 2536
rect 6039 2484 6051 2536
rect 6103 2484 6126 2536
rect 5964 2467 6126 2484
rect 5964 2415 5987 2467
rect 6039 2415 6051 2467
rect 6103 2415 6126 2467
rect 5964 2398 6126 2415
rect 5964 2346 5987 2398
rect 6039 2346 6051 2398
rect 6103 2346 6126 2398
rect 5964 2340 6126 2346
rect 5988 2205 6127 2212
rect 5988 2153 5994 2205
rect 6046 2153 6069 2205
rect 6121 2153 6127 2205
rect 5988 2146 6127 2153
rect 513 1323 519 1503
rect 635 1323 641 1503
rect 1228 1323 1234 1503
rect 1350 1323 1356 1503
rect 1855 1323 1861 1503
rect 1977 1323 1983 1503
rect 2567 1323 2573 1503
rect 2689 1323 2695 1503
rect 3022 1195 3150 2056
rect 8541 1740 8737 1746
rect 5964 1705 6126 1711
rect 5964 1653 5987 1705
rect 6039 1653 6051 1705
rect 6103 1653 6126 1705
rect 5964 1625 6126 1653
rect 5964 1573 5987 1625
rect 6039 1573 6051 1625
rect 6103 1573 6126 1625
rect 5964 1567 6126 1573
rect 8541 1688 8549 1740
rect 8601 1688 8613 1740
rect 8665 1688 8677 1740
rect 8729 1688 8737 1740
rect 8541 1671 8737 1688
rect 8541 1619 8549 1671
rect 8601 1619 8613 1671
rect 8665 1619 8677 1671
rect 8729 1619 8737 1671
rect 8541 1602 8737 1619
rect 8541 1550 8549 1602
rect 8601 1550 8613 1602
rect 8665 1550 8677 1602
rect 8729 1550 8737 1602
rect 8541 1544 8737 1550
<< rmetal1 >>
rect 18341 6480 18343 6647
<< via1 >>
rect -2502 43637 -2450 43689
rect -2438 43637 -2386 43689
rect -2374 43637 -2322 43689
rect -2310 43637 -2258 43689
rect -2246 43637 -2194 43689
rect -2182 43637 -2130 43689
rect -2118 43637 -2066 43689
rect -2054 43637 -2002 43689
rect -1990 43637 -1938 43689
rect -1926 43637 -1874 43689
rect -1862 43637 -1810 43689
rect -1798 43637 -1746 43689
rect -1734 43637 -1682 43689
rect -1670 43637 -1618 43689
rect -1606 43637 -1554 43689
rect -1542 43637 -1490 43689
rect -1478 43637 -1426 43689
rect -1414 43637 -1362 43689
rect -1350 43637 -1298 43689
rect -1286 43637 -1234 43689
rect -1222 43637 -1170 43689
rect -1158 43637 -1106 43689
rect -1094 43637 -1042 43689
rect -1030 43637 -978 43689
rect -966 43637 -914 43689
rect -902 43637 -850 43689
rect -838 43637 -786 43689
rect -774 43637 -722 43689
rect -710 43637 -658 43689
rect -2502 43571 -2450 43623
rect -2438 43571 -2386 43623
rect -2374 43571 -2322 43623
rect -2310 43571 -2258 43623
rect -2246 43571 -2194 43623
rect -2182 43571 -2130 43623
rect -2118 43571 -2066 43623
rect -2054 43571 -2002 43623
rect -1990 43571 -1938 43623
rect -1926 43571 -1874 43623
rect -1862 43571 -1810 43623
rect -1798 43571 -1746 43623
rect -1734 43571 -1682 43623
rect -1670 43571 -1618 43623
rect -1606 43571 -1554 43623
rect -1542 43571 -1490 43623
rect -1478 43571 -1426 43623
rect -1414 43571 -1362 43623
rect -1350 43571 -1298 43623
rect -1286 43571 -1234 43623
rect -1222 43571 -1170 43623
rect -1158 43571 -1106 43623
rect -1094 43571 -1042 43623
rect -1030 43571 -978 43623
rect -966 43571 -914 43623
rect -902 43571 -850 43623
rect -838 43571 -786 43623
rect -774 43571 -722 43623
rect -710 43571 -658 43623
rect -2502 43505 -2450 43557
rect -2438 43505 -2386 43557
rect -2374 43505 -2322 43557
rect -2310 43505 -2258 43557
rect -2246 43505 -2194 43557
rect -2182 43505 -2130 43557
rect -2118 43505 -2066 43557
rect -2054 43505 -2002 43557
rect -1990 43505 -1938 43557
rect -1926 43505 -1874 43557
rect -1862 43505 -1810 43557
rect -1798 43505 -1746 43557
rect -1734 43505 -1682 43557
rect -1670 43505 -1618 43557
rect -1606 43505 -1554 43557
rect -1542 43505 -1490 43557
rect -1478 43505 -1426 43557
rect -1414 43505 -1362 43557
rect -1350 43505 -1298 43557
rect -1286 43505 -1234 43557
rect -1222 43505 -1170 43557
rect -1158 43505 -1106 43557
rect -1094 43505 -1042 43557
rect -1030 43505 -978 43557
rect -966 43505 -914 43557
rect -902 43505 -850 43557
rect -838 43505 -786 43557
rect -774 43505 -722 43557
rect -710 43505 -658 43557
rect -2502 43439 -2450 43491
rect -2438 43439 -2386 43491
rect -2374 43439 -2322 43491
rect -2310 43439 -2258 43491
rect -2246 43439 -2194 43491
rect -2182 43439 -2130 43491
rect -2118 43439 -2066 43491
rect -2054 43439 -2002 43491
rect -1990 43439 -1938 43491
rect -1926 43439 -1874 43491
rect -1862 43439 -1810 43491
rect -1798 43439 -1746 43491
rect -1734 43439 -1682 43491
rect -1670 43439 -1618 43491
rect -1606 43439 -1554 43491
rect -1542 43439 -1490 43491
rect -1478 43439 -1426 43491
rect -1414 43439 -1362 43491
rect -1350 43439 -1298 43491
rect -1286 43439 -1234 43491
rect -1222 43439 -1170 43491
rect -1158 43439 -1106 43491
rect -1094 43439 -1042 43491
rect -1030 43439 -978 43491
rect -966 43439 -914 43491
rect -902 43439 -850 43491
rect -838 43439 -786 43491
rect -774 43439 -722 43491
rect -710 43439 -658 43491
rect -2502 43373 -2450 43425
rect -2438 43373 -2386 43425
rect -2374 43373 -2322 43425
rect -2310 43373 -2258 43425
rect -2246 43373 -2194 43425
rect -2182 43373 -2130 43425
rect -2118 43373 -2066 43425
rect -2054 43373 -2002 43425
rect -1990 43373 -1938 43425
rect -1926 43373 -1874 43425
rect -1862 43373 -1810 43425
rect -1798 43373 -1746 43425
rect -1734 43373 -1682 43425
rect -1670 43373 -1618 43425
rect -1606 43373 -1554 43425
rect -1542 43373 -1490 43425
rect -1478 43373 -1426 43425
rect -1414 43373 -1362 43425
rect -1350 43373 -1298 43425
rect -1286 43373 -1234 43425
rect -1222 43373 -1170 43425
rect -1158 43373 -1106 43425
rect -1094 43373 -1042 43425
rect -1030 43373 -978 43425
rect -966 43373 -914 43425
rect -902 43373 -850 43425
rect -838 43373 -786 43425
rect -774 43373 -722 43425
rect -710 43373 -658 43425
rect -2502 43307 -2450 43359
rect -2438 43307 -2386 43359
rect -2374 43307 -2322 43359
rect -2310 43307 -2258 43359
rect -2246 43307 -2194 43359
rect -2182 43307 -2130 43359
rect -2118 43307 -2066 43359
rect -2054 43307 -2002 43359
rect -1990 43307 -1938 43359
rect -1926 43307 -1874 43359
rect -1862 43307 -1810 43359
rect -1798 43307 -1746 43359
rect -1734 43307 -1682 43359
rect -1670 43307 -1618 43359
rect -1606 43307 -1554 43359
rect -1542 43307 -1490 43359
rect -1478 43307 -1426 43359
rect -1414 43307 -1362 43359
rect -1350 43307 -1298 43359
rect -1286 43307 -1234 43359
rect -1222 43307 -1170 43359
rect -1158 43307 -1106 43359
rect -1094 43307 -1042 43359
rect -1030 43307 -978 43359
rect -966 43307 -914 43359
rect -902 43307 -850 43359
rect -838 43307 -786 43359
rect -774 43307 -722 43359
rect -710 43307 -658 43359
rect -2502 43241 -2450 43293
rect -2438 43241 -2386 43293
rect -2374 43241 -2322 43293
rect -2310 43241 -2258 43293
rect -2246 43241 -2194 43293
rect -2182 43241 -2130 43293
rect -2118 43241 -2066 43293
rect -2054 43241 -2002 43293
rect -1990 43241 -1938 43293
rect -1926 43241 -1874 43293
rect -1862 43241 -1810 43293
rect -1798 43241 -1746 43293
rect -1734 43241 -1682 43293
rect -1670 43241 -1618 43293
rect -1606 43241 -1554 43293
rect -1542 43241 -1490 43293
rect -1478 43241 -1426 43293
rect -1414 43241 -1362 43293
rect -1350 43241 -1298 43293
rect -1286 43241 -1234 43293
rect -1222 43241 -1170 43293
rect -1158 43241 -1106 43293
rect -1094 43241 -1042 43293
rect -1030 43241 -978 43293
rect -966 43241 -914 43293
rect -902 43241 -850 43293
rect -838 43241 -786 43293
rect -774 43241 -722 43293
rect -710 43241 -658 43293
rect -2502 43174 -2450 43226
rect -2438 43174 -2386 43226
rect -2374 43174 -2322 43226
rect -2310 43174 -2258 43226
rect -2246 43174 -2194 43226
rect -2182 43174 -2130 43226
rect -2118 43174 -2066 43226
rect -2054 43174 -2002 43226
rect -1990 43174 -1938 43226
rect -1926 43174 -1874 43226
rect -1862 43174 -1810 43226
rect -1798 43174 -1746 43226
rect -1734 43174 -1682 43226
rect -1670 43174 -1618 43226
rect -1606 43174 -1554 43226
rect -1542 43174 -1490 43226
rect -1478 43174 -1426 43226
rect -1414 43174 -1362 43226
rect -1350 43174 -1298 43226
rect -1286 43174 -1234 43226
rect -1222 43174 -1170 43226
rect -1158 43174 -1106 43226
rect -1094 43174 -1042 43226
rect -1030 43174 -978 43226
rect -966 43174 -914 43226
rect -902 43174 -850 43226
rect -838 43174 -786 43226
rect -774 43174 -722 43226
rect -710 43174 -658 43226
rect 646 43637 698 43689
rect 710 43637 762 43689
rect 774 43637 826 43689
rect 838 43637 890 43689
rect 902 43637 954 43689
rect 966 43637 1018 43689
rect 1030 43637 1082 43689
rect 646 43571 698 43623
rect 710 43571 762 43623
rect 774 43571 826 43623
rect 838 43571 890 43623
rect 902 43571 954 43623
rect 966 43571 1018 43623
rect 1030 43571 1082 43623
rect 646 43505 698 43557
rect 710 43505 762 43557
rect 774 43505 826 43557
rect 838 43505 890 43557
rect 902 43505 954 43557
rect 966 43505 1018 43557
rect 1030 43505 1082 43557
rect 646 43439 698 43491
rect 710 43439 762 43491
rect 774 43439 826 43491
rect 838 43439 890 43491
rect 902 43439 954 43491
rect 966 43439 1018 43491
rect 1030 43439 1082 43491
rect 646 43373 698 43425
rect 710 43373 762 43425
rect 774 43373 826 43425
rect 838 43373 890 43425
rect 902 43373 954 43425
rect 966 43373 1018 43425
rect 1030 43373 1082 43425
rect 646 43307 698 43359
rect 710 43307 762 43359
rect 774 43307 826 43359
rect 838 43307 890 43359
rect 902 43307 954 43359
rect 966 43307 1018 43359
rect 1030 43307 1082 43359
rect 646 43241 698 43293
rect 710 43241 762 43293
rect 774 43241 826 43293
rect 838 43241 890 43293
rect 902 43241 954 43293
rect 966 43241 1018 43293
rect 1030 43241 1082 43293
rect 646 43174 698 43226
rect 710 43174 762 43226
rect 774 43174 826 43226
rect 838 43174 890 43226
rect 902 43174 954 43226
rect 966 43174 1018 43226
rect 1030 43174 1082 43226
rect 31413 40072 31529 40188
rect 31599 39827 31715 39943
rect -1188 25109 -1136 25161
rect -1120 25109 -1068 25161
rect -1052 25109 -1000 25161
rect -984 25109 -932 25161
rect -916 25109 -864 25161
rect -848 25109 -796 25161
rect -780 25109 -728 25161
rect -712 25109 -660 25161
rect -644 25109 -592 25161
rect -1188 25045 -1136 25097
rect -1120 25045 -1068 25097
rect -1052 25045 -1000 25097
rect -984 25045 -932 25097
rect -916 25045 -864 25097
rect -848 25045 -796 25097
rect -780 25045 -728 25097
rect -712 25045 -660 25097
rect -644 25045 -592 25097
rect -1188 24981 -1136 25033
rect -1120 24981 -1068 25033
rect -1052 24981 -1000 25033
rect -984 24981 -932 25033
rect -916 24981 -864 25033
rect -848 24981 -796 25033
rect -780 24981 -728 25033
rect -712 24981 -660 25033
rect -644 24981 -592 25033
rect -1188 24917 -1136 24969
rect -1120 24917 -1068 24969
rect -1052 24917 -1000 24969
rect -984 24917 -932 24969
rect -916 24917 -864 24969
rect -848 24917 -796 24969
rect -780 24917 -728 24969
rect -712 24917 -660 24969
rect -644 24917 -592 24969
rect -1188 24853 -1136 24905
rect -1120 24853 -1068 24905
rect -1052 24853 -1000 24905
rect -984 24853 -932 24905
rect -916 24853 -864 24905
rect -848 24853 -796 24905
rect -780 24853 -728 24905
rect -712 24853 -660 24905
rect -644 24853 -592 24905
rect -1188 24789 -1136 24841
rect -1120 24789 -1068 24841
rect -1052 24789 -1000 24841
rect -984 24789 -932 24841
rect -916 24789 -864 24841
rect -848 24789 -796 24841
rect -780 24789 -728 24841
rect -712 24789 -660 24841
rect -644 24789 -592 24841
rect -1188 24725 -1136 24777
rect -1120 24725 -1068 24777
rect -1052 24725 -1000 24777
rect -984 24725 -932 24777
rect -916 24725 -864 24777
rect -848 24725 -796 24777
rect -780 24725 -728 24777
rect -712 24725 -660 24777
rect -644 24725 -592 24777
rect -1188 24661 -1136 24713
rect -1120 24661 -1068 24713
rect -1052 24661 -1000 24713
rect -984 24661 -932 24713
rect -916 24661 -864 24713
rect -848 24661 -796 24713
rect -780 24661 -728 24713
rect -712 24661 -660 24713
rect -644 24661 -592 24713
rect -1188 24597 -1136 24649
rect -1120 24597 -1068 24649
rect -1052 24597 -1000 24649
rect -984 24597 -932 24649
rect -916 24597 -864 24649
rect -848 24597 -796 24649
rect -780 24597 -728 24649
rect -712 24597 -660 24649
rect -644 24597 -592 24649
rect -1188 24533 -1136 24585
rect -1120 24533 -1068 24585
rect -1052 24533 -1000 24585
rect -984 24533 -932 24585
rect -916 24533 -864 24585
rect -848 24533 -796 24585
rect -780 24533 -728 24585
rect -712 24533 -660 24585
rect -644 24533 -592 24585
rect -1188 24469 -1136 24521
rect -1120 24469 -1068 24521
rect -1052 24469 -1000 24521
rect -984 24469 -932 24521
rect -916 24469 -864 24521
rect -848 24469 -796 24521
rect -780 24469 -728 24521
rect -712 24469 -660 24521
rect -644 24469 -592 24521
rect -1188 24405 -1136 24457
rect -1120 24405 -1068 24457
rect -1052 24405 -1000 24457
rect -984 24405 -932 24457
rect -916 24405 -864 24457
rect -848 24405 -796 24457
rect -780 24405 -728 24457
rect -712 24405 -660 24457
rect -644 24405 -592 24457
rect -1188 24341 -1136 24393
rect -1120 24341 -1068 24393
rect -1052 24341 -1000 24393
rect -984 24341 -932 24393
rect -916 24341 -864 24393
rect -848 24341 -796 24393
rect -780 24341 -728 24393
rect -712 24341 -660 24393
rect -644 24341 -592 24393
rect -1188 24277 -1136 24329
rect -1120 24277 -1068 24329
rect -1052 24277 -1000 24329
rect -984 24277 -932 24329
rect -916 24277 -864 24329
rect -848 24277 -796 24329
rect -780 24277 -728 24329
rect -712 24277 -660 24329
rect -644 24277 -592 24329
rect -1188 24213 -1136 24265
rect -1120 24213 -1068 24265
rect -1052 24213 -1000 24265
rect -984 24213 -932 24265
rect -916 24213 -864 24265
rect -848 24213 -796 24265
rect -780 24213 -728 24265
rect -712 24213 -660 24265
rect -644 24213 -592 24265
rect -1188 24149 -1136 24201
rect -1120 24149 -1068 24201
rect -1052 24149 -1000 24201
rect -984 24149 -932 24201
rect -916 24149 -864 24201
rect -848 24149 -796 24201
rect -780 24149 -728 24201
rect -712 24149 -660 24201
rect -644 24149 -592 24201
rect -1188 24085 -1136 24137
rect -1120 24085 -1068 24137
rect -1052 24085 -1000 24137
rect -984 24085 -932 24137
rect -916 24085 -864 24137
rect -848 24085 -796 24137
rect -780 24085 -728 24137
rect -712 24085 -660 24137
rect -644 24085 -592 24137
rect -1188 24021 -1136 24073
rect -1120 24021 -1068 24073
rect -1052 24021 -1000 24073
rect -984 24021 -932 24073
rect -916 24021 -864 24073
rect -848 24021 -796 24073
rect -780 24021 -728 24073
rect -712 24021 -660 24073
rect -644 24021 -592 24073
rect -1188 23957 -1136 24009
rect -1120 23957 -1068 24009
rect -1052 23957 -1000 24009
rect -984 23957 -932 24009
rect -916 23957 -864 24009
rect -848 23957 -796 24009
rect -780 23957 -728 24009
rect -712 23957 -660 24009
rect -644 23957 -592 24009
rect -1188 23893 -1136 23945
rect -1120 23893 -1068 23945
rect -1052 23893 -1000 23945
rect -984 23893 -932 23945
rect -916 23893 -864 23945
rect -848 23893 -796 23945
rect -780 23893 -728 23945
rect -712 23893 -660 23945
rect -644 23893 -592 23945
rect -1188 23828 -1136 23880
rect -1120 23828 -1068 23880
rect -1052 23828 -1000 23880
rect -984 23828 -932 23880
rect -916 23828 -864 23880
rect -848 23828 -796 23880
rect -780 23828 -728 23880
rect -712 23828 -660 23880
rect -644 23828 -592 23880
rect -1188 23763 -1136 23815
rect -1120 23763 -1068 23815
rect -1052 23763 -1000 23815
rect -984 23763 -932 23815
rect -916 23763 -864 23815
rect -848 23763 -796 23815
rect -780 23763 -728 23815
rect -712 23763 -660 23815
rect -644 23763 -592 23815
rect -1188 23698 -1136 23750
rect -1120 23698 -1068 23750
rect -1052 23698 -1000 23750
rect -984 23698 -932 23750
rect -916 23698 -864 23750
rect -848 23698 -796 23750
rect -780 23698 -728 23750
rect -712 23698 -660 23750
rect -644 23698 -592 23750
rect -1188 23633 -1136 23685
rect -1120 23633 -1068 23685
rect -1052 23633 -1000 23685
rect -984 23633 -932 23685
rect -916 23633 -864 23685
rect -848 23633 -796 23685
rect -780 23633 -728 23685
rect -712 23633 -660 23685
rect -644 23633 -592 23685
rect -1188 23568 -1136 23620
rect -1120 23568 -1068 23620
rect -1052 23568 -1000 23620
rect -984 23568 -932 23620
rect -916 23568 -864 23620
rect -848 23568 -796 23620
rect -780 23568 -728 23620
rect -712 23568 -660 23620
rect -644 23568 -592 23620
rect -1188 23503 -1136 23555
rect -1120 23503 -1068 23555
rect -1052 23503 -1000 23555
rect -984 23503 -932 23555
rect -916 23503 -864 23555
rect -848 23503 -796 23555
rect -780 23503 -728 23555
rect -712 23503 -660 23555
rect -644 23503 -592 23555
rect -1188 23438 -1136 23490
rect -1120 23438 -1068 23490
rect -1052 23438 -1000 23490
rect -984 23438 -932 23490
rect -916 23438 -864 23490
rect -848 23438 -796 23490
rect -780 23438 -728 23490
rect -712 23438 -660 23490
rect -644 23438 -592 23490
rect -1188 23373 -1136 23425
rect -1120 23373 -1068 23425
rect -1052 23373 -1000 23425
rect -984 23373 -932 23425
rect -916 23373 -864 23425
rect -848 23373 -796 23425
rect -780 23373 -728 23425
rect -712 23373 -660 23425
rect -644 23373 -592 23425
rect -1188 23308 -1136 23360
rect -1120 23308 -1068 23360
rect -1052 23308 -1000 23360
rect -984 23308 -932 23360
rect -916 23308 -864 23360
rect -848 23308 -796 23360
rect -780 23308 -728 23360
rect -712 23308 -660 23360
rect -644 23308 -592 23360
rect -1188 23243 -1136 23295
rect -1120 23243 -1068 23295
rect -1052 23243 -1000 23295
rect -984 23243 -932 23295
rect -916 23243 -864 23295
rect -848 23243 -796 23295
rect -780 23243 -728 23295
rect -712 23243 -660 23295
rect -644 23243 -592 23295
rect -1188 23178 -1136 23230
rect -1120 23178 -1068 23230
rect -1052 23178 -1000 23230
rect -984 23178 -932 23230
rect -916 23178 -864 23230
rect -848 23178 -796 23230
rect -780 23178 -728 23230
rect -712 23178 -660 23230
rect -644 23178 -592 23230
rect -1188 23113 -1136 23165
rect -1120 23113 -1068 23165
rect -1052 23113 -1000 23165
rect -984 23113 -932 23165
rect -916 23113 -864 23165
rect -848 23113 -796 23165
rect -780 23113 -728 23165
rect -712 23113 -660 23165
rect -644 23113 -592 23165
rect -1188 23048 -1136 23100
rect -1120 23048 -1068 23100
rect -1052 23048 -1000 23100
rect -984 23048 -932 23100
rect -916 23048 -864 23100
rect -848 23048 -796 23100
rect -780 23048 -728 23100
rect -712 23048 -660 23100
rect -644 23048 -592 23100
rect -1188 22983 -1136 23035
rect -1120 22983 -1068 23035
rect -1052 22983 -1000 23035
rect -984 22983 -932 23035
rect -916 22983 -864 23035
rect -848 22983 -796 23035
rect -780 22983 -728 23035
rect -712 22983 -660 23035
rect -644 22983 -592 23035
rect -1188 22918 -1136 22970
rect -1120 22918 -1068 22970
rect -1052 22918 -1000 22970
rect -984 22918 -932 22970
rect -916 22918 -864 22970
rect -848 22918 -796 22970
rect -780 22918 -728 22970
rect -712 22918 -660 22970
rect -644 22918 -592 22970
rect -1188 22853 -1136 22905
rect -1120 22853 -1068 22905
rect -1052 22853 -1000 22905
rect -984 22853 -932 22905
rect -916 22853 -864 22905
rect -848 22853 -796 22905
rect -780 22853 -728 22905
rect -712 22853 -660 22905
rect -644 22853 -592 22905
rect -1188 22788 -1136 22840
rect -1120 22788 -1068 22840
rect -1052 22788 -1000 22840
rect -984 22788 -932 22840
rect -916 22788 -864 22840
rect -848 22788 -796 22840
rect -780 22788 -728 22840
rect -712 22788 -660 22840
rect -644 22788 -592 22840
rect 31469 14014 31521 14066
rect 31545 14014 31597 14066
rect 31621 14014 31673 14066
rect 31469 13950 31521 14002
rect 31545 13950 31597 14002
rect 31621 13950 31673 14002
rect 31469 13886 31521 13938
rect 31545 13886 31597 13938
rect 31621 13886 31673 13938
rect 31469 13822 31521 13874
rect 31545 13822 31597 13874
rect 31621 13822 31673 13874
rect 31469 13758 31521 13810
rect 31545 13758 31597 13810
rect 31621 13758 31673 13810
rect 31469 13693 31521 13745
rect 31545 13693 31597 13745
rect 31621 13693 31673 13745
rect 31469 13628 31521 13680
rect 31545 13628 31597 13680
rect 31621 13628 31673 13680
rect 31469 13563 31521 13615
rect 31545 13563 31597 13615
rect 31621 13563 31673 13615
rect 31469 13498 31521 13550
rect 31545 13498 31597 13550
rect 31621 13498 31673 13550
rect 31469 13433 31521 13485
rect 31545 13433 31597 13485
rect 31621 13433 31673 13485
rect 31469 13368 31521 13420
rect 31545 13368 31597 13420
rect 31621 13368 31673 13420
rect 31469 13303 31521 13355
rect 31545 13303 31597 13355
rect 31621 13303 31673 13355
rect 31469 13238 31521 13290
rect 31545 13238 31597 13290
rect 31621 13238 31673 13290
rect 31469 13173 31521 13225
rect 31545 13173 31597 13225
rect 31621 13173 31673 13225
rect 31469 13108 31521 13160
rect 31545 13108 31597 13160
rect 31621 13108 31673 13160
rect 31469 13043 31521 13095
rect 31545 13043 31597 13095
rect 31621 13043 31673 13095
rect 15149 12980 15201 13032
rect 15213 12980 15265 13032
rect 15277 12980 15329 13032
rect 15341 12980 15393 13032
rect 15405 12980 15457 13032
rect 15149 12910 15201 12962
rect 15213 12910 15265 12962
rect 15277 12910 15329 12962
rect 15341 12910 15393 12962
rect 15405 12910 15457 12962
rect 15149 12840 15201 12892
rect 15213 12840 15265 12892
rect 15277 12840 15329 12892
rect 15341 12840 15393 12892
rect 15405 12840 15457 12892
rect 15149 12770 15201 12822
rect 15213 12770 15265 12822
rect 15277 12770 15329 12822
rect 15341 12770 15393 12822
rect 15405 12770 15457 12822
rect 31469 12978 31521 13030
rect 31545 12978 31597 13030
rect 31621 12978 31673 13030
rect 31469 12913 31521 12965
rect 31545 12913 31597 12965
rect 31621 12913 31673 12965
rect 31469 12848 31521 12900
rect 31545 12848 31597 12900
rect 31621 12848 31673 12900
rect 31469 12783 31521 12835
rect 31545 12783 31597 12835
rect 31621 12783 31673 12835
rect 31469 12718 31521 12770
rect 31545 12718 31597 12770
rect 31621 12718 31673 12770
rect 31469 12653 31521 12705
rect 31545 12653 31597 12705
rect 31621 12653 31673 12705
rect 31469 12588 31521 12640
rect 31545 12588 31597 12640
rect 31621 12588 31673 12640
rect 31469 12523 31521 12575
rect 31545 12523 31597 12575
rect 31621 12523 31673 12575
rect 31469 12458 31521 12510
rect 31545 12458 31597 12510
rect 31621 12458 31673 12510
rect 31469 12393 31521 12445
rect 31545 12393 31597 12445
rect 31621 12393 31673 12445
rect 31469 12328 31521 12380
rect 31545 12328 31597 12380
rect 31621 12328 31673 12380
rect 31469 12263 31521 12315
rect 31545 12263 31597 12315
rect 31621 12263 31673 12315
rect 31469 12198 31521 12250
rect 31545 12198 31597 12250
rect 31621 12198 31673 12250
rect 31469 12133 31521 12185
rect 31545 12133 31597 12185
rect 31621 12133 31673 12185
rect 31469 12068 31521 12120
rect 31545 12068 31597 12120
rect 31621 12068 31673 12120
rect 17617 11985 17669 12037
rect 17685 11985 17737 12037
rect 17752 11985 17804 12037
rect 17819 11985 17871 12037
rect 17886 11985 17938 12037
rect 17953 11985 18005 12037
rect 18020 11985 18072 12037
rect 18087 11985 18139 12037
rect 18154 11985 18206 12037
rect 18221 11985 18273 12037
rect 18288 11985 18340 12037
rect 18355 11985 18407 12037
rect 17617 11913 17669 11965
rect 17685 11913 17737 11965
rect 17752 11913 17804 11965
rect 17819 11913 17871 11965
rect 17886 11913 17938 11965
rect 17953 11913 18005 11965
rect 18020 11913 18072 11965
rect 18087 11913 18139 11965
rect 18154 11913 18206 11965
rect 18221 11913 18273 11965
rect 18288 11913 18340 11965
rect 18355 11913 18407 11965
rect 17617 11841 17669 11893
rect 17685 11841 17737 11893
rect 17752 11841 17804 11893
rect 17819 11841 17871 11893
rect 17886 11841 17938 11893
rect 17953 11841 18005 11893
rect 18020 11841 18072 11893
rect 18087 11841 18139 11893
rect 18154 11841 18206 11893
rect 18221 11841 18273 11893
rect 18288 11841 18340 11893
rect 18355 11841 18407 11893
rect 17617 11769 17669 11821
rect 17685 11769 17737 11821
rect 17752 11769 17804 11821
rect 17819 11769 17871 11821
rect 17886 11769 17938 11821
rect 17953 11769 18005 11821
rect 18020 11769 18072 11821
rect 18087 11769 18139 11821
rect 18154 11769 18206 11821
rect 18221 11769 18273 11821
rect 18288 11769 18340 11821
rect 18355 11769 18407 11821
rect 31469 12003 31521 12055
rect 31545 12003 31597 12055
rect 31621 12003 31673 12055
rect 31469 11938 31521 11990
rect 31545 11938 31597 11990
rect 31621 11938 31673 11990
rect 31469 11873 31521 11925
rect 31545 11873 31597 11925
rect 31621 11873 31673 11925
rect 31469 11808 31521 11860
rect 31545 11808 31597 11860
rect 31621 11808 31673 11860
rect 31469 11743 31521 11795
rect 31545 11743 31597 11795
rect 31621 11743 31673 11795
rect 4079 11653 4131 11705
rect 4143 11653 4195 11705
rect 5115 11653 5167 11705
rect 5179 11653 5231 11705
rect 31469 11678 31521 11730
rect 31545 11678 31597 11730
rect 31621 11678 31673 11730
rect 31469 11613 31521 11665
rect 31545 11613 31597 11665
rect 31621 11613 31673 11665
rect 19836 11530 19888 11582
rect 19908 11530 19960 11582
rect 19979 11530 20031 11582
rect 20050 11530 20102 11582
rect 20121 11530 20173 11582
rect 20192 11530 20244 11582
rect 20263 11530 20315 11582
rect 19836 11462 19888 11514
rect 19908 11462 19960 11514
rect 19979 11462 20031 11514
rect 20050 11462 20102 11514
rect 20121 11462 20173 11514
rect 20192 11462 20244 11514
rect 20263 11462 20315 11514
rect 19836 11394 19888 11446
rect 19908 11394 19960 11446
rect 19979 11394 20031 11446
rect 20050 11394 20102 11446
rect 20121 11394 20173 11446
rect 20192 11394 20244 11446
rect 20263 11394 20315 11446
rect 19836 11326 19888 11378
rect 19908 11326 19960 11378
rect 19979 11326 20031 11378
rect 20050 11326 20102 11378
rect 20121 11326 20173 11378
rect 20192 11326 20244 11378
rect 20263 11326 20315 11378
rect 31469 11548 31521 11600
rect 31545 11548 31597 11600
rect 31621 11548 31673 11600
rect 31469 11483 31521 11535
rect 31545 11483 31597 11535
rect 31621 11483 31673 11535
rect 31469 11418 31521 11470
rect 31545 11418 31597 11470
rect 31621 11418 31673 11470
rect 31469 11353 31521 11405
rect 31545 11353 31597 11405
rect 31621 11353 31673 11405
rect 13890 11265 13942 11274
rect 13981 11265 14033 11274
rect 14071 11265 14123 11274
rect 14424 11265 14476 11274
rect 14489 11265 14541 11274
rect 14553 11265 14605 11274
rect 13890 11231 13921 11265
rect 13921 11231 13942 11265
rect 13981 11231 13994 11265
rect 13994 11231 14033 11265
rect 14071 11231 14106 11265
rect 14106 11231 14123 11265
rect 14424 11231 14432 11265
rect 14432 11231 14471 11265
rect 14471 11231 14476 11265
rect 14489 11231 14505 11265
rect 14505 11231 14541 11265
rect 14553 11231 14578 11265
rect 14578 11231 14605 11265
rect 13890 11222 13942 11231
rect 13981 11222 14033 11231
rect 14071 11222 14123 11231
rect 14424 11222 14476 11231
rect 14489 11222 14541 11231
rect 14553 11222 14605 11231
rect 14617 11265 14669 11274
rect 14617 11231 14651 11265
rect 14651 11231 14669 11265
rect 14617 11222 14669 11231
rect 14681 11265 14733 11274
rect 14681 11231 14690 11265
rect 14690 11231 14724 11265
rect 14724 11231 14733 11265
rect 14681 11222 14733 11231
rect 31469 11288 31521 11340
rect 31545 11288 31597 11340
rect 31621 11288 31673 11340
rect 31469 11223 31521 11275
rect 31545 11223 31597 11275
rect 31621 11223 31673 11275
rect 31469 11158 31521 11210
rect 31545 11158 31597 11210
rect 31621 11158 31673 11210
rect 4085 11090 4137 11142
rect 4149 11090 4201 11142
rect 31469 11093 31521 11145
rect 31545 11093 31597 11145
rect 31621 11093 31673 11145
rect 13890 10542 13942 10551
rect 13981 10542 14033 10551
rect 14071 10542 14123 10551
rect 14424 10542 14476 10551
rect 14489 10542 14541 10551
rect 14553 10542 14605 10551
rect 14617 10542 14669 10551
rect 14681 10542 14733 10551
rect 13890 10508 13930 10542
rect 13930 10508 13942 10542
rect 13981 10508 14004 10542
rect 14004 10508 14033 10542
rect 14071 10508 14078 10542
rect 14078 10508 14112 10542
rect 14112 10508 14123 10542
rect 14424 10508 14448 10542
rect 14448 10508 14476 10542
rect 14489 10508 14522 10542
rect 14522 10508 14541 10542
rect 14553 10508 14556 10542
rect 14556 10508 14596 10542
rect 14596 10508 14605 10542
rect 14617 10508 14630 10542
rect 14630 10508 14669 10542
rect 14681 10508 14704 10542
rect 14704 10508 14733 10542
rect 13890 10499 13942 10508
rect 13981 10499 14033 10508
rect 14071 10499 14123 10508
rect 14424 10499 14476 10508
rect 14489 10499 14541 10508
rect 14553 10499 14605 10508
rect 14617 10499 14669 10508
rect 14681 10499 14733 10508
rect 6025 9871 6077 9923
rect 6089 9871 6141 9923
rect 5623 9169 5675 9221
rect 6123 9195 6175 9247
rect 6187 9195 6239 9247
rect 10054 9195 10106 9247
rect 10118 9195 10170 9247
rect 10785 9204 10837 9256
rect 10849 9204 10901 9256
rect 5623 9105 5675 9157
rect 18537 8371 18589 8423
rect 18601 8371 18653 8423
rect 18665 8371 18717 8423
rect 18729 8371 18781 8423
rect 18793 8371 18845 8423
rect 18857 8371 18909 8423
rect 5298 7436 5350 7488
rect 6123 7429 6175 7481
rect 6187 7429 6239 7481
rect 5298 7372 5350 7424
rect 13259 7327 13311 7379
rect 13323 7327 13375 7379
rect -587 7009 -535 7061
rect -505 7009 -453 7061
rect -423 7009 -371 7061
rect -341 7009 -289 7061
rect -259 7009 -207 7061
rect -587 6945 -535 6997
rect -505 6945 -453 6997
rect -423 6945 -371 6997
rect -341 6945 -289 6997
rect -259 6945 -207 6997
rect 23958 6302 24010 6354
rect 24042 6302 24094 6354
rect 24126 6302 24178 6354
rect 24209 6302 24261 6354
rect 23958 6236 24010 6288
rect 24042 6236 24094 6288
rect 24126 6236 24178 6288
rect 24209 6236 24261 6288
rect 23958 6170 24010 6222
rect 24042 6170 24094 6222
rect 24126 6170 24178 6222
rect 24209 6170 24261 6222
rect 76 5648 192 5764
rect 2145 5647 2261 5763
rect -594 4764 -542 4816
rect -510 4764 -458 4816
rect -426 4764 -374 4816
rect -342 4764 -290 4816
rect -258 4764 -206 4816
rect 4847 3200 4899 3252
rect 4847 3136 4899 3188
rect 5987 2484 6039 2536
rect 6051 2484 6103 2536
rect 5987 2415 6039 2467
rect 6051 2415 6103 2467
rect 5987 2346 6039 2398
rect 6051 2346 6103 2398
rect 5994 2153 6046 2205
rect 6069 2153 6121 2205
rect 519 1323 635 1503
rect 1234 1323 1350 1503
rect 1861 1323 1977 1503
rect 2573 1323 2689 1503
rect 5987 1653 6039 1705
rect 6051 1653 6103 1705
rect 5987 1573 6039 1625
rect 6051 1573 6103 1625
rect 8549 1688 8601 1740
rect 8613 1688 8665 1740
rect 8677 1688 8729 1740
rect 8549 1619 8601 1671
rect 8613 1619 8665 1671
rect 8677 1619 8729 1671
rect 8549 1550 8601 1602
rect 8613 1550 8665 1602
rect 8677 1550 8729 1602
<< metal2 >>
rect -2519 43689 1083 43695
rect -2519 43637 -2502 43689
rect -2450 43637 -2438 43689
rect -2386 43637 -2374 43689
rect -2322 43637 -2310 43689
rect -2258 43637 -2246 43689
rect -2194 43637 -2182 43689
rect -2130 43637 -2118 43689
rect -2066 43637 -2054 43689
rect -2002 43637 -1990 43689
rect -1938 43637 -1926 43689
rect -1874 43637 -1862 43689
rect -1810 43637 -1798 43689
rect -1746 43637 -1734 43689
rect -1682 43637 -1670 43689
rect -1618 43637 -1606 43689
rect -1554 43637 -1542 43689
rect -1490 43637 -1478 43689
rect -1426 43637 -1414 43689
rect -1362 43637 -1350 43689
rect -1298 43637 -1286 43689
rect -1234 43637 -1222 43689
rect -1170 43637 -1158 43689
rect -1106 43637 -1094 43689
rect -1042 43637 -1030 43689
rect -978 43637 -966 43689
rect -914 43637 -902 43689
rect -850 43637 -838 43689
rect -786 43637 -774 43689
rect -722 43637 -710 43689
rect -658 43637 646 43689
rect 698 43637 710 43689
rect 762 43637 774 43689
rect 826 43637 838 43689
rect 890 43637 902 43689
rect 954 43637 966 43689
rect 1018 43637 1030 43689
rect 1082 43637 1083 43689
rect -2519 43623 1083 43637
rect -2519 43571 -2502 43623
rect -2450 43571 -2438 43623
rect -2386 43571 -2374 43623
rect -2322 43571 -2310 43623
rect -2258 43571 -2246 43623
rect -2194 43571 -2182 43623
rect -2130 43571 -2118 43623
rect -2066 43571 -2054 43623
rect -2002 43571 -1990 43623
rect -1938 43571 -1926 43623
rect -1874 43571 -1862 43623
rect -1810 43571 -1798 43623
rect -1746 43571 -1734 43623
rect -1682 43571 -1670 43623
rect -1618 43571 -1606 43623
rect -1554 43571 -1542 43623
rect -1490 43571 -1478 43623
rect -1426 43571 -1414 43623
rect -1362 43571 -1350 43623
rect -1298 43571 -1286 43623
rect -1234 43571 -1222 43623
rect -1170 43571 -1158 43623
rect -1106 43571 -1094 43623
rect -1042 43571 -1030 43623
rect -978 43571 -966 43623
rect -914 43571 -902 43623
rect -850 43571 -838 43623
rect -786 43571 -774 43623
rect -722 43571 -710 43623
rect -658 43571 646 43623
rect 698 43571 710 43623
rect 762 43571 774 43623
rect 826 43571 838 43623
rect 890 43571 902 43623
rect 954 43571 966 43623
rect 1018 43571 1030 43623
rect 1082 43571 1083 43623
rect -2519 43557 1083 43571
rect -2519 43505 -2502 43557
rect -2450 43505 -2438 43557
rect -2386 43505 -2374 43557
rect -2322 43505 -2310 43557
rect -2258 43505 -2246 43557
rect -2194 43505 -2182 43557
rect -2130 43505 -2118 43557
rect -2066 43505 -2054 43557
rect -2002 43505 -1990 43557
rect -1938 43505 -1926 43557
rect -1874 43505 -1862 43557
rect -1810 43505 -1798 43557
rect -1746 43505 -1734 43557
rect -1682 43505 -1670 43557
rect -1618 43505 -1606 43557
rect -1554 43505 -1542 43557
rect -1490 43505 -1478 43557
rect -1426 43505 -1414 43557
rect -1362 43505 -1350 43557
rect -1298 43505 -1286 43557
rect -1234 43505 -1222 43557
rect -1170 43505 -1158 43557
rect -1106 43505 -1094 43557
rect -1042 43505 -1030 43557
rect -978 43505 -966 43557
rect -914 43505 -902 43557
rect -850 43505 -838 43557
rect -786 43505 -774 43557
rect -722 43505 -710 43557
rect -658 43505 646 43557
rect 698 43505 710 43557
rect 762 43505 774 43557
rect 826 43505 838 43557
rect 890 43505 902 43557
rect 954 43505 966 43557
rect 1018 43505 1030 43557
rect 1082 43505 1083 43557
rect -2519 43491 1083 43505
rect -2519 43439 -2502 43491
rect -2450 43439 -2438 43491
rect -2386 43439 -2374 43491
rect -2322 43439 -2310 43491
rect -2258 43439 -2246 43491
rect -2194 43439 -2182 43491
rect -2130 43439 -2118 43491
rect -2066 43439 -2054 43491
rect -2002 43439 -1990 43491
rect -1938 43439 -1926 43491
rect -1874 43439 -1862 43491
rect -1810 43439 -1798 43491
rect -1746 43439 -1734 43491
rect -1682 43439 -1670 43491
rect -1618 43439 -1606 43491
rect -1554 43439 -1542 43491
rect -1490 43439 -1478 43491
rect -1426 43439 -1414 43491
rect -1362 43439 -1350 43491
rect -1298 43439 -1286 43491
rect -1234 43439 -1222 43491
rect -1170 43439 -1158 43491
rect -1106 43439 -1094 43491
rect -1042 43439 -1030 43491
rect -978 43439 -966 43491
rect -914 43439 -902 43491
rect -850 43439 -838 43491
rect -786 43439 -774 43491
rect -722 43439 -710 43491
rect -658 43439 646 43491
rect 698 43439 710 43491
rect 762 43439 774 43491
rect 826 43439 838 43491
rect 890 43439 902 43491
rect 954 43439 966 43491
rect 1018 43439 1030 43491
rect 1082 43439 1083 43491
rect -2519 43425 1083 43439
rect -2519 43373 -2502 43425
rect -2450 43373 -2438 43425
rect -2386 43373 -2374 43425
rect -2322 43373 -2310 43425
rect -2258 43373 -2246 43425
rect -2194 43373 -2182 43425
rect -2130 43373 -2118 43425
rect -2066 43373 -2054 43425
rect -2002 43373 -1990 43425
rect -1938 43373 -1926 43425
rect -1874 43373 -1862 43425
rect -1810 43373 -1798 43425
rect -1746 43373 -1734 43425
rect -1682 43373 -1670 43425
rect -1618 43373 -1606 43425
rect -1554 43373 -1542 43425
rect -1490 43373 -1478 43425
rect -1426 43373 -1414 43425
rect -1362 43373 -1350 43425
rect -1298 43373 -1286 43425
rect -1234 43373 -1222 43425
rect -1170 43373 -1158 43425
rect -1106 43373 -1094 43425
rect -1042 43373 -1030 43425
rect -978 43373 -966 43425
rect -914 43373 -902 43425
rect -850 43373 -838 43425
rect -786 43373 -774 43425
rect -722 43373 -710 43425
rect -658 43373 646 43425
rect 698 43373 710 43425
rect 762 43373 774 43425
rect 826 43373 838 43425
rect 890 43373 902 43425
rect 954 43373 966 43425
rect 1018 43373 1030 43425
rect 1082 43373 1083 43425
rect -2519 43359 1083 43373
rect -2519 43307 -2502 43359
rect -2450 43307 -2438 43359
rect -2386 43307 -2374 43359
rect -2322 43307 -2310 43359
rect -2258 43307 -2246 43359
rect -2194 43307 -2182 43359
rect -2130 43307 -2118 43359
rect -2066 43307 -2054 43359
rect -2002 43307 -1990 43359
rect -1938 43307 -1926 43359
rect -1874 43307 -1862 43359
rect -1810 43307 -1798 43359
rect -1746 43307 -1734 43359
rect -1682 43307 -1670 43359
rect -1618 43307 -1606 43359
rect -1554 43307 -1542 43359
rect -1490 43307 -1478 43359
rect -1426 43307 -1414 43359
rect -1362 43307 -1350 43359
rect -1298 43307 -1286 43359
rect -1234 43307 -1222 43359
rect -1170 43307 -1158 43359
rect -1106 43307 -1094 43359
rect -1042 43307 -1030 43359
rect -978 43307 -966 43359
rect -914 43307 -902 43359
rect -850 43307 -838 43359
rect -786 43307 -774 43359
rect -722 43307 -710 43359
rect -658 43307 646 43359
rect 698 43307 710 43359
rect 762 43307 774 43359
rect 826 43307 838 43359
rect 890 43307 902 43359
rect 954 43307 966 43359
rect 1018 43307 1030 43359
rect 1082 43307 1083 43359
rect -2519 43293 1083 43307
rect -2519 43241 -2502 43293
rect -2450 43241 -2438 43293
rect -2386 43241 -2374 43293
rect -2322 43241 -2310 43293
rect -2258 43241 -2246 43293
rect -2194 43241 -2182 43293
rect -2130 43241 -2118 43293
rect -2066 43241 -2054 43293
rect -2002 43241 -1990 43293
rect -1938 43241 -1926 43293
rect -1874 43241 -1862 43293
rect -1810 43241 -1798 43293
rect -1746 43241 -1734 43293
rect -1682 43241 -1670 43293
rect -1618 43241 -1606 43293
rect -1554 43241 -1542 43293
rect -1490 43241 -1478 43293
rect -1426 43241 -1414 43293
rect -1362 43241 -1350 43293
rect -1298 43241 -1286 43293
rect -1234 43241 -1222 43293
rect -1170 43241 -1158 43293
rect -1106 43241 -1094 43293
rect -1042 43241 -1030 43293
rect -978 43241 -966 43293
rect -914 43241 -902 43293
rect -850 43241 -838 43293
rect -786 43241 -774 43293
rect -722 43241 -710 43293
rect -658 43241 646 43293
rect 698 43241 710 43293
rect 762 43241 774 43293
rect 826 43241 838 43293
rect 890 43241 902 43293
rect 954 43241 966 43293
rect 1018 43241 1030 43293
rect 1082 43241 1083 43293
rect -2519 43226 1083 43241
rect -2519 43174 -2502 43226
rect -2450 43174 -2438 43226
rect -2386 43174 -2374 43226
rect -2322 43174 -2310 43226
rect -2258 43174 -2246 43226
rect -2194 43174 -2182 43226
rect -2130 43174 -2118 43226
rect -2066 43174 -2054 43226
rect -2002 43174 -1990 43226
rect -1938 43174 -1926 43226
rect -1874 43174 -1862 43226
rect -1810 43174 -1798 43226
rect -1746 43174 -1734 43226
rect -1682 43174 -1670 43226
rect -1618 43174 -1606 43226
rect -1554 43174 -1542 43226
rect -1490 43174 -1478 43226
rect -1426 43174 -1414 43226
rect -1362 43174 -1350 43226
rect -1298 43174 -1286 43226
rect -1234 43174 -1222 43226
rect -1170 43174 -1158 43226
rect -1106 43174 -1094 43226
rect -1042 43174 -1030 43226
rect -978 43174 -966 43226
rect -914 43174 -902 43226
rect -850 43174 -838 43226
rect -786 43174 -774 43226
rect -722 43174 -710 43226
rect -658 43174 646 43226
rect 698 43174 710 43226
rect 762 43174 774 43226
rect 826 43174 838 43226
rect 890 43174 902 43226
rect 954 43174 966 43226
rect 1018 43174 1030 43226
rect 1082 43174 1083 43226
rect -2519 43168 1083 43174
tri 1702 40810 2123 41231 se
rect 2123 40810 2389 41231
rect 1702 40707 2389 40810
rect 1702 40257 2028 40707
tri 2028 40563 2172 40707 nw
rect 31407 40072 31413 40188
rect 31529 40072 31535 40188
rect 31407 32050 31535 40072
rect 31593 39827 31599 39943
rect 31715 39827 31721 39943
rect 31593 32050 31721 39827
rect -1190 25161 -590 26406
rect -1190 25109 -1188 25161
rect -1136 25109 -1120 25161
rect -1068 25109 -1052 25161
rect -1000 25109 -984 25161
rect -932 25109 -916 25161
rect -864 25109 -848 25161
rect -796 25109 -780 25161
rect -728 25109 -712 25161
rect -660 25109 -644 25161
rect -592 25109 -590 25161
rect -1190 25097 -590 25109
rect -1190 25045 -1188 25097
rect -1136 25045 -1120 25097
rect -1068 25045 -1052 25097
rect -1000 25045 -984 25097
rect -932 25045 -916 25097
rect -864 25045 -848 25097
rect -796 25045 -780 25097
rect -728 25045 -712 25097
rect -660 25045 -644 25097
rect -592 25045 -590 25097
rect -1190 25033 -590 25045
rect -1190 24981 -1188 25033
rect -1136 24981 -1120 25033
rect -1068 24981 -1052 25033
rect -1000 24981 -984 25033
rect -932 24981 -916 25033
rect -864 24981 -848 25033
rect -796 24981 -780 25033
rect -728 24981 -712 25033
rect -660 24981 -644 25033
rect -592 24981 -590 25033
rect 14796 25012 14850 25111
rect -1190 24969 -590 24981
rect -1190 24917 -1188 24969
rect -1136 24917 -1120 24969
rect -1068 24917 -1052 24969
rect -1000 24917 -984 24969
rect -932 24917 -916 24969
rect -864 24917 -848 24969
rect -796 24917 -780 24969
rect -728 24917 -712 24969
rect -660 24917 -644 24969
rect -592 24917 -590 24969
rect -1190 24905 -590 24917
rect -1190 24853 -1188 24905
rect -1136 24853 -1120 24905
rect -1068 24853 -1052 24905
rect -1000 24853 -984 24905
rect -932 24853 -916 24905
rect -864 24853 -848 24905
rect -796 24853 -780 24905
rect -728 24853 -712 24905
rect -660 24853 -644 24905
rect -592 24853 -590 24905
rect -1190 24841 -590 24853
rect -1190 24789 -1188 24841
rect -1136 24789 -1120 24841
rect -1068 24789 -1052 24841
rect -1000 24789 -984 24841
rect -932 24789 -916 24841
rect -864 24789 -848 24841
rect -796 24789 -780 24841
rect -728 24789 -712 24841
rect -660 24789 -644 24841
rect -592 24789 -590 24841
rect -1190 24777 -590 24789
rect -1190 24725 -1188 24777
rect -1136 24725 -1120 24777
rect -1068 24725 -1052 24777
rect -1000 24725 -984 24777
rect -932 24725 -916 24777
rect -864 24725 -848 24777
rect -796 24725 -780 24777
rect -728 24725 -712 24777
rect -660 24725 -644 24777
rect -592 24725 -590 24777
rect -1190 24713 -590 24725
rect -1190 24661 -1188 24713
rect -1136 24661 -1120 24713
rect -1068 24661 -1052 24713
rect -1000 24661 -984 24713
rect -932 24661 -916 24713
rect -864 24661 -848 24713
rect -796 24661 -780 24713
rect -728 24661 -712 24713
rect -660 24661 -644 24713
rect -592 24661 -590 24713
rect -1190 24649 -590 24661
rect -1190 24597 -1188 24649
rect -1136 24597 -1120 24649
rect -1068 24597 -1052 24649
rect -1000 24597 -984 24649
rect -932 24597 -916 24649
rect -864 24597 -848 24649
rect -796 24597 -780 24649
rect -728 24597 -712 24649
rect -660 24597 -644 24649
rect -592 24597 -590 24649
rect -1190 24585 -590 24597
rect -1190 24533 -1188 24585
rect -1136 24533 -1120 24585
rect -1068 24533 -1052 24585
rect -1000 24533 -984 24585
rect -932 24533 -916 24585
rect -864 24533 -848 24585
rect -796 24533 -780 24585
rect -728 24533 -712 24585
rect -660 24533 -644 24585
rect -592 24533 -590 24585
rect -1190 24521 -590 24533
rect -1190 24469 -1188 24521
rect -1136 24469 -1120 24521
rect -1068 24469 -1052 24521
rect -1000 24469 -984 24521
rect -932 24469 -916 24521
rect -864 24469 -848 24521
rect -796 24469 -780 24521
rect -728 24469 -712 24521
rect -660 24469 -644 24521
rect -592 24469 -590 24521
rect -1190 24457 -590 24469
rect -1190 24405 -1188 24457
rect -1136 24405 -1120 24457
rect -1068 24405 -1052 24457
rect -1000 24405 -984 24457
rect -932 24405 -916 24457
rect -864 24405 -848 24457
rect -796 24405 -780 24457
rect -728 24405 -712 24457
rect -660 24405 -644 24457
rect -592 24405 -590 24457
rect -1190 24393 -590 24405
rect -1190 24341 -1188 24393
rect -1136 24341 -1120 24393
rect -1068 24341 -1052 24393
rect -1000 24341 -984 24393
rect -932 24341 -916 24393
rect -864 24341 -848 24393
rect -796 24341 -780 24393
rect -728 24341 -712 24393
rect -660 24341 -644 24393
rect -592 24341 -590 24393
rect -1190 24329 -590 24341
rect -1190 24277 -1188 24329
rect -1136 24277 -1120 24329
rect -1068 24277 -1052 24329
rect -1000 24277 -984 24329
rect -932 24277 -916 24329
rect -864 24277 -848 24329
rect -796 24277 -780 24329
rect -728 24277 -712 24329
rect -660 24277 -644 24329
rect -592 24277 -590 24329
rect -1190 24265 -590 24277
rect -1190 24213 -1188 24265
rect -1136 24213 -1120 24265
rect -1068 24213 -1052 24265
rect -1000 24213 -984 24265
rect -932 24213 -916 24265
rect -864 24213 -848 24265
rect -796 24213 -780 24265
rect -728 24213 -712 24265
rect -660 24213 -644 24265
rect -592 24213 -590 24265
rect -1190 24201 -590 24213
rect -1190 24149 -1188 24201
rect -1136 24149 -1120 24201
rect -1068 24149 -1052 24201
rect -1000 24149 -984 24201
rect -932 24149 -916 24201
rect -864 24149 -848 24201
rect -796 24149 -780 24201
rect -728 24149 -712 24201
rect -660 24149 -644 24201
rect -592 24149 -590 24201
rect -1190 24137 -590 24149
rect -1190 24085 -1188 24137
rect -1136 24085 -1120 24137
rect -1068 24085 -1052 24137
rect -1000 24085 -984 24137
rect -932 24085 -916 24137
rect -864 24085 -848 24137
rect -796 24085 -780 24137
rect -728 24085 -712 24137
rect -660 24085 -644 24137
rect -592 24085 -590 24137
rect -1190 24073 -590 24085
rect -1190 24021 -1188 24073
rect -1136 24021 -1120 24073
rect -1068 24021 -1052 24073
rect -1000 24021 -984 24073
rect -932 24021 -916 24073
rect -864 24021 -848 24073
rect -796 24021 -780 24073
rect -728 24021 -712 24073
rect -660 24021 -644 24073
rect -592 24021 -590 24073
rect -1190 24009 -590 24021
rect -1190 23957 -1188 24009
rect -1136 23957 -1120 24009
rect -1068 23957 -1052 24009
rect -1000 23957 -984 24009
rect -932 23957 -916 24009
rect -864 23957 -848 24009
rect -796 23957 -780 24009
rect -728 23957 -712 24009
rect -660 23957 -644 24009
rect -592 23957 -590 24009
rect -1190 23945 -590 23957
rect -1190 23893 -1188 23945
rect -1136 23893 -1120 23945
rect -1068 23893 -1052 23945
rect -1000 23893 -984 23945
rect -932 23893 -916 23945
rect -864 23893 -848 23945
rect -796 23893 -780 23945
rect -728 23893 -712 23945
rect -660 23893 -644 23945
rect -592 23893 -590 23945
rect -1190 23880 -590 23893
rect -1190 23828 -1188 23880
rect -1136 23828 -1120 23880
rect -1068 23828 -1052 23880
rect -1000 23828 -984 23880
rect -932 23828 -916 23880
rect -864 23828 -848 23880
rect -796 23828 -780 23880
rect -728 23828 -712 23880
rect -660 23828 -644 23880
rect -592 23828 -590 23880
rect -1190 23815 -590 23828
rect -1190 23763 -1188 23815
rect -1136 23763 -1120 23815
rect -1068 23763 -1052 23815
rect -1000 23763 -984 23815
rect -932 23763 -916 23815
rect -864 23763 -848 23815
rect -796 23763 -780 23815
rect -728 23763 -712 23815
rect -660 23763 -644 23815
rect -592 23763 -590 23815
rect -1190 23750 -590 23763
rect -1190 23698 -1188 23750
rect -1136 23698 -1120 23750
rect -1068 23698 -1052 23750
rect -1000 23698 -984 23750
rect -932 23698 -916 23750
rect -864 23698 -848 23750
rect -796 23698 -780 23750
rect -728 23698 -712 23750
rect -660 23698 -644 23750
rect -592 23698 -590 23750
rect -1190 23685 -590 23698
rect -1190 23633 -1188 23685
rect -1136 23633 -1120 23685
rect -1068 23633 -1052 23685
rect -1000 23633 -984 23685
rect -932 23633 -916 23685
rect -864 23633 -848 23685
rect -796 23633 -780 23685
rect -728 23633 -712 23685
rect -660 23633 -644 23685
rect -592 23633 -590 23685
rect -1190 23620 -590 23633
rect -1190 23568 -1188 23620
rect -1136 23568 -1120 23620
rect -1068 23568 -1052 23620
rect -1000 23568 -984 23620
rect -932 23568 -916 23620
rect -864 23568 -848 23620
rect -796 23568 -780 23620
rect -728 23568 -712 23620
rect -660 23568 -644 23620
rect -592 23568 -590 23620
rect -1190 23555 -590 23568
rect -1190 23503 -1188 23555
rect -1136 23503 -1120 23555
rect -1068 23503 -1052 23555
rect -1000 23503 -984 23555
rect -932 23503 -916 23555
rect -864 23503 -848 23555
rect -796 23503 -780 23555
rect -728 23503 -712 23555
rect -660 23503 -644 23555
rect -592 23503 -590 23555
rect -1190 23490 -590 23503
rect -1190 23438 -1188 23490
rect -1136 23438 -1120 23490
rect -1068 23438 -1052 23490
rect -1000 23438 -984 23490
rect -932 23438 -916 23490
rect -864 23438 -848 23490
rect -796 23438 -780 23490
rect -728 23438 -712 23490
rect -660 23438 -644 23490
rect -592 23438 -590 23490
rect -1190 23425 -590 23438
rect -1190 23373 -1188 23425
rect -1136 23373 -1120 23425
rect -1068 23373 -1052 23425
rect -1000 23373 -984 23425
rect -932 23373 -916 23425
rect -864 23373 -848 23425
rect -796 23373 -780 23425
rect -728 23373 -712 23425
rect -660 23373 -644 23425
rect -592 23373 -590 23425
rect -1190 23360 -590 23373
rect -1190 23308 -1188 23360
rect -1136 23308 -1120 23360
rect -1068 23308 -1052 23360
rect -1000 23308 -984 23360
rect -932 23308 -916 23360
rect -864 23308 -848 23360
rect -796 23308 -780 23360
rect -728 23308 -712 23360
rect -660 23308 -644 23360
rect -592 23308 -590 23360
rect -1190 23295 -590 23308
rect -1190 23243 -1188 23295
rect -1136 23243 -1120 23295
rect -1068 23243 -1052 23295
rect -1000 23243 -984 23295
rect -932 23243 -916 23295
rect -864 23243 -848 23295
rect -796 23243 -780 23295
rect -728 23243 -712 23295
rect -660 23243 -644 23295
rect -592 23243 -590 23295
rect -1190 23230 -590 23243
rect -1190 23178 -1188 23230
rect -1136 23178 -1120 23230
rect -1068 23178 -1052 23230
rect -1000 23178 -984 23230
rect -932 23178 -916 23230
rect -864 23178 -848 23230
rect -796 23178 -780 23230
rect -728 23178 -712 23230
rect -660 23178 -644 23230
rect -592 23178 -590 23230
rect -1190 23165 -590 23178
rect -1190 23113 -1188 23165
rect -1136 23113 -1120 23165
rect -1068 23113 -1052 23165
rect -1000 23113 -984 23165
rect -932 23113 -916 23165
rect -864 23113 -848 23165
rect -796 23113 -780 23165
rect -728 23113 -712 23165
rect -660 23113 -644 23165
rect -592 23113 -590 23165
rect -1190 23100 -590 23113
rect -1190 23048 -1188 23100
rect -1136 23048 -1120 23100
rect -1068 23048 -1052 23100
rect -1000 23048 -984 23100
rect -932 23048 -916 23100
rect -864 23048 -848 23100
rect -796 23048 -780 23100
rect -728 23048 -712 23100
rect -660 23048 -644 23100
rect -592 23048 -590 23100
rect -1190 23035 -590 23048
rect -1190 22983 -1188 23035
rect -1136 22983 -1120 23035
rect -1068 22983 -1052 23035
rect -1000 22983 -984 23035
rect -932 22983 -916 23035
rect -864 22983 -848 23035
rect -796 22983 -780 23035
rect -728 22983 -712 23035
rect -660 22983 -644 23035
rect -592 22983 -590 23035
rect -1190 22970 -590 22983
rect -1190 22918 -1188 22970
rect -1136 22918 -1120 22970
rect -1068 22918 -1052 22970
rect -1000 22918 -984 22970
rect -932 22918 -916 22970
rect -864 22918 -848 22970
rect -796 22918 -780 22970
rect -728 22918 -712 22970
rect -660 22918 -644 22970
rect -592 22918 -590 22970
rect -1190 22905 -590 22918
rect -1190 22853 -1188 22905
rect -1136 22853 -1120 22905
rect -1068 22853 -1052 22905
rect -1000 22853 -984 22905
rect -932 22853 -916 22905
rect -864 22853 -848 22905
rect -796 22853 -780 22905
rect -728 22853 -712 22905
rect -660 22853 -644 22905
rect -592 22853 -590 22905
rect -1190 22840 -590 22853
rect -1190 22788 -1188 22840
rect -1136 22788 -1120 22840
rect -1068 22788 -1052 22840
rect -1000 22788 -984 22840
rect -932 22788 -916 22840
rect -864 22788 -848 22840
rect -796 22788 -780 22840
rect -728 22788 -712 22840
rect -660 22788 -644 22840
rect -592 22788 -590 22840
rect -1190 21856 -590 22788
tri -590 21856 -426 22020 sw
rect -1190 21677 -426 21856
tri -1190 21439 -952 21677 ne
rect -952 17351 -426 21677
tri -426 17351 -201 17576 sw
rect -952 17243 -201 17351
tri -952 16884 -593 17243 ne
rect -593 7061 -201 17243
rect 31468 14066 31674 14072
rect 31468 14014 31469 14066
rect 31521 14014 31545 14066
rect 31597 14014 31621 14066
rect 31673 14014 31674 14066
rect 31468 14002 31674 14014
rect 31468 13950 31469 14002
rect 31521 13950 31545 14002
rect 31597 13950 31621 14002
rect 31673 13950 31674 14002
rect 31468 13938 31674 13950
rect 31468 13886 31469 13938
rect 31521 13886 31545 13938
rect 31597 13886 31621 13938
rect 31673 13886 31674 13938
rect 31468 13874 31674 13886
rect 31468 13822 31469 13874
rect 31521 13822 31545 13874
rect 31597 13822 31621 13874
rect 31673 13822 31674 13874
rect 31468 13810 31674 13822
rect 31468 13758 31469 13810
rect 31521 13758 31545 13810
rect 31597 13758 31621 13810
rect 31673 13758 31674 13810
rect 31468 13745 31674 13758
rect 31468 13693 31469 13745
rect 31521 13693 31545 13745
rect 31597 13693 31621 13745
rect 31673 13693 31674 13745
rect 31468 13680 31674 13693
rect 31468 13628 31469 13680
rect 31521 13628 31545 13680
rect 31597 13628 31621 13680
rect 31673 13628 31674 13680
rect 31468 13615 31674 13628
rect 31468 13563 31469 13615
rect 31521 13563 31545 13615
rect 31597 13563 31621 13615
rect 31673 13563 31674 13615
rect 31468 13550 31674 13563
rect 31468 13498 31469 13550
rect 31521 13498 31545 13550
rect 31597 13498 31621 13550
rect 31673 13498 31674 13550
rect 31468 13485 31674 13498
rect 31468 13433 31469 13485
rect 31521 13433 31545 13485
rect 31597 13433 31621 13485
rect 31673 13433 31674 13485
rect 31468 13420 31674 13433
rect 31468 13368 31469 13420
rect 31521 13368 31545 13420
rect 31597 13368 31621 13420
rect 31673 13368 31674 13420
rect 31468 13355 31674 13368
rect 31468 13303 31469 13355
rect 31521 13303 31545 13355
rect 31597 13303 31621 13355
rect 31673 13303 31674 13355
rect 31468 13290 31674 13303
rect 31468 13238 31469 13290
rect 31521 13238 31545 13290
rect 31597 13238 31621 13290
rect 31673 13238 31674 13290
rect 31468 13225 31674 13238
rect 31468 13173 31469 13225
rect 31521 13173 31545 13225
rect 31597 13173 31621 13225
rect 31673 13173 31674 13225
rect 31468 13160 31674 13173
rect 31468 13108 31469 13160
rect 31521 13108 31545 13160
rect 31597 13108 31621 13160
rect 31673 13108 31674 13160
rect 31468 13095 31674 13108
rect 31468 13043 31469 13095
rect 31521 13043 31545 13095
rect 31597 13043 31621 13095
rect 31673 13043 31674 13095
rect 15143 13032 15463 13033
rect 15143 12980 15149 13032
rect 15201 12980 15213 13032
rect 15265 12980 15277 13032
rect 15329 12980 15341 13032
rect 15393 12980 15405 13032
rect 15457 12980 15463 13032
rect 15143 12962 15463 12980
rect 15143 12910 15149 12962
rect 15201 12910 15213 12962
rect 15265 12910 15277 12962
rect 15329 12910 15341 12962
rect 15393 12910 15405 12962
rect 15457 12910 15463 12962
rect 15143 12892 15463 12910
rect 15143 12840 15149 12892
rect 15201 12840 15213 12892
rect 15265 12840 15277 12892
rect 15329 12840 15341 12892
rect 15393 12840 15405 12892
rect 15457 12840 15463 12892
rect 15143 12822 15463 12840
rect 15143 12770 15149 12822
rect 15201 12770 15213 12822
rect 15265 12770 15277 12822
rect 15329 12770 15341 12822
rect 15393 12770 15405 12822
rect 15457 12770 15463 12822
rect 4073 11653 4079 11705
rect 4131 11653 4143 11705
rect 4195 11653 4201 11705
rect 5109 11653 5115 11705
rect 5167 11653 5179 11705
rect 5231 11653 5237 11705
rect 4073 11142 4201 11653
tri 5160 11628 5185 11653 ne
rect 4073 11090 4085 11142
rect 4137 11090 4149 11142
rect 4073 11084 4201 11090
tri 2927 9678 3003 9754 ne
tri 4657 7307 4664 7314 sw
rect -593 7009 -587 7061
rect -535 7009 -505 7061
rect -453 7009 -423 7061
rect -371 7009 -341 7061
rect -289 7009 -259 7061
rect -207 7009 -201 7061
rect -593 6997 -201 7009
rect -593 6945 -587 6997
rect -535 6945 -505 6997
rect -453 6945 -423 6997
rect -371 6945 -341 6997
rect -289 6945 -259 6997
rect -207 6945 -201 6997
tri 3842 6669 3846 6673 nw
tri 4660 6669 4664 6673 nw
tri 5159 6302 5185 6328 se
rect 5185 6302 5237 11653
rect 7390 11104 7518 11865
rect 15143 11703 15463 12770
rect 31468 13030 31674 13043
rect 31468 12978 31469 13030
rect 31521 12978 31545 13030
rect 31597 12978 31621 13030
rect 31673 12978 31674 13030
rect 31468 12965 31674 12978
rect 31468 12913 31469 12965
rect 31521 12913 31545 12965
rect 31597 12913 31621 12965
rect 31673 12913 31674 12965
rect 31468 12900 31674 12913
rect 31468 12848 31469 12900
rect 31521 12848 31545 12900
rect 31597 12848 31621 12900
rect 31673 12848 31674 12900
rect 31468 12835 31674 12848
rect 31468 12783 31469 12835
rect 31521 12783 31545 12835
rect 31597 12783 31621 12835
rect 31673 12783 31674 12835
rect 31468 12770 31674 12783
rect 31468 12718 31469 12770
rect 31521 12718 31545 12770
rect 31597 12718 31621 12770
rect 31673 12718 31674 12770
rect 31468 12705 31674 12718
rect 31468 12653 31469 12705
rect 31521 12653 31545 12705
rect 31597 12653 31621 12705
rect 31673 12653 31674 12705
rect 31468 12640 31674 12653
rect 31468 12588 31469 12640
rect 31521 12588 31545 12640
rect 31597 12588 31621 12640
rect 31673 12588 31674 12640
rect 31468 12575 31674 12588
rect 31468 12523 31469 12575
rect 31521 12523 31545 12575
rect 31597 12523 31621 12575
rect 31673 12523 31674 12575
rect 31468 12510 31674 12523
rect 31468 12458 31469 12510
rect 31521 12458 31545 12510
rect 31597 12458 31621 12510
rect 31673 12458 31674 12510
rect 31468 12445 31674 12458
rect 31468 12393 31469 12445
rect 31521 12393 31545 12445
rect 31597 12393 31621 12445
rect 31673 12393 31674 12445
rect 31468 12380 31674 12393
rect 31468 12328 31469 12380
rect 31521 12328 31545 12380
rect 31597 12328 31621 12380
rect 31673 12328 31674 12380
rect 31468 12315 31674 12328
rect 31468 12263 31469 12315
rect 31521 12263 31545 12315
rect 31597 12263 31621 12315
rect 31673 12263 31674 12315
rect 31468 12250 31674 12263
rect 31468 12198 31469 12250
rect 31521 12198 31545 12250
rect 31597 12198 31621 12250
rect 31673 12198 31674 12250
rect 31468 12185 31674 12198
rect 31468 12133 31469 12185
rect 31521 12133 31545 12185
rect 31597 12133 31621 12185
rect 31673 12133 31674 12185
rect 31468 12120 31674 12133
rect 31468 12068 31469 12120
rect 31521 12068 31545 12120
rect 31597 12068 31621 12120
rect 31673 12068 31674 12120
rect 31468 12055 31674 12068
rect 17611 12037 18413 12039
rect 17611 11985 17617 12037
rect 17669 11985 17685 12037
rect 17737 11985 17752 12037
rect 17804 11985 17819 12037
rect 17871 11985 17886 12037
rect 17938 11985 17953 12037
rect 18005 11985 18020 12037
rect 18072 11985 18087 12037
rect 18139 11985 18154 12037
rect 18206 11985 18221 12037
rect 18273 11985 18288 12037
rect 18340 11985 18355 12037
rect 18407 11985 18413 12037
rect 17611 11965 18413 11985
rect 17611 11913 17617 11965
rect 17669 11913 17685 11965
rect 17737 11913 17752 11965
rect 17804 11913 17819 11965
rect 17871 11913 17886 11965
rect 17938 11913 17953 11965
rect 18005 11913 18020 11965
rect 18072 11913 18087 11965
rect 18139 11913 18154 11965
rect 18206 11913 18221 11965
rect 18273 11913 18288 11965
rect 18340 11913 18355 11965
rect 18407 11913 18413 11965
rect 17611 11893 18413 11913
rect 17611 11841 17617 11893
rect 17669 11841 17685 11893
rect 17737 11841 17752 11893
rect 17804 11841 17819 11893
rect 17871 11841 17886 11893
rect 17938 11841 17953 11893
rect 18005 11841 18020 11893
rect 18072 11841 18087 11893
rect 18139 11841 18154 11893
rect 18206 11841 18221 11893
rect 18273 11841 18288 11893
rect 18340 11841 18355 11893
rect 18407 11841 18413 11893
rect 17611 11821 18413 11841
rect 17611 11769 17617 11821
rect 17669 11769 17685 11821
rect 17737 11769 17752 11821
rect 17804 11769 17819 11821
rect 17871 11769 17886 11821
rect 17938 11769 17953 11821
rect 18005 11769 18020 11821
rect 18072 11769 18087 11821
rect 18139 11769 18154 11821
rect 18206 11769 18221 11821
rect 18273 11769 18288 11821
rect 18340 11769 18355 11821
rect 18407 11769 18413 11821
rect 17611 11767 18413 11769
rect 31468 12003 31469 12055
rect 31521 12003 31545 12055
rect 31597 12003 31621 12055
rect 31673 12003 31674 12055
rect 31468 11990 31674 12003
rect 31468 11938 31469 11990
rect 31521 11938 31545 11990
rect 31597 11938 31621 11990
rect 31673 11938 31674 11990
rect 31468 11925 31674 11938
rect 31468 11873 31469 11925
rect 31521 11873 31545 11925
rect 31597 11873 31621 11925
rect 31673 11873 31674 11925
rect 31468 11860 31674 11873
rect 31468 11808 31469 11860
rect 31521 11808 31545 11860
rect 31597 11808 31621 11860
rect 31673 11808 31674 11860
rect 31468 11795 31674 11808
rect 31468 11743 31469 11795
rect 31521 11743 31545 11795
rect 31597 11743 31621 11795
rect 31673 11743 31674 11795
rect 31468 11730 31674 11743
rect 31468 11678 31469 11730
rect 31521 11678 31545 11730
rect 31597 11678 31621 11730
rect 31673 11678 31674 11730
rect 31468 11665 31674 11678
rect 31468 11613 31469 11665
rect 31521 11613 31545 11665
rect 31597 11613 31621 11665
rect 31673 11613 31674 11665
rect 31468 11600 31674 11613
rect 19830 11582 20321 11583
rect 19830 11530 19836 11582
rect 19888 11530 19908 11582
rect 19960 11530 19979 11582
rect 20031 11530 20050 11582
rect 20102 11530 20121 11582
rect 20173 11530 20192 11582
rect 20244 11530 20263 11582
rect 20315 11530 20321 11582
rect 19830 11514 20321 11530
rect 19830 11462 19836 11514
rect 19888 11462 19908 11514
rect 19960 11462 19979 11514
rect 20031 11462 20050 11514
rect 20102 11462 20121 11514
rect 20173 11462 20192 11514
rect 20244 11462 20263 11514
rect 20315 11462 20321 11514
rect 19830 11446 20321 11462
rect 19830 11394 19836 11446
rect 19888 11394 19908 11446
rect 19960 11394 19979 11446
rect 20031 11394 20050 11446
rect 20102 11394 20121 11446
rect 20173 11394 20192 11446
rect 20244 11394 20263 11446
rect 20315 11394 20321 11446
rect 19830 11378 20321 11394
rect 19830 11326 19836 11378
rect 19888 11326 19908 11378
rect 19960 11326 19979 11378
rect 20031 11326 20050 11378
rect 20102 11326 20121 11378
rect 20173 11326 20192 11378
rect 20244 11326 20263 11378
rect 20315 11326 20321 11378
rect 19830 11325 20321 11326
rect 31468 11548 31469 11600
rect 31521 11548 31545 11600
rect 31597 11548 31621 11600
rect 31673 11548 31674 11600
rect 31468 11535 31674 11548
rect 31468 11483 31469 11535
rect 31521 11483 31545 11535
rect 31597 11483 31621 11535
rect 31673 11483 31674 11535
rect 31468 11470 31674 11483
rect 31468 11418 31469 11470
rect 31521 11418 31545 11470
rect 31597 11418 31621 11470
rect 31673 11418 31674 11470
rect 31468 11405 31674 11418
rect 31468 11353 31469 11405
rect 31521 11353 31545 11405
rect 31597 11353 31621 11405
rect 31673 11353 31674 11405
rect 31468 11340 31674 11353
rect 31468 11288 31469 11340
rect 31521 11288 31545 11340
rect 31597 11288 31621 11340
rect 31673 11288 31674 11340
rect 31468 11275 31674 11288
rect 13884 11222 13890 11274
rect 13942 11222 13981 11274
rect 14033 11222 14071 11274
rect 14123 11222 14129 11274
rect 14418 11222 14424 11274
rect 14476 11222 14489 11274
rect 14541 11222 14553 11274
rect 14605 11222 14617 11274
rect 14669 11222 14681 11274
rect 14733 11222 14739 11274
tri 9196 10801 9230 10835 ne
rect 9230 10499 9262 10835
tri 9262 10801 9296 10835 nw
rect 14418 10551 14739 11222
rect 31468 11223 31469 11275
rect 31521 11223 31545 11275
rect 31597 11223 31621 11275
rect 31673 11223 31674 11275
rect 31468 11210 31674 11223
rect 31468 11158 31469 11210
rect 31521 11158 31545 11210
rect 31597 11158 31621 11210
rect 31673 11158 31674 11210
rect 31468 11145 31674 11158
rect 31468 11093 31469 11145
rect 31521 11093 31545 11145
rect 31597 11093 31621 11145
rect 31673 11093 31674 11145
rect 31468 11087 31674 11093
tri 9262 10499 9273 10510 sw
rect 13884 10499 13890 10551
rect 13942 10499 13981 10551
rect 14033 10499 14071 10551
rect 14123 10499 14129 10551
rect 14418 10499 14424 10551
rect 14476 10499 14489 10551
rect 14541 10499 14553 10551
rect 14605 10499 14617 10551
rect 14669 10499 14681 10551
rect 14733 10499 14739 10551
rect 9230 10496 9273 10499
tri 9230 10475 9251 10496 ne
rect 9251 10475 9273 10496
tri 9273 10475 9297 10499 sw
tri 9251 10464 9262 10475 ne
rect 9262 10464 9297 10475
tri 9262 10429 9297 10464 ne
tri 9297 10429 9343 10475 sw
tri 9297 10383 9343 10429 ne
tri 9343 10383 9389 10429 sw
tri 9343 10337 9389 10383 ne
tri 9389 10369 9403 10383 sw
rect 9389 10337 9403 10369
tri 9403 10337 9435 10369 sw
tri 9389 10323 9403 10337 ne
rect 6019 9871 6025 9923
rect 6077 9871 6089 9923
rect 6141 9871 6147 9923
rect 5623 9221 5675 9227
rect 5623 9157 5675 9169
rect 5298 7488 5350 7497
rect 5298 7424 5350 7436
rect 5298 7366 5350 7372
tri 5298 7356 5308 7366 ne
tri 5145 6288 5159 6302 se
rect 5159 6288 5237 6302
tri 5110 6253 5145 6288 se
rect 5145 6253 5237 6288
tri 5093 6236 5110 6253 se
rect 5110 6236 5220 6253
tri 5220 6236 5237 6253 nw
tri 5079 6222 5093 6236 se
rect 5093 6222 5206 6236
tri 5206 6222 5220 6236 nw
tri 5077 6220 5079 6222 se
rect 5079 6220 5181 6222
rect 5077 6197 5181 6220
tri 5181 6197 5206 6222 nw
rect 5077 6170 5154 6197
tri 5154 6170 5181 6197 nw
tri 5281 6170 5308 6197 se
rect 5308 6183 5340 7366
tri 5340 7356 5350 7366 nw
rect 5308 6170 5327 6183
tri 5327 6170 5340 6183 nw
rect 5077 6151 5135 6170
tri 5135 6151 5154 6170 nw
tri 5262 6151 5281 6170 se
rect 5281 6151 5308 6170
tri 5308 6151 5327 6170 nw
rect 74 5764 194 5770
rect 74 5648 76 5764
rect 192 5648 194 5764
rect 74 5470 194 5648
rect 2145 5763 2261 5769
rect 5077 5683 5129 6151
tri 5129 6145 5135 6151 nw
tri 5256 6145 5262 6151 se
tri 5216 6105 5256 6145 se
rect 5256 6105 5262 6145
tri 5262 6105 5308 6151 nw
tri 5174 6063 5216 6105 se
rect 5216 6063 5220 6105
tri 5220 6063 5262 6105 nw
rect 5174 5898 5206 6063
tri 5206 6049 5220 6063 nw
tri 5206 5898 5220 5912 sw
tri 5174 5852 5220 5898 ne
tri 5220 5852 5266 5898 sw
tri 5220 5806 5266 5852 ne
tri 5266 5816 5302 5852 sw
rect 5266 5806 5302 5816
tri 5266 5802 5270 5806 ne
tri 5077 5650 5110 5683 ne
rect 5110 5650 5129 5683
tri 5129 5650 5237 5758 sw
rect 2145 5641 2261 5647
tri 5110 5641 5119 5650 ne
rect 5119 5641 5237 5650
tri 5119 5631 5129 5641 ne
rect 5129 5631 5237 5641
tri 5129 5627 5133 5631 ne
rect 5133 5627 5237 5631
tri 4739 5626 4740 5627 nw
tri 5133 5626 5134 5627 ne
rect 5134 5626 5237 5627
tri 5134 5613 5147 5626 ne
rect 5147 5613 5237 5626
rect -600 4816 -200 4846
rect -600 4764 -594 4816
rect -542 4764 -510 4816
rect -458 4764 -426 4816
rect -374 4764 -342 4816
rect -290 4764 -258 4816
rect -206 4764 -200 4816
rect -600 0 -200 4764
rect 512 1323 519 1503
rect 635 1323 1234 1503
rect 1350 1323 1861 1503
rect 1977 1323 2573 1503
rect 2689 1323 3586 1503
rect 512 1195 3586 1323
rect 3870 0 3922 5613
rect 3950 0 4002 5613
rect 4384 0 4436 5613
rect 4464 0 4516 5613
tri 5147 5575 5185 5613 ne
rect 4847 3252 4899 3258
rect 4847 3188 4899 3200
rect 4847 3130 4899 3136
rect 5185 0 5237 5613
rect 5270 1120 5302 5806
rect 5623 0 5675 9105
tri 5945 5626 6019 5700 se
rect 6019 5678 6071 9871
tri 6071 9846 6096 9871 nw
rect 9403 9275 9435 10337
rect 9987 9804 10128 10369
rect 10015 9478 10067 9794
tri 11626 9735 11665 9774 se
tri 12462 9678 12519 9735 ne
rect 12839 9678 12862 9735
tri 12862 9678 12919 9735 nw
tri 12839 9655 12862 9678 nw
tri 13412 9494 13432 9514 se
rect 13432 9494 13484 9798
tri 10067 9478 10083 9494 sw
tri 13396 9478 13412 9494 se
rect 13412 9492 13484 9494
rect 13412 9478 13432 9492
rect 10015 9472 10083 9478
tri 10015 9404 10083 9472 ne
tri 10083 9404 10157 9478 sw
tri 13358 9440 13396 9478 se
rect 13396 9440 13432 9478
tri 13432 9440 13484 9492 nw
tri 13335 9417 13358 9440 se
tri 10506 9409 10514 9417 ne
tri 13327 9409 13335 9417 se
rect 13335 9409 13358 9417
tri 13322 9404 13327 9409 se
rect 13327 9404 13358 9409
tri 10083 9330 10157 9404 ne
tri 10157 9330 10231 9404 sw
tri 13284 9366 13322 9404 se
rect 13322 9366 13358 9404
tri 13358 9366 13432 9440 nw
tri 13253 9335 13284 9366 se
rect 13284 9335 13327 9366
tri 13327 9335 13358 9366 nw
rect 13253 9330 13322 9335
tri 13322 9330 13327 9335 nw
tri 10157 9289 10198 9330 ne
rect 10198 9289 10231 9330
tri 9403 9256 9422 9275 ne
rect 9422 9256 9435 9275
tri 9435 9256 9468 9289 sw
tri 10198 9256 10231 9289 ne
tri 10231 9256 10305 9330 sw
tri 9422 9247 9431 9256 ne
rect 9431 9247 9468 9256
tri 9468 9247 9477 9256 sw
tri 10231 9247 10240 9256 ne
rect 10240 9247 10785 9256
rect 6114 9195 6123 9247
rect 6175 9195 6187 9247
rect 6239 9195 6245 9247
tri 9431 9243 9435 9247 ne
rect 9435 9243 9477 9247
tri 9477 9243 9481 9247 sw
tri 10044 9243 10048 9247 se
rect 10048 9243 10054 9247
tri 9435 9200 9478 9243 ne
rect 9478 9200 10054 9243
tri 10043 9195 10048 9200 ne
rect 10048 9195 10054 9200
rect 10106 9195 10118 9247
rect 10170 9195 10176 9247
tri 10240 9204 10283 9247 ne
rect 10283 9204 10785 9247
rect 10837 9204 10849 9256
rect 10901 9204 10907 9256
tri 10819 9195 10828 9204 ne
rect 10828 9195 10907 9204
rect 6114 9194 6201 9195
tri 6114 9158 6150 9194 ne
tri 6116 7481 6150 7515 se
rect 6150 7481 6201 9194
tri 6201 9158 6238 9195 nw
tri 10828 9168 10855 9195 ne
tri 6280 8426 6282 8428 se
tri 6598 8426 6600 8428 sw
tri 9457 7995 9494 8032 ne
tri 6201 7481 6235 7515 sw
rect 6114 7429 6123 7481
rect 6175 7429 6187 7481
rect 6239 7429 6245 7481
tri 8861 7307 8865 7311 sw
tri 8686 7211 8699 7224 sw
tri 8861 6669 8865 6673 nw
tri 8294 6049 8319 6074 se
tri 8217 5994 8272 6049 se
rect 8272 5997 8319 6049
rect 8272 5994 8291 5997
tri 8291 5994 8294 5997 nw
tri 8143 5822 8217 5896 se
rect 8217 5874 8269 5994
tri 8269 5972 8291 5994 nw
tri 8217 5822 8269 5874 nw
tri 6019 5626 6071 5678 nw
tri 8111 5790 8143 5822 se
rect 8143 5790 8185 5822
tri 8185 5790 8217 5822 nw
rect 8111 5770 8165 5790
tri 8165 5770 8185 5790 nw
rect 8111 5769 8164 5770
tri 8164 5769 8165 5770 nw
tri 5871 5552 5945 5626 se
tri 5945 5552 6019 5626 nw
tri 5797 5478 5871 5552 se
tri 5871 5478 5945 5552 nw
tri 5723 5404 5797 5478 se
tri 5797 5404 5871 5478 nw
tri 5703 5384 5723 5404 se
rect 5723 5384 5777 5404
tri 5777 5384 5797 5404 nw
rect 5703 0 5755 5384
tri 5755 5362 5777 5384 nw
tri 5940 2542 6125 2727 sw
rect 5940 2541 6126 2542
rect 5824 2540 6126 2541
tri 6126 2540 6127 2541 sw
rect 5824 2536 6127 2540
rect 5824 2484 5987 2536
rect 6039 2484 6051 2536
rect 6103 2484 6127 2536
rect 5824 2467 6127 2484
rect 5824 2415 5987 2467
rect 6039 2415 6051 2467
rect 6103 2415 6127 2467
rect 5824 2398 6127 2415
rect 5824 2346 5987 2398
rect 6039 2346 6051 2398
rect 6103 2346 6127 2398
rect 5824 2205 6127 2346
rect 5824 2153 5994 2205
rect 6046 2153 6069 2205
rect 6121 2153 6127 2205
rect 5824 1705 6127 2153
rect 5824 1653 5987 1705
rect 6039 1653 6051 1705
rect 6103 1653 6127 1705
rect 5824 1625 6127 1653
rect 5824 1573 5987 1625
rect 6039 1573 6051 1625
rect 6103 1573 6127 1625
rect 5824 1524 6127 1573
rect 6665 0 6717 454
rect 6745 0 6797 454
tri 6871 399 6889 417 ne
rect 6889 399 6981 417
tri 6981 399 6999 417 nw
rect 6889 0 6958 399
tri 6958 376 6981 399 nw
rect 8031 0 8083 5613
rect 8111 0 8163 5769
tri 8163 5768 8164 5769 nw
rect 9574 4853 9626 5613
tri 10179 5597 10195 5613 nw
tri 9574 4829 9598 4853 ne
rect 9598 4829 9626 4853
tri 9626 4829 9672 4875 sw
tri 9598 4801 9626 4829 ne
rect 9626 4801 9672 4829
tri 9626 4755 9672 4801 ne
tri 9672 4755 9746 4829 sw
tri 9672 4733 9694 4755 ne
tri 9620 2134 9694 2208 se
rect 9694 2186 9746 4755
tri 9694 2134 9746 2186 nw
tri 9546 2060 9620 2134 se
tri 9620 2060 9694 2134 nw
tri 9521 2035 9546 2060 se
rect 9546 2035 9595 2060
tri 9595 2035 9620 2060 nw
rect 8541 1740 8737 1746
rect 8541 1688 8549 1740
rect 8601 1688 8613 1740
rect 8665 1688 8677 1740
rect 8729 1688 8737 1740
rect 8541 1671 8737 1688
rect 8541 1619 8549 1671
rect 8601 1619 8613 1671
rect 8665 1619 8677 1671
rect 8729 1619 8737 1671
rect 8541 1602 8737 1619
rect 8541 1550 8549 1602
rect 8601 1550 8613 1602
rect 8665 1550 8677 1602
rect 8729 1550 8737 1602
rect 8541 228 8737 1550
rect 9521 0 9573 2035
tri 9573 2013 9595 2035 nw
rect 10855 0 10907 9195
tri 13179 9118 13253 9192 se
rect 13253 9170 13305 9330
tri 13305 9313 13322 9330 nw
tri 13253 9118 13305 9170 nw
rect 13179 7282 13231 9118
tri 13231 9096 13253 9118 nw
rect 18531 8371 18537 8423
rect 18589 8371 18601 8423
rect 18653 8371 18665 8423
rect 18717 8371 18729 8423
rect 18781 8371 18793 8423
rect 18845 8371 18857 8423
rect 18909 8371 18915 8423
rect 13259 7379 13375 7385
rect 13311 7327 13323 7379
rect 13259 7321 13375 7327
tri 13231 7282 13235 7286 sw
rect 13179 7264 13235 7282
tri 13179 7260 13183 7264 ne
tri 13128 3493 13183 3548 se
rect 13183 3526 13235 7264
rect 18531 6575 18931 8109
rect 21680 7536 22220 7545
rect 21680 6600 21682 7536
rect 22218 6600 22220 7536
rect 21680 6575 22220 6600
rect 21680 6519 21682 6575
rect 21738 6519 21762 6575
rect 21818 6519 21842 6575
rect 21898 6519 21922 6575
rect 21978 6519 22002 6575
rect 22058 6519 22082 6575
rect 22138 6519 22162 6575
rect 22218 6519 22220 6575
rect 21680 6494 22220 6519
rect 21680 6438 21682 6494
rect 21738 6438 21762 6494
rect 21818 6438 21842 6494
rect 21898 6438 21922 6494
rect 21978 6438 22002 6494
rect 22058 6438 22082 6494
rect 22138 6438 22162 6494
rect 22218 6438 22220 6494
rect 27764 7482 28018 7491
rect 27764 7426 27765 7482
rect 27821 7426 27863 7482
rect 27919 7426 27961 7482
rect 28017 7426 28018 7482
rect 27764 7397 28018 7426
rect 27764 7341 27765 7397
rect 27821 7341 27863 7397
rect 27919 7341 27961 7397
rect 28017 7341 28018 7397
rect 27764 7312 28018 7341
rect 27764 7256 27765 7312
rect 27821 7256 27863 7312
rect 27919 7256 27961 7312
rect 28017 7256 28018 7312
rect 27764 7226 28018 7256
rect 27764 7170 27765 7226
rect 27821 7170 27863 7226
rect 27919 7170 27961 7226
rect 28017 7170 28018 7226
rect 27764 7140 28018 7170
rect 27764 7084 27765 7140
rect 27821 7084 27863 7140
rect 27919 7084 27961 7140
rect 28017 7084 28018 7140
rect 27764 7054 28018 7084
rect 27764 6998 27765 7054
rect 27821 6998 27863 7054
rect 27919 6998 27961 7054
rect 28017 6998 28018 7054
rect 27764 6968 28018 6998
rect 27764 6912 27765 6968
rect 27821 6912 27863 6968
rect 27919 6912 27961 6968
rect 28017 6912 28018 6968
rect 27764 6882 28018 6912
rect 27764 6826 27765 6882
rect 27821 6826 27863 6882
rect 27919 6826 27961 6882
rect 28017 6826 28018 6882
rect 27764 6796 28018 6826
rect 27764 6740 27765 6796
rect 27821 6740 27863 6796
rect 27919 6740 27961 6796
rect 28017 6740 28018 6796
rect 27764 6710 28018 6740
rect 27764 6654 27765 6710
rect 27821 6654 27863 6710
rect 27919 6654 27961 6710
rect 28017 6654 28018 6710
rect 27764 6624 28018 6654
rect 27764 6568 27765 6624
rect 27821 6568 27863 6624
rect 27919 6568 27961 6624
rect 28017 6568 28018 6624
rect 27764 6538 28018 6568
rect 27764 6482 27765 6538
rect 27821 6482 27863 6538
rect 27919 6482 27961 6538
rect 28017 6482 28018 6538
rect 27764 6473 28018 6482
rect 21680 6429 22220 6438
rect 23952 6302 23958 6354
rect 24010 6302 24042 6354
rect 24094 6302 24126 6354
rect 24178 6302 24209 6354
rect 24261 6302 24267 6354
rect 23952 6288 24267 6302
rect 23952 6236 23958 6288
rect 24010 6236 24042 6288
rect 24094 6236 24126 6288
rect 24178 6236 24209 6288
rect 24261 6236 24267 6288
tri 30272 6283 30273 6284 se
rect 23952 6222 24267 6236
rect 23952 6170 23958 6222
rect 24010 6170 24042 6222
rect 24094 6170 24126 6222
rect 24178 6170 24209 6222
rect 24261 6170 24267 6222
rect 13661 5613 13713 5781
tri 30586 5507 30617 5538 nw
rect 13183 3493 13202 3526
tri 13202 3493 13235 3526 nw
rect 32404 3563 32724 3573
rect 32460 3507 32492 3563
rect 32548 3507 32580 3563
rect 32636 3507 32668 3563
rect 13128 0 13180 3493
tri 13180 3471 13202 3493 nw
rect 32404 3480 32724 3507
rect 32460 3424 32492 3480
rect 32548 3424 32580 3480
rect 32636 3424 32668 3480
rect 32404 3397 32724 3424
rect 32460 3341 32492 3397
rect 32548 3341 32580 3397
rect 32636 3341 32668 3397
rect 32404 3314 32724 3341
rect 32460 3258 32492 3314
rect 32548 3258 32580 3314
rect 32636 3258 32668 3314
rect 32404 3231 32724 3258
rect 32460 3175 32492 3231
rect 32548 3175 32580 3231
rect 32636 3175 32668 3231
rect 32404 3148 32724 3175
rect 32460 3092 32492 3148
rect 32548 3092 32580 3148
rect 32636 3092 32668 3148
rect 32404 3065 32724 3092
rect 32460 3009 32492 3065
rect 32548 3009 32580 3065
rect 32636 3009 32668 3065
rect 32404 2982 32724 3009
rect 32460 2926 32492 2982
rect 32548 2926 32580 2982
rect 32636 2926 32668 2982
rect 32404 2899 32724 2926
rect 32460 2843 32492 2899
rect 32548 2843 32580 2899
rect 32636 2843 32668 2899
rect 32404 2816 32724 2843
rect 32460 2760 32492 2816
rect 32548 2760 32580 2816
rect 32636 2760 32668 2816
rect 32404 2733 32724 2760
rect 32460 2677 32492 2733
rect 32548 2677 32580 2733
rect 32636 2677 32668 2733
rect 32404 2650 32724 2677
rect 32460 2594 32492 2650
rect 32548 2594 32580 2650
rect 32636 2594 32668 2650
rect 32404 2567 32724 2594
rect 32460 2511 32492 2567
rect 32548 2511 32580 2567
rect 32636 2511 32668 2567
rect 32404 2483 32724 2511
rect 32460 2427 32492 2483
rect 32548 2427 32580 2483
rect 32636 2427 32668 2483
rect 32404 2399 32724 2427
rect 32460 2343 32492 2399
rect 32548 2343 32580 2399
rect 32636 2343 32668 2399
rect 32404 2205 32724 2343
rect 32460 2149 32492 2205
rect 32548 2149 32580 2205
rect 32636 2149 32668 2205
rect 32404 2124 32724 2149
rect 32460 2068 32492 2124
rect 32548 2068 32580 2124
rect 32636 2068 32668 2124
rect 32404 2043 32724 2068
rect 32460 1987 32492 2043
rect 32548 1987 32580 2043
rect 32636 1987 32668 2043
rect 32404 1962 32724 1987
rect 32460 1906 32492 1962
rect 32548 1906 32580 1962
rect 32636 1906 32668 1962
rect 32404 1881 32724 1906
rect 32460 1825 32492 1881
rect 32548 1825 32580 1881
rect 32636 1825 32668 1881
rect 32404 1800 32724 1825
rect 32460 1744 32492 1800
rect 32548 1744 32580 1800
rect 32636 1744 32668 1800
rect 32404 1719 32724 1744
rect 32460 1663 32492 1719
rect 32548 1663 32580 1719
rect 32636 1663 32668 1719
rect 32404 1638 32724 1663
rect 32460 1582 32492 1638
rect 32548 1582 32580 1638
rect 32636 1582 32668 1638
rect 32404 1557 32724 1582
rect 32460 1501 32492 1557
rect 32548 1501 32580 1557
rect 32636 1501 32668 1557
rect 32404 1476 32724 1501
rect 32460 1420 32492 1476
rect 32548 1420 32580 1476
rect 32636 1420 32668 1476
rect 32404 1395 32724 1420
rect 32460 1339 32492 1395
rect 32548 1339 32580 1395
rect 32636 1339 32668 1395
rect 32404 1313 32724 1339
rect 32460 1257 32492 1313
rect 32548 1257 32580 1313
rect 32636 1257 32668 1313
rect 32404 1231 32724 1257
rect 32460 1175 32492 1231
rect 32548 1175 32580 1231
rect 32636 1175 32668 1231
rect 32404 1159 32724 1175
rect 13804 0 13856 75
rect 14433 0 14582 517
tri 14642 379 14690 427 se
rect 14690 379 14892 517
rect 14642 174 14892 379
tri 14642 126 14690 174 ne
rect 14690 0 14892 174
rect 15021 0 15073 517
rect 15237 0 15289 517
rect 15332 0 15652 517
rect 15713 0 16033 517
rect 17779 0 17949 454
rect 17977 0 18146 454
<< via2 >>
rect 21682 6600 22218 7536
rect 21682 6519 21738 6575
rect 21762 6519 21818 6575
rect 21842 6519 21898 6575
rect 21922 6519 21978 6575
rect 22002 6519 22058 6575
rect 22082 6519 22138 6575
rect 22162 6519 22218 6575
rect 21682 6438 21738 6494
rect 21762 6438 21818 6494
rect 21842 6438 21898 6494
rect 21922 6438 21978 6494
rect 22002 6438 22058 6494
rect 22082 6438 22138 6494
rect 22162 6438 22218 6494
rect 27765 7426 27821 7482
rect 27863 7426 27919 7482
rect 27961 7426 28017 7482
rect 27765 7341 27821 7397
rect 27863 7341 27919 7397
rect 27961 7341 28017 7397
rect 27765 7256 27821 7312
rect 27863 7256 27919 7312
rect 27961 7256 28017 7312
rect 27765 7170 27821 7226
rect 27863 7170 27919 7226
rect 27961 7170 28017 7226
rect 27765 7084 27821 7140
rect 27863 7084 27919 7140
rect 27961 7084 28017 7140
rect 27765 6998 27821 7054
rect 27863 6998 27919 7054
rect 27961 6998 28017 7054
rect 27765 6912 27821 6968
rect 27863 6912 27919 6968
rect 27961 6912 28017 6968
rect 27765 6826 27821 6882
rect 27863 6826 27919 6882
rect 27961 6826 28017 6882
rect 27765 6740 27821 6796
rect 27863 6740 27919 6796
rect 27961 6740 28017 6796
rect 27765 6654 27821 6710
rect 27863 6654 27919 6710
rect 27961 6654 28017 6710
rect 27765 6568 27821 6624
rect 27863 6568 27919 6624
rect 27961 6568 28017 6624
rect 27765 6482 27821 6538
rect 27863 6482 27919 6538
rect 27961 6482 28017 6538
rect 32404 3507 32460 3563
rect 32492 3507 32548 3563
rect 32580 3507 32636 3563
rect 32668 3507 32724 3563
rect 32404 3424 32460 3480
rect 32492 3424 32548 3480
rect 32580 3424 32636 3480
rect 32668 3424 32724 3480
rect 32404 3341 32460 3397
rect 32492 3341 32548 3397
rect 32580 3341 32636 3397
rect 32668 3341 32724 3397
rect 32404 3258 32460 3314
rect 32492 3258 32548 3314
rect 32580 3258 32636 3314
rect 32668 3258 32724 3314
rect 32404 3175 32460 3231
rect 32492 3175 32548 3231
rect 32580 3175 32636 3231
rect 32668 3175 32724 3231
rect 32404 3092 32460 3148
rect 32492 3092 32548 3148
rect 32580 3092 32636 3148
rect 32668 3092 32724 3148
rect 32404 3009 32460 3065
rect 32492 3009 32548 3065
rect 32580 3009 32636 3065
rect 32668 3009 32724 3065
rect 32404 2926 32460 2982
rect 32492 2926 32548 2982
rect 32580 2926 32636 2982
rect 32668 2926 32724 2982
rect 32404 2843 32460 2899
rect 32492 2843 32548 2899
rect 32580 2843 32636 2899
rect 32668 2843 32724 2899
rect 32404 2760 32460 2816
rect 32492 2760 32548 2816
rect 32580 2760 32636 2816
rect 32668 2760 32724 2816
rect 32404 2677 32460 2733
rect 32492 2677 32548 2733
rect 32580 2677 32636 2733
rect 32668 2677 32724 2733
rect 32404 2594 32460 2650
rect 32492 2594 32548 2650
rect 32580 2594 32636 2650
rect 32668 2594 32724 2650
rect 32404 2511 32460 2567
rect 32492 2511 32548 2567
rect 32580 2511 32636 2567
rect 32668 2511 32724 2567
rect 32404 2427 32460 2483
rect 32492 2427 32548 2483
rect 32580 2427 32636 2483
rect 32668 2427 32724 2483
rect 32404 2343 32460 2399
rect 32492 2343 32548 2399
rect 32580 2343 32636 2399
rect 32668 2343 32724 2399
rect 32404 2149 32460 2205
rect 32492 2149 32548 2205
rect 32580 2149 32636 2205
rect 32668 2149 32724 2205
rect 32404 2068 32460 2124
rect 32492 2068 32548 2124
rect 32580 2068 32636 2124
rect 32668 2068 32724 2124
rect 32404 1987 32460 2043
rect 32492 1987 32548 2043
rect 32580 1987 32636 2043
rect 32668 1987 32724 2043
rect 32404 1906 32460 1962
rect 32492 1906 32548 1962
rect 32580 1906 32636 1962
rect 32668 1906 32724 1962
rect 32404 1825 32460 1881
rect 32492 1825 32548 1881
rect 32580 1825 32636 1881
rect 32668 1825 32724 1881
rect 32404 1744 32460 1800
rect 32492 1744 32548 1800
rect 32580 1744 32636 1800
rect 32668 1744 32724 1800
rect 32404 1663 32460 1719
rect 32492 1663 32548 1719
rect 32580 1663 32636 1719
rect 32668 1663 32724 1719
rect 32404 1582 32460 1638
rect 32492 1582 32548 1638
rect 32580 1582 32636 1638
rect 32668 1582 32724 1638
rect 32404 1501 32460 1557
rect 32492 1501 32548 1557
rect 32580 1501 32636 1557
rect 32668 1501 32724 1557
rect 32404 1420 32460 1476
rect 32492 1420 32548 1476
rect 32580 1420 32636 1476
rect 32668 1420 32724 1476
rect 32404 1339 32460 1395
rect 32492 1339 32548 1395
rect 32580 1339 32636 1395
rect 32668 1339 32724 1395
rect 32404 1257 32460 1313
rect 32492 1257 32548 1313
rect 32580 1257 32636 1313
rect 32668 1257 32724 1313
rect 32404 1175 32460 1231
rect 32492 1175 32548 1231
rect 32580 1175 32636 1231
rect 32668 1175 32724 1231
<< metal3 >>
tri 3004 40058 3005 40059 sw
tri 2447 40056 2449 40058 se
rect 3004 40056 3005 40058
tri 3005 40056 3007 40058 sw
rect 112 22362 142 22392
rect 15909 20847 28761 24635
rect 112 19224 142 19254
rect 16482 18527 29018 20387
rect 112 16446 142 16476
rect 16640 15195 28558 18029
rect 112 13717 142 13747
rect 112 12366 142 12396
rect 112 11029 142 11059
rect 725 9638 755 9668
rect 112 8358 142 8388
rect 21675 7536 22225 7541
rect 725 6905 755 6935
rect 21675 6600 21682 7536
rect 22218 6600 22225 7536
rect 21675 6575 22225 6600
rect 21675 6519 21682 6575
rect 21738 6519 21762 6575
rect 21818 6519 21842 6575
rect 21898 6519 21922 6575
rect 21978 6519 22002 6575
rect 22058 6519 22082 6575
rect 22138 6519 22162 6575
rect 22218 6519 22225 6575
rect 21675 6494 22225 6519
rect 21675 6438 21682 6494
rect 21738 6438 21762 6494
rect 21818 6438 21842 6494
rect 21898 6438 21922 6494
rect 21978 6438 22002 6494
rect 22058 6438 22082 6494
rect 22138 6438 22162 6494
rect 22218 6438 22225 6494
rect 27759 7482 28023 7487
rect 27759 7426 27765 7482
rect 27821 7426 27863 7482
rect 27919 7426 27961 7482
rect 28017 7426 28023 7482
rect 27759 7397 28023 7426
rect 27759 7341 27765 7397
rect 27821 7341 27863 7397
rect 27919 7341 27961 7397
rect 28017 7341 28023 7397
rect 27759 7312 28023 7341
rect 27759 7256 27765 7312
rect 27821 7256 27863 7312
rect 27919 7256 27961 7312
rect 28017 7256 28023 7312
rect 27759 7226 28023 7256
rect 27759 7170 27765 7226
rect 27821 7170 27863 7226
rect 27919 7170 27961 7226
rect 28017 7170 28023 7226
rect 27759 7140 28023 7170
rect 27759 7084 27765 7140
rect 27821 7084 27863 7140
rect 27919 7084 27961 7140
rect 28017 7084 28023 7140
rect 27759 7054 28023 7084
rect 27759 6998 27765 7054
rect 27821 6998 27863 7054
rect 27919 6998 27961 7054
rect 28017 6998 28023 7054
rect 27759 6968 28023 6998
rect 27759 6912 27765 6968
rect 27821 6912 27863 6968
rect 27919 6912 27961 6968
rect 28017 6912 28023 6968
rect 27759 6882 28023 6912
rect 27759 6826 27765 6882
rect 27821 6826 27863 6882
rect 27919 6826 27961 6882
rect 28017 6826 28023 6882
rect 27759 6796 28023 6826
rect 27759 6740 27765 6796
rect 27821 6740 27863 6796
rect 27919 6740 27961 6796
rect 28017 6740 28023 6796
rect 27759 6710 28023 6740
rect 27759 6654 27765 6710
rect 27821 6654 27863 6710
rect 27919 6654 27961 6710
rect 28017 6654 28023 6710
rect 27759 6624 28023 6654
rect 27759 6568 27765 6624
rect 27821 6568 27863 6624
rect 27919 6568 27961 6624
rect 28017 6568 28023 6624
rect 27759 6538 28023 6568
rect 27759 6482 27765 6538
rect 27821 6482 27863 6538
rect 27919 6482 27961 6538
rect 28017 6482 28023 6538
rect 27759 6477 28023 6482
rect 21675 6433 22225 6438
rect 112 5593 142 5623
rect 725 4184 755 4214
rect 32000 3563 32729 3572
rect 32000 3507 32404 3563
rect 32460 3507 32492 3563
rect 32548 3507 32580 3563
rect 32636 3507 32668 3563
rect 32724 3507 32729 3563
rect 32000 3480 32729 3507
rect 32000 3424 32404 3480
rect 32460 3424 32492 3480
rect 32548 3424 32580 3480
rect 32636 3424 32668 3480
rect 32724 3424 32729 3480
rect 32000 3397 32729 3424
rect 32000 3341 32404 3397
rect 32460 3341 32492 3397
rect 32548 3341 32580 3397
rect 32636 3341 32668 3397
rect 32724 3341 32729 3397
rect 32000 3314 32729 3341
rect 32000 3258 32404 3314
rect 32460 3258 32492 3314
rect 32548 3258 32580 3314
rect 32636 3258 32668 3314
rect 32724 3258 32729 3314
rect 32000 3231 32729 3258
rect 32000 3175 32404 3231
rect 32460 3175 32492 3231
rect 32548 3175 32580 3231
rect 32636 3175 32668 3231
rect 32724 3175 32729 3231
rect 32000 3148 32729 3175
rect 32000 3092 32404 3148
rect 32460 3092 32492 3148
rect 32548 3092 32580 3148
rect 32636 3092 32668 3148
rect 32724 3092 32729 3148
rect 32000 3065 32729 3092
rect 32000 3009 32404 3065
rect 32460 3009 32492 3065
rect 32548 3009 32580 3065
rect 32636 3009 32668 3065
rect 32724 3009 32729 3065
rect 32000 2982 32729 3009
rect 32000 2926 32404 2982
rect 32460 2926 32492 2982
rect 32548 2926 32580 2982
rect 32636 2926 32668 2982
rect 32724 2926 32729 2982
rect 32000 2899 32729 2926
rect 32000 2843 32404 2899
rect 32460 2843 32492 2899
rect 32548 2843 32580 2899
rect 32636 2843 32668 2899
rect 32724 2843 32729 2899
rect 32000 2816 32729 2843
rect 725 2754 755 2784
rect 32000 2760 32404 2816
rect 32460 2760 32492 2816
rect 32548 2760 32580 2816
rect 32636 2760 32668 2816
rect 32724 2760 32729 2816
rect 32000 2733 32729 2760
rect 32000 2677 32404 2733
rect 32460 2677 32492 2733
rect 32548 2677 32580 2733
rect 32636 2677 32668 2733
rect 32724 2677 32729 2733
rect 32000 2650 32729 2677
rect 32000 2594 32404 2650
rect 32460 2594 32492 2650
rect 32548 2594 32580 2650
rect 32636 2594 32668 2650
rect 32724 2594 32729 2650
rect 32000 2567 32729 2594
rect 32000 2511 32404 2567
rect 32460 2511 32492 2567
rect 32548 2511 32580 2567
rect 32636 2511 32668 2567
rect 32724 2511 32729 2567
rect 32000 2483 32729 2511
rect 32000 2427 32404 2483
rect 32460 2427 32492 2483
rect 32548 2427 32580 2483
rect 32636 2427 32668 2483
rect 32724 2427 32729 2483
rect 32000 2399 32729 2427
rect 32000 2343 32404 2399
rect 32460 2343 32492 2399
rect 32548 2343 32580 2399
rect 32636 2343 32668 2399
rect 32724 2343 32729 2399
rect 32000 2334 32729 2343
rect 32000 2205 32730 2214
rect 32000 2149 32404 2205
rect 32460 2149 32492 2205
rect 32548 2149 32580 2205
rect 32636 2149 32668 2205
rect 32724 2149 32730 2205
rect 32000 2124 32730 2149
rect 32000 2068 32404 2124
rect 32460 2068 32492 2124
rect 32548 2068 32580 2124
rect 32636 2068 32668 2124
rect 32724 2068 32730 2124
rect 32000 2043 32730 2068
rect 32000 1987 32404 2043
rect 32460 1987 32492 2043
rect 32548 1987 32580 2043
rect 32636 1987 32668 2043
rect 32724 1987 32730 2043
rect 32000 1962 32730 1987
rect 32000 1906 32404 1962
rect 32460 1906 32492 1962
rect 32548 1906 32580 1962
rect 32636 1906 32668 1962
rect 32724 1906 32730 1962
rect 32000 1881 32730 1906
rect 32000 1825 32404 1881
rect 32460 1825 32492 1881
rect 32548 1825 32580 1881
rect 32636 1825 32668 1881
rect 32724 1825 32730 1881
rect 32000 1800 32730 1825
rect 32000 1744 32404 1800
rect 32460 1744 32492 1800
rect 32548 1744 32580 1800
rect 32636 1744 32668 1800
rect 32724 1744 32730 1800
rect 32000 1719 32730 1744
rect 32000 1663 32404 1719
rect 32460 1663 32492 1719
rect 32548 1663 32580 1719
rect 32636 1663 32668 1719
rect 32724 1663 32730 1719
rect 32000 1638 32730 1663
rect 725 1595 755 1625
rect 32000 1582 32404 1638
rect 32460 1582 32492 1638
rect 32548 1582 32580 1638
rect 32636 1582 32668 1638
rect 32724 1582 32730 1638
rect 32000 1557 32730 1582
rect 32000 1501 32404 1557
rect 32460 1501 32492 1557
rect 32548 1501 32580 1557
rect 32636 1501 32668 1557
rect 32724 1501 32730 1557
rect 32000 1476 32730 1501
rect 32000 1420 32404 1476
rect 32460 1420 32492 1476
rect 32548 1420 32580 1476
rect 32636 1420 32668 1476
rect 32724 1420 32730 1476
rect 32000 1395 32730 1420
rect 32000 1339 32404 1395
rect 32460 1339 32492 1395
rect 32548 1339 32580 1395
rect 32636 1339 32668 1395
rect 32724 1339 32730 1395
rect 32000 1313 32730 1339
rect 32000 1257 32404 1313
rect 32460 1257 32492 1313
rect 32548 1257 32580 1313
rect 32636 1257 32668 1313
rect 32724 1257 32730 1313
rect 32000 1231 32730 1257
rect 32000 1175 32404 1231
rect 32460 1175 32492 1231
rect 32548 1175 32580 1231
rect 32636 1175 32668 1231
rect 32724 1175 32730 1231
rect 32000 1166 32730 1175
<< metal4 >>
rect 27658 22390 29608 23280
<< metal5 >>
rect 3685 28901 10710 31756
<< glass >>
rect 3685 28901 10710 31756
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 10176 0 1 9195
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 10907 0 1 9204
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 5675 1 0 9099
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 1 0 6019 0 1 9871
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 1 0 4073 0 1 11653
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 1 0 5109 0 1 11653
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 2145 -1 0 5769
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform 0 1 76 -1 0 5770
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 1 0 31407 0 1 40072
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 31593 0 1 39827
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 1 0 2567 0 1 1323
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 1 0 1228 0 1 1323
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1707688321
transform 1 0 1855 0 1 1323
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1707688321
transform 1 0 513 0 1 1323
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1707688321
transform 1 0 18531 0 1 8371
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 4085 1 0 11084
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 0 -1 13375 1 0 7321
box 0 0 1 1
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_0
timestamp 1707688321
transform 1 0 3022 0 1 1195
box 0 0 128 308
use M1M2_CDNS_524688791851176  M1M2_CDNS_524688791851176_0
timestamp 1707688321
transform 1 0 3586 0 1 1195
box 0 0 256 308
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 18531 0 -1 6691
box 0 0 384 116
use M1short_CDNS_524688791851666  M1short_CDNS_524688791851666_0
timestamp 1707688321
transform 1 0 18328 0 1 6480
box 0 0 1 1
use M2M3_CDNS_524688791851174  M2M3_CDNS_524688791851174_0
timestamp 1707688321
transform 1 0 1719 0 1 40257
box -5 0 301 154
use M3M4_CDNS_524688791851178  M3M4_CDNS_524688791851178_0
timestamp 1707688321
transform 0 1 960 1 0 36490
box -1 0 945 476
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1707688321
transform 0 1 18530 -1 0 8423
box 0 0 2270 404
use s8_esd_res250only_small  s8_esd_res250only_small_1
timestamp 1707688321
transform 0 1 -601 -1 0 7001
box 0 0 2270 404
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_0
timestamp 1707688321
transform 1 0 15311 0 1 2525
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_1
timestamp 1707688321
transform 1 0 15693 0 1 1167
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_2
timestamp 1707688321
transform 1 0 26804 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_3
timestamp 1707688321
transform 1 0 27471 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_4
timestamp 1707688321
transform 1 0 25912 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_5
timestamp 1707688321
transform 1 0 24823 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_6
timestamp 1707688321
transform 1 0 21740 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_7
timestamp 1707688321
transform 1 0 23322 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_8
timestamp 1707688321
transform 1 0 22129 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_9
timestamp 1707688321
transform 1 0 19979 0 1 21955
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_10
timestamp 1707688321
transform 1 0 20675 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_11
timestamp 1707688321
transform 1 0 30869 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_12
timestamp 1707688321
transform 1 0 23167 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_13
timestamp 1707688321
transform 1 0 25912 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_14
timestamp 1707688321
transform 1 0 19794 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_15
timestamp 1707688321
transform 1 0 29345 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_16
timestamp 1707688321
transform 1 0 20288 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_17
timestamp 1707688321
transform 1 0 18890 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_18
timestamp 1707688321
transform 1 0 19384 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_19
timestamp 1707688321
transform 1 0 27103 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_20
timestamp 1707688321
transform 1 0 28202 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_21
timestamp 1707688321
transform 1 0 19979 0 1 22943
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_22
timestamp 1707688321
transform 1 0 25006 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_23
timestamp 1707688321
transform 1 0 17330 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_24
timestamp 1707688321
transform 1 0 26900 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_25
timestamp 1707688321
transform 1 0 28696 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_26
timestamp 1707688321
transform 1 0 30248 0 1 3882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_27
timestamp 1707688321
transform 1 0 31379 0 1 3747
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_28
timestamp 1707688321
transform 1 0 30246 0 1 5468
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_29
timestamp 1707688321
transform 1 0 18077 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_30
timestamp 1707688321
transform 1 0 17583 0 1 13467
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_31
timestamp 1707688321
transform 1 0 24924 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_32
timestamp 1707688321
transform 1 0 24430 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_33
timestamp 1707688321
transform 1 0 23755 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_34
timestamp 1707688321
transform 1 0 22407 0 1 6677
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_35
timestamp 1707688321
transform 1 0 28851 0 1 12109
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_36
timestamp 1707688321
transform 1 0 24517 0 1 3917
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_37
timestamp 1707688321
transform 1 0 25011 0 1 3912
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_38
timestamp 1707688321
transform 1 0 23755 0 1 3882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_39
timestamp 1707688321
transform 1 0 22558 0 1 3979
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_40
timestamp 1707688321
transform 1 0 21712 0 1 3924
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_41
timestamp 1707688321
transform 1 0 21239 0 1 3882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_42
timestamp 1707688321
transform 1 0 19954 0 1 3882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_43
timestamp 1707688321
transform 1 0 18581 0 1 5240
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_44
timestamp 1707688321
transform 1 0 18233 0 1 5240
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_45
timestamp 1707688321
transform 1 0 17330 0 1 3882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_46
timestamp 1707688321
transform 1 0 16525 0 1 5240
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_47
timestamp 1707688321
transform 1 0 29199 0 1 6882
box 26 34 340 820
use sky130_fd_io__com_m2m3_strap  sky130_fd_io__com_m2m3_strap_48
timestamp 1707688321
transform 1 0 19979 0 1 20967
box 26 34 340 820
use sky130_fd_io__sio_busses  sky130_fd_io__sio_busses_0
timestamp 1707688321
transform 1 0 15000 0 1 916
box 0 80 17000 23759
use sky130_fd_io__sio_busses  sky130_fd_io__sio_busses_1
timestamp 1707688321
transform 1 0 0 0 1 916
box 0 80 17000 23759
use sky130_fd_io__sio_ctl  sky130_fd_io__sio_ctl_0
timestamp 1707688321
transform 1 0 55 0 1 5613
box -53 -5613 15322 4638
use sky130_fd_io__sio_ipath_tsg4  sky130_fd_io__sio_ipath_tsg4_0
timestamp 1707688321
transform 1 0 -3815 0 1 504
box 3870 -504 36901 13672
use sky130_fd_io__sio_opath  sky130_fd_io__sio_opath_0
timestamp 1707688321
transform 1 0 -423 0 1 8544
box -2893 -1422 34075 42403
use sky130_fd_io__sio_top_pad  sky130_fd_io__sio_top_pad_0
timestamp 1707688321
transform 1 0 0 0 1 916
box 960 24219 14040 39299
<< labels >>
flabel comment s 1572 3253 1572 3253 0 FreeSans 440 0 0 0 lv_net
flabel comment s 7369 10378 7369 10378 0 FreeSans 500 90 0 0 no_jumper_check
flabel comment s 11871 10391 11871 10391 0 FreeSans 500 90 0 0 no_jumper_check
flabel comment s 1788 12553 1788 12553 0 FreeSans 8000 0 0 0 vssd
flabel comment s 1788 11286 1788 11286 0 FreeSans 8000 0 0 0 vccd
flabel comment s -421 5882 -421 5882 0 FreeSans 1600 90 0 0 leaker
flabel comment s 1788 13967 1788 13967 0 FreeSans 8000 0 0 0 vccio
flabel comment s 30461 50597 30461 50597 0 FreeSans 500 0 0 0 li_jumper_ok
flabel comment s 4477 22438 4477 22438 0 FreeSans 440 0 0 0 leaker
flabel comment s 21217 42912 21217 42912 0 FreeSans 1000 0 0 0 switched_power
flabel comment s 1788 16670 1788 16670 0 FreeSans 8000 0 0 0 vssio
flabel comment s 18684 7202 18684 7202 0 FreeSans 1600 90 0 0 leaker
flabel comment s 17353 15424 17353 15424 0 FreeSans 1600 90 0 0 leaker
flabel comment s 23251 32032 23251 32032 3 FreeSans 200 270 0 0 oe_hs_h
flabel comment s 23158 32032 23158 32032 3 FreeSans 200 270 0 0 od_h
flabel comment s 8130 975 8130 975 0 FreeSans 200 90 0 0 ibuf_sel
flabel comment s 5648 955 5648 955 0 FreeSans 200 90 0 0 slow
flabel comment s 10717 1008 10717 1008 0 FreeSans 200 90 0 0 force_h<1>
flabel comment s 10800 1008 10800 1008 0 FreeSans 200 90 0 0 force_h<0>
flabel comment s 11465 1112 11465 1112 0 FreeSans 200 90 0 0 sio_diff_hyst_en
flabel comment s 3892 979 3892 979 0 FreeSans 200 90 0 0 dm<0>
flabel comment s 3975 979 3975 979 0 FreeSans 200 90 0 0 dm<1>
flabel comment s 4409 979 4409 979 0 FreeSans 200 90 0 0 dm<2>
flabel comment s 5727 956 5727 956 0 FreeSans 200 90 0 0 oe_n
flabel comment s 4483 966 4483 966 0 FreeSans 200 90 0 0 od_h
flabel comment s 10882 935 10882 935 0 FreeSans 200 0 0 0 in
flabel comment s 8056 973 8056 973 0 FreeSans 200 90 0 0 hld_h_n
flabel comment s 13267 1031 13267 1031 0 FreeSans 200 90 0 0 force_lovol_h
flabel comment s 13342 1005 13342 1005 0 FreeSans 200 90 0 0 tie_lo_esd
flabel comment s 9544 980 9544 980 0 FreeSans 200 90 0 0 vtrip_sel
flabel comment s 4790 1035 4790 1035 0 FreeSans 200 90 0 0 sio_reg_hifreq
flabel comment s 5209 976 5209 976 0 FreeSans 200 90 0 0 vreg_en
flabel metal1 s 32729 5699 32781 5750 3 FreeSans 520 0 0 0 vinref
port 2 nsew
flabel metal1 s 32247 39897 32301 39943 7 FreeSans 200 0 0 0 refleak_bias
port 3 nsew
flabel metal1 s 32241 40136 32301 40188 7 FreeSans 200 0 0 0 voutref
port 4 nsew
flabel metal1 s 10922 8137 10922 8137 0 FreeSans 1000 0 0 0 sio_diff_hyst_en_h_n
flabel metal1 s 15679 6867 15679 6867 0 FreeSans 1000 0 0 0 sio_diff_hyst_en_h
flabel metal1 s 32271 40162 32271 40162 7 FreeSans 200 0 0 0 voutref
flabel metal5 s 3685 28901 10710 31756 0 FreeSans 3000 0 0 0 pad
port 5 nsew
flabel metal4 s 28852 22697 29186 22968 0 FreeSans 96 0 0 0 vssio_q
port 6 nsew
flabel metal3 s 112 11029 142 11059 3 FreeSans 3000 0 0 0 vccd
port 7 nsew
flabel metal3 s 725 4184 755 4214 3 FreeSans 3000 0 0 0 vssd
port 8 nsew
flabel metal3 s 725 6905 755 6935 3 FreeSans 3000 0 0 0 vssd
port 8 nsew
flabel metal3 s 112 8358 142 8388 3 FreeSans 3000 0 0 0 vddio_q
port 9 nsew
flabel metal3 s 725 9638 755 9668 3 FreeSans 3000 0 0 0 vccd
port 7 nsew
flabel metal3 s 112 22362 142 22392 3 FreeSans 3000 0 0 0 vssio
port 10 nsew
flabel metal3 s 112 13717 142 13747 3 FreeSans 3000 0 0 0 vddio
port 11 nsew
flabel metal3 s 112 12366 142 12396 3 FreeSans 3000 0 0 0 vssd
port 8 nsew
flabel metal3 s 112 16446 142 16476 3 FreeSans 3000 0 0 0 vssio
port 10 nsew
flabel metal3 s 112 19224 142 19254 3 FreeSans 3000 0 0 0 vddio
port 11 nsew
flabel metal3 s 725 2754 755 2784 3 FreeSans 3000 0 0 0 vcchib
port 12 nsew
flabel metal3 s 112 5593 142 5623 3 FreeSans 3000 0 0 0 vddio_q
port 9 nsew
flabel metal3 s 725 1595 755 1625 3 FreeSans 3000 0 0 0 vcchib
port 12 nsew
flabel metal2 s -498 0 -329 80 3 FreeSans 400 90 0 0 pad_a_esd_1_h
port 13 nsew
flabel metal2 s 6665 0 6717 62 3 FreeSans 520 90 0 0 in_h
port 14 nsew
flabel metal2 s 4896 9781 4896 9781 3 FreeSans 1000 90 0 0 hld_i_h_n
flabel metal2 s 1527 9938 1527 9938 3 FreeSans 1000 90 0 0 dm_h<0>
flabel metal2 s 2628 9840 2628 9840 3 FreeSans 1000 90 0 0 dm_h<1>
flabel metal2 s 5741 9137 5741 9137 3 FreeSans 1000 90 0 0 dm_h<2>
flabel metal2 s 1008 9916 1008 9916 3 FreeSans 1000 90 0 0 dm_h_n<0>
flabel metal2 s 2393 9848 2393 9848 3 FreeSans 1000 90 0 0 dm_h_n<1>
flabel metal2 s 5961 9899 5961 9899 3 FreeSans 1000 90 0 0 dm_h_n<2>
flabel metal2 s 9913 5874 9913 5874 3 FreeSans 1000 90 0 0 trip_sel_h
flabel metal2 s 10158 5880 10158 5880 3 FreeSans 1000 90 0 0 trip_sel_h_n
flabel metal2 s 6677 5808 6677 5808 3 FreeSans 1000 90 0 0 ibuf_sel_h
flabel metal2 s 13128 0 13180 75 3 FreeSans 400 90 0 0 tie_lo_esd
port 15 nsew
flabel metal2 s 5623 0 5675 80 3 FreeSans 400 90 0 0 slow
port 16 nsew
flabel metal2 s 17779 0 17949 80 3 FreeSans 400 90 0 0 pad_a_noesd_h
port 17 nsew
flabel metal2 s 17977 0 18146 80 3 FreeSans 400 90 0 0 pad_a_esd_0_h
port 18 nsew
flabel metal2 s 6745 0 6797 75 3 FreeSans 400 90 0 0 in
port 19 nsew
flabel metal2 s 5703 0 5755 75 3 FreeSans 400 90 0 0 oe_n
port 20 nsew
flabel metal2 s 4464 0 4516 75 3 FreeSans 400 90 0 0 enable_h
port 21 nsew
flabel metal2 s 13804 0 13856 75 3 FreeSans 400 90 0 0 inp_dis
port 22 nsew
flabel metal2 s 10855 0 10907 75 0 FreeSans 400 90 0 0 out
port 23 nsew
flabel metal2 s 8111 0 8163 75 3 FreeSans 400 90 0 0 ibuf_sel
port 24 nsew
flabel metal2 s 8031 0 8083 75 3 FreeSans 400 90 0 0 hld_h_n
port 25 nsew
flabel metal2 s 4384 0 4436 75 3 FreeSans 400 90 0 0 dm<2>
port 26 nsew
flabel metal2 s 3950 0 4002 75 3 FreeSans 400 90 0 0 dm<1>
port 27 nsew
flabel metal2 s 3870 0 3922 75 3 FreeSans 400 90 0 0 dm<0>
port 28 nsew
flabel metal2 s 6757 5804 6757 5804 3 FreeSans 1000 90 0 0 ibuf_sel_h_n
flabel metal2 s 9521 0 9573 62 3 FreeSans 400 90 0 0 vtrip_sel
port 29 nsew
flabel metal2 s 5185 0 5237 61 3 FreeSans 400 90 0 0 vreg_en
port 30 nsew
flabel metal2 s 6889 0 6958 75 3 FreeSans 200 90 0 0 hld_ovr
port 31 nsew
<< properties >>
string GDS_END 102516344
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 100633364
string path 814.100 29.150 814.100 55.350 
<< end >>
