magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 0 976 806
<< pmoslvt >>
rect 204 102 304 704
rect 360 102 460 704
rect 516 102 616 704
rect 672 102 772 704
<< pdiff >>
rect 148 692 204 704
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 304 692 360 704
rect 304 658 315 692
rect 349 658 360 692
rect 304 624 360 658
rect 304 590 315 624
rect 349 590 360 624
rect 304 556 360 590
rect 304 522 315 556
rect 349 522 360 556
rect 304 488 360 522
rect 304 454 315 488
rect 349 454 360 488
rect 304 420 360 454
rect 304 386 315 420
rect 349 386 360 420
rect 304 352 360 386
rect 304 318 315 352
rect 349 318 360 352
rect 304 284 360 318
rect 304 250 315 284
rect 349 250 360 284
rect 304 216 360 250
rect 304 182 315 216
rect 349 182 360 216
rect 304 148 360 182
rect 304 114 315 148
rect 349 114 360 148
rect 304 102 360 114
rect 460 692 516 704
rect 460 658 471 692
rect 505 658 516 692
rect 460 624 516 658
rect 460 590 471 624
rect 505 590 516 624
rect 460 556 516 590
rect 460 522 471 556
rect 505 522 516 556
rect 460 488 516 522
rect 460 454 471 488
rect 505 454 516 488
rect 460 420 516 454
rect 460 386 471 420
rect 505 386 516 420
rect 460 352 516 386
rect 460 318 471 352
rect 505 318 516 352
rect 460 284 516 318
rect 460 250 471 284
rect 505 250 516 284
rect 460 216 516 250
rect 460 182 471 216
rect 505 182 516 216
rect 460 148 516 182
rect 460 114 471 148
rect 505 114 516 148
rect 460 102 516 114
rect 616 692 672 704
rect 616 658 627 692
rect 661 658 672 692
rect 616 624 672 658
rect 616 590 627 624
rect 661 590 672 624
rect 616 556 672 590
rect 616 522 627 556
rect 661 522 672 556
rect 616 488 672 522
rect 616 454 627 488
rect 661 454 672 488
rect 616 420 672 454
rect 616 386 627 420
rect 661 386 672 420
rect 616 352 672 386
rect 616 318 627 352
rect 661 318 672 352
rect 616 284 672 318
rect 616 250 627 284
rect 661 250 672 284
rect 616 216 672 250
rect 616 182 627 216
rect 661 182 672 216
rect 616 148 672 182
rect 616 114 627 148
rect 661 114 672 148
rect 616 102 672 114
rect 772 692 828 704
rect 772 658 783 692
rect 817 658 828 692
rect 772 624 828 658
rect 772 590 783 624
rect 817 590 828 624
rect 772 556 828 590
rect 772 522 783 556
rect 817 522 828 556
rect 772 488 828 522
rect 772 454 783 488
rect 817 454 828 488
rect 772 420 828 454
rect 772 386 783 420
rect 817 386 828 420
rect 772 352 828 386
rect 772 318 783 352
rect 817 318 828 352
rect 772 284 828 318
rect 772 250 783 284
rect 817 250 828 284
rect 772 216 828 250
rect 772 182 783 216
rect 817 182 828 216
rect 772 148 828 182
rect 772 114 783 148
rect 817 114 828 148
rect 772 102 828 114
<< pdiffc >>
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 315 658 349 692
rect 315 590 349 624
rect 315 522 349 556
rect 315 454 349 488
rect 315 386 349 420
rect 315 318 349 352
rect 315 250 349 284
rect 315 182 349 216
rect 315 114 349 148
rect 471 658 505 692
rect 471 590 505 624
rect 471 522 505 556
rect 471 454 505 488
rect 471 386 505 420
rect 471 318 505 352
rect 471 250 505 284
rect 471 182 505 216
rect 471 114 505 148
rect 627 658 661 692
rect 627 590 661 624
rect 627 522 661 556
rect 627 454 661 488
rect 627 386 661 420
rect 627 318 661 352
rect 627 250 661 284
rect 627 182 661 216
rect 627 114 661 148
rect 783 658 817 692
rect 783 590 817 624
rect 783 522 817 556
rect 783 454 817 488
rect 783 386 817 420
rect 783 318 817 352
rect 783 250 817 284
rect 783 182 817 216
rect 783 114 817 148
<< nsubdiff >>
rect 36 658 94 704
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 882 658 940 704
rect 882 624 894 658
rect 928 624 940 658
rect 882 590 940 624
rect 882 556 894 590
rect 928 556 940 590
rect 882 522 940 556
rect 882 488 894 522
rect 928 488 940 522
rect 882 454 940 488
rect 882 420 894 454
rect 928 420 940 454
rect 882 386 940 420
rect 882 352 894 386
rect 928 352 940 386
rect 882 318 940 352
rect 882 284 894 318
rect 928 284 940 318
rect 882 250 940 284
rect 882 216 894 250
rect 928 216 940 250
rect 882 182 940 216
rect 882 148 894 182
rect 928 148 940 182
rect 882 102 940 148
<< nsubdiffcont >>
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 894 624 928 658
rect 894 556 928 590
rect 894 488 928 522
rect 894 420 928 454
rect 894 352 928 386
rect 894 284 928 318
rect 894 216 928 250
rect 894 148 928 182
<< poly >>
rect 183 786 793 806
rect 183 752 199 786
rect 233 752 267 786
rect 301 752 335 786
rect 369 752 403 786
rect 437 752 471 786
rect 505 752 539 786
rect 573 752 607 786
rect 641 752 675 786
rect 709 752 743 786
rect 777 752 793 786
rect 183 736 793 752
rect 204 704 304 736
rect 360 704 460 736
rect 516 704 616 736
rect 672 704 772 736
rect 204 70 304 102
rect 360 70 460 102
rect 516 70 616 102
rect 672 70 772 102
rect 183 54 793 70
rect 183 20 199 54
rect 233 20 267 54
rect 301 20 335 54
rect 369 20 403 54
rect 437 20 471 54
rect 505 20 539 54
rect 573 20 607 54
rect 641 20 675 54
rect 709 20 743 54
rect 777 20 793 54
rect 183 0 793 20
<< polycont >>
rect 199 752 233 786
rect 267 752 301 786
rect 335 752 369 786
rect 403 752 437 786
rect 471 752 505 786
rect 539 752 573 786
rect 607 752 641 786
rect 675 752 709 786
rect 743 752 777 786
rect 199 20 233 54
rect 267 20 301 54
rect 335 20 369 54
rect 403 20 437 54
rect 471 20 505 54
rect 539 20 573 54
rect 607 20 641 54
rect 675 20 709 54
rect 743 20 777 54
<< locali >>
rect 233 752 255 786
rect 301 752 327 786
rect 369 752 399 786
rect 437 752 471 786
rect 505 752 539 786
rect 577 752 607 786
rect 649 752 675 786
rect 721 752 743 786
rect 159 692 193 708
rect 48 672 82 674
rect 48 600 82 624
rect 48 528 82 556
rect 48 456 82 488
rect 48 386 82 420
rect 48 318 82 350
rect 48 250 82 278
rect 48 182 82 206
rect 48 132 82 134
rect 159 624 193 638
rect 159 556 193 566
rect 159 488 193 494
rect 159 420 193 422
rect 159 384 193 386
rect 159 312 193 318
rect 159 240 193 250
rect 159 168 193 182
rect 159 98 193 114
rect 315 692 349 708
rect 315 624 349 638
rect 315 556 349 566
rect 315 488 349 494
rect 315 420 349 422
rect 315 384 349 386
rect 315 312 349 318
rect 315 240 349 250
rect 315 168 349 182
rect 315 98 349 114
rect 471 692 505 708
rect 471 624 505 638
rect 471 556 505 566
rect 471 488 505 494
rect 471 420 505 422
rect 471 384 505 386
rect 471 312 505 318
rect 471 240 505 250
rect 471 168 505 182
rect 471 98 505 114
rect 627 692 661 708
rect 627 624 661 638
rect 627 556 661 566
rect 627 488 661 494
rect 627 420 661 422
rect 627 384 661 386
rect 627 312 661 318
rect 627 240 661 250
rect 627 168 661 182
rect 627 98 661 114
rect 783 692 817 708
rect 783 624 817 638
rect 783 556 817 566
rect 783 488 817 494
rect 783 420 817 422
rect 783 384 817 386
rect 783 312 817 318
rect 783 240 817 250
rect 783 168 817 182
rect 894 672 928 674
rect 894 600 928 624
rect 894 528 928 556
rect 894 456 928 488
rect 894 386 928 420
rect 894 318 928 350
rect 894 250 928 278
rect 894 182 928 206
rect 894 132 928 134
rect 783 98 817 114
rect 233 20 255 54
rect 301 20 327 54
rect 369 20 399 54
rect 437 20 471 54
rect 505 20 539 54
rect 577 20 607 54
rect 649 20 675 54
rect 721 20 743 54
<< viali >>
rect 183 752 199 786
rect 199 752 217 786
rect 255 752 267 786
rect 267 752 289 786
rect 327 752 335 786
rect 335 752 361 786
rect 399 752 403 786
rect 403 752 433 786
rect 471 752 505 786
rect 543 752 573 786
rect 573 752 577 786
rect 615 752 641 786
rect 641 752 649 786
rect 687 752 709 786
rect 709 752 721 786
rect 759 752 777 786
rect 777 752 793 786
rect 48 658 82 672
rect 48 638 82 658
rect 48 590 82 600
rect 48 566 82 590
rect 48 522 82 528
rect 48 494 82 522
rect 48 454 82 456
rect 48 422 82 454
rect 48 352 82 384
rect 48 350 82 352
rect 48 284 82 312
rect 48 278 82 284
rect 48 216 82 240
rect 48 206 82 216
rect 48 148 82 168
rect 48 134 82 148
rect 159 658 193 672
rect 159 638 193 658
rect 159 590 193 600
rect 159 566 193 590
rect 159 522 193 528
rect 159 494 193 522
rect 159 454 193 456
rect 159 422 193 454
rect 159 352 193 384
rect 159 350 193 352
rect 159 284 193 312
rect 159 278 193 284
rect 159 216 193 240
rect 159 206 193 216
rect 159 148 193 168
rect 159 134 193 148
rect 315 658 349 672
rect 315 638 349 658
rect 315 590 349 600
rect 315 566 349 590
rect 315 522 349 528
rect 315 494 349 522
rect 315 454 349 456
rect 315 422 349 454
rect 315 352 349 384
rect 315 350 349 352
rect 315 284 349 312
rect 315 278 349 284
rect 315 216 349 240
rect 315 206 349 216
rect 315 148 349 168
rect 315 134 349 148
rect 471 658 505 672
rect 471 638 505 658
rect 471 590 505 600
rect 471 566 505 590
rect 471 522 505 528
rect 471 494 505 522
rect 471 454 505 456
rect 471 422 505 454
rect 471 352 505 384
rect 471 350 505 352
rect 471 284 505 312
rect 471 278 505 284
rect 471 216 505 240
rect 471 206 505 216
rect 471 148 505 168
rect 471 134 505 148
rect 627 658 661 672
rect 627 638 661 658
rect 627 590 661 600
rect 627 566 661 590
rect 627 522 661 528
rect 627 494 661 522
rect 627 454 661 456
rect 627 422 661 454
rect 627 352 661 384
rect 627 350 661 352
rect 627 284 661 312
rect 627 278 661 284
rect 627 216 661 240
rect 627 206 661 216
rect 627 148 661 168
rect 627 134 661 148
rect 783 658 817 672
rect 783 638 817 658
rect 783 590 817 600
rect 783 566 817 590
rect 783 522 817 528
rect 783 494 817 522
rect 783 454 817 456
rect 783 422 817 454
rect 783 352 817 384
rect 783 350 817 352
rect 783 284 817 312
rect 783 278 817 284
rect 783 216 817 240
rect 783 206 817 216
rect 783 148 817 168
rect 783 134 817 148
rect 894 658 928 672
rect 894 638 928 658
rect 894 590 928 600
rect 894 566 928 590
rect 894 522 928 528
rect 894 494 928 522
rect 894 454 928 456
rect 894 422 928 454
rect 894 352 928 384
rect 894 350 928 352
rect 894 284 928 312
rect 894 278 928 284
rect 894 216 928 240
rect 894 206 928 216
rect 894 148 928 168
rect 894 134 928 148
rect 183 20 199 54
rect 199 20 217 54
rect 255 20 267 54
rect 267 20 289 54
rect 327 20 335 54
rect 335 20 361 54
rect 399 20 403 54
rect 403 20 433 54
rect 471 20 505 54
rect 543 20 573 54
rect 573 20 577 54
rect 615 20 641 54
rect 641 20 649 54
rect 687 20 709 54
rect 709 20 721 54
rect 759 20 777 54
rect 777 20 793 54
<< metal1 >>
rect 171 786 805 806
rect 171 752 183 786
rect 217 752 255 786
rect 289 752 327 786
rect 361 752 399 786
rect 433 752 471 786
rect 505 752 543 786
rect 577 752 615 786
rect 649 752 687 786
rect 721 752 759 786
rect 793 752 805 786
rect 171 740 805 752
rect 36 672 94 684
rect 36 638 48 672
rect 82 638 94 672
rect 36 600 94 638
rect 36 566 48 600
rect 82 566 94 600
rect 36 528 94 566
rect 36 494 48 528
rect 82 494 94 528
rect 36 456 94 494
rect 36 422 48 456
rect 82 422 94 456
rect 36 384 94 422
rect 36 350 48 384
rect 82 350 94 384
rect 36 312 94 350
rect 36 278 48 312
rect 82 278 94 312
rect 36 240 94 278
rect 36 206 48 240
rect 82 206 94 240
rect 36 168 94 206
rect 36 134 48 168
rect 82 134 94 168
rect 36 122 94 134
rect 150 672 202 684
rect 150 638 159 672
rect 193 638 202 672
rect 150 600 202 638
rect 150 566 159 600
rect 193 566 202 600
rect 150 528 202 566
rect 150 494 159 528
rect 193 494 202 528
rect 150 456 202 494
rect 150 422 159 456
rect 193 422 202 456
rect 150 384 202 422
rect 150 372 159 384
rect 193 372 202 384
rect 150 312 202 320
rect 150 308 159 312
rect 193 308 202 312
rect 150 244 202 256
rect 150 180 202 192
rect 150 122 202 128
rect 306 678 358 684
rect 306 614 358 626
rect 306 550 358 562
rect 306 494 315 498
rect 349 494 358 498
rect 306 486 358 494
rect 306 422 315 434
rect 349 422 358 434
rect 306 384 358 422
rect 306 350 315 384
rect 349 350 358 384
rect 306 312 358 350
rect 306 278 315 312
rect 349 278 358 312
rect 306 240 358 278
rect 306 206 315 240
rect 349 206 358 240
rect 306 168 358 206
rect 306 134 315 168
rect 349 134 358 168
rect 306 122 358 134
rect 462 672 514 684
rect 462 638 471 672
rect 505 638 514 672
rect 462 600 514 638
rect 462 566 471 600
rect 505 566 514 600
rect 462 528 514 566
rect 462 494 471 528
rect 505 494 514 528
rect 462 456 514 494
rect 462 422 471 456
rect 505 422 514 456
rect 462 384 514 422
rect 462 372 471 384
rect 505 372 514 384
rect 462 312 514 320
rect 462 308 471 312
rect 505 308 514 312
rect 462 244 514 256
rect 462 180 514 192
rect 462 122 514 128
rect 618 678 670 684
rect 618 614 670 626
rect 618 550 670 562
rect 618 494 627 498
rect 661 494 670 498
rect 618 486 670 494
rect 618 422 627 434
rect 661 422 670 434
rect 618 384 670 422
rect 618 350 627 384
rect 661 350 670 384
rect 618 312 670 350
rect 618 278 627 312
rect 661 278 670 312
rect 618 240 670 278
rect 618 206 627 240
rect 661 206 670 240
rect 618 168 670 206
rect 618 134 627 168
rect 661 134 670 168
rect 618 122 670 134
rect 774 672 826 684
rect 774 638 783 672
rect 817 638 826 672
rect 774 600 826 638
rect 774 566 783 600
rect 817 566 826 600
rect 774 528 826 566
rect 774 494 783 528
rect 817 494 826 528
rect 774 456 826 494
rect 774 422 783 456
rect 817 422 826 456
rect 774 384 826 422
rect 774 372 783 384
rect 817 372 826 384
rect 774 312 826 320
rect 774 308 783 312
rect 817 308 826 312
rect 774 244 826 256
rect 774 180 826 192
rect 774 122 826 128
rect 882 672 940 684
rect 882 638 894 672
rect 928 638 940 672
rect 882 600 940 638
rect 882 566 894 600
rect 928 566 940 600
rect 882 528 940 566
rect 882 494 894 528
rect 928 494 940 528
rect 882 456 940 494
rect 882 422 894 456
rect 928 422 940 456
rect 882 384 940 422
rect 882 350 894 384
rect 928 350 940 384
rect 882 312 940 350
rect 882 278 894 312
rect 928 278 940 312
rect 882 240 940 278
rect 882 206 894 240
rect 928 206 940 240
rect 882 168 940 206
rect 882 134 894 168
rect 928 134 940 168
rect 882 122 940 134
rect 171 54 805 66
rect 171 20 183 54
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
rect 793 20 805 54
rect 171 0 805 20
<< via1 >>
rect 150 350 159 372
rect 159 350 193 372
rect 193 350 202 372
rect 150 320 202 350
rect 150 278 159 308
rect 159 278 193 308
rect 193 278 202 308
rect 150 256 202 278
rect 150 240 202 244
rect 150 206 159 240
rect 159 206 193 240
rect 193 206 202 240
rect 150 192 202 206
rect 150 168 202 180
rect 150 134 159 168
rect 159 134 193 168
rect 193 134 202 168
rect 150 128 202 134
rect 306 672 358 678
rect 306 638 315 672
rect 315 638 349 672
rect 349 638 358 672
rect 306 626 358 638
rect 306 600 358 614
rect 306 566 315 600
rect 315 566 349 600
rect 349 566 358 600
rect 306 562 358 566
rect 306 528 358 550
rect 306 498 315 528
rect 315 498 349 528
rect 349 498 358 528
rect 306 456 358 486
rect 306 434 315 456
rect 315 434 349 456
rect 349 434 358 456
rect 462 350 471 372
rect 471 350 505 372
rect 505 350 514 372
rect 462 320 514 350
rect 462 278 471 308
rect 471 278 505 308
rect 505 278 514 308
rect 462 256 514 278
rect 462 240 514 244
rect 462 206 471 240
rect 471 206 505 240
rect 505 206 514 240
rect 462 192 514 206
rect 462 168 514 180
rect 462 134 471 168
rect 471 134 505 168
rect 505 134 514 168
rect 462 128 514 134
rect 618 672 670 678
rect 618 638 627 672
rect 627 638 661 672
rect 661 638 670 672
rect 618 626 670 638
rect 618 600 670 614
rect 618 566 627 600
rect 627 566 661 600
rect 661 566 670 600
rect 618 562 670 566
rect 618 528 670 550
rect 618 498 627 528
rect 627 498 661 528
rect 661 498 670 528
rect 618 456 670 486
rect 618 434 627 456
rect 627 434 661 456
rect 661 434 670 456
rect 774 350 783 372
rect 783 350 817 372
rect 817 350 826 372
rect 774 320 826 350
rect 774 278 783 308
rect 783 278 817 308
rect 817 278 826 308
rect 774 256 826 278
rect 774 240 826 244
rect 774 206 783 240
rect 783 206 817 240
rect 817 206 826 240
rect 774 192 826 206
rect 774 168 826 180
rect 774 134 783 168
rect 783 134 817 168
rect 817 134 826 168
rect 774 128 826 134
<< metal2 >>
rect 10 678 966 684
rect 10 626 306 678
rect 358 626 618 678
rect 670 626 966 678
rect 10 614 966 626
rect 10 562 306 614
rect 358 562 618 614
rect 670 562 966 614
rect 10 550 966 562
rect 10 498 306 550
rect 358 498 618 550
rect 670 498 966 550
rect 10 486 966 498
rect 10 434 306 486
rect 358 434 618 486
rect 670 434 966 486
rect 10 428 966 434
rect 10 372 966 378
rect 10 320 150 372
rect 202 320 462 372
rect 514 320 774 372
rect 826 320 966 372
rect 10 308 966 320
rect 10 256 150 308
rect 202 256 462 308
rect 514 256 774 308
rect 826 256 966 308
rect 10 244 966 256
rect 10 192 150 244
rect 202 192 462 244
rect 514 192 774 244
rect 826 192 966 244
rect 10 180 966 192
rect 10 128 150 180
rect 202 128 462 180
rect 514 128 774 180
rect 826 128 966 180
rect 10 122 966 128
<< labels >>
flabel metal2 s 10 428 30 684 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 122 30 378 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 882 122 940 138 3 FreeSans 300 90 0 0 BULK
port 4 nsew
flabel metal1 s 36 122 94 138 3 FreeSans 300 90 0 0 BULK
port 4 nsew
flabel metal1 s 171 0 805 66 0 FreeSans 300 0 0 0 GATE
port 5 nsew
flabel metal1 s 171 740 805 806 0 FreeSans 300 0 0 0 GATE
port 5 nsew
<< properties >>
string GDS_END 9947904
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9931888
<< end >>
