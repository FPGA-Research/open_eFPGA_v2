magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal3 >>
rect 380 10164 616 10165
rect 711 10164 947 10165
rect 1048 10164 1284 10165
rect 1380 10164 1616 10165
rect 1711 10164 1947 10165
rect 2048 10164 2284 10165
rect 2380 10164 2616 10165
rect 2711 10164 2947 10165
rect 3048 10164 3284 10165
rect 3380 10164 3616 10165
rect 3711 10164 3947 10165
rect 4048 10164 4284 10165
rect 4380 10164 4616 10165
rect 4711 10164 4947 10165
rect 100 9930 4947 10164
rect 380 9929 616 9930
rect 711 9929 947 9930
rect 1048 9929 1284 9930
rect 1380 9929 1616 9930
rect 1711 9929 1947 9930
rect 2048 9929 2284 9930
rect 2380 9929 2616 9930
rect 2711 9929 2947 9930
rect 3048 9929 3284 9930
rect 3380 9929 3616 9930
rect 3711 9929 3947 9930
rect 4048 9929 4284 9930
rect 4380 9929 4616 9930
rect 4711 9929 4947 9930
rect 10048 10164 10284 10165
rect 10380 10164 10616 10165
rect 10711 10164 10947 10165
rect 11048 10164 11284 10165
rect 11380 10164 11616 10165
rect 11711 10164 11947 10165
rect 12048 10164 12284 10165
rect 12380 10164 12616 10165
rect 12711 10164 12947 10165
rect 13048 10164 13284 10165
rect 13380 10164 13616 10165
rect 13711 10164 13947 10165
rect 14048 10164 14284 10165
rect 14380 10164 14616 10165
rect 10048 9930 14931 10164
rect 10048 9929 10284 9930
rect 10380 9929 10616 9930
rect 10711 9929 10947 9930
rect 11048 9929 11284 9930
rect 11380 9929 11616 9930
rect 11711 9929 11947 9930
rect 12048 9929 12284 9930
rect 12380 9929 12616 9930
rect 12711 9929 12947 9930
rect 13048 9929 13284 9930
rect 13380 9929 13616 9930
rect 13711 9929 13947 9930
rect 14048 9929 14284 9930
rect 14380 9929 14616 9930
rect 10151 7593 14931 7636
rect 10111 7357 14931 7593
rect 10151 7227 14931 7357
rect 10111 6991 14931 7227
rect 10151 6948 14931 6991
<< obsm3 >>
rect 100 6948 4880 7636
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 380 9929 616 10165
rect 711 9929 947 10165
rect 1048 9929 1284 10165
rect 1380 9929 1616 10165
rect 1711 9929 1947 10165
rect 2048 9929 2284 10165
rect 2380 9929 2616 10165
rect 2711 9929 2947 10165
rect 3048 9929 3284 10165
rect 3380 9929 3616 10165
rect 3711 9929 3947 10165
rect 4048 9929 4284 10165
rect 4380 9929 4616 10165
rect 4711 9929 4947 10165
rect 10048 9929 10284 10165
rect 10380 9929 10616 10165
rect 10711 9929 10947 10165
rect 11048 9929 11284 10165
rect 11380 9929 11616 10165
rect 11711 9929 11947 10165
rect 12048 9929 12284 10165
rect 12380 9929 12616 10165
rect 12711 9929 12947 10165
rect 13048 9929 13284 10165
rect 13380 9929 13616 10165
rect 13711 9929 13947 10165
rect 14048 9929 14284 10165
rect 14380 9929 14616 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 270 7568 334 7632
rect 352 7568 416 7632
rect 434 7568 498 7632
rect 516 7568 580 7632
rect 598 7568 662 7632
rect 679 7568 743 7632
rect 760 7568 824 7632
rect 841 7568 905 7632
rect 922 7568 986 7632
rect 1003 7568 1067 7632
rect 1084 7568 1148 7632
rect 1165 7568 1229 7632
rect 1246 7568 1310 7632
rect 1327 7568 1391 7632
rect 1408 7568 1472 7632
rect 1489 7568 1553 7632
rect 1570 7568 1634 7632
rect 1651 7568 1715 7632
rect 1732 7568 1796 7632
rect 1813 7568 1877 7632
rect 1894 7568 1958 7632
rect 1975 7568 2039 7632
rect 2056 7568 2120 7632
rect 2137 7568 2201 7632
rect 2218 7568 2282 7632
rect 2299 7568 2363 7632
rect 2380 7568 2444 7632
rect 2461 7568 2525 7632
rect 2542 7568 2606 7632
rect 2623 7568 2687 7632
rect 2704 7568 2768 7632
rect 2785 7568 2849 7632
rect 2866 7568 2930 7632
rect 2947 7568 3011 7632
rect 3028 7568 3092 7632
rect 3109 7568 3173 7632
rect 3190 7568 3254 7632
rect 3271 7568 3335 7632
rect 3352 7568 3416 7632
rect 3433 7568 3497 7632
rect 3514 7568 3578 7632
rect 3595 7568 3659 7632
rect 3676 7568 3740 7632
rect 3757 7568 3821 7632
rect 3838 7568 3902 7632
rect 3919 7568 3983 7632
rect 4000 7568 4064 7632
rect 4081 7568 4145 7632
rect 4162 7568 4226 7632
rect 4243 7568 4307 7632
rect 4324 7568 4388 7632
rect 4405 7568 4469 7632
rect 4486 7568 4550 7632
rect 4567 7568 4631 7632
rect 4648 7568 4712 7632
rect 4729 7568 4793 7632
rect 4810 7568 4874 7632
rect 14746 7593 15000 7637
rect 270 7480 334 7544
rect 352 7480 416 7544
rect 434 7480 498 7544
rect 516 7480 580 7544
rect 598 7480 662 7544
rect 679 7480 743 7544
rect 760 7480 824 7544
rect 841 7480 905 7544
rect 922 7480 986 7544
rect 1003 7480 1067 7544
rect 1084 7480 1148 7544
rect 1165 7480 1229 7544
rect 1246 7480 1310 7544
rect 1327 7480 1391 7544
rect 1408 7480 1472 7544
rect 1489 7480 1553 7544
rect 1570 7480 1634 7544
rect 1651 7480 1715 7544
rect 1732 7480 1796 7544
rect 1813 7480 1877 7544
rect 1894 7480 1958 7544
rect 1975 7480 2039 7544
rect 2056 7480 2120 7544
rect 2137 7480 2201 7544
rect 2218 7480 2282 7544
rect 2299 7480 2363 7544
rect 2380 7480 2444 7544
rect 2461 7480 2525 7544
rect 2542 7480 2606 7544
rect 2623 7480 2687 7544
rect 2704 7480 2768 7544
rect 2785 7480 2849 7544
rect 2866 7480 2930 7544
rect 2947 7480 3011 7544
rect 3028 7480 3092 7544
rect 3109 7480 3173 7544
rect 3190 7480 3254 7544
rect 3271 7480 3335 7544
rect 3352 7480 3416 7544
rect 3433 7480 3497 7544
rect 3514 7480 3578 7544
rect 3595 7480 3659 7544
rect 3676 7480 3740 7544
rect 3757 7480 3821 7544
rect 3838 7480 3902 7544
rect 3919 7480 3983 7544
rect 4000 7480 4064 7544
rect 4081 7480 4145 7544
rect 4162 7480 4226 7544
rect 4243 7480 4307 7544
rect 4324 7480 4388 7544
rect 4405 7480 4469 7544
rect 4486 7480 4550 7544
rect 4567 7480 4631 7544
rect 4648 7480 4712 7544
rect 4729 7480 4793 7544
rect 4810 7480 4874 7544
rect 270 7392 334 7456
rect 352 7392 416 7456
rect 434 7392 498 7456
rect 516 7392 580 7456
rect 598 7392 662 7456
rect 679 7392 743 7456
rect 760 7392 824 7456
rect 841 7392 905 7456
rect 922 7392 986 7456
rect 1003 7392 1067 7456
rect 1084 7392 1148 7456
rect 1165 7392 1229 7456
rect 1246 7392 1310 7456
rect 1327 7392 1391 7456
rect 1408 7392 1472 7456
rect 1489 7392 1553 7456
rect 1570 7392 1634 7456
rect 1651 7392 1715 7456
rect 1732 7392 1796 7456
rect 1813 7392 1877 7456
rect 1894 7392 1958 7456
rect 1975 7392 2039 7456
rect 2056 7392 2120 7456
rect 2137 7392 2201 7456
rect 2218 7392 2282 7456
rect 2299 7392 2363 7456
rect 2380 7392 2444 7456
rect 2461 7392 2525 7456
rect 2542 7392 2606 7456
rect 2623 7392 2687 7456
rect 2704 7392 2768 7456
rect 2785 7392 2849 7456
rect 2866 7392 2930 7456
rect 2947 7392 3011 7456
rect 3028 7392 3092 7456
rect 3109 7392 3173 7456
rect 3190 7392 3254 7456
rect 3271 7392 3335 7456
rect 3352 7392 3416 7456
rect 3433 7392 3497 7456
rect 3514 7392 3578 7456
rect 3595 7392 3659 7456
rect 3676 7392 3740 7456
rect 3757 7392 3821 7456
rect 3838 7392 3902 7456
rect 3919 7392 3983 7456
rect 4000 7392 4064 7456
rect 4081 7392 4145 7456
rect 4162 7392 4226 7456
rect 4243 7392 4307 7456
rect 4324 7392 4388 7456
rect 4405 7392 4469 7456
rect 4486 7392 4550 7456
rect 4567 7392 4631 7456
rect 4648 7392 4712 7456
rect 4729 7392 4793 7456
rect 4810 7392 4874 7456
rect 270 7304 334 7368
rect 352 7304 416 7368
rect 434 7304 498 7368
rect 516 7304 580 7368
rect 598 7304 662 7368
rect 679 7304 743 7368
rect 760 7304 824 7368
rect 841 7304 905 7368
rect 922 7304 986 7368
rect 1003 7304 1067 7368
rect 1084 7304 1148 7368
rect 1165 7304 1229 7368
rect 1246 7304 1310 7368
rect 1327 7304 1391 7368
rect 1408 7304 1472 7368
rect 1489 7304 1553 7368
rect 1570 7304 1634 7368
rect 1651 7304 1715 7368
rect 1732 7304 1796 7368
rect 1813 7304 1877 7368
rect 1894 7304 1958 7368
rect 1975 7304 2039 7368
rect 2056 7304 2120 7368
rect 2137 7304 2201 7368
rect 2218 7304 2282 7368
rect 2299 7304 2363 7368
rect 2380 7304 2444 7368
rect 2461 7304 2525 7368
rect 2542 7304 2606 7368
rect 2623 7304 2687 7368
rect 2704 7304 2768 7368
rect 2785 7304 2849 7368
rect 2866 7304 2930 7368
rect 2947 7304 3011 7368
rect 3028 7304 3092 7368
rect 3109 7304 3173 7368
rect 3190 7304 3254 7368
rect 3271 7304 3335 7368
rect 3352 7304 3416 7368
rect 3433 7304 3497 7368
rect 3514 7304 3578 7368
rect 3595 7304 3659 7368
rect 3676 7304 3740 7368
rect 3757 7304 3821 7368
rect 3838 7304 3902 7368
rect 3919 7304 3983 7368
rect 4000 7304 4064 7368
rect 4081 7304 4145 7368
rect 4162 7304 4226 7368
rect 4243 7304 4307 7368
rect 4324 7304 4388 7368
rect 4405 7304 4469 7368
rect 4486 7304 4550 7368
rect 4567 7304 4631 7368
rect 4648 7304 4712 7368
rect 4729 7304 4793 7368
rect 4810 7304 4874 7368
rect 10111 7357 10347 7593
rect 10432 7357 10668 7593
rect 10753 7357 10989 7593
rect 11074 7357 11310 7593
rect 11395 7357 11631 7593
rect 11716 7357 11952 7593
rect 12037 7357 12273 7593
rect 12358 7357 12594 7593
rect 12679 7357 12915 7593
rect 13000 7357 13236 7593
rect 13321 7357 13557 7593
rect 13642 7357 13878 7593
rect 13963 7357 14199 7593
rect 14284 7357 14520 7593
rect 14605 7357 15000 7593
rect 270 7216 334 7280
rect 352 7216 416 7280
rect 434 7216 498 7280
rect 516 7216 580 7280
rect 598 7216 662 7280
rect 679 7216 743 7280
rect 760 7216 824 7280
rect 841 7216 905 7280
rect 922 7216 986 7280
rect 1003 7216 1067 7280
rect 1084 7216 1148 7280
rect 1165 7216 1229 7280
rect 1246 7216 1310 7280
rect 1327 7216 1391 7280
rect 1408 7216 1472 7280
rect 1489 7216 1553 7280
rect 1570 7216 1634 7280
rect 1651 7216 1715 7280
rect 1732 7216 1796 7280
rect 1813 7216 1877 7280
rect 1894 7216 1958 7280
rect 1975 7216 2039 7280
rect 2056 7216 2120 7280
rect 2137 7216 2201 7280
rect 2218 7216 2282 7280
rect 2299 7216 2363 7280
rect 2380 7216 2444 7280
rect 2461 7216 2525 7280
rect 2542 7216 2606 7280
rect 2623 7216 2687 7280
rect 2704 7216 2768 7280
rect 2785 7216 2849 7280
rect 2866 7216 2930 7280
rect 2947 7216 3011 7280
rect 3028 7216 3092 7280
rect 3109 7216 3173 7280
rect 3190 7216 3254 7280
rect 3271 7216 3335 7280
rect 3352 7216 3416 7280
rect 3433 7216 3497 7280
rect 3514 7216 3578 7280
rect 3595 7216 3659 7280
rect 3676 7216 3740 7280
rect 3757 7216 3821 7280
rect 3838 7216 3902 7280
rect 3919 7216 3983 7280
rect 4000 7216 4064 7280
rect 4081 7216 4145 7280
rect 4162 7216 4226 7280
rect 4243 7216 4307 7280
rect 4324 7216 4388 7280
rect 4405 7216 4469 7280
rect 4486 7216 4550 7280
rect 4567 7216 4631 7280
rect 4648 7216 4712 7280
rect 4729 7216 4793 7280
rect 4810 7216 4874 7280
rect 14746 7227 15000 7357
rect 270 7128 334 7192
rect 352 7128 416 7192
rect 434 7128 498 7192
rect 516 7128 580 7192
rect 598 7128 662 7192
rect 679 7128 743 7192
rect 760 7128 824 7192
rect 841 7128 905 7192
rect 922 7128 986 7192
rect 1003 7128 1067 7192
rect 1084 7128 1148 7192
rect 1165 7128 1229 7192
rect 1246 7128 1310 7192
rect 1327 7128 1391 7192
rect 1408 7128 1472 7192
rect 1489 7128 1553 7192
rect 1570 7128 1634 7192
rect 1651 7128 1715 7192
rect 1732 7128 1796 7192
rect 1813 7128 1877 7192
rect 1894 7128 1958 7192
rect 1975 7128 2039 7192
rect 2056 7128 2120 7192
rect 2137 7128 2201 7192
rect 2218 7128 2282 7192
rect 2299 7128 2363 7192
rect 2380 7128 2444 7192
rect 2461 7128 2525 7192
rect 2542 7128 2606 7192
rect 2623 7128 2687 7192
rect 2704 7128 2768 7192
rect 2785 7128 2849 7192
rect 2866 7128 2930 7192
rect 2947 7128 3011 7192
rect 3028 7128 3092 7192
rect 3109 7128 3173 7192
rect 3190 7128 3254 7192
rect 3271 7128 3335 7192
rect 3352 7128 3416 7192
rect 3433 7128 3497 7192
rect 3514 7128 3578 7192
rect 3595 7128 3659 7192
rect 3676 7128 3740 7192
rect 3757 7128 3821 7192
rect 3838 7128 3902 7192
rect 3919 7128 3983 7192
rect 4000 7128 4064 7192
rect 4081 7128 4145 7192
rect 4162 7128 4226 7192
rect 4243 7128 4307 7192
rect 4324 7128 4388 7192
rect 4405 7128 4469 7192
rect 4486 7128 4550 7192
rect 4567 7128 4631 7192
rect 4648 7128 4712 7192
rect 4729 7128 4793 7192
rect 4810 7128 4874 7192
rect 270 7040 334 7104
rect 352 7040 416 7104
rect 434 7040 498 7104
rect 516 7040 580 7104
rect 598 7040 662 7104
rect 679 7040 743 7104
rect 760 7040 824 7104
rect 841 7040 905 7104
rect 922 7040 986 7104
rect 1003 7040 1067 7104
rect 1084 7040 1148 7104
rect 1165 7040 1229 7104
rect 1246 7040 1310 7104
rect 1327 7040 1391 7104
rect 1408 7040 1472 7104
rect 1489 7040 1553 7104
rect 1570 7040 1634 7104
rect 1651 7040 1715 7104
rect 1732 7040 1796 7104
rect 1813 7040 1877 7104
rect 1894 7040 1958 7104
rect 1975 7040 2039 7104
rect 2056 7040 2120 7104
rect 2137 7040 2201 7104
rect 2218 7040 2282 7104
rect 2299 7040 2363 7104
rect 2380 7040 2444 7104
rect 2461 7040 2525 7104
rect 2542 7040 2606 7104
rect 2623 7040 2687 7104
rect 2704 7040 2768 7104
rect 2785 7040 2849 7104
rect 2866 7040 2930 7104
rect 2947 7040 3011 7104
rect 3028 7040 3092 7104
rect 3109 7040 3173 7104
rect 3190 7040 3254 7104
rect 3271 7040 3335 7104
rect 3352 7040 3416 7104
rect 3433 7040 3497 7104
rect 3514 7040 3578 7104
rect 3595 7040 3659 7104
rect 3676 7040 3740 7104
rect 3757 7040 3821 7104
rect 3838 7040 3902 7104
rect 3919 7040 3983 7104
rect 4000 7040 4064 7104
rect 4081 7040 4145 7104
rect 4162 7040 4226 7104
rect 4243 7040 4307 7104
rect 4324 7040 4388 7104
rect 4405 7040 4469 7104
rect 4486 7040 4550 7104
rect 4567 7040 4631 7104
rect 4648 7040 4712 7104
rect 4729 7040 4793 7104
rect 4810 7040 4874 7104
rect 270 6952 334 7016
rect 352 6952 416 7016
rect 434 6952 498 7016
rect 516 6952 580 7016
rect 598 6952 662 7016
rect 679 6952 743 7016
rect 760 6952 824 7016
rect 841 6952 905 7016
rect 922 6952 986 7016
rect 1003 6952 1067 7016
rect 1084 6952 1148 7016
rect 1165 6952 1229 7016
rect 1246 6952 1310 7016
rect 1327 6952 1391 7016
rect 1408 6952 1472 7016
rect 1489 6952 1553 7016
rect 1570 6952 1634 7016
rect 1651 6952 1715 7016
rect 1732 6952 1796 7016
rect 1813 6952 1877 7016
rect 1894 6952 1958 7016
rect 1975 6952 2039 7016
rect 2056 6952 2120 7016
rect 2137 6952 2201 7016
rect 2218 6952 2282 7016
rect 2299 6952 2363 7016
rect 2380 6952 2444 7016
rect 2461 6952 2525 7016
rect 2542 6952 2606 7016
rect 2623 6952 2687 7016
rect 2704 6952 2768 7016
rect 2785 6952 2849 7016
rect 2866 6952 2930 7016
rect 2947 6952 3011 7016
rect 3028 6952 3092 7016
rect 3109 6952 3173 7016
rect 3190 6952 3254 7016
rect 3271 6952 3335 7016
rect 3352 6952 3416 7016
rect 3433 6952 3497 7016
rect 3514 6952 3578 7016
rect 3595 6952 3659 7016
rect 3676 6952 3740 7016
rect 3757 6952 3821 7016
rect 3838 6952 3902 7016
rect 3919 6952 3983 7016
rect 4000 6952 4064 7016
rect 4081 6952 4145 7016
rect 4162 6952 4226 7016
rect 4243 6952 4307 7016
rect 4324 6952 4388 7016
rect 4405 6952 4469 7016
rect 4486 6952 4550 7016
rect 4567 6952 4631 7016
rect 4648 6952 4712 7016
rect 4729 6952 4793 7016
rect 4810 6952 4874 7016
rect 10111 6991 10347 7227
rect 10432 6991 10668 7227
rect 10753 6991 10989 7227
rect 11074 6991 11310 7227
rect 11395 6991 11631 7227
rect 11716 6991 11952 7227
rect 12037 6991 12273 7227
rect 12358 6991 12594 7227
rect 12679 6991 12915 7227
rect 13000 6991 13236 7227
rect 13321 6991 13557 7227
rect 13642 6991 13878 7227
rect 13963 6991 14199 7227
rect 14284 6991 14520 7227
rect 14605 6991 15000 7227
rect 14746 6947 15000 6991
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 380 10145
rect 616 9949 711 10145
rect 947 9949 1048 10145
rect 1284 9949 1380 10145
rect 1616 9949 1711 10145
rect 1947 9949 2048 10145
rect 2284 9949 2380 10145
rect 2616 9949 2711 10145
rect 2947 9949 3048 10145
rect 3284 9949 3380 10145
rect 3616 9949 3711 10145
rect 3947 9949 4048 10145
rect 4284 9949 4380 10145
rect 4616 9949 4711 10145
rect 4947 9949 10048 10145
rect 10284 9949 10380 10145
rect 10616 9949 10711 10145
rect 10947 9949 11048 10145
rect 11284 9949 11380 10145
rect 11616 9949 11711 10145
rect 11947 9949 12048 10145
rect 12284 9949 12380 10145
rect 12616 9949 12711 10145
rect 12947 9949 13048 10145
rect 13284 9949 13380 10145
rect 13616 9949 13711 10145
rect 13947 9949 14048 10145
rect 14284 9949 14380 10145
rect 14616 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 7632 14666 7717
rect 334 7568 352 7632
rect 416 7568 434 7632
rect 498 7568 516 7632
rect 580 7568 598 7632
rect 662 7568 679 7632
rect 743 7568 760 7632
rect 824 7568 841 7632
rect 905 7568 922 7632
rect 986 7568 1003 7632
rect 1067 7568 1084 7632
rect 1148 7568 1165 7632
rect 1229 7568 1246 7632
rect 1310 7568 1327 7632
rect 1391 7568 1408 7632
rect 1472 7568 1489 7632
rect 1553 7568 1570 7632
rect 1634 7568 1651 7632
rect 1715 7568 1732 7632
rect 1796 7568 1813 7632
rect 1877 7568 1894 7632
rect 1958 7568 1975 7632
rect 2039 7568 2056 7632
rect 2120 7568 2137 7632
rect 2201 7568 2218 7632
rect 2282 7568 2299 7632
rect 2363 7568 2380 7632
rect 2444 7568 2461 7632
rect 2525 7568 2542 7632
rect 2606 7568 2623 7632
rect 2687 7568 2704 7632
rect 2768 7568 2785 7632
rect 2849 7568 2866 7632
rect 2930 7568 2947 7632
rect 3011 7568 3028 7632
rect 3092 7568 3109 7632
rect 3173 7568 3190 7632
rect 3254 7568 3271 7632
rect 3335 7568 3352 7632
rect 3416 7568 3433 7632
rect 3497 7568 3514 7632
rect 3578 7568 3595 7632
rect 3659 7568 3676 7632
rect 3740 7568 3757 7632
rect 3821 7568 3838 7632
rect 3902 7568 3919 7632
rect 3983 7568 4000 7632
rect 4064 7568 4081 7632
rect 4145 7568 4162 7632
rect 4226 7568 4243 7632
rect 4307 7568 4324 7632
rect 4388 7568 4405 7632
rect 4469 7568 4486 7632
rect 4550 7568 4567 7632
rect 4631 7568 4648 7632
rect 4712 7568 4729 7632
rect 4793 7568 4810 7632
rect 4874 7593 14666 7632
rect 4874 7568 10111 7593
rect 334 7544 10111 7568
rect 334 7480 352 7544
rect 416 7480 434 7544
rect 498 7480 516 7544
rect 580 7480 598 7544
rect 662 7480 679 7544
rect 743 7480 760 7544
rect 824 7480 841 7544
rect 905 7480 922 7544
rect 986 7480 1003 7544
rect 1067 7480 1084 7544
rect 1148 7480 1165 7544
rect 1229 7480 1246 7544
rect 1310 7480 1327 7544
rect 1391 7480 1408 7544
rect 1472 7480 1489 7544
rect 1553 7480 1570 7544
rect 1634 7480 1651 7544
rect 1715 7480 1732 7544
rect 1796 7480 1813 7544
rect 1877 7480 1894 7544
rect 1958 7480 1975 7544
rect 2039 7480 2056 7544
rect 2120 7480 2137 7544
rect 2201 7480 2218 7544
rect 2282 7480 2299 7544
rect 2363 7480 2380 7544
rect 2444 7480 2461 7544
rect 2525 7480 2542 7544
rect 2606 7480 2623 7544
rect 2687 7480 2704 7544
rect 2768 7480 2785 7544
rect 2849 7480 2866 7544
rect 2930 7480 2947 7544
rect 3011 7480 3028 7544
rect 3092 7480 3109 7544
rect 3173 7480 3190 7544
rect 3254 7480 3271 7544
rect 3335 7480 3352 7544
rect 3416 7480 3433 7544
rect 3497 7480 3514 7544
rect 3578 7480 3595 7544
rect 3659 7480 3676 7544
rect 3740 7480 3757 7544
rect 3821 7480 3838 7544
rect 3902 7480 3919 7544
rect 3983 7480 4000 7544
rect 4064 7480 4081 7544
rect 4145 7480 4162 7544
rect 4226 7480 4243 7544
rect 4307 7480 4324 7544
rect 4388 7480 4405 7544
rect 4469 7480 4486 7544
rect 4550 7480 4567 7544
rect 4631 7480 4648 7544
rect 4712 7480 4729 7544
rect 4793 7480 4810 7544
rect 4874 7480 10111 7544
rect 334 7456 10111 7480
rect 334 7392 352 7456
rect 416 7392 434 7456
rect 498 7392 516 7456
rect 580 7392 598 7456
rect 662 7392 679 7456
rect 743 7392 760 7456
rect 824 7392 841 7456
rect 905 7392 922 7456
rect 986 7392 1003 7456
rect 1067 7392 1084 7456
rect 1148 7392 1165 7456
rect 1229 7392 1246 7456
rect 1310 7392 1327 7456
rect 1391 7392 1408 7456
rect 1472 7392 1489 7456
rect 1553 7392 1570 7456
rect 1634 7392 1651 7456
rect 1715 7392 1732 7456
rect 1796 7392 1813 7456
rect 1877 7392 1894 7456
rect 1958 7392 1975 7456
rect 2039 7392 2056 7456
rect 2120 7392 2137 7456
rect 2201 7392 2218 7456
rect 2282 7392 2299 7456
rect 2363 7392 2380 7456
rect 2444 7392 2461 7456
rect 2525 7392 2542 7456
rect 2606 7392 2623 7456
rect 2687 7392 2704 7456
rect 2768 7392 2785 7456
rect 2849 7392 2866 7456
rect 2930 7392 2947 7456
rect 3011 7392 3028 7456
rect 3092 7392 3109 7456
rect 3173 7392 3190 7456
rect 3254 7392 3271 7456
rect 3335 7392 3352 7456
rect 3416 7392 3433 7456
rect 3497 7392 3514 7456
rect 3578 7392 3595 7456
rect 3659 7392 3676 7456
rect 3740 7392 3757 7456
rect 3821 7392 3838 7456
rect 3902 7392 3919 7456
rect 3983 7392 4000 7456
rect 4064 7392 4081 7456
rect 4145 7392 4162 7456
rect 4226 7392 4243 7456
rect 4307 7392 4324 7456
rect 4388 7392 4405 7456
rect 4469 7392 4486 7456
rect 4550 7392 4567 7456
rect 4631 7392 4648 7456
rect 4712 7392 4729 7456
rect 4793 7392 4810 7456
rect 4874 7392 10111 7456
rect 334 7368 10111 7392
rect 334 7304 352 7368
rect 416 7304 434 7368
rect 498 7304 516 7368
rect 580 7304 598 7368
rect 662 7304 679 7368
rect 743 7304 760 7368
rect 824 7304 841 7368
rect 905 7304 922 7368
rect 986 7304 1003 7368
rect 1067 7304 1084 7368
rect 1148 7304 1165 7368
rect 1229 7304 1246 7368
rect 1310 7304 1327 7368
rect 1391 7304 1408 7368
rect 1472 7304 1489 7368
rect 1553 7304 1570 7368
rect 1634 7304 1651 7368
rect 1715 7304 1732 7368
rect 1796 7304 1813 7368
rect 1877 7304 1894 7368
rect 1958 7304 1975 7368
rect 2039 7304 2056 7368
rect 2120 7304 2137 7368
rect 2201 7304 2218 7368
rect 2282 7304 2299 7368
rect 2363 7304 2380 7368
rect 2444 7304 2461 7368
rect 2525 7304 2542 7368
rect 2606 7304 2623 7368
rect 2687 7304 2704 7368
rect 2768 7304 2785 7368
rect 2849 7304 2866 7368
rect 2930 7304 2947 7368
rect 3011 7304 3028 7368
rect 3092 7304 3109 7368
rect 3173 7304 3190 7368
rect 3254 7304 3271 7368
rect 3335 7304 3352 7368
rect 3416 7304 3433 7368
rect 3497 7304 3514 7368
rect 3578 7304 3595 7368
rect 3659 7304 3676 7368
rect 3740 7304 3757 7368
rect 3821 7304 3838 7368
rect 3902 7304 3919 7368
rect 3983 7304 4000 7368
rect 4064 7304 4081 7368
rect 4145 7304 4162 7368
rect 4226 7304 4243 7368
rect 4307 7304 4324 7368
rect 4388 7304 4405 7368
rect 4469 7304 4486 7368
rect 4550 7304 4567 7368
rect 4631 7304 4648 7368
rect 4712 7304 4729 7368
rect 4793 7304 4810 7368
rect 4874 7357 10111 7368
rect 10347 7357 10432 7593
rect 10668 7357 10753 7593
rect 10989 7357 11074 7593
rect 11310 7357 11395 7593
rect 11631 7357 11716 7593
rect 11952 7357 12037 7593
rect 12273 7357 12358 7593
rect 12594 7357 12679 7593
rect 12915 7357 13000 7593
rect 13236 7357 13321 7593
rect 13557 7357 13642 7593
rect 13878 7357 13963 7593
rect 14199 7357 14284 7593
rect 14520 7357 14605 7593
rect 4874 7304 14666 7357
rect 334 7280 14666 7304
rect 334 7216 352 7280
rect 416 7216 434 7280
rect 498 7216 516 7280
rect 580 7216 598 7280
rect 662 7216 679 7280
rect 743 7216 760 7280
rect 824 7216 841 7280
rect 905 7216 922 7280
rect 986 7216 1003 7280
rect 1067 7216 1084 7280
rect 1148 7216 1165 7280
rect 1229 7216 1246 7280
rect 1310 7216 1327 7280
rect 1391 7216 1408 7280
rect 1472 7216 1489 7280
rect 1553 7216 1570 7280
rect 1634 7216 1651 7280
rect 1715 7216 1732 7280
rect 1796 7216 1813 7280
rect 1877 7216 1894 7280
rect 1958 7216 1975 7280
rect 2039 7216 2056 7280
rect 2120 7216 2137 7280
rect 2201 7216 2218 7280
rect 2282 7216 2299 7280
rect 2363 7216 2380 7280
rect 2444 7216 2461 7280
rect 2525 7216 2542 7280
rect 2606 7216 2623 7280
rect 2687 7216 2704 7280
rect 2768 7216 2785 7280
rect 2849 7216 2866 7280
rect 2930 7216 2947 7280
rect 3011 7216 3028 7280
rect 3092 7216 3109 7280
rect 3173 7216 3190 7280
rect 3254 7216 3271 7280
rect 3335 7216 3352 7280
rect 3416 7216 3433 7280
rect 3497 7216 3514 7280
rect 3578 7216 3595 7280
rect 3659 7216 3676 7280
rect 3740 7216 3757 7280
rect 3821 7216 3838 7280
rect 3902 7216 3919 7280
rect 3983 7216 4000 7280
rect 4064 7216 4081 7280
rect 4145 7216 4162 7280
rect 4226 7216 4243 7280
rect 4307 7216 4324 7280
rect 4388 7216 4405 7280
rect 4469 7216 4486 7280
rect 4550 7216 4567 7280
rect 4631 7216 4648 7280
rect 4712 7216 4729 7280
rect 4793 7216 4810 7280
rect 4874 7227 14666 7280
rect 4874 7216 10111 7227
rect 334 7192 10111 7216
rect 334 7128 352 7192
rect 416 7128 434 7192
rect 498 7128 516 7192
rect 580 7128 598 7192
rect 662 7128 679 7192
rect 743 7128 760 7192
rect 824 7128 841 7192
rect 905 7128 922 7192
rect 986 7128 1003 7192
rect 1067 7128 1084 7192
rect 1148 7128 1165 7192
rect 1229 7128 1246 7192
rect 1310 7128 1327 7192
rect 1391 7128 1408 7192
rect 1472 7128 1489 7192
rect 1553 7128 1570 7192
rect 1634 7128 1651 7192
rect 1715 7128 1732 7192
rect 1796 7128 1813 7192
rect 1877 7128 1894 7192
rect 1958 7128 1975 7192
rect 2039 7128 2056 7192
rect 2120 7128 2137 7192
rect 2201 7128 2218 7192
rect 2282 7128 2299 7192
rect 2363 7128 2380 7192
rect 2444 7128 2461 7192
rect 2525 7128 2542 7192
rect 2606 7128 2623 7192
rect 2687 7128 2704 7192
rect 2768 7128 2785 7192
rect 2849 7128 2866 7192
rect 2930 7128 2947 7192
rect 3011 7128 3028 7192
rect 3092 7128 3109 7192
rect 3173 7128 3190 7192
rect 3254 7128 3271 7192
rect 3335 7128 3352 7192
rect 3416 7128 3433 7192
rect 3497 7128 3514 7192
rect 3578 7128 3595 7192
rect 3659 7128 3676 7192
rect 3740 7128 3757 7192
rect 3821 7128 3838 7192
rect 3902 7128 3919 7192
rect 3983 7128 4000 7192
rect 4064 7128 4081 7192
rect 4145 7128 4162 7192
rect 4226 7128 4243 7192
rect 4307 7128 4324 7192
rect 4388 7128 4405 7192
rect 4469 7128 4486 7192
rect 4550 7128 4567 7192
rect 4631 7128 4648 7192
rect 4712 7128 4729 7192
rect 4793 7128 4810 7192
rect 4874 7128 10111 7192
rect 334 7104 10111 7128
rect 334 7040 352 7104
rect 416 7040 434 7104
rect 498 7040 516 7104
rect 580 7040 598 7104
rect 662 7040 679 7104
rect 743 7040 760 7104
rect 824 7040 841 7104
rect 905 7040 922 7104
rect 986 7040 1003 7104
rect 1067 7040 1084 7104
rect 1148 7040 1165 7104
rect 1229 7040 1246 7104
rect 1310 7040 1327 7104
rect 1391 7040 1408 7104
rect 1472 7040 1489 7104
rect 1553 7040 1570 7104
rect 1634 7040 1651 7104
rect 1715 7040 1732 7104
rect 1796 7040 1813 7104
rect 1877 7040 1894 7104
rect 1958 7040 1975 7104
rect 2039 7040 2056 7104
rect 2120 7040 2137 7104
rect 2201 7040 2218 7104
rect 2282 7040 2299 7104
rect 2363 7040 2380 7104
rect 2444 7040 2461 7104
rect 2525 7040 2542 7104
rect 2606 7040 2623 7104
rect 2687 7040 2704 7104
rect 2768 7040 2785 7104
rect 2849 7040 2866 7104
rect 2930 7040 2947 7104
rect 3011 7040 3028 7104
rect 3092 7040 3109 7104
rect 3173 7040 3190 7104
rect 3254 7040 3271 7104
rect 3335 7040 3352 7104
rect 3416 7040 3433 7104
rect 3497 7040 3514 7104
rect 3578 7040 3595 7104
rect 3659 7040 3676 7104
rect 3740 7040 3757 7104
rect 3821 7040 3838 7104
rect 3902 7040 3919 7104
rect 3983 7040 4000 7104
rect 4064 7040 4081 7104
rect 4145 7040 4162 7104
rect 4226 7040 4243 7104
rect 4307 7040 4324 7104
rect 4388 7040 4405 7104
rect 4469 7040 4486 7104
rect 4550 7040 4567 7104
rect 4631 7040 4648 7104
rect 4712 7040 4729 7104
rect 4793 7040 4810 7104
rect 4874 7040 10111 7104
rect 334 7016 10111 7040
rect 334 6952 352 7016
rect 416 6952 434 7016
rect 498 6952 516 7016
rect 580 6952 598 7016
rect 662 6952 679 7016
rect 743 6952 760 7016
rect 824 6952 841 7016
rect 905 6952 922 7016
rect 986 6952 1003 7016
rect 1067 6952 1084 7016
rect 1148 6952 1165 7016
rect 1229 6952 1246 7016
rect 1310 6952 1327 7016
rect 1391 6952 1408 7016
rect 1472 6952 1489 7016
rect 1553 6952 1570 7016
rect 1634 6952 1651 7016
rect 1715 6952 1732 7016
rect 1796 6952 1813 7016
rect 1877 6952 1894 7016
rect 1958 6952 1975 7016
rect 2039 6952 2056 7016
rect 2120 6952 2137 7016
rect 2201 6952 2218 7016
rect 2282 6952 2299 7016
rect 2363 6952 2380 7016
rect 2444 6952 2461 7016
rect 2525 6952 2542 7016
rect 2606 6952 2623 7016
rect 2687 6952 2704 7016
rect 2768 6952 2785 7016
rect 2849 6952 2866 7016
rect 2930 6952 2947 7016
rect 3011 6952 3028 7016
rect 3092 6952 3109 7016
rect 3173 6952 3190 7016
rect 3254 6952 3271 7016
rect 3335 6952 3352 7016
rect 3416 6952 3433 7016
rect 3497 6952 3514 7016
rect 3578 6952 3595 7016
rect 3659 6952 3676 7016
rect 3740 6952 3757 7016
rect 3821 6952 3838 7016
rect 3902 6952 3919 7016
rect 3983 6952 4000 7016
rect 4064 6952 4081 7016
rect 4145 6952 4162 7016
rect 4226 6952 4243 7016
rect 4307 6952 4324 7016
rect 4388 6952 4405 7016
rect 4469 6952 4486 7016
rect 4550 6952 4567 7016
rect 4631 6952 4648 7016
rect 4712 6952 4729 7016
rect 4793 6952 4810 7016
rect 4874 6991 10111 7016
rect 10347 6991 10432 7227
rect 10668 6991 10753 7227
rect 10989 6991 11074 7227
rect 11310 6991 11395 7227
rect 11631 6991 11716 7227
rect 11952 6991 12037 7227
rect 12273 6991 12358 7227
rect 12594 6991 12679 7227
rect 12915 6991 13000 7227
rect 13236 6991 13321 7227
rect 13557 6991 13642 7227
rect 13878 6991 13963 7227
rect 14199 6991 14284 7227
rect 14520 6991 14605 7227
rect 4874 6952 14666 6991
rect 334 6867 14666 6952
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 380 9929 616 10165
rect 711 9929 947 10165
rect 1048 9929 1284 10165
rect 1380 9929 1616 10165
rect 1711 9929 1947 10165
rect 2048 9929 2284 10165
rect 2380 9929 2616 10165
rect 2711 9929 2947 10165
rect 3048 9929 3284 10165
rect 3380 9929 3616 10165
rect 3711 9929 3947 10165
rect 4048 9929 4284 10165
rect 4380 9929 4616 10165
rect 4711 9929 4947 10165
rect 10048 9929 10284 10165
rect 10380 9929 10616 10165
rect 10711 9929 10947 10165
rect 11048 9929 11284 10165
rect 11380 9929 11616 10165
rect 11711 9929 11947 10165
rect 12048 9929 12284 10165
rect 12380 9929 12616 10165
rect 12711 9929 12947 10165
rect 13048 9929 13284 10165
rect 13380 9929 13616 10165
rect 13711 9929 13947 10165
rect 14048 9929 14284 10165
rect 14380 9929 14616 10165
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 7593 15000 7617
rect 10111 7357 10347 7593
rect 10432 7357 10668 7593
rect 10753 7357 10989 7593
rect 11074 7357 11310 7593
rect 11395 7357 11631 7593
rect 11716 7357 11952 7593
rect 12037 7357 12273 7593
rect 12358 7357 12594 7593
rect 12679 7357 12915 7593
rect 13000 7357 13236 7593
rect 13321 7357 13557 7593
rect 13642 7357 13878 7593
rect 13963 7357 14199 7593
rect 14284 7357 14520 7593
rect 14605 7357 15000 7593
rect 14746 7227 15000 7357
rect 10111 6991 10347 7227
rect 10432 6991 10668 7227
rect 10753 6991 10989 7227
rect 11074 6991 11310 7227
rect 11395 6991 11631 7227
rect 11716 6991 11952 7227
rect 12037 6991 12273 7227
rect 12358 6991 12594 7227
rect 12679 6991 12915 7227
rect 13000 6991 13236 7227
rect 13321 6991 13557 7227
rect 13642 6991 13878 7227
rect 13963 6991 14199 7227
rect 14284 6991 14520 7227
rect 14605 6991 15000 7227
rect 14746 6968 15000 6991
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 10165 14426 18917
rect 616 9929 711 10165
rect 947 9929 1048 10165
rect 1284 9929 1380 10165
rect 1616 9929 1711 10165
rect 1947 9929 2048 10165
rect 2284 9929 2380 10165
rect 2616 9929 2711 10165
rect 2947 9929 3048 10165
rect 3284 9929 3380 10165
rect 3616 9929 3711 10165
rect 3947 9929 4048 10165
rect 4284 9929 4380 10165
rect 4616 9929 4711 10165
rect 4947 9929 10048 10165
rect 10284 9929 10380 10165
rect 10616 9929 10711 10165
rect 10947 9929 11048 10165
rect 11284 9929 11380 10165
rect 11616 9929 11711 10165
rect 11947 9929 12048 10165
rect 12284 9929 12380 10165
rect 12616 9929 12711 10165
rect 12947 9929 13048 10165
rect 13284 9929 13380 10165
rect 13616 9929 13711 10165
rect 13947 9929 14048 10165
rect 14284 9929 14380 10165
rect 574 7593 14426 9929
rect 574 7357 10111 7593
rect 10347 7357 10432 7593
rect 10668 7357 10753 7593
rect 10989 7357 11074 7593
rect 11310 7357 11395 7593
rect 11631 7357 11716 7593
rect 11952 7357 12037 7593
rect 12273 7357 12358 7593
rect 12594 7357 12679 7593
rect 12915 7357 13000 7593
rect 13236 7357 13321 7593
rect 13557 7357 13642 7593
rect 13878 7357 13963 7593
rect 14199 7357 14284 7593
rect 574 7227 14426 7357
rect 574 6991 10111 7227
rect 10347 6991 10432 7227
rect 10668 6991 10753 7227
rect 10989 6991 11074 7227
rect 11310 6991 11395 7227
rect 11631 6991 11716 7227
rect 11952 6991 12037 7227
rect 12273 6991 12358 7227
rect 12594 6991 12679 7227
rect 12915 6991 13000 7227
rect 13236 6991 13321 7227
rect 13557 6991 13642 7227
rect 13878 6991 13963 7227
rect 14199 6991 14284 7227
rect 574 6968 14426 6991
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 2 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 2 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 2 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 2 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 3 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 3 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 3 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 100 9930 4880 10164 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10151 6948 14931 7636 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10151 9930 14931 10164 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 10111 14913 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 10027 14913 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 9943 14913 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7580 14913 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7492 14913 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7404 14913 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7316 14913 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7228 14913 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7140 14913 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 7052 14913 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14873 6964 14913 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 10111 14832 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 10027 14832 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 9943 14832 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7580 14832 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7492 14832 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7404 14832 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7316 14832 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7228 14832 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7140 14832 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 7052 14832 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14792 6964 14832 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 10111 14751 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 10027 14751 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 9943 14751 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7580 14751 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7492 14751 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7404 14751 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7316 14751 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7228 14751 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7140 14751 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 7052 14751 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14711 6964 14751 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 10111 14670 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 10027 14670 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 9943 14670 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 7580 14670 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14605 7357 14746 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14605 7357 14746 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14605 7357 14746 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 7316 14670 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14630 7228 14670 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14605 6991 14746 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14605 6991 14746 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14605 6991 14746 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14380 9929 14616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14380 9929 14616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14380 9929 14616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7580 14589 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7492 14589 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7404 14589 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7316 14589 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7228 14589 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7140 14589 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 7052 14589 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14549 6964 14589 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14468 7580 14508 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14284 7357 14520 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14284 7357 14520 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14284 7357 14520 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14468 7316 14508 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14468 7228 14508 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14284 6991 14520 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14284 6991 14520 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14284 6991 14520 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14387 7316 14427 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14387 7228 14427 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14306 10111 14346 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14306 10027 14346 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14306 9943 14346 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14306 7316 14346 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14306 7228 14346 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14048 9929 14284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 14048 9929 14284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14048 9929 14284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7580 14265 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7492 14265 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7404 14265 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7316 14265 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7228 14265 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7140 14265 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 7052 14265 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14225 6964 14265 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14144 7580 14184 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13963 7357 14199 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13963 7357 14199 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13963 7357 14199 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14144 7316 14184 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14144 7228 14184 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13963 6991 14199 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13963 6991 14199 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13963 6991 14199 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14063 7316 14103 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 14063 7228 14103 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13982 10111 14022 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13982 10027 14022 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13982 9943 14022 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13982 7316 14022 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13982 7228 14022 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13711 9929 13947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13711 9929 13947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13711 9929 13947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7580 13941 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7492 13941 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7404 13941 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7316 13941 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7228 13941 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7140 13941 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 7052 13941 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13901 6964 13941 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13820 7580 13860 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13642 7357 13878 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13642 7357 13878 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13642 7357 13878 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13820 7316 13860 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13820 7228 13860 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13642 6991 13878 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13642 6991 13878 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13642 6991 13878 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13739 7316 13779 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13739 7228 13779 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13658 10111 13698 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13658 10027 13698 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13658 9943 13698 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13658 7316 13698 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13658 7228 13698 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 10111 13617 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 10027 13617 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 9943 13617 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7580 13617 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7492 13617 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7404 13617 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7316 13617 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7228 13617 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7140 13617 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 7052 13617 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13577 6964 13617 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13380 9929 13616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13380 9929 13616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13380 9929 13616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13496 7580 13536 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13321 7357 13557 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13321 7357 13557 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13321 7357 13557 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13496 7316 13536 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13496 7228 13536 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13321 6991 13557 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13321 6991 13557 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13321 6991 13557 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13415 7316 13455 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13415 7228 13455 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13334 10111 13374 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13334 10027 13374 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13334 9943 13374 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13334 7316 13374 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13334 7228 13374 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 10111 13293 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 10027 13293 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 9943 13293 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7580 13293 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7492 13293 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7404 13293 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7316 13293 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7228 13293 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7140 13293 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 7052 13293 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13253 6964 13293 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13048 9929 13284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13048 9929 13284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13048 9929 13284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13172 7580 13212 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13000 7357 13236 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13000 7357 13236 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13000 7357 13236 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13172 7316 13212 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13172 7228 13212 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 13000 6991 13236 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 13000 6991 13236 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13000 6991 13236 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13091 7316 13131 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13091 7228 13131 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13010 7316 13050 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 13010 7228 13050 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 10111 12969 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 10027 12969 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 9943 12969 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7580 12969 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7492 12969 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7404 12969 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7316 12969 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7228 12969 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7140 12969 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 7052 12969 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12929 6964 12969 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12711 9929 12947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12711 9929 12947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12711 9929 12947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12848 7580 12888 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12679 7357 12915 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12679 7357 12915 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12679 7357 12915 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12848 7316 12888 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12848 7228 12888 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12679 6991 12915 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12679 6991 12915 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12679 6991 12915 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12767 7316 12807 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12767 7228 12807 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12686 7316 12726 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12686 7228 12726 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 10111 12645 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 10027 12645 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 9943 12645 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7580 12645 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7492 12645 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7404 12645 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7316 12645 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7228 12645 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7140 12645 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 7052 12645 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12605 6964 12645 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12380 9929 12616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12380 9929 12616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12380 9929 12616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12524 7580 12564 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12358 7357 12594 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12358 7357 12594 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12358 7357 12594 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12524 7316 12564 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12524 7228 12564 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12358 6991 12594 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12358 6991 12594 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12358 6991 12594 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12443 7316 12483 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12443 7228 12483 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12362 7316 12402 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12362 7228 12402 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 10111 12321 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 10027 12321 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 9943 12321 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7580 12321 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7492 12321 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7404 12321 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7316 12321 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7228 12321 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7140 12321 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 7052 12321 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12281 6964 12321 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12048 9929 12284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12048 9929 12284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12048 9929 12284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12200 7580 12240 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12037 7357 12273 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12037 7357 12273 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12037 7357 12273 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12200 7316 12240 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12200 7228 12240 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 12037 6991 12273 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 12037 6991 12273 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12037 6991 12273 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12119 7316 12159 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12119 7228 12159 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12038 7316 12078 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 12038 7228 12078 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 10111 11997 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 10027 11997 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 9943 11997 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7580 11997 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7492 11997 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7404 11997 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7316 11997 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7228 11997 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7140 11997 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 7052 11997 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11957 6964 11997 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11711 9929 11947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11711 9929 11947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11711 9929 11947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11876 7580 11916 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11716 7357 11952 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11716 7357 11952 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11716 7357 11952 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11876 7316 11916 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11876 7228 11916 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11716 6991 11952 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11716 6991 11952 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11716 6991 11952 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11795 7316 11835 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11795 7228 11835 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11714 7316 11754 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11714 7228 11754 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 10111 11673 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 10027 11673 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 9943 11673 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7580 11673 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7492 11673 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7404 11673 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7316 11673 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7228 11673 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7140 11673 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 7052 11673 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11633 6964 11673 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11380 9929 11616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11380 9929 11616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11380 9929 11616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11552 7580 11592 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11395 7357 11631 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11395 7357 11631 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11395 7357 11631 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11552 7316 11592 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11552 7228 11592 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11395 6991 11631 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11395 6991 11631 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11395 6991 11631 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11471 7316 11511 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11471 7228 11511 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11390 7316 11430 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11390 7228 11430 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 10111 11349 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 10027 11349 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 9943 11349 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7580 11349 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7492 11349 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7404 11349 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7316 11349 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7228 11349 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7140 11349 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 7052 11349 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11309 6964 11349 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11048 9929 11284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11048 9929 11284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11048 9929 11284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11228 7580 11268 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11074 7357 11310 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11074 7357 11310 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11074 7357 11310 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11228 7316 11268 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11228 7228 11268 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 11074 6991 11310 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 11074 6991 11310 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11074 6991 11310 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11147 7316 11187 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11147 7228 11187 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11066 7316 11106 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 11066 7228 11106 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 10111 11025 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 10027 11025 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 9943 11025 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7580 11025 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7492 11025 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7404 11025 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7316 11025 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7228 11025 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7140 11025 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 7052 11025 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10985 6964 11025 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10711 9929 10947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10711 9929 10947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10711 9929 10947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10904 7580 10944 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10753 7357 10989 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10753 7357 10989 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10753 7357 10989 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10904 7316 10944 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10904 7228 10944 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10753 6991 10989 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10753 6991 10989 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10753 6991 10989 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10823 7316 10863 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10823 7228 10863 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10742 7316 10782 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10742 7228 10782 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 10111 10701 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 10027 10701 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 9943 10701 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7580 10701 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7492 10701 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7404 10701 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7316 10701 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7228 10701 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7140 10701 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 7052 10701 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10661 6964 10701 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 10111 10619 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 10027 10619 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 9943 10619 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 7580 10619 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10432 7357 10668 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10432 7357 10668 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10432 7357 10668 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 7316 10619 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10579 7228 10619 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10432 6991 10668 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10432 6991 10668 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10432 6991 10668 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10380 9929 10616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10380 9929 10616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10380 9929 10616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10497 7316 10537 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10497 7228 10537 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10415 7316 10455 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10415 7228 10455 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 10111 10373 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 10027 10373 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 9943 10373 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7580 10373 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7492 10373 7532 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7404 10373 7444 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7316 10373 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7228 10373 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7140 10373 7180 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 7052 10373 7092 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10333 6964 10373 7004 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 10111 10291 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 10027 10291 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 9943 10291 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 7580 10291 7620 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10111 7357 10347 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10111 7357 10347 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10111 7357 10347 7593 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 7316 10291 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10251 7228 10291 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10111 6991 10347 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10111 6991 10347 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10111 6991 10347 7227 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 10048 9929 10284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 10048 9929 10284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10048 9929 10284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10169 7316 10209 7356 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 10169 7228 10209 7268 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 4711 9929 4947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4711 9929 4947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4711 9929 4947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7568 4874 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7568 4874 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7480 4874 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7480 4874 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7392 4874 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7392 4874 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7304 4874 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7304 4874 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7216 4874 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7216 4874 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7128 4874 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7128 4874 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 7040 4874 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 7040 4874 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4810 6952 4874 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4810 6952 4874 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7568 4793 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7568 4793 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7480 4793 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7480 4793 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7392 4793 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7392 4793 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7304 4793 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7304 4793 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7216 4793 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7216 4793 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7128 4793 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7128 4793 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 7040 4793 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 7040 4793 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4729 6952 4793 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4729 6952 4793 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4660 10111 4700 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4660 10027 4700 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4660 9943 4700 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7568 4712 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7568 4712 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7480 4712 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7480 4712 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7392 4712 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7392 4712 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7304 4712 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7304 4712 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7216 4712 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7216 4712 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7128 4712 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7128 4712 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 7040 4712 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 7040 4712 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4648 6952 4712 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4648 6952 4712 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4579 10111 4619 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4579 10027 4619 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4579 9943 4619 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7568 4631 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7568 4631 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7480 4631 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7480 4631 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7392 4631 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7392 4631 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7304 4631 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7304 4631 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7216 4631 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7216 4631 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7128 4631 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7128 4631 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 7040 4631 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 7040 4631 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4567 6952 4631 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4567 6952 4631 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 4380 9929 4616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4380 9929 4616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4380 9929 4616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7568 4550 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7568 4550 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7480 4550 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7480 4550 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7392 4550 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7392 4550 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7304 4550 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7304 4550 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7216 4550 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7216 4550 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7128 4550 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7128 4550 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 7040 4550 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 7040 4550 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4486 6952 4550 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4486 6952 4550 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7568 4469 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7568 4469 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7480 4469 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7480 4469 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7392 4469 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7392 4469 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7304 4469 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7304 4469 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7216 4469 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7216 4469 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7128 4469 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7128 4469 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 7040 4469 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 7040 4469 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4405 6952 4469 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4405 6952 4469 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4336 10111 4376 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4336 10027 4376 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4336 9943 4376 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7568 4388 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7568 4388 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7480 4388 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7480 4388 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7392 4388 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7392 4388 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7304 4388 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7304 4388 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7216 4388 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7216 4388 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7128 4388 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7128 4388 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 7040 4388 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 7040 4388 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4324 6952 4388 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4324 6952 4388 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4255 10111 4295 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4255 10027 4295 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4255 9943 4295 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7568 4307 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7568 4307 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7480 4307 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7480 4307 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7392 4307 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7392 4307 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7304 4307 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7304 4307 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7216 4307 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7216 4307 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7128 4307 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7128 4307 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 7040 4307 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 7040 4307 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4243 6952 4307 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4243 6952 4307 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 4048 9929 4284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4048 9929 4284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4048 9929 4284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7568 4226 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7568 4226 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7480 4226 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7480 4226 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7392 4226 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7392 4226 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7304 4226 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7304 4226 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7216 4226 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7216 4226 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7128 4226 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7128 4226 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 7040 4226 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 7040 4226 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4162 6952 4226 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4162 6952 4226 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7568 4145 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7568 4145 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7480 4145 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7480 4145 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7392 4145 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7392 4145 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7304 4145 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7304 4145 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7216 4145 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7216 4145 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7128 4145 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7128 4145 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 7040 4145 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 7040 4145 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4081 6952 4145 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4081 6952 4145 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7568 4064 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7568 4064 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7480 4064 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7480 4064 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7392 4064 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7392 4064 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7304 4064 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7304 4064 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7216 4064 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7216 4064 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7128 4064 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7128 4064 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 7040 4064 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 7040 4064 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 4000 6952 4064 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 4000 6952 4064 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3931 10111 3971 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3931 10027 3971 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3931 9943 3971 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7568 3983 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7568 3983 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7480 3983 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7480 3983 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7392 3983 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7392 3983 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7304 3983 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7304 3983 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7216 3983 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7216 3983 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7128 3983 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7128 3983 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 7040 3983 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 7040 3983 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3919 6952 3983 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3919 6952 3983 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 3711 9929 3947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3711 9929 3947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3711 9929 3947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7568 3902 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7568 3902 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7480 3902 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7480 3902 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7392 3902 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7392 3902 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7304 3902 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7304 3902 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7216 3902 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7216 3902 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7128 3902 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7128 3902 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 7040 3902 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 7040 3902 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3838 6952 3902 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3838 6952 3902 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7568 3821 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7568 3821 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7480 3821 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7480 3821 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7392 3821 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7392 3821 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7304 3821 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7304 3821 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7216 3821 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7216 3821 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7128 3821 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7128 3821 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 7040 3821 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 7040 3821 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3757 6952 3821 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3757 6952 3821 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7568 3740 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7568 3740 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7480 3740 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7480 3740 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7392 3740 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7392 3740 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7304 3740 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7304 3740 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7216 3740 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7216 3740 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7128 3740 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7128 3740 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 7040 3740 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 7040 3740 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3676 6952 3740 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3676 6952 3740 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3607 10111 3647 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3607 10027 3647 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3607 9943 3647 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7568 3659 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7568 3659 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7480 3659 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7480 3659 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7392 3659 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7392 3659 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7304 3659 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7304 3659 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7216 3659 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7216 3659 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7128 3659 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7128 3659 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 7040 3659 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 7040 3659 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3595 6952 3659 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3595 6952 3659 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 3380 9929 3616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3380 9929 3616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3380 9929 3616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7568 3578 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7568 3578 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7480 3578 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7480 3578 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7392 3578 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7392 3578 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7304 3578 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7304 3578 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7216 3578 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7216 3578 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7128 3578 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7128 3578 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 7040 3578 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 7040 3578 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3514 6952 3578 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3514 6952 3578 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7568 3497 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7568 3497 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7480 3497 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7480 3497 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7392 3497 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7392 3497 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7304 3497 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7304 3497 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7216 3497 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7216 3497 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7128 3497 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7128 3497 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 7040 3497 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 7040 3497 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3433 6952 3497 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3433 6952 3497 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7568 3416 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7568 3416 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7480 3416 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7480 3416 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7392 3416 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7392 3416 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7304 3416 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7304 3416 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7216 3416 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7216 3416 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7128 3416 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7128 3416 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 7040 3416 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 7040 3416 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3352 6952 3416 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3352 6952 3416 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3283 10111 3323 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3283 10027 3323 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3283 9943 3323 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7568 3335 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7568 3335 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7480 3335 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7480 3335 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7392 3335 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7392 3335 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7304 3335 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7304 3335 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7216 3335 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7216 3335 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7128 3335 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7128 3335 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 7040 3335 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 7040 3335 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3271 6952 3335 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3271 6952 3335 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 3048 9929 3284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3048 9929 3284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3048 9929 3284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7568 3254 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7568 3254 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7480 3254 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7480 3254 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7392 3254 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7392 3254 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7304 3254 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7304 3254 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7216 3254 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7216 3254 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7128 3254 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7128 3254 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 7040 3254 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 7040 3254 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3190 6952 3254 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3190 6952 3254 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7568 3173 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7568 3173 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7480 3173 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7480 3173 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7392 3173 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7392 3173 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7304 3173 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7304 3173 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7216 3173 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7216 3173 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7128 3173 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7128 3173 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 7040 3173 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 7040 3173 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3109 6952 3173 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3109 6952 3173 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7568 3092 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7568 3092 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7480 3092 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7480 3092 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7392 3092 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7392 3092 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7304 3092 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7304 3092 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7216 3092 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7216 3092 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7128 3092 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7128 3092 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 7040 3092 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 7040 3092 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 3028 6952 3092 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 3028 6952 3092 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2959 10111 2999 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2959 10027 2999 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2959 9943 2999 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7568 3011 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7568 3011 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7480 3011 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7480 3011 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7392 3011 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7392 3011 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7304 3011 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7304 3011 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7216 3011 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7216 3011 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7128 3011 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7128 3011 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 7040 3011 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 7040 3011 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2947 6952 3011 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2947 6952 3011 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 2711 9929 2947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2711 9929 2947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2711 9929 2947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7568 2930 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7568 2930 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7480 2930 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7480 2930 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7392 2930 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7392 2930 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7304 2930 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7304 2930 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7216 2930 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7216 2930 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7128 2930 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7128 2930 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 7040 2930 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 7040 2930 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2866 6952 2930 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2866 6952 2930 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7568 2849 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7568 2849 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7480 2849 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7480 2849 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7392 2849 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7392 2849 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7304 2849 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7304 2849 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7216 2849 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7216 2849 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7128 2849 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7128 2849 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 7040 2849 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 7040 2849 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2785 6952 2849 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2785 6952 2849 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7568 2768 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7568 2768 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7480 2768 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7480 2768 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7392 2768 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7392 2768 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7304 2768 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7304 2768 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7216 2768 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7216 2768 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7128 2768 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7128 2768 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 7040 2768 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 7040 2768 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2704 6952 2768 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2704 6952 2768 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2635 10111 2675 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2635 10027 2675 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2635 9943 2675 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7568 2687 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7568 2687 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7480 2687 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7480 2687 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7392 2687 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7392 2687 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7304 2687 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7304 2687 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7216 2687 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7216 2687 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7128 2687 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7128 2687 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 7040 2687 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 7040 2687 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2623 6952 2687 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2623 6952 2687 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 2380 9929 2616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 9929 2616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 9929 2616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7568 2606 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7568 2606 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7480 2606 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7480 2606 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7392 2606 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7392 2606 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7304 2606 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7304 2606 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7216 2606 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7216 2606 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7128 2606 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7128 2606 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 7040 2606 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 7040 2606 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2542 6952 2606 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2542 6952 2606 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7568 2525 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7568 2525 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7480 2525 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7480 2525 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7392 2525 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7392 2525 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7304 2525 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7304 2525 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7216 2525 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7216 2525 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7128 2525 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7128 2525 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 7040 2525 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 7040 2525 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2461 6952 2525 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2461 6952 2525 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7568 2444 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7568 2444 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7480 2444 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7480 2444 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7392 2444 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7392 2444 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7304 2444 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7304 2444 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7216 2444 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7216 2444 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7128 2444 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7128 2444 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 7040 2444 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 7040 2444 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2380 6952 2444 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2380 6952 2444 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2311 10111 2351 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2311 10027 2351 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2311 9943 2351 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7568 2363 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7568 2363 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7480 2363 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7480 2363 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7392 2363 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7392 2363 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7304 2363 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7304 2363 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7216 2363 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7216 2363 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7128 2363 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7128 2363 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 7040 2363 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 7040 2363 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2299 6952 2363 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2299 6952 2363 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 2048 9929 2284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2048 9929 2284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2048 9929 2284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7568 2282 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7568 2282 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7480 2282 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7480 2282 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7392 2282 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7392 2282 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7304 2282 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7304 2282 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7216 2282 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7216 2282 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7128 2282 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7128 2282 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 7040 2282 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 7040 2282 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2218 6952 2282 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2218 6952 2282 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7568 2201 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7568 2201 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7480 2201 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7480 2201 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7392 2201 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7392 2201 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7304 2201 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7304 2201 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7216 2201 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7216 2201 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7128 2201 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7128 2201 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 7040 2201 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 7040 2201 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2137 6952 2201 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2137 6952 2201 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7568 2120 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7568 2120 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7480 2120 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7480 2120 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7392 2120 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7392 2120 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7304 2120 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7304 2120 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7216 2120 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7216 2120 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7128 2120 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7128 2120 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 7040 2120 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 7040 2120 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 2056 6952 2120 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 2056 6952 2120 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1987 10111 2027 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1987 10027 2027 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1987 9943 2027 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7568 2039 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7568 2039 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7480 2039 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7480 2039 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7392 2039 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7392 2039 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7304 2039 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7304 2039 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7216 2039 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7216 2039 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7128 2039 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7128 2039 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 7040 2039 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 7040 2039 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1975 6952 2039 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1975 6952 2039 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 1711 9929 1947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1711 9929 1947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1711 9929 1947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7568 1958 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7568 1958 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7480 1958 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7480 1958 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7392 1958 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7392 1958 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7304 1958 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7304 1958 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7216 1958 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7216 1958 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7128 1958 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7128 1958 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 7040 1958 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 7040 1958 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1894 6952 1958 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1894 6952 1958 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7568 1877 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7568 1877 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7480 1877 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7480 1877 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7392 1877 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7392 1877 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7304 1877 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7304 1877 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7216 1877 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7216 1877 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7128 1877 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7128 1877 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 7040 1877 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 7040 1877 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1813 6952 1877 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1813 6952 1877 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7568 1796 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7568 1796 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7480 1796 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7480 1796 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7392 1796 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7392 1796 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7304 1796 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7304 1796 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7216 1796 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7216 1796 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7128 1796 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7128 1796 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 7040 1796 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 7040 1796 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1732 6952 1796 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1732 6952 1796 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1663 10111 1703 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1663 10027 1703 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1663 9943 1703 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7568 1715 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7568 1715 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7480 1715 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7480 1715 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7392 1715 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7392 1715 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7304 1715 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7304 1715 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7216 1715 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7216 1715 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7128 1715 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7128 1715 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 7040 1715 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 7040 1715 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1651 6952 1715 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1651 6952 1715 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1582 10111 1622 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1582 10027 1622 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1582 9943 1622 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7568 1634 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7568 1634 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7480 1634 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7480 1634 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7392 1634 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7392 1634 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7304 1634 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7304 1634 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7216 1634 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7216 1634 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7128 1634 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7128 1634 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 7040 1634 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 7040 1634 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1570 6952 1634 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1570 6952 1634 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 1380 9929 1616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1380 9929 1616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1380 9929 1616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7568 1553 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7568 1553 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7480 1553 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7480 1553 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7392 1553 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7392 1553 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7304 1553 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7304 1553 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7216 1553 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7216 1553 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7128 1553 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7128 1553 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 7040 1553 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 7040 1553 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1489 6952 1553 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1489 6952 1553 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7568 1472 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7568 1472 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7480 1472 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7480 1472 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7392 1472 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7392 1472 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7304 1472 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7304 1472 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7216 1472 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7216 1472 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7128 1472 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7128 1472 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 7040 1472 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 7040 1472 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1408 6952 1472 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1408 6952 1472 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1339 10111 1379 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1339 10027 1379 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1339 9943 1379 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7568 1391 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7568 1391 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7480 1391 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7480 1391 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7392 1391 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7392 1391 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7304 1391 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7304 1391 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7216 1391 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7216 1391 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7128 1391 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7128 1391 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 7040 1391 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 7040 1391 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1327 6952 1391 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1327 6952 1391 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1258 10111 1298 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1258 10027 1298 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1258 9943 1298 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7568 1310 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7568 1310 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7480 1310 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7480 1310 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7392 1310 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7392 1310 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7304 1310 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7304 1310 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7216 1310 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7216 1310 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7128 1310 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7128 1310 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 7040 1310 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 7040 1310 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1246 6952 1310 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1246 6952 1310 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 1048 9929 1284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1048 9929 1284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1048 9929 1284 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7568 1229 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7568 1229 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7480 1229 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7480 1229 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7392 1229 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7392 1229 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7304 1229 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7304 1229 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7216 1229 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7216 1229 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7128 1229 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7128 1229 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 7040 1229 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 7040 1229 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1165 6952 1229 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1165 6952 1229 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7568 1148 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7568 1148 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7480 1148 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7480 1148 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7392 1148 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7392 1148 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7304 1148 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7304 1148 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7216 1148 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7216 1148 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7128 1148 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7128 1148 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 7040 1148 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 7040 1148 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1084 6952 1148 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1084 6952 1148 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7568 1067 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7568 1067 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7480 1067 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7480 1067 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7392 1067 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7392 1067 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7304 1067 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7304 1067 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7216 1067 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7216 1067 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7128 1067 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7128 1067 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 7040 1067 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 7040 1067 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 1003 6952 1067 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 1003 6952 1067 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 934 10111 974 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 934 10027 974 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 934 9943 974 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7568 986 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7568 986 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7480 986 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7480 986 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7392 986 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7392 986 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7304 986 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7304 986 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7216 986 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7216 986 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7128 986 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7128 986 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 7040 986 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 7040 986 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 922 6952 986 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 922 6952 986 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 711 9929 947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 711 9929 947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 711 9929 947 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7568 905 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7568 905 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7480 905 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7480 905 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7392 905 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7392 905 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7304 905 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7304 905 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7216 905 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7216 905 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7128 905 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7128 905 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 7040 905 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 7040 905 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 841 6952 905 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 841 6952 905 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7568 824 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7568 824 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7480 824 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7480 824 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7392 824 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7392 824 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7304 824 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7304 824 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7216 824 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7216 824 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7128 824 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7128 824 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 7040 824 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 7040 824 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 760 6952 824 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 760 6952 824 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7568 743 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7568 743 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7480 743 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7480 743 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7392 743 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7392 743 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7304 743 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7304 743 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7216 743 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7216 743 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7128 743 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7128 743 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 7040 743 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 7040 743 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 679 6952 743 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 679 6952 743 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 610 10111 650 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 610 10027 650 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 610 9943 650 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7568 662 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7568 662 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7480 662 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7480 662 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7392 662 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7392 662 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7304 662 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7304 662 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7216 662 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7216 662 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7128 662 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7128 662 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 7040 662 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 7040 662 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 598 6952 662 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 598 6952 662 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 380 9929 616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 380 9929 616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 380 9929 616 10165 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7568 580 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7568 580 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7480 580 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7480 580 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7392 580 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7392 580 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7304 580 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7304 580 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7216 580 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7216 580 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7128 580 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7128 580 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 7040 580 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 7040 580 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 516 6952 580 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 516 6952 580 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7568 498 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7568 498 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7480 498 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7480 498 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7392 498 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7392 498 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7304 498 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7304 498 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7216 498 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7216 498 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7128 498 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7128 498 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 7040 498 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 7040 498 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 434 6952 498 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 434 6952 498 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7568 416 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7568 416 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7480 416 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7480 416 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7392 416 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7392 416 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7304 416 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7304 416 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7216 416 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7216 416 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7128 416 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7128 416 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 7040 416 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 7040 416 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 352 6952 416 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 352 6952 416 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 282 10111 322 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 282 10027 322 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 282 9943 322 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7568 334 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7568 334 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7480 334 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7480 334 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7392 334 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7392 334 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7304 334 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7304 334 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7216 334 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7216 334 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7128 334 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7128 334 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 7040 334 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 7040 334 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal4 s 270 6952 334 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 270 6952 334 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 200 10111 240 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 200 10027 240 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 200 9943 240 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7568 252 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7480 252 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7392 252 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7304 252 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7216 252 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7128 252 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 7040 252 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 188 6952 252 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 118 10111 158 10151 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 118 10027 158 10067 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 118 9943 158 9983 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7568 170 7632 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7480 170 7544 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7392 170 7456 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7304 170 7368 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7216 170 7280 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7128 170 7192 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 7040 170 7104 6 VSSA
port 4 nsew ground bidirectional
rlabel metal3 s 106 6952 170 7016 6 VSSA
port 4 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 5 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 5 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 5 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 6 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 8 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 9 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 9 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 10 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 10 nsew power bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 12 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 11749940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11658148
<< end >>
