magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 2136 91 4159 2085
<< nwell >>
rect 2056 1805 4239 2165
rect 3879 371 4239 1805
rect 7827 433 8377 1383
rect 2056 11 4239 371
rect 7757 27 8377 433
<< pwell >>
rect 2243 1659 3819 1745
rect 3733 517 3819 1659
rect 2243 431 3819 517
<< nsubdiff >>
rect 7863 1313 7887 1347
rect 7921 1313 7967 1347
rect 8001 1313 8046 1347
rect 8080 1313 8125 1347
rect 8159 1313 8204 1347
rect 8238 1313 8283 1347
rect 8317 1313 8341 1347
rect 7863 1279 7897 1313
rect 8307 1279 8341 1313
rect 7863 1210 7897 1245
rect 8307 1210 8341 1245
rect 7863 1141 7897 1176
rect 7863 1073 7897 1107
rect 7863 1005 7897 1039
rect 7863 937 7897 971
rect 7863 869 7897 903
rect 7863 801 7897 835
rect 7863 733 7897 767
rect 7863 665 7897 699
rect 7863 597 7897 631
rect 7863 529 7897 563
rect 7863 461 7897 495
rect 7863 393 7897 427
rect 7863 325 7897 359
rect 7863 257 7897 291
rect 7863 189 7897 223
rect 7863 121 7897 155
rect 8307 1141 8341 1176
rect 8307 1073 8341 1107
rect 8307 1005 8341 1039
rect 8307 937 8341 971
rect 8307 869 8341 903
rect 8307 801 8341 835
rect 8307 733 8341 767
rect 8307 665 8341 699
rect 8307 597 8341 631
rect 8307 529 8341 563
rect 8307 461 8341 495
rect 8307 393 8341 427
rect 8307 325 8341 359
rect 8307 257 8341 291
rect 8307 189 8341 223
rect 8307 121 8341 155
rect 7897 87 7931 97
rect 7863 63 7931 87
rect 7965 63 8033 97
rect 8067 63 8146 97
rect 8180 63 8228 97
rect 8262 87 8307 97
rect 8262 63 8341 87
<< mvpsubdiff >>
rect 2269 1685 2303 1719
rect 2337 1685 2371 1719
rect 2405 1685 2439 1719
rect 2473 1685 2507 1719
rect 2541 1685 2575 1719
rect 2609 1685 2643 1719
rect 2677 1685 2711 1719
rect 2745 1685 2779 1719
rect 2813 1685 2847 1719
rect 2881 1685 3000 1719
rect 3034 1685 3068 1719
rect 3102 1685 3136 1719
rect 3170 1685 3204 1719
rect 3238 1685 3272 1719
rect 3306 1685 3340 1719
rect 3374 1685 3408 1719
rect 3442 1685 3476 1719
rect 3510 1685 3544 1719
rect 3578 1685 3612 1719
rect 3646 1685 3680 1719
rect 3714 1685 3793 1719
rect 3759 1617 3793 1651
rect 3759 1549 3793 1583
rect 3759 1481 3793 1515
rect 3759 1413 3793 1447
rect 3759 1345 3793 1379
rect 3759 1277 3793 1311
rect 3759 1209 3793 1243
rect 3759 1141 3793 1175
rect 3759 1073 3793 1107
rect 3759 1005 3793 1039
rect 3759 937 3793 971
rect 3759 869 3793 903
rect 3759 801 3793 835
rect 3759 733 3793 767
rect 3759 665 3793 699
rect 3759 597 3793 631
rect 2269 457 2365 491
rect 2399 457 2433 491
rect 2467 457 2501 491
rect 2535 457 2569 491
rect 2603 457 2637 491
rect 2671 457 2705 491
rect 2739 457 2773 491
rect 2807 457 2841 491
rect 2875 457 2909 491
rect 2943 457 2977 491
rect 3011 457 3045 491
rect 3079 457 3113 491
rect 3147 457 3181 491
rect 3215 457 3249 491
rect 3283 457 3317 491
rect 3351 457 3385 491
rect 3419 457 3453 491
rect 3487 457 3521 491
rect 3555 457 3589 491
rect 3623 457 3657 491
rect 3691 457 3725 491
rect 3759 457 3793 563
<< mvnsubdiff >>
rect 2196 2042 4116 2076
rect 2196 1872 2230 2042
rect 3964 2008 3998 2042
rect 4032 2008 4116 2042
rect 3964 1974 4082 2008
rect 3964 1940 4014 1974
rect 4048 1940 4116 1974
rect 3896 1906 4082 1940
rect 3896 1872 4116 1906
rect 3945 1848 4116 1872
rect 3979 1814 4116 1848
rect 3945 1806 4116 1814
rect 3945 1780 4042 1806
rect 3979 1772 4042 1780
rect 4076 1772 4116 1806
rect 3979 1746 4116 1772
rect 3945 1738 4116 1746
rect 3945 1712 4042 1738
rect 3979 1704 4042 1712
rect 4076 1704 4116 1738
rect 3979 1678 4116 1704
rect 3945 1670 4116 1678
rect 3945 1644 4042 1670
rect 3979 1636 4042 1644
rect 4076 1636 4116 1670
rect 3979 1610 4116 1636
rect 3945 1602 4116 1610
rect 3945 1576 4042 1602
rect 3979 1568 4042 1576
rect 4076 1568 4116 1602
rect 3979 1542 4116 1568
rect 3945 1534 4116 1542
rect 3945 1508 4042 1534
rect 3979 1500 4042 1508
rect 4076 1500 4116 1534
rect 3979 1474 4116 1500
rect 3945 1466 4116 1474
rect 3945 1440 4042 1466
rect 3979 1432 4042 1440
rect 4076 1432 4116 1466
rect 3979 1406 4116 1432
rect 3945 1398 4116 1406
rect 3945 1372 4042 1398
rect 3979 1364 4042 1372
rect 4076 1364 4116 1398
rect 3979 1338 4116 1364
rect 3945 1330 4116 1338
rect 3945 1304 4042 1330
rect 3979 1296 4042 1304
rect 4076 1296 4116 1330
rect 3979 1270 4116 1296
rect 3945 1262 4116 1270
rect 3945 1236 4042 1262
rect 3979 1228 4042 1236
rect 4076 1228 4116 1262
rect 3979 1202 4116 1228
rect 3945 1194 4116 1202
rect 3945 1167 4042 1194
rect 3979 1160 4042 1167
rect 4076 1160 4116 1194
rect 3979 1133 4116 1160
rect 3945 1126 4116 1133
rect 3945 1098 4042 1126
rect 3979 1092 4042 1098
rect 4076 1092 4116 1126
rect 3979 1064 4116 1092
rect 3945 1058 4116 1064
rect 3945 1029 4042 1058
rect 3979 1024 4042 1029
rect 4076 1024 4116 1058
rect 3979 995 4116 1024
rect 3945 990 4116 995
rect 3945 960 4042 990
rect 3979 956 4042 960
rect 4076 956 4116 990
rect 3979 926 4116 956
rect 3945 922 4116 926
rect 3945 891 4042 922
rect 3979 888 4042 891
rect 4076 888 4116 922
rect 3979 857 4116 888
rect 3945 854 4116 857
rect 3945 822 4042 854
rect 3979 820 4042 822
rect 4076 820 4116 854
rect 3979 788 4116 820
rect 3945 786 4116 788
rect 3945 753 4042 786
rect 3979 752 4042 753
rect 4076 752 4116 786
rect 3979 719 4116 752
rect 3945 718 4116 719
rect 3945 684 4042 718
rect 4076 684 4116 718
rect 3979 650 4116 684
rect 3945 616 4042 650
rect 4076 616 4116 650
rect 3945 615 4116 616
rect 3979 582 4116 615
rect 3979 581 4042 582
rect 3945 548 4042 581
rect 4076 548 4116 582
rect 3945 546 4116 548
rect 3979 514 4116 546
rect 3979 512 4042 514
rect 3945 480 4042 512
rect 4076 480 4116 514
rect 3945 477 4116 480
rect 3979 446 4116 477
rect 3979 443 4042 446
rect 3945 412 4042 443
rect 4076 412 4116 446
rect 3945 408 4116 412
rect 3979 378 4116 408
rect 3979 374 4042 378
rect 3945 344 4042 374
rect 4076 344 4116 378
rect 3945 339 4116 344
rect 3979 310 4116 339
rect 3979 305 4042 310
rect 2214 271 2238 305
rect 2272 271 2308 305
rect 2342 271 2378 305
rect 2412 271 2448 305
rect 2482 271 2518 305
rect 2552 271 2588 305
rect 2622 271 2658 305
rect 2692 271 2728 305
rect 2762 271 2798 305
rect 2832 271 2868 305
rect 2902 271 2938 305
rect 2972 271 3008 305
rect 3042 271 3078 305
rect 3112 271 3148 305
rect 3182 271 3218 305
rect 3252 271 3288 305
rect 3322 271 3358 305
rect 3392 271 3427 305
rect 3461 271 3496 305
rect 3530 271 3565 305
rect 3599 271 3634 305
rect 3668 271 3703 305
rect 3737 271 3772 305
rect 3806 271 3841 305
rect 3875 276 4042 305
rect 4076 276 4116 310
rect 3875 271 4116 276
rect 2214 242 4116 271
rect 2214 208 4042 242
rect 4076 208 4116 242
rect 2214 174 2248 208
rect 2282 174 2316 208
rect 2350 174 2384 208
rect 2418 174 2452 208
rect 2486 174 2520 208
rect 2554 174 2588 208
rect 2622 174 2656 208
rect 2690 174 2724 208
rect 2758 174 2792 208
rect 2826 174 2860 208
rect 2894 174 2928 208
rect 2962 174 2996 208
rect 3030 174 3064 208
rect 3098 174 3132 208
rect 3166 174 3200 208
rect 3234 174 3268 208
rect 3302 174 3336 208
rect 3370 174 3404 208
rect 3438 174 3472 208
rect 3506 174 3540 208
rect 3574 174 3608 208
rect 3642 174 3676 208
rect 3710 174 3744 208
rect 3778 174 3812 208
rect 3846 174 3880 208
rect 3914 174 3948 208
rect 3982 174 4116 208
<< nsubdiffcont >>
rect 7887 1313 7921 1347
rect 7967 1313 8001 1347
rect 8046 1313 8080 1347
rect 8125 1313 8159 1347
rect 8204 1313 8238 1347
rect 8283 1313 8317 1347
rect 7863 1245 7897 1279
rect 7863 1176 7897 1210
rect 8307 1245 8341 1279
rect 7863 1107 7897 1141
rect 7863 1039 7897 1073
rect 7863 971 7897 1005
rect 7863 903 7897 937
rect 7863 835 7897 869
rect 7863 767 7897 801
rect 7863 699 7897 733
rect 7863 631 7897 665
rect 7863 563 7897 597
rect 7863 495 7897 529
rect 7863 427 7897 461
rect 7863 359 7897 393
rect 7863 291 7897 325
rect 7863 223 7897 257
rect 7863 155 7897 189
rect 7863 87 7897 121
rect 8307 1176 8341 1210
rect 8307 1107 8341 1141
rect 8307 1039 8341 1073
rect 8307 971 8341 1005
rect 8307 903 8341 937
rect 8307 835 8341 869
rect 8307 767 8341 801
rect 8307 699 8341 733
rect 8307 631 8341 665
rect 8307 563 8341 597
rect 8307 495 8341 529
rect 8307 427 8341 461
rect 8307 359 8341 393
rect 8307 291 8341 325
rect 8307 223 8341 257
rect 8307 155 8341 189
rect 7931 63 7965 97
rect 8033 63 8067 97
rect 8146 63 8180 97
rect 8228 63 8262 97
rect 8307 87 8341 121
<< mvpsubdiffcont >>
rect 2303 1685 2337 1719
rect 2371 1685 2405 1719
rect 2439 1685 2473 1719
rect 2507 1685 2541 1719
rect 2575 1685 2609 1719
rect 2643 1685 2677 1719
rect 2711 1685 2745 1719
rect 2779 1685 2813 1719
rect 2847 1685 2881 1719
rect 3000 1685 3034 1719
rect 3068 1685 3102 1719
rect 3136 1685 3170 1719
rect 3204 1685 3238 1719
rect 3272 1685 3306 1719
rect 3340 1685 3374 1719
rect 3408 1685 3442 1719
rect 3476 1685 3510 1719
rect 3544 1685 3578 1719
rect 3612 1685 3646 1719
rect 3680 1685 3714 1719
rect 3759 1651 3793 1685
rect 3759 1583 3793 1617
rect 3759 1515 3793 1549
rect 3759 1447 3793 1481
rect 3759 1379 3793 1413
rect 3759 1311 3793 1345
rect 3759 1243 3793 1277
rect 3759 1175 3793 1209
rect 3759 1107 3793 1141
rect 3759 1039 3793 1073
rect 3759 971 3793 1005
rect 3759 903 3793 937
rect 3759 835 3793 869
rect 3759 767 3793 801
rect 3759 699 3793 733
rect 3759 631 3793 665
rect 3759 563 3793 597
rect 2365 457 2399 491
rect 2433 457 2467 491
rect 2501 457 2535 491
rect 2569 457 2603 491
rect 2637 457 2671 491
rect 2705 457 2739 491
rect 2773 457 2807 491
rect 2841 457 2875 491
rect 2909 457 2943 491
rect 2977 457 3011 491
rect 3045 457 3079 491
rect 3113 457 3147 491
rect 3181 457 3215 491
rect 3249 457 3283 491
rect 3317 457 3351 491
rect 3385 457 3419 491
rect 3453 457 3487 491
rect 3521 457 3555 491
rect 3589 457 3623 491
rect 3657 457 3691 491
rect 3725 457 3759 491
<< mvnsubdiffcont >>
rect 2230 1940 3964 2042
rect 3998 2008 4032 2042
rect 4082 1974 4116 2008
rect 4014 1940 4048 1974
rect 2230 1872 3896 1940
rect 4082 1906 4116 1940
rect 3945 1814 3979 1848
rect 3945 1746 3979 1780
rect 4042 1772 4076 1806
rect 3945 1678 3979 1712
rect 4042 1704 4076 1738
rect 3945 1610 3979 1644
rect 4042 1636 4076 1670
rect 3945 1542 3979 1576
rect 4042 1568 4076 1602
rect 3945 1474 3979 1508
rect 4042 1500 4076 1534
rect 3945 1406 3979 1440
rect 4042 1432 4076 1466
rect 3945 1338 3979 1372
rect 4042 1364 4076 1398
rect 3945 1270 3979 1304
rect 4042 1296 4076 1330
rect 3945 1202 3979 1236
rect 4042 1228 4076 1262
rect 3945 1133 3979 1167
rect 4042 1160 4076 1194
rect 3945 1064 3979 1098
rect 4042 1092 4076 1126
rect 3945 995 3979 1029
rect 4042 1024 4076 1058
rect 3945 926 3979 960
rect 4042 956 4076 990
rect 3945 857 3979 891
rect 4042 888 4076 922
rect 3945 788 3979 822
rect 4042 820 4076 854
rect 3945 719 3979 753
rect 4042 752 4076 786
rect 4042 684 4076 718
rect 3945 650 3979 684
rect 4042 616 4076 650
rect 3945 581 3979 615
rect 4042 548 4076 582
rect 3945 512 3979 546
rect 4042 480 4076 514
rect 3945 443 3979 477
rect 4042 412 4076 446
rect 3945 374 3979 408
rect 4042 344 4076 378
rect 3945 305 3979 339
rect 2238 271 2272 305
rect 2308 271 2342 305
rect 2378 271 2412 305
rect 2448 271 2482 305
rect 2518 271 2552 305
rect 2588 271 2622 305
rect 2658 271 2692 305
rect 2728 271 2762 305
rect 2798 271 2832 305
rect 2868 271 2902 305
rect 2938 271 2972 305
rect 3008 271 3042 305
rect 3078 271 3112 305
rect 3148 271 3182 305
rect 3218 271 3252 305
rect 3288 271 3322 305
rect 3358 271 3392 305
rect 3427 271 3461 305
rect 3496 271 3530 305
rect 3565 271 3599 305
rect 3634 271 3668 305
rect 3703 271 3737 305
rect 3772 271 3806 305
rect 3841 271 3875 305
rect 4042 276 4076 310
rect 4042 208 4076 242
rect 2248 174 2282 208
rect 2316 174 2350 208
rect 2384 174 2418 208
rect 2452 174 2486 208
rect 2520 174 2554 208
rect 2588 174 2622 208
rect 2656 174 2690 208
rect 2724 174 2758 208
rect 2792 174 2826 208
rect 2860 174 2894 208
rect 2928 174 2962 208
rect 2996 174 3030 208
rect 3064 174 3098 208
rect 3132 174 3166 208
rect 3200 174 3234 208
rect 3268 174 3302 208
rect 3336 174 3370 208
rect 3404 174 3438 208
rect 3472 174 3506 208
rect 3540 174 3574 208
rect 3608 174 3642 208
rect 3676 174 3710 208
rect 3744 174 3778 208
rect 3812 174 3846 208
rect 3880 174 3914 208
rect 3948 174 3982 208
<< poly >>
rect 8909 22229 10821 22245
rect 8909 22213 9005 22229
rect 8909 22179 8925 22213
rect 8959 22195 9005 22213
rect 9039 22195 9075 22229
rect 9109 22195 9145 22229
rect 9179 22195 9215 22229
rect 9249 22195 9285 22229
rect 9319 22195 9355 22229
rect 9389 22195 9425 22229
rect 9459 22195 9495 22229
rect 9529 22195 9565 22229
rect 9599 22195 9635 22229
rect 9669 22195 9705 22229
rect 9739 22195 9775 22229
rect 9809 22195 9845 22229
rect 9879 22195 9915 22229
rect 9949 22195 9985 22229
rect 10019 22195 10056 22229
rect 10090 22195 10127 22229
rect 10161 22195 10198 22229
rect 10232 22195 10269 22229
rect 10303 22195 10340 22229
rect 10374 22195 10411 22229
rect 10445 22195 10482 22229
rect 10516 22195 10553 22229
rect 10587 22195 10624 22229
rect 10658 22195 10695 22229
rect 10729 22213 10821 22229
rect 10729 22195 10771 22213
rect 8959 22179 10771 22195
rect 10805 22179 10821 22213
rect 8909 22145 8975 22179
rect 8909 22111 8925 22145
rect 8959 22111 8975 22145
rect 8909 22077 8975 22111
rect 8909 22043 8925 22077
rect 8959 22043 8975 22077
rect 8909 22009 8975 22043
rect 8909 21975 8925 22009
rect 8959 21975 8975 22009
rect 8909 21941 8975 21975
rect 8909 21907 8925 21941
rect 8959 21907 8975 21941
rect 8909 21873 8975 21907
rect 8909 21839 8925 21873
rect 8959 21839 8975 21873
rect 8909 21805 8975 21839
rect 8909 21771 8925 21805
rect 8959 21771 8975 21805
rect 8909 21737 8975 21771
rect 8909 21703 8925 21737
rect 8959 21703 8975 21737
rect 8909 21669 8975 21703
rect 8909 21635 8925 21669
rect 8959 21635 8975 21669
rect 8909 21601 8975 21635
rect 8909 21567 8925 21601
rect 8959 21567 8975 21601
rect 8909 21533 8975 21567
rect 8909 21499 8925 21533
rect 8959 21499 8975 21533
rect 8909 21465 8975 21499
rect 8909 21431 8925 21465
rect 8959 21431 8975 21465
rect 8909 21397 8975 21431
rect 8909 21363 8925 21397
rect 8959 21363 8975 21397
rect 8909 21329 8975 21363
rect 8909 21295 8925 21329
rect 8959 21295 8975 21329
rect 8909 21261 8975 21295
rect 8909 21227 8925 21261
rect 8959 21227 8975 21261
rect 8909 21193 8975 21227
rect 8909 21159 8925 21193
rect 8959 21159 8975 21193
rect 8909 21125 8975 21159
rect 8909 21091 8925 21125
rect 8959 21091 8975 21125
rect 8909 21057 8975 21091
rect 8909 21023 8925 21057
rect 8959 21023 8975 21057
rect 8909 20989 8975 21023
rect 8909 20955 8925 20989
rect 8959 20955 8975 20989
rect 8909 20921 8975 20955
rect 8909 20887 8925 20921
rect 8959 20887 8975 20921
rect 8909 20853 8975 20887
rect 8909 20819 8925 20853
rect 8959 20819 8975 20853
rect 8909 20785 8975 20819
rect 8909 20751 8925 20785
rect 8959 20751 8975 20785
rect 8909 20717 8975 20751
rect 8909 20683 8925 20717
rect 8959 20683 8975 20717
rect 8909 20649 8975 20683
rect 8909 20615 8925 20649
rect 8959 20615 8975 20649
rect 8909 20581 8975 20615
rect 8909 20547 8925 20581
rect 8959 20547 8975 20581
rect 8909 20513 8975 20547
rect 8909 20479 8925 20513
rect 8959 20479 8975 20513
rect 8909 20445 8975 20479
rect 8909 20411 8925 20445
rect 8959 20411 8975 20445
rect 8909 20377 8975 20411
rect 8909 20343 8925 20377
rect 8959 20343 8975 20377
rect 8909 20309 8975 20343
rect 8909 20275 8925 20309
rect 8959 20275 8975 20309
rect 8909 20241 8975 20275
rect 8909 20207 8925 20241
rect 8959 20207 8975 20241
rect 8909 20173 8975 20207
rect 8909 20139 8925 20173
rect 8959 20139 8975 20173
rect 8909 20105 8975 20139
rect 8909 20071 8925 20105
rect 8959 20071 8975 20105
rect 8909 20037 8975 20071
rect 8909 20003 8925 20037
rect 8959 20003 8975 20037
rect 8909 19969 8975 20003
rect 8909 19935 8925 19969
rect 8959 19935 8975 19969
rect 8909 19901 8975 19935
rect 8909 19867 8925 19901
rect 8959 19867 8975 19901
rect 8909 19833 8975 19867
rect 8909 19799 8925 19833
rect 8959 19799 8975 19833
rect 8909 19765 8975 19799
rect 8909 19731 8925 19765
rect 8959 19731 8975 19765
rect 8909 19697 8975 19731
rect 8909 19663 8925 19697
rect 8959 19663 8975 19697
rect 8909 19629 8975 19663
rect 8909 19595 8925 19629
rect 8959 19595 8975 19629
rect 8909 19561 8975 19595
rect 8909 19527 8925 19561
rect 8959 19527 8975 19561
rect 8909 19493 8975 19527
rect 8909 19459 8925 19493
rect 8959 19459 8975 19493
rect 8909 19425 8975 19459
rect 8909 19391 8925 19425
rect 8959 19391 8975 19425
rect 8909 19357 8975 19391
rect 8909 19323 8925 19357
rect 8959 19323 8975 19357
rect 8909 19289 8975 19323
rect 8909 19255 8925 19289
rect 8959 19255 8975 19289
rect 8909 19221 8975 19255
rect 8909 19187 8925 19221
rect 8959 19187 8975 19221
rect 8909 19153 8975 19187
rect 8909 19119 8925 19153
rect 8959 19119 8975 19153
rect 8909 19085 8975 19119
rect 8909 19051 8925 19085
rect 8959 19051 8975 19085
rect 8909 19017 8975 19051
rect 8909 18983 8925 19017
rect 8959 18983 8975 19017
rect 8909 18949 8975 18983
rect 8909 18915 8925 18949
rect 8959 18915 8975 18949
rect 8909 18881 8975 18915
rect 8909 18847 8925 18881
rect 8959 18847 8975 18881
rect 8909 18813 8975 18847
rect 8909 18779 8925 18813
rect 8959 18779 8975 18813
rect 8909 18745 8975 18779
rect 8909 18711 8925 18745
rect 8959 18711 8975 18745
rect 8909 18677 8975 18711
rect 8909 18643 8925 18677
rect 8959 18643 8975 18677
rect 8909 18609 8975 18643
rect 8909 18575 8925 18609
rect 8959 18575 8975 18609
rect 8909 18541 8975 18575
rect 8909 18507 8925 18541
rect 8959 18507 8975 18541
rect 8909 18473 8975 18507
rect 8909 18439 8925 18473
rect 8959 18439 8975 18473
rect 8909 18405 8975 18439
rect 8909 18371 8925 18405
rect 8959 18371 8975 18405
rect 8909 18337 8975 18371
rect 8909 18303 8925 18337
rect 8959 18303 8975 18337
rect 8909 18269 8975 18303
rect 8909 18235 8925 18269
rect 8959 18235 8975 18269
rect 8909 18201 8975 18235
rect 8909 18167 8925 18201
rect 8959 18167 8975 18201
rect 8909 18133 8975 18167
rect 8909 18099 8925 18133
rect 8959 18099 8975 18133
rect 8909 18065 8975 18099
rect 8909 18031 8925 18065
rect 8959 18031 8975 18065
rect 8909 17997 8975 18031
rect 8909 17963 8925 17997
rect 8959 17963 8975 17997
rect 8909 17929 8975 17963
rect 8909 17895 8925 17929
rect 8959 17895 8975 17929
rect 8909 17861 8975 17895
rect 8909 17827 8925 17861
rect 8959 17827 8975 17861
rect 8909 17793 8975 17827
rect 8909 17759 8925 17793
rect 8959 17759 8975 17793
rect 8909 17725 8975 17759
rect 8909 17691 8925 17725
rect 8959 17691 8975 17725
rect 8909 17657 8975 17691
rect 8909 17623 8925 17657
rect 8959 17623 8975 17657
rect 8909 17589 8975 17623
rect 8909 17555 8925 17589
rect 8959 17555 8975 17589
rect 8909 17521 8975 17555
rect 8909 17487 8925 17521
rect 8959 17487 8975 17521
rect 8909 17453 8975 17487
rect 8909 17419 8925 17453
rect 8959 17419 8975 17453
rect 8909 17385 8975 17419
rect 8909 17351 8925 17385
rect 8959 17351 8975 17385
rect 8909 17317 8975 17351
rect 8909 17283 8925 17317
rect 8959 17283 8975 17317
rect 8909 17249 8975 17283
rect 8909 17215 8925 17249
rect 8959 17215 8975 17249
rect 8909 17181 8975 17215
rect 8909 17147 8925 17181
rect 8959 17147 8975 17181
rect 8909 17113 8975 17147
rect 8909 17079 8925 17113
rect 8959 17079 8975 17113
rect 8909 17045 8975 17079
rect 8909 17011 8925 17045
rect 8959 17011 8975 17045
rect 8909 16977 8975 17011
rect 8909 16943 8925 16977
rect 8959 16943 8975 16977
rect 8909 16909 8975 16943
rect 8909 16875 8925 16909
rect 8959 16875 8975 16909
rect 8909 16841 8975 16875
rect 8909 16807 8925 16841
rect 8959 16807 8975 16841
rect 8909 16773 8975 16807
rect 8909 16739 8925 16773
rect 8959 16739 8975 16773
rect 8909 16705 8975 16739
rect 8909 16671 8925 16705
rect 8959 16671 8975 16705
rect 8909 16637 8975 16671
rect 8909 16603 8925 16637
rect 8959 16603 8975 16637
rect 8909 16569 8975 16603
rect 8909 16535 8925 16569
rect 8959 16535 8975 16569
rect 8909 16501 8975 16535
rect 8909 16467 8925 16501
rect 8959 16467 8975 16501
rect 8909 16433 8975 16467
rect 8909 16399 8925 16433
rect 8959 16399 8975 16433
rect 8909 16365 8975 16399
rect 8909 16331 8925 16365
rect 8959 16331 8975 16365
rect 8909 16297 8975 16331
rect 8909 16263 8925 16297
rect 8959 16263 8975 16297
rect 8909 16229 8975 16263
rect 8909 16195 8925 16229
rect 8959 16195 8975 16229
rect 8909 16161 8975 16195
rect 8909 16127 8925 16161
rect 8959 16127 8975 16161
rect 8909 16093 8975 16127
rect 8909 16059 8925 16093
rect 8959 16059 8975 16093
rect 8909 16025 8975 16059
rect 8909 15991 8925 16025
rect 8959 15991 8975 16025
rect 8909 15957 8975 15991
rect 8909 15923 8925 15957
rect 8959 15923 8975 15957
rect 8909 15889 8975 15923
rect 8909 15855 8925 15889
rect 8959 15855 8975 15889
rect 8909 15821 8975 15855
rect 8909 15787 8925 15821
rect 8959 15787 8975 15821
rect 8909 15753 8975 15787
rect 8909 15719 8925 15753
rect 8959 15719 8975 15753
rect 8909 15685 8975 15719
rect 8909 15651 8925 15685
rect 8959 15651 8975 15685
rect 8909 15617 8975 15651
rect 8909 15583 8925 15617
rect 8959 15583 8975 15617
rect 8909 15549 8975 15583
rect 8909 15515 8925 15549
rect 8959 15515 8975 15549
rect 8909 15481 8975 15515
rect 8909 15447 8925 15481
rect 8959 15447 8975 15481
rect 8909 15413 8975 15447
rect 8909 15379 8925 15413
rect 8959 15379 8975 15413
rect 8909 15345 8975 15379
rect 8909 15311 8925 15345
rect 8959 15311 8975 15345
rect 8909 15277 8975 15311
rect 8909 15243 8925 15277
rect 8959 15243 8975 15277
rect 8909 15209 8975 15243
rect 8909 15175 8925 15209
rect 8959 15175 8975 15209
rect 8909 15141 8975 15175
rect 8909 15107 8925 15141
rect 8959 15107 8975 15141
rect 8909 15073 8975 15107
rect 8909 15039 8925 15073
rect 8959 15039 8975 15073
rect 8909 15005 8975 15039
rect 8909 14971 8925 15005
rect 8959 14971 8975 15005
rect 8909 14937 8975 14971
rect 8909 14903 8925 14937
rect 8959 14903 8975 14937
rect 8909 14869 8975 14903
rect 8909 14835 8925 14869
rect 8959 14835 8975 14869
rect 8909 14801 8975 14835
rect 8909 14767 8925 14801
rect 8959 14767 8975 14801
rect 8909 14733 8975 14767
rect 8909 14699 8925 14733
rect 8959 14699 8975 14733
rect 8909 14665 8975 14699
rect 8909 14631 8925 14665
rect 8959 14631 8975 14665
rect 8909 14597 8975 14631
rect 8909 14563 8925 14597
rect 8959 14563 8975 14597
rect 8909 14529 8975 14563
rect 8909 14495 8925 14529
rect 8959 14495 8975 14529
rect 8909 14461 8975 14495
rect 8909 14427 8925 14461
rect 8959 14427 8975 14461
rect 8909 14393 8975 14427
rect 8909 14359 8925 14393
rect 8959 14359 8975 14393
rect 8909 14325 8975 14359
rect 8909 14291 8925 14325
rect 8959 14291 8975 14325
rect 8909 14257 8975 14291
rect 8909 14223 8925 14257
rect 8959 14223 8975 14257
rect 8909 14189 8975 14223
rect 8909 14155 8925 14189
rect 8959 14155 8975 14189
rect 8909 14121 8975 14155
rect 8909 14087 8925 14121
rect 8959 14087 8975 14121
rect 8909 14053 8975 14087
rect 8909 14019 8925 14053
rect 8959 14019 8975 14053
rect 8909 13985 8975 14019
rect 8909 13951 8925 13985
rect 8959 13951 8975 13985
rect 8909 13917 8975 13951
rect 8909 13883 8925 13917
rect 8959 13883 8975 13917
rect 8909 13849 8975 13883
rect 8909 13815 8925 13849
rect 8959 13815 8975 13849
rect 8909 13781 8975 13815
rect 8909 13747 8925 13781
rect 8959 13747 8975 13781
rect 8909 13713 8975 13747
rect 8909 13679 8925 13713
rect 8959 13679 8975 13713
rect 8909 13645 8975 13679
rect 8909 13611 8925 13645
rect 8959 13611 8975 13645
rect 8909 13577 8975 13611
rect 8909 13543 8925 13577
rect 8959 13543 8975 13577
rect 8909 13509 8975 13543
rect 8909 13475 8925 13509
rect 8959 13475 8975 13509
rect 8909 13441 8975 13475
rect 8909 13407 8925 13441
rect 8959 13407 8975 13441
rect 8909 13373 8975 13407
rect 8909 13339 8925 13373
rect 8959 13339 8975 13373
rect 8909 13305 8975 13339
rect 8909 13271 8925 13305
rect 8959 13271 8975 13305
rect 8909 13237 8975 13271
rect 8909 13203 8925 13237
rect 8959 13203 8975 13237
rect 8909 13169 8975 13203
rect 8909 13135 8925 13169
rect 8959 13135 8975 13169
rect 8909 13101 8975 13135
rect 8909 13067 8925 13101
rect 8959 13067 8975 13101
rect 8909 13033 8975 13067
rect 8909 12999 8925 13033
rect 8959 12999 8975 13033
rect 8909 12965 8975 12999
rect 8909 12931 8925 12965
rect 8959 12931 8975 12965
rect 8909 12897 8975 12931
rect 8909 12863 8925 12897
rect 8959 12863 8975 12897
rect 8909 12829 8975 12863
rect 8909 12795 8925 12829
rect 8959 12795 8975 12829
rect 8909 12761 8975 12795
rect 8909 12727 8925 12761
rect 8959 12727 8975 12761
rect 8909 12693 8975 12727
rect 8909 12659 8925 12693
rect 8959 12659 8975 12693
rect 8909 12625 8975 12659
rect 8909 12591 8925 12625
rect 8959 12591 8975 12625
rect 8909 12557 8975 12591
rect 8909 12523 8925 12557
rect 8959 12523 8975 12557
rect 8909 12489 8975 12523
rect 8909 12455 8925 12489
rect 8959 12455 8975 12489
rect 8909 12421 8975 12455
rect 8909 12387 8925 12421
rect 8959 12387 8975 12421
rect 8909 12353 8975 12387
rect 8909 12319 8925 12353
rect 8959 12319 8975 12353
rect 8909 12285 8975 12319
rect 8909 12251 8925 12285
rect 8959 12251 8975 12285
rect 8909 12217 8975 12251
rect 8909 12183 8925 12217
rect 8959 12183 8975 12217
rect 8909 12149 8975 12183
rect 8909 12115 8925 12149
rect 8959 12115 8975 12149
rect 8909 12081 8975 12115
rect 8909 12047 8925 12081
rect 8959 12047 8975 12081
rect 8909 12013 8975 12047
rect 8909 11979 8925 12013
rect 8959 11979 8975 12013
rect 8909 11945 8975 11979
rect 8909 11911 8925 11945
rect 8959 11911 8975 11945
rect 8909 11877 8975 11911
rect 8909 11843 8925 11877
rect 8959 11843 8975 11877
rect 8909 11809 8975 11843
rect 8909 11775 8925 11809
rect 8959 11775 8975 11809
rect 8909 11741 8975 11775
rect 8909 11707 8925 11741
rect 8959 11707 8975 11741
rect 8909 11673 8975 11707
rect 8909 11639 8925 11673
rect 8959 11639 8975 11673
rect 8909 11605 8975 11639
rect 8909 11571 8925 11605
rect 8959 11571 8975 11605
rect 8909 11537 8975 11571
rect 8909 11503 8925 11537
rect 8959 11503 8975 11537
rect 8909 11469 8975 11503
rect 8909 11435 8925 11469
rect 8959 11435 8975 11469
rect 8909 11401 8975 11435
rect 8909 11367 8925 11401
rect 8959 11367 8975 11401
rect 8909 11333 8975 11367
rect 8909 11299 8925 11333
rect 8959 11299 8975 11333
rect 8909 11265 8975 11299
rect 8909 11231 8925 11265
rect 8959 11231 8975 11265
rect 8909 11197 8975 11231
rect 8909 11163 8925 11197
rect 8959 11163 8975 11197
rect 8909 11129 8975 11163
rect 8909 11095 8925 11129
rect 8959 11095 8975 11129
rect 8909 11061 8975 11095
rect 8909 11027 8925 11061
rect 8959 11027 8975 11061
rect 8909 10993 8975 11027
rect 8909 10959 8925 10993
rect 8959 10959 8975 10993
rect 8909 10925 8975 10959
rect 8909 10891 8925 10925
rect 8959 10891 8975 10925
rect 8909 10857 8975 10891
rect 8909 10823 8925 10857
rect 8959 10823 8975 10857
rect 8909 10789 8975 10823
rect 8909 10755 8925 10789
rect 8959 10755 8975 10789
rect 8909 10721 8975 10755
rect 8909 10687 8925 10721
rect 8959 10687 8975 10721
rect 8909 10653 8975 10687
rect 8909 10619 8925 10653
rect 8959 10619 8975 10653
rect 8909 10585 8975 10619
rect 8909 10551 8925 10585
rect 8959 10551 8975 10585
rect 8909 10517 8975 10551
rect 8909 10483 8925 10517
rect 8959 10483 8975 10517
rect 8909 10449 8975 10483
rect 8909 10415 8925 10449
rect 8959 10415 8975 10449
rect 8909 10381 8975 10415
rect 8909 10347 8925 10381
rect 8959 10347 8975 10381
rect 8909 10313 8975 10347
rect 8909 10279 8925 10313
rect 8959 10279 8975 10313
rect 8909 10245 8975 10279
rect 8909 10211 8925 10245
rect 8959 10211 8975 10245
rect 8909 10177 8975 10211
rect 8909 10143 8925 10177
rect 8959 10143 8975 10177
rect 8909 10109 8975 10143
rect 8909 10075 8925 10109
rect 8959 10075 8975 10109
rect 8909 10041 8975 10075
rect 8909 10007 8925 10041
rect 8959 10007 8975 10041
rect 8909 9973 8975 10007
rect 8909 9939 8925 9973
rect 8959 9939 8975 9973
rect 8909 9905 8975 9939
rect 8909 9871 8925 9905
rect 8959 9871 8975 9905
rect 8909 9837 8975 9871
rect 8909 9803 8925 9837
rect 8959 9803 8975 9837
rect 8909 9769 8975 9803
rect 8909 9735 8925 9769
rect 8959 9735 8975 9769
rect 8909 9701 8975 9735
rect 8909 9667 8925 9701
rect 8959 9667 8975 9701
rect 8909 9633 8975 9667
rect 8909 9599 8925 9633
rect 8959 9599 8975 9633
rect 8909 9565 8975 9599
rect 8909 9531 8925 9565
rect 8959 9531 8975 9565
rect 8909 9497 8975 9531
rect 8909 9463 8925 9497
rect 8959 9463 8975 9497
rect 8909 9429 8975 9463
rect 8909 9395 8925 9429
rect 8959 9395 8975 9429
rect 8909 9361 8975 9395
rect 8909 9327 8925 9361
rect 8959 9327 8975 9361
rect 8909 9293 8975 9327
rect 8909 9259 8925 9293
rect 8959 9259 8975 9293
rect 8909 9225 8975 9259
rect 8909 9191 8925 9225
rect 8959 9191 8975 9225
rect 8909 9157 8975 9191
rect 8909 9123 8925 9157
rect 8959 9123 8975 9157
rect 8909 9089 8975 9123
rect 8909 9055 8925 9089
rect 8959 9055 8975 9089
rect 8909 9021 8975 9055
rect 8909 8987 8925 9021
rect 8959 8987 8975 9021
rect 8909 8953 8975 8987
rect 8909 8919 8925 8953
rect 8959 8919 8975 8953
rect 8909 8885 8975 8919
rect 8909 8851 8925 8885
rect 8959 8851 8975 8885
rect 8909 8817 8975 8851
rect 8909 8783 8925 8817
rect 8959 8783 8975 8817
rect 8909 8749 8975 8783
rect 8909 8715 8925 8749
rect 8959 8715 8975 8749
rect 8909 8681 8975 8715
rect 8909 8647 8925 8681
rect 8959 8647 8975 8681
rect 8909 8613 8975 8647
rect 8909 8579 8925 8613
rect 8959 8579 8975 8613
rect 8909 8545 8975 8579
rect 8909 8511 8925 8545
rect 8959 8511 8975 8545
rect 8909 8477 8975 8511
rect 8909 8443 8925 8477
rect 8959 8443 8975 8477
rect 8909 8409 8975 8443
rect 8909 8375 8925 8409
rect 8959 8375 8975 8409
rect 8909 8341 8975 8375
rect 8909 8307 8925 8341
rect 8959 8307 8975 8341
rect 8909 8273 8975 8307
rect 8909 8239 8925 8273
rect 8959 8239 8975 8273
rect 8909 8205 8975 8239
rect 8909 8171 8925 8205
rect 8959 8171 8975 8205
rect 8909 8137 8975 8171
rect 8909 8103 8925 8137
rect 8959 8103 8975 8137
rect 8909 8069 8975 8103
rect 8909 8035 8925 8069
rect 8959 8035 8975 8069
rect 8909 8001 8975 8035
rect 8909 7967 8925 8001
rect 8959 7967 8975 8001
rect 8909 7933 8975 7967
rect 8909 7899 8925 7933
rect 8959 7899 8975 7933
rect 8909 7865 8975 7899
rect 8909 7831 8925 7865
rect 8959 7831 8975 7865
rect 8909 7797 8975 7831
rect 8909 7763 8925 7797
rect 8959 7763 8975 7797
rect 8909 7729 8975 7763
rect 8909 7695 8925 7729
rect 8959 7695 8975 7729
rect 8909 7661 8975 7695
rect 8909 7627 8925 7661
rect 8959 7627 8975 7661
rect 8909 7593 8975 7627
rect 8909 7559 8925 7593
rect 8959 7559 8975 7593
rect 8909 7525 8975 7559
rect 8909 7491 8925 7525
rect 8959 7491 8975 7525
rect 8909 7457 8975 7491
rect 8909 7423 8925 7457
rect 8959 7423 8975 7457
rect 8909 7389 8975 7423
rect 8909 7355 8925 7389
rect 8959 7355 8975 7389
rect 8909 7321 8975 7355
rect 8909 7287 8925 7321
rect 8959 7287 8975 7321
rect 8909 7253 8975 7287
rect 8909 7219 8925 7253
rect 8959 7219 8975 7253
rect 8909 7185 8975 7219
rect 8909 7151 8925 7185
rect 8959 7151 8975 7185
rect 8909 7117 8975 7151
rect 8909 7083 8925 7117
rect 8959 7083 8975 7117
rect 8909 7049 8975 7083
rect 8909 7015 8925 7049
rect 8959 7015 8975 7049
rect 8909 6981 8975 7015
rect 8909 6947 8925 6981
rect 8959 6947 8975 6981
rect 8909 6913 8975 6947
rect 8909 6879 8925 6913
rect 8959 6879 8975 6913
rect 8909 6845 8975 6879
rect 8909 6811 8925 6845
rect 8959 6811 8975 6845
rect 8909 6777 8975 6811
rect 8909 6743 8925 6777
rect 8959 6743 8975 6777
rect 8909 6709 8975 6743
rect 8909 6675 8925 6709
rect 8959 6675 8975 6709
rect 8909 6641 8975 6675
rect 8909 6607 8925 6641
rect 8959 6607 8975 6641
rect 8909 6573 8975 6607
rect 8909 6539 8925 6573
rect 8959 6539 8975 6573
rect 8909 6505 8975 6539
rect 8909 6471 8925 6505
rect 8959 6471 8975 6505
rect 8909 6437 8975 6471
rect 8909 6403 8925 6437
rect 8959 6403 8975 6437
rect 8909 6369 8975 6403
rect 8909 6335 8925 6369
rect 8959 6335 8975 6369
rect 8909 6301 8975 6335
rect 8909 6267 8925 6301
rect 8959 6267 8975 6301
rect 8909 6233 8975 6267
rect 8909 6199 8925 6233
rect 8959 6199 8975 6233
rect 8909 6165 8975 6199
rect 8909 6131 8925 6165
rect 8959 6131 8975 6165
rect 8909 6097 8975 6131
rect 8909 6063 8925 6097
rect 8959 6063 8975 6097
rect 8909 6029 8975 6063
rect 8909 5995 8925 6029
rect 8959 5995 8975 6029
rect 8909 5961 8975 5995
rect 8909 5927 8925 5961
rect 8959 5927 8975 5961
rect 8909 5893 8975 5927
rect 8909 5859 8925 5893
rect 8959 5859 8975 5893
rect 8909 5825 8975 5859
rect 8909 5791 8925 5825
rect 8959 5791 8975 5825
rect 8909 5757 8975 5791
rect 8909 5723 8925 5757
rect 8959 5723 8975 5757
rect 8909 5689 8975 5723
rect 8909 5655 8925 5689
rect 8959 5655 8975 5689
rect 8909 5621 8975 5655
rect 8909 5587 8925 5621
rect 8959 5587 8975 5621
rect 8909 5553 8975 5587
rect 8909 5519 8925 5553
rect 8959 5519 8975 5553
rect 8909 5485 8975 5519
rect 8909 5451 8925 5485
rect 8959 5451 8975 5485
rect 8909 5417 8975 5451
rect 8909 5383 8925 5417
rect 8959 5383 8975 5417
rect 8909 5349 8975 5383
rect 8909 5315 8925 5349
rect 8959 5315 8975 5349
rect 8909 5281 8975 5315
rect 8909 5247 8925 5281
rect 8959 5247 8975 5281
rect 8909 5213 8975 5247
rect 8909 5179 8925 5213
rect 8959 5179 8975 5213
rect 8909 5145 8975 5179
rect 8909 5111 8925 5145
rect 8959 5111 8975 5145
rect 8909 5077 8975 5111
rect 8909 5043 8925 5077
rect 8959 5043 8975 5077
rect 8909 5009 8975 5043
rect 8909 4975 8925 5009
rect 8959 4975 8975 5009
rect 8909 4941 8975 4975
rect 8909 4907 8925 4941
rect 8959 4907 8975 4941
rect 8909 4873 8975 4907
rect 8909 4839 8925 4873
rect 8959 4839 8975 4873
rect 8909 4805 8975 4839
rect 8909 4771 8925 4805
rect 8959 4771 8975 4805
rect 8909 4737 8975 4771
rect 8909 4703 8925 4737
rect 8959 4703 8975 4737
rect 8909 4669 8975 4703
rect 8909 4635 8925 4669
rect 8959 4635 8975 4669
rect 8909 4601 8975 4635
rect 8909 4567 8925 4601
rect 8959 4567 8975 4601
rect 8909 4533 8975 4567
rect 8909 4499 8925 4533
rect 8959 4499 8975 4533
rect 8909 4465 8975 4499
rect 8909 4431 8925 4465
rect 8959 4431 8975 4465
rect 8909 4397 8975 4431
rect 8909 4363 8925 4397
rect 8959 4363 8975 4397
rect 8909 4329 8975 4363
rect 8909 4295 8925 4329
rect 8959 4295 8975 4329
rect 8909 4261 8975 4295
rect 8909 4227 8925 4261
rect 8959 4227 8975 4261
rect 8909 4193 8975 4227
rect 8909 4159 8925 4193
rect 8959 4159 8975 4193
rect 8909 4125 8975 4159
rect 8909 4091 8925 4125
rect 8959 4091 8975 4125
rect 8909 4057 8975 4091
rect 8909 4023 8925 4057
rect 8959 4023 8975 4057
rect 8909 3989 8975 4023
rect 8909 3955 8925 3989
rect 8959 3955 8975 3989
rect 8909 3921 8975 3955
rect 8909 3887 8925 3921
rect 8959 3887 8975 3921
rect 8909 3853 8975 3887
rect 8909 3819 8925 3853
rect 8959 3819 8975 3853
rect 8909 3785 8975 3819
rect 8909 3751 8925 3785
rect 8959 3751 8975 3785
rect 8909 3717 8975 3751
rect 8909 3683 8925 3717
rect 8959 3683 8975 3717
rect 8909 3649 8975 3683
rect 8909 3615 8925 3649
rect 8959 3615 8975 3649
rect 8909 3581 8975 3615
rect 8909 3547 8925 3581
rect 8959 3547 8975 3581
rect 8909 3513 8975 3547
rect 8909 3479 8925 3513
rect 8959 3479 8975 3513
rect 8909 3445 8975 3479
rect 8909 3411 8925 3445
rect 8959 3411 8975 3445
rect 8909 3377 8975 3411
rect 8909 3343 8925 3377
rect 8959 3343 8975 3377
rect 8909 3309 8975 3343
rect 8909 3275 8925 3309
rect 8959 3275 8975 3309
rect 8909 3241 8975 3275
rect 8909 3207 8925 3241
rect 8959 3207 8975 3241
rect 8909 3173 8975 3207
rect 8909 3139 8925 3173
rect 8959 3139 8975 3173
rect 8909 3105 8975 3139
rect 8909 3071 8925 3105
rect 8959 3071 8975 3105
rect 8909 3037 8975 3071
rect 8909 3003 8925 3037
rect 8959 3003 8975 3037
rect 8909 2969 8975 3003
rect 8909 2935 8925 2969
rect 8959 2935 8975 2969
rect 8909 2901 8975 2935
rect 8909 2867 8925 2901
rect 8959 2867 8975 2901
rect 8909 2833 8975 2867
rect 8909 2799 8925 2833
rect 8959 2799 8975 2833
rect 8909 2765 8975 2799
rect 8909 2731 8925 2765
rect 8959 2731 8975 2765
rect 8909 2697 8975 2731
rect 8909 2663 8925 2697
rect 8959 2663 8975 2697
rect 8909 2629 8975 2663
rect 8909 2595 8925 2629
rect 8959 2595 8975 2629
rect 8909 2561 8975 2595
rect 8909 2527 8925 2561
rect 8959 2527 8975 2561
rect 8909 2493 8975 2527
rect 8909 2459 8925 2493
rect 8959 2459 8975 2493
rect 8909 2425 8975 2459
rect 8909 2391 8925 2425
rect 8959 2391 8975 2425
rect 8909 2357 8975 2391
rect 8909 2323 8925 2357
rect 8959 2323 8975 2357
rect 8909 2289 8975 2323
rect 8909 2255 8925 2289
rect 8959 2255 8975 2289
rect 8909 2221 8975 2255
rect 8909 2187 8925 2221
rect 8959 2187 8975 2221
rect 8909 2153 8975 2187
rect 8909 2119 8925 2153
rect 8959 2119 8975 2153
rect 8909 2085 8975 2119
rect 2310 1637 2452 1653
rect 2310 1603 2326 1637
rect 2360 1603 2402 1637
rect 2436 1603 2452 1637
rect 2310 1587 2452 1603
rect 2508 1637 2708 1653
rect 2508 1603 2524 1637
rect 2558 1603 2658 1637
rect 2692 1603 2708 1637
rect 2508 1587 2708 1603
rect 2764 1637 2964 1653
rect 2764 1603 2780 1637
rect 2814 1603 2914 1637
rect 2948 1603 2964 1637
rect 2764 1587 2964 1603
rect 3020 1637 3220 1653
rect 3020 1603 3036 1637
rect 3070 1603 3170 1637
rect 3204 1603 3220 1637
rect 3020 1587 3220 1603
rect 3276 1637 3476 1653
rect 3276 1603 3292 1637
rect 3326 1603 3426 1637
rect 3460 1603 3476 1637
rect 3276 1587 3476 1603
rect 3532 1637 3674 1653
rect 3532 1603 3548 1637
rect 3582 1603 3624 1637
rect 3658 1603 3674 1637
rect 3532 1587 3674 1603
rect 8909 2051 8925 2085
rect 8959 2051 8975 2085
rect 8909 2017 8975 2051
rect 8909 1983 8925 2017
rect 8959 1983 8975 2017
rect 8909 1949 8975 1983
rect 8909 1915 8925 1949
rect 8959 1915 8975 1949
rect 8909 1881 8975 1915
rect 8909 1847 8925 1881
rect 8959 1847 8975 1881
rect 8909 1813 8975 1847
rect 8909 1779 8925 1813
rect 8959 1779 8975 1813
rect 8909 1745 8975 1779
rect 8909 1711 8925 1745
rect 8959 1711 8975 1745
rect 8909 1677 8975 1711
rect 8909 1643 8925 1677
rect 8959 1643 8975 1677
rect 8909 1609 8975 1643
rect 8909 1575 8925 1609
rect 8959 1575 8975 1609
rect 8909 1541 8975 1575
rect 8909 1507 8925 1541
rect 8959 1507 8975 1541
rect 8909 1473 8975 1507
rect 8909 1439 8925 1473
rect 8959 1439 8975 1473
rect 8909 1405 8975 1439
rect 8909 1371 8925 1405
rect 8959 1371 8975 1405
rect 8024 1253 8180 1269
rect 8024 1219 8050 1253
rect 8084 1219 8126 1253
rect 8160 1219 8180 1253
rect 8024 1203 8180 1219
rect 8024 1197 8074 1203
rect 8130 1197 8180 1203
rect 8909 1337 8975 1371
rect 8909 1303 8925 1337
rect 8959 1303 8975 1337
rect 8909 1269 8975 1303
rect 8909 1235 8925 1269
rect 8959 1235 8975 1269
rect 8909 1201 8975 1235
rect 8909 1167 8925 1201
rect 8959 1167 8975 1201
rect 8909 1133 8975 1167
rect 8909 1099 8925 1133
rect 8959 1099 8975 1133
rect 8909 1065 8975 1099
rect 8909 1031 8925 1065
rect 8959 1031 8975 1065
rect 8909 997 8975 1031
rect 8909 963 8925 997
rect 8959 963 8975 997
rect 8909 929 8975 963
rect 8909 895 8925 929
rect 8959 895 8975 929
rect 8909 861 8975 895
rect 8909 827 8925 861
rect 8959 827 8975 861
rect 8909 793 8975 827
rect 8909 759 8925 793
rect 8959 759 8975 793
rect 8909 725 8975 759
rect 8909 691 8925 725
rect 8959 691 8975 725
rect 8909 657 8975 691
rect 8909 623 8925 657
rect 8959 623 8975 657
rect 8909 589 8975 623
rect 8909 555 8925 589
rect 8959 555 8975 589
rect 8909 521 8975 555
rect 8909 487 8925 521
rect 8959 487 8975 521
rect 8909 453 8975 487
rect 8909 419 8925 453
rect 8959 419 8975 453
rect 8909 385 8975 419
rect 8909 351 8925 385
rect 8959 351 8975 385
rect 8909 317 8975 351
rect 8909 283 8925 317
rect 8959 283 8975 317
rect 8909 249 8975 283
rect 8909 215 8925 249
rect 8959 215 8975 249
rect 8909 181 8975 215
rect 8909 147 8925 181
rect 8959 147 8975 181
rect 8909 113 8975 147
rect 8909 79 8925 113
rect 8959 79 8975 113
rect 8909 45 8975 79
rect 8909 11 8925 45
rect 8959 11 8975 45
rect 8909 -23 8975 11
rect 8909 -57 8925 -23
rect 8959 -57 8975 -23
rect 8909 -91 8975 -57
rect 8909 -125 8925 -91
rect 8959 -125 8975 -91
rect 8909 -159 8975 -125
rect 8909 -193 8925 -159
rect 8959 -193 8975 -159
rect 8909 -227 8975 -193
rect 8909 -261 8925 -227
rect 8959 -261 8975 -227
rect 8909 -295 8975 -261
rect 8909 -329 8925 -295
rect 8959 -329 8975 -295
rect 8909 -363 8975 -329
rect 8909 -397 8925 -363
rect 8959 -397 8975 -363
rect 8909 -431 8975 -397
rect 8909 -465 8925 -431
rect 8959 -465 8975 -431
rect 8909 -499 8975 -465
rect 8909 -533 8925 -499
rect 8959 -533 8975 -499
rect 8909 -567 8975 -533
rect 8909 -601 8925 -567
rect 8959 -601 8975 -567
rect 8909 -635 8975 -601
rect 8909 -669 8925 -635
rect 8959 -669 8975 -635
rect 8909 -703 8975 -669
rect 8909 -737 8925 -703
rect 8959 -737 8975 -703
rect 8909 -771 8975 -737
rect 8909 -805 8925 -771
rect 8959 -805 8975 -771
rect 8909 -839 8975 -805
rect 8909 -873 8925 -839
rect 8959 -873 8975 -839
rect 8909 -907 8975 -873
rect 8909 -941 8925 -907
rect 8959 -941 8975 -907
rect 8909 -975 8975 -941
rect 8909 -1009 8925 -975
rect 8959 -1009 8975 -975
rect 8909 -1043 8975 -1009
rect 8909 -1077 8925 -1043
rect 8959 -1077 8975 -1043
rect 8909 -1111 8975 -1077
rect 8909 -1145 8925 -1111
rect 8959 -1145 8975 -1111
rect 8909 -1179 8975 -1145
rect 8909 -1213 8925 -1179
rect 8959 -1213 8975 -1179
rect 8909 -1247 8975 -1213
rect 8909 -1281 8925 -1247
rect 8959 -1281 8975 -1247
rect 8909 -1315 8975 -1281
rect 8909 -1349 8925 -1315
rect 8959 -1349 8975 -1315
rect 8909 -1383 8975 -1349
rect 8909 -1417 8925 -1383
rect 8959 -1417 8975 -1383
rect 8909 -1451 8975 -1417
rect 8909 -1485 8925 -1451
rect 8959 -1485 8975 -1451
rect 8909 -1519 8975 -1485
rect 8909 -1553 8925 -1519
rect 8959 -1553 8975 -1519
rect 8909 -1587 8975 -1553
rect 8909 -1621 8925 -1587
rect 8959 -1621 8975 -1587
rect 8909 -1655 8975 -1621
rect 8909 -1689 8925 -1655
rect 8959 -1689 8975 -1655
rect 8909 -1723 8975 -1689
rect 8909 -1757 8925 -1723
rect 8959 -1757 8975 -1723
rect 8909 -1791 8975 -1757
rect 8909 -1825 8925 -1791
rect 8959 -1825 8975 -1791
rect 8909 -1859 8975 -1825
rect 8909 -1893 8925 -1859
rect 8959 -1893 8975 -1859
rect 8909 -1927 8975 -1893
rect 8909 -1961 8925 -1927
rect 8959 -1961 8975 -1927
rect 8909 -1995 8975 -1961
rect 8909 -2029 8925 -1995
rect 8959 -2029 8975 -1995
rect 8909 -2064 8975 -2029
rect 8909 -2098 8925 -2064
rect 8959 -2098 8975 -2064
rect 8909 -2133 8975 -2098
rect 8909 -2167 8925 -2133
rect 8959 -2167 8975 -2133
rect 8909 -2202 8975 -2167
rect 8909 -2236 8925 -2202
rect 8959 -2236 8975 -2202
rect 8909 -2271 8975 -2236
rect 8909 -2305 8925 -2271
rect 8959 -2305 8975 -2271
rect 8909 -2340 8975 -2305
rect 8909 -2374 8925 -2340
rect 8959 -2374 8975 -2340
rect 8909 -2409 8975 -2374
rect 8909 -2443 8925 -2409
rect 8959 -2443 8975 -2409
rect 8909 -2478 8975 -2443
rect 8909 -2512 8925 -2478
rect 8959 -2512 8975 -2478
rect 8909 -2547 8975 -2512
rect 8909 -2581 8925 -2547
rect 8959 -2581 8975 -2547
rect 8909 -2616 8975 -2581
rect 8909 -2650 8925 -2616
rect 8959 -2650 8975 -2616
rect 8909 -2685 8975 -2650
rect 8909 -2719 8925 -2685
rect 8959 -2719 8975 -2685
rect 8909 -2754 8975 -2719
rect 8909 -2788 8925 -2754
rect 8959 -2788 8975 -2754
rect 8909 -2823 8975 -2788
rect 8909 -2857 8925 -2823
rect 8959 -2857 8975 -2823
rect 8909 -2892 8975 -2857
rect 8909 -2926 8925 -2892
rect 8959 -2926 8975 -2892
rect 8909 -2961 8975 -2926
rect 8909 -2995 8925 -2961
rect 8959 -2995 8975 -2961
rect 8909 -3030 8975 -2995
rect 8909 -3064 8925 -3030
rect 8959 -3064 8975 -3030
rect 8909 -3099 8975 -3064
rect 8909 -3133 8925 -3099
rect 8959 -3133 8975 -3099
rect 8909 -3168 8975 -3133
rect 8909 -3202 8925 -3168
rect 8959 -3202 8975 -3168
rect 8909 -3237 8975 -3202
rect 8909 -3271 8925 -3237
rect 8959 -3271 8975 -3237
rect 8909 -3306 8975 -3271
rect 8909 -3340 8925 -3306
rect 8959 -3340 8975 -3306
rect 8909 -3375 8975 -3340
rect 8909 -3409 8925 -3375
rect 8959 -3409 8975 -3375
rect 8909 -3444 8975 -3409
rect 8909 -3478 8925 -3444
rect 8959 -3478 8975 -3444
rect 8909 -3513 8975 -3478
rect 8909 -3547 8925 -3513
rect 8959 -3547 8975 -3513
rect 8909 -3582 8975 -3547
rect 8909 -3616 8925 -3582
rect 8959 -3616 8975 -3582
rect 8909 -3651 8975 -3616
rect 8909 -3685 8925 -3651
rect 8959 -3685 8975 -3651
rect 8909 -3720 8975 -3685
rect 8909 -3754 8925 -3720
rect 8959 -3754 8975 -3720
rect 8909 -3789 8975 -3754
rect 8909 -3823 8925 -3789
rect 8959 -3823 8975 -3789
rect 8909 -3858 8975 -3823
rect 8909 -3892 8925 -3858
rect 8959 -3892 8975 -3858
rect 8909 -3927 8975 -3892
rect 8909 -3961 8925 -3927
rect 8959 -3929 8975 -3927
rect 10755 22145 10821 22179
rect 10755 22111 10771 22145
rect 10805 22111 10821 22145
rect 10755 22077 10821 22111
rect 10755 22043 10771 22077
rect 10805 22043 10821 22077
rect 10755 22009 10821 22043
rect 10755 21975 10771 22009
rect 10805 21975 10821 22009
rect 10755 21941 10821 21975
rect 10755 21907 10771 21941
rect 10805 21907 10821 21941
rect 10755 21873 10821 21907
rect 10755 21839 10771 21873
rect 10805 21839 10821 21873
rect 10755 21805 10821 21839
rect 10755 21771 10771 21805
rect 10805 21771 10821 21805
rect 10755 21737 10821 21771
rect 10755 21703 10771 21737
rect 10805 21703 10821 21737
rect 10755 21669 10821 21703
rect 10755 21635 10771 21669
rect 10805 21635 10821 21669
rect 10755 21601 10821 21635
rect 10755 21567 10771 21601
rect 10805 21567 10821 21601
rect 10755 21533 10821 21567
rect 10755 21499 10771 21533
rect 10805 21499 10821 21533
rect 10755 21465 10821 21499
rect 10755 21431 10771 21465
rect 10805 21431 10821 21465
rect 10755 21397 10821 21431
rect 10755 21363 10771 21397
rect 10805 21363 10821 21397
rect 10755 21329 10821 21363
rect 10755 21295 10771 21329
rect 10805 21295 10821 21329
rect 10755 21261 10821 21295
rect 10755 21227 10771 21261
rect 10805 21227 10821 21261
rect 10755 21193 10821 21227
rect 10755 21159 10771 21193
rect 10805 21159 10821 21193
rect 10755 21125 10821 21159
rect 10755 21091 10771 21125
rect 10805 21091 10821 21125
rect 10755 21057 10821 21091
rect 10755 21023 10771 21057
rect 10805 21023 10821 21057
rect 10755 20989 10821 21023
rect 10755 20955 10771 20989
rect 10805 20955 10821 20989
rect 10755 20921 10821 20955
rect 10755 20887 10771 20921
rect 10805 20887 10821 20921
rect 10755 20853 10821 20887
rect 10755 20819 10771 20853
rect 10805 20819 10821 20853
rect 10755 20785 10821 20819
rect 10755 20751 10771 20785
rect 10805 20751 10821 20785
rect 10755 20717 10821 20751
rect 10755 20683 10771 20717
rect 10805 20683 10821 20717
rect 10755 20649 10821 20683
rect 10755 20615 10771 20649
rect 10805 20615 10821 20649
rect 10755 20581 10821 20615
rect 10755 20547 10771 20581
rect 10805 20547 10821 20581
rect 10755 20513 10821 20547
rect 10755 20479 10771 20513
rect 10805 20479 10821 20513
rect 10755 20445 10821 20479
rect 10755 20411 10771 20445
rect 10805 20411 10821 20445
rect 10755 20377 10821 20411
rect 10755 20343 10771 20377
rect 10805 20343 10821 20377
rect 10755 20309 10821 20343
rect 10755 20275 10771 20309
rect 10805 20275 10821 20309
rect 10755 20241 10821 20275
rect 10755 20207 10771 20241
rect 10805 20207 10821 20241
rect 10755 20173 10821 20207
rect 10755 20139 10771 20173
rect 10805 20139 10821 20173
rect 10755 20105 10821 20139
rect 10755 20071 10771 20105
rect 10805 20071 10821 20105
rect 10755 20037 10821 20071
rect 10755 20003 10771 20037
rect 10805 20003 10821 20037
rect 10755 19969 10821 20003
rect 10755 19935 10771 19969
rect 10805 19935 10821 19969
rect 10755 19901 10821 19935
rect 10755 19867 10771 19901
rect 10805 19867 10821 19901
rect 10755 19833 10821 19867
rect 10755 19799 10771 19833
rect 10805 19799 10821 19833
rect 10755 19765 10821 19799
rect 10755 19731 10771 19765
rect 10805 19731 10821 19765
rect 10755 19697 10821 19731
rect 10755 19663 10771 19697
rect 10805 19663 10821 19697
rect 10755 19629 10821 19663
rect 10755 19595 10771 19629
rect 10805 19595 10821 19629
rect 10755 19561 10821 19595
rect 10755 19527 10771 19561
rect 10805 19527 10821 19561
rect 10755 19493 10821 19527
rect 10755 19459 10771 19493
rect 10805 19459 10821 19493
rect 10755 19425 10821 19459
rect 10755 19391 10771 19425
rect 10805 19391 10821 19425
rect 10755 19357 10821 19391
rect 10755 19323 10771 19357
rect 10805 19323 10821 19357
rect 10755 19289 10821 19323
rect 10755 19255 10771 19289
rect 10805 19255 10821 19289
rect 10755 19221 10821 19255
rect 10755 19187 10771 19221
rect 10805 19187 10821 19221
rect 10755 19153 10821 19187
rect 10755 19119 10771 19153
rect 10805 19119 10821 19153
rect 10755 19085 10821 19119
rect 10755 19051 10771 19085
rect 10805 19051 10821 19085
rect 10755 19017 10821 19051
rect 10755 18983 10771 19017
rect 10805 18983 10821 19017
rect 10755 18949 10821 18983
rect 10755 18915 10771 18949
rect 10805 18915 10821 18949
rect 10755 18881 10821 18915
rect 10755 18847 10771 18881
rect 10805 18847 10821 18881
rect 10755 18813 10821 18847
rect 10755 18779 10771 18813
rect 10805 18779 10821 18813
rect 10755 18745 10821 18779
rect 10755 18711 10771 18745
rect 10805 18711 10821 18745
rect 10755 18677 10821 18711
rect 10755 18643 10771 18677
rect 10805 18643 10821 18677
rect 10755 18609 10821 18643
rect 10755 18575 10771 18609
rect 10805 18575 10821 18609
rect 10755 18541 10821 18575
rect 10755 18507 10771 18541
rect 10805 18507 10821 18541
rect 10755 18473 10821 18507
rect 10755 18439 10771 18473
rect 10805 18439 10821 18473
rect 10755 18405 10821 18439
rect 10755 18371 10771 18405
rect 10805 18371 10821 18405
rect 10755 18337 10821 18371
rect 10755 18303 10771 18337
rect 10805 18303 10821 18337
rect 10755 18269 10821 18303
rect 10755 18235 10771 18269
rect 10805 18235 10821 18269
rect 10755 18201 10821 18235
rect 10755 18167 10771 18201
rect 10805 18167 10821 18201
rect 10755 18133 10821 18167
rect 10755 18099 10771 18133
rect 10805 18099 10821 18133
rect 10755 18065 10821 18099
rect 10755 18031 10771 18065
rect 10805 18031 10821 18065
rect 10755 17997 10821 18031
rect 10755 17963 10771 17997
rect 10805 17963 10821 17997
rect 10755 17929 10821 17963
rect 10755 17895 10771 17929
rect 10805 17895 10821 17929
rect 10755 17861 10821 17895
rect 10755 17827 10771 17861
rect 10805 17827 10821 17861
rect 10755 17793 10821 17827
rect 10755 17759 10771 17793
rect 10805 17759 10821 17793
rect 10755 17725 10821 17759
rect 10755 17691 10771 17725
rect 10805 17691 10821 17725
rect 10755 17657 10821 17691
rect 10755 17623 10771 17657
rect 10805 17623 10821 17657
rect 10755 17589 10821 17623
rect 10755 17555 10771 17589
rect 10805 17555 10821 17589
rect 10755 17521 10821 17555
rect 10755 17487 10771 17521
rect 10805 17487 10821 17521
rect 10755 17453 10821 17487
rect 10755 17419 10771 17453
rect 10805 17419 10821 17453
rect 10755 17385 10821 17419
rect 10755 17351 10771 17385
rect 10805 17351 10821 17385
rect 10755 17317 10821 17351
rect 10755 17283 10771 17317
rect 10805 17283 10821 17317
rect 10755 17249 10821 17283
rect 10755 17215 10771 17249
rect 10805 17215 10821 17249
rect 10755 17181 10821 17215
rect 10755 17147 10771 17181
rect 10805 17147 10821 17181
rect 10755 17113 10821 17147
rect 10755 17079 10771 17113
rect 10805 17079 10821 17113
rect 10755 17045 10821 17079
rect 10755 17011 10771 17045
rect 10805 17011 10821 17045
rect 10755 16977 10821 17011
rect 10755 16943 10771 16977
rect 10805 16943 10821 16977
rect 10755 16909 10821 16943
rect 10755 16875 10771 16909
rect 10805 16875 10821 16909
rect 10755 16841 10821 16875
rect 10755 16807 10771 16841
rect 10805 16807 10821 16841
rect 10755 16773 10821 16807
rect 10755 16739 10771 16773
rect 10805 16739 10821 16773
rect 10755 16705 10821 16739
rect 10755 16671 10771 16705
rect 10805 16671 10821 16705
rect 10755 16637 10821 16671
rect 10755 16603 10771 16637
rect 10805 16603 10821 16637
rect 10755 16569 10821 16603
rect 10755 16535 10771 16569
rect 10805 16535 10821 16569
rect 10755 16501 10821 16535
rect 10755 16467 10771 16501
rect 10805 16467 10821 16501
rect 10755 16433 10821 16467
rect 10755 16399 10771 16433
rect 10805 16399 10821 16433
rect 10755 16365 10821 16399
rect 10755 16331 10771 16365
rect 10805 16331 10821 16365
rect 10755 16297 10821 16331
rect 10755 16263 10771 16297
rect 10805 16263 10821 16297
rect 10755 16229 10821 16263
rect 10755 16195 10771 16229
rect 10805 16195 10821 16229
rect 10755 16161 10821 16195
rect 10755 16127 10771 16161
rect 10805 16127 10821 16161
rect 10755 16093 10821 16127
rect 10755 16059 10771 16093
rect 10805 16059 10821 16093
rect 10755 16025 10821 16059
rect 10755 15991 10771 16025
rect 10805 15991 10821 16025
rect 10755 15957 10821 15991
rect 10755 15923 10771 15957
rect 10805 15923 10821 15957
rect 10755 15889 10821 15923
rect 10755 15855 10771 15889
rect 10805 15855 10821 15889
rect 10755 15821 10821 15855
rect 10755 15787 10771 15821
rect 10805 15787 10821 15821
rect 10755 15753 10821 15787
rect 10755 15719 10771 15753
rect 10805 15719 10821 15753
rect 10755 15685 10821 15719
rect 10755 15651 10771 15685
rect 10805 15651 10821 15685
rect 10755 15617 10821 15651
rect 10755 15583 10771 15617
rect 10805 15583 10821 15617
rect 10755 15549 10821 15583
rect 10755 15515 10771 15549
rect 10805 15515 10821 15549
rect 10755 15481 10821 15515
rect 10755 15447 10771 15481
rect 10805 15447 10821 15481
rect 10755 15413 10821 15447
rect 10755 15379 10771 15413
rect 10805 15379 10821 15413
rect 10755 15345 10821 15379
rect 10755 15311 10771 15345
rect 10805 15311 10821 15345
rect 10755 15277 10821 15311
rect 10755 15243 10771 15277
rect 10805 15243 10821 15277
rect 10755 15209 10821 15243
rect 10755 15175 10771 15209
rect 10805 15175 10821 15209
rect 10755 15141 10821 15175
rect 10755 15107 10771 15141
rect 10805 15107 10821 15141
rect 10755 15073 10821 15107
rect 10755 15039 10771 15073
rect 10805 15039 10821 15073
rect 10755 15005 10821 15039
rect 10755 14971 10771 15005
rect 10805 14971 10821 15005
rect 10755 14937 10821 14971
rect 10755 14903 10771 14937
rect 10805 14903 10821 14937
rect 10755 14869 10821 14903
rect 10755 14835 10771 14869
rect 10805 14835 10821 14869
rect 10755 14801 10821 14835
rect 10755 14767 10771 14801
rect 10805 14767 10821 14801
rect 10755 14733 10821 14767
rect 10755 14699 10771 14733
rect 10805 14699 10821 14733
rect 10755 14665 10821 14699
rect 10755 14631 10771 14665
rect 10805 14631 10821 14665
rect 10755 14597 10821 14631
rect 10755 14563 10771 14597
rect 10805 14563 10821 14597
rect 10755 14529 10821 14563
rect 10755 14495 10771 14529
rect 10805 14495 10821 14529
rect 10755 14461 10821 14495
rect 10755 14427 10771 14461
rect 10805 14427 10821 14461
rect 10755 14393 10821 14427
rect 10755 14359 10771 14393
rect 10805 14359 10821 14393
rect 10755 14325 10821 14359
rect 10755 14291 10771 14325
rect 10805 14291 10821 14325
rect 10755 14257 10821 14291
rect 10755 14223 10771 14257
rect 10805 14223 10821 14257
rect 10755 14189 10821 14223
rect 10755 14155 10771 14189
rect 10805 14155 10821 14189
rect 10755 14121 10821 14155
rect 10755 14087 10771 14121
rect 10805 14087 10821 14121
rect 10755 14053 10821 14087
rect 10755 14019 10771 14053
rect 10805 14019 10821 14053
rect 10755 13985 10821 14019
rect 10755 13951 10771 13985
rect 10805 13951 10821 13985
rect 10755 13917 10821 13951
rect 10755 13883 10771 13917
rect 10805 13883 10821 13917
rect 10755 13849 10821 13883
rect 10755 13815 10771 13849
rect 10805 13815 10821 13849
rect 10755 13781 10821 13815
rect 10755 13747 10771 13781
rect 10805 13747 10821 13781
rect 10755 13713 10821 13747
rect 10755 13679 10771 13713
rect 10805 13679 10821 13713
rect 10755 13645 10821 13679
rect 10755 13611 10771 13645
rect 10805 13611 10821 13645
rect 10755 13577 10821 13611
rect 10755 13543 10771 13577
rect 10805 13543 10821 13577
rect 10755 13509 10821 13543
rect 10755 13475 10771 13509
rect 10805 13475 10821 13509
rect 10755 13441 10821 13475
rect 10755 13407 10771 13441
rect 10805 13407 10821 13441
rect 10755 13373 10821 13407
rect 10755 13339 10771 13373
rect 10805 13339 10821 13373
rect 10755 13305 10821 13339
rect 10755 13271 10771 13305
rect 10805 13271 10821 13305
rect 10755 13237 10821 13271
rect 10755 13203 10771 13237
rect 10805 13203 10821 13237
rect 10755 13169 10821 13203
rect 10755 13135 10771 13169
rect 10805 13135 10821 13169
rect 10755 13101 10821 13135
rect 10755 13067 10771 13101
rect 10805 13067 10821 13101
rect 10755 13033 10821 13067
rect 10755 12999 10771 13033
rect 10805 12999 10821 13033
rect 10755 12965 10821 12999
rect 10755 12931 10771 12965
rect 10805 12931 10821 12965
rect 10755 12897 10821 12931
rect 10755 12863 10771 12897
rect 10805 12863 10821 12897
rect 10755 12829 10821 12863
rect 10755 12795 10771 12829
rect 10805 12795 10821 12829
rect 10755 12761 10821 12795
rect 10755 12727 10771 12761
rect 10805 12727 10821 12761
rect 10755 12693 10821 12727
rect 10755 12659 10771 12693
rect 10805 12659 10821 12693
rect 10755 12625 10821 12659
rect 10755 12591 10771 12625
rect 10805 12591 10821 12625
rect 10755 12557 10821 12591
rect 10755 12523 10771 12557
rect 10805 12523 10821 12557
rect 10755 12489 10821 12523
rect 10755 12455 10771 12489
rect 10805 12455 10821 12489
rect 10755 12421 10821 12455
rect 10755 12387 10771 12421
rect 10805 12387 10821 12421
rect 10755 12353 10821 12387
rect 10755 12319 10771 12353
rect 10805 12319 10821 12353
rect 10755 12285 10821 12319
rect 10755 12251 10771 12285
rect 10805 12251 10821 12285
rect 10755 12217 10821 12251
rect 10755 12183 10771 12217
rect 10805 12183 10821 12217
rect 10755 12149 10821 12183
rect 10755 12115 10771 12149
rect 10805 12115 10821 12149
rect 10755 12081 10821 12115
rect 10755 12047 10771 12081
rect 10805 12047 10821 12081
rect 10755 12013 10821 12047
rect 10755 11979 10771 12013
rect 10805 11979 10821 12013
rect 10755 11945 10821 11979
rect 10755 11911 10771 11945
rect 10805 11911 10821 11945
rect 10755 11877 10821 11911
rect 10755 11843 10771 11877
rect 10805 11843 10821 11877
rect 10755 11809 10821 11843
rect 10755 11775 10771 11809
rect 10805 11775 10821 11809
rect 10755 11741 10821 11775
rect 10755 11707 10771 11741
rect 10805 11707 10821 11741
rect 10755 11673 10821 11707
rect 10755 11639 10771 11673
rect 10805 11639 10821 11673
rect 10755 11605 10821 11639
rect 10755 11571 10771 11605
rect 10805 11571 10821 11605
rect 10755 11537 10821 11571
rect 10755 11503 10771 11537
rect 10805 11503 10821 11537
rect 10755 11469 10821 11503
rect 10755 11435 10771 11469
rect 10805 11435 10821 11469
rect 10755 11401 10821 11435
rect 10755 11367 10771 11401
rect 10805 11367 10821 11401
rect 10755 11333 10821 11367
rect 10755 11299 10771 11333
rect 10805 11299 10821 11333
rect 10755 11265 10821 11299
rect 10755 11231 10771 11265
rect 10805 11231 10821 11265
rect 10755 11197 10821 11231
rect 10755 11163 10771 11197
rect 10805 11163 10821 11197
rect 10755 11129 10821 11163
rect 10755 11095 10771 11129
rect 10805 11095 10821 11129
rect 10755 11061 10821 11095
rect 10755 11027 10771 11061
rect 10805 11027 10821 11061
rect 10755 10993 10821 11027
rect 10755 10959 10771 10993
rect 10805 10959 10821 10993
rect 10755 10925 10821 10959
rect 10755 10891 10771 10925
rect 10805 10891 10821 10925
rect 10755 10857 10821 10891
rect 10755 10823 10771 10857
rect 10805 10823 10821 10857
rect 10755 10789 10821 10823
rect 10755 10755 10771 10789
rect 10805 10755 10821 10789
rect 10755 10721 10821 10755
rect 10755 10687 10771 10721
rect 10805 10687 10821 10721
rect 10755 10653 10821 10687
rect 10755 10619 10771 10653
rect 10805 10619 10821 10653
rect 10755 10585 10821 10619
rect 10755 10551 10771 10585
rect 10805 10551 10821 10585
rect 10755 10517 10821 10551
rect 10755 10483 10771 10517
rect 10805 10483 10821 10517
rect 10755 10449 10821 10483
rect 10755 10415 10771 10449
rect 10805 10415 10821 10449
rect 10755 10381 10821 10415
rect 10755 10347 10771 10381
rect 10805 10347 10821 10381
rect 10755 10313 10821 10347
rect 10755 10279 10771 10313
rect 10805 10279 10821 10313
rect 10755 10245 10821 10279
rect 10755 10211 10771 10245
rect 10805 10211 10821 10245
rect 10755 10177 10821 10211
rect 10755 10143 10771 10177
rect 10805 10143 10821 10177
rect 10755 10109 10821 10143
rect 10755 10075 10771 10109
rect 10805 10075 10821 10109
rect 10755 10041 10821 10075
rect 10755 10007 10771 10041
rect 10805 10007 10821 10041
rect 10755 9973 10821 10007
rect 10755 9939 10771 9973
rect 10805 9939 10821 9973
rect 10755 9905 10821 9939
rect 10755 9871 10771 9905
rect 10805 9871 10821 9905
rect 10755 9837 10821 9871
rect 10755 9803 10771 9837
rect 10805 9803 10821 9837
rect 10755 9769 10821 9803
rect 10755 9735 10771 9769
rect 10805 9735 10821 9769
rect 10755 9701 10821 9735
rect 10755 9667 10771 9701
rect 10805 9667 10821 9701
rect 10755 9633 10821 9667
rect 10755 9599 10771 9633
rect 10805 9599 10821 9633
rect 10755 9565 10821 9599
rect 10755 9531 10771 9565
rect 10805 9531 10821 9565
rect 10755 9497 10821 9531
rect 10755 9463 10771 9497
rect 10805 9463 10821 9497
rect 10755 9429 10821 9463
rect 10755 9395 10771 9429
rect 10805 9395 10821 9429
rect 10755 9361 10821 9395
rect 10755 9327 10771 9361
rect 10805 9327 10821 9361
rect 10755 9293 10821 9327
rect 10755 9259 10771 9293
rect 10805 9259 10821 9293
rect 10755 9225 10821 9259
rect 10755 9191 10771 9225
rect 10805 9191 10821 9225
rect 10755 9157 10821 9191
rect 10755 9123 10771 9157
rect 10805 9123 10821 9157
rect 10755 9089 10821 9123
rect 10755 9055 10771 9089
rect 10805 9055 10821 9089
rect 10755 9021 10821 9055
rect 10755 8987 10771 9021
rect 10805 8987 10821 9021
rect 10755 8953 10821 8987
rect 10755 8919 10771 8953
rect 10805 8919 10821 8953
rect 10755 8885 10821 8919
rect 10755 8851 10771 8885
rect 10805 8851 10821 8885
rect 10755 8817 10821 8851
rect 10755 8783 10771 8817
rect 10805 8783 10821 8817
rect 10755 8749 10821 8783
rect 10755 8715 10771 8749
rect 10805 8715 10821 8749
rect 10755 8681 10821 8715
rect 10755 8647 10771 8681
rect 10805 8647 10821 8681
rect 10755 8613 10821 8647
rect 10755 8579 10771 8613
rect 10805 8579 10821 8613
rect 10755 8545 10821 8579
rect 10755 8511 10771 8545
rect 10805 8511 10821 8545
rect 10755 8477 10821 8511
rect 10755 8443 10771 8477
rect 10805 8443 10821 8477
rect 10755 8409 10821 8443
rect 10755 8375 10771 8409
rect 10805 8375 10821 8409
rect 10755 8341 10821 8375
rect 10755 8307 10771 8341
rect 10805 8307 10821 8341
rect 10755 8273 10821 8307
rect 10755 8239 10771 8273
rect 10805 8239 10821 8273
rect 10755 8205 10821 8239
rect 10755 8171 10771 8205
rect 10805 8171 10821 8205
rect 10755 8137 10821 8171
rect 10755 8103 10771 8137
rect 10805 8103 10821 8137
rect 10755 8069 10821 8103
rect 10755 8035 10771 8069
rect 10805 8035 10821 8069
rect 10755 8001 10821 8035
rect 10755 7967 10771 8001
rect 10805 7967 10821 8001
rect 10755 7933 10821 7967
rect 10755 7899 10771 7933
rect 10805 7899 10821 7933
rect 10755 7865 10821 7899
rect 10755 7831 10771 7865
rect 10805 7831 10821 7865
rect 10755 7797 10821 7831
rect 10755 7763 10771 7797
rect 10805 7763 10821 7797
rect 10755 7729 10821 7763
rect 10755 7695 10771 7729
rect 10805 7695 10821 7729
rect 10755 7661 10821 7695
rect 10755 7627 10771 7661
rect 10805 7627 10821 7661
rect 10755 7593 10821 7627
rect 10755 7559 10771 7593
rect 10805 7559 10821 7593
rect 10755 7525 10821 7559
rect 10755 7491 10771 7525
rect 10805 7491 10821 7525
rect 10755 7457 10821 7491
rect 10755 7423 10771 7457
rect 10805 7423 10821 7457
rect 10755 7389 10821 7423
rect 10755 7355 10771 7389
rect 10805 7355 10821 7389
rect 10755 7321 10821 7355
rect 10755 7287 10771 7321
rect 10805 7287 10821 7321
rect 10755 7253 10821 7287
rect 10755 7219 10771 7253
rect 10805 7219 10821 7253
rect 10755 7185 10821 7219
rect 10755 7151 10771 7185
rect 10805 7151 10821 7185
rect 10755 7117 10821 7151
rect 10755 7083 10771 7117
rect 10805 7083 10821 7117
rect 10755 7049 10821 7083
rect 10755 7015 10771 7049
rect 10805 7015 10821 7049
rect 10755 6981 10821 7015
rect 10755 6947 10771 6981
rect 10805 6947 10821 6981
rect 10755 6913 10821 6947
rect 10755 6879 10771 6913
rect 10805 6879 10821 6913
rect 10755 6845 10821 6879
rect 10755 6811 10771 6845
rect 10805 6811 10821 6845
rect 10755 6777 10821 6811
rect 10755 6743 10771 6777
rect 10805 6743 10821 6777
rect 10755 6709 10821 6743
rect 10755 6675 10771 6709
rect 10805 6675 10821 6709
rect 10755 6641 10821 6675
rect 10755 6607 10771 6641
rect 10805 6607 10821 6641
rect 10755 6573 10821 6607
rect 10755 6539 10771 6573
rect 10805 6539 10821 6573
rect 10755 6505 10821 6539
rect 10755 6471 10771 6505
rect 10805 6471 10821 6505
rect 10755 6437 10821 6471
rect 10755 6403 10771 6437
rect 10805 6403 10821 6437
rect 10755 6369 10821 6403
rect 10755 6335 10771 6369
rect 10805 6335 10821 6369
rect 10755 6301 10821 6335
rect 10755 6267 10771 6301
rect 10805 6267 10821 6301
rect 10755 6233 10821 6267
rect 10755 6199 10771 6233
rect 10805 6199 10821 6233
rect 10755 6165 10821 6199
rect 10755 6131 10771 6165
rect 10805 6131 10821 6165
rect 10755 6097 10821 6131
rect 10755 6063 10771 6097
rect 10805 6063 10821 6097
rect 10755 6029 10821 6063
rect 10755 5995 10771 6029
rect 10805 5995 10821 6029
rect 10755 5961 10821 5995
rect 10755 5927 10771 5961
rect 10805 5927 10821 5961
rect 10755 5893 10821 5927
rect 10755 5859 10771 5893
rect 10805 5859 10821 5893
rect 10755 5825 10821 5859
rect 10755 5791 10771 5825
rect 10805 5791 10821 5825
rect 10755 5757 10821 5791
rect 10755 5723 10771 5757
rect 10805 5723 10821 5757
rect 10755 5689 10821 5723
rect 10755 5655 10771 5689
rect 10805 5655 10821 5689
rect 10755 5621 10821 5655
rect 10755 5587 10771 5621
rect 10805 5587 10821 5621
rect 10755 5553 10821 5587
rect 10755 5519 10771 5553
rect 10805 5519 10821 5553
rect 10755 5485 10821 5519
rect 10755 5451 10771 5485
rect 10805 5451 10821 5485
rect 10755 5417 10821 5451
rect 10755 5383 10771 5417
rect 10805 5383 10821 5417
rect 10755 5349 10821 5383
rect 10755 5315 10771 5349
rect 10805 5315 10821 5349
rect 10755 5281 10821 5315
rect 10755 5247 10771 5281
rect 10805 5247 10821 5281
rect 10755 5213 10821 5247
rect 10755 5179 10771 5213
rect 10805 5179 10821 5213
rect 10755 5145 10821 5179
rect 10755 5111 10771 5145
rect 10805 5111 10821 5145
rect 10755 5077 10821 5111
rect 10755 5043 10771 5077
rect 10805 5043 10821 5077
rect 10755 5009 10821 5043
rect 10755 4975 10771 5009
rect 10805 4975 10821 5009
rect 10755 4941 10821 4975
rect 10755 4907 10771 4941
rect 10805 4907 10821 4941
rect 10755 4873 10821 4907
rect 10755 4839 10771 4873
rect 10805 4839 10821 4873
rect 10755 4805 10821 4839
rect 10755 4771 10771 4805
rect 10805 4771 10821 4805
rect 10755 4737 10821 4771
rect 10755 4703 10771 4737
rect 10805 4703 10821 4737
rect 10755 4669 10821 4703
rect 10755 4635 10771 4669
rect 10805 4635 10821 4669
rect 10755 4601 10821 4635
rect 10755 4567 10771 4601
rect 10805 4567 10821 4601
rect 10755 4533 10821 4567
rect 10755 4499 10771 4533
rect 10805 4499 10821 4533
rect 10755 4465 10821 4499
rect 10755 4431 10771 4465
rect 10805 4431 10821 4465
rect 10755 4397 10821 4431
rect 10755 4363 10771 4397
rect 10805 4363 10821 4397
rect 10755 4329 10821 4363
rect 10755 4295 10771 4329
rect 10805 4295 10821 4329
rect 10755 4261 10821 4295
rect 10755 4227 10771 4261
rect 10805 4227 10821 4261
rect 10755 4193 10821 4227
rect 10755 4159 10771 4193
rect 10805 4159 10821 4193
rect 10755 4125 10821 4159
rect 10755 4091 10771 4125
rect 10805 4091 10821 4125
rect 10755 4057 10821 4091
rect 10755 4023 10771 4057
rect 10805 4023 10821 4057
rect 10755 3989 10821 4023
rect 10755 3955 10771 3989
rect 10805 3955 10821 3989
rect 10755 3921 10821 3955
rect 10755 3887 10771 3921
rect 10805 3887 10821 3921
rect 10755 3853 10821 3887
rect 10755 3819 10771 3853
rect 10805 3819 10821 3853
rect 10755 3785 10821 3819
rect 10755 3751 10771 3785
rect 10805 3751 10821 3785
rect 10755 3717 10821 3751
rect 10755 3683 10771 3717
rect 10805 3683 10821 3717
rect 10755 3649 10821 3683
rect 10755 3615 10771 3649
rect 10805 3615 10821 3649
rect 10755 3581 10821 3615
rect 10755 3547 10771 3581
rect 10805 3547 10821 3581
rect 10755 3513 10821 3547
rect 10755 3479 10771 3513
rect 10805 3479 10821 3513
rect 10755 3445 10821 3479
rect 10755 3411 10771 3445
rect 10805 3411 10821 3445
rect 10755 3377 10821 3411
rect 10755 3343 10771 3377
rect 10805 3343 10821 3377
rect 10755 3309 10821 3343
rect 10755 3275 10771 3309
rect 10805 3275 10821 3309
rect 10755 3241 10821 3275
rect 10755 3207 10771 3241
rect 10805 3207 10821 3241
rect 10755 3173 10821 3207
rect 10755 3139 10771 3173
rect 10805 3139 10821 3173
rect 10755 3105 10821 3139
rect 10755 3071 10771 3105
rect 10805 3071 10821 3105
rect 10755 3037 10821 3071
rect 10755 3003 10771 3037
rect 10805 3003 10821 3037
rect 10755 2969 10821 3003
rect 10755 2935 10771 2969
rect 10805 2935 10821 2969
rect 10755 2901 10821 2935
rect 10755 2867 10771 2901
rect 10805 2867 10821 2901
rect 10755 2833 10821 2867
rect 10755 2799 10771 2833
rect 10805 2799 10821 2833
rect 10755 2765 10821 2799
rect 10755 2731 10771 2765
rect 10805 2731 10821 2765
rect 10755 2697 10821 2731
rect 10755 2663 10771 2697
rect 10805 2663 10821 2697
rect 10755 2629 10821 2663
rect 10755 2595 10771 2629
rect 10805 2595 10821 2629
rect 10755 2561 10821 2595
rect 10755 2527 10771 2561
rect 10805 2527 10821 2561
rect 10755 2493 10821 2527
rect 10755 2459 10771 2493
rect 10805 2459 10821 2493
rect 10755 2425 10821 2459
rect 10755 2391 10771 2425
rect 10805 2391 10821 2425
rect 10755 2357 10821 2391
rect 10755 2323 10771 2357
rect 10805 2323 10821 2357
rect 10755 2289 10821 2323
rect 10755 2255 10771 2289
rect 10805 2255 10821 2289
rect 10755 2221 10821 2255
rect 10755 2187 10771 2221
rect 10805 2187 10821 2221
rect 10755 2153 10821 2187
rect 10755 2119 10771 2153
rect 10805 2119 10821 2153
rect 10755 2085 10821 2119
rect 10755 2051 10771 2085
rect 10805 2051 10821 2085
rect 10755 2017 10821 2051
rect 10755 1983 10771 2017
rect 10805 1983 10821 2017
rect 10755 1949 10821 1983
rect 10755 1915 10771 1949
rect 10805 1915 10821 1949
rect 10755 1881 10821 1915
rect 10755 1847 10771 1881
rect 10805 1847 10821 1881
rect 10755 1813 10821 1847
rect 10755 1779 10771 1813
rect 10805 1779 10821 1813
rect 10755 1745 10821 1779
rect 10755 1711 10771 1745
rect 10805 1711 10821 1745
rect 10755 1677 10821 1711
rect 10755 1643 10771 1677
rect 10805 1643 10821 1677
rect 10755 1609 10821 1643
rect 10755 1575 10771 1609
rect 10805 1575 10821 1609
rect 10755 1541 10821 1575
rect 10755 1507 10771 1541
rect 10805 1507 10821 1541
rect 10755 1473 10821 1507
rect 10755 1439 10771 1473
rect 10805 1439 10821 1473
rect 10755 1405 10821 1439
rect 10755 1371 10771 1405
rect 10805 1371 10821 1405
rect 10755 1337 10821 1371
rect 10755 1303 10771 1337
rect 10805 1303 10821 1337
rect 10755 1269 10821 1303
rect 10755 1235 10771 1269
rect 10805 1235 10821 1269
rect 10755 1201 10821 1235
rect 10755 1167 10771 1201
rect 10805 1167 10821 1201
rect 10755 1133 10821 1167
rect 10755 1099 10771 1133
rect 10805 1099 10821 1133
rect 10755 1065 10821 1099
rect 10755 1031 10771 1065
rect 10805 1031 10821 1065
rect 10755 997 10821 1031
rect 10755 963 10771 997
rect 10805 963 10821 997
rect 10755 929 10821 963
rect 10755 895 10771 929
rect 10805 895 10821 929
rect 10755 861 10821 895
rect 10755 827 10771 861
rect 10805 827 10821 861
rect 10755 793 10821 827
rect 10755 759 10771 793
rect 10805 759 10821 793
rect 10755 725 10821 759
rect 10755 691 10771 725
rect 10805 691 10821 725
rect 10755 657 10821 691
rect 10755 623 10771 657
rect 10805 623 10821 657
rect 10755 589 10821 623
rect 10755 555 10771 589
rect 10805 555 10821 589
rect 10755 521 10821 555
rect 10755 487 10771 521
rect 10805 487 10821 521
rect 10755 453 10821 487
rect 10755 419 10771 453
rect 10805 419 10821 453
rect 10755 385 10821 419
rect 10755 351 10771 385
rect 10805 351 10821 385
rect 10755 317 10821 351
rect 10755 283 10771 317
rect 10805 283 10821 317
rect 10755 249 10821 283
rect 10755 215 10771 249
rect 10805 215 10821 249
rect 10755 181 10821 215
rect 10755 147 10771 181
rect 10805 147 10821 181
rect 10755 113 10821 147
rect 10755 79 10771 113
rect 10805 79 10821 113
rect 10755 45 10821 79
rect 10755 11 10771 45
rect 10805 11 10821 45
rect 10755 -23 10821 11
rect 10755 -57 10771 -23
rect 10805 -57 10821 -23
rect 10755 -91 10821 -57
rect 10755 -125 10771 -91
rect 10805 -125 10821 -91
rect 10755 -159 10821 -125
rect 10755 -193 10771 -159
rect 10805 -193 10821 -159
rect 10755 -227 10821 -193
rect 10755 -261 10771 -227
rect 10805 -261 10821 -227
rect 10755 -295 10821 -261
rect 10755 -329 10771 -295
rect 10805 -329 10821 -295
rect 10755 -363 10821 -329
rect 10755 -397 10771 -363
rect 10805 -397 10821 -363
rect 10755 -431 10821 -397
rect 10755 -465 10771 -431
rect 10805 -465 10821 -431
rect 10755 -499 10821 -465
rect 10755 -533 10771 -499
rect 10805 -533 10821 -499
rect 10755 -567 10821 -533
rect 10755 -601 10771 -567
rect 10805 -601 10821 -567
rect 10755 -635 10821 -601
rect 10755 -669 10771 -635
rect 10805 -669 10821 -635
rect 10755 -703 10821 -669
rect 10755 -737 10771 -703
rect 10805 -737 10821 -703
rect 10755 -771 10821 -737
rect 10755 -805 10771 -771
rect 10805 -805 10821 -771
rect 10755 -839 10821 -805
rect 10755 -873 10771 -839
rect 10805 -873 10821 -839
rect 10755 -907 10821 -873
rect 10755 -941 10771 -907
rect 10805 -941 10821 -907
rect 10755 -975 10821 -941
rect 10755 -1009 10771 -975
rect 10805 -1009 10821 -975
rect 10755 -1043 10821 -1009
rect 10755 -1077 10771 -1043
rect 10805 -1077 10821 -1043
rect 10755 -1111 10821 -1077
rect 10755 -1145 10771 -1111
rect 10805 -1145 10821 -1111
rect 10755 -1179 10821 -1145
rect 10755 -1213 10771 -1179
rect 10805 -1213 10821 -1179
rect 10755 -1247 10821 -1213
rect 10755 -1281 10771 -1247
rect 10805 -1281 10821 -1247
rect 10755 -1315 10821 -1281
rect 10755 -1349 10771 -1315
rect 10805 -1349 10821 -1315
rect 10755 -1383 10821 -1349
rect 10755 -1417 10771 -1383
rect 10805 -1417 10821 -1383
rect 10755 -1451 10821 -1417
rect 10755 -1485 10771 -1451
rect 10805 -1485 10821 -1451
rect 10755 -1519 10821 -1485
rect 10755 -1553 10771 -1519
rect 10805 -1553 10821 -1519
rect 10755 -1587 10821 -1553
rect 10755 -1621 10771 -1587
rect 10805 -1621 10821 -1587
rect 10755 -1655 10821 -1621
rect 10755 -1689 10771 -1655
rect 10805 -1689 10821 -1655
rect 10755 -1723 10821 -1689
rect 10755 -1757 10771 -1723
rect 10805 -1757 10821 -1723
rect 10755 -1791 10821 -1757
rect 10755 -1825 10771 -1791
rect 10805 -1825 10821 -1791
rect 10755 -1859 10821 -1825
rect 10755 -1893 10771 -1859
rect 10805 -1893 10821 -1859
rect 10755 -1927 10821 -1893
rect 10755 -1961 10771 -1927
rect 10805 -1961 10821 -1927
rect 10755 -1995 10821 -1961
rect 10755 -2029 10771 -1995
rect 10805 -2029 10821 -1995
rect 10755 -2063 10821 -2029
rect 10755 -2097 10771 -2063
rect 10805 -2097 10821 -2063
rect 10755 -2131 10821 -2097
rect 10755 -2165 10771 -2131
rect 10805 -2165 10821 -2131
rect 10755 -2199 10821 -2165
rect 10755 -2233 10771 -2199
rect 10805 -2233 10821 -2199
rect 10755 -2267 10821 -2233
rect 10755 -2301 10771 -2267
rect 10805 -2301 10821 -2267
rect 10755 -2335 10821 -2301
rect 10755 -2369 10771 -2335
rect 10805 -2369 10821 -2335
rect 10755 -2403 10821 -2369
rect 10755 -2437 10771 -2403
rect 10805 -2437 10821 -2403
rect 10755 -2471 10821 -2437
rect 10755 -2505 10771 -2471
rect 10805 -2505 10821 -2471
rect 10755 -2539 10821 -2505
rect 10755 -2573 10771 -2539
rect 10805 -2573 10821 -2539
rect 10755 -2607 10821 -2573
rect 10755 -2641 10771 -2607
rect 10805 -2641 10821 -2607
rect 10755 -2675 10821 -2641
rect 10755 -2709 10771 -2675
rect 10805 -2709 10821 -2675
rect 10755 -2743 10821 -2709
rect 10755 -2777 10771 -2743
rect 10805 -2777 10821 -2743
rect 10755 -2811 10821 -2777
rect 10755 -2845 10771 -2811
rect 10805 -2845 10821 -2811
rect 10755 -2879 10821 -2845
rect 10755 -2913 10771 -2879
rect 10805 -2913 10821 -2879
rect 10755 -2947 10821 -2913
rect 10755 -2981 10771 -2947
rect 10805 -2981 10821 -2947
rect 10755 -3015 10821 -2981
rect 10755 -3049 10771 -3015
rect 10805 -3049 10821 -3015
rect 10755 -3083 10821 -3049
rect 10755 -3117 10771 -3083
rect 10805 -3117 10821 -3083
rect 10755 -3151 10821 -3117
rect 10755 -3185 10771 -3151
rect 10805 -3185 10821 -3151
rect 10755 -3219 10821 -3185
rect 10755 -3253 10771 -3219
rect 10805 -3253 10821 -3219
rect 10755 -3287 10821 -3253
rect 10755 -3321 10771 -3287
rect 10805 -3321 10821 -3287
rect 10755 -3355 10821 -3321
rect 10755 -3389 10771 -3355
rect 10805 -3389 10821 -3355
rect 10755 -3424 10821 -3389
rect 10755 -3458 10771 -3424
rect 10805 -3458 10821 -3424
rect 10755 -3493 10821 -3458
rect 10755 -3527 10771 -3493
rect 10805 -3527 10821 -3493
rect 10755 -3562 10821 -3527
rect 10755 -3596 10771 -3562
rect 10805 -3596 10821 -3562
rect 10755 -3631 10821 -3596
rect 10755 -3665 10771 -3631
rect 10805 -3665 10821 -3631
rect 10755 -3700 10821 -3665
rect 10755 -3734 10771 -3700
rect 10805 -3734 10821 -3700
rect 10755 -3769 10821 -3734
rect 10755 -3803 10771 -3769
rect 10805 -3803 10821 -3769
rect 10755 -3838 10821 -3803
rect 10755 -3872 10771 -3838
rect 10805 -3872 10821 -3838
rect 10755 -3907 10821 -3872
rect 8959 -3945 9363 -3929
rect 8959 -3961 9015 -3945
rect 8909 -3979 9015 -3961
rect 9049 -3979 9085 -3945
rect 9119 -3979 9155 -3945
rect 9189 -3979 9225 -3945
rect 9259 -3979 9295 -3945
rect 9329 -3979 9363 -3945
rect 8909 -3995 9363 -3979
rect 9297 -4033 9363 -3995
rect 9297 -4067 9313 -4033
rect 9347 -4067 9363 -4033
rect 9297 -4102 9363 -4067
rect 9297 -4136 9313 -4102
rect 9347 -4136 9363 -4102
rect 9297 -4171 9363 -4136
rect 9297 -4205 9313 -4171
rect 9347 -4205 9363 -4171
rect 9297 -4240 9363 -4205
rect 9297 -4274 9313 -4240
rect 9347 -4274 9363 -4240
rect 9297 -4309 9363 -4274
rect 9297 -4343 9313 -4309
rect 9347 -4343 9363 -4309
rect 9297 -4378 9363 -4343
rect 9297 -4412 9313 -4378
rect 9347 -4412 9363 -4378
rect 9297 -4447 9363 -4412
rect 9297 -4481 9313 -4447
rect 9347 -4481 9363 -4447
rect 9297 -4516 9363 -4481
rect 9297 -4550 9313 -4516
rect 9347 -4550 9363 -4516
rect 9297 -4585 9363 -4550
rect 9297 -4619 9313 -4585
rect 9347 -4619 9363 -4585
rect 9297 -4654 9363 -4619
rect 9297 -4688 9313 -4654
rect 9347 -4688 9363 -4654
rect 9297 -4723 9363 -4688
rect 9297 -4757 9313 -4723
rect 9347 -4757 9363 -4723
rect 9297 -4792 9363 -4757
rect 9297 -4826 9313 -4792
rect 9347 -4826 9363 -4792
rect 9297 -4861 9363 -4826
rect 9297 -4895 9313 -4861
rect 9347 -4895 9363 -4861
rect 9297 -4930 9363 -4895
rect 9297 -4964 9313 -4930
rect 9347 -4964 9363 -4930
rect 9297 -4999 9363 -4964
rect 9297 -5033 9313 -4999
rect 9347 -5033 9363 -4999
rect 9297 -5068 9363 -5033
rect 9297 -5102 9313 -5068
rect 9347 -5102 9363 -5068
rect 9297 -5137 9363 -5102
rect 9297 -5171 9313 -5137
rect 9347 -5171 9363 -5137
rect 9297 -5206 9363 -5171
rect 9297 -5240 9313 -5206
rect 9347 -5240 9363 -5206
rect 9297 -5275 9363 -5240
rect 9297 -5309 9313 -5275
rect 9347 -5309 9363 -5275
rect 9297 -5344 9363 -5309
rect 9297 -5378 9313 -5344
rect 9347 -5378 9363 -5344
rect 9297 -5413 9363 -5378
rect 9297 -5447 9313 -5413
rect 9347 -5447 9363 -5413
rect 9297 -5482 9363 -5447
rect 9297 -5516 9313 -5482
rect 9347 -5516 9363 -5482
rect 9297 -5551 9363 -5516
rect 9297 -5585 9313 -5551
rect 9347 -5585 9363 -5551
rect 9297 -5620 9363 -5585
rect 9297 -5654 9313 -5620
rect 9347 -5654 9363 -5620
rect 9297 -5689 9363 -5654
rect 9297 -5723 9313 -5689
rect 9347 -5723 9363 -5689
rect 9297 -5759 9363 -5723
rect 9297 -5793 9313 -5759
rect 9347 -5793 9363 -5759
rect 9297 -5829 9363 -5793
rect 9297 -5863 9313 -5829
rect 9347 -5863 9363 -5829
rect 9297 -5899 9363 -5863
rect 9297 -5933 9313 -5899
rect 9347 -5933 9363 -5899
rect 9297 -5969 9363 -5933
rect 9297 -6003 9313 -5969
rect 9347 -6003 9363 -5969
rect 9297 -6039 9363 -6003
rect 9297 -6073 9313 -6039
rect 9347 -6073 9363 -6039
rect 9297 -6109 9363 -6073
rect 9297 -6143 9313 -6109
rect 9347 -6111 9363 -6109
rect 10755 -3941 10771 -3907
rect 10805 -3941 10821 -3907
rect 10755 -3976 10821 -3941
rect 10755 -4010 10771 -3976
rect 10805 -4010 10821 -3976
rect 10755 -4045 10821 -4010
rect 10755 -4079 10771 -4045
rect 10805 -4079 10821 -4045
rect 10755 -4114 10821 -4079
rect 10755 -4148 10771 -4114
rect 10805 -4148 10821 -4114
rect 10755 -4183 10821 -4148
rect 10755 -4217 10771 -4183
rect 10805 -4217 10821 -4183
rect 10755 -4252 10821 -4217
rect 10755 -4286 10771 -4252
rect 10805 -4286 10821 -4252
rect 10755 -4321 10821 -4286
rect 10755 -4355 10771 -4321
rect 10805 -4355 10821 -4321
rect 10755 -4390 10821 -4355
rect 10755 -4424 10771 -4390
rect 10805 -4424 10821 -4390
rect 10755 -4459 10821 -4424
rect 10755 -4493 10771 -4459
rect 10805 -4493 10821 -4459
rect 10755 -4528 10821 -4493
rect 10755 -4562 10771 -4528
rect 10805 -4562 10821 -4528
rect 10755 -4597 10821 -4562
rect 10755 -4631 10771 -4597
rect 10805 -4631 10821 -4597
rect 10755 -4666 10821 -4631
rect 10755 -4700 10771 -4666
rect 10805 -4700 10821 -4666
rect 10755 -4735 10821 -4700
rect 10755 -4769 10771 -4735
rect 10805 -4769 10821 -4735
rect 10755 -4804 10821 -4769
rect 10755 -4838 10771 -4804
rect 10805 -4838 10821 -4804
rect 10755 -4873 10821 -4838
rect 10755 -4907 10771 -4873
rect 10805 -4907 10821 -4873
rect 10755 -4942 10821 -4907
rect 10755 -4976 10771 -4942
rect 10805 -4976 10821 -4942
rect 10755 -5011 10821 -4976
rect 10755 -5045 10771 -5011
rect 10805 -5045 10821 -5011
rect 10755 -5080 10821 -5045
rect 10755 -5114 10771 -5080
rect 10805 -5114 10821 -5080
rect 10755 -5149 10821 -5114
rect 10755 -5183 10771 -5149
rect 10805 -5183 10821 -5149
rect 10755 -5218 10821 -5183
rect 10755 -5252 10771 -5218
rect 10805 -5252 10821 -5218
rect 10755 -5287 10821 -5252
rect 10755 -5321 10771 -5287
rect 10805 -5321 10821 -5287
rect 10755 -5356 10821 -5321
rect 10755 -5390 10771 -5356
rect 10805 -5390 10821 -5356
rect 10755 -5425 10821 -5390
rect 10755 -5459 10771 -5425
rect 10805 -5459 10821 -5425
rect 10755 -5494 10821 -5459
rect 10755 -5528 10771 -5494
rect 10805 -5528 10821 -5494
rect 10755 -5563 10821 -5528
rect 10755 -5597 10771 -5563
rect 10805 -5597 10821 -5563
rect 10755 -5632 10821 -5597
rect 10755 -5666 10771 -5632
rect 10805 -5666 10821 -5632
rect 10755 -5701 10821 -5666
rect 10755 -5735 10771 -5701
rect 10805 -5735 10821 -5701
rect 10755 -5770 10821 -5735
rect 10755 -5804 10771 -5770
rect 10805 -5804 10821 -5770
rect 10755 -5839 10821 -5804
rect 10755 -5873 10771 -5839
rect 10805 -5873 10821 -5839
rect 10755 -5908 10821 -5873
rect 10755 -5942 10771 -5908
rect 10805 -5942 10821 -5908
rect 10755 -5977 10821 -5942
rect 10755 -6011 10771 -5977
rect 10805 -6011 10821 -5977
rect 10755 -6046 10821 -6011
rect 10755 -6080 10771 -6046
rect 10805 -6080 10821 -6046
rect 9347 -6127 9521 -6111
rect 9347 -6143 9453 -6127
rect 9297 -6161 9453 -6143
rect 9487 -6161 9521 -6127
rect 9297 -6177 9521 -6161
rect 9455 -6238 9521 -6177
rect 9455 -6272 9471 -6238
rect 9505 -6272 9521 -6238
rect 9455 -6324 9521 -6272
rect 10755 -6115 10821 -6080
rect 10755 -6149 10771 -6115
rect 10805 -6149 10821 -6115
rect 10755 -6184 10821 -6149
rect 10755 -6218 10771 -6184
rect 10805 -6218 10821 -6184
rect 10755 -6253 10821 -6218
rect 10755 -6287 10771 -6253
rect 10805 -6287 10821 -6253
rect 10755 -6322 10821 -6287
rect 10755 -6324 10771 -6322
rect 9455 -6340 10771 -6324
rect 9455 -6374 9489 -6340
rect 9523 -6374 9560 -6340
rect 9594 -6374 9631 -6340
rect 9665 -6374 9701 -6340
rect 9735 -6374 9771 -6340
rect 9805 -6374 9841 -6340
rect 9875 -6374 9911 -6340
rect 9945 -6374 9981 -6340
rect 10015 -6374 10051 -6340
rect 10085 -6374 10121 -6340
rect 10155 -6374 10191 -6340
rect 10225 -6374 10261 -6340
rect 10295 -6374 10331 -6340
rect 10365 -6374 10401 -6340
rect 10435 -6374 10471 -6340
rect 10505 -6374 10541 -6340
rect 10575 -6374 10611 -6340
rect 10645 -6374 10681 -6340
rect 10715 -6356 10771 -6340
rect 10805 -6356 10821 -6322
rect 10715 -6374 10821 -6356
rect 9455 -6390 10821 -6374
<< polycont >>
rect 8925 22179 8959 22213
rect 9005 22195 9039 22229
rect 9075 22195 9109 22229
rect 9145 22195 9179 22229
rect 9215 22195 9249 22229
rect 9285 22195 9319 22229
rect 9355 22195 9389 22229
rect 9425 22195 9459 22229
rect 9495 22195 9529 22229
rect 9565 22195 9599 22229
rect 9635 22195 9669 22229
rect 9705 22195 9739 22229
rect 9775 22195 9809 22229
rect 9845 22195 9879 22229
rect 9915 22195 9949 22229
rect 9985 22195 10019 22229
rect 10056 22195 10090 22229
rect 10127 22195 10161 22229
rect 10198 22195 10232 22229
rect 10269 22195 10303 22229
rect 10340 22195 10374 22229
rect 10411 22195 10445 22229
rect 10482 22195 10516 22229
rect 10553 22195 10587 22229
rect 10624 22195 10658 22229
rect 10695 22195 10729 22229
rect 10771 22179 10805 22213
rect 8925 22111 8959 22145
rect 8925 22043 8959 22077
rect 8925 21975 8959 22009
rect 8925 21907 8959 21941
rect 8925 21839 8959 21873
rect 8925 21771 8959 21805
rect 8925 21703 8959 21737
rect 8925 21635 8959 21669
rect 8925 21567 8959 21601
rect 8925 21499 8959 21533
rect 8925 21431 8959 21465
rect 8925 21363 8959 21397
rect 8925 21295 8959 21329
rect 8925 21227 8959 21261
rect 8925 21159 8959 21193
rect 8925 21091 8959 21125
rect 8925 21023 8959 21057
rect 8925 20955 8959 20989
rect 8925 20887 8959 20921
rect 8925 20819 8959 20853
rect 8925 20751 8959 20785
rect 8925 20683 8959 20717
rect 8925 20615 8959 20649
rect 8925 20547 8959 20581
rect 8925 20479 8959 20513
rect 8925 20411 8959 20445
rect 8925 20343 8959 20377
rect 8925 20275 8959 20309
rect 8925 20207 8959 20241
rect 8925 20139 8959 20173
rect 8925 20071 8959 20105
rect 8925 20003 8959 20037
rect 8925 19935 8959 19969
rect 8925 19867 8959 19901
rect 8925 19799 8959 19833
rect 8925 19731 8959 19765
rect 8925 19663 8959 19697
rect 8925 19595 8959 19629
rect 8925 19527 8959 19561
rect 8925 19459 8959 19493
rect 8925 19391 8959 19425
rect 8925 19323 8959 19357
rect 8925 19255 8959 19289
rect 8925 19187 8959 19221
rect 8925 19119 8959 19153
rect 8925 19051 8959 19085
rect 8925 18983 8959 19017
rect 8925 18915 8959 18949
rect 8925 18847 8959 18881
rect 8925 18779 8959 18813
rect 8925 18711 8959 18745
rect 8925 18643 8959 18677
rect 8925 18575 8959 18609
rect 8925 18507 8959 18541
rect 8925 18439 8959 18473
rect 8925 18371 8959 18405
rect 8925 18303 8959 18337
rect 8925 18235 8959 18269
rect 8925 18167 8959 18201
rect 8925 18099 8959 18133
rect 8925 18031 8959 18065
rect 8925 17963 8959 17997
rect 8925 17895 8959 17929
rect 8925 17827 8959 17861
rect 8925 17759 8959 17793
rect 8925 17691 8959 17725
rect 8925 17623 8959 17657
rect 8925 17555 8959 17589
rect 8925 17487 8959 17521
rect 8925 17419 8959 17453
rect 8925 17351 8959 17385
rect 8925 17283 8959 17317
rect 8925 17215 8959 17249
rect 8925 17147 8959 17181
rect 8925 17079 8959 17113
rect 8925 17011 8959 17045
rect 8925 16943 8959 16977
rect 8925 16875 8959 16909
rect 8925 16807 8959 16841
rect 8925 16739 8959 16773
rect 8925 16671 8959 16705
rect 8925 16603 8959 16637
rect 8925 16535 8959 16569
rect 8925 16467 8959 16501
rect 8925 16399 8959 16433
rect 8925 16331 8959 16365
rect 8925 16263 8959 16297
rect 8925 16195 8959 16229
rect 8925 16127 8959 16161
rect 8925 16059 8959 16093
rect 8925 15991 8959 16025
rect 8925 15923 8959 15957
rect 8925 15855 8959 15889
rect 8925 15787 8959 15821
rect 8925 15719 8959 15753
rect 8925 15651 8959 15685
rect 8925 15583 8959 15617
rect 8925 15515 8959 15549
rect 8925 15447 8959 15481
rect 8925 15379 8959 15413
rect 8925 15311 8959 15345
rect 8925 15243 8959 15277
rect 8925 15175 8959 15209
rect 8925 15107 8959 15141
rect 8925 15039 8959 15073
rect 8925 14971 8959 15005
rect 8925 14903 8959 14937
rect 8925 14835 8959 14869
rect 8925 14767 8959 14801
rect 8925 14699 8959 14733
rect 8925 14631 8959 14665
rect 8925 14563 8959 14597
rect 8925 14495 8959 14529
rect 8925 14427 8959 14461
rect 8925 14359 8959 14393
rect 8925 14291 8959 14325
rect 8925 14223 8959 14257
rect 8925 14155 8959 14189
rect 8925 14087 8959 14121
rect 8925 14019 8959 14053
rect 8925 13951 8959 13985
rect 8925 13883 8959 13917
rect 8925 13815 8959 13849
rect 8925 13747 8959 13781
rect 8925 13679 8959 13713
rect 8925 13611 8959 13645
rect 8925 13543 8959 13577
rect 8925 13475 8959 13509
rect 8925 13407 8959 13441
rect 8925 13339 8959 13373
rect 8925 13271 8959 13305
rect 8925 13203 8959 13237
rect 8925 13135 8959 13169
rect 8925 13067 8959 13101
rect 8925 12999 8959 13033
rect 8925 12931 8959 12965
rect 8925 12863 8959 12897
rect 8925 12795 8959 12829
rect 8925 12727 8959 12761
rect 8925 12659 8959 12693
rect 8925 12591 8959 12625
rect 8925 12523 8959 12557
rect 8925 12455 8959 12489
rect 8925 12387 8959 12421
rect 8925 12319 8959 12353
rect 8925 12251 8959 12285
rect 8925 12183 8959 12217
rect 8925 12115 8959 12149
rect 8925 12047 8959 12081
rect 8925 11979 8959 12013
rect 8925 11911 8959 11945
rect 8925 11843 8959 11877
rect 8925 11775 8959 11809
rect 8925 11707 8959 11741
rect 8925 11639 8959 11673
rect 8925 11571 8959 11605
rect 8925 11503 8959 11537
rect 8925 11435 8959 11469
rect 8925 11367 8959 11401
rect 8925 11299 8959 11333
rect 8925 11231 8959 11265
rect 8925 11163 8959 11197
rect 8925 11095 8959 11129
rect 8925 11027 8959 11061
rect 8925 10959 8959 10993
rect 8925 10891 8959 10925
rect 8925 10823 8959 10857
rect 8925 10755 8959 10789
rect 8925 10687 8959 10721
rect 8925 10619 8959 10653
rect 8925 10551 8959 10585
rect 8925 10483 8959 10517
rect 8925 10415 8959 10449
rect 8925 10347 8959 10381
rect 8925 10279 8959 10313
rect 8925 10211 8959 10245
rect 8925 10143 8959 10177
rect 8925 10075 8959 10109
rect 8925 10007 8959 10041
rect 8925 9939 8959 9973
rect 8925 9871 8959 9905
rect 8925 9803 8959 9837
rect 8925 9735 8959 9769
rect 8925 9667 8959 9701
rect 8925 9599 8959 9633
rect 8925 9531 8959 9565
rect 8925 9463 8959 9497
rect 8925 9395 8959 9429
rect 8925 9327 8959 9361
rect 8925 9259 8959 9293
rect 8925 9191 8959 9225
rect 8925 9123 8959 9157
rect 8925 9055 8959 9089
rect 8925 8987 8959 9021
rect 8925 8919 8959 8953
rect 8925 8851 8959 8885
rect 8925 8783 8959 8817
rect 8925 8715 8959 8749
rect 8925 8647 8959 8681
rect 8925 8579 8959 8613
rect 8925 8511 8959 8545
rect 8925 8443 8959 8477
rect 8925 8375 8959 8409
rect 8925 8307 8959 8341
rect 8925 8239 8959 8273
rect 8925 8171 8959 8205
rect 8925 8103 8959 8137
rect 8925 8035 8959 8069
rect 8925 7967 8959 8001
rect 8925 7899 8959 7933
rect 8925 7831 8959 7865
rect 8925 7763 8959 7797
rect 8925 7695 8959 7729
rect 8925 7627 8959 7661
rect 8925 7559 8959 7593
rect 8925 7491 8959 7525
rect 8925 7423 8959 7457
rect 8925 7355 8959 7389
rect 8925 7287 8959 7321
rect 8925 7219 8959 7253
rect 8925 7151 8959 7185
rect 8925 7083 8959 7117
rect 8925 7015 8959 7049
rect 8925 6947 8959 6981
rect 8925 6879 8959 6913
rect 8925 6811 8959 6845
rect 8925 6743 8959 6777
rect 8925 6675 8959 6709
rect 8925 6607 8959 6641
rect 8925 6539 8959 6573
rect 8925 6471 8959 6505
rect 8925 6403 8959 6437
rect 8925 6335 8959 6369
rect 8925 6267 8959 6301
rect 8925 6199 8959 6233
rect 8925 6131 8959 6165
rect 8925 6063 8959 6097
rect 8925 5995 8959 6029
rect 8925 5927 8959 5961
rect 8925 5859 8959 5893
rect 8925 5791 8959 5825
rect 8925 5723 8959 5757
rect 8925 5655 8959 5689
rect 8925 5587 8959 5621
rect 8925 5519 8959 5553
rect 8925 5451 8959 5485
rect 8925 5383 8959 5417
rect 8925 5315 8959 5349
rect 8925 5247 8959 5281
rect 8925 5179 8959 5213
rect 8925 5111 8959 5145
rect 8925 5043 8959 5077
rect 8925 4975 8959 5009
rect 8925 4907 8959 4941
rect 8925 4839 8959 4873
rect 8925 4771 8959 4805
rect 8925 4703 8959 4737
rect 8925 4635 8959 4669
rect 8925 4567 8959 4601
rect 8925 4499 8959 4533
rect 8925 4431 8959 4465
rect 8925 4363 8959 4397
rect 8925 4295 8959 4329
rect 8925 4227 8959 4261
rect 8925 4159 8959 4193
rect 8925 4091 8959 4125
rect 8925 4023 8959 4057
rect 8925 3955 8959 3989
rect 8925 3887 8959 3921
rect 8925 3819 8959 3853
rect 8925 3751 8959 3785
rect 8925 3683 8959 3717
rect 8925 3615 8959 3649
rect 8925 3547 8959 3581
rect 8925 3479 8959 3513
rect 8925 3411 8959 3445
rect 8925 3343 8959 3377
rect 8925 3275 8959 3309
rect 8925 3207 8959 3241
rect 8925 3139 8959 3173
rect 8925 3071 8959 3105
rect 8925 3003 8959 3037
rect 8925 2935 8959 2969
rect 8925 2867 8959 2901
rect 8925 2799 8959 2833
rect 8925 2731 8959 2765
rect 8925 2663 8959 2697
rect 8925 2595 8959 2629
rect 8925 2527 8959 2561
rect 8925 2459 8959 2493
rect 8925 2391 8959 2425
rect 8925 2323 8959 2357
rect 8925 2255 8959 2289
rect 8925 2187 8959 2221
rect 8925 2119 8959 2153
rect 2326 1603 2360 1637
rect 2402 1603 2436 1637
rect 2524 1603 2558 1637
rect 2658 1603 2692 1637
rect 2780 1603 2814 1637
rect 2914 1603 2948 1637
rect 3036 1603 3070 1637
rect 3170 1603 3204 1637
rect 3292 1603 3326 1637
rect 3426 1603 3460 1637
rect 3548 1603 3582 1637
rect 3624 1603 3658 1637
rect 8925 2051 8959 2085
rect 8925 1983 8959 2017
rect 8925 1915 8959 1949
rect 8925 1847 8959 1881
rect 8925 1779 8959 1813
rect 8925 1711 8959 1745
rect 8925 1643 8959 1677
rect 8925 1575 8959 1609
rect 8925 1507 8959 1541
rect 8925 1439 8959 1473
rect 8925 1371 8959 1405
rect 8050 1219 8084 1253
rect 8126 1219 8160 1253
rect 8925 1303 8959 1337
rect 8925 1235 8959 1269
rect 8925 1167 8959 1201
rect 8925 1099 8959 1133
rect 8925 1031 8959 1065
rect 8925 963 8959 997
rect 8925 895 8959 929
rect 8925 827 8959 861
rect 8925 759 8959 793
rect 8925 691 8959 725
rect 8925 623 8959 657
rect 8925 555 8959 589
rect 8925 487 8959 521
rect 8925 419 8959 453
rect 8925 351 8959 385
rect 8925 283 8959 317
rect 8925 215 8959 249
rect 8925 147 8959 181
rect 8925 79 8959 113
rect 8925 11 8959 45
rect 8925 -57 8959 -23
rect 8925 -125 8959 -91
rect 8925 -193 8959 -159
rect 8925 -261 8959 -227
rect 8925 -329 8959 -295
rect 8925 -397 8959 -363
rect 8925 -465 8959 -431
rect 8925 -533 8959 -499
rect 8925 -601 8959 -567
rect 8925 -669 8959 -635
rect 8925 -737 8959 -703
rect 8925 -805 8959 -771
rect 8925 -873 8959 -839
rect 8925 -941 8959 -907
rect 8925 -1009 8959 -975
rect 8925 -1077 8959 -1043
rect 8925 -1145 8959 -1111
rect 8925 -1213 8959 -1179
rect 8925 -1281 8959 -1247
rect 8925 -1349 8959 -1315
rect 8925 -1417 8959 -1383
rect 8925 -1485 8959 -1451
rect 8925 -1553 8959 -1519
rect 8925 -1621 8959 -1587
rect 8925 -1689 8959 -1655
rect 8925 -1757 8959 -1723
rect 8925 -1825 8959 -1791
rect 8925 -1893 8959 -1859
rect 8925 -1961 8959 -1927
rect 8925 -2029 8959 -1995
rect 8925 -2098 8959 -2064
rect 8925 -2167 8959 -2133
rect 8925 -2236 8959 -2202
rect 8925 -2305 8959 -2271
rect 8925 -2374 8959 -2340
rect 8925 -2443 8959 -2409
rect 8925 -2512 8959 -2478
rect 8925 -2581 8959 -2547
rect 8925 -2650 8959 -2616
rect 8925 -2719 8959 -2685
rect 8925 -2788 8959 -2754
rect 8925 -2857 8959 -2823
rect 8925 -2926 8959 -2892
rect 8925 -2995 8959 -2961
rect 8925 -3064 8959 -3030
rect 8925 -3133 8959 -3099
rect 8925 -3202 8959 -3168
rect 8925 -3271 8959 -3237
rect 8925 -3340 8959 -3306
rect 8925 -3409 8959 -3375
rect 8925 -3478 8959 -3444
rect 8925 -3547 8959 -3513
rect 8925 -3616 8959 -3582
rect 8925 -3685 8959 -3651
rect 8925 -3754 8959 -3720
rect 8925 -3823 8959 -3789
rect 8925 -3892 8959 -3858
rect 8925 -3961 8959 -3927
rect 10771 22111 10805 22145
rect 10771 22043 10805 22077
rect 10771 21975 10805 22009
rect 10771 21907 10805 21941
rect 10771 21839 10805 21873
rect 10771 21771 10805 21805
rect 10771 21703 10805 21737
rect 10771 21635 10805 21669
rect 10771 21567 10805 21601
rect 10771 21499 10805 21533
rect 10771 21431 10805 21465
rect 10771 21363 10805 21397
rect 10771 21295 10805 21329
rect 10771 21227 10805 21261
rect 10771 21159 10805 21193
rect 10771 21091 10805 21125
rect 10771 21023 10805 21057
rect 10771 20955 10805 20989
rect 10771 20887 10805 20921
rect 10771 20819 10805 20853
rect 10771 20751 10805 20785
rect 10771 20683 10805 20717
rect 10771 20615 10805 20649
rect 10771 20547 10805 20581
rect 10771 20479 10805 20513
rect 10771 20411 10805 20445
rect 10771 20343 10805 20377
rect 10771 20275 10805 20309
rect 10771 20207 10805 20241
rect 10771 20139 10805 20173
rect 10771 20071 10805 20105
rect 10771 20003 10805 20037
rect 10771 19935 10805 19969
rect 10771 19867 10805 19901
rect 10771 19799 10805 19833
rect 10771 19731 10805 19765
rect 10771 19663 10805 19697
rect 10771 19595 10805 19629
rect 10771 19527 10805 19561
rect 10771 19459 10805 19493
rect 10771 19391 10805 19425
rect 10771 19323 10805 19357
rect 10771 19255 10805 19289
rect 10771 19187 10805 19221
rect 10771 19119 10805 19153
rect 10771 19051 10805 19085
rect 10771 18983 10805 19017
rect 10771 18915 10805 18949
rect 10771 18847 10805 18881
rect 10771 18779 10805 18813
rect 10771 18711 10805 18745
rect 10771 18643 10805 18677
rect 10771 18575 10805 18609
rect 10771 18507 10805 18541
rect 10771 18439 10805 18473
rect 10771 18371 10805 18405
rect 10771 18303 10805 18337
rect 10771 18235 10805 18269
rect 10771 18167 10805 18201
rect 10771 18099 10805 18133
rect 10771 18031 10805 18065
rect 10771 17963 10805 17997
rect 10771 17895 10805 17929
rect 10771 17827 10805 17861
rect 10771 17759 10805 17793
rect 10771 17691 10805 17725
rect 10771 17623 10805 17657
rect 10771 17555 10805 17589
rect 10771 17487 10805 17521
rect 10771 17419 10805 17453
rect 10771 17351 10805 17385
rect 10771 17283 10805 17317
rect 10771 17215 10805 17249
rect 10771 17147 10805 17181
rect 10771 17079 10805 17113
rect 10771 17011 10805 17045
rect 10771 16943 10805 16977
rect 10771 16875 10805 16909
rect 10771 16807 10805 16841
rect 10771 16739 10805 16773
rect 10771 16671 10805 16705
rect 10771 16603 10805 16637
rect 10771 16535 10805 16569
rect 10771 16467 10805 16501
rect 10771 16399 10805 16433
rect 10771 16331 10805 16365
rect 10771 16263 10805 16297
rect 10771 16195 10805 16229
rect 10771 16127 10805 16161
rect 10771 16059 10805 16093
rect 10771 15991 10805 16025
rect 10771 15923 10805 15957
rect 10771 15855 10805 15889
rect 10771 15787 10805 15821
rect 10771 15719 10805 15753
rect 10771 15651 10805 15685
rect 10771 15583 10805 15617
rect 10771 15515 10805 15549
rect 10771 15447 10805 15481
rect 10771 15379 10805 15413
rect 10771 15311 10805 15345
rect 10771 15243 10805 15277
rect 10771 15175 10805 15209
rect 10771 15107 10805 15141
rect 10771 15039 10805 15073
rect 10771 14971 10805 15005
rect 10771 14903 10805 14937
rect 10771 14835 10805 14869
rect 10771 14767 10805 14801
rect 10771 14699 10805 14733
rect 10771 14631 10805 14665
rect 10771 14563 10805 14597
rect 10771 14495 10805 14529
rect 10771 14427 10805 14461
rect 10771 14359 10805 14393
rect 10771 14291 10805 14325
rect 10771 14223 10805 14257
rect 10771 14155 10805 14189
rect 10771 14087 10805 14121
rect 10771 14019 10805 14053
rect 10771 13951 10805 13985
rect 10771 13883 10805 13917
rect 10771 13815 10805 13849
rect 10771 13747 10805 13781
rect 10771 13679 10805 13713
rect 10771 13611 10805 13645
rect 10771 13543 10805 13577
rect 10771 13475 10805 13509
rect 10771 13407 10805 13441
rect 10771 13339 10805 13373
rect 10771 13271 10805 13305
rect 10771 13203 10805 13237
rect 10771 13135 10805 13169
rect 10771 13067 10805 13101
rect 10771 12999 10805 13033
rect 10771 12931 10805 12965
rect 10771 12863 10805 12897
rect 10771 12795 10805 12829
rect 10771 12727 10805 12761
rect 10771 12659 10805 12693
rect 10771 12591 10805 12625
rect 10771 12523 10805 12557
rect 10771 12455 10805 12489
rect 10771 12387 10805 12421
rect 10771 12319 10805 12353
rect 10771 12251 10805 12285
rect 10771 12183 10805 12217
rect 10771 12115 10805 12149
rect 10771 12047 10805 12081
rect 10771 11979 10805 12013
rect 10771 11911 10805 11945
rect 10771 11843 10805 11877
rect 10771 11775 10805 11809
rect 10771 11707 10805 11741
rect 10771 11639 10805 11673
rect 10771 11571 10805 11605
rect 10771 11503 10805 11537
rect 10771 11435 10805 11469
rect 10771 11367 10805 11401
rect 10771 11299 10805 11333
rect 10771 11231 10805 11265
rect 10771 11163 10805 11197
rect 10771 11095 10805 11129
rect 10771 11027 10805 11061
rect 10771 10959 10805 10993
rect 10771 10891 10805 10925
rect 10771 10823 10805 10857
rect 10771 10755 10805 10789
rect 10771 10687 10805 10721
rect 10771 10619 10805 10653
rect 10771 10551 10805 10585
rect 10771 10483 10805 10517
rect 10771 10415 10805 10449
rect 10771 10347 10805 10381
rect 10771 10279 10805 10313
rect 10771 10211 10805 10245
rect 10771 10143 10805 10177
rect 10771 10075 10805 10109
rect 10771 10007 10805 10041
rect 10771 9939 10805 9973
rect 10771 9871 10805 9905
rect 10771 9803 10805 9837
rect 10771 9735 10805 9769
rect 10771 9667 10805 9701
rect 10771 9599 10805 9633
rect 10771 9531 10805 9565
rect 10771 9463 10805 9497
rect 10771 9395 10805 9429
rect 10771 9327 10805 9361
rect 10771 9259 10805 9293
rect 10771 9191 10805 9225
rect 10771 9123 10805 9157
rect 10771 9055 10805 9089
rect 10771 8987 10805 9021
rect 10771 8919 10805 8953
rect 10771 8851 10805 8885
rect 10771 8783 10805 8817
rect 10771 8715 10805 8749
rect 10771 8647 10805 8681
rect 10771 8579 10805 8613
rect 10771 8511 10805 8545
rect 10771 8443 10805 8477
rect 10771 8375 10805 8409
rect 10771 8307 10805 8341
rect 10771 8239 10805 8273
rect 10771 8171 10805 8205
rect 10771 8103 10805 8137
rect 10771 8035 10805 8069
rect 10771 7967 10805 8001
rect 10771 7899 10805 7933
rect 10771 7831 10805 7865
rect 10771 7763 10805 7797
rect 10771 7695 10805 7729
rect 10771 7627 10805 7661
rect 10771 7559 10805 7593
rect 10771 7491 10805 7525
rect 10771 7423 10805 7457
rect 10771 7355 10805 7389
rect 10771 7287 10805 7321
rect 10771 7219 10805 7253
rect 10771 7151 10805 7185
rect 10771 7083 10805 7117
rect 10771 7015 10805 7049
rect 10771 6947 10805 6981
rect 10771 6879 10805 6913
rect 10771 6811 10805 6845
rect 10771 6743 10805 6777
rect 10771 6675 10805 6709
rect 10771 6607 10805 6641
rect 10771 6539 10805 6573
rect 10771 6471 10805 6505
rect 10771 6403 10805 6437
rect 10771 6335 10805 6369
rect 10771 6267 10805 6301
rect 10771 6199 10805 6233
rect 10771 6131 10805 6165
rect 10771 6063 10805 6097
rect 10771 5995 10805 6029
rect 10771 5927 10805 5961
rect 10771 5859 10805 5893
rect 10771 5791 10805 5825
rect 10771 5723 10805 5757
rect 10771 5655 10805 5689
rect 10771 5587 10805 5621
rect 10771 5519 10805 5553
rect 10771 5451 10805 5485
rect 10771 5383 10805 5417
rect 10771 5315 10805 5349
rect 10771 5247 10805 5281
rect 10771 5179 10805 5213
rect 10771 5111 10805 5145
rect 10771 5043 10805 5077
rect 10771 4975 10805 5009
rect 10771 4907 10805 4941
rect 10771 4839 10805 4873
rect 10771 4771 10805 4805
rect 10771 4703 10805 4737
rect 10771 4635 10805 4669
rect 10771 4567 10805 4601
rect 10771 4499 10805 4533
rect 10771 4431 10805 4465
rect 10771 4363 10805 4397
rect 10771 4295 10805 4329
rect 10771 4227 10805 4261
rect 10771 4159 10805 4193
rect 10771 4091 10805 4125
rect 10771 4023 10805 4057
rect 10771 3955 10805 3989
rect 10771 3887 10805 3921
rect 10771 3819 10805 3853
rect 10771 3751 10805 3785
rect 10771 3683 10805 3717
rect 10771 3615 10805 3649
rect 10771 3547 10805 3581
rect 10771 3479 10805 3513
rect 10771 3411 10805 3445
rect 10771 3343 10805 3377
rect 10771 3275 10805 3309
rect 10771 3207 10805 3241
rect 10771 3139 10805 3173
rect 10771 3071 10805 3105
rect 10771 3003 10805 3037
rect 10771 2935 10805 2969
rect 10771 2867 10805 2901
rect 10771 2799 10805 2833
rect 10771 2731 10805 2765
rect 10771 2663 10805 2697
rect 10771 2595 10805 2629
rect 10771 2527 10805 2561
rect 10771 2459 10805 2493
rect 10771 2391 10805 2425
rect 10771 2323 10805 2357
rect 10771 2255 10805 2289
rect 10771 2187 10805 2221
rect 10771 2119 10805 2153
rect 10771 2051 10805 2085
rect 10771 1983 10805 2017
rect 10771 1915 10805 1949
rect 10771 1847 10805 1881
rect 10771 1779 10805 1813
rect 10771 1711 10805 1745
rect 10771 1643 10805 1677
rect 10771 1575 10805 1609
rect 10771 1507 10805 1541
rect 10771 1439 10805 1473
rect 10771 1371 10805 1405
rect 10771 1303 10805 1337
rect 10771 1235 10805 1269
rect 10771 1167 10805 1201
rect 10771 1099 10805 1133
rect 10771 1031 10805 1065
rect 10771 963 10805 997
rect 10771 895 10805 929
rect 10771 827 10805 861
rect 10771 759 10805 793
rect 10771 691 10805 725
rect 10771 623 10805 657
rect 10771 555 10805 589
rect 10771 487 10805 521
rect 10771 419 10805 453
rect 10771 351 10805 385
rect 10771 283 10805 317
rect 10771 215 10805 249
rect 10771 147 10805 181
rect 10771 79 10805 113
rect 10771 11 10805 45
rect 10771 -57 10805 -23
rect 10771 -125 10805 -91
rect 10771 -193 10805 -159
rect 10771 -261 10805 -227
rect 10771 -329 10805 -295
rect 10771 -397 10805 -363
rect 10771 -465 10805 -431
rect 10771 -533 10805 -499
rect 10771 -601 10805 -567
rect 10771 -669 10805 -635
rect 10771 -737 10805 -703
rect 10771 -805 10805 -771
rect 10771 -873 10805 -839
rect 10771 -941 10805 -907
rect 10771 -1009 10805 -975
rect 10771 -1077 10805 -1043
rect 10771 -1145 10805 -1111
rect 10771 -1213 10805 -1179
rect 10771 -1281 10805 -1247
rect 10771 -1349 10805 -1315
rect 10771 -1417 10805 -1383
rect 10771 -1485 10805 -1451
rect 10771 -1553 10805 -1519
rect 10771 -1621 10805 -1587
rect 10771 -1689 10805 -1655
rect 10771 -1757 10805 -1723
rect 10771 -1825 10805 -1791
rect 10771 -1893 10805 -1859
rect 10771 -1961 10805 -1927
rect 10771 -2029 10805 -1995
rect 10771 -2097 10805 -2063
rect 10771 -2165 10805 -2131
rect 10771 -2233 10805 -2199
rect 10771 -2301 10805 -2267
rect 10771 -2369 10805 -2335
rect 10771 -2437 10805 -2403
rect 10771 -2505 10805 -2471
rect 10771 -2573 10805 -2539
rect 10771 -2641 10805 -2607
rect 10771 -2709 10805 -2675
rect 10771 -2777 10805 -2743
rect 10771 -2845 10805 -2811
rect 10771 -2913 10805 -2879
rect 10771 -2981 10805 -2947
rect 10771 -3049 10805 -3015
rect 10771 -3117 10805 -3083
rect 10771 -3185 10805 -3151
rect 10771 -3253 10805 -3219
rect 10771 -3321 10805 -3287
rect 10771 -3389 10805 -3355
rect 10771 -3458 10805 -3424
rect 10771 -3527 10805 -3493
rect 10771 -3596 10805 -3562
rect 10771 -3665 10805 -3631
rect 10771 -3734 10805 -3700
rect 10771 -3803 10805 -3769
rect 10771 -3872 10805 -3838
rect 9015 -3979 9049 -3945
rect 9085 -3979 9119 -3945
rect 9155 -3979 9189 -3945
rect 9225 -3979 9259 -3945
rect 9295 -3979 9329 -3945
rect 9313 -4067 9347 -4033
rect 9313 -4136 9347 -4102
rect 9313 -4205 9347 -4171
rect 9313 -4274 9347 -4240
rect 9313 -4343 9347 -4309
rect 9313 -4412 9347 -4378
rect 9313 -4481 9347 -4447
rect 9313 -4550 9347 -4516
rect 9313 -4619 9347 -4585
rect 9313 -4688 9347 -4654
rect 9313 -4757 9347 -4723
rect 9313 -4826 9347 -4792
rect 9313 -4895 9347 -4861
rect 9313 -4964 9347 -4930
rect 9313 -5033 9347 -4999
rect 9313 -5102 9347 -5068
rect 9313 -5171 9347 -5137
rect 9313 -5240 9347 -5206
rect 9313 -5309 9347 -5275
rect 9313 -5378 9347 -5344
rect 9313 -5447 9347 -5413
rect 9313 -5516 9347 -5482
rect 9313 -5585 9347 -5551
rect 9313 -5654 9347 -5620
rect 9313 -5723 9347 -5689
rect 9313 -5793 9347 -5759
rect 9313 -5863 9347 -5829
rect 9313 -5933 9347 -5899
rect 9313 -6003 9347 -5969
rect 9313 -6073 9347 -6039
rect 9313 -6143 9347 -6109
rect 10771 -3941 10805 -3907
rect 10771 -4010 10805 -3976
rect 10771 -4079 10805 -4045
rect 10771 -4148 10805 -4114
rect 10771 -4217 10805 -4183
rect 10771 -4286 10805 -4252
rect 10771 -4355 10805 -4321
rect 10771 -4424 10805 -4390
rect 10771 -4493 10805 -4459
rect 10771 -4562 10805 -4528
rect 10771 -4631 10805 -4597
rect 10771 -4700 10805 -4666
rect 10771 -4769 10805 -4735
rect 10771 -4838 10805 -4804
rect 10771 -4907 10805 -4873
rect 10771 -4976 10805 -4942
rect 10771 -5045 10805 -5011
rect 10771 -5114 10805 -5080
rect 10771 -5183 10805 -5149
rect 10771 -5252 10805 -5218
rect 10771 -5321 10805 -5287
rect 10771 -5390 10805 -5356
rect 10771 -5459 10805 -5425
rect 10771 -5528 10805 -5494
rect 10771 -5597 10805 -5563
rect 10771 -5666 10805 -5632
rect 10771 -5735 10805 -5701
rect 10771 -5804 10805 -5770
rect 10771 -5873 10805 -5839
rect 10771 -5942 10805 -5908
rect 10771 -6011 10805 -5977
rect 10771 -6080 10805 -6046
rect 9453 -6161 9487 -6127
rect 9471 -6272 9505 -6238
rect 10771 -6149 10805 -6115
rect 10771 -6218 10805 -6184
rect 10771 -6287 10805 -6253
rect 9489 -6374 9523 -6340
rect 9560 -6374 9594 -6340
rect 9631 -6374 9665 -6340
rect 9701 -6374 9735 -6340
rect 9771 -6374 9805 -6340
rect 9841 -6374 9875 -6340
rect 9911 -6374 9945 -6340
rect 9981 -6374 10015 -6340
rect 10051 -6374 10085 -6340
rect 10121 -6374 10155 -6340
rect 10191 -6374 10225 -6340
rect 10261 -6374 10295 -6340
rect 10331 -6374 10365 -6340
rect 10401 -6374 10435 -6340
rect 10471 -6374 10505 -6340
rect 10541 -6374 10575 -6340
rect 10611 -6374 10645 -6340
rect 10681 -6374 10715 -6340
rect 10771 -6356 10805 -6322
<< locali >>
rect 8919 22229 10811 22235
rect 8919 22213 8931 22229
rect 8919 22179 8925 22213
rect 8965 22195 9003 22229
rect 9039 22195 9075 22229
rect 9109 22195 9145 22229
rect 9181 22195 9215 22229
rect 9253 22195 9285 22229
rect 9325 22195 9355 22229
rect 9397 22195 9425 22229
rect 9469 22195 9495 22229
rect 9541 22195 9565 22229
rect 9613 22195 9635 22229
rect 9685 22195 9705 22229
rect 9757 22195 9775 22229
rect 9829 22195 9845 22229
rect 9901 22195 9915 22229
rect 9973 22195 9985 22229
rect 10045 22195 10056 22229
rect 10117 22195 10127 22229
rect 10189 22195 10198 22229
rect 10261 22195 10269 22229
rect 10333 22195 10340 22229
rect 10405 22195 10411 22229
rect 10477 22195 10482 22229
rect 10549 22195 10553 22229
rect 10621 22195 10624 22229
rect 10658 22195 10659 22229
rect 10693 22195 10695 22229
rect 10729 22223 10811 22229
rect 10729 22195 10771 22223
rect 8959 22189 10771 22195
rect 8959 22179 8965 22189
rect 8919 22145 8965 22179
rect 8919 22098 8925 22145
rect 8959 22098 8965 22145
rect 8919 22077 8965 22098
rect 8919 22026 8925 22077
rect 8959 22026 8965 22077
rect 8919 22009 8965 22026
rect 8919 21954 8925 22009
rect 8959 21954 8965 22009
rect 10765 22179 10771 22189
rect 10805 22179 10811 22223
rect 10765 22151 10811 22179
rect 10765 22111 10771 22151
rect 10805 22111 10811 22151
rect 10765 22079 10811 22111
rect 10765 22043 10771 22079
rect 10805 22043 10811 22079
rect 10765 22009 10811 22043
rect 8919 21941 8965 21954
rect 8919 21882 8925 21941
rect 8959 21882 8965 21941
rect 8919 21873 8965 21882
rect 8919 21810 8925 21873
rect 8959 21810 8965 21873
rect 9459 21980 9525 21989
rect 9459 21946 9482 21980
rect 9516 21946 9525 21980
rect 9459 21908 9525 21946
rect 9459 21874 9482 21908
rect 9516 21874 9525 21908
rect 9459 21871 9525 21874
rect 9621 21980 9687 21989
rect 9621 21946 9637 21980
rect 9671 21946 9687 21980
rect 9621 21908 9687 21946
rect 9621 21874 9637 21908
rect 9671 21874 9687 21908
rect 9621 21871 9687 21874
rect 9783 21980 9849 21989
rect 9783 21946 9809 21980
rect 9843 21946 9849 21980
rect 9783 21908 9849 21946
rect 9783 21874 9809 21908
rect 9843 21874 9849 21908
rect 9783 21871 9849 21874
rect 9945 21980 10011 21989
rect 9945 21946 9951 21980
rect 9985 21946 10011 21980
rect 9945 21908 10011 21946
rect 9945 21874 9951 21908
rect 9985 21874 10011 21908
rect 9945 21871 10011 21874
rect 10107 21980 10173 21989
rect 10107 21946 10123 21980
rect 10157 21946 10173 21980
rect 10107 21908 10173 21946
rect 10107 21874 10123 21908
rect 10157 21874 10173 21908
rect 10107 21871 10173 21874
rect 10269 21980 10335 21989
rect 10269 21946 10284 21980
rect 10318 21946 10335 21980
rect 10269 21908 10335 21946
rect 10269 21874 10284 21908
rect 10318 21874 10335 21908
rect 10269 21871 10335 21874
rect 10765 21973 10771 22009
rect 10805 21973 10811 22009
rect 10765 21941 10811 21973
rect 10765 21901 10771 21941
rect 10805 21901 10811 21941
rect 10765 21873 10811 21901
rect 8919 21805 8965 21810
rect 8919 21738 8925 21805
rect 8959 21738 8965 21805
rect 8919 21737 8965 21738
rect 8919 21703 8925 21737
rect 8959 21703 8965 21737
rect 8919 21700 8965 21703
rect 8919 21635 8925 21700
rect 8959 21635 8965 21700
rect 8919 21628 8965 21635
rect 8919 21567 8925 21628
rect 8959 21567 8965 21628
rect 8919 21556 8965 21567
rect 8919 21499 8925 21556
rect 8959 21499 8965 21556
rect 8919 21484 8965 21499
rect 8919 21431 8925 21484
rect 8959 21431 8965 21484
rect 8919 21412 8965 21431
rect 8919 21363 8925 21412
rect 8959 21363 8965 21412
rect 8919 21340 8965 21363
rect 8919 21295 8925 21340
rect 8959 21295 8965 21340
rect 8919 21268 8965 21295
rect 8919 21227 8925 21268
rect 8959 21227 8965 21268
rect 8919 21196 8965 21227
rect 8919 21159 8925 21196
rect 8959 21159 8965 21196
rect 8919 21125 8965 21159
rect 8919 21090 8925 21125
rect 8959 21090 8965 21125
rect 8919 21057 8965 21090
rect 8919 21018 8925 21057
rect 8959 21018 8965 21057
rect 8919 20989 8965 21018
rect 8919 20946 8925 20989
rect 8959 20946 8965 20989
rect 8919 20921 8965 20946
rect 8919 20874 8925 20921
rect 8959 20874 8965 20921
rect 8919 20853 8965 20874
rect 8919 20802 8925 20853
rect 8959 20802 8965 20853
rect 8919 20785 8965 20802
rect 8919 20730 8925 20785
rect 8959 20730 8965 20785
rect 8919 20717 8965 20730
rect 8919 20658 8925 20717
rect 8959 20658 8965 20717
rect 8919 20649 8965 20658
rect 8919 20586 8925 20649
rect 8959 20586 8965 20649
rect 8919 20581 8965 20586
rect 8919 20514 8925 20581
rect 8959 20514 8965 20581
rect 8919 20513 8965 20514
rect 8919 20479 8925 20513
rect 8959 20479 8965 20513
rect 8919 20476 8965 20479
rect 8919 20411 8925 20476
rect 8959 20411 8965 20476
rect 8919 20404 8965 20411
rect 8919 20343 8925 20404
rect 8959 20343 8965 20404
rect 8919 20332 8965 20343
rect 8919 20275 8925 20332
rect 8959 20275 8965 20332
rect 8919 20260 8965 20275
rect 8919 20207 8925 20260
rect 8959 20207 8965 20260
rect 8919 20188 8965 20207
rect 8919 20139 8925 20188
rect 8959 20139 8965 20188
rect 8919 20116 8965 20139
rect 8919 20071 8925 20116
rect 8959 20071 8965 20116
rect 8919 20044 8965 20071
rect 8919 20003 8925 20044
rect 8959 20003 8965 20044
rect 8919 19972 8965 20003
rect 8919 19935 8925 19972
rect 8959 19935 8965 19972
rect 8919 19901 8965 19935
rect 8919 19866 8925 19901
rect 8959 19866 8965 19901
rect 8919 19833 8965 19866
rect 8919 19794 8925 19833
rect 8959 19794 8965 19833
rect 8919 19765 8965 19794
rect 8919 19722 8925 19765
rect 8959 19722 8965 19765
rect 8919 19697 8965 19722
rect 8919 19650 8925 19697
rect 8959 19650 8965 19697
rect 8919 19629 8965 19650
rect 8919 19578 8925 19629
rect 8959 19578 8965 19629
rect 8919 19561 8965 19578
rect 8919 19506 8925 19561
rect 8959 19506 8965 19561
rect 8919 19493 8965 19506
rect 8919 19434 8925 19493
rect 8959 19434 8965 19493
rect 8919 19425 8965 19434
rect 8919 19362 8925 19425
rect 8959 19362 8965 19425
rect 8919 19357 8965 19362
rect 8919 19290 8925 19357
rect 8959 19290 8965 19357
rect 8919 19289 8965 19290
rect 8919 19255 8925 19289
rect 8959 19255 8965 19289
rect 8919 19252 8965 19255
rect 8919 19187 8925 19252
rect 8959 19187 8965 19252
rect 8919 19180 8965 19187
rect 8919 19119 8925 19180
rect 8959 19119 8965 19180
rect 8919 19108 8965 19119
rect 8919 19051 8925 19108
rect 8959 19051 8965 19108
rect 8919 19036 8965 19051
rect 8919 18983 8925 19036
rect 8959 18983 8965 19036
rect 8919 18964 8965 18983
rect 8919 18915 8925 18964
rect 8959 18915 8965 18964
rect 8919 18892 8965 18915
rect 8919 18847 8925 18892
rect 8959 18847 8965 18892
rect 8919 18820 8965 18847
rect 8919 18779 8925 18820
rect 8959 18779 8965 18820
rect 8919 18748 8965 18779
rect 8919 18711 8925 18748
rect 8959 18711 8965 18748
rect 8919 18677 8965 18711
rect 8919 18642 8925 18677
rect 8959 18642 8965 18677
rect 8919 18609 8965 18642
rect 8919 18570 8925 18609
rect 8959 18570 8965 18609
rect 8919 18541 8965 18570
rect 8919 18498 8925 18541
rect 8959 18498 8965 18541
rect 8919 18473 8965 18498
rect 8919 18426 8925 18473
rect 8959 18426 8965 18473
rect 8919 18405 8965 18426
rect 8919 18354 8925 18405
rect 8959 18354 8965 18405
rect 8919 18337 8965 18354
rect 8919 18282 8925 18337
rect 8959 18282 8965 18337
rect 8919 18269 8965 18282
rect 8919 18210 8925 18269
rect 8959 18210 8965 18269
rect 8919 18201 8965 18210
rect 8919 18138 8925 18201
rect 8959 18138 8965 18201
rect 8919 18133 8965 18138
rect 8919 18066 8925 18133
rect 8959 18066 8965 18133
rect 8919 18065 8965 18066
rect 8919 18031 8925 18065
rect 8959 18031 8965 18065
rect 8919 18028 8965 18031
rect 8919 17963 8925 18028
rect 8959 17963 8965 18028
rect 8919 17956 8965 17963
rect 8919 17895 8925 17956
rect 8959 17895 8965 17956
rect 8919 17884 8965 17895
rect 8919 17827 8925 17884
rect 8959 17827 8965 17884
rect 8919 17812 8965 17827
rect 8919 17759 8925 17812
rect 8959 17759 8965 17812
rect 8919 17740 8965 17759
rect 8919 17691 8925 17740
rect 8959 17691 8965 17740
rect 8919 17668 8965 17691
rect 8919 17623 8925 17668
rect 8959 17623 8965 17668
rect 8919 17596 8965 17623
rect 8919 17555 8925 17596
rect 8959 17555 8965 17596
rect 8919 17524 8965 17555
rect 8919 17487 8925 17524
rect 8959 17487 8965 17524
rect 8919 17453 8965 17487
rect 8919 17418 8925 17453
rect 8959 17418 8965 17453
rect 8919 17385 8965 17418
rect 8919 17346 8925 17385
rect 8959 17346 8965 17385
rect 8919 17317 8965 17346
rect 8919 17274 8925 17317
rect 8959 17274 8965 17317
rect 8919 17249 8965 17274
rect 8919 17202 8925 17249
rect 8959 17202 8965 17249
rect 8919 17181 8965 17202
rect 8919 17130 8925 17181
rect 8959 17130 8965 17181
rect 8919 17113 8965 17130
rect 8919 17058 8925 17113
rect 8959 17058 8965 17113
rect 8919 17045 8965 17058
rect 8919 16986 8925 17045
rect 8959 16986 8965 17045
rect 8919 16977 8965 16986
rect 8919 16914 8925 16977
rect 8959 16914 8965 16977
rect 8919 16909 8965 16914
rect 8919 16842 8925 16909
rect 8959 16842 8965 16909
rect 8919 16841 8965 16842
rect 8919 16807 8925 16841
rect 8959 16807 8965 16841
rect 8919 16804 8965 16807
rect 8919 16739 8925 16804
rect 8959 16739 8965 16804
rect 8919 16732 8965 16739
rect 8919 16671 8925 16732
rect 8959 16671 8965 16732
rect 8919 16660 8965 16671
rect 8919 16603 8925 16660
rect 8959 16603 8965 16660
rect 8919 16588 8965 16603
rect 8919 16535 8925 16588
rect 8959 16535 8965 16588
rect 8919 16516 8965 16535
rect 8919 16467 8925 16516
rect 8959 16467 8965 16516
rect 8919 16444 8965 16467
rect 8919 16399 8925 16444
rect 8959 16399 8965 16444
rect 8919 16372 8965 16399
rect 8919 16331 8925 16372
rect 8959 16331 8965 16372
rect 8919 16300 8965 16331
rect 8919 16263 8925 16300
rect 8959 16263 8965 16300
rect 8919 16229 8965 16263
rect 8919 16194 8925 16229
rect 8959 16194 8965 16229
rect 8919 16161 8965 16194
rect 8919 16122 8925 16161
rect 8959 16122 8965 16161
rect 8919 16093 8965 16122
rect 8919 16050 8925 16093
rect 8959 16050 8965 16093
rect 8919 16025 8965 16050
rect 8919 15978 8925 16025
rect 8959 15978 8965 16025
rect 8919 15957 8965 15978
rect 8919 15906 8925 15957
rect 8959 15906 8965 15957
rect 8919 15889 8965 15906
rect 8919 15834 8925 15889
rect 8959 15834 8965 15889
rect 8919 15821 8965 15834
rect 8919 15762 8925 15821
rect 8959 15762 8965 15821
rect 8919 15753 8965 15762
rect 8919 15690 8925 15753
rect 8959 15690 8965 15753
rect 8919 15685 8965 15690
rect 8919 15618 8925 15685
rect 8959 15618 8965 15685
rect 8919 15617 8965 15618
rect 8919 15583 8925 15617
rect 8959 15583 8965 15617
rect 8919 15580 8965 15583
rect 8919 15515 8925 15580
rect 8959 15515 8965 15580
rect 8919 15508 8965 15515
rect 8919 15447 8925 15508
rect 8959 15447 8965 15508
rect 8919 15436 8965 15447
rect 8919 15379 8925 15436
rect 8959 15379 8965 15436
rect 8919 15364 8965 15379
rect 8919 15311 8925 15364
rect 8959 15311 8965 15364
rect 8919 15292 8965 15311
rect 8919 15243 8925 15292
rect 8959 15243 8965 15292
rect 8919 15220 8965 15243
rect 8919 15175 8925 15220
rect 8959 15175 8965 15220
rect 8919 15148 8965 15175
rect 8919 15107 8925 15148
rect 8959 15107 8965 15148
rect 8919 15076 8965 15107
rect 8919 15039 8925 15076
rect 8959 15039 8965 15076
rect 8919 15005 8965 15039
rect 8919 14970 8925 15005
rect 8959 14970 8965 15005
rect 8919 14937 8965 14970
rect 8919 14898 8925 14937
rect 8959 14898 8965 14937
rect 8919 14869 8965 14898
rect 8919 14826 8925 14869
rect 8959 14826 8965 14869
rect 8919 14801 8965 14826
rect 8919 14754 8925 14801
rect 8959 14754 8965 14801
rect 8919 14733 8965 14754
rect 8919 14682 8925 14733
rect 8959 14682 8965 14733
rect 8919 14665 8965 14682
rect 8919 14610 8925 14665
rect 8959 14610 8965 14665
rect 8919 14597 8965 14610
rect 8919 14538 8925 14597
rect 8959 14538 8965 14597
rect 8919 14529 8965 14538
rect 8919 14466 8925 14529
rect 8959 14466 8965 14529
rect 8919 14461 8965 14466
rect 8919 14394 8925 14461
rect 8959 14394 8965 14461
rect 8919 14393 8965 14394
rect 8919 14359 8925 14393
rect 8959 14359 8965 14393
rect 8919 14356 8965 14359
rect 8919 14291 8925 14356
rect 8959 14291 8965 14356
rect 8919 14284 8965 14291
rect 8919 14223 8925 14284
rect 8959 14223 8965 14284
rect 8919 14212 8965 14223
rect 8919 14155 8925 14212
rect 8959 14155 8965 14212
rect 8919 14140 8965 14155
rect 8919 14087 8925 14140
rect 8959 14087 8965 14140
rect 8919 14068 8965 14087
rect 8919 14019 8925 14068
rect 8959 14019 8965 14068
rect 8919 13996 8965 14019
rect 8919 13951 8925 13996
rect 8959 13951 8965 13996
rect 8919 13924 8965 13951
rect 8919 13883 8925 13924
rect 8959 13883 8965 13924
rect 8919 13852 8965 13883
rect 8919 13815 8925 13852
rect 8959 13815 8965 13852
rect 8919 13781 8965 13815
rect 8919 13746 8925 13781
rect 8959 13746 8965 13781
rect 8919 13713 8965 13746
rect 8919 13674 8925 13713
rect 8959 13674 8965 13713
rect 8919 13645 8965 13674
rect 8919 13602 8925 13645
rect 8959 13602 8965 13645
rect 8919 13577 8965 13602
rect 8919 13530 8925 13577
rect 8959 13530 8965 13577
rect 8919 13509 8965 13530
rect 8919 13458 8925 13509
rect 8959 13458 8965 13509
rect 8919 13441 8965 13458
rect 8919 13386 8925 13441
rect 8959 13386 8965 13441
rect 8919 13373 8965 13386
rect 8919 13314 8925 13373
rect 8959 13314 8965 13373
rect 8919 13305 8965 13314
rect 8919 13242 8925 13305
rect 8959 13242 8965 13305
rect 8919 13237 8965 13242
rect 8919 13170 8925 13237
rect 8959 13170 8965 13237
rect 8919 13169 8965 13170
rect 8919 13135 8925 13169
rect 8959 13135 8965 13169
rect 8919 13132 8965 13135
rect 8919 13067 8925 13132
rect 8959 13067 8965 13132
rect 8919 13060 8965 13067
rect 8919 12999 8925 13060
rect 8959 12999 8965 13060
rect 8919 12988 8965 12999
rect 8919 12931 8925 12988
rect 8959 12931 8965 12988
rect 8919 12916 8965 12931
rect 8919 12863 8925 12916
rect 8959 12863 8965 12916
rect 8919 12844 8965 12863
rect 8919 12795 8925 12844
rect 8959 12795 8965 12844
rect 8919 12772 8965 12795
rect 8919 12727 8925 12772
rect 8959 12727 8965 12772
rect 8919 12700 8965 12727
rect 8919 12659 8925 12700
rect 8959 12659 8965 12700
rect 8919 12628 8965 12659
rect 8919 12591 8925 12628
rect 8959 12591 8965 12628
rect 10765 21829 10771 21873
rect 10805 21829 10811 21873
rect 10765 21805 10811 21829
rect 10765 21757 10771 21805
rect 10805 21757 10811 21805
rect 10765 21737 10811 21757
rect 10765 21685 10771 21737
rect 10805 21685 10811 21737
rect 10765 21669 10811 21685
rect 10765 21613 10771 21669
rect 10805 21613 10811 21669
rect 10765 21601 10811 21613
rect 10765 21541 10771 21601
rect 10805 21541 10811 21601
rect 10765 21533 10811 21541
rect 10765 21469 10771 21533
rect 10805 21469 10811 21533
rect 10765 21465 10811 21469
rect 10765 21363 10771 21465
rect 10805 21363 10811 21465
rect 10765 21359 10811 21363
rect 10765 21295 10771 21359
rect 10805 21295 10811 21359
rect 10765 21287 10811 21295
rect 10765 21227 10771 21287
rect 10805 21227 10811 21287
rect 10765 21215 10811 21227
rect 10765 21159 10771 21215
rect 10805 21159 10811 21215
rect 10765 21143 10811 21159
rect 10765 21091 10771 21143
rect 10805 21091 10811 21143
rect 10765 21071 10811 21091
rect 10765 21023 10771 21071
rect 10805 21023 10811 21071
rect 10765 20999 10811 21023
rect 10765 20955 10771 20999
rect 10805 20955 10811 20999
rect 10765 20927 10811 20955
rect 10765 20887 10771 20927
rect 10805 20887 10811 20927
rect 10765 20855 10811 20887
rect 10765 20819 10771 20855
rect 10805 20819 10811 20855
rect 10765 20785 10811 20819
rect 10765 20749 10771 20785
rect 10805 20749 10811 20785
rect 10765 20717 10811 20749
rect 10765 20677 10771 20717
rect 10805 20677 10811 20717
rect 10765 20649 10811 20677
rect 10765 20605 10771 20649
rect 10805 20605 10811 20649
rect 10765 20581 10811 20605
rect 10765 20533 10771 20581
rect 10805 20533 10811 20581
rect 10765 20513 10811 20533
rect 10765 20461 10771 20513
rect 10805 20461 10811 20513
rect 10765 20445 10811 20461
rect 10765 20389 10771 20445
rect 10805 20389 10811 20445
rect 10765 20377 10811 20389
rect 10765 20317 10771 20377
rect 10805 20317 10811 20377
rect 10765 20309 10811 20317
rect 10765 20245 10771 20309
rect 10805 20245 10811 20309
rect 10765 20241 10811 20245
rect 10765 20139 10771 20241
rect 10805 20139 10811 20241
rect 10765 20135 10811 20139
rect 10765 20071 10771 20135
rect 10805 20071 10811 20135
rect 10765 20063 10811 20071
rect 10765 20003 10771 20063
rect 10805 20003 10811 20063
rect 10765 19991 10811 20003
rect 10765 19935 10771 19991
rect 10805 19935 10811 19991
rect 10765 19919 10811 19935
rect 10765 19867 10771 19919
rect 10805 19867 10811 19919
rect 10765 19847 10811 19867
rect 10765 19799 10771 19847
rect 10805 19799 10811 19847
rect 10765 19775 10811 19799
rect 10765 19731 10771 19775
rect 10805 19731 10811 19775
rect 10765 19703 10811 19731
rect 10765 19663 10771 19703
rect 10805 19663 10811 19703
rect 10765 19631 10811 19663
rect 10765 19595 10771 19631
rect 10805 19595 10811 19631
rect 10765 19561 10811 19595
rect 10765 19525 10771 19561
rect 10805 19525 10811 19561
rect 10765 19493 10811 19525
rect 10765 19453 10771 19493
rect 10805 19453 10811 19493
rect 10765 19425 10811 19453
rect 10765 19381 10771 19425
rect 10805 19381 10811 19425
rect 10765 19357 10811 19381
rect 10765 19309 10771 19357
rect 10805 19309 10811 19357
rect 10765 19289 10811 19309
rect 10765 19237 10771 19289
rect 10805 19237 10811 19289
rect 10765 19221 10811 19237
rect 10765 19165 10771 19221
rect 10805 19165 10811 19221
rect 10765 19153 10811 19165
rect 10765 19093 10771 19153
rect 10805 19093 10811 19153
rect 10765 19085 10811 19093
rect 10765 19021 10771 19085
rect 10805 19021 10811 19085
rect 10765 19017 10811 19021
rect 10765 18915 10771 19017
rect 10805 18915 10811 19017
rect 10765 18911 10811 18915
rect 10765 18847 10771 18911
rect 10805 18847 10811 18911
rect 10765 18839 10811 18847
rect 10765 18779 10771 18839
rect 10805 18779 10811 18839
rect 10765 18767 10811 18779
rect 10765 18711 10771 18767
rect 10805 18711 10811 18767
rect 10765 18695 10811 18711
rect 10765 18643 10771 18695
rect 10805 18643 10811 18695
rect 10765 18623 10811 18643
rect 10765 18575 10771 18623
rect 10805 18575 10811 18623
rect 10765 18551 10811 18575
rect 10765 18507 10771 18551
rect 10805 18507 10811 18551
rect 10765 18479 10811 18507
rect 10765 18439 10771 18479
rect 10805 18439 10811 18479
rect 10765 18407 10811 18439
rect 10765 18371 10771 18407
rect 10805 18371 10811 18407
rect 10765 18337 10811 18371
rect 10765 18301 10771 18337
rect 10805 18301 10811 18337
rect 10765 18269 10811 18301
rect 10765 18229 10771 18269
rect 10805 18229 10811 18269
rect 10765 18201 10811 18229
rect 10765 18157 10771 18201
rect 10805 18157 10811 18201
rect 10765 18133 10811 18157
rect 10765 18085 10771 18133
rect 10805 18085 10811 18133
rect 10765 18065 10811 18085
rect 10765 18013 10771 18065
rect 10805 18013 10811 18065
rect 10765 17997 10811 18013
rect 10765 17941 10771 17997
rect 10805 17941 10811 17997
rect 10765 17929 10811 17941
rect 10765 17869 10771 17929
rect 10805 17869 10811 17929
rect 10765 17861 10811 17869
rect 10765 17797 10771 17861
rect 10805 17797 10811 17861
rect 10765 17793 10811 17797
rect 10765 17691 10771 17793
rect 10805 17691 10811 17793
rect 10765 17687 10811 17691
rect 10765 17623 10771 17687
rect 10805 17623 10811 17687
rect 10765 17615 10811 17623
rect 10765 17555 10771 17615
rect 10805 17555 10811 17615
rect 10765 17543 10811 17555
rect 10765 17487 10771 17543
rect 10805 17487 10811 17543
rect 10765 17471 10811 17487
rect 10765 17419 10771 17471
rect 10805 17419 10811 17471
rect 10765 17399 10811 17419
rect 10765 17351 10771 17399
rect 10805 17351 10811 17399
rect 10765 17327 10811 17351
rect 10765 17283 10771 17327
rect 10805 17283 10811 17327
rect 10765 17255 10811 17283
rect 10765 17215 10771 17255
rect 10805 17215 10811 17255
rect 10765 17183 10811 17215
rect 10765 17147 10771 17183
rect 10805 17147 10811 17183
rect 10765 17113 10811 17147
rect 10765 17077 10771 17113
rect 10805 17077 10811 17113
rect 10765 17045 10811 17077
rect 10765 17005 10771 17045
rect 10805 17005 10811 17045
rect 10765 16977 10811 17005
rect 10765 16933 10771 16977
rect 10805 16933 10811 16977
rect 10765 16909 10811 16933
rect 10765 16861 10771 16909
rect 10805 16861 10811 16909
rect 10765 16841 10811 16861
rect 10765 16789 10771 16841
rect 10805 16789 10811 16841
rect 10765 16773 10811 16789
rect 10765 16717 10771 16773
rect 10805 16717 10811 16773
rect 10765 16705 10811 16717
rect 10765 16645 10771 16705
rect 10805 16645 10811 16705
rect 10765 16637 10811 16645
rect 10765 16573 10771 16637
rect 10805 16573 10811 16637
rect 10765 16569 10811 16573
rect 10765 16467 10771 16569
rect 10805 16467 10811 16569
rect 10765 16463 10811 16467
rect 10765 16399 10771 16463
rect 10805 16399 10811 16463
rect 10765 16391 10811 16399
rect 10765 16331 10771 16391
rect 10805 16331 10811 16391
rect 10765 16319 10811 16331
rect 10765 16263 10771 16319
rect 10805 16263 10811 16319
rect 10765 16247 10811 16263
rect 10765 16195 10771 16247
rect 10805 16195 10811 16247
rect 10765 16175 10811 16195
rect 10765 16127 10771 16175
rect 10805 16127 10811 16175
rect 10765 16103 10811 16127
rect 10765 16059 10771 16103
rect 10805 16059 10811 16103
rect 10765 16031 10811 16059
rect 10765 15991 10771 16031
rect 10805 15991 10811 16031
rect 10765 15959 10811 15991
rect 10765 15923 10771 15959
rect 10805 15923 10811 15959
rect 10765 15889 10811 15923
rect 10765 15853 10771 15889
rect 10805 15853 10811 15889
rect 10765 15821 10811 15853
rect 10765 15781 10771 15821
rect 10805 15781 10811 15821
rect 10765 15753 10811 15781
rect 10765 15709 10771 15753
rect 10805 15709 10811 15753
rect 10765 15685 10811 15709
rect 10765 15637 10771 15685
rect 10805 15637 10811 15685
rect 10765 15617 10811 15637
rect 10765 15565 10771 15617
rect 10805 15565 10811 15617
rect 10765 15549 10811 15565
rect 10765 15493 10771 15549
rect 10805 15493 10811 15549
rect 10765 15481 10811 15493
rect 10765 15421 10771 15481
rect 10805 15421 10811 15481
rect 10765 15413 10811 15421
rect 10765 15349 10771 15413
rect 10805 15349 10811 15413
rect 10765 15345 10811 15349
rect 10765 15243 10771 15345
rect 10805 15243 10811 15345
rect 10765 15239 10811 15243
rect 10765 15175 10771 15239
rect 10805 15175 10811 15239
rect 10765 15167 10811 15175
rect 10765 15107 10771 15167
rect 10805 15107 10811 15167
rect 10765 15095 10811 15107
rect 10765 15039 10771 15095
rect 10805 15039 10811 15095
rect 10765 15023 10811 15039
rect 10765 14971 10771 15023
rect 10805 14971 10811 15023
rect 10765 14951 10811 14971
rect 10765 14903 10771 14951
rect 10805 14903 10811 14951
rect 10765 14879 10811 14903
rect 10765 14835 10771 14879
rect 10805 14835 10811 14879
rect 10765 14807 10811 14835
rect 10765 14767 10771 14807
rect 10805 14767 10811 14807
rect 10765 14735 10811 14767
rect 10765 14699 10771 14735
rect 10805 14699 10811 14735
rect 10765 14665 10811 14699
rect 10765 14629 10771 14665
rect 10805 14629 10811 14665
rect 10765 14597 10811 14629
rect 10765 14557 10771 14597
rect 10805 14557 10811 14597
rect 10765 14529 10811 14557
rect 10765 14485 10771 14529
rect 10805 14485 10811 14529
rect 10765 14461 10811 14485
rect 10765 14413 10771 14461
rect 10805 14413 10811 14461
rect 10765 14393 10811 14413
rect 10765 14341 10771 14393
rect 10805 14341 10811 14393
rect 10765 14325 10811 14341
rect 10765 14269 10771 14325
rect 10805 14269 10811 14325
rect 10765 14257 10811 14269
rect 10765 14197 10771 14257
rect 10805 14197 10811 14257
rect 10765 14189 10811 14197
rect 10765 14125 10771 14189
rect 10805 14125 10811 14189
rect 10765 14121 10811 14125
rect 10765 14019 10771 14121
rect 10805 14019 10811 14121
rect 10765 14015 10811 14019
rect 10765 13951 10771 14015
rect 10805 13951 10811 14015
rect 10765 13943 10811 13951
rect 10765 13883 10771 13943
rect 10805 13883 10811 13943
rect 10765 13871 10811 13883
rect 10765 13815 10771 13871
rect 10805 13815 10811 13871
rect 10765 13799 10811 13815
rect 10765 13747 10771 13799
rect 10805 13747 10811 13799
rect 10765 13727 10811 13747
rect 10765 13679 10771 13727
rect 10805 13679 10811 13727
rect 10765 13655 10811 13679
rect 10765 13611 10771 13655
rect 10805 13611 10811 13655
rect 10765 13583 10811 13611
rect 10765 13543 10771 13583
rect 10805 13543 10811 13583
rect 10765 13511 10811 13543
rect 10765 13475 10771 13511
rect 10805 13475 10811 13511
rect 10765 13441 10811 13475
rect 10765 13405 10771 13441
rect 10805 13405 10811 13441
rect 10765 13373 10811 13405
rect 10765 13333 10771 13373
rect 10805 13333 10811 13373
rect 10765 13305 10811 13333
rect 10765 13261 10771 13305
rect 10805 13261 10811 13305
rect 10765 13237 10811 13261
rect 10765 13189 10771 13237
rect 10805 13189 10811 13237
rect 10765 13169 10811 13189
rect 10765 13117 10771 13169
rect 10805 13117 10811 13169
rect 10765 13101 10811 13117
rect 10765 13045 10771 13101
rect 10805 13045 10811 13101
rect 10765 13033 10811 13045
rect 10765 12973 10771 13033
rect 10805 12973 10811 13033
rect 10765 12965 10811 12973
rect 10765 12901 10771 12965
rect 10805 12901 10811 12965
rect 10765 12897 10811 12901
rect 10765 12795 10771 12897
rect 10805 12795 10811 12897
rect 10765 12791 10811 12795
rect 10765 12727 10771 12791
rect 10805 12727 10811 12791
rect 10765 12719 10811 12727
rect 10765 12659 10771 12719
rect 10805 12659 10811 12719
rect 10765 12647 10811 12659
rect 8919 12557 8965 12591
rect 8919 12522 8925 12557
rect 8959 12522 8965 12557
rect 8919 12489 8965 12522
rect 10269 12593 10284 12627
rect 10318 12593 10335 12627
rect 10269 12555 10335 12593
rect 10269 12521 10284 12555
rect 10318 12521 10335 12555
rect 10269 12509 10335 12521
rect 10765 12591 10771 12647
rect 10805 12591 10811 12647
rect 10765 12575 10811 12591
rect 10765 12523 10771 12575
rect 10805 12523 10811 12575
rect 8919 12450 8925 12489
rect 8959 12450 8965 12489
rect 8919 12421 8965 12450
rect 8919 12378 8925 12421
rect 8959 12378 8965 12421
rect 8919 12353 8965 12378
rect 8919 12306 8925 12353
rect 8959 12306 8965 12353
rect 8919 12285 8965 12306
rect 8919 12234 8925 12285
rect 8959 12234 8965 12285
rect 8919 12217 8965 12234
rect 8919 12162 8925 12217
rect 8959 12162 8965 12217
rect 8919 12149 8965 12162
rect 8919 12090 8925 12149
rect 8959 12090 8965 12149
rect 8919 12081 8965 12090
rect 8919 12018 8925 12081
rect 8959 12018 8965 12081
rect 8919 12013 8965 12018
rect 8919 11946 8925 12013
rect 8959 11946 8965 12013
rect 8919 11945 8965 11946
rect 8919 11911 8925 11945
rect 8959 11911 8965 11945
rect 8919 11908 8965 11911
rect 8919 11843 8925 11908
rect 8959 11843 8965 11908
rect 8919 11836 8965 11843
rect 8919 11775 8925 11836
rect 8959 11775 8965 11836
rect 8919 11764 8965 11775
rect 8919 11707 8925 11764
rect 8959 11707 8965 11764
rect 8919 11692 8965 11707
rect 8919 11639 8925 11692
rect 8959 11639 8965 11692
rect 8919 11620 8965 11639
rect 8919 11571 8925 11620
rect 8959 11571 8965 11620
rect 8919 11548 8965 11571
rect 8919 11503 8925 11548
rect 8959 11503 8965 11548
rect 8919 11476 8965 11503
rect 8919 11435 8925 11476
rect 8959 11435 8965 11476
rect 8919 11404 8965 11435
rect 8919 11367 8925 11404
rect 8959 11367 8965 11404
rect 8919 11333 8965 11367
rect 8919 11298 8925 11333
rect 8959 11298 8965 11333
rect 8919 11265 8965 11298
rect 8919 11226 8925 11265
rect 8959 11226 8965 11265
rect 8919 11197 8965 11226
rect 8919 11154 8925 11197
rect 8959 11154 8965 11197
rect 8919 11129 8965 11154
rect 8919 11082 8925 11129
rect 8959 11082 8965 11129
rect 8919 11061 8965 11082
rect 8919 11010 8925 11061
rect 8959 11010 8965 11061
rect 8919 10993 8965 11010
rect 8919 10938 8925 10993
rect 8959 10938 8965 10993
rect 8919 10925 8965 10938
rect 8919 10866 8925 10925
rect 8959 10866 8965 10925
rect 8919 10857 8965 10866
rect 8919 10794 8925 10857
rect 8959 10794 8965 10857
rect 8919 10789 8965 10794
rect 8919 10722 8925 10789
rect 8959 10722 8965 10789
rect 8919 10721 8965 10722
rect 8919 10687 8925 10721
rect 8959 10687 8965 10721
rect 8919 10684 8965 10687
rect 8919 10619 8925 10684
rect 8959 10619 8965 10684
rect 8919 10612 8965 10619
rect 8919 10551 8925 10612
rect 8959 10551 8965 10612
rect 8919 10540 8965 10551
rect 8919 10483 8925 10540
rect 8959 10483 8965 10540
rect 8919 10468 8965 10483
rect 8919 10415 8925 10468
rect 8959 10415 8965 10468
rect 8919 10396 8965 10415
rect 8919 10347 8925 10396
rect 8959 10347 8965 10396
rect 8919 10324 8965 10347
rect 8919 10279 8925 10324
rect 8959 10279 8965 10324
rect 8919 10252 8965 10279
rect 8919 10211 8925 10252
rect 8959 10211 8965 10252
rect 8919 10180 8965 10211
rect 8919 10143 8925 10180
rect 8959 10143 8965 10180
rect 8919 10109 8965 10143
rect 8919 10074 8925 10109
rect 8959 10074 8965 10109
rect 8919 10041 8965 10074
rect 8919 10002 8925 10041
rect 8959 10002 8965 10041
rect 8919 9973 8965 10002
rect 8919 9930 8925 9973
rect 8959 9930 8965 9973
rect 8919 9905 8965 9930
rect 8919 9858 8925 9905
rect 8959 9858 8965 9905
rect 8919 9837 8965 9858
rect 8919 9786 8925 9837
rect 8959 9786 8965 9837
rect 8919 9769 8965 9786
rect 8919 9714 8925 9769
rect 8959 9714 8965 9769
rect 8919 9701 8965 9714
rect 8919 9642 8925 9701
rect 8959 9642 8965 9701
rect 8919 9633 8965 9642
rect 8919 9570 8925 9633
rect 8959 9570 8965 9633
rect 8919 9565 8965 9570
rect 8919 9498 8925 9565
rect 8959 9498 8965 9565
rect 8919 9497 8965 9498
rect 8919 9463 8925 9497
rect 8959 9463 8965 9497
rect 8919 9460 8965 9463
rect 8919 9395 8925 9460
rect 8959 9395 8965 9460
rect 8919 9388 8965 9395
rect 8919 9327 8925 9388
rect 8959 9327 8965 9388
rect 8919 9316 8965 9327
rect 8919 9259 8925 9316
rect 8959 9259 8965 9316
rect 8919 9244 8965 9259
rect 8919 9191 8925 9244
rect 8959 9191 8965 9244
rect 8919 9172 8965 9191
rect 8919 9123 8925 9172
rect 8959 9123 8965 9172
rect 8919 9100 8965 9123
rect 8919 9055 8925 9100
rect 8959 9055 8965 9100
rect 8919 9028 8965 9055
rect 8919 8987 8925 9028
rect 8959 8987 8965 9028
rect 8919 8956 8965 8987
rect 8919 8919 8925 8956
rect 8959 8919 8965 8956
rect 8919 8885 8965 8919
rect 8919 8850 8925 8885
rect 8959 8850 8965 8885
rect 8919 8817 8965 8850
rect 8919 8778 8925 8817
rect 8959 8778 8965 8817
rect 8919 8749 8965 8778
rect 8919 8706 8925 8749
rect 8959 8706 8965 8749
rect 8919 8681 8965 8706
rect 8919 8634 8925 8681
rect 8959 8634 8965 8681
rect 8919 8613 8965 8634
rect 8919 8562 8925 8613
rect 8959 8562 8965 8613
rect 8919 8545 8965 8562
rect 8919 8490 8925 8545
rect 8959 8490 8965 8545
rect 8919 8477 8965 8490
rect 8919 8418 8925 8477
rect 8959 8418 8965 8477
rect 8919 8409 8965 8418
rect 8919 8346 8925 8409
rect 8959 8346 8965 8409
rect 8919 8341 8965 8346
rect 8919 8274 8925 8341
rect 8959 8274 8965 8341
rect 8919 8273 8965 8274
rect 8919 8239 8925 8273
rect 8959 8239 8965 8273
rect 8919 8236 8965 8239
rect 8919 8171 8925 8236
rect 8959 8171 8965 8236
rect 8919 8164 8965 8171
rect 8919 8103 8925 8164
rect 8959 8103 8965 8164
rect 8919 8092 8965 8103
rect 8919 8035 8925 8092
rect 8959 8035 8965 8092
rect 8919 8020 8965 8035
rect 8919 7967 8925 8020
rect 8959 7967 8965 8020
rect 8919 7948 8965 7967
rect 8919 7899 8925 7948
rect 8959 7899 8965 7948
rect 8919 7876 8965 7899
rect 8919 7831 8925 7876
rect 8959 7831 8965 7876
rect 8919 7804 8965 7831
rect 8919 7763 8925 7804
rect 8959 7763 8965 7804
rect 8919 7732 8965 7763
rect 8919 7695 8925 7732
rect 8959 7695 8965 7732
rect 8919 7661 8965 7695
rect 8919 7626 8925 7661
rect 8959 7626 8965 7661
rect 8919 7593 8965 7626
rect 8919 7554 8925 7593
rect 8959 7554 8965 7593
rect 8919 7525 8965 7554
rect 8919 7482 8925 7525
rect 8959 7482 8965 7525
rect 8919 7457 8965 7482
rect 8919 7410 8925 7457
rect 8959 7410 8965 7457
rect 8919 7389 8965 7410
rect 8919 7338 8925 7389
rect 8959 7338 8965 7389
rect 8919 7321 8965 7338
rect 8919 7266 8925 7321
rect 8959 7266 8965 7321
rect 8919 7253 8965 7266
rect 8919 7194 8925 7253
rect 8959 7194 8965 7253
rect 8919 7185 8965 7194
rect 8919 7122 8925 7185
rect 8959 7122 8965 7185
rect 8919 7117 8965 7122
rect 8919 7050 8925 7117
rect 8959 7050 8965 7117
rect 8919 7049 8965 7050
rect 8919 7015 8925 7049
rect 8959 7015 8965 7049
rect 8919 7012 8965 7015
rect 8919 6947 8925 7012
rect 8959 6947 8965 7012
rect 8919 6940 8965 6947
rect 8919 6879 8925 6940
rect 8959 6879 8965 6940
rect 8919 6868 8965 6879
rect 8919 6811 8925 6868
rect 8959 6811 8965 6868
rect 8919 6796 8965 6811
rect 8919 6743 8925 6796
rect 8959 6743 8965 6796
rect 8919 6724 8965 6743
rect 8919 6675 8925 6724
rect 8959 6675 8965 6724
rect 8919 6652 8965 6675
rect 8919 6607 8925 6652
rect 8959 6607 8965 6652
rect 8919 6580 8965 6607
rect 8919 6539 8925 6580
rect 8959 6539 8965 6580
rect 8919 6508 8965 6539
rect 8919 6471 8925 6508
rect 8959 6471 8965 6508
rect 8919 6437 8965 6471
rect 8919 6402 8925 6437
rect 8959 6402 8965 6437
rect 8919 6369 8965 6402
rect 8919 6330 8925 6369
rect 8959 6330 8965 6369
rect 8919 6301 8965 6330
rect 8919 6258 8925 6301
rect 8959 6258 8965 6301
rect 8919 6233 8965 6258
rect 8919 6186 8925 6233
rect 8959 6186 8965 6233
rect 8919 6165 8965 6186
rect 8919 6114 8925 6165
rect 8959 6114 8965 6165
rect 8919 6097 8965 6114
rect 8919 6042 8925 6097
rect 8959 6042 8965 6097
rect 8919 6029 8965 6042
rect 8919 5970 8925 6029
rect 8959 5970 8965 6029
rect 8919 5961 8965 5970
rect 8919 5898 8925 5961
rect 8959 5898 8965 5961
rect 8919 5893 8965 5898
rect 8919 5826 8925 5893
rect 8959 5826 8965 5893
rect 8919 5825 8965 5826
rect 8919 5791 8925 5825
rect 8959 5791 8965 5825
rect 8919 5788 8965 5791
rect 8919 5723 8925 5788
rect 8959 5723 8965 5788
rect 8919 5716 8965 5723
rect 8919 5655 8925 5716
rect 8959 5655 8965 5716
rect 8919 5644 8965 5655
rect 8919 5587 8925 5644
rect 8959 5587 8965 5644
rect 8919 5572 8965 5587
rect 8919 5519 8925 5572
rect 8959 5519 8965 5572
rect 8919 5500 8965 5519
rect 8919 5451 8925 5500
rect 8959 5451 8965 5500
rect 8919 5428 8965 5451
rect 8919 5383 8925 5428
rect 8959 5383 8965 5428
rect 8919 5356 8965 5383
rect 8919 5315 8925 5356
rect 8959 5315 8965 5356
rect 8919 5284 8965 5315
rect 8919 5247 8925 5284
rect 8959 5247 8965 5284
rect 8919 5213 8965 5247
rect 8919 5178 8925 5213
rect 8959 5178 8965 5213
rect 8919 5145 8965 5178
rect 8919 5106 8925 5145
rect 8959 5106 8965 5145
rect 8919 5077 8965 5106
rect 8919 5034 8925 5077
rect 8959 5034 8965 5077
rect 8919 5009 8965 5034
rect 8919 4962 8925 5009
rect 8959 4962 8965 5009
rect 8919 4941 8965 4962
rect 8919 4890 8925 4941
rect 8959 4890 8965 4941
rect 8919 4873 8965 4890
rect 8919 4818 8925 4873
rect 8959 4818 8965 4873
rect 8919 4805 8965 4818
rect 8919 4746 8925 4805
rect 8959 4746 8965 4805
rect 8919 4737 8965 4746
rect 8919 4674 8925 4737
rect 8959 4674 8965 4737
rect 8919 4669 8965 4674
rect 8919 4602 8925 4669
rect 8959 4602 8965 4669
rect 8919 4601 8965 4602
rect 8919 4567 8925 4601
rect 8959 4567 8965 4601
rect 8919 4564 8965 4567
rect 8919 4499 8925 4564
rect 8959 4499 8965 4564
rect 8919 4492 8965 4499
rect 8919 4431 8925 4492
rect 8959 4431 8965 4492
rect 8919 4420 8965 4431
rect 8919 4363 8925 4420
rect 8959 4363 8965 4420
rect 8919 4348 8965 4363
rect 8919 4295 8925 4348
rect 8959 4295 8965 4348
rect 8919 4276 8965 4295
rect 8919 4227 8925 4276
rect 8959 4227 8965 4276
rect 8919 4204 8965 4227
rect 8919 4159 8925 4204
rect 8959 4159 8965 4204
rect 8919 4132 8965 4159
rect 8919 4091 8925 4132
rect 8959 4091 8965 4132
rect 8919 4060 8965 4091
rect 8919 4023 8925 4060
rect 8959 4023 8965 4060
rect 8919 3989 8965 4023
rect 8919 3954 8925 3989
rect 8959 3954 8965 3989
rect 8919 3921 8965 3954
rect 8919 3882 8925 3921
rect 8959 3882 8965 3921
rect 8919 3853 8965 3882
rect 8919 3810 8925 3853
rect 8959 3810 8965 3853
rect 8919 3785 8965 3810
rect 8919 3738 8925 3785
rect 8959 3738 8965 3785
rect 8919 3717 8965 3738
rect 8919 3666 8925 3717
rect 8959 3666 8965 3717
rect 8919 3649 8965 3666
rect 8919 3594 8925 3649
rect 8959 3594 8965 3649
rect 8919 3581 8965 3594
rect 8919 3522 8925 3581
rect 8959 3522 8965 3581
rect 8919 3513 8965 3522
rect 8919 3450 8925 3513
rect 8959 3450 8965 3513
rect 8919 3445 8965 3450
rect 8919 3378 8925 3445
rect 8959 3378 8965 3445
rect 8919 3377 8965 3378
rect 8919 3343 8925 3377
rect 8959 3343 8965 3377
rect 8919 3340 8965 3343
rect 8919 3275 8925 3340
rect 8959 3275 8965 3340
rect 8919 3268 8965 3275
rect 8919 3207 8925 3268
rect 8959 3207 8965 3268
rect 8919 3196 8965 3207
rect 8919 3139 8925 3196
rect 8959 3139 8965 3196
rect 8919 3124 8965 3139
rect 8919 3071 8925 3124
rect 8959 3071 8965 3124
rect 8919 3052 8965 3071
rect 8919 3003 8925 3052
rect 8959 3003 8965 3052
rect 8919 2980 8965 3003
rect 8919 2935 8925 2980
rect 8959 2935 8965 2980
rect 8919 2908 8965 2935
rect 8919 2867 8925 2908
rect 8959 2867 8965 2908
rect 8919 2836 8965 2867
rect 8919 2799 8925 2836
rect 8959 2799 8965 2836
rect 8919 2765 8965 2799
rect 8919 2730 8925 2765
rect 8959 2730 8965 2765
rect 8919 2697 8965 2730
rect 8919 2658 8925 2697
rect 8959 2658 8965 2697
rect 8919 2629 8965 2658
rect 8919 2586 8925 2629
rect 8959 2586 8965 2629
rect 8919 2561 8965 2586
rect 8919 2514 8925 2561
rect 8959 2514 8965 2561
rect 8919 2493 8965 2514
rect 8919 2442 8925 2493
rect 8959 2442 8965 2493
rect 8919 2425 8965 2442
rect 8919 2370 8925 2425
rect 8959 2370 8965 2425
rect 8919 2357 8965 2370
rect 8919 2298 8925 2357
rect 8959 2298 8965 2357
rect 8919 2289 8965 2298
rect 8919 2226 8925 2289
rect 8959 2226 8965 2289
rect 8919 2221 8965 2226
rect 8919 2154 8925 2221
rect 8959 2154 8965 2221
rect 8919 2153 8965 2154
rect 8919 2119 8925 2153
rect 8959 2119 8965 2153
rect 8919 2116 8965 2119
rect 2196 2042 4116 2076
rect 2196 2025 2230 2042
rect 2196 1991 2208 2025
rect 3964 2008 3998 2042
rect 4032 2025 4116 2042
rect 3964 1991 4000 2008
rect 4034 1991 4074 2025
rect 4108 2008 4116 2025
rect 2196 1953 2230 1991
rect 3964 1974 4082 1991
rect 3964 1953 4014 1974
rect 4048 1953 4116 1974
rect 2196 1919 2208 1953
rect 3964 1940 4000 1953
rect 4048 1940 4074 1953
rect 4108 1940 4116 1953
rect 3896 1919 3926 1940
rect 3960 1919 4000 1940
rect 4034 1919 4074 1940
rect 2196 1872 2230 1919
rect 3896 1906 4082 1919
rect 3896 1872 4116 1906
rect 3945 1848 4116 1872
rect 3979 1814 4116 1848
rect 3945 1806 4116 1814
rect 3945 1780 4042 1806
rect 3979 1772 4042 1780
rect 4076 1772 4116 1806
rect 8919 2051 8925 2116
rect 8959 2051 8965 2116
rect 8919 2044 8965 2051
rect 8919 1983 8925 2044
rect 8959 1983 8965 2044
rect 8919 1972 8965 1983
rect 8919 1915 8925 1972
rect 8959 1915 8965 1972
rect 8919 1900 8965 1915
rect 8919 1847 8925 1900
rect 8959 1847 8965 1900
rect 8919 1828 8965 1847
rect 8919 1782 8925 1828
rect 3979 1746 4116 1772
rect 3945 1738 4116 1746
rect 2269 1685 2303 1719
rect 2337 1685 2371 1719
rect 2406 1685 2439 1719
rect 2479 1685 2507 1719
rect 2552 1685 2575 1719
rect 2625 1685 2643 1719
rect 2698 1685 2711 1719
rect 2771 1685 2779 1719
rect 2844 1685 2847 1719
rect 2881 1685 2883 1719
rect 2917 1685 2956 1719
rect 2990 1685 3000 1719
rect 3063 1685 3068 1719
rect 3170 1685 3175 1719
rect 3238 1685 3248 1719
rect 3306 1685 3321 1719
rect 3374 1685 3394 1719
rect 3442 1685 3467 1719
rect 3510 1685 3540 1719
rect 3578 1685 3612 1719
rect 3647 1685 3680 1719
rect 3720 1685 3759 1719
rect 2508 1637 3476 1648
rect 2307 1603 2326 1637
rect 2360 1603 2402 1637
rect 2436 1603 2452 1637
rect 2508 1603 2524 1637
rect 2558 1603 2658 1637
rect 2692 1603 2780 1637
rect 2814 1603 2914 1637
rect 2948 1603 3036 1637
rect 3070 1603 3170 1637
rect 3204 1603 3292 1637
rect 3326 1603 3426 1637
rect 3460 1603 3476 1637
rect 3532 1603 3548 1637
rect 3582 1603 3624 1637
rect 3658 1603 3674 1637
rect 3759 1617 3793 1651
rect 2307 1511 2341 1603
rect 2508 1592 3476 1603
rect 2719 1511 2753 1592
rect 3231 1511 3265 1592
rect 3563 1563 3597 1603
rect 3563 1491 3597 1529
rect 2304 1419 2307 1453
rect 2341 1419 2344 1453
rect 2304 1381 2344 1419
rect 2304 1347 2307 1381
rect 2341 1347 2344 1381
rect 2304 1309 2344 1347
rect 2304 1275 2307 1309
rect 2341 1275 2344 1309
rect 2304 1236 2344 1275
rect 2304 1202 2307 1236
rect 2341 1202 2344 1236
rect 2304 1163 2344 1202
rect 2304 1129 2307 1163
rect 2341 1129 2344 1163
rect 2304 1090 2344 1129
rect 2304 1056 2307 1090
rect 2341 1056 2344 1090
rect 2304 1017 2344 1056
rect 2304 983 2307 1017
rect 2341 983 2344 1017
rect 2304 944 2344 983
rect 2304 910 2307 944
rect 2341 910 2344 944
rect 2304 871 2344 910
rect 2304 837 2307 871
rect 2341 837 2344 871
rect 2304 798 2344 837
rect 2304 764 2307 798
rect 2341 764 2344 798
rect 2304 725 2344 764
rect 2304 691 2307 725
rect 2341 691 2344 725
rect 2460 1419 2463 1453
rect 2497 1419 2500 1453
rect 2460 1381 2500 1419
rect 2460 1347 2463 1381
rect 2497 1347 2500 1381
rect 2460 1309 2500 1347
rect 2460 1275 2463 1309
rect 2497 1275 2500 1309
rect 2460 1236 2500 1275
rect 2460 1202 2463 1236
rect 2497 1202 2500 1236
rect 2460 1163 2500 1202
rect 2460 1129 2463 1163
rect 2497 1129 2500 1163
rect 2460 1090 2500 1129
rect 2460 1056 2463 1090
rect 2497 1056 2500 1090
rect 2460 1017 2500 1056
rect 2460 983 2463 1017
rect 2497 983 2500 1017
rect 2460 944 2500 983
rect 2460 910 2463 944
rect 2497 910 2500 944
rect 2460 871 2500 910
rect 2460 837 2463 871
rect 2497 837 2500 871
rect 2460 798 2500 837
rect 2460 764 2463 798
rect 2497 764 2500 798
rect 2460 725 2500 764
rect 2460 691 2463 725
rect 2497 691 2500 725
rect 2716 1431 2719 1465
rect 2753 1431 2756 1465
rect 2716 1393 2756 1431
rect 2716 1359 2719 1393
rect 2753 1359 2756 1393
rect 2716 1321 2756 1359
rect 2716 1287 2719 1321
rect 2753 1287 2756 1321
rect 2716 1248 2756 1287
rect 2716 1214 2719 1248
rect 2753 1214 2756 1248
rect 2716 1175 2756 1214
rect 2716 1141 2719 1175
rect 2753 1141 2756 1175
rect 2716 1102 2756 1141
rect 2716 1068 2719 1102
rect 2753 1068 2756 1102
rect 2716 1029 2756 1068
rect 2716 995 2719 1029
rect 2753 995 2756 1029
rect 2716 956 2756 995
rect 2716 922 2719 956
rect 2753 922 2756 956
rect 2716 883 2756 922
rect 2716 849 2719 883
rect 2753 849 2756 883
rect 2716 810 2756 849
rect 2716 776 2719 810
rect 2753 776 2756 810
rect 2716 737 2756 776
rect 2716 703 2719 737
rect 2753 703 2756 737
rect 2972 1419 2975 1453
rect 3009 1419 3012 1453
rect 2972 1381 3012 1419
rect 2972 1347 2975 1381
rect 3009 1347 3012 1381
rect 2972 1309 3012 1347
rect 2972 1275 2975 1309
rect 3009 1275 3012 1309
rect 2972 1236 3012 1275
rect 2972 1202 2975 1236
rect 3009 1202 3012 1236
rect 2972 1163 3012 1202
rect 2972 1129 2975 1163
rect 3009 1129 3012 1163
rect 2972 1090 3012 1129
rect 2972 1056 2975 1090
rect 3009 1056 3012 1090
rect 2972 1017 3012 1056
rect 2972 983 2975 1017
rect 3009 983 3012 1017
rect 2972 944 3012 983
rect 2972 910 2975 944
rect 3009 910 3012 944
rect 2972 871 3012 910
rect 2972 837 2975 871
rect 3009 837 3012 871
rect 2972 798 3012 837
rect 2972 764 2975 798
rect 3009 764 3012 798
rect 2972 725 3012 764
rect 2972 691 2975 725
rect 3009 691 3012 725
rect 3228 1431 3231 1465
rect 3265 1431 3268 1465
rect 3759 1549 3793 1583
rect 3759 1481 3793 1515
rect 3228 1393 3268 1431
rect 3759 1413 3793 1447
rect 3945 1712 4042 1738
rect 3979 1704 4042 1712
rect 4076 1704 4116 1738
rect 3979 1678 4116 1704
rect 3945 1670 4116 1678
rect 3945 1644 4042 1670
rect 3979 1636 4042 1644
rect 4076 1636 4116 1670
rect 3979 1610 4116 1636
rect 3945 1602 4116 1610
rect 3945 1576 4042 1602
rect 3979 1568 4042 1576
rect 4076 1568 4116 1602
rect 3979 1542 4116 1568
rect 3945 1534 4116 1542
rect 3945 1508 4042 1534
rect 3979 1500 4042 1508
rect 4076 1500 4116 1534
rect 3979 1474 4116 1500
rect 3945 1466 4116 1474
rect 3945 1440 4042 1466
rect 3228 1359 3231 1393
rect 3265 1359 3268 1393
rect 3228 1321 3268 1359
rect 3640 1377 3643 1411
rect 3677 1377 3680 1411
rect 3640 1337 3680 1377
rect 3228 1287 3231 1321
rect 3265 1287 3268 1321
rect 3228 1248 3268 1287
rect 3228 1214 3231 1248
rect 3265 1214 3268 1248
rect 3228 1175 3268 1214
rect 3228 1141 3231 1175
rect 3265 1141 3268 1175
rect 3228 1102 3268 1141
rect 3228 1068 3231 1102
rect 3265 1068 3268 1102
rect 3228 1029 3268 1068
rect 3228 995 3231 1029
rect 3265 995 3268 1029
rect 3228 956 3268 995
rect 3228 922 3231 956
rect 3265 922 3268 956
rect 3228 883 3268 922
rect 3228 849 3231 883
rect 3265 849 3268 883
rect 3228 810 3268 849
rect 3228 776 3231 810
rect 3265 776 3268 810
rect 3228 737 3268 776
rect 3228 703 3231 737
rect 3265 703 3268 737
rect 3480 1297 3483 1331
rect 3517 1297 3520 1331
rect 3480 1256 3520 1297
rect 3480 1222 3483 1256
rect 3517 1222 3520 1256
rect 3480 1181 3520 1222
rect 3480 1147 3483 1181
rect 3517 1147 3520 1181
rect 3480 1105 3520 1147
rect 3480 1071 3483 1105
rect 3517 1071 3520 1105
rect 3480 1029 3520 1071
rect 3480 995 3483 1029
rect 3517 995 3520 1029
rect 3480 953 3520 995
rect 3480 919 3483 953
rect 3517 919 3520 953
rect 3480 877 3520 919
rect 3480 843 3483 877
rect 3517 843 3520 877
rect 3480 801 3520 843
rect 3480 767 3483 801
rect 3517 767 3520 801
rect 3480 725 3520 767
rect 3480 691 3483 725
rect 3517 691 3520 725
rect 3640 1303 3643 1337
rect 3677 1303 3680 1337
rect 3640 1262 3680 1303
rect 3640 1228 3643 1262
rect 3677 1228 3680 1262
rect 3640 1187 3680 1228
rect 3640 1153 3643 1187
rect 3677 1153 3680 1187
rect 3640 1112 3680 1153
rect 3640 1078 3643 1112
rect 3677 1078 3680 1112
rect 3640 1037 3680 1078
rect 3640 1003 3643 1037
rect 3677 1003 3680 1037
rect 3640 962 3680 1003
rect 3640 928 3643 962
rect 3677 928 3680 962
rect 3640 887 3680 928
rect 3640 853 3643 887
rect 3677 853 3680 887
rect 3640 812 3680 853
rect 3640 778 3643 812
rect 3677 778 3680 812
rect 3640 737 3680 778
rect 3640 703 3643 737
rect 3677 703 3680 737
rect 3756 1377 3759 1411
rect 3793 1377 3796 1411
rect 3756 1345 3796 1377
rect 3756 1303 3759 1345
rect 3793 1303 3796 1345
rect 3756 1277 3796 1303
rect 3756 1228 3759 1277
rect 3793 1228 3796 1277
rect 3756 1209 3796 1228
rect 3756 1153 3759 1209
rect 3793 1153 3796 1209
rect 3756 1141 3796 1153
rect 3756 1078 3759 1141
rect 3793 1078 3796 1141
rect 3756 1073 3796 1078
rect 3756 1039 3759 1073
rect 3793 1039 3796 1073
rect 3756 1037 3796 1039
rect 3756 971 3759 1037
rect 3793 971 3796 1037
rect 3756 962 3796 971
rect 3756 903 3759 962
rect 3793 903 3796 962
rect 3756 887 3796 903
rect 3756 835 3759 887
rect 3793 835 3796 887
rect 3756 812 3796 835
rect 3756 767 3759 812
rect 3793 767 3796 812
rect 3756 737 3796 767
rect 3756 703 3759 737
rect 3793 703 3796 737
rect 3979 1432 4042 1440
rect 4076 1432 4116 1466
rect 3979 1406 4116 1432
rect 3945 1399 4116 1406
rect 3945 1372 3986 1399
rect 3979 1365 3986 1372
rect 4020 1398 4058 1399
rect 4020 1365 4042 1398
rect 4092 1365 4116 1399
rect 3979 1364 4042 1365
rect 4076 1364 4116 1365
rect 3979 1338 4116 1364
rect 8959 1782 8965 1828
rect 10765 12503 10811 12523
rect 10765 12455 10771 12503
rect 10805 12455 10811 12503
rect 10765 12431 10811 12455
rect 10765 12387 10771 12431
rect 10805 12387 10811 12431
rect 10765 12359 10811 12387
rect 10765 12319 10771 12359
rect 10805 12319 10811 12359
rect 10765 12287 10811 12319
rect 10765 12251 10771 12287
rect 10805 12251 10811 12287
rect 10765 12217 10811 12251
rect 10765 12181 10771 12217
rect 10805 12181 10811 12217
rect 10765 12149 10811 12181
rect 10765 12109 10771 12149
rect 10805 12109 10811 12149
rect 10765 12081 10811 12109
rect 10765 12037 10771 12081
rect 10805 12037 10811 12081
rect 10765 12013 10811 12037
rect 10765 11965 10771 12013
rect 10805 11965 10811 12013
rect 10765 11945 10811 11965
rect 10765 11893 10771 11945
rect 10805 11893 10811 11945
rect 10765 11877 10811 11893
rect 10765 11821 10771 11877
rect 10805 11821 10811 11877
rect 10765 11809 10811 11821
rect 10765 11749 10771 11809
rect 10805 11749 10811 11809
rect 10765 11741 10811 11749
rect 10765 11677 10771 11741
rect 10805 11677 10811 11741
rect 10765 11673 10811 11677
rect 10765 11571 10771 11673
rect 10805 11571 10811 11673
rect 10765 11567 10811 11571
rect 10765 11503 10771 11567
rect 10805 11503 10811 11567
rect 10765 11495 10811 11503
rect 10765 11435 10771 11495
rect 10805 11435 10811 11495
rect 10765 11423 10811 11435
rect 10765 11367 10771 11423
rect 10805 11367 10811 11423
rect 10765 11351 10811 11367
rect 10765 11299 10771 11351
rect 10805 11299 10811 11351
rect 10765 11279 10811 11299
rect 10765 11231 10771 11279
rect 10805 11231 10811 11279
rect 10765 11207 10811 11231
rect 10765 11163 10771 11207
rect 10805 11163 10811 11207
rect 10765 11135 10811 11163
rect 10765 11095 10771 11135
rect 10805 11095 10811 11135
rect 10765 11063 10811 11095
rect 10765 11027 10771 11063
rect 10805 11027 10811 11063
rect 10765 10993 10811 11027
rect 10765 10957 10771 10993
rect 10805 10957 10811 10993
rect 10765 10925 10811 10957
rect 10765 10885 10771 10925
rect 10805 10885 10811 10925
rect 10765 10857 10811 10885
rect 10765 10813 10771 10857
rect 10805 10813 10811 10857
rect 10765 10789 10811 10813
rect 10765 10741 10771 10789
rect 10805 10741 10811 10789
rect 10765 10721 10811 10741
rect 10765 10669 10771 10721
rect 10805 10669 10811 10721
rect 10765 10653 10811 10669
rect 10765 10597 10771 10653
rect 10805 10597 10811 10653
rect 10765 10585 10811 10597
rect 10765 10525 10771 10585
rect 10805 10525 10811 10585
rect 10765 10517 10811 10525
rect 10765 10453 10771 10517
rect 10805 10453 10811 10517
rect 10765 10449 10811 10453
rect 10765 10347 10771 10449
rect 10805 10347 10811 10449
rect 10765 10343 10811 10347
rect 10765 10279 10771 10343
rect 10805 10279 10811 10343
rect 10765 10271 10811 10279
rect 10765 10211 10771 10271
rect 10805 10211 10811 10271
rect 10765 10199 10811 10211
rect 10765 10143 10771 10199
rect 10805 10143 10811 10199
rect 10765 10127 10811 10143
rect 10765 10075 10771 10127
rect 10805 10075 10811 10127
rect 10765 10055 10811 10075
rect 10765 10007 10771 10055
rect 10805 10007 10811 10055
rect 10765 9983 10811 10007
rect 10765 9939 10771 9983
rect 10805 9939 10811 9983
rect 10765 9911 10811 9939
rect 10765 9871 10771 9911
rect 10805 9871 10811 9911
rect 10765 9839 10811 9871
rect 10765 9803 10771 9839
rect 10805 9803 10811 9839
rect 10765 9769 10811 9803
rect 10765 9733 10771 9769
rect 10805 9733 10811 9769
rect 10765 9701 10811 9733
rect 10765 9661 10771 9701
rect 10805 9661 10811 9701
rect 10765 9633 10811 9661
rect 10765 9589 10771 9633
rect 10805 9589 10811 9633
rect 10765 9565 10811 9589
rect 10765 9517 10771 9565
rect 10805 9517 10811 9565
rect 10765 9497 10811 9517
rect 10765 9445 10771 9497
rect 10805 9445 10811 9497
rect 10765 9429 10811 9445
rect 10765 9373 10771 9429
rect 10805 9373 10811 9429
rect 10765 9361 10811 9373
rect 10765 9301 10771 9361
rect 10805 9301 10811 9361
rect 10765 9293 10811 9301
rect 10765 9229 10771 9293
rect 10805 9229 10811 9293
rect 10765 9225 10811 9229
rect 10765 9123 10771 9225
rect 10805 9123 10811 9225
rect 10765 9119 10811 9123
rect 10765 9055 10771 9119
rect 10805 9055 10811 9119
rect 10765 9047 10811 9055
rect 10765 8987 10771 9047
rect 10805 8987 10811 9047
rect 10765 8975 10811 8987
rect 10765 8919 10771 8975
rect 10805 8919 10811 8975
rect 10765 8903 10811 8919
rect 10765 8851 10771 8903
rect 10805 8851 10811 8903
rect 10765 8831 10811 8851
rect 10765 8783 10771 8831
rect 10805 8783 10811 8831
rect 10765 8759 10811 8783
rect 10765 8715 10771 8759
rect 10805 8715 10811 8759
rect 10765 8687 10811 8715
rect 10765 8647 10771 8687
rect 10805 8647 10811 8687
rect 10765 8615 10811 8647
rect 10765 8579 10771 8615
rect 10805 8579 10811 8615
rect 10765 8545 10811 8579
rect 10765 8509 10771 8545
rect 10805 8509 10811 8545
rect 10765 8477 10811 8509
rect 10765 8437 10771 8477
rect 10805 8437 10811 8477
rect 10765 8409 10811 8437
rect 10765 8365 10771 8409
rect 10805 8365 10811 8409
rect 10765 8341 10811 8365
rect 10765 8293 10771 8341
rect 10805 8293 10811 8341
rect 10765 8273 10811 8293
rect 10765 8221 10771 8273
rect 10805 8221 10811 8273
rect 10765 8205 10811 8221
rect 10765 8149 10771 8205
rect 10805 8149 10811 8205
rect 10765 8137 10811 8149
rect 10765 8077 10771 8137
rect 10805 8077 10811 8137
rect 10765 8069 10811 8077
rect 10765 8005 10771 8069
rect 10805 8005 10811 8069
rect 10765 8001 10811 8005
rect 10765 7899 10771 8001
rect 10805 7899 10811 8001
rect 10765 7895 10811 7899
rect 10765 7831 10771 7895
rect 10805 7831 10811 7895
rect 10765 7823 10811 7831
rect 10765 7763 10771 7823
rect 10805 7763 10811 7823
rect 10765 7751 10811 7763
rect 10765 7695 10771 7751
rect 10805 7695 10811 7751
rect 10765 7679 10811 7695
rect 10765 7627 10771 7679
rect 10805 7627 10811 7679
rect 10765 7607 10811 7627
rect 10765 7559 10771 7607
rect 10805 7559 10811 7607
rect 10765 7535 10811 7559
rect 10765 7491 10771 7535
rect 10805 7491 10811 7535
rect 10765 7463 10811 7491
rect 10765 7423 10771 7463
rect 10805 7423 10811 7463
rect 10765 7391 10811 7423
rect 10765 7355 10771 7391
rect 10805 7355 10811 7391
rect 10765 7321 10811 7355
rect 10765 7285 10771 7321
rect 10805 7285 10811 7321
rect 10765 7253 10811 7285
rect 10765 7213 10771 7253
rect 10805 7213 10811 7253
rect 10765 7185 10811 7213
rect 10765 7141 10771 7185
rect 10805 7141 10811 7185
rect 10765 7117 10811 7141
rect 10765 7069 10771 7117
rect 10805 7069 10811 7117
rect 10765 7049 10811 7069
rect 10765 6997 10771 7049
rect 10805 6997 10811 7049
rect 10765 6981 10811 6997
rect 10765 6925 10771 6981
rect 10805 6925 10811 6981
rect 10765 6913 10811 6925
rect 10765 6853 10771 6913
rect 10805 6853 10811 6913
rect 10765 6845 10811 6853
rect 10765 6781 10771 6845
rect 10805 6781 10811 6845
rect 10765 6777 10811 6781
rect 10765 6675 10771 6777
rect 10805 6675 10811 6777
rect 10765 6671 10811 6675
rect 10765 6607 10771 6671
rect 10805 6607 10811 6671
rect 10765 6599 10811 6607
rect 10765 6539 10771 6599
rect 10805 6539 10811 6599
rect 10765 6527 10811 6539
rect 10765 6471 10771 6527
rect 10805 6471 10811 6527
rect 10765 6455 10811 6471
rect 10765 6403 10771 6455
rect 10805 6403 10811 6455
rect 10765 6383 10811 6403
rect 10765 6335 10771 6383
rect 10805 6335 10811 6383
rect 10765 6311 10811 6335
rect 10765 6267 10771 6311
rect 10805 6267 10811 6311
rect 10765 6239 10811 6267
rect 10765 6199 10771 6239
rect 10805 6199 10811 6239
rect 10765 6167 10811 6199
rect 10765 6131 10771 6167
rect 10805 6131 10811 6167
rect 10765 6097 10811 6131
rect 10765 6061 10771 6097
rect 10805 6061 10811 6097
rect 10765 6029 10811 6061
rect 10765 5989 10771 6029
rect 10805 5989 10811 6029
rect 10765 5961 10811 5989
rect 10765 5917 10771 5961
rect 10805 5917 10811 5961
rect 10765 5893 10811 5917
rect 10765 5845 10771 5893
rect 10805 5845 10811 5893
rect 10765 5825 10811 5845
rect 10765 5773 10771 5825
rect 10805 5773 10811 5825
rect 10765 5757 10811 5773
rect 10765 5701 10771 5757
rect 10805 5701 10811 5757
rect 10765 5689 10811 5701
rect 10765 5629 10771 5689
rect 10805 5629 10811 5689
rect 10765 5621 10811 5629
rect 10765 5557 10771 5621
rect 10805 5557 10811 5621
rect 10765 5553 10811 5557
rect 10765 5451 10771 5553
rect 10805 5451 10811 5553
rect 10765 5447 10811 5451
rect 10765 5383 10771 5447
rect 10805 5383 10811 5447
rect 10765 5375 10811 5383
rect 10765 5315 10771 5375
rect 10805 5315 10811 5375
rect 10765 5303 10811 5315
rect 10765 5247 10771 5303
rect 10805 5247 10811 5303
rect 10765 5231 10811 5247
rect 10765 5179 10771 5231
rect 10805 5179 10811 5231
rect 10765 5159 10811 5179
rect 10765 5111 10771 5159
rect 10805 5111 10811 5159
rect 10765 5087 10811 5111
rect 10765 5043 10771 5087
rect 10805 5043 10811 5087
rect 10765 5015 10811 5043
rect 10765 4975 10771 5015
rect 10805 4975 10811 5015
rect 10765 4943 10811 4975
rect 10765 4907 10771 4943
rect 10805 4907 10811 4943
rect 10765 4873 10811 4907
rect 10765 4837 10771 4873
rect 10805 4837 10811 4873
rect 10765 4805 10811 4837
rect 10765 4765 10771 4805
rect 10805 4765 10811 4805
rect 10765 4737 10811 4765
rect 10765 4693 10771 4737
rect 10805 4693 10811 4737
rect 10765 4669 10811 4693
rect 10765 4621 10771 4669
rect 10805 4621 10811 4669
rect 10765 4601 10811 4621
rect 10765 4549 10771 4601
rect 10805 4549 10811 4601
rect 10765 4533 10811 4549
rect 10765 4477 10771 4533
rect 10805 4477 10811 4533
rect 10765 4465 10811 4477
rect 10765 4405 10771 4465
rect 10805 4405 10811 4465
rect 10765 4397 10811 4405
rect 10765 4333 10771 4397
rect 10805 4333 10811 4397
rect 10765 4329 10811 4333
rect 10765 4227 10771 4329
rect 10805 4227 10811 4329
rect 10765 4223 10811 4227
rect 10765 4159 10771 4223
rect 10805 4159 10811 4223
rect 10765 4151 10811 4159
rect 10765 4091 10771 4151
rect 10805 4091 10811 4151
rect 10765 4079 10811 4091
rect 10765 4023 10771 4079
rect 10805 4023 10811 4079
rect 10765 4007 10811 4023
rect 10765 3955 10771 4007
rect 10805 3955 10811 4007
rect 10765 3935 10811 3955
rect 10765 3887 10771 3935
rect 10805 3887 10811 3935
rect 10765 3863 10811 3887
rect 10765 3819 10771 3863
rect 10805 3819 10811 3863
rect 10765 3791 10811 3819
rect 10765 3751 10771 3791
rect 10805 3751 10811 3791
rect 10765 3719 10811 3751
rect 10765 3683 10771 3719
rect 10805 3683 10811 3719
rect 10765 3649 10811 3683
rect 10765 3613 10771 3649
rect 10805 3613 10811 3649
rect 10765 3581 10811 3613
rect 10765 3541 10771 3581
rect 10805 3541 10811 3581
rect 10765 3513 10811 3541
rect 10765 3469 10771 3513
rect 10805 3469 10811 3513
rect 10765 3445 10811 3469
rect 10765 3397 10771 3445
rect 10805 3397 10811 3445
rect 10765 3377 10811 3397
rect 10765 3325 10771 3377
rect 10805 3325 10811 3377
rect 10765 3309 10811 3325
rect 10765 3253 10771 3309
rect 10805 3253 10811 3309
rect 10765 3241 10811 3253
rect 10765 3181 10771 3241
rect 10805 3181 10811 3241
rect 10765 3173 10811 3181
rect 10765 3109 10771 3173
rect 10805 3109 10811 3173
rect 10765 3105 10811 3109
rect 10765 3003 10771 3105
rect 10805 3003 10811 3105
rect 10765 2999 10811 3003
rect 10765 2935 10771 2999
rect 10805 2935 10811 2999
rect 10765 2927 10811 2935
rect 10765 2867 10771 2927
rect 10805 2867 10811 2927
rect 10765 2855 10811 2867
rect 10765 2799 10771 2855
rect 10805 2799 10811 2855
rect 10765 2783 10811 2799
rect 10765 2731 10771 2783
rect 10805 2731 10811 2783
rect 10765 2711 10811 2731
rect 10765 2663 10771 2711
rect 10805 2663 10811 2711
rect 10765 2639 10811 2663
rect 10765 2595 10771 2639
rect 10805 2595 10811 2639
rect 10765 2567 10811 2595
rect 10765 2527 10771 2567
rect 10805 2527 10811 2567
rect 10765 2495 10811 2527
rect 10765 2459 10771 2495
rect 10805 2459 10811 2495
rect 10765 2425 10811 2459
rect 10765 2389 10771 2425
rect 10805 2389 10811 2425
rect 10765 2357 10811 2389
rect 10765 2317 10771 2357
rect 10805 2317 10811 2357
rect 10765 2289 10811 2317
rect 10765 2245 10771 2289
rect 10805 2245 10811 2289
rect 10765 2221 10811 2245
rect 10765 2173 10771 2221
rect 10805 2173 10811 2221
rect 10765 2153 10811 2173
rect 10765 2101 10771 2153
rect 10805 2101 10811 2153
rect 10765 2085 10811 2101
rect 10765 2029 10771 2085
rect 10805 2029 10811 2085
rect 10765 2017 10811 2029
rect 10765 1957 10771 2017
rect 10805 1957 10811 2017
rect 10765 1949 10811 1957
rect 10765 1885 10771 1949
rect 10805 1885 10811 1949
rect 10765 1881 10811 1885
rect 8925 1745 8959 1779
rect 8925 1677 8959 1711
rect 8925 1609 8959 1643
rect 8925 1541 8959 1575
rect 8925 1473 8959 1507
rect 8925 1405 8959 1439
rect 3945 1330 4116 1338
rect 3945 1324 4042 1330
rect 4076 1324 4116 1330
rect 3945 1304 3986 1324
rect 3979 1290 3986 1304
rect 4020 1296 4042 1324
rect 4020 1290 4058 1296
rect 4092 1290 4116 1324
rect 3979 1270 4116 1290
rect 3945 1262 4116 1270
rect 3945 1249 4042 1262
rect 4076 1249 4116 1262
rect 3945 1236 3986 1249
rect 3979 1215 3986 1236
rect 4020 1228 4042 1249
rect 4020 1215 4058 1228
rect 4092 1215 4116 1249
rect 3979 1202 4116 1215
rect 3945 1194 4116 1202
rect 3945 1174 4042 1194
rect 4076 1174 4116 1194
rect 3945 1167 3986 1174
rect 3979 1140 3986 1167
rect 4020 1160 4042 1174
rect 4020 1140 4058 1160
rect 4092 1140 4116 1174
rect 3979 1133 4116 1140
rect 3945 1126 4116 1133
rect 3945 1099 4042 1126
rect 4076 1099 4116 1126
rect 3945 1098 3986 1099
rect 3979 1065 3986 1098
rect 4020 1092 4042 1099
rect 4020 1065 4058 1092
rect 4092 1065 4116 1099
rect 3979 1064 4116 1065
rect 3945 1058 4116 1064
rect 3945 1029 4042 1058
rect 3979 1024 4042 1029
rect 4076 1024 4116 1058
rect 3979 995 3986 1024
rect 3945 990 3986 995
rect 4020 990 4058 1024
rect 4092 990 4116 1024
rect 3945 960 4042 990
rect 3979 956 4042 960
rect 4076 956 4116 990
rect 3979 949 4116 956
rect 3979 926 3986 949
rect 3945 915 3986 926
rect 4020 922 4058 949
rect 4020 915 4042 922
rect 4092 915 4116 949
rect 3945 891 4042 915
rect 3979 888 4042 891
rect 4076 888 4116 915
rect 3979 874 4116 888
rect 3979 857 3986 874
rect 3945 840 3986 857
rect 4020 854 4058 874
rect 4020 840 4042 854
rect 4092 840 4116 874
rect 3945 822 4042 840
rect 3979 820 4042 822
rect 4076 820 4116 840
rect 3979 799 4116 820
rect 3979 788 3986 799
rect 3945 765 3986 788
rect 4020 786 4058 799
rect 4020 765 4042 786
rect 4092 765 4116 799
rect 3945 753 4042 765
rect 3979 752 4042 753
rect 4076 752 4116 765
rect 3979 724 4116 752
rect 3979 719 3986 724
rect 3759 665 3793 699
rect 3759 597 3793 631
rect 3759 491 3793 563
rect 2269 457 2365 491
rect 2406 457 2433 491
rect 2479 457 2501 491
rect 2552 457 2569 491
rect 2625 457 2637 491
rect 2698 457 2705 491
rect 2771 457 2773 491
rect 2807 457 2810 491
rect 2875 457 2882 491
rect 2943 457 2954 491
rect 3011 457 3026 491
rect 3079 457 3098 491
rect 3147 457 3170 491
rect 3215 457 3242 491
rect 3283 457 3314 491
rect 3351 457 3385 491
rect 3420 457 3453 491
rect 3492 457 3521 491
rect 3564 457 3589 491
rect 3636 457 3657 491
rect 3708 457 3725 491
rect 3780 457 3793 491
rect 3945 690 3986 719
rect 4020 718 4058 724
rect 4020 690 4042 718
rect 4092 690 4116 724
rect 3945 684 4042 690
rect 4076 684 4116 690
rect 3979 650 4116 684
rect 3945 649 4042 650
rect 4076 649 4116 650
rect 3945 615 3986 649
rect 4020 616 4042 649
rect 4020 615 4058 616
rect 4092 615 4116 649
rect 3979 582 4116 615
rect 3979 581 4042 582
rect 3945 574 4042 581
rect 4076 574 4116 582
rect 3945 546 3986 574
rect 3979 540 3986 546
rect 4020 548 4042 574
rect 4020 540 4058 548
rect 4092 540 4116 574
rect 3979 514 4116 540
rect 3979 512 4042 514
rect 3945 500 4042 512
rect 4076 500 4116 514
rect 3945 477 3986 500
rect 3979 466 3986 477
rect 4020 480 4042 500
rect 4020 466 4058 480
rect 4092 466 4116 500
rect 3979 446 4116 466
rect 3979 443 4042 446
rect 3945 426 4042 443
rect 4076 426 4116 446
rect 3945 408 3986 426
rect 3979 392 3986 408
rect 4020 412 4042 426
rect 4020 392 4058 412
rect 4092 392 4116 426
rect 3979 378 4116 392
rect 3979 374 4042 378
rect 3945 352 4042 374
rect 4076 352 4116 378
rect 3945 339 3986 352
rect 3979 318 3986 339
rect 4020 344 4042 352
rect 4020 318 4058 344
rect 4092 318 4116 352
rect 3979 310 4116 318
rect 3979 305 4042 310
rect 2214 280 2238 305
rect 2272 280 2308 305
rect 2342 280 2378 305
rect 2412 280 2448 305
rect 2214 246 2226 280
rect 2272 271 2300 280
rect 2342 271 2373 280
rect 2412 271 2446 280
rect 2482 271 2518 305
rect 2552 280 2588 305
rect 2622 280 2658 305
rect 2692 280 2728 305
rect 2762 280 2798 305
rect 2832 280 2868 305
rect 2902 280 2938 305
rect 2972 280 3008 305
rect 3042 280 3078 305
rect 3112 280 3148 305
rect 3182 280 3218 305
rect 3252 280 3288 305
rect 2553 271 2588 280
rect 2626 271 2658 280
rect 2699 271 2728 280
rect 2772 271 2798 280
rect 2845 271 2868 280
rect 2918 271 2938 280
rect 2991 271 3008 280
rect 3064 271 3078 280
rect 3137 271 3148 280
rect 3210 271 3218 280
rect 3283 271 3288 280
rect 3322 280 3358 305
rect 2260 246 2300 271
rect 2334 246 2373 271
rect 2407 246 2446 271
rect 2480 246 2519 271
rect 2553 246 2592 271
rect 2626 246 2665 271
rect 2699 246 2738 271
rect 2772 246 2811 271
rect 2845 246 2884 271
rect 2918 246 2957 271
rect 2991 246 3030 271
rect 3064 246 3103 271
rect 3137 246 3176 271
rect 3210 246 3249 271
rect 3283 246 3322 271
rect 3356 271 3358 280
rect 3392 280 3427 305
rect 3461 280 3496 305
rect 3530 280 3565 305
rect 3599 280 3634 305
rect 3668 280 3703 305
rect 3737 280 3772 305
rect 3806 280 3841 305
rect 3875 280 4042 305
rect 4076 280 4116 310
rect 3392 271 3395 280
rect 3461 271 3468 280
rect 3530 271 3541 280
rect 3599 271 3614 280
rect 3668 271 3687 280
rect 3737 271 3760 280
rect 3806 271 3833 280
rect 3875 271 3906 280
rect 3356 246 3395 271
rect 3429 246 3468 271
rect 3502 246 3541 271
rect 3575 246 3614 271
rect 3648 246 3687 271
rect 3721 246 3760 271
rect 3794 246 3833 271
rect 3867 246 3906 271
rect 3940 246 3979 280
rect 4013 276 4042 280
rect 4013 246 4052 276
rect 4086 246 4116 280
rect 2214 242 4116 246
rect 2214 208 4042 242
rect 4076 208 4116 242
rect 2214 174 2226 208
rect 2282 174 2300 208
rect 2350 174 2373 208
rect 2418 174 2446 208
rect 2486 174 2519 208
rect 2554 174 2588 208
rect 2626 174 2656 208
rect 2699 174 2724 208
rect 2772 174 2792 208
rect 2845 174 2860 208
rect 2918 174 2928 208
rect 2991 174 2996 208
rect 3098 174 3103 208
rect 3166 174 3176 208
rect 3234 174 3249 208
rect 3302 174 3322 208
rect 3370 174 3395 208
rect 3438 174 3468 208
rect 3506 174 3540 208
rect 3575 174 3608 208
rect 3648 174 3676 208
rect 3721 174 3744 208
rect 3794 174 3812 208
rect 3867 174 3880 208
rect 3940 174 3948 208
rect 4013 174 4052 208
rect 4086 174 4116 208
rect 7863 1313 7887 1347
rect 7921 1313 7967 1347
rect 8001 1313 8046 1347
rect 8080 1313 8125 1347
rect 8159 1313 8197 1347
rect 8238 1313 8283 1347
rect 8335 1313 8341 1347
rect 7863 1279 7897 1313
rect 8307 1279 8341 1313
rect 7863 1210 7897 1245
rect 7965 1219 8003 1253
rect 8037 1219 8050 1253
rect 8084 1219 8126 1253
rect 8160 1219 8176 1253
rect 7863 1161 7897 1176
rect 8307 1210 8341 1241
rect 7863 1085 7897 1107
rect 7863 1009 7897 1039
rect 7863 937 7897 971
rect 7863 869 7897 899
rect 7863 801 7897 823
rect 7863 733 7897 747
rect 7863 665 7897 671
rect 7863 629 7897 631
rect 7863 553 7897 563
rect 7863 478 7897 495
rect 7863 403 7897 427
rect 7863 328 7897 359
rect 7863 257 7897 291
rect 7863 189 7897 219
rect 7979 1088 8013 1127
rect 7979 1015 8013 1054
rect 8191 1088 8225 1127
rect 8191 1015 8225 1054
rect 7979 942 8013 981
rect 7979 869 8013 908
rect 7979 796 8013 835
rect 7979 723 8013 762
rect 7979 650 8013 689
rect 7979 577 8013 616
rect 7979 505 8013 543
rect 7979 433 8013 471
rect 7979 361 8013 399
rect 7979 289 8013 327
rect 7979 217 8013 255
rect 8085 922 8119 961
rect 8085 849 8119 888
rect 8085 776 8119 815
rect 8085 703 8119 742
rect 8085 631 8119 669
rect 8085 559 8119 597
rect 8085 487 8119 525
rect 8085 415 8119 453
rect 8085 343 8119 381
rect 8085 271 8119 309
rect 8191 942 8225 981
rect 8191 869 8225 908
rect 8191 796 8225 835
rect 8191 723 8225 762
rect 8191 650 8225 689
rect 8191 577 8225 616
rect 8191 505 8225 543
rect 8191 433 8225 471
rect 8191 361 8225 399
rect 8191 289 8225 327
rect 8191 217 8225 255
rect 8307 1141 8341 1167
rect 8307 1073 8341 1093
rect 8307 1005 8341 1019
rect 8307 937 8341 945
rect 8307 869 8341 872
rect 8307 833 8341 835
rect 8307 760 8341 767
rect 8307 687 8341 699
rect 8307 614 8341 631
rect 8307 541 8341 563
rect 8307 468 8341 495
rect 8307 395 8341 427
rect 8307 325 8341 359
rect 8307 257 8341 288
rect 8307 189 8341 215
rect 7863 121 7897 144
rect 8307 121 8341 142
rect 7897 69 7931 97
rect 7863 63 7931 69
rect 7965 63 8005 97
rect 8067 63 8146 97
rect 8199 63 8228 97
rect 8262 69 8307 97
rect 8262 63 8341 69
rect 8925 1337 8959 1371
rect 8925 1269 8959 1303
rect 8925 1201 8959 1235
rect 8925 1133 8959 1167
rect 8925 1065 8959 1099
rect 8925 997 8959 1031
rect 8925 929 8959 963
rect 8925 861 8959 895
rect 8925 793 8959 827
rect 8925 725 8959 759
rect 8925 657 8959 691
rect 8925 589 8959 623
rect 8925 521 8959 555
rect 8925 453 8959 487
rect 8925 385 8959 419
rect 8925 317 8959 351
rect 8925 249 8959 283
rect 8925 181 8959 215
rect 8925 113 8959 147
rect 8925 45 8959 79
rect 8925 -23 8959 11
rect 8925 -91 8959 -57
rect 8925 -159 8959 -125
rect 8925 -227 8959 -193
rect 8925 -295 8959 -261
rect 8925 -363 8959 -329
rect 8925 -431 8959 -397
rect 8925 -499 8959 -465
rect 8925 -567 8959 -533
rect 8925 -635 8959 -601
rect 8925 -703 8959 -669
rect 8925 -771 8959 -737
rect 8925 -839 8959 -805
rect 8925 -907 8959 -873
rect 8925 -975 8959 -941
rect 8925 -1043 8959 -1009
rect 8925 -1111 8959 -1077
rect 8925 -1179 8959 -1145
rect 8925 -1247 8959 -1213
rect 8925 -1315 8959 -1281
rect 8925 -1383 8959 -1349
rect 8925 -1451 8959 -1417
rect 8925 -1519 8959 -1485
rect 10765 1779 10771 1881
rect 10805 1779 10811 1881
rect 10765 1775 10811 1779
rect 10765 1711 10771 1775
rect 10805 1711 10811 1775
rect 10765 1703 10811 1711
rect 10765 1643 10771 1703
rect 10805 1643 10811 1703
rect 10765 1631 10811 1643
rect 10765 1575 10771 1631
rect 10805 1575 10811 1631
rect 10765 1559 10811 1575
rect 10765 1507 10771 1559
rect 10805 1507 10811 1559
rect 10765 1487 10811 1507
rect 10765 1439 10771 1487
rect 10805 1439 10811 1487
rect 10765 1415 10811 1439
rect 10765 1371 10771 1415
rect 10805 1371 10811 1415
rect 10765 1343 10811 1371
rect 10765 1303 10771 1343
rect 10805 1303 10811 1343
rect 10765 1271 10811 1303
rect 10765 1235 10771 1271
rect 10805 1235 10811 1271
rect 10765 1201 10811 1235
rect 10765 1165 10771 1201
rect 10805 1165 10811 1201
rect 10765 1133 10811 1165
rect 10765 1093 10771 1133
rect 10805 1093 10811 1133
rect 10765 1065 10811 1093
rect 10765 1021 10771 1065
rect 10805 1021 10811 1065
rect 10765 997 10811 1021
rect 10765 949 10771 997
rect 10805 949 10811 997
rect 10765 929 10811 949
rect 10765 877 10771 929
rect 10805 877 10811 929
rect 10765 861 10811 877
rect 10765 805 10771 861
rect 10805 805 10811 861
rect 10765 793 10811 805
rect 10765 733 10771 793
rect 10805 733 10811 793
rect 10765 725 10811 733
rect 10765 661 10771 725
rect 10805 661 10811 725
rect 10765 657 10811 661
rect 10765 555 10771 657
rect 10805 555 10811 657
rect 10765 551 10811 555
rect 10765 487 10771 551
rect 10805 487 10811 551
rect 10765 479 10811 487
rect 10765 419 10771 479
rect 10805 419 10811 479
rect 10765 407 10811 419
rect 10765 351 10771 407
rect 10805 351 10811 407
rect 10765 335 10811 351
rect 10765 283 10771 335
rect 10805 283 10811 335
rect 10765 263 10811 283
rect 10765 215 10771 263
rect 10805 215 10811 263
rect 10765 191 10811 215
rect 10765 147 10771 191
rect 10805 147 10811 191
rect 10765 119 10811 147
rect 10765 79 10771 119
rect 10805 79 10811 119
rect 10765 47 10811 79
rect 10765 11 10771 47
rect 10805 11 10811 47
rect 10765 -23 10811 11
rect 10765 -59 10771 -23
rect 10805 -59 10811 -23
rect 10765 -91 10811 -59
rect 10765 -131 10771 -91
rect 10805 -131 10811 -91
rect 10765 -159 10811 -131
rect 10765 -203 10771 -159
rect 10805 -203 10811 -159
rect 10765 -227 10811 -203
rect 10765 -275 10771 -227
rect 10805 -275 10811 -227
rect 10765 -295 10811 -275
rect 10765 -347 10771 -295
rect 10805 -347 10811 -295
rect 10765 -363 10811 -347
rect 10765 -419 10771 -363
rect 10805 -419 10811 -363
rect 10765 -431 10811 -419
rect 10765 -491 10771 -431
rect 10805 -491 10811 -431
rect 10765 -499 10811 -491
rect 10765 -563 10771 -499
rect 10805 -563 10811 -499
rect 10765 -567 10811 -563
rect 10765 -669 10771 -567
rect 10805 -669 10811 -567
rect 10765 -673 10811 -669
rect 10765 -737 10771 -673
rect 10805 -737 10811 -673
rect 10765 -745 10811 -737
rect 10765 -805 10771 -745
rect 10805 -805 10811 -745
rect 10765 -817 10811 -805
rect 10765 -873 10771 -817
rect 10805 -873 10811 -817
rect 10765 -889 10811 -873
rect 10765 -941 10771 -889
rect 10805 -941 10811 -889
rect 10765 -961 10811 -941
rect 10765 -1009 10771 -961
rect 10805 -1009 10811 -961
rect 10765 -1033 10811 -1009
rect 10765 -1077 10771 -1033
rect 10805 -1077 10811 -1033
rect 10765 -1105 10811 -1077
rect 10765 -1145 10771 -1105
rect 10805 -1145 10811 -1105
rect 10765 -1177 10811 -1145
rect 10765 -1213 10771 -1177
rect 10805 -1213 10811 -1177
rect 10765 -1247 10811 -1213
rect 10765 -1283 10771 -1247
rect 10805 -1283 10811 -1247
rect 10765 -1315 10811 -1283
rect 10765 -1355 10771 -1315
rect 10805 -1355 10811 -1315
rect 10765 -1383 10811 -1355
rect 10765 -1427 10771 -1383
rect 10805 -1427 10811 -1383
rect 10765 -1451 10811 -1427
rect 10765 -1499 10771 -1451
rect 10805 -1499 10811 -1451
rect 10765 -1519 10811 -1499
rect 8925 -1587 8959 -1553
rect 8925 -1655 8959 -1621
rect 10431 -1555 10497 -1546
rect 10431 -1589 10446 -1555
rect 10480 -1589 10497 -1555
rect 10431 -1627 10497 -1589
rect 10431 -1661 10446 -1627
rect 10480 -1661 10497 -1627
rect 10431 -1664 10497 -1661
rect 10593 -1556 10676 -1546
rect 10593 -1590 10642 -1556
rect 10593 -1628 10676 -1590
rect 10593 -1662 10642 -1628
rect 10593 -1664 10676 -1662
rect 10765 -1571 10771 -1519
rect 10805 -1571 10811 -1519
rect 10765 -1587 10811 -1571
rect 10765 -1643 10771 -1587
rect 10805 -1643 10811 -1587
rect 10765 -1655 10811 -1643
rect 8925 -1723 8959 -1689
rect 8925 -1791 8959 -1757
rect 8925 -1859 8959 -1825
rect 8925 -1927 8959 -1893
rect 8925 -1995 8959 -1961
rect 8925 -2064 8959 -2029
rect 8925 -2133 8959 -2098
rect 8925 -2202 8959 -2167
rect 8925 -2271 8959 -2236
rect 8925 -2340 8959 -2305
rect 8925 -2409 8959 -2374
rect 8925 -2478 8959 -2443
rect 8925 -2547 8959 -2512
rect 8925 -2616 8959 -2581
rect 8925 -2685 8959 -2650
rect 8925 -2754 8959 -2719
rect 8925 -2823 8959 -2788
rect 8925 -2892 8959 -2857
rect 8925 -2961 8959 -2926
rect 8925 -3030 8959 -2995
rect 10765 -1715 10771 -1655
rect 10805 -1715 10811 -1655
rect 10765 -1723 10811 -1715
rect 10765 -1787 10771 -1723
rect 10805 -1787 10811 -1723
rect 10765 -1791 10811 -1787
rect 10765 -1893 10771 -1791
rect 10805 -1893 10811 -1791
rect 10765 -1897 10811 -1893
rect 10765 -1961 10771 -1897
rect 10805 -1961 10811 -1897
rect 10765 -1969 10811 -1961
rect 10765 -2029 10771 -1969
rect 10805 -2029 10811 -1969
rect 10765 -2041 10811 -2029
rect 10765 -2097 10771 -2041
rect 10805 -2097 10811 -2041
rect 10765 -2113 10811 -2097
rect 10765 -2165 10771 -2113
rect 10805 -2165 10811 -2113
rect 10765 -2185 10811 -2165
rect 10765 -2233 10771 -2185
rect 10805 -2233 10811 -2185
rect 10765 -2257 10811 -2233
rect 10765 -2301 10771 -2257
rect 10805 -2301 10811 -2257
rect 10765 -2329 10811 -2301
rect 10765 -2369 10771 -2329
rect 10805 -2369 10811 -2329
rect 10765 -2401 10811 -2369
rect 10765 -2437 10771 -2401
rect 10805 -2437 10811 -2401
rect 10765 -2471 10811 -2437
rect 10765 -2507 10771 -2471
rect 10805 -2507 10811 -2471
rect 10765 -2539 10811 -2507
rect 10765 -2579 10771 -2539
rect 10805 -2579 10811 -2539
rect 10765 -2607 10811 -2579
rect 10765 -2651 10771 -2607
rect 10805 -2651 10811 -2607
rect 10765 -2675 10811 -2651
rect 10765 -2723 10771 -2675
rect 10805 -2723 10811 -2675
rect 10765 -2743 10811 -2723
rect 10765 -2795 10771 -2743
rect 10805 -2795 10811 -2743
rect 10765 -2811 10811 -2795
rect 10765 -2867 10771 -2811
rect 10805 -2867 10811 -2811
rect 10765 -2879 10811 -2867
rect 10765 -2939 10771 -2879
rect 10805 -2939 10811 -2879
rect 10765 -2947 10811 -2939
rect 10765 -3011 10771 -2947
rect 10805 -3011 10811 -2947
rect 10765 -3015 10811 -3011
rect 8925 -3099 8959 -3064
rect 8925 -3168 8959 -3133
rect 8925 -3237 8959 -3202
rect 8925 -3306 8959 -3271
rect 8925 -3375 8959 -3340
rect 9071 -3093 9087 -3059
rect 9121 -3093 9137 -3059
rect 9071 -3131 9137 -3093
rect 9071 -3165 9087 -3131
rect 9121 -3165 9137 -3131
rect 9071 -3377 9137 -3165
rect 9233 -3143 9277 -3109
rect 9311 -3143 9339 -3109
rect 9233 -3181 9339 -3143
rect 9233 -3215 9277 -3181
rect 9311 -3215 9339 -3181
rect 9233 -3377 9339 -3215
rect 8925 -3444 8959 -3409
rect 8925 -3513 8959 -3478
rect 8925 -3582 8959 -3547
rect 8925 -3651 8959 -3616
rect 8925 -3720 8959 -3685
rect 8925 -3789 8959 -3754
rect 8925 -3858 8959 -3823
rect 9209 -3835 9339 -3377
rect 9209 -3869 9221 -3835
rect 9255 -3869 9293 -3835
rect 9327 -3869 9339 -3835
rect 9209 -3886 9339 -3869
rect 10765 -3117 10771 -3015
rect 10805 -3117 10811 -3015
rect 10765 -3121 10811 -3117
rect 10765 -3185 10771 -3121
rect 10805 -3185 10811 -3121
rect 10765 -3193 10811 -3185
rect 10765 -3253 10771 -3193
rect 10805 -3253 10811 -3193
rect 10765 -3265 10811 -3253
rect 10765 -3321 10771 -3265
rect 10805 -3321 10811 -3265
rect 10765 -3337 10811 -3321
rect 10765 -3389 10771 -3337
rect 10805 -3389 10811 -3337
rect 10765 -3409 10811 -3389
rect 10765 -3458 10771 -3409
rect 10805 -3458 10811 -3409
rect 10765 -3481 10811 -3458
rect 10765 -3527 10771 -3481
rect 10805 -3527 10811 -3481
rect 10765 -3553 10811 -3527
rect 10765 -3596 10771 -3553
rect 10805 -3596 10811 -3553
rect 10765 -3625 10811 -3596
rect 10765 -3665 10771 -3625
rect 10805 -3665 10811 -3625
rect 10765 -3697 10811 -3665
rect 10765 -3734 10771 -3697
rect 10805 -3734 10811 -3697
rect 10765 -3769 10811 -3734
rect 10765 -3803 10771 -3769
rect 10805 -3803 10811 -3769
rect 10765 -3838 10811 -3803
rect 10765 -3875 10771 -3838
rect 10805 -3875 10811 -3838
rect 8925 -3927 8959 -3892
rect 10765 -3907 10811 -3875
rect 8959 -3961 9015 -3945
rect 8925 -3979 9015 -3961
rect 9049 -3979 9085 -3945
rect 9119 -3979 9155 -3945
rect 9189 -3979 9225 -3945
rect 9259 -3979 9295 -3945
rect 9329 -3979 9347 -3945
rect 9313 -4033 9347 -3979
rect 9313 -4102 9347 -4067
rect 9313 -4171 9347 -4136
rect 9313 -4240 9347 -4205
rect 9313 -4309 9347 -4274
rect 9313 -4378 9347 -4343
rect 9313 -4447 9347 -4412
rect 9313 -4516 9347 -4481
rect 9313 -4585 9347 -4550
rect 9313 -4654 9347 -4619
rect 9313 -4723 9347 -4688
rect 9313 -4792 9347 -4757
rect 9313 -4861 9347 -4826
rect 9313 -4930 9347 -4895
rect 9313 -4999 9347 -4964
rect 9313 -5068 9347 -5033
rect 9313 -5137 9347 -5102
rect 9313 -5206 9347 -5171
rect 9313 -5275 9347 -5240
rect 9313 -5344 9347 -5309
rect 9313 -5413 9347 -5378
rect 9313 -5482 9347 -5447
rect 9313 -5551 9347 -5516
rect 9313 -5620 9347 -5585
rect 9313 -5689 9347 -5654
rect 9313 -5759 9347 -5723
rect 9313 -5829 9347 -5793
rect 9313 -5899 9347 -5863
rect 10765 -3947 10771 -3907
rect 10805 -3947 10811 -3907
rect 10765 -3976 10811 -3947
rect 10765 -4019 10771 -3976
rect 10805 -4019 10811 -3976
rect 10765 -4045 10811 -4019
rect 10765 -4091 10771 -4045
rect 10805 -4091 10811 -4045
rect 10765 -4114 10811 -4091
rect 10765 -4163 10771 -4114
rect 10805 -4163 10811 -4114
rect 10765 -4183 10811 -4163
rect 10765 -4235 10771 -4183
rect 10805 -4235 10811 -4183
rect 10765 -4252 10811 -4235
rect 10765 -4307 10771 -4252
rect 10805 -4307 10811 -4252
rect 10765 -4321 10811 -4307
rect 10765 -4379 10771 -4321
rect 10805 -4379 10811 -4321
rect 10765 -4390 10811 -4379
rect 10765 -4451 10771 -4390
rect 10805 -4451 10811 -4390
rect 10765 -4459 10811 -4451
rect 10765 -4523 10771 -4459
rect 10805 -4523 10811 -4459
rect 10765 -4528 10811 -4523
rect 10765 -4595 10771 -4528
rect 10805 -4595 10811 -4528
rect 10765 -4597 10811 -4595
rect 10765 -4631 10771 -4597
rect 10805 -4631 10811 -4597
rect 10765 -4633 10811 -4631
rect 10765 -4700 10771 -4633
rect 10805 -4700 10811 -4633
rect 10765 -4705 10811 -4700
rect 10765 -4769 10771 -4705
rect 10805 -4769 10811 -4705
rect 10765 -4777 10811 -4769
rect 10765 -4838 10771 -4777
rect 10805 -4838 10811 -4777
rect 10765 -4849 10811 -4838
rect 10765 -4907 10771 -4849
rect 10805 -4907 10811 -4849
rect 10765 -4921 10811 -4907
rect 10765 -4976 10771 -4921
rect 10805 -4976 10811 -4921
rect 10765 -4993 10811 -4976
rect 10765 -5045 10771 -4993
rect 10805 -5045 10811 -4993
rect 10765 -5065 10811 -5045
rect 10765 -5114 10771 -5065
rect 10805 -5114 10811 -5065
rect 10765 -5137 10811 -5114
rect 10765 -5183 10771 -5137
rect 10805 -5183 10811 -5137
rect 10765 -5209 10811 -5183
rect 10765 -5252 10771 -5209
rect 10805 -5252 10811 -5209
rect 10765 -5281 10811 -5252
rect 10765 -5321 10771 -5281
rect 10805 -5321 10811 -5281
rect 10765 -5353 10811 -5321
rect 10765 -5390 10771 -5353
rect 10805 -5390 10811 -5353
rect 10765 -5425 10811 -5390
rect 10765 -5459 10771 -5425
rect 10805 -5459 10811 -5425
rect 10765 -5494 10811 -5459
rect 10765 -5531 10771 -5494
rect 10805 -5531 10811 -5494
rect 10765 -5563 10811 -5531
rect 10765 -5603 10771 -5563
rect 10805 -5603 10811 -5563
rect 10765 -5632 10811 -5603
rect 10765 -5675 10771 -5632
rect 10805 -5675 10811 -5632
rect 10765 -5701 10811 -5675
rect 10765 -5747 10771 -5701
rect 10805 -5747 10811 -5701
rect 10765 -5770 10811 -5747
rect 10765 -5819 10771 -5770
rect 10805 -5819 10811 -5770
rect 10765 -5839 10811 -5819
rect 10765 -5891 10771 -5839
rect 10805 -5891 10811 -5839
rect 10765 -5908 10811 -5891
rect 9313 -5969 9347 -5933
rect 9313 -6039 9347 -6003
rect 9459 -5950 9477 -5916
rect 9511 -5950 9525 -5916
rect 9459 -5988 9525 -5950
rect 9459 -6022 9477 -5988
rect 9511 -6022 9525 -5988
rect 9459 -6034 9525 -6022
rect 10765 -5963 10771 -5908
rect 10805 -5963 10811 -5908
rect 10765 -5977 10811 -5963
rect 9313 -6109 9347 -6073
rect 10765 -6035 10771 -5977
rect 10805 -6035 10811 -5977
rect 10765 -6046 10811 -6035
rect 10765 -6107 10771 -6046
rect 10805 -6107 10811 -6046
rect 10765 -6115 10811 -6107
rect 9347 -6143 9453 -6127
rect 9313 -6161 9453 -6143
rect 9487 -6161 9505 -6127
rect 9471 -6238 9505 -6161
rect 9471 -6340 9505 -6272
rect 10765 -6179 10771 -6115
rect 10805 -6179 10811 -6115
rect 10765 -6184 10811 -6179
rect 10765 -6251 10771 -6184
rect 10805 -6251 10811 -6184
rect 10765 -6253 10811 -6251
rect 10765 -6287 10771 -6253
rect 10805 -6287 10811 -6253
rect 10765 -6322 10811 -6287
rect 10765 -6334 10771 -6322
rect 10031 -6340 10771 -6334
rect 9471 -6374 9489 -6340
rect 9523 -6374 9560 -6340
rect 9594 -6374 9631 -6340
rect 9665 -6374 9701 -6340
rect 9735 -6374 9771 -6340
rect 9805 -6374 9841 -6340
rect 9875 -6374 9911 -6340
rect 9945 -6374 9981 -6340
rect 10015 -6374 10045 -6340
rect 10085 -6374 10117 -6340
rect 10155 -6374 10189 -6340
rect 10225 -6374 10261 -6340
rect 10295 -6374 10331 -6340
rect 10367 -6374 10401 -6340
rect 10439 -6374 10471 -6340
rect 10511 -6374 10541 -6340
rect 10583 -6374 10611 -6340
rect 10655 -6374 10681 -6340
rect 10727 -6374 10765 -6340
rect 10805 -6356 10811 -6322
rect 10799 -6374 10811 -6356
rect 10031 -6380 10811 -6374
<< viali >>
rect 8931 22213 8965 22229
rect 8931 22195 8959 22213
rect 8959 22195 8965 22213
rect 9003 22195 9005 22229
rect 9005 22195 9037 22229
rect 9075 22195 9109 22229
rect 9147 22195 9179 22229
rect 9179 22195 9181 22229
rect 9219 22195 9249 22229
rect 9249 22195 9253 22229
rect 9291 22195 9319 22229
rect 9319 22195 9325 22229
rect 9363 22195 9389 22229
rect 9389 22195 9397 22229
rect 9435 22195 9459 22229
rect 9459 22195 9469 22229
rect 9507 22195 9529 22229
rect 9529 22195 9541 22229
rect 9579 22195 9599 22229
rect 9599 22195 9613 22229
rect 9651 22195 9669 22229
rect 9669 22195 9685 22229
rect 9723 22195 9739 22229
rect 9739 22195 9757 22229
rect 9795 22195 9809 22229
rect 9809 22195 9829 22229
rect 9867 22195 9879 22229
rect 9879 22195 9901 22229
rect 9939 22195 9949 22229
rect 9949 22195 9973 22229
rect 10011 22195 10019 22229
rect 10019 22195 10045 22229
rect 10083 22195 10090 22229
rect 10090 22195 10117 22229
rect 10155 22195 10161 22229
rect 10161 22195 10189 22229
rect 10227 22195 10232 22229
rect 10232 22195 10261 22229
rect 10299 22195 10303 22229
rect 10303 22195 10333 22229
rect 10371 22195 10374 22229
rect 10374 22195 10405 22229
rect 10443 22195 10445 22229
rect 10445 22195 10477 22229
rect 10515 22195 10516 22229
rect 10516 22195 10549 22229
rect 10587 22195 10621 22229
rect 10659 22195 10693 22229
rect 10771 22213 10805 22223
rect 10771 22189 10805 22213
rect 8925 22111 8959 22132
rect 8925 22098 8959 22111
rect 8925 22043 8959 22060
rect 8925 22026 8959 22043
rect 8925 21975 8959 21988
rect 8925 21954 8959 21975
rect 10771 22145 10805 22151
rect 10771 22117 10805 22145
rect 10771 22077 10805 22079
rect 10771 22045 10805 22077
rect 8925 21907 8959 21916
rect 8925 21882 8959 21907
rect 8925 21839 8959 21844
rect 8925 21810 8959 21839
rect 9482 21946 9516 21980
rect 9482 21874 9516 21908
rect 9637 21946 9671 21980
rect 9637 21874 9671 21908
rect 9809 21946 9843 21980
rect 9809 21874 9843 21908
rect 9951 21946 9985 21980
rect 9951 21874 9985 21908
rect 10123 21946 10157 21980
rect 10123 21874 10157 21908
rect 10284 21946 10318 21980
rect 10284 21874 10318 21908
rect 10771 21975 10805 22007
rect 10771 21973 10805 21975
rect 10771 21907 10805 21935
rect 10771 21901 10805 21907
rect 8925 21771 8959 21772
rect 8925 21738 8959 21771
rect 8925 21669 8959 21700
rect 8925 21666 8959 21669
rect 8925 21601 8959 21628
rect 8925 21594 8959 21601
rect 8925 21533 8959 21556
rect 8925 21522 8959 21533
rect 8925 21465 8959 21484
rect 8925 21450 8959 21465
rect 8925 21397 8959 21412
rect 8925 21378 8959 21397
rect 8925 21329 8959 21340
rect 8925 21306 8959 21329
rect 8925 21261 8959 21268
rect 8925 21234 8959 21261
rect 8925 21193 8959 21196
rect 8925 21162 8959 21193
rect 8925 21091 8959 21124
rect 8925 21090 8959 21091
rect 8925 21023 8959 21052
rect 8925 21018 8959 21023
rect 8925 20955 8959 20980
rect 8925 20946 8959 20955
rect 8925 20887 8959 20908
rect 8925 20874 8959 20887
rect 8925 20819 8959 20836
rect 8925 20802 8959 20819
rect 8925 20751 8959 20764
rect 8925 20730 8959 20751
rect 8925 20683 8959 20692
rect 8925 20658 8959 20683
rect 8925 20615 8959 20620
rect 8925 20586 8959 20615
rect 8925 20547 8959 20548
rect 8925 20514 8959 20547
rect 8925 20445 8959 20476
rect 8925 20442 8959 20445
rect 8925 20377 8959 20404
rect 8925 20370 8959 20377
rect 8925 20309 8959 20332
rect 8925 20298 8959 20309
rect 8925 20241 8959 20260
rect 8925 20226 8959 20241
rect 8925 20173 8959 20188
rect 8925 20154 8959 20173
rect 8925 20105 8959 20116
rect 8925 20082 8959 20105
rect 8925 20037 8959 20044
rect 8925 20010 8959 20037
rect 8925 19969 8959 19972
rect 8925 19938 8959 19969
rect 8925 19867 8959 19900
rect 8925 19866 8959 19867
rect 8925 19799 8959 19828
rect 8925 19794 8959 19799
rect 8925 19731 8959 19756
rect 8925 19722 8959 19731
rect 8925 19663 8959 19684
rect 8925 19650 8959 19663
rect 8925 19595 8959 19612
rect 8925 19578 8959 19595
rect 8925 19527 8959 19540
rect 8925 19506 8959 19527
rect 8925 19459 8959 19468
rect 8925 19434 8959 19459
rect 8925 19391 8959 19396
rect 8925 19362 8959 19391
rect 8925 19323 8959 19324
rect 8925 19290 8959 19323
rect 8925 19221 8959 19252
rect 8925 19218 8959 19221
rect 8925 19153 8959 19180
rect 8925 19146 8959 19153
rect 8925 19085 8959 19108
rect 8925 19074 8959 19085
rect 8925 19017 8959 19036
rect 8925 19002 8959 19017
rect 8925 18949 8959 18964
rect 8925 18930 8959 18949
rect 8925 18881 8959 18892
rect 8925 18858 8959 18881
rect 8925 18813 8959 18820
rect 8925 18786 8959 18813
rect 8925 18745 8959 18748
rect 8925 18714 8959 18745
rect 8925 18643 8959 18676
rect 8925 18642 8959 18643
rect 8925 18575 8959 18604
rect 8925 18570 8959 18575
rect 8925 18507 8959 18532
rect 8925 18498 8959 18507
rect 8925 18439 8959 18460
rect 8925 18426 8959 18439
rect 8925 18371 8959 18388
rect 8925 18354 8959 18371
rect 8925 18303 8959 18316
rect 8925 18282 8959 18303
rect 8925 18235 8959 18244
rect 8925 18210 8959 18235
rect 8925 18167 8959 18172
rect 8925 18138 8959 18167
rect 8925 18099 8959 18100
rect 8925 18066 8959 18099
rect 8925 17997 8959 18028
rect 8925 17994 8959 17997
rect 8925 17929 8959 17956
rect 8925 17922 8959 17929
rect 8925 17861 8959 17884
rect 8925 17850 8959 17861
rect 8925 17793 8959 17812
rect 8925 17778 8959 17793
rect 8925 17725 8959 17740
rect 8925 17706 8959 17725
rect 8925 17657 8959 17668
rect 8925 17634 8959 17657
rect 8925 17589 8959 17596
rect 8925 17562 8959 17589
rect 8925 17521 8959 17524
rect 8925 17490 8959 17521
rect 8925 17419 8959 17452
rect 8925 17418 8959 17419
rect 8925 17351 8959 17380
rect 8925 17346 8959 17351
rect 8925 17283 8959 17308
rect 8925 17274 8959 17283
rect 8925 17215 8959 17236
rect 8925 17202 8959 17215
rect 8925 17147 8959 17164
rect 8925 17130 8959 17147
rect 8925 17079 8959 17092
rect 8925 17058 8959 17079
rect 8925 17011 8959 17020
rect 8925 16986 8959 17011
rect 8925 16943 8959 16948
rect 8925 16914 8959 16943
rect 8925 16875 8959 16876
rect 8925 16842 8959 16875
rect 8925 16773 8959 16804
rect 8925 16770 8959 16773
rect 8925 16705 8959 16732
rect 8925 16698 8959 16705
rect 8925 16637 8959 16660
rect 8925 16626 8959 16637
rect 8925 16569 8959 16588
rect 8925 16554 8959 16569
rect 8925 16501 8959 16516
rect 8925 16482 8959 16501
rect 8925 16433 8959 16444
rect 8925 16410 8959 16433
rect 8925 16365 8959 16372
rect 8925 16338 8959 16365
rect 8925 16297 8959 16300
rect 8925 16266 8959 16297
rect 8925 16195 8959 16228
rect 8925 16194 8959 16195
rect 8925 16127 8959 16156
rect 8925 16122 8959 16127
rect 8925 16059 8959 16084
rect 8925 16050 8959 16059
rect 8925 15991 8959 16012
rect 8925 15978 8959 15991
rect 8925 15923 8959 15940
rect 8925 15906 8959 15923
rect 8925 15855 8959 15868
rect 8925 15834 8959 15855
rect 8925 15787 8959 15796
rect 8925 15762 8959 15787
rect 8925 15719 8959 15724
rect 8925 15690 8959 15719
rect 8925 15651 8959 15652
rect 8925 15618 8959 15651
rect 8925 15549 8959 15580
rect 8925 15546 8959 15549
rect 8925 15481 8959 15508
rect 8925 15474 8959 15481
rect 8925 15413 8959 15436
rect 8925 15402 8959 15413
rect 8925 15345 8959 15364
rect 8925 15330 8959 15345
rect 8925 15277 8959 15292
rect 8925 15258 8959 15277
rect 8925 15209 8959 15220
rect 8925 15186 8959 15209
rect 8925 15141 8959 15148
rect 8925 15114 8959 15141
rect 8925 15073 8959 15076
rect 8925 15042 8959 15073
rect 8925 14971 8959 15004
rect 8925 14970 8959 14971
rect 8925 14903 8959 14932
rect 8925 14898 8959 14903
rect 8925 14835 8959 14860
rect 8925 14826 8959 14835
rect 8925 14767 8959 14788
rect 8925 14754 8959 14767
rect 8925 14699 8959 14716
rect 8925 14682 8959 14699
rect 8925 14631 8959 14644
rect 8925 14610 8959 14631
rect 8925 14563 8959 14572
rect 8925 14538 8959 14563
rect 8925 14495 8959 14500
rect 8925 14466 8959 14495
rect 8925 14427 8959 14428
rect 8925 14394 8959 14427
rect 8925 14325 8959 14356
rect 8925 14322 8959 14325
rect 8925 14257 8959 14284
rect 8925 14250 8959 14257
rect 8925 14189 8959 14212
rect 8925 14178 8959 14189
rect 8925 14121 8959 14140
rect 8925 14106 8959 14121
rect 8925 14053 8959 14068
rect 8925 14034 8959 14053
rect 8925 13985 8959 13996
rect 8925 13962 8959 13985
rect 8925 13917 8959 13924
rect 8925 13890 8959 13917
rect 8925 13849 8959 13852
rect 8925 13818 8959 13849
rect 8925 13747 8959 13780
rect 8925 13746 8959 13747
rect 8925 13679 8959 13708
rect 8925 13674 8959 13679
rect 8925 13611 8959 13636
rect 8925 13602 8959 13611
rect 8925 13543 8959 13564
rect 8925 13530 8959 13543
rect 8925 13475 8959 13492
rect 8925 13458 8959 13475
rect 8925 13407 8959 13420
rect 8925 13386 8959 13407
rect 8925 13339 8959 13348
rect 8925 13314 8959 13339
rect 8925 13271 8959 13276
rect 8925 13242 8959 13271
rect 8925 13203 8959 13204
rect 8925 13170 8959 13203
rect 8925 13101 8959 13132
rect 8925 13098 8959 13101
rect 8925 13033 8959 13060
rect 8925 13026 8959 13033
rect 8925 12965 8959 12988
rect 8925 12954 8959 12965
rect 8925 12897 8959 12916
rect 8925 12882 8959 12897
rect 8925 12829 8959 12844
rect 8925 12810 8959 12829
rect 8925 12761 8959 12772
rect 8925 12738 8959 12761
rect 8925 12693 8959 12700
rect 8925 12666 8959 12693
rect 8925 12625 8959 12628
rect 8925 12594 8959 12625
rect 10771 21839 10805 21863
rect 10771 21829 10805 21839
rect 10771 21771 10805 21791
rect 10771 21757 10805 21771
rect 10771 21703 10805 21719
rect 10771 21685 10805 21703
rect 10771 21635 10805 21647
rect 10771 21613 10805 21635
rect 10771 21567 10805 21575
rect 10771 21541 10805 21567
rect 10771 21499 10805 21503
rect 10771 21469 10805 21499
rect 10771 21397 10805 21431
rect 10771 21329 10805 21359
rect 10771 21325 10805 21329
rect 10771 21261 10805 21287
rect 10771 21253 10805 21261
rect 10771 21193 10805 21215
rect 10771 21181 10805 21193
rect 10771 21125 10805 21143
rect 10771 21109 10805 21125
rect 10771 21057 10805 21071
rect 10771 21037 10805 21057
rect 10771 20989 10805 20999
rect 10771 20965 10805 20989
rect 10771 20921 10805 20927
rect 10771 20893 10805 20921
rect 10771 20853 10805 20855
rect 10771 20821 10805 20853
rect 10771 20751 10805 20783
rect 10771 20749 10805 20751
rect 10771 20683 10805 20711
rect 10771 20677 10805 20683
rect 10771 20615 10805 20639
rect 10771 20605 10805 20615
rect 10771 20547 10805 20567
rect 10771 20533 10805 20547
rect 10771 20479 10805 20495
rect 10771 20461 10805 20479
rect 10771 20411 10805 20423
rect 10771 20389 10805 20411
rect 10771 20343 10805 20351
rect 10771 20317 10805 20343
rect 10771 20275 10805 20279
rect 10771 20245 10805 20275
rect 10771 20173 10805 20207
rect 10771 20105 10805 20135
rect 10771 20101 10805 20105
rect 10771 20037 10805 20063
rect 10771 20029 10805 20037
rect 10771 19969 10805 19991
rect 10771 19957 10805 19969
rect 10771 19901 10805 19919
rect 10771 19885 10805 19901
rect 10771 19833 10805 19847
rect 10771 19813 10805 19833
rect 10771 19765 10805 19775
rect 10771 19741 10805 19765
rect 10771 19697 10805 19703
rect 10771 19669 10805 19697
rect 10771 19629 10805 19631
rect 10771 19597 10805 19629
rect 10771 19527 10805 19559
rect 10771 19525 10805 19527
rect 10771 19459 10805 19487
rect 10771 19453 10805 19459
rect 10771 19391 10805 19415
rect 10771 19381 10805 19391
rect 10771 19323 10805 19343
rect 10771 19309 10805 19323
rect 10771 19255 10805 19271
rect 10771 19237 10805 19255
rect 10771 19187 10805 19199
rect 10771 19165 10805 19187
rect 10771 19119 10805 19127
rect 10771 19093 10805 19119
rect 10771 19051 10805 19055
rect 10771 19021 10805 19051
rect 10771 18949 10805 18983
rect 10771 18881 10805 18911
rect 10771 18877 10805 18881
rect 10771 18813 10805 18839
rect 10771 18805 10805 18813
rect 10771 18745 10805 18767
rect 10771 18733 10805 18745
rect 10771 18677 10805 18695
rect 10771 18661 10805 18677
rect 10771 18609 10805 18623
rect 10771 18589 10805 18609
rect 10771 18541 10805 18551
rect 10771 18517 10805 18541
rect 10771 18473 10805 18479
rect 10771 18445 10805 18473
rect 10771 18405 10805 18407
rect 10771 18373 10805 18405
rect 10771 18303 10805 18335
rect 10771 18301 10805 18303
rect 10771 18235 10805 18263
rect 10771 18229 10805 18235
rect 10771 18167 10805 18191
rect 10771 18157 10805 18167
rect 10771 18099 10805 18119
rect 10771 18085 10805 18099
rect 10771 18031 10805 18047
rect 10771 18013 10805 18031
rect 10771 17963 10805 17975
rect 10771 17941 10805 17963
rect 10771 17895 10805 17903
rect 10771 17869 10805 17895
rect 10771 17827 10805 17831
rect 10771 17797 10805 17827
rect 10771 17725 10805 17759
rect 10771 17657 10805 17687
rect 10771 17653 10805 17657
rect 10771 17589 10805 17615
rect 10771 17581 10805 17589
rect 10771 17521 10805 17543
rect 10771 17509 10805 17521
rect 10771 17453 10805 17471
rect 10771 17437 10805 17453
rect 10771 17385 10805 17399
rect 10771 17365 10805 17385
rect 10771 17317 10805 17327
rect 10771 17293 10805 17317
rect 10771 17249 10805 17255
rect 10771 17221 10805 17249
rect 10771 17181 10805 17183
rect 10771 17149 10805 17181
rect 10771 17079 10805 17111
rect 10771 17077 10805 17079
rect 10771 17011 10805 17039
rect 10771 17005 10805 17011
rect 10771 16943 10805 16967
rect 10771 16933 10805 16943
rect 10771 16875 10805 16895
rect 10771 16861 10805 16875
rect 10771 16807 10805 16823
rect 10771 16789 10805 16807
rect 10771 16739 10805 16751
rect 10771 16717 10805 16739
rect 10771 16671 10805 16679
rect 10771 16645 10805 16671
rect 10771 16603 10805 16607
rect 10771 16573 10805 16603
rect 10771 16501 10805 16535
rect 10771 16433 10805 16463
rect 10771 16429 10805 16433
rect 10771 16365 10805 16391
rect 10771 16357 10805 16365
rect 10771 16297 10805 16319
rect 10771 16285 10805 16297
rect 10771 16229 10805 16247
rect 10771 16213 10805 16229
rect 10771 16161 10805 16175
rect 10771 16141 10805 16161
rect 10771 16093 10805 16103
rect 10771 16069 10805 16093
rect 10771 16025 10805 16031
rect 10771 15997 10805 16025
rect 10771 15957 10805 15959
rect 10771 15925 10805 15957
rect 10771 15855 10805 15887
rect 10771 15853 10805 15855
rect 10771 15787 10805 15815
rect 10771 15781 10805 15787
rect 10771 15719 10805 15743
rect 10771 15709 10805 15719
rect 10771 15651 10805 15671
rect 10771 15637 10805 15651
rect 10771 15583 10805 15599
rect 10771 15565 10805 15583
rect 10771 15515 10805 15527
rect 10771 15493 10805 15515
rect 10771 15447 10805 15455
rect 10771 15421 10805 15447
rect 10771 15379 10805 15383
rect 10771 15349 10805 15379
rect 10771 15277 10805 15311
rect 10771 15209 10805 15239
rect 10771 15205 10805 15209
rect 10771 15141 10805 15167
rect 10771 15133 10805 15141
rect 10771 15073 10805 15095
rect 10771 15061 10805 15073
rect 10771 15005 10805 15023
rect 10771 14989 10805 15005
rect 10771 14937 10805 14951
rect 10771 14917 10805 14937
rect 10771 14869 10805 14879
rect 10771 14845 10805 14869
rect 10771 14801 10805 14807
rect 10771 14773 10805 14801
rect 10771 14733 10805 14735
rect 10771 14701 10805 14733
rect 10771 14631 10805 14663
rect 10771 14629 10805 14631
rect 10771 14563 10805 14591
rect 10771 14557 10805 14563
rect 10771 14495 10805 14519
rect 10771 14485 10805 14495
rect 10771 14427 10805 14447
rect 10771 14413 10805 14427
rect 10771 14359 10805 14375
rect 10771 14341 10805 14359
rect 10771 14291 10805 14303
rect 10771 14269 10805 14291
rect 10771 14223 10805 14231
rect 10771 14197 10805 14223
rect 10771 14155 10805 14159
rect 10771 14125 10805 14155
rect 10771 14053 10805 14087
rect 10771 13985 10805 14015
rect 10771 13981 10805 13985
rect 10771 13917 10805 13943
rect 10771 13909 10805 13917
rect 10771 13849 10805 13871
rect 10771 13837 10805 13849
rect 10771 13781 10805 13799
rect 10771 13765 10805 13781
rect 10771 13713 10805 13727
rect 10771 13693 10805 13713
rect 10771 13645 10805 13655
rect 10771 13621 10805 13645
rect 10771 13577 10805 13583
rect 10771 13549 10805 13577
rect 10771 13509 10805 13511
rect 10771 13477 10805 13509
rect 10771 13407 10805 13439
rect 10771 13405 10805 13407
rect 10771 13339 10805 13367
rect 10771 13333 10805 13339
rect 10771 13271 10805 13295
rect 10771 13261 10805 13271
rect 10771 13203 10805 13223
rect 10771 13189 10805 13203
rect 10771 13135 10805 13151
rect 10771 13117 10805 13135
rect 10771 13067 10805 13079
rect 10771 13045 10805 13067
rect 10771 12999 10805 13007
rect 10771 12973 10805 12999
rect 10771 12931 10805 12935
rect 10771 12901 10805 12931
rect 10771 12829 10805 12863
rect 10771 12761 10805 12791
rect 10771 12757 10805 12761
rect 10771 12693 10805 12719
rect 10771 12685 10805 12693
rect 8925 12523 8959 12556
rect 8925 12522 8959 12523
rect 10284 12593 10318 12627
rect 10284 12521 10318 12555
rect 10771 12625 10805 12647
rect 10771 12613 10805 12625
rect 10771 12557 10805 12575
rect 10771 12541 10805 12557
rect 8925 12455 8959 12484
rect 8925 12450 8959 12455
rect 8925 12387 8959 12412
rect 8925 12378 8959 12387
rect 8925 12319 8959 12340
rect 8925 12306 8959 12319
rect 8925 12251 8959 12268
rect 8925 12234 8959 12251
rect 8925 12183 8959 12196
rect 8925 12162 8959 12183
rect 8925 12115 8959 12124
rect 8925 12090 8959 12115
rect 8925 12047 8959 12052
rect 8925 12018 8959 12047
rect 8925 11979 8959 11980
rect 8925 11946 8959 11979
rect 8925 11877 8959 11908
rect 8925 11874 8959 11877
rect 8925 11809 8959 11836
rect 8925 11802 8959 11809
rect 8925 11741 8959 11764
rect 8925 11730 8959 11741
rect 8925 11673 8959 11692
rect 8925 11658 8959 11673
rect 8925 11605 8959 11620
rect 8925 11586 8959 11605
rect 8925 11537 8959 11548
rect 8925 11514 8959 11537
rect 8925 11469 8959 11476
rect 8925 11442 8959 11469
rect 8925 11401 8959 11404
rect 8925 11370 8959 11401
rect 8925 11299 8959 11332
rect 8925 11298 8959 11299
rect 8925 11231 8959 11260
rect 8925 11226 8959 11231
rect 8925 11163 8959 11188
rect 8925 11154 8959 11163
rect 8925 11095 8959 11116
rect 8925 11082 8959 11095
rect 8925 11027 8959 11044
rect 8925 11010 8959 11027
rect 8925 10959 8959 10972
rect 8925 10938 8959 10959
rect 8925 10891 8959 10900
rect 8925 10866 8959 10891
rect 8925 10823 8959 10828
rect 8925 10794 8959 10823
rect 8925 10755 8959 10756
rect 8925 10722 8959 10755
rect 8925 10653 8959 10684
rect 8925 10650 8959 10653
rect 8925 10585 8959 10612
rect 8925 10578 8959 10585
rect 8925 10517 8959 10540
rect 8925 10506 8959 10517
rect 8925 10449 8959 10468
rect 8925 10434 8959 10449
rect 8925 10381 8959 10396
rect 8925 10362 8959 10381
rect 8925 10313 8959 10324
rect 8925 10290 8959 10313
rect 8925 10245 8959 10252
rect 8925 10218 8959 10245
rect 8925 10177 8959 10180
rect 8925 10146 8959 10177
rect 8925 10075 8959 10108
rect 8925 10074 8959 10075
rect 8925 10007 8959 10036
rect 8925 10002 8959 10007
rect 8925 9939 8959 9964
rect 8925 9930 8959 9939
rect 8925 9871 8959 9892
rect 8925 9858 8959 9871
rect 8925 9803 8959 9820
rect 8925 9786 8959 9803
rect 8925 9735 8959 9748
rect 8925 9714 8959 9735
rect 8925 9667 8959 9676
rect 8925 9642 8959 9667
rect 8925 9599 8959 9604
rect 8925 9570 8959 9599
rect 8925 9531 8959 9532
rect 8925 9498 8959 9531
rect 8925 9429 8959 9460
rect 8925 9426 8959 9429
rect 8925 9361 8959 9388
rect 8925 9354 8959 9361
rect 8925 9293 8959 9316
rect 8925 9282 8959 9293
rect 8925 9225 8959 9244
rect 8925 9210 8959 9225
rect 8925 9157 8959 9172
rect 8925 9138 8959 9157
rect 8925 9089 8959 9100
rect 8925 9066 8959 9089
rect 8925 9021 8959 9028
rect 8925 8994 8959 9021
rect 8925 8953 8959 8956
rect 8925 8922 8959 8953
rect 8925 8851 8959 8884
rect 8925 8850 8959 8851
rect 8925 8783 8959 8812
rect 8925 8778 8959 8783
rect 8925 8715 8959 8740
rect 8925 8706 8959 8715
rect 8925 8647 8959 8668
rect 8925 8634 8959 8647
rect 8925 8579 8959 8596
rect 8925 8562 8959 8579
rect 8925 8511 8959 8524
rect 8925 8490 8959 8511
rect 8925 8443 8959 8452
rect 8925 8418 8959 8443
rect 8925 8375 8959 8380
rect 8925 8346 8959 8375
rect 8925 8307 8959 8308
rect 8925 8274 8959 8307
rect 8925 8205 8959 8236
rect 8925 8202 8959 8205
rect 8925 8137 8959 8164
rect 8925 8130 8959 8137
rect 8925 8069 8959 8092
rect 8925 8058 8959 8069
rect 8925 8001 8959 8020
rect 8925 7986 8959 8001
rect 8925 7933 8959 7948
rect 8925 7914 8959 7933
rect 8925 7865 8959 7876
rect 8925 7842 8959 7865
rect 8925 7797 8959 7804
rect 8925 7770 8959 7797
rect 8925 7729 8959 7732
rect 8925 7698 8959 7729
rect 8925 7627 8959 7660
rect 8925 7626 8959 7627
rect 8925 7559 8959 7588
rect 8925 7554 8959 7559
rect 8925 7491 8959 7516
rect 8925 7482 8959 7491
rect 8925 7423 8959 7444
rect 8925 7410 8959 7423
rect 8925 7355 8959 7372
rect 8925 7338 8959 7355
rect 8925 7287 8959 7300
rect 8925 7266 8959 7287
rect 8925 7219 8959 7228
rect 8925 7194 8959 7219
rect 8925 7151 8959 7156
rect 8925 7122 8959 7151
rect 8925 7083 8959 7084
rect 8925 7050 8959 7083
rect 8925 6981 8959 7012
rect 8925 6978 8959 6981
rect 8925 6913 8959 6940
rect 8925 6906 8959 6913
rect 8925 6845 8959 6868
rect 8925 6834 8959 6845
rect 8925 6777 8959 6796
rect 8925 6762 8959 6777
rect 8925 6709 8959 6724
rect 8925 6690 8959 6709
rect 8925 6641 8959 6652
rect 8925 6618 8959 6641
rect 8925 6573 8959 6580
rect 8925 6546 8959 6573
rect 8925 6505 8959 6508
rect 8925 6474 8959 6505
rect 8925 6403 8959 6436
rect 8925 6402 8959 6403
rect 8925 6335 8959 6364
rect 8925 6330 8959 6335
rect 8925 6267 8959 6292
rect 8925 6258 8959 6267
rect 8925 6199 8959 6220
rect 8925 6186 8959 6199
rect 8925 6131 8959 6148
rect 8925 6114 8959 6131
rect 8925 6063 8959 6076
rect 8925 6042 8959 6063
rect 8925 5995 8959 6004
rect 8925 5970 8959 5995
rect 8925 5927 8959 5932
rect 8925 5898 8959 5927
rect 8925 5859 8959 5860
rect 8925 5826 8959 5859
rect 8925 5757 8959 5788
rect 8925 5754 8959 5757
rect 8925 5689 8959 5716
rect 8925 5682 8959 5689
rect 8925 5621 8959 5644
rect 8925 5610 8959 5621
rect 8925 5553 8959 5572
rect 8925 5538 8959 5553
rect 8925 5485 8959 5500
rect 8925 5466 8959 5485
rect 8925 5417 8959 5428
rect 8925 5394 8959 5417
rect 8925 5349 8959 5356
rect 8925 5322 8959 5349
rect 8925 5281 8959 5284
rect 8925 5250 8959 5281
rect 8925 5179 8959 5212
rect 8925 5178 8959 5179
rect 8925 5111 8959 5140
rect 8925 5106 8959 5111
rect 8925 5043 8959 5068
rect 8925 5034 8959 5043
rect 8925 4975 8959 4996
rect 8925 4962 8959 4975
rect 8925 4907 8959 4924
rect 8925 4890 8959 4907
rect 8925 4839 8959 4852
rect 8925 4818 8959 4839
rect 8925 4771 8959 4780
rect 8925 4746 8959 4771
rect 8925 4703 8959 4708
rect 8925 4674 8959 4703
rect 8925 4635 8959 4636
rect 8925 4602 8959 4635
rect 8925 4533 8959 4564
rect 8925 4530 8959 4533
rect 8925 4465 8959 4492
rect 8925 4458 8959 4465
rect 8925 4397 8959 4420
rect 8925 4386 8959 4397
rect 8925 4329 8959 4348
rect 8925 4314 8959 4329
rect 8925 4261 8959 4276
rect 8925 4242 8959 4261
rect 8925 4193 8959 4204
rect 8925 4170 8959 4193
rect 8925 4125 8959 4132
rect 8925 4098 8959 4125
rect 8925 4057 8959 4060
rect 8925 4026 8959 4057
rect 8925 3955 8959 3988
rect 8925 3954 8959 3955
rect 8925 3887 8959 3916
rect 8925 3882 8959 3887
rect 8925 3819 8959 3844
rect 8925 3810 8959 3819
rect 8925 3751 8959 3772
rect 8925 3738 8959 3751
rect 8925 3683 8959 3700
rect 8925 3666 8959 3683
rect 8925 3615 8959 3628
rect 8925 3594 8959 3615
rect 8925 3547 8959 3556
rect 8925 3522 8959 3547
rect 8925 3479 8959 3484
rect 8925 3450 8959 3479
rect 8925 3411 8959 3412
rect 8925 3378 8959 3411
rect 8925 3309 8959 3340
rect 8925 3306 8959 3309
rect 8925 3241 8959 3268
rect 8925 3234 8959 3241
rect 8925 3173 8959 3196
rect 8925 3162 8959 3173
rect 8925 3105 8959 3124
rect 8925 3090 8959 3105
rect 8925 3037 8959 3052
rect 8925 3018 8959 3037
rect 8925 2969 8959 2980
rect 8925 2946 8959 2969
rect 8925 2901 8959 2908
rect 8925 2874 8959 2901
rect 8925 2833 8959 2836
rect 8925 2802 8959 2833
rect 8925 2731 8959 2764
rect 8925 2730 8959 2731
rect 8925 2663 8959 2692
rect 8925 2658 8959 2663
rect 8925 2595 8959 2620
rect 8925 2586 8959 2595
rect 8925 2527 8959 2548
rect 8925 2514 8959 2527
rect 8925 2459 8959 2476
rect 8925 2442 8959 2459
rect 8925 2391 8959 2404
rect 8925 2370 8959 2391
rect 8925 2323 8959 2332
rect 8925 2298 8959 2323
rect 8925 2255 8959 2260
rect 8925 2226 8959 2255
rect 8925 2187 8959 2188
rect 8925 2154 8959 2187
rect 2208 1991 2230 2025
rect 2230 1991 2242 2025
rect 2283 1991 2317 2025
rect 2358 1991 2392 2025
rect 2433 1991 2467 2025
rect 2508 1991 2542 2025
rect 2583 1991 2617 2025
rect 2658 1991 2692 2025
rect 2733 1991 2767 2025
rect 2808 1991 2842 2025
rect 2883 1991 2917 2025
rect 2958 1991 2992 2025
rect 3033 1991 3067 2025
rect 3108 1991 3142 2025
rect 3183 1991 3217 2025
rect 3258 1991 3292 2025
rect 3333 1991 3367 2025
rect 3408 1991 3442 2025
rect 3482 1991 3516 2025
rect 3556 1991 3590 2025
rect 3630 1991 3664 2025
rect 3704 1991 3738 2025
rect 3778 1991 3812 2025
rect 3852 1991 3886 2025
rect 3926 1991 3960 2025
rect 4000 2008 4032 2025
rect 4032 2008 4034 2025
rect 4000 1991 4034 2008
rect 4074 2008 4108 2025
rect 4074 1991 4082 2008
rect 4082 1991 4108 2008
rect 2208 1919 2230 1953
rect 2230 1919 2242 1953
rect 2283 1919 2317 1953
rect 2358 1919 2392 1953
rect 2433 1919 2467 1953
rect 2508 1919 2542 1953
rect 2583 1919 2617 1953
rect 2658 1919 2692 1953
rect 2733 1919 2767 1953
rect 2808 1919 2842 1953
rect 2883 1919 2917 1953
rect 2958 1919 2992 1953
rect 3033 1919 3067 1953
rect 3108 1919 3142 1953
rect 3183 1919 3217 1953
rect 3258 1919 3292 1953
rect 3333 1919 3367 1953
rect 3408 1919 3442 1953
rect 3482 1919 3516 1953
rect 3556 1919 3590 1953
rect 3630 1919 3664 1953
rect 3704 1919 3738 1953
rect 3778 1919 3812 1953
rect 3852 1919 3886 1953
rect 3926 1940 3960 1953
rect 4000 1940 4014 1953
rect 4014 1940 4034 1953
rect 4074 1940 4108 1953
rect 3926 1919 3960 1940
rect 4000 1919 4034 1940
rect 4074 1919 4082 1940
rect 4082 1919 4108 1940
rect 8925 2085 8959 2116
rect 8925 2082 8959 2085
rect 8925 2017 8959 2044
rect 8925 2010 8959 2017
rect 8925 1949 8959 1972
rect 8925 1938 8959 1949
rect 8925 1881 8959 1900
rect 8925 1866 8959 1881
rect 8925 1813 8959 1828
rect 8925 1794 8959 1813
rect 2372 1685 2405 1719
rect 2405 1685 2406 1719
rect 2445 1685 2473 1719
rect 2473 1685 2479 1719
rect 2518 1685 2541 1719
rect 2541 1685 2552 1719
rect 2591 1685 2609 1719
rect 2609 1685 2625 1719
rect 2664 1685 2677 1719
rect 2677 1685 2698 1719
rect 2737 1685 2745 1719
rect 2745 1685 2771 1719
rect 2810 1685 2813 1719
rect 2813 1685 2844 1719
rect 2883 1685 2917 1719
rect 2956 1685 2990 1719
rect 3029 1685 3034 1719
rect 3034 1685 3063 1719
rect 3102 1685 3136 1719
rect 3175 1685 3204 1719
rect 3204 1685 3209 1719
rect 3248 1685 3272 1719
rect 3272 1685 3282 1719
rect 3321 1685 3340 1719
rect 3340 1685 3355 1719
rect 3394 1685 3408 1719
rect 3408 1685 3428 1719
rect 3467 1685 3476 1719
rect 3476 1685 3501 1719
rect 3540 1685 3544 1719
rect 3544 1685 3574 1719
rect 3613 1685 3646 1719
rect 3646 1685 3647 1719
rect 3686 1685 3714 1719
rect 3714 1685 3720 1719
rect 3759 1685 3793 1719
rect 3563 1529 3597 1563
rect 2307 1419 2341 1453
rect 2307 1347 2341 1381
rect 2307 1275 2341 1309
rect 2307 1202 2341 1236
rect 2307 1129 2341 1163
rect 2307 1056 2341 1090
rect 2307 983 2341 1017
rect 2307 910 2341 944
rect 2307 837 2341 871
rect 2307 764 2341 798
rect 2307 691 2341 725
rect 2463 1419 2497 1453
rect 2463 1347 2497 1381
rect 2463 1275 2497 1309
rect 2463 1202 2497 1236
rect 2463 1129 2497 1163
rect 2463 1056 2497 1090
rect 2463 983 2497 1017
rect 2463 910 2497 944
rect 2463 837 2497 871
rect 2463 764 2497 798
rect 2463 691 2497 725
rect 2719 1431 2753 1465
rect 2719 1359 2753 1393
rect 2719 1287 2753 1321
rect 2719 1214 2753 1248
rect 2719 1141 2753 1175
rect 2719 1068 2753 1102
rect 2719 995 2753 1029
rect 2719 922 2753 956
rect 2719 849 2753 883
rect 2719 776 2753 810
rect 2719 703 2753 737
rect 2975 1419 3009 1453
rect 2975 1347 3009 1381
rect 2975 1275 3009 1309
rect 2975 1202 3009 1236
rect 2975 1129 3009 1163
rect 2975 1056 3009 1090
rect 2975 983 3009 1017
rect 2975 910 3009 944
rect 2975 837 3009 871
rect 2975 764 3009 798
rect 2975 691 3009 725
rect 3231 1431 3265 1465
rect 3563 1457 3597 1491
rect 3231 1359 3265 1393
rect 3643 1377 3677 1411
rect 3231 1287 3265 1321
rect 3231 1214 3265 1248
rect 3231 1141 3265 1175
rect 3231 1068 3265 1102
rect 3231 995 3265 1029
rect 3231 922 3265 956
rect 3231 849 3265 883
rect 3231 776 3265 810
rect 3231 703 3265 737
rect 3483 1297 3517 1331
rect 3483 1222 3517 1256
rect 3483 1147 3517 1181
rect 3483 1071 3517 1105
rect 3483 995 3517 1029
rect 3483 919 3517 953
rect 3483 843 3517 877
rect 3483 767 3517 801
rect 3483 691 3517 725
rect 3643 1303 3677 1337
rect 3643 1228 3677 1262
rect 3643 1153 3677 1187
rect 3643 1078 3677 1112
rect 3643 1003 3677 1037
rect 3643 928 3677 962
rect 3643 853 3677 887
rect 3643 778 3677 812
rect 3643 703 3677 737
rect 3759 1379 3793 1411
rect 3759 1377 3793 1379
rect 3759 1311 3793 1337
rect 3759 1303 3793 1311
rect 3759 1243 3793 1262
rect 3759 1228 3793 1243
rect 3759 1175 3793 1187
rect 3759 1153 3793 1175
rect 3759 1107 3793 1112
rect 3759 1078 3793 1107
rect 3759 1005 3793 1037
rect 3759 1003 3793 1005
rect 3759 937 3793 962
rect 3759 928 3793 937
rect 3759 869 3793 887
rect 3759 853 3793 869
rect 3759 801 3793 812
rect 3759 778 3793 801
rect 3759 733 3793 737
rect 3759 703 3793 733
rect 3986 1365 4020 1399
rect 4058 1398 4092 1399
rect 4058 1365 4076 1398
rect 4076 1365 4092 1398
rect 10771 12489 10805 12503
rect 10771 12469 10805 12489
rect 10771 12421 10805 12431
rect 10771 12397 10805 12421
rect 10771 12353 10805 12359
rect 10771 12325 10805 12353
rect 10771 12285 10805 12287
rect 10771 12253 10805 12285
rect 10771 12183 10805 12215
rect 10771 12181 10805 12183
rect 10771 12115 10805 12143
rect 10771 12109 10805 12115
rect 10771 12047 10805 12071
rect 10771 12037 10805 12047
rect 10771 11979 10805 11999
rect 10771 11965 10805 11979
rect 10771 11911 10805 11927
rect 10771 11893 10805 11911
rect 10771 11843 10805 11855
rect 10771 11821 10805 11843
rect 10771 11775 10805 11783
rect 10771 11749 10805 11775
rect 10771 11707 10805 11711
rect 10771 11677 10805 11707
rect 10771 11605 10805 11639
rect 10771 11537 10805 11567
rect 10771 11533 10805 11537
rect 10771 11469 10805 11495
rect 10771 11461 10805 11469
rect 10771 11401 10805 11423
rect 10771 11389 10805 11401
rect 10771 11333 10805 11351
rect 10771 11317 10805 11333
rect 10771 11265 10805 11279
rect 10771 11245 10805 11265
rect 10771 11197 10805 11207
rect 10771 11173 10805 11197
rect 10771 11129 10805 11135
rect 10771 11101 10805 11129
rect 10771 11061 10805 11063
rect 10771 11029 10805 11061
rect 10771 10959 10805 10991
rect 10771 10957 10805 10959
rect 10771 10891 10805 10919
rect 10771 10885 10805 10891
rect 10771 10823 10805 10847
rect 10771 10813 10805 10823
rect 10771 10755 10805 10775
rect 10771 10741 10805 10755
rect 10771 10687 10805 10703
rect 10771 10669 10805 10687
rect 10771 10619 10805 10631
rect 10771 10597 10805 10619
rect 10771 10551 10805 10559
rect 10771 10525 10805 10551
rect 10771 10483 10805 10487
rect 10771 10453 10805 10483
rect 10771 10381 10805 10415
rect 10771 10313 10805 10343
rect 10771 10309 10805 10313
rect 10771 10245 10805 10271
rect 10771 10237 10805 10245
rect 10771 10177 10805 10199
rect 10771 10165 10805 10177
rect 10771 10109 10805 10127
rect 10771 10093 10805 10109
rect 10771 10041 10805 10055
rect 10771 10021 10805 10041
rect 10771 9973 10805 9983
rect 10771 9949 10805 9973
rect 10771 9905 10805 9911
rect 10771 9877 10805 9905
rect 10771 9837 10805 9839
rect 10771 9805 10805 9837
rect 10771 9735 10805 9767
rect 10771 9733 10805 9735
rect 10771 9667 10805 9695
rect 10771 9661 10805 9667
rect 10771 9599 10805 9623
rect 10771 9589 10805 9599
rect 10771 9531 10805 9551
rect 10771 9517 10805 9531
rect 10771 9463 10805 9479
rect 10771 9445 10805 9463
rect 10771 9395 10805 9407
rect 10771 9373 10805 9395
rect 10771 9327 10805 9335
rect 10771 9301 10805 9327
rect 10771 9259 10805 9263
rect 10771 9229 10805 9259
rect 10771 9157 10805 9191
rect 10771 9089 10805 9119
rect 10771 9085 10805 9089
rect 10771 9021 10805 9047
rect 10771 9013 10805 9021
rect 10771 8953 10805 8975
rect 10771 8941 10805 8953
rect 10771 8885 10805 8903
rect 10771 8869 10805 8885
rect 10771 8817 10805 8831
rect 10771 8797 10805 8817
rect 10771 8749 10805 8759
rect 10771 8725 10805 8749
rect 10771 8681 10805 8687
rect 10771 8653 10805 8681
rect 10771 8613 10805 8615
rect 10771 8581 10805 8613
rect 10771 8511 10805 8543
rect 10771 8509 10805 8511
rect 10771 8443 10805 8471
rect 10771 8437 10805 8443
rect 10771 8375 10805 8399
rect 10771 8365 10805 8375
rect 10771 8307 10805 8327
rect 10771 8293 10805 8307
rect 10771 8239 10805 8255
rect 10771 8221 10805 8239
rect 10771 8171 10805 8183
rect 10771 8149 10805 8171
rect 10771 8103 10805 8111
rect 10771 8077 10805 8103
rect 10771 8035 10805 8039
rect 10771 8005 10805 8035
rect 10771 7933 10805 7967
rect 10771 7865 10805 7895
rect 10771 7861 10805 7865
rect 10771 7797 10805 7823
rect 10771 7789 10805 7797
rect 10771 7729 10805 7751
rect 10771 7717 10805 7729
rect 10771 7661 10805 7679
rect 10771 7645 10805 7661
rect 10771 7593 10805 7607
rect 10771 7573 10805 7593
rect 10771 7525 10805 7535
rect 10771 7501 10805 7525
rect 10771 7457 10805 7463
rect 10771 7429 10805 7457
rect 10771 7389 10805 7391
rect 10771 7357 10805 7389
rect 10771 7287 10805 7319
rect 10771 7285 10805 7287
rect 10771 7219 10805 7247
rect 10771 7213 10805 7219
rect 10771 7151 10805 7175
rect 10771 7141 10805 7151
rect 10771 7083 10805 7103
rect 10771 7069 10805 7083
rect 10771 7015 10805 7031
rect 10771 6997 10805 7015
rect 10771 6947 10805 6959
rect 10771 6925 10805 6947
rect 10771 6879 10805 6887
rect 10771 6853 10805 6879
rect 10771 6811 10805 6815
rect 10771 6781 10805 6811
rect 10771 6709 10805 6743
rect 10771 6641 10805 6671
rect 10771 6637 10805 6641
rect 10771 6573 10805 6599
rect 10771 6565 10805 6573
rect 10771 6505 10805 6527
rect 10771 6493 10805 6505
rect 10771 6437 10805 6455
rect 10771 6421 10805 6437
rect 10771 6369 10805 6383
rect 10771 6349 10805 6369
rect 10771 6301 10805 6311
rect 10771 6277 10805 6301
rect 10771 6233 10805 6239
rect 10771 6205 10805 6233
rect 10771 6165 10805 6167
rect 10771 6133 10805 6165
rect 10771 6063 10805 6095
rect 10771 6061 10805 6063
rect 10771 5995 10805 6023
rect 10771 5989 10805 5995
rect 10771 5927 10805 5951
rect 10771 5917 10805 5927
rect 10771 5859 10805 5879
rect 10771 5845 10805 5859
rect 10771 5791 10805 5807
rect 10771 5773 10805 5791
rect 10771 5723 10805 5735
rect 10771 5701 10805 5723
rect 10771 5655 10805 5663
rect 10771 5629 10805 5655
rect 10771 5587 10805 5591
rect 10771 5557 10805 5587
rect 10771 5485 10805 5519
rect 10771 5417 10805 5447
rect 10771 5413 10805 5417
rect 10771 5349 10805 5375
rect 10771 5341 10805 5349
rect 10771 5281 10805 5303
rect 10771 5269 10805 5281
rect 10771 5213 10805 5231
rect 10771 5197 10805 5213
rect 10771 5145 10805 5159
rect 10771 5125 10805 5145
rect 10771 5077 10805 5087
rect 10771 5053 10805 5077
rect 10771 5009 10805 5015
rect 10771 4981 10805 5009
rect 10771 4941 10805 4943
rect 10771 4909 10805 4941
rect 10771 4839 10805 4871
rect 10771 4837 10805 4839
rect 10771 4771 10805 4799
rect 10771 4765 10805 4771
rect 10771 4703 10805 4727
rect 10771 4693 10805 4703
rect 10771 4635 10805 4655
rect 10771 4621 10805 4635
rect 10771 4567 10805 4583
rect 10771 4549 10805 4567
rect 10771 4499 10805 4511
rect 10771 4477 10805 4499
rect 10771 4431 10805 4439
rect 10771 4405 10805 4431
rect 10771 4363 10805 4367
rect 10771 4333 10805 4363
rect 10771 4261 10805 4295
rect 10771 4193 10805 4223
rect 10771 4189 10805 4193
rect 10771 4125 10805 4151
rect 10771 4117 10805 4125
rect 10771 4057 10805 4079
rect 10771 4045 10805 4057
rect 10771 3989 10805 4007
rect 10771 3973 10805 3989
rect 10771 3921 10805 3935
rect 10771 3901 10805 3921
rect 10771 3853 10805 3863
rect 10771 3829 10805 3853
rect 10771 3785 10805 3791
rect 10771 3757 10805 3785
rect 10771 3717 10805 3719
rect 10771 3685 10805 3717
rect 10771 3615 10805 3647
rect 10771 3613 10805 3615
rect 10771 3547 10805 3575
rect 10771 3541 10805 3547
rect 10771 3479 10805 3503
rect 10771 3469 10805 3479
rect 10771 3411 10805 3431
rect 10771 3397 10805 3411
rect 10771 3343 10805 3359
rect 10771 3325 10805 3343
rect 10771 3275 10805 3287
rect 10771 3253 10805 3275
rect 10771 3207 10805 3215
rect 10771 3181 10805 3207
rect 10771 3139 10805 3143
rect 10771 3109 10805 3139
rect 10771 3037 10805 3071
rect 10771 2969 10805 2999
rect 10771 2965 10805 2969
rect 10771 2901 10805 2927
rect 10771 2893 10805 2901
rect 10771 2833 10805 2855
rect 10771 2821 10805 2833
rect 10771 2765 10805 2783
rect 10771 2749 10805 2765
rect 10771 2697 10805 2711
rect 10771 2677 10805 2697
rect 10771 2629 10805 2639
rect 10771 2605 10805 2629
rect 10771 2561 10805 2567
rect 10771 2533 10805 2561
rect 10771 2493 10805 2495
rect 10771 2461 10805 2493
rect 10771 2391 10805 2423
rect 10771 2389 10805 2391
rect 10771 2323 10805 2351
rect 10771 2317 10805 2323
rect 10771 2255 10805 2279
rect 10771 2245 10805 2255
rect 10771 2187 10805 2207
rect 10771 2173 10805 2187
rect 10771 2119 10805 2135
rect 10771 2101 10805 2119
rect 10771 2051 10805 2063
rect 10771 2029 10805 2051
rect 10771 1983 10805 1991
rect 10771 1957 10805 1983
rect 10771 1915 10805 1919
rect 10771 1885 10805 1915
rect 3986 1290 4020 1324
rect 4058 1296 4076 1324
rect 4076 1296 4092 1324
rect 4058 1290 4092 1296
rect 3986 1215 4020 1249
rect 4058 1228 4076 1249
rect 4076 1228 4092 1249
rect 4058 1215 4092 1228
rect 3986 1140 4020 1174
rect 4058 1160 4076 1174
rect 4076 1160 4092 1174
rect 4058 1140 4092 1160
rect 3986 1065 4020 1099
rect 4058 1092 4076 1099
rect 4076 1092 4092 1099
rect 4058 1065 4092 1092
rect 3986 990 4020 1024
rect 4058 990 4092 1024
rect 3986 915 4020 949
rect 4058 922 4092 949
rect 4058 915 4076 922
rect 4076 915 4092 922
rect 3986 840 4020 874
rect 4058 854 4092 874
rect 4058 840 4076 854
rect 4076 840 4092 854
rect 3986 765 4020 799
rect 4058 786 4092 799
rect 4058 765 4076 786
rect 4076 765 4092 786
rect 2372 457 2399 491
rect 2399 457 2406 491
rect 2445 457 2467 491
rect 2467 457 2479 491
rect 2518 457 2535 491
rect 2535 457 2552 491
rect 2591 457 2603 491
rect 2603 457 2625 491
rect 2664 457 2671 491
rect 2671 457 2698 491
rect 2737 457 2739 491
rect 2739 457 2771 491
rect 2810 457 2841 491
rect 2841 457 2844 491
rect 2882 457 2909 491
rect 2909 457 2916 491
rect 2954 457 2977 491
rect 2977 457 2988 491
rect 3026 457 3045 491
rect 3045 457 3060 491
rect 3098 457 3113 491
rect 3113 457 3132 491
rect 3170 457 3181 491
rect 3181 457 3204 491
rect 3242 457 3249 491
rect 3249 457 3276 491
rect 3314 457 3317 491
rect 3317 457 3348 491
rect 3386 457 3419 491
rect 3419 457 3420 491
rect 3458 457 3487 491
rect 3487 457 3492 491
rect 3530 457 3555 491
rect 3555 457 3564 491
rect 3602 457 3623 491
rect 3623 457 3636 491
rect 3674 457 3691 491
rect 3691 457 3708 491
rect 3746 457 3759 491
rect 3759 457 3780 491
rect 3986 690 4020 724
rect 4058 718 4092 724
rect 4058 690 4076 718
rect 4076 690 4092 718
rect 3986 615 4020 649
rect 4058 616 4076 649
rect 4076 616 4092 649
rect 4058 615 4092 616
rect 3986 540 4020 574
rect 4058 548 4076 574
rect 4076 548 4092 574
rect 4058 540 4092 548
rect 3986 466 4020 500
rect 4058 480 4076 500
rect 4076 480 4092 500
rect 4058 466 4092 480
rect 3986 392 4020 426
rect 4058 412 4076 426
rect 4076 412 4092 426
rect 4058 392 4092 412
rect 3986 318 4020 352
rect 4058 344 4076 352
rect 4076 344 4092 352
rect 4058 318 4092 344
rect 2226 271 2238 280
rect 2238 271 2260 280
rect 2300 271 2308 280
rect 2308 271 2334 280
rect 2373 271 2378 280
rect 2378 271 2407 280
rect 2446 271 2448 280
rect 2448 271 2480 280
rect 2519 271 2552 280
rect 2552 271 2553 280
rect 2592 271 2622 280
rect 2622 271 2626 280
rect 2665 271 2692 280
rect 2692 271 2699 280
rect 2738 271 2762 280
rect 2762 271 2772 280
rect 2811 271 2832 280
rect 2832 271 2845 280
rect 2884 271 2902 280
rect 2902 271 2918 280
rect 2957 271 2972 280
rect 2972 271 2991 280
rect 3030 271 3042 280
rect 3042 271 3064 280
rect 3103 271 3112 280
rect 3112 271 3137 280
rect 3176 271 3182 280
rect 3182 271 3210 280
rect 3249 271 3252 280
rect 3252 271 3283 280
rect 2226 246 2260 271
rect 2300 246 2334 271
rect 2373 246 2407 271
rect 2446 246 2480 271
rect 2519 246 2553 271
rect 2592 246 2626 271
rect 2665 246 2699 271
rect 2738 246 2772 271
rect 2811 246 2845 271
rect 2884 246 2918 271
rect 2957 246 2991 271
rect 3030 246 3064 271
rect 3103 246 3137 271
rect 3176 246 3210 271
rect 3249 246 3283 271
rect 3322 246 3356 280
rect 3395 271 3427 280
rect 3427 271 3429 280
rect 3468 271 3496 280
rect 3496 271 3502 280
rect 3541 271 3565 280
rect 3565 271 3575 280
rect 3614 271 3634 280
rect 3634 271 3648 280
rect 3687 271 3703 280
rect 3703 271 3721 280
rect 3760 271 3772 280
rect 3772 271 3794 280
rect 3833 271 3841 280
rect 3841 271 3867 280
rect 3395 246 3429 271
rect 3468 246 3502 271
rect 3541 246 3575 271
rect 3614 246 3648 271
rect 3687 246 3721 271
rect 3760 246 3794 271
rect 3833 246 3867 271
rect 3906 246 3940 280
rect 3979 246 4013 280
rect 4052 276 4076 280
rect 4076 276 4086 280
rect 4052 246 4086 276
rect 2226 174 2248 208
rect 2248 174 2260 208
rect 2300 174 2316 208
rect 2316 174 2334 208
rect 2373 174 2384 208
rect 2384 174 2407 208
rect 2446 174 2452 208
rect 2452 174 2480 208
rect 2519 174 2520 208
rect 2520 174 2553 208
rect 2592 174 2622 208
rect 2622 174 2626 208
rect 2665 174 2690 208
rect 2690 174 2699 208
rect 2738 174 2758 208
rect 2758 174 2772 208
rect 2811 174 2826 208
rect 2826 174 2845 208
rect 2884 174 2894 208
rect 2894 174 2918 208
rect 2957 174 2962 208
rect 2962 174 2991 208
rect 3030 174 3064 208
rect 3103 174 3132 208
rect 3132 174 3137 208
rect 3176 174 3200 208
rect 3200 174 3210 208
rect 3249 174 3268 208
rect 3268 174 3283 208
rect 3322 174 3336 208
rect 3336 174 3356 208
rect 3395 174 3404 208
rect 3404 174 3429 208
rect 3468 174 3472 208
rect 3472 174 3502 208
rect 3541 174 3574 208
rect 3574 174 3575 208
rect 3614 174 3642 208
rect 3642 174 3648 208
rect 3687 174 3710 208
rect 3710 174 3721 208
rect 3760 174 3778 208
rect 3778 174 3794 208
rect 3833 174 3846 208
rect 3846 174 3867 208
rect 3906 174 3914 208
rect 3914 174 3940 208
rect 3979 174 3982 208
rect 3982 174 4013 208
rect 4052 174 4086 208
rect 8197 1313 8204 1347
rect 8204 1313 8231 1347
rect 8301 1313 8317 1347
rect 8317 1313 8335 1347
rect 7931 1219 7965 1253
rect 8003 1219 8037 1253
rect 8307 1245 8341 1275
rect 8307 1241 8341 1245
rect 8307 1176 8341 1201
rect 8307 1167 8341 1176
rect 7863 1141 7897 1161
rect 7863 1127 7897 1141
rect 7863 1073 7897 1085
rect 7863 1051 7897 1073
rect 7863 1005 7897 1009
rect 7863 975 7897 1005
rect 7863 903 7897 933
rect 7863 899 7897 903
rect 7863 835 7897 857
rect 7863 823 7897 835
rect 7863 767 7897 781
rect 7863 747 7897 767
rect 7863 699 7897 705
rect 7863 671 7897 699
rect 7863 597 7897 629
rect 7863 595 7897 597
rect 7863 529 7897 553
rect 7863 519 7897 529
rect 7863 461 7897 478
rect 7863 444 7897 461
rect 7863 393 7897 403
rect 7863 369 7897 393
rect 7863 325 7897 328
rect 7863 294 7897 325
rect 7863 223 7897 253
rect 7863 219 7897 223
rect 7979 1127 8013 1161
rect 7979 1054 8013 1088
rect 7979 981 8013 1015
rect 8191 1127 8225 1161
rect 8191 1054 8225 1088
rect 7979 908 8013 942
rect 7979 835 8013 869
rect 7979 762 8013 796
rect 7979 689 8013 723
rect 7979 616 8013 650
rect 7979 543 8013 577
rect 7979 471 8013 505
rect 7979 399 8013 433
rect 7979 327 8013 361
rect 7979 255 8013 289
rect 8085 961 8119 995
rect 8085 888 8119 922
rect 8085 815 8119 849
rect 8085 742 8119 776
rect 8085 669 8119 703
rect 8085 597 8119 631
rect 8085 525 8119 559
rect 8085 453 8119 487
rect 8085 381 8119 415
rect 8085 309 8119 343
rect 8085 237 8119 271
rect 8191 981 8225 1015
rect 8191 908 8225 942
rect 8191 835 8225 869
rect 8191 762 8225 796
rect 8191 689 8225 723
rect 8191 616 8225 650
rect 8191 543 8225 577
rect 8191 471 8225 505
rect 8191 399 8225 433
rect 8191 327 8225 361
rect 8191 255 8225 289
rect 7979 183 8013 217
rect 8191 183 8225 217
rect 8307 1107 8341 1127
rect 8307 1093 8341 1107
rect 8307 1039 8341 1053
rect 8307 1019 8341 1039
rect 8307 971 8341 979
rect 8307 945 8341 971
rect 8307 903 8341 906
rect 8307 872 8341 903
rect 8307 801 8341 833
rect 8307 799 8341 801
rect 8307 733 8341 760
rect 8307 726 8341 733
rect 8307 665 8341 687
rect 8307 653 8341 665
rect 8307 597 8341 614
rect 8307 580 8341 597
rect 8307 529 8341 541
rect 8307 507 8341 529
rect 8307 461 8341 468
rect 8307 434 8341 461
rect 8307 393 8341 395
rect 8307 361 8341 393
rect 8307 291 8341 322
rect 8307 288 8341 291
rect 8307 223 8341 249
rect 8307 215 8341 223
rect 7863 155 7897 178
rect 7863 144 7897 155
rect 7863 87 7897 103
rect 8307 155 8341 176
rect 8307 142 8341 155
rect 7863 69 7897 87
rect 8005 63 8033 97
rect 8033 63 8039 97
rect 8165 63 8180 97
rect 8180 63 8199 97
rect 8307 87 8341 103
rect 8307 69 8341 87
rect 10771 1813 10805 1847
rect 10771 1745 10805 1775
rect 10771 1741 10805 1745
rect 10771 1677 10805 1703
rect 10771 1669 10805 1677
rect 10771 1609 10805 1631
rect 10771 1597 10805 1609
rect 10771 1541 10805 1559
rect 10771 1525 10805 1541
rect 10771 1473 10805 1487
rect 10771 1453 10805 1473
rect 10771 1405 10805 1415
rect 10771 1381 10805 1405
rect 10771 1337 10805 1343
rect 10771 1309 10805 1337
rect 10771 1269 10805 1271
rect 10771 1237 10805 1269
rect 10771 1167 10805 1199
rect 10771 1165 10805 1167
rect 10771 1099 10805 1127
rect 10771 1093 10805 1099
rect 10771 1031 10805 1055
rect 10771 1021 10805 1031
rect 10771 963 10805 983
rect 10771 949 10805 963
rect 10771 895 10805 911
rect 10771 877 10805 895
rect 10771 827 10805 839
rect 10771 805 10805 827
rect 10771 759 10805 767
rect 10771 733 10805 759
rect 10771 691 10805 695
rect 10771 661 10805 691
rect 10771 589 10805 623
rect 10771 521 10805 551
rect 10771 517 10805 521
rect 10771 453 10805 479
rect 10771 445 10805 453
rect 10771 385 10805 407
rect 10771 373 10805 385
rect 10771 317 10805 335
rect 10771 301 10805 317
rect 10771 249 10805 263
rect 10771 229 10805 249
rect 10771 181 10805 191
rect 10771 157 10805 181
rect 10771 113 10805 119
rect 10771 85 10805 113
rect 10771 45 10805 47
rect 10771 13 10805 45
rect 10771 -57 10805 -25
rect 10771 -59 10805 -57
rect 10771 -125 10805 -97
rect 10771 -131 10805 -125
rect 10771 -193 10805 -169
rect 10771 -203 10805 -193
rect 10771 -261 10805 -241
rect 10771 -275 10805 -261
rect 10771 -329 10805 -313
rect 10771 -347 10805 -329
rect 10771 -397 10805 -385
rect 10771 -419 10805 -397
rect 10771 -465 10805 -457
rect 10771 -491 10805 -465
rect 10771 -533 10805 -529
rect 10771 -563 10805 -533
rect 10771 -635 10805 -601
rect 10771 -703 10805 -673
rect 10771 -707 10805 -703
rect 10771 -771 10805 -745
rect 10771 -779 10805 -771
rect 10771 -839 10805 -817
rect 10771 -851 10805 -839
rect 10771 -907 10805 -889
rect 10771 -923 10805 -907
rect 10771 -975 10805 -961
rect 10771 -995 10805 -975
rect 10771 -1043 10805 -1033
rect 10771 -1067 10805 -1043
rect 10771 -1111 10805 -1105
rect 10771 -1139 10805 -1111
rect 10771 -1179 10805 -1177
rect 10771 -1211 10805 -1179
rect 10771 -1281 10805 -1249
rect 10771 -1283 10805 -1281
rect 10771 -1349 10805 -1321
rect 10771 -1355 10805 -1349
rect 10771 -1417 10805 -1393
rect 10771 -1427 10805 -1417
rect 10771 -1485 10805 -1465
rect 10771 -1499 10805 -1485
rect 10446 -1589 10480 -1555
rect 10446 -1661 10480 -1627
rect 10642 -1590 10676 -1556
rect 10642 -1662 10676 -1628
rect 10771 -1553 10805 -1537
rect 10771 -1571 10805 -1553
rect 10771 -1621 10805 -1609
rect 10771 -1643 10805 -1621
rect 10771 -1689 10805 -1681
rect 10771 -1715 10805 -1689
rect 10771 -1757 10805 -1753
rect 10771 -1787 10805 -1757
rect 10771 -1859 10805 -1825
rect 10771 -1927 10805 -1897
rect 10771 -1931 10805 -1927
rect 10771 -1995 10805 -1969
rect 10771 -2003 10805 -1995
rect 10771 -2063 10805 -2041
rect 10771 -2075 10805 -2063
rect 10771 -2131 10805 -2113
rect 10771 -2147 10805 -2131
rect 10771 -2199 10805 -2185
rect 10771 -2219 10805 -2199
rect 10771 -2267 10805 -2257
rect 10771 -2291 10805 -2267
rect 10771 -2335 10805 -2329
rect 10771 -2363 10805 -2335
rect 10771 -2403 10805 -2401
rect 10771 -2435 10805 -2403
rect 10771 -2505 10805 -2473
rect 10771 -2507 10805 -2505
rect 10771 -2573 10805 -2545
rect 10771 -2579 10805 -2573
rect 10771 -2641 10805 -2617
rect 10771 -2651 10805 -2641
rect 10771 -2709 10805 -2689
rect 10771 -2723 10805 -2709
rect 10771 -2777 10805 -2761
rect 10771 -2795 10805 -2777
rect 10771 -2845 10805 -2833
rect 10771 -2867 10805 -2845
rect 10771 -2913 10805 -2905
rect 10771 -2939 10805 -2913
rect 10771 -2981 10805 -2977
rect 10771 -3011 10805 -2981
rect 9087 -3093 9121 -3059
rect 9087 -3165 9121 -3131
rect 9277 -3143 9311 -3109
rect 9277 -3215 9311 -3181
rect 9221 -3869 9255 -3835
rect 9293 -3869 9327 -3835
rect 10771 -3083 10805 -3049
rect 10771 -3151 10805 -3121
rect 10771 -3155 10805 -3151
rect 10771 -3219 10805 -3193
rect 10771 -3227 10805 -3219
rect 10771 -3287 10805 -3265
rect 10771 -3299 10805 -3287
rect 10771 -3355 10805 -3337
rect 10771 -3371 10805 -3355
rect 10771 -3424 10805 -3409
rect 10771 -3443 10805 -3424
rect 10771 -3493 10805 -3481
rect 10771 -3515 10805 -3493
rect 10771 -3562 10805 -3553
rect 10771 -3587 10805 -3562
rect 10771 -3631 10805 -3625
rect 10771 -3659 10805 -3631
rect 10771 -3700 10805 -3697
rect 10771 -3731 10805 -3700
rect 10771 -3803 10805 -3769
rect 10771 -3872 10805 -3841
rect 10771 -3875 10805 -3872
rect 10771 -3941 10805 -3913
rect 10771 -3947 10805 -3941
rect 10771 -4010 10805 -3985
rect 10771 -4019 10805 -4010
rect 10771 -4079 10805 -4057
rect 10771 -4091 10805 -4079
rect 10771 -4148 10805 -4129
rect 10771 -4163 10805 -4148
rect 10771 -4217 10805 -4201
rect 10771 -4235 10805 -4217
rect 10771 -4286 10805 -4273
rect 10771 -4307 10805 -4286
rect 10771 -4355 10805 -4345
rect 10771 -4379 10805 -4355
rect 10771 -4424 10805 -4417
rect 10771 -4451 10805 -4424
rect 10771 -4493 10805 -4489
rect 10771 -4523 10805 -4493
rect 10771 -4562 10805 -4561
rect 10771 -4595 10805 -4562
rect 10771 -4666 10805 -4633
rect 10771 -4667 10805 -4666
rect 10771 -4735 10805 -4705
rect 10771 -4739 10805 -4735
rect 10771 -4804 10805 -4777
rect 10771 -4811 10805 -4804
rect 10771 -4873 10805 -4849
rect 10771 -4883 10805 -4873
rect 10771 -4942 10805 -4921
rect 10771 -4955 10805 -4942
rect 10771 -5011 10805 -4993
rect 10771 -5027 10805 -5011
rect 10771 -5080 10805 -5065
rect 10771 -5099 10805 -5080
rect 10771 -5149 10805 -5137
rect 10771 -5171 10805 -5149
rect 10771 -5218 10805 -5209
rect 10771 -5243 10805 -5218
rect 10771 -5287 10805 -5281
rect 10771 -5315 10805 -5287
rect 10771 -5356 10805 -5353
rect 10771 -5387 10805 -5356
rect 10771 -5459 10805 -5425
rect 10771 -5528 10805 -5497
rect 10771 -5531 10805 -5528
rect 10771 -5597 10805 -5569
rect 10771 -5603 10805 -5597
rect 10771 -5666 10805 -5641
rect 10771 -5675 10805 -5666
rect 10771 -5735 10805 -5713
rect 10771 -5747 10805 -5735
rect 10771 -5804 10805 -5785
rect 10771 -5819 10805 -5804
rect 10771 -5873 10805 -5857
rect 10771 -5891 10805 -5873
rect 9477 -5950 9511 -5916
rect 9477 -6022 9511 -5988
rect 10771 -5942 10805 -5929
rect 10771 -5963 10805 -5942
rect 10771 -6011 10805 -6001
rect 10771 -6035 10805 -6011
rect 10771 -6080 10805 -6073
rect 10771 -6107 10805 -6080
rect 10771 -6149 10805 -6145
rect 10771 -6179 10805 -6149
rect 10771 -6218 10805 -6217
rect 10771 -6251 10805 -6218
rect 10045 -6374 10051 -6340
rect 10051 -6374 10079 -6340
rect 10117 -6374 10121 -6340
rect 10121 -6374 10151 -6340
rect 10189 -6374 10191 -6340
rect 10191 -6374 10223 -6340
rect 10261 -6374 10295 -6340
rect 10333 -6374 10365 -6340
rect 10365 -6374 10367 -6340
rect 10405 -6374 10435 -6340
rect 10435 -6374 10439 -6340
rect 10477 -6374 10505 -6340
rect 10505 -6374 10511 -6340
rect 10549 -6374 10575 -6340
rect 10575 -6374 10583 -6340
rect 10621 -6374 10645 -6340
rect 10645 -6374 10655 -6340
rect 10693 -6374 10715 -6340
rect 10715 -6374 10727 -6340
rect 10765 -6356 10771 -6340
rect 10771 -6356 10799 -6340
rect 10765 -6374 10799 -6356
<< metal1 >>
rect 8919 22229 10811 22235
rect 8919 22195 8931 22229
rect 8965 22195 9003 22229
rect 9037 22195 9075 22229
rect 9109 22195 9147 22229
rect 9181 22195 9219 22229
rect 9253 22195 9291 22229
rect 9325 22195 9363 22229
rect 9397 22195 9435 22229
rect 9469 22195 9507 22229
rect 9541 22195 9579 22229
rect 9613 22195 9651 22229
rect 9685 22195 9723 22229
rect 9757 22195 9795 22229
rect 9829 22195 9867 22229
rect 9901 22195 9939 22229
rect 9973 22195 10011 22229
rect 10045 22195 10083 22229
rect 10117 22195 10155 22229
rect 10189 22195 10227 22229
rect 10261 22195 10299 22229
rect 10333 22195 10371 22229
rect 10405 22195 10443 22229
rect 10477 22195 10515 22229
rect 10549 22195 10587 22229
rect 10621 22195 10659 22229
rect 10693 22223 10811 22229
rect 10693 22195 10771 22223
rect 8919 22189 10771 22195
rect 10805 22189 10811 22223
rect 8919 22151 8978 22189
tri 8978 22151 9016 22189 nw
tri 10714 22151 10752 22189 ne
rect 10752 22151 10811 22189
rect 8919 22132 8965 22151
tri 8965 22138 8978 22151 nw
tri 10752 22138 10765 22151 ne
rect 8919 22098 8925 22132
rect 8959 22098 8965 22132
rect 8919 22060 8965 22098
rect 8919 22026 8925 22060
rect 8959 22026 8965 22060
rect 8919 21988 8965 22026
rect 10765 22117 10771 22151
rect 10805 22117 10811 22151
rect 10765 22079 10811 22117
rect 10765 22045 10771 22079
rect 10805 22045 10811 22079
rect 10765 22007 10811 22045
rect 8919 21954 8925 21988
rect 8959 21954 8965 21988
rect 8919 21916 8965 21954
rect 8919 21882 8925 21916
rect 8959 21882 8965 21916
rect 8919 21844 8965 21882
rect 9459 21980 9677 21992
tri 9677 21980 9683 21986 sw
tri 9797 21980 9803 21986 se
rect 9803 21980 9991 21992
tri 9991 21980 9997 21986 sw
tri 10111 21980 10117 21986 se
rect 10117 21980 10324 21992
rect 9459 21946 9482 21980
rect 9516 21946 9637 21980
rect 9671 21950 9683 21980
tri 9683 21950 9713 21980 sw
tri 9767 21950 9797 21980 se
rect 9797 21950 9809 21980
rect 9671 21946 9719 21950
rect 9459 21908 9719 21946
rect 9459 21874 9482 21908
rect 9516 21874 9637 21908
rect 9671 21898 9719 21908
rect 9720 21899 9721 21949
rect 9757 21899 9758 21949
rect 9759 21946 9809 21950
rect 9843 21946 9951 21980
rect 9985 21950 9997 21980
tri 9997 21950 10027 21980 sw
tri 10081 21950 10111 21980 se
rect 10111 21950 10123 21980
rect 9985 21946 10033 21950
rect 9759 21908 10033 21946
rect 9759 21898 9809 21908
rect 9671 21874 9689 21898
tri 9689 21874 9713 21898 nw
tri 9767 21874 9791 21898 ne
rect 9791 21874 9809 21898
rect 9843 21874 9951 21908
rect 9985 21898 10033 21908
rect 10034 21899 10035 21949
rect 10071 21899 10072 21949
rect 10073 21946 10123 21950
rect 10157 21946 10284 21980
rect 10318 21946 10324 21980
rect 10073 21908 10324 21946
rect 10073 21898 10123 21908
rect 9985 21874 10003 21898
tri 10003 21874 10027 21898 nw
tri 10081 21874 10105 21898 ne
rect 10105 21874 10123 21898
rect 10157 21874 10284 21908
rect 10318 21874 10324 21908
rect 9459 21863 9678 21874
tri 9678 21863 9689 21874 nw
tri 9791 21863 9802 21874 ne
rect 9802 21863 9992 21874
tri 9992 21863 10003 21874 nw
tri 10105 21863 10116 21874 ne
rect 10116 21863 10324 21874
rect 9459 21862 9677 21863
tri 9677 21862 9678 21863 nw
tri 9802 21862 9803 21863 ne
rect 9803 21862 9991 21863
tri 9991 21862 9992 21863 nw
tri 10116 21862 10117 21863 ne
rect 10117 21862 10324 21863
rect 8919 21810 8925 21844
rect 8959 21810 8965 21844
tri 9475 21837 9500 21862 ne
rect 8919 21772 8965 21810
rect 8919 21738 8925 21772
rect 8959 21738 8965 21772
rect 8919 21700 8965 21738
rect 8919 21666 8925 21700
rect 8959 21666 8965 21700
rect 8919 21628 8965 21666
rect 8919 21594 8925 21628
rect 8959 21594 8965 21628
rect 8919 21556 8965 21594
rect 8919 21522 8925 21556
rect 8959 21522 8965 21556
rect 8919 21484 8965 21522
rect 8919 21450 8925 21484
rect 8959 21450 8965 21484
rect 8919 21412 8965 21450
rect 8919 21378 8925 21412
rect 8959 21378 8965 21412
rect 8919 21340 8965 21378
rect 8919 21306 8925 21340
rect 8959 21306 8965 21340
rect 8919 21268 8965 21306
rect 8919 21234 8925 21268
rect 8959 21234 8965 21268
rect 8919 21196 8965 21234
rect 8919 21162 8925 21196
rect 8959 21162 8965 21196
rect 8919 21124 8965 21162
rect 8919 21090 8925 21124
rect 8959 21090 8965 21124
rect 8919 21052 8965 21090
rect 8919 21018 8925 21052
rect 8959 21018 8965 21052
rect 8919 20980 8965 21018
rect 8919 20946 8925 20980
rect 8959 20946 8965 20980
rect 8919 20908 8965 20946
rect 8919 20874 8925 20908
rect 8959 20874 8965 20908
rect 8919 20836 8965 20874
rect 8919 20802 8925 20836
rect 8959 20802 8965 20836
rect 8919 20764 8965 20802
rect 8919 20730 8925 20764
rect 8959 20730 8965 20764
rect 8919 20692 8965 20730
rect 8919 20658 8925 20692
rect 8959 20658 8965 20692
rect 8919 20620 8965 20658
rect 8919 20586 8925 20620
rect 8959 20586 8965 20620
rect 8919 20548 8965 20586
rect 8919 20514 8925 20548
rect 8959 20514 8965 20548
rect 8919 20476 8965 20514
rect 8919 20442 8925 20476
rect 8959 20442 8965 20476
rect 8919 20404 8965 20442
rect 8919 20370 8925 20404
rect 8959 20370 8965 20404
rect 8919 20332 8965 20370
rect 8919 20298 8925 20332
rect 8959 20298 8965 20332
rect 8919 20260 8965 20298
rect 8919 20226 8925 20260
rect 8959 20226 8965 20260
rect 8919 20188 8965 20226
rect 8919 20154 8925 20188
rect 8959 20154 8965 20188
rect 8919 20116 8965 20154
rect 8919 20082 8925 20116
rect 8959 20082 8965 20116
rect 8919 20044 8965 20082
rect 8919 20010 8925 20044
rect 8959 20010 8965 20044
rect 8919 19972 8965 20010
rect 8919 19938 8925 19972
rect 8959 19938 8965 19972
rect 8919 19900 8965 19938
rect 8919 19866 8925 19900
rect 8959 19866 8965 19900
rect 8919 19828 8965 19866
rect 8919 19794 8925 19828
rect 8959 19794 8965 19828
rect 8919 19756 8965 19794
rect 8919 19722 8925 19756
rect 8959 19722 8965 19756
rect 8919 19684 8965 19722
rect 8919 19650 8925 19684
rect 8959 19650 8965 19684
rect 8919 19612 8965 19650
rect 8919 19578 8925 19612
rect 8959 19578 8965 19612
rect 8919 19540 8965 19578
rect 8919 19506 8925 19540
rect 8959 19506 8965 19540
rect 8919 19468 8965 19506
rect 8919 19434 8925 19468
rect 8959 19434 8965 19468
rect 8919 19396 8965 19434
rect 8919 19362 8925 19396
rect 8959 19362 8965 19396
rect 8919 19324 8965 19362
rect 8919 19290 8925 19324
rect 8959 19290 8965 19324
rect 8919 19252 8965 19290
rect 8919 19218 8925 19252
rect 8959 19218 8965 19252
rect 8919 19180 8965 19218
rect 8919 19146 8925 19180
rect 8959 19146 8965 19180
rect 8919 19108 8965 19146
rect 8919 19074 8925 19108
rect 8959 19074 8965 19108
rect 8919 19036 8965 19074
rect 8919 19002 8925 19036
rect 8959 19002 8965 19036
rect 8919 18964 8965 19002
rect 8919 18930 8925 18964
rect 8959 18930 8965 18964
rect 8919 18892 8965 18930
rect 8919 18858 8925 18892
rect 8959 18858 8965 18892
rect 8919 18820 8965 18858
rect 8919 18786 8925 18820
rect 8959 18786 8965 18820
rect 8919 18748 8965 18786
rect 8919 18714 8925 18748
rect 8959 18714 8965 18748
rect 8919 18676 8965 18714
rect 8919 18642 8925 18676
rect 8959 18642 8965 18676
rect 8919 18604 8965 18642
rect 8919 18570 8925 18604
rect 8959 18570 8965 18604
rect 8919 18532 8965 18570
rect 8919 18498 8925 18532
rect 8959 18498 8965 18532
rect 8919 18460 8965 18498
rect 8919 18426 8925 18460
rect 8959 18426 8965 18460
rect 8919 18388 8965 18426
rect 8919 18354 8925 18388
rect 8959 18354 8965 18388
rect 8919 18316 8965 18354
rect 8919 18282 8925 18316
rect 8959 18282 8965 18316
rect 8919 18244 8965 18282
rect 8919 18210 8925 18244
rect 8959 18210 8965 18244
rect 8919 18172 8965 18210
rect 8919 18138 8925 18172
rect 8959 18138 8965 18172
rect 8919 18100 8965 18138
rect 8919 18066 8925 18100
rect 8959 18066 8965 18100
rect 8919 18028 8965 18066
rect 8919 17994 8925 18028
rect 8959 17994 8965 18028
rect 8919 17956 8965 17994
rect 8919 17922 8925 17956
rect 8959 17922 8965 17956
rect 8919 17884 8965 17922
rect 8919 17850 8925 17884
rect 8959 17850 8965 17884
rect 8919 17812 8965 17850
rect 8919 17778 8925 17812
rect 8959 17778 8965 17812
rect 8919 17740 8965 17778
rect 8919 17706 8925 17740
rect 8959 17706 8965 17740
rect 8919 17668 8965 17706
rect 8919 17634 8925 17668
rect 8959 17634 8965 17668
rect 8919 17596 8965 17634
rect 8919 17562 8925 17596
rect 8959 17562 8965 17596
rect 8919 17524 8965 17562
rect 8919 17490 8925 17524
rect 8959 17490 8965 17524
rect 8919 17452 8965 17490
rect 8919 17418 8925 17452
rect 8959 17418 8965 17452
rect 8919 17380 8965 17418
rect 8919 17346 8925 17380
rect 8959 17346 8965 17380
rect 8919 17308 8965 17346
rect 8919 17274 8925 17308
rect 8959 17274 8965 17308
rect 8919 17236 8965 17274
rect 8919 17202 8925 17236
rect 8959 17202 8965 17236
rect 8919 17164 8965 17202
rect 8919 17130 8925 17164
rect 8959 17130 8965 17164
rect 8919 17092 8965 17130
rect 8919 17058 8925 17092
rect 8959 17058 8965 17092
rect 8919 17020 8965 17058
rect 8919 16986 8925 17020
rect 8959 16986 8965 17020
rect 8919 16948 8965 16986
rect 8919 16914 8925 16948
rect 8959 16914 8965 16948
rect 8919 16876 8965 16914
rect 8919 16842 8925 16876
rect 8959 16842 8965 16876
rect 8919 16804 8965 16842
rect 8919 16770 8925 16804
rect 8959 16770 8965 16804
rect 8919 16732 8965 16770
rect 8919 16698 8925 16732
rect 8959 16698 8965 16732
rect 8919 16660 8965 16698
rect 8919 16626 8925 16660
rect 8959 16626 8965 16660
rect 8919 16588 8965 16626
rect 8919 16554 8925 16588
rect 8959 16554 8965 16588
rect 8919 16516 8965 16554
rect 8919 16482 8925 16516
rect 8959 16482 8965 16516
rect 8919 16444 8965 16482
rect 8919 16410 8925 16444
rect 8959 16410 8965 16444
rect 8919 16372 8965 16410
rect 8919 16338 8925 16372
rect 8959 16338 8965 16372
rect 8919 16300 8965 16338
rect 8919 16266 8925 16300
rect 8959 16266 8965 16300
rect 8919 16228 8965 16266
rect 8919 16194 8925 16228
rect 8959 16194 8965 16228
rect 8919 16156 8965 16194
rect 8919 16122 8925 16156
rect 8959 16122 8965 16156
rect 8919 16084 8965 16122
rect 8919 16050 8925 16084
rect 8959 16050 8965 16084
rect 8919 16012 8965 16050
rect 8919 15978 8925 16012
rect 8959 15978 8965 16012
rect 8919 15940 8965 15978
rect 8919 15906 8925 15940
rect 8959 15906 8965 15940
rect 8919 15868 8965 15906
rect 8919 15834 8925 15868
rect 8959 15834 8965 15868
rect 8919 15796 8965 15834
rect 8919 15762 8925 15796
rect 8959 15762 8965 15796
rect 8919 15724 8965 15762
rect 8919 15690 8925 15724
rect 8959 15690 8965 15724
rect 8919 15652 8965 15690
rect 8919 15618 8925 15652
rect 8959 15618 8965 15652
rect 8919 15580 8965 15618
rect 8919 15546 8925 15580
rect 8959 15546 8965 15580
rect 8919 15508 8965 15546
rect 8919 15474 8925 15508
rect 8959 15474 8965 15508
rect 8919 15436 8965 15474
rect 8919 15402 8925 15436
rect 8959 15402 8965 15436
rect 8919 15364 8965 15402
rect 8919 15330 8925 15364
rect 8959 15330 8965 15364
rect 8919 15292 8965 15330
rect 8919 15258 8925 15292
rect 8959 15258 8965 15292
rect 8919 15220 8965 15258
rect 8919 15186 8925 15220
rect 8959 15186 8965 15220
rect 8919 15148 8965 15186
rect 8919 15114 8925 15148
rect 8959 15114 8965 15148
rect 8919 15076 8965 15114
rect 8919 15042 8925 15076
rect 8959 15042 8965 15076
rect 8919 15004 8965 15042
rect 8919 14970 8925 15004
rect 8959 14970 8965 15004
rect 8919 14932 8965 14970
rect 8919 14898 8925 14932
rect 8959 14898 8965 14932
rect 8919 14860 8965 14898
rect 8919 14826 8925 14860
rect 8959 14826 8965 14860
rect 8919 14788 8965 14826
rect 8919 14754 8925 14788
rect 8959 14754 8965 14788
rect 8919 14716 8965 14754
rect 8919 14682 8925 14716
rect 8959 14682 8965 14716
rect 8919 14644 8965 14682
rect 8919 14610 8925 14644
rect 8959 14610 8965 14644
rect 8919 14572 8965 14610
rect 8919 14538 8925 14572
rect 8959 14538 8965 14572
rect 8919 14500 8965 14538
rect 8919 14466 8925 14500
rect 8959 14466 8965 14500
rect 8919 14428 8965 14466
rect 8919 14394 8925 14428
rect 8959 14394 8965 14428
rect 8919 14356 8965 14394
rect 8919 14322 8925 14356
rect 8959 14322 8965 14356
rect 8919 14284 8965 14322
rect 8919 14250 8925 14284
rect 8959 14250 8965 14284
rect 8919 14212 8965 14250
rect 8919 14178 8925 14212
rect 8959 14178 8965 14212
rect 8919 14140 8965 14178
rect 8919 14106 8925 14140
rect 8959 14106 8965 14140
rect 8919 14068 8965 14106
rect 8919 14034 8925 14068
rect 8959 14034 8965 14068
rect 8919 13996 8965 14034
rect 8919 13962 8925 13996
rect 8959 13962 8965 13996
rect 8919 13924 8965 13962
rect 8919 13890 8925 13924
rect 8959 13890 8965 13924
rect 8919 13852 8965 13890
rect 8919 13818 8925 13852
rect 8959 13818 8965 13852
rect 8919 13780 8965 13818
rect 8919 13746 8925 13780
rect 8959 13746 8965 13780
tri 8913 13727 8919 13733 se
rect 8919 13727 8965 13746
tri 8894 13708 8913 13727 se
rect 8913 13708 8965 13727
tri 8860 13674 8894 13708 se
rect 8894 13674 8925 13708
rect 8959 13674 8965 13708
tri 8841 13655 8860 13674 se
rect 8860 13655 8965 13674
tri 8822 13636 8841 13655 se
rect 8841 13636 8965 13655
tri 8788 13602 8822 13636 se
rect 8822 13602 8925 13636
rect 8959 13602 8965 13636
tri 8773 13587 8788 13602 se
rect 8788 13587 8965 13602
rect 8818 13564 8965 13587
rect 8818 13530 8925 13564
rect 8959 13530 8965 13564
rect 8818 13492 8965 13530
rect 8818 13458 8925 13492
rect 8959 13458 8965 13492
rect 8818 13420 8965 13458
rect 8818 13386 8925 13420
rect 8959 13386 8965 13420
rect 8818 13348 8965 13386
rect 8818 13314 8925 13348
rect 8959 13314 8965 13348
rect 8818 13276 8965 13314
rect 8818 13242 8925 13276
rect 8959 13242 8965 13276
rect 8818 13204 8965 13242
rect 8818 13170 8925 13204
rect 8959 13170 8965 13204
rect 8818 13132 8965 13170
rect 8818 13098 8925 13132
rect 8959 13098 8965 13132
rect 8818 13060 8965 13098
rect 8818 13026 8925 13060
rect 8959 13026 8965 13060
rect 8818 12988 8965 13026
rect 8818 12954 8925 12988
rect 8959 12954 8965 12988
rect 8818 12916 8965 12954
rect 8818 12882 8925 12916
rect 8959 12882 8965 12916
rect 8818 12844 8965 12882
rect 8818 12810 8925 12844
rect 8959 12810 8965 12844
rect 8818 12772 8965 12810
rect 8818 12738 8925 12772
rect 8959 12738 8965 12772
rect 8818 12700 8965 12738
rect 8818 12666 8925 12700
rect 8959 12666 8965 12700
rect 8818 12628 8965 12666
rect 8818 12594 8925 12628
rect 8959 12594 8965 12628
rect 8818 12587 8965 12594
tri 8773 12575 8785 12587 ne
rect 8785 12575 8965 12587
tri 8785 12556 8804 12575 ne
rect 8804 12556 8965 12575
tri 8804 12522 8838 12556 ne
rect 8838 12522 8925 12556
rect 8959 12522 8965 12556
tri 8838 12521 8839 12522 ne
rect 8839 12521 8965 12522
tri 8839 12503 8857 12521 ne
rect 8857 12503 8965 12521
tri 8857 12484 8876 12503 ne
rect 8876 12484 8965 12503
tri 8876 12450 8910 12484 ne
rect 8910 12450 8925 12484
rect 8959 12450 8965 12484
tri 8910 12441 8919 12450 ne
rect 8919 12412 8965 12450
rect 8919 12378 8925 12412
rect 8959 12378 8965 12412
rect 8919 12340 8965 12378
rect 8919 12306 8925 12340
rect 8959 12306 8965 12340
rect 8919 12268 8965 12306
rect 8919 12234 8925 12268
rect 8959 12234 8965 12268
rect 8919 12196 8965 12234
rect 8919 12162 8925 12196
rect 8959 12162 8965 12196
rect 8919 12124 8965 12162
rect 8919 12090 8925 12124
rect 8959 12090 8965 12124
rect 8919 12052 8965 12090
rect 8919 12018 8925 12052
rect 8959 12018 8965 12052
rect 8919 11980 8965 12018
rect 8919 11946 8925 11980
rect 8959 11946 8965 11980
rect 8919 11908 8965 11946
rect 8919 11874 8925 11908
rect 8959 11874 8965 11908
rect 8919 11836 8965 11874
rect 8919 11802 8925 11836
rect 8959 11802 8965 11836
rect 8919 11764 8965 11802
rect 8919 11730 8925 11764
rect 8959 11730 8965 11764
rect 8919 11692 8965 11730
rect 8919 11658 8925 11692
rect 8959 11658 8965 11692
rect 8919 11620 8965 11658
rect 8919 11586 8925 11620
rect 8959 11586 8965 11620
rect 8919 11548 8965 11586
rect 8919 11514 8925 11548
rect 8959 11514 8965 11548
rect 8919 11476 8965 11514
rect 8919 11442 8925 11476
rect 8959 11442 8965 11476
rect 8919 11404 8965 11442
rect 8919 11370 8925 11404
rect 8959 11370 8965 11404
rect 8919 11332 8965 11370
rect 8919 11298 8925 11332
rect 8959 11298 8965 11332
rect 8919 11260 8965 11298
rect 8919 11226 8925 11260
rect 8959 11226 8965 11260
rect 8919 11188 8965 11226
rect 8919 11154 8925 11188
rect 8959 11154 8965 11188
rect 8919 11116 8965 11154
rect 8919 11082 8925 11116
rect 8959 11082 8965 11116
rect 8919 11044 8965 11082
rect 8919 11010 8925 11044
rect 8959 11010 8965 11044
rect 8919 10972 8965 11010
rect 8919 10938 8925 10972
rect 8959 10938 8965 10972
rect 8919 10900 8965 10938
rect 8919 10866 8925 10900
rect 8959 10866 8965 10900
rect 8919 10828 8965 10866
rect 8919 10794 8925 10828
rect 8959 10794 8965 10828
rect 8919 10756 8965 10794
rect 8919 10722 8925 10756
rect 8959 10722 8965 10756
rect 8919 10684 8965 10722
rect 8919 10650 8925 10684
rect 8959 10650 8965 10684
rect 8919 10612 8965 10650
rect 8919 10578 8925 10612
rect 8959 10578 8965 10612
rect 8919 10540 8965 10578
rect 8919 10506 8925 10540
rect 8959 10506 8965 10540
rect 8919 10468 8965 10506
rect 8919 10434 8925 10468
rect 8959 10434 8965 10468
rect 8919 10396 8965 10434
rect 8919 10362 8925 10396
rect 8959 10362 8965 10396
rect 8919 10324 8965 10362
rect 8919 10290 8925 10324
rect 8959 10290 8965 10324
rect 8919 10252 8965 10290
rect 8919 10218 8925 10252
rect 8959 10218 8965 10252
rect 8919 10180 8965 10218
rect 8919 10146 8925 10180
rect 8959 10146 8965 10180
rect 8919 10108 8965 10146
rect 8919 10074 8925 10108
rect 8959 10074 8965 10108
rect 8919 10036 8965 10074
rect 8919 10002 8925 10036
rect 8959 10002 8965 10036
rect 8919 9964 8965 10002
rect 8919 9930 8925 9964
rect 8959 9930 8965 9964
rect 8919 9892 8965 9930
rect 8919 9858 8925 9892
rect 8959 9858 8965 9892
rect 8919 9820 8965 9858
rect 8919 9786 8925 9820
rect 8959 9786 8965 9820
rect 8919 9748 8965 9786
rect 8919 9714 8925 9748
rect 8959 9714 8965 9748
rect 8919 9676 8965 9714
rect 8919 9642 8925 9676
rect 8959 9642 8965 9676
rect 8919 9604 8965 9642
rect 8919 9570 8925 9604
rect 8959 9570 8965 9604
rect 8919 9532 8965 9570
rect 8919 9498 8925 9532
rect 8959 9498 8965 9532
rect 8919 9460 8965 9498
rect 8919 9426 8925 9460
rect 8959 9426 8965 9460
rect 8919 9388 8965 9426
rect 8919 9354 8925 9388
rect 8959 9354 8965 9388
rect 8919 9316 8965 9354
rect 8919 9282 8925 9316
rect 8959 9282 8965 9316
rect 8919 9244 8965 9282
rect 8919 9210 8925 9244
rect 8959 9210 8965 9244
rect 8919 9172 8965 9210
rect 8919 9138 8925 9172
rect 8959 9138 8965 9172
rect 8919 9100 8965 9138
rect 8919 9066 8925 9100
rect 8959 9066 8965 9100
rect 8919 9028 8965 9066
rect 8919 8994 8925 9028
rect 8959 8994 8965 9028
rect 8919 8956 8965 8994
rect 8919 8922 8925 8956
rect 8959 8922 8965 8956
rect 8919 8884 8965 8922
rect 8919 8850 8925 8884
rect 8959 8850 8965 8884
rect 8919 8812 8965 8850
rect 8919 8778 8925 8812
rect 8959 8778 8965 8812
rect 8919 8740 8965 8778
rect 8919 8706 8925 8740
rect 8959 8706 8965 8740
rect 8919 8668 8965 8706
rect 8919 8634 8925 8668
rect 8959 8634 8965 8668
rect 8919 8596 8965 8634
rect 8919 8562 8925 8596
rect 8959 8562 8965 8596
rect 8919 8524 8965 8562
rect 8919 8490 8925 8524
rect 8959 8490 8965 8524
rect 8919 8452 8965 8490
rect 8919 8418 8925 8452
rect 8959 8418 8965 8452
rect 8919 8380 8965 8418
rect 8919 8346 8925 8380
rect 8959 8346 8965 8380
rect 8919 8308 8965 8346
rect 8919 8274 8925 8308
rect 8959 8274 8965 8308
rect 8919 8236 8965 8274
rect 8919 8202 8925 8236
rect 8959 8202 8965 8236
rect 8919 8164 8965 8202
rect 8919 8130 8925 8164
rect 8959 8130 8965 8164
rect 8919 8092 8965 8130
rect 8919 8058 8925 8092
rect 8959 8058 8965 8092
rect 8919 8020 8965 8058
rect 8919 7986 8925 8020
rect 8959 7986 8965 8020
rect 8919 7948 8965 7986
rect 8919 7914 8925 7948
rect 8959 7914 8965 7948
rect 8919 7876 8965 7914
rect 8919 7842 8925 7876
rect 8959 7842 8965 7876
rect 8919 7804 8965 7842
rect 8919 7770 8925 7804
rect 8959 7770 8965 7804
rect 8919 7732 8965 7770
rect 8919 7698 8925 7732
rect 8959 7698 8965 7732
rect 8919 7660 8965 7698
rect 8919 7626 8925 7660
rect 8959 7626 8965 7660
rect 8919 7588 8965 7626
rect 8919 7554 8925 7588
rect 8959 7554 8965 7588
rect 8919 7516 8965 7554
rect 8919 7482 8925 7516
rect 8959 7482 8965 7516
rect 8919 7444 8965 7482
rect 8919 7410 8925 7444
rect 8959 7410 8965 7444
rect 8919 7372 8965 7410
rect 8919 7338 8925 7372
rect 8959 7338 8965 7372
rect 8919 7300 8965 7338
rect 8919 7266 8925 7300
rect 8959 7266 8965 7300
rect 8919 7228 8965 7266
rect 8919 7194 8925 7228
rect 8959 7194 8965 7228
rect 8919 7156 8965 7194
rect 8919 7122 8925 7156
rect 8959 7122 8965 7156
rect 8919 7084 8965 7122
rect 8919 7050 8925 7084
rect 8959 7050 8965 7084
rect 8919 7012 8965 7050
rect 8919 6978 8925 7012
rect 8959 6978 8965 7012
rect 8919 6940 8965 6978
rect 8919 6906 8925 6940
rect 8959 6906 8965 6940
rect 8919 6868 8965 6906
rect 8919 6834 8925 6868
rect 8959 6834 8965 6868
rect 8919 6796 8965 6834
rect 8919 6762 8925 6796
rect 8959 6762 8965 6796
rect 8919 6724 8965 6762
rect 8919 6690 8925 6724
rect 8959 6690 8965 6724
rect 8919 6652 8965 6690
rect 8919 6618 8925 6652
rect 8959 6618 8965 6652
rect 8919 6580 8965 6618
rect 8919 6546 8925 6580
rect 8959 6546 8965 6580
rect 8919 6508 8965 6546
rect 8919 6474 8925 6508
rect 8959 6474 8965 6508
rect 8919 6436 8965 6474
rect 8919 6402 8925 6436
rect 8959 6402 8965 6436
rect 8919 6364 8965 6402
rect 8919 6330 8925 6364
rect 8959 6330 8965 6364
rect 8919 6292 8965 6330
rect 8919 6258 8925 6292
rect 8959 6258 8965 6292
rect 8919 6220 8965 6258
rect 8919 6186 8925 6220
rect 8959 6186 8965 6220
rect 8919 6148 8965 6186
rect 8919 6114 8925 6148
rect 8959 6114 8965 6148
rect 8919 6076 8965 6114
rect 8919 6042 8925 6076
rect 8959 6042 8965 6076
rect 8919 6004 8965 6042
rect 8919 5970 8925 6004
rect 8959 5970 8965 6004
rect 8919 5932 8965 5970
rect 8919 5898 8925 5932
rect 8959 5898 8965 5932
rect 8919 5860 8965 5898
rect 8919 5826 8925 5860
rect 8959 5826 8965 5860
rect 8919 5788 8965 5826
rect 8919 5754 8925 5788
rect 8959 5754 8965 5788
rect 8919 5716 8965 5754
rect 8919 5682 8925 5716
rect 8959 5682 8965 5716
rect 8919 5644 8965 5682
rect 8919 5610 8925 5644
rect 8959 5610 8965 5644
rect 8919 5572 8965 5610
rect 8919 5538 8925 5572
rect 8959 5538 8965 5572
rect 8919 5500 8965 5538
rect 8919 5466 8925 5500
rect 8959 5466 8965 5500
rect 8919 5428 8965 5466
rect 8919 5394 8925 5428
rect 8959 5394 8965 5428
rect 8919 5356 8965 5394
rect 8919 5322 8925 5356
rect 8959 5322 8965 5356
rect 8919 5284 8965 5322
rect 8919 5250 8925 5284
rect 8959 5250 8965 5284
rect 8919 5212 8965 5250
rect 8919 5178 8925 5212
rect 8959 5178 8965 5212
rect 8919 5140 8965 5178
rect 8919 5106 8925 5140
rect 8959 5106 8965 5140
rect 8919 5068 8965 5106
rect 8919 5034 8925 5068
rect 8959 5034 8965 5068
rect 8919 4996 8965 5034
rect 8919 4962 8925 4996
rect 8959 4962 8965 4996
rect 8919 4924 8965 4962
rect 8919 4890 8925 4924
rect 8959 4890 8965 4924
rect 8919 4852 8965 4890
rect 8919 4818 8925 4852
rect 8959 4818 8965 4852
rect 8919 4780 8965 4818
rect 8919 4746 8925 4780
rect 8959 4746 8965 4780
rect 8919 4708 8965 4746
rect 8919 4674 8925 4708
rect 8959 4674 8965 4708
rect 8919 4636 8965 4674
rect 8919 4602 8925 4636
rect 8959 4602 8965 4636
rect 8919 4564 8965 4602
rect 8919 4530 8925 4564
rect 8959 4530 8965 4564
rect 8919 4492 8965 4530
rect 8919 4458 8925 4492
rect 8959 4458 8965 4492
rect 8919 4420 8965 4458
rect 8919 4386 8925 4420
rect 8959 4386 8965 4420
rect 8919 4348 8965 4386
rect 8919 4314 8925 4348
rect 8959 4314 8965 4348
rect 8919 4276 8965 4314
rect 8919 4242 8925 4276
rect 8959 4242 8965 4276
rect 8919 4204 8965 4242
rect 8919 4170 8925 4204
rect 8959 4170 8965 4204
rect 8919 4132 8965 4170
rect 8919 4098 8925 4132
rect 8959 4098 8965 4132
rect 8919 4060 8965 4098
rect 8919 4026 8925 4060
rect 8959 4026 8965 4060
rect 8919 3988 8965 4026
rect 8919 3954 8925 3988
rect 8959 3954 8965 3988
rect 8919 3916 8965 3954
rect 8919 3882 8925 3916
rect 8959 3882 8965 3916
rect 8919 3844 8965 3882
rect 8919 3810 8925 3844
rect 8959 3810 8965 3844
rect 8919 3772 8965 3810
rect 8919 3738 8925 3772
rect 8959 3738 8965 3772
rect 8919 3700 8965 3738
rect 8919 3666 8925 3700
rect 8959 3666 8965 3700
rect 8919 3628 8965 3666
rect 8919 3594 8925 3628
rect 8959 3594 8965 3628
rect 8919 3556 8965 3594
rect 8919 3522 8925 3556
rect 8959 3522 8965 3556
rect 8919 3484 8965 3522
rect 8919 3450 8925 3484
rect 8959 3450 8965 3484
rect 8919 3412 8965 3450
rect 8919 3378 8925 3412
rect 8959 3378 8965 3412
rect 8919 3340 8965 3378
rect 8919 3306 8925 3340
rect 8959 3306 8965 3340
rect 8919 3268 8965 3306
rect 8919 3234 8925 3268
rect 8959 3234 8965 3268
rect 8919 3196 8965 3234
rect 8919 3162 8925 3196
rect 8959 3162 8965 3196
rect 8919 3124 8965 3162
rect 8919 3090 8925 3124
rect 8959 3090 8965 3124
rect 8919 3052 8965 3090
rect 8919 3018 8925 3052
rect 8959 3018 8965 3052
rect 8919 2980 8965 3018
rect 8919 2946 8925 2980
rect 8959 2946 8965 2980
rect 8919 2908 8965 2946
rect 8919 2874 8925 2908
rect 8959 2874 8965 2908
rect 8919 2836 8965 2874
rect 8919 2802 8925 2836
rect 8959 2802 8965 2836
rect 8919 2764 8965 2802
rect 8919 2730 8925 2764
rect 8959 2730 8965 2764
rect 8919 2692 8965 2730
rect 8919 2658 8925 2692
rect 8959 2658 8965 2692
tri 866 2639 884 2657 se
tri 847 2620 866 2639 se
rect 866 2620 884 2639
tri 844 2617 847 2620 se
rect 847 2617 884 2620
tri 936 2639 954 2657 sw
rect 936 2620 954 2639
tri 954 2620 973 2639 sw
rect 8919 2620 8965 2658
rect 936 2617 973 2620
tri 973 2617 976 2620 sw
rect 8919 2586 8925 2620
rect 8959 2586 8965 2620
rect 8919 2548 8965 2586
rect 8919 2514 8925 2548
rect 8959 2514 8965 2548
rect 8919 2476 8965 2514
rect 8919 2442 8925 2476
rect 8959 2442 8965 2476
rect 8919 2404 8965 2442
rect 8919 2370 8925 2404
rect 8959 2370 8965 2404
rect 8919 2332 8965 2370
rect 8919 2298 8925 2332
rect 8959 2298 8965 2332
rect 8919 2260 8965 2298
rect 8919 2226 8925 2260
rect 8959 2226 8965 2260
rect 8919 2188 8965 2226
rect 8919 2154 8925 2188
rect 8959 2154 8965 2188
rect 8919 2116 8965 2154
rect 2196 2093 4610 2104
rect 2196 2025 3987 2093
rect 4103 2076 4610 2093
rect 4103 2063 4597 2076
tri 4597 2063 4610 2076 nw
rect 8919 2082 8925 2116
rect 8959 2082 8965 2116
rect 4103 2044 4578 2063
tri 4578 2044 4597 2063 nw
rect 8919 2044 8965 2082
rect 4103 2031 4565 2044
tri 4565 2031 4578 2044 nw
rect 4103 2025 4544 2031
rect 2196 1991 2208 2025
rect 2242 1991 2283 2025
rect 2317 1991 2358 2025
rect 2392 1991 2433 2025
rect 2467 1991 2508 2025
rect 2542 1991 2583 2025
rect 2617 1991 2658 2025
rect 2692 1991 2733 2025
rect 2767 1991 2808 2025
rect 2842 1991 2883 2025
rect 2917 1991 2958 2025
rect 2992 1991 3033 2025
rect 3067 1991 3108 2025
rect 3142 1991 3183 2025
rect 3217 1991 3258 2025
rect 3292 1991 3333 2025
rect 3367 1991 3408 2025
rect 3442 1991 3482 2025
rect 3516 1991 3556 2025
rect 3590 1991 3630 2025
rect 3664 1991 3704 2025
rect 3738 1991 3778 2025
rect 3812 1991 3852 2025
rect 3886 1991 3926 2025
rect 3960 1991 3987 2025
rect 4108 2010 4544 2025
tri 4544 2010 4565 2031 nw
rect 8919 2010 8925 2044
rect 8959 2010 8965 2044
rect 4108 1991 4525 2010
tri 4525 1991 4544 2010 nw
rect 2196 1953 3987 1991
rect 4103 1972 4506 1991
tri 4506 1972 4525 1991 nw
rect 8919 1972 8965 2010
rect 4103 1953 4472 1972
rect 2196 1919 2208 1953
rect 2242 1919 2283 1953
rect 2317 1919 2358 1953
rect 2392 1919 2433 1953
rect 2467 1919 2508 1953
rect 2542 1919 2583 1953
rect 2617 1919 2658 1953
rect 2692 1919 2733 1953
rect 2767 1919 2808 1953
rect 2842 1919 2883 1953
rect 2917 1919 2958 1953
rect 2992 1919 3033 1953
rect 3067 1919 3108 1953
rect 3142 1919 3183 1953
rect 3217 1919 3258 1953
rect 3292 1919 3333 1953
rect 3367 1919 3408 1953
rect 3442 1919 3482 1953
rect 3516 1919 3556 1953
rect 3590 1919 3630 1953
rect 3664 1919 3704 1953
rect 3738 1919 3778 1953
rect 3812 1919 3852 1953
rect 3886 1919 3926 1953
rect 3960 1919 3987 1953
rect 4108 1938 4472 1953
tri 4472 1938 4506 1972 nw
rect 8919 1938 8925 1972
rect 8959 1938 8965 1972
rect 4108 1919 4453 1938
tri 4453 1919 4472 1938 nw
rect 2196 1913 3987 1919
rect 4103 1913 4447 1919
tri 4447 1913 4453 1919 nw
rect 8919 1900 8965 1938
rect 8919 1866 8925 1900
rect 8959 1866 8965 1900
rect 8919 1828 8965 1866
rect 8919 1794 8925 1828
rect 8959 1794 8965 1828
rect 8919 1782 8965 1794
rect 2253 1719 3755 1725
rect 2253 1685 2372 1719
rect 2406 1685 2445 1719
rect 2479 1685 2518 1719
rect 2552 1685 2591 1719
rect 2625 1685 2664 1719
rect 2698 1685 2737 1719
rect 2771 1685 2810 1719
rect 2844 1685 2883 1719
rect 2917 1685 2956 1719
rect 2990 1685 3029 1719
rect 3063 1685 3102 1719
rect 3136 1685 3175 1719
rect 3209 1685 3248 1719
rect 3282 1685 3321 1719
rect 3355 1685 3394 1719
rect 3428 1685 3467 1719
rect 3501 1685 3540 1719
rect 3574 1685 3613 1719
rect 3647 1685 3686 1719
rect 3720 1685 3755 1719
rect 2253 1679 3755 1685
tri 3743 1673 3749 1679 ne
rect 3749 1673 3755 1679
rect 3807 1673 3819 1725
rect 3871 1673 3877 1725
tri 3317 1645 3322 1650 se
rect 3322 1645 3732 1650
tri 3732 1645 3737 1650 sw
tri 3889 1645 3894 1650 se
rect 3894 1645 9061 1650
tri 3303 1631 3317 1645 se
rect 3317 1631 9061 1645
tri 3270 1598 3303 1631 se
rect 3303 1598 9061 1631
rect 9113 1598 9125 1650
rect 9177 1598 9183 1650
tri 3269 1597 3270 1598 se
rect 3270 1597 3343 1598
tri 3343 1597 3344 1598 nw
tri 3248 1576 3269 1597 se
rect 3269 1576 3322 1597
tri 3322 1576 3343 1597 nw
tri 3241 1569 3248 1576 se
rect 3248 1569 3315 1576
tri 3315 1569 3322 1576 nw
tri 3235 1563 3241 1569 se
rect 3241 1563 3309 1569
tri 3309 1563 3315 1569 nw
rect 3551 1563 3609 1569
tri 3229 1557 3235 1563 se
rect 3235 1557 3303 1563
tri 3303 1557 3309 1563 nw
rect 2269 1505 3296 1557
tri 3296 1550 3303 1557 nw
tri 2682 1491 2696 1505 ne
rect 2696 1491 2776 1505
tri 2776 1491 2790 1505 nw
tri 3194 1491 3208 1505 ne
rect 3208 1491 3296 1505
tri 2696 1477 2710 1491 ne
rect 2710 1465 2762 1491
tri 2762 1477 2776 1491 nw
tri 3208 1477 3222 1491 ne
rect 3222 1465 3296 1491
rect 3551 1529 3563 1563
rect 3597 1529 3609 1563
rect 3551 1497 3609 1529
tri 3609 1497 3634 1522 sw
rect 3551 1491 7335 1497
rect 2298 1453 2350 1465
rect 2298 1419 2307 1453
rect 2341 1419 2350 1453
rect 2298 1381 2350 1419
rect 2298 1347 2307 1381
rect 2341 1347 2350 1381
rect 2298 1309 2350 1347
rect 2298 1275 2307 1309
rect 2341 1275 2350 1309
rect 2298 1236 2350 1275
rect 2298 1202 2307 1236
rect 2341 1202 2350 1236
rect 2298 1163 2350 1202
rect 2298 1129 2307 1163
rect 2341 1129 2350 1163
rect 2298 1090 2350 1129
rect 2298 1056 2307 1090
rect 2341 1056 2350 1090
rect 2298 1017 2350 1056
rect 2298 983 2307 1017
rect 2341 983 2350 1017
rect 2298 944 2350 983
rect 2298 910 2307 944
rect 2341 910 2350 944
rect 2298 871 2350 910
rect 2298 837 2307 871
rect 2341 837 2350 871
rect 2298 798 2350 837
rect 2298 764 2307 798
rect 2341 764 2350 798
rect 2298 725 2350 764
rect 2298 691 2307 725
rect 2341 691 2350 725
tri 2290 671 2298 679 se
rect 2298 671 2350 691
rect 2454 1453 2506 1465
rect 2454 1419 2463 1453
rect 2497 1419 2506 1453
rect 2454 1381 2506 1419
rect 2454 1347 2463 1381
rect 2497 1347 2506 1381
rect 2454 1309 2506 1347
rect 2454 1275 2463 1309
rect 2497 1275 2506 1309
rect 2454 1236 2506 1275
rect 2454 1202 2463 1236
rect 2497 1202 2506 1236
rect 2454 1163 2506 1202
rect 2454 1129 2463 1163
rect 2497 1129 2506 1163
rect 2454 1090 2506 1129
rect 2454 1056 2463 1090
rect 2497 1056 2506 1090
rect 2454 1017 2506 1056
rect 2454 983 2463 1017
rect 2497 983 2506 1017
rect 2454 944 2506 983
rect 2454 910 2463 944
rect 2497 910 2506 944
rect 2454 871 2506 910
rect 2454 837 2463 871
rect 2497 837 2506 871
rect 2454 798 2506 837
rect 2454 764 2463 798
rect 2497 764 2506 798
rect 2454 725 2506 764
rect 2454 691 2463 725
rect 2497 691 2506 725
rect 2710 1431 2719 1465
rect 2753 1431 2762 1465
rect 2710 1393 2762 1431
rect 2710 1359 2719 1393
rect 2753 1359 2762 1393
rect 2710 1321 2762 1359
rect 2710 1287 2719 1321
rect 2753 1287 2762 1321
rect 2710 1248 2762 1287
rect 2710 1214 2719 1248
rect 2753 1214 2762 1248
rect 2710 1175 2762 1214
rect 2710 1141 2719 1175
rect 2753 1141 2762 1175
rect 2710 1102 2762 1141
rect 2710 1068 2719 1102
rect 2753 1068 2762 1102
rect 2710 1029 2762 1068
rect 2710 995 2719 1029
rect 2753 995 2762 1029
rect 2710 956 2762 995
rect 2710 922 2719 956
rect 2753 922 2762 956
rect 2710 883 2762 922
rect 2710 849 2719 883
rect 2753 849 2762 883
rect 2710 810 2762 849
rect 2710 776 2719 810
rect 2753 776 2762 810
rect 2710 737 2762 776
rect 2710 703 2719 737
rect 2753 703 2762 737
rect 2710 691 2762 703
rect 2966 1453 3018 1465
rect 2966 1419 2975 1453
rect 3009 1419 3018 1453
rect 2966 1381 3018 1419
rect 2966 1347 2975 1381
rect 3009 1347 3018 1381
rect 2966 1309 3018 1347
rect 2966 1275 2975 1309
rect 3009 1275 3018 1309
rect 2966 1236 3018 1275
rect 2966 1202 2975 1236
rect 3009 1202 3018 1236
rect 2966 1163 3018 1202
rect 2966 1129 2975 1163
rect 3009 1129 3018 1163
rect 2966 1090 3018 1129
rect 2966 1056 2975 1090
rect 3009 1056 3018 1090
rect 2966 1017 3018 1056
rect 2966 983 2975 1017
rect 3009 983 3018 1017
rect 2966 944 3018 983
rect 2966 910 2975 944
rect 3009 910 3018 944
rect 2966 871 3018 910
rect 2966 837 2975 871
rect 3009 837 3018 871
rect 2966 798 3018 837
rect 2966 764 2975 798
rect 3009 764 3018 798
rect 2966 725 3018 764
rect 2966 691 2975 725
rect 3009 691 3018 725
rect 3222 1431 3231 1465
rect 3265 1457 3296 1465
tri 3296 1457 3316 1477 sw
rect 3551 1457 3563 1491
rect 3597 1457 7335 1491
rect 3265 1453 3316 1457
tri 3316 1453 3320 1457 sw
rect 3265 1451 3320 1453
tri 3320 1451 3322 1453 sw
rect 3551 1451 7335 1457
rect 3265 1445 3322 1451
tri 3322 1445 3328 1451 sw
tri 7323 1445 7329 1451 ne
rect 7329 1445 7335 1451
rect 7387 1445 7399 1497
rect 7451 1487 7755 1497
tri 7755 1487 7765 1497 sw
rect 7451 1481 7765 1487
tri 7765 1481 7771 1487 sw
rect 7451 1453 7771 1481
tri 7771 1453 7799 1481 sw
rect 7451 1451 7799 1453
rect 7451 1445 7457 1451
tri 7457 1445 7463 1451 nw
tri 7727 1445 7733 1451 ne
rect 7733 1445 7799 1451
tri 7799 1445 7807 1453 sw
rect 3265 1431 3328 1445
rect 3222 1423 3328 1431
tri 3328 1423 3350 1445 sw
tri 7733 1423 7755 1445 ne
rect 7755 1423 7807 1445
rect 3222 1411 3686 1423
rect 3222 1393 3643 1411
rect 3222 1359 3231 1393
rect 3265 1377 3643 1393
rect 3677 1377 3686 1411
rect 3265 1371 3686 1377
rect 3265 1365 3296 1371
tri 3296 1365 3302 1371 nw
tri 3606 1365 3612 1371 ne
rect 3612 1365 3686 1371
rect 3265 1359 3278 1365
rect 3222 1347 3278 1359
tri 3278 1347 3296 1365 nw
tri 3612 1347 3630 1365 ne
rect 3630 1347 3686 1365
rect 3222 1321 3274 1347
tri 3274 1343 3278 1347 nw
tri 3630 1343 3634 1347 ne
rect 3222 1287 3231 1321
rect 3265 1287 3274 1321
rect 3222 1248 3274 1287
rect 3222 1214 3231 1248
rect 3265 1214 3274 1248
rect 3222 1175 3274 1214
rect 3222 1141 3231 1175
rect 3265 1141 3274 1175
rect 3222 1102 3274 1141
rect 3222 1068 3231 1102
rect 3265 1068 3274 1102
rect 3222 1029 3274 1068
rect 3222 995 3231 1029
rect 3265 995 3274 1029
rect 3222 956 3274 995
rect 3222 922 3231 956
rect 3265 922 3274 956
rect 3222 883 3274 922
rect 3222 849 3231 883
rect 3265 849 3274 883
rect 3222 810 3274 849
rect 3222 776 3231 810
rect 3265 776 3274 810
rect 3222 737 3274 776
rect 3222 703 3231 737
rect 3265 703 3274 737
rect 3222 691 3274 703
rect 3474 1331 3526 1343
rect 3474 1297 3483 1331
rect 3517 1297 3526 1331
rect 3474 1256 3526 1297
rect 3474 1222 3483 1256
rect 3517 1222 3526 1256
rect 3474 1181 3526 1222
rect 3474 1147 3483 1181
rect 3517 1147 3526 1181
rect 3474 1105 3526 1147
rect 3474 1071 3483 1105
rect 3517 1071 3526 1105
rect 3474 1029 3526 1071
rect 3474 995 3483 1029
rect 3517 995 3526 1029
rect 3474 953 3526 995
rect 3474 919 3483 953
rect 3517 919 3526 953
rect 3474 877 3526 919
rect 3474 843 3483 877
rect 3517 843 3526 877
rect 3474 801 3526 843
rect 3474 767 3483 801
rect 3517 767 3526 801
rect 3474 725 3526 767
rect 3474 691 3483 725
rect 3517 691 3526 725
rect 3634 1337 3686 1347
rect 3634 1303 3643 1337
rect 3677 1303 3686 1337
rect 3634 1262 3686 1303
rect 3634 1228 3643 1262
rect 3677 1228 3686 1262
rect 3634 1187 3686 1228
rect 3634 1153 3643 1187
rect 3677 1153 3686 1187
rect 3634 1112 3686 1153
rect 3634 1078 3643 1112
rect 3677 1078 3686 1112
rect 3634 1037 3686 1078
rect 3634 1003 3643 1037
rect 3677 1003 3686 1037
rect 3634 962 3686 1003
rect 3634 928 3643 962
rect 3677 928 3686 962
rect 3634 887 3686 928
rect 3634 853 3643 887
rect 3677 853 3686 887
rect 3634 812 3686 853
rect 3634 778 3643 812
rect 3677 778 3686 812
rect 3634 737 3686 778
rect 3634 703 3643 737
rect 3677 703 3686 737
rect 3634 691 3686 703
rect 3750 1411 3802 1423
tri 7755 1415 7763 1423 ne
rect 7763 1415 7807 1423
tri 7807 1415 7837 1445 sw
tri 7763 1411 7767 1415 ne
rect 7767 1411 7837 1415
tri 7837 1411 7841 1415 sw
rect 3750 1377 3759 1411
rect 3793 1377 3802 1411
rect 3750 1337 3802 1377
rect 3750 1303 3759 1337
rect 3793 1303 3802 1337
rect 3750 1262 3802 1303
rect 3750 1228 3759 1262
rect 3793 1228 3802 1262
rect 3750 1187 3802 1228
rect 3750 1153 3759 1187
rect 3793 1153 3802 1187
rect 3750 1112 3802 1153
rect 3750 1078 3759 1112
rect 3793 1078 3802 1112
rect 3750 1037 3802 1078
rect 3750 1003 3759 1037
rect 3793 1003 3802 1037
rect 3750 962 3802 1003
rect 3750 928 3759 962
rect 3793 928 3802 962
rect 3750 887 3802 928
rect 3750 853 3759 887
rect 3793 853 3802 887
rect 3750 812 3802 853
rect 3750 778 3759 812
rect 3793 778 3802 812
rect 3750 737 3802 778
rect 3750 703 3759 737
rect 3793 703 3802 737
rect 3980 1405 4098 1411
tri 7767 1407 7771 1411 ne
rect 7771 1407 7841 1411
tri 7841 1407 7845 1411 sw
rect 3980 1353 3981 1405
rect 4033 1353 4045 1405
rect 4097 1353 4098 1405
tri 7771 1381 7797 1407 ne
rect 7797 1381 7845 1407
tri 7845 1381 7871 1407 sw
rect 3980 1340 4098 1353
tri 7797 1347 7831 1381 ne
rect 7831 1353 7871 1381
tri 7871 1353 7899 1381 sw
rect 7831 1347 7899 1353
tri 7899 1347 7905 1353 sw
rect 8185 1347 8418 1353
rect 3980 1288 3981 1340
rect 4033 1288 4045 1340
rect 4097 1288 4098 1340
tri 7831 1333 7845 1347 ne
rect 7845 1333 7905 1347
tri 7905 1333 7919 1347 sw
tri 7845 1313 7865 1333 ne
rect 7865 1313 7919 1333
tri 7919 1313 7939 1333 sw
rect 8185 1313 8197 1347
rect 8231 1313 8301 1347
tri 7865 1309 7869 1313 ne
rect 7869 1309 7939 1313
tri 7939 1309 7943 1313 sw
rect 3980 1275 4098 1288
tri 7869 1275 7903 1309 ne
rect 7903 1307 7943 1309
tri 7943 1307 7945 1309 sw
rect 8185 1307 8302 1313
rect 7903 1287 7945 1307
tri 7945 1287 7965 1307 sw
rect 7903 1275 7965 1287
tri 7965 1275 7977 1287 sw
rect 3980 1223 3981 1275
rect 4033 1223 4045 1275
rect 4097 1223 4098 1275
tri 7903 1259 7919 1275 ne
rect 7919 1259 7977 1275
tri 7977 1259 7993 1275 sw
rect 3980 1215 3986 1223
rect 4020 1215 4058 1223
rect 4092 1215 4098 1223
rect 3980 1210 4098 1215
rect 7919 1253 8049 1259
rect 7919 1219 7931 1253
rect 7965 1219 8003 1253
rect 8037 1219 8049 1253
rect 7919 1213 8049 1219
rect 3980 1158 3981 1210
rect 4033 1158 4045 1210
rect 4097 1158 4098 1210
tri 8160 1173 8185 1198 se
rect 8185 1173 8239 1197
rect 3980 1145 3986 1158
rect 4020 1145 4058 1158
rect 4092 1145 4098 1158
rect 3980 1093 3981 1145
rect 4033 1093 4045 1145
rect 4097 1093 4098 1145
rect 3980 1080 3986 1093
rect 4020 1080 4058 1093
rect 4092 1080 4098 1093
rect 3980 1028 3981 1080
rect 4033 1028 4045 1080
rect 4097 1028 4098 1080
rect 3980 1024 4098 1028
rect 3980 1015 3986 1024
rect 4020 1015 4058 1024
rect 4092 1015 4098 1024
rect 3980 963 3981 1015
rect 4033 963 4045 1015
rect 4097 963 4098 1015
rect 7857 1161 7903 1173
rect 7857 1127 7863 1161
rect 7897 1127 7903 1161
rect 7857 1085 7903 1127
rect 7857 1051 7863 1085
rect 7897 1051 7903 1085
rect 7857 1009 7903 1051
rect 3980 950 4098 963
rect 3980 898 3981 950
rect 4033 898 4045 950
rect 4097 898 4098 950
rect 3980 885 4098 898
rect 3980 833 3981 885
rect 4033 833 4045 885
rect 4097 833 4098 885
rect 6275 870 6281 986
rect 6461 870 6467 986
rect 7857 975 7863 1009
rect 7897 975 7903 1009
rect 7857 933 7903 975
rect 7857 899 7863 933
rect 7897 899 7903 933
rect 3980 820 4098 833
rect 3980 768 3981 820
rect 4033 768 4045 820
rect 4097 768 4098 820
rect 7857 857 7903 899
rect 7857 823 7863 857
rect 7897 823 7903 857
rect 3980 765 3986 768
rect 4020 765 4058 768
rect 4092 765 4098 768
rect 3980 754 4098 765
tri 2350 671 2358 679 sw
tri 2446 671 2454 679 se
rect 2454 671 2506 691
tri 2506 671 2514 679 sw
tri 2958 671 2966 679 se
rect 2966 671 3018 691
tri 3018 671 3026 679 sw
tri 3466 671 3474 679 se
rect 3474 678 3526 691
rect 3750 690 3802 703
tri 3802 690 3818 706 sw
rect 3980 702 3981 754
rect 4033 702 4045 754
rect 4097 702 4098 754
rect 3980 690 3986 702
rect 4020 690 4058 702
rect 4092 690 4098 702
rect 3750 685 3818 690
tri 3818 685 3823 690 sw
rect 3980 688 4098 690
rect 3750 681 3823 685
tri 3823 681 3827 685 sw
tri 3526 678 3529 681 sw
rect 3750 678 3827 681
tri 3827 678 3830 681 sw
rect 3474 671 3529 678
tri 3529 671 3536 678 sw
tri 3742 671 3749 678 se
tri 3749 675 3750 676 se
rect 3750 675 3830 678
rect 3749 671 3830 675
tri 3830 671 3837 678 sw
tri 2288 669 2290 671 se
rect 2290 669 2358 671
tri 2358 669 2360 671 sw
tri 2444 669 2446 671 se
rect 2446 669 2514 671
tri 2514 669 2516 671 sw
tri 2956 669 2958 671 se
rect 2958 669 3026 671
tri 3026 669 3028 671 sw
tri 3464 669 3466 671 se
rect 3466 669 3536 671
tri 3536 669 3538 671 sw
tri 3740 669 3742 671 se
rect 3742 669 3837 671
tri 3837 669 3839 671 sw
tri 2272 653 2288 669 se
rect 2288 653 2360 669
tri 2360 653 2376 669 sw
tri 2428 653 2444 669 se
rect 2444 653 2516 669
tri 2516 653 2532 669 sw
tri 2940 653 2956 669 se
rect 2956 653 3028 669
tri 3028 653 3044 669 sw
tri 3448 653 3464 669 se
rect 3464 653 3538 669
tri 3538 653 3554 669 sw
tri 3724 653 3740 669 se
rect 3740 653 3839 669
tri 3839 653 3855 669 sw
tri 2270 651 2272 653 se
rect 2272 651 2376 653
tri 2376 651 2378 653 sw
tri 2426 651 2428 653 se
rect 2428 651 2532 653
tri 2532 651 2534 653 sw
tri 2938 651 2940 653 se
rect 2940 651 3044 653
tri 3044 651 3046 653 sw
tri 3446 651 3448 653 se
rect 3448 651 3855 653
rect 2253 650 3855 651
tri 3855 650 3858 653 sw
rect 2253 649 3858 650
tri 3858 649 3859 650 sw
rect 2253 647 3859 649
rect 2253 531 3593 647
rect 3709 631 3859 647
tri 3859 631 3877 649 sw
rect 3709 531 3755 631
rect 2253 491 3755 531
rect 2253 457 2372 491
rect 2406 457 2445 491
rect 2479 457 2518 491
rect 2552 457 2591 491
rect 2625 457 2664 491
rect 2698 457 2737 491
rect 2771 457 2810 491
rect 2844 457 2882 491
rect 2916 457 2954 491
rect 2988 457 3026 491
rect 3060 457 3098 491
rect 3132 457 3170 491
rect 3204 457 3242 491
rect 3276 457 3314 491
rect 3348 457 3386 491
rect 3420 457 3458 491
rect 3492 457 3530 491
rect 3564 457 3602 491
rect 3636 457 3674 491
rect 3708 457 3746 491
rect 2253 451 3755 457
rect 3871 451 3877 631
rect 3980 636 3981 688
rect 4033 636 4045 688
rect 4097 636 4098 688
rect 7329 807 7381 813
rect 7329 743 7381 755
rect 7329 685 7381 691
tri 7329 679 7335 685 ne
rect 7335 679 7375 685
tri 7375 679 7381 685 nw
rect 7857 781 7903 823
rect 7857 747 7863 781
rect 7897 747 7903 781
rect 7857 705 7903 747
rect 3980 622 3986 636
rect 4020 622 4058 636
rect 4092 622 4098 636
rect 3980 570 3981 622
rect 4033 570 4045 622
rect 4097 570 4098 622
rect 3980 556 3986 570
rect 4020 556 4058 570
rect 4092 556 4098 570
rect 3980 504 3981 556
rect 4033 504 4045 556
rect 4097 504 4098 556
rect 3980 500 4098 504
rect 3980 490 3986 500
rect 4020 490 4058 500
rect 4092 490 4098 500
rect 3980 438 3981 490
rect 4033 438 4045 490
rect 4097 438 4098 490
rect 3980 426 4098 438
rect 3980 424 3986 426
rect 4020 424 4058 426
rect 4092 424 4098 426
rect 3980 372 3981 424
rect 4033 372 4045 424
rect 4097 372 4098 424
rect 3980 358 4098 372
tri 3963 294 3980 311 se
rect 3980 306 3981 358
rect 4033 306 4045 358
rect 4097 306 4098 358
rect 3980 294 4098 306
tri 3958 289 3963 294 se
rect 3963 292 4098 294
rect 3963 289 3981 292
tri 3955 286 3958 289 se
rect 3958 286 3981 289
tri 2208 280 2214 286 se
rect 2214 280 3981 286
tri 2174 246 2208 280 se
rect 2208 246 2226 280
rect 2260 246 2300 280
rect 2334 246 2373 280
rect 2407 246 2446 280
rect 2480 246 2519 280
rect 2553 246 2592 280
rect 2626 246 2665 280
rect 2699 246 2738 280
rect 2772 246 2811 280
rect 2845 246 2884 280
rect 2918 246 2957 280
rect 2991 246 3030 280
rect 3064 246 3103 280
rect 3137 246 3176 280
rect 3210 246 3249 280
rect 3283 246 3322 280
rect 3356 246 3395 280
rect 3429 246 3468 280
rect 3502 246 3541 280
rect 3575 246 3614 280
rect 3648 246 3687 280
rect 3721 246 3760 280
rect 3794 246 3833 280
rect 3867 246 3906 280
rect 3940 246 3979 280
tri 2153 225 2174 246 se
rect 2174 240 3981 246
rect 4033 240 4045 292
rect 4097 240 4098 292
rect 2174 226 4098 240
rect 2174 225 3981 226
tri 2147 219 2153 225 se
rect 2153 219 3981 225
tri 2145 217 2147 219 se
rect 2147 217 3981 219
tri 2142 214 2145 217 se
rect 2145 214 3981 217
rect 2142 208 3981 214
rect 2142 174 2226 208
rect 2260 174 2300 208
rect 2334 174 2373 208
rect 2407 174 2446 208
rect 2480 174 2519 208
rect 2553 174 2592 208
rect 2626 174 2665 208
rect 2699 174 2738 208
rect 2772 174 2811 208
rect 2845 174 2884 208
rect 2918 174 2957 208
rect 2991 174 3030 208
rect 3064 174 3103 208
rect 3137 174 3176 208
rect 3210 174 3249 208
rect 3283 174 3322 208
rect 3356 174 3395 208
rect 3429 174 3468 208
rect 3502 174 3541 208
rect 3575 174 3614 208
rect 3648 174 3687 208
rect 3721 174 3760 208
rect 3794 174 3833 208
rect 3867 174 3906 208
rect 3940 174 3979 208
rect 4033 174 4045 226
rect 4097 174 4098 226
rect 2142 168 4098 174
rect 7857 671 7863 705
rect 7897 671 7903 705
rect 7857 629 7903 671
rect 7857 595 7863 629
rect 7897 595 7903 629
rect 7857 553 7903 595
rect 7857 519 7863 553
rect 7897 519 7903 553
rect 7857 478 7903 519
rect 7857 444 7863 478
rect 7897 444 7903 478
rect 7857 403 7903 444
rect 7857 369 7863 403
rect 7897 369 7903 403
rect 7857 328 7903 369
rect 7857 294 7863 328
rect 7897 294 7903 328
rect 7857 253 7903 294
rect 7857 219 7863 253
rect 7897 219 7903 253
rect 7857 178 7903 219
rect 7857 144 7863 178
rect 7897 144 7903 178
rect 7857 119 7903 144
rect 7931 1161 8239 1173
rect 7931 1127 7979 1161
rect 8013 1127 8191 1161
rect 8225 1127 8239 1161
rect 7931 1088 8239 1127
rect 7931 1054 7979 1088
rect 8013 1063 8191 1088
rect 8013 1054 8035 1063
tri 8035 1054 8044 1063 nw
tri 8160 1054 8169 1063 ne
rect 8169 1054 8191 1063
rect 8225 1054 8239 1088
rect 7931 1053 8034 1054
tri 8034 1053 8035 1054 nw
tri 8169 1053 8170 1054 ne
rect 8170 1053 8239 1054
rect 7931 1015 8019 1053
tri 8019 1038 8034 1053 nw
tri 8170 1038 8185 1053 ne
rect 7931 981 7979 1015
rect 8013 981 8019 1015
rect 8185 1015 8239 1053
rect 7931 942 8019 981
rect 7931 908 7979 942
rect 8013 908 8019 942
rect 7931 869 8019 908
rect 7931 835 7979 869
rect 8013 835 8019 869
rect 7931 796 8019 835
rect 7931 762 7979 796
rect 8013 762 8019 796
rect 7931 723 8019 762
rect 7931 689 7979 723
rect 8013 689 8019 723
rect 7931 650 8019 689
rect 7931 616 7979 650
rect 8013 616 8019 650
rect 7931 577 8019 616
rect 7931 543 7979 577
rect 8013 543 8019 577
rect 7931 505 8019 543
rect 7931 471 7979 505
rect 8013 471 8019 505
rect 7931 433 8019 471
rect 7931 399 7979 433
rect 8013 399 8019 433
rect 7931 361 8019 399
rect 7931 327 7979 361
rect 8013 327 8019 361
rect 7931 289 8019 327
rect 7931 255 7979 289
rect 8013 255 8019 289
rect 7931 217 8019 255
rect 7931 183 7979 217
rect 8013 183 8019 217
rect 7931 141 8019 183
tri 7931 131 7941 141 ne
rect 7941 131 8019 141
rect 8079 995 8125 1007
rect 8079 961 8085 995
rect 8119 961 8125 995
rect 8079 922 8125 961
rect 8079 888 8085 922
rect 8119 888 8125 922
rect 8079 849 8125 888
rect 8079 815 8085 849
rect 8119 815 8125 849
rect 8079 776 8125 815
rect 8079 742 8085 776
rect 8119 742 8125 776
rect 8079 703 8125 742
rect 8079 669 8085 703
rect 8119 669 8125 703
rect 8079 631 8125 669
rect 8079 597 8085 631
rect 8119 597 8125 631
rect 8079 559 8125 597
rect 8079 525 8085 559
rect 8119 525 8125 559
rect 8079 487 8125 525
rect 8079 453 8085 487
rect 8119 453 8125 487
rect 8079 415 8125 453
rect 8079 381 8085 415
rect 8119 381 8125 415
rect 8079 343 8125 381
rect 8079 309 8085 343
rect 8119 309 8125 343
rect 8079 271 8125 309
rect 8079 237 8085 271
rect 8119 237 8125 271
tri 7903 119 7912 128 sw
rect 2253 57 3415 109
rect 3467 57 3481 109
rect 3533 57 3539 109
rect 7857 103 7912 119
tri 7912 103 7928 119 sw
rect 7857 69 7863 103
rect 7897 97 8051 103
rect 7897 69 8005 97
rect 7857 63 8005 69
rect 8039 63 8051 97
rect 7857 57 8051 63
rect 2253 -35 6748 17
rect 6800 -35 6814 17
rect 6866 -35 6872 17
rect 2253 -169 5026 -117
rect 5078 -169 5092 -117
rect 5144 -169 5150 -117
rect 8079 -131 8125 237
rect 8185 981 8191 1015
rect 8225 981 8239 1015
rect 8185 942 8239 981
rect 8185 908 8191 942
rect 8225 908 8239 942
rect 8185 869 8239 908
rect 8185 835 8191 869
rect 8225 835 8239 869
rect 8185 796 8239 835
rect 8185 762 8191 796
rect 8225 762 8239 796
rect 8185 723 8239 762
rect 8185 689 8191 723
rect 8225 689 8239 723
rect 8185 650 8239 689
rect 8185 616 8191 650
rect 8225 616 8239 650
rect 8185 577 8239 616
rect 8185 543 8191 577
rect 8225 543 8239 577
rect 8185 505 8239 543
rect 8185 471 8191 505
rect 8225 471 8239 505
rect 8185 433 8239 471
rect 8185 399 8191 433
rect 8225 399 8239 433
rect 8185 361 8239 399
rect 8185 327 8191 361
rect 8225 327 8239 361
rect 8185 289 8239 327
rect 8185 255 8191 289
rect 8225 255 8239 289
rect 8185 217 8239 255
tri 8158 183 8185 210 se
rect 8185 183 8191 217
rect 8225 183 8239 217
tri 8153 178 8158 183 se
rect 8158 178 8239 183
rect 8153 122 8239 178
rect 8301 1103 8302 1307
rect 8301 1093 8307 1103
rect 8341 1093 8418 1103
rect 8301 1090 8418 1093
rect 8301 1038 8302 1090
rect 8354 1038 8366 1090
rect 8301 1025 8307 1038
rect 8341 1025 8418 1038
rect 8301 973 8302 1025
rect 8354 973 8366 1025
rect 8301 960 8307 973
rect 8341 960 8418 973
rect 8301 908 8302 960
rect 8354 908 8366 960
rect 8301 906 8418 908
rect 8301 895 8307 906
rect 8341 895 8418 906
rect 8301 843 8302 895
rect 8354 843 8366 895
rect 8301 833 8418 843
rect 8301 830 8307 833
rect 8341 830 8418 833
rect 8301 778 8302 830
rect 8354 778 8366 830
rect 8301 765 8418 778
rect 8301 713 8302 765
rect 8354 713 8366 765
rect 8301 700 8418 713
rect 8301 648 8302 700
rect 8354 648 8366 700
rect 8301 635 8418 648
rect 8301 583 8302 635
rect 8354 583 8366 635
rect 8301 580 8307 583
rect 8341 580 8418 583
rect 8301 570 8418 580
rect 8301 518 8302 570
rect 8354 518 8366 570
rect 8301 507 8307 518
rect 8341 507 8418 518
rect 8301 505 8418 507
rect 8301 453 8302 505
rect 8354 453 8366 505
rect 8301 440 8307 453
rect 8341 440 8418 453
rect 8301 388 8302 440
rect 8354 388 8366 440
rect 8301 375 8307 388
rect 8341 375 8418 388
rect 8301 323 8302 375
rect 8354 323 8366 375
rect 8301 322 8418 323
rect 8301 310 8307 322
rect 8341 310 8418 322
rect 8301 258 8302 310
rect 8354 258 8366 310
rect 8301 249 8418 258
rect 8301 245 8307 249
rect 8341 245 8418 249
rect 8301 193 8302 245
rect 8354 193 8366 245
rect 8301 180 8418 193
rect 8301 128 8302 180
rect 8354 128 8366 180
rect 8301 115 8418 128
rect 8301 103 8302 115
rect 8153 97 8302 103
rect 8153 63 8165 97
rect 8199 63 8302 97
rect 8354 63 8366 115
rect 8153 57 8418 63
tri 8125 -131 8150 -106 sw
rect 8079 -143 8150 -131
tri 8150 -143 8162 -131 sw
rect 8079 -165 9142 -143
tri 8079 -169 8083 -165 ne
rect 8083 -169 9142 -165
tri 8083 -197 8111 -169 ne
rect 8111 -197 9142 -169
rect 2253 -249 7111 -197
rect 7163 -249 7177 -197
rect 7229 -249 7235 -197
tri 8111 -202 8116 -197 ne
rect 8116 -202 9142 -197
tri 9018 -203 9019 -202 ne
rect 9019 -203 9142 -202
tri 9019 -241 9057 -203 ne
rect 9057 -241 9142 -203
tri 9057 -249 9065 -241 ne
rect 9065 -249 9142 -241
tri 9065 -253 9069 -249 ne
tri 3590 -318 3593 -315 se
rect 3593 -318 3599 -315
rect 3590 -364 3599 -318
tri 3590 -367 3593 -364 ne
rect 3593 -367 3599 -364
rect 3651 -367 3663 -315
rect 3715 -367 3755 -315
rect 3807 -367 3819 -315
rect 3871 -318 3877 -315
tri 3877 -318 3880 -315 sw
rect 3871 -364 3880 -318
rect 3871 -367 3877 -364
tri 3877 -367 3880 -364 nw
rect 9069 -3049 9142 -249
tri 9142 -3049 9144 -3047 sw
rect 9069 -3059 9144 -3049
rect 9069 -3093 9087 -3059
rect 9121 -3076 9144 -3059
tri 9144 -3076 9171 -3049 sw
tri 9473 -3076 9500 -3049 se
rect 9500 -3076 9546 21862
tri 9546 21837 9571 21862 nw
tri 10227 21837 10252 21862 ne
rect 10252 21837 10324 21862
tri 10252 21829 10260 21837 ne
rect 10260 21829 10324 21837
tri 10260 21817 10272 21829 ne
rect 10272 21816 10324 21829
rect 10272 21765 10273 21815
rect 10274 21764 10322 21816
rect 10323 21765 10324 21815
tri 10250 21591 10272 21613 se
rect 10272 21591 10324 21764
tri 10241 21582 10250 21591 se
rect 10250 21582 10315 21591
tri 10315 21582 10324 21591 nw
rect 10765 21973 10771 22007
rect 10805 21973 10811 22007
rect 10765 21935 10811 21973
rect 10765 21901 10771 21935
rect 10805 21901 10811 21935
rect 10765 21863 10811 21901
rect 10765 21829 10771 21863
rect 10805 21829 10811 21863
rect 10765 21791 10811 21829
rect 10765 21757 10771 21791
rect 10805 21757 10811 21791
rect 10765 21719 10811 21757
rect 10765 21685 10771 21719
rect 10805 21685 10811 21719
rect 10765 21647 10811 21685
rect 10765 21613 10771 21647
rect 10805 21613 10811 21647
tri 10234 21575 10241 21582 se
rect 10241 21575 10308 21582
tri 10308 21575 10315 21582 nw
rect 10765 21575 10811 21613
tri 10200 21541 10234 21575 se
rect 10234 21541 10274 21575
tri 10274 21541 10308 21575 nw
rect 10765 21541 10771 21575
rect 10805 21541 10811 21575
tri 10167 21508 10200 21541 se
rect 10200 21508 10241 21541
tri 10241 21508 10274 21541 nw
tri 10162 21503 10167 21508 se
rect 10167 21503 10236 21508
tri 10236 21503 10241 21508 nw
rect 10765 21503 10811 21541
tri 10128 21469 10162 21503 se
rect 10162 21469 10202 21503
tri 10202 21469 10236 21503 nw
rect 10765 21469 10771 21503
rect 10805 21469 10811 21503
tri 10093 21434 10128 21469 se
rect 10128 21434 10167 21469
tri 10167 21434 10202 21469 nw
tri 10090 21431 10093 21434 se
rect 10093 21431 10164 21434
tri 10164 21431 10167 21434 nw
rect 10765 21431 10811 21469
tri 10056 21397 10090 21431 se
rect 10090 21397 10130 21431
tri 10130 21397 10164 21431 nw
rect 10765 21397 10771 21431
rect 10805 21397 10811 21431
tri 10019 21360 10056 21397 se
rect 10056 21360 10093 21397
tri 10093 21360 10130 21397 nw
tri 10018 21359 10019 21360 se
rect 10019 21359 10092 21360
tri 10092 21359 10093 21360 nw
rect 10765 21359 10811 21397
tri 9984 21325 10018 21359 se
rect 10018 21325 10058 21359
tri 10058 21325 10092 21359 nw
rect 10765 21325 10771 21359
rect 10805 21325 10811 21359
tri 9946 21287 9984 21325 se
rect 9984 21287 10020 21325
tri 10020 21287 10058 21325 nw
rect 10765 21287 10811 21325
tri 9945 21286 9946 21287 se
rect 9946 21286 10019 21287
tri 10019 21286 10020 21287 nw
tri 9912 21253 9945 21286 se
rect 9945 21253 9986 21286
tri 9986 21253 10019 21286 nw
rect 10765 21253 10771 21287
rect 10805 21253 10811 21287
tri 9893 21234 9912 21253 se
rect 9912 21234 9948 21253
rect 9893 21215 9948 21234
tri 9948 21215 9986 21253 nw
rect 10765 21215 10811 21253
rect 9893 12791 9945 21215
tri 9945 21212 9948 21215 nw
rect 10765 21181 10771 21215
rect 10805 21181 10811 21215
rect 10765 21143 10811 21181
rect 10765 21109 10771 21143
rect 10805 21109 10811 21143
rect 10765 21071 10811 21109
rect 10765 21037 10771 21071
rect 10805 21037 10811 21071
rect 10765 20999 10811 21037
rect 10765 20965 10771 20999
rect 10805 20965 10811 20999
rect 10765 20927 10811 20965
rect 10765 20893 10771 20927
rect 10805 20893 10811 20927
rect 10765 20855 10811 20893
rect 10765 20821 10771 20855
rect 10805 20821 10811 20855
rect 10765 20783 10811 20821
rect 10765 20749 10771 20783
rect 10805 20749 10811 20783
rect 10765 20711 10811 20749
rect 10765 20677 10771 20711
rect 10805 20677 10811 20711
rect 10765 20639 10811 20677
rect 10765 20605 10771 20639
rect 10805 20605 10811 20639
rect 10765 20567 10811 20605
rect 10765 20533 10771 20567
rect 10805 20533 10811 20567
rect 10765 20495 10811 20533
rect 10765 20461 10771 20495
rect 10805 20461 10811 20495
rect 10765 20423 10811 20461
rect 10765 20389 10771 20423
rect 10805 20389 10811 20423
rect 10765 20351 10811 20389
rect 10765 20317 10771 20351
rect 10805 20317 10811 20351
rect 10765 20279 10811 20317
rect 10765 20245 10771 20279
rect 10805 20245 10811 20279
rect 10765 20207 10811 20245
rect 10765 20173 10771 20207
rect 10805 20173 10811 20207
rect 10765 20135 10811 20173
rect 10765 20101 10771 20135
rect 10805 20101 10811 20135
rect 10765 20063 10811 20101
rect 10765 20029 10771 20063
rect 10805 20029 10811 20063
rect 10765 19991 10811 20029
rect 10765 19957 10771 19991
rect 10805 19957 10811 19991
rect 10765 19919 10811 19957
rect 10765 19885 10771 19919
rect 10805 19885 10811 19919
rect 10765 19847 10811 19885
rect 10765 19813 10771 19847
rect 10805 19813 10811 19847
rect 10765 19775 10811 19813
rect 10765 19741 10771 19775
rect 10805 19741 10811 19775
rect 10765 19703 10811 19741
rect 10765 19669 10771 19703
rect 10805 19669 10811 19703
rect 10765 19631 10811 19669
rect 10765 19597 10771 19631
rect 10805 19597 10811 19631
rect 10765 19559 10811 19597
rect 10765 19525 10771 19559
rect 10805 19525 10811 19559
rect 10765 19487 10811 19525
rect 10765 19453 10771 19487
rect 10805 19453 10811 19487
rect 10765 19415 10811 19453
rect 10765 19381 10771 19415
rect 10805 19381 10811 19415
rect 10765 19343 10811 19381
rect 10765 19309 10771 19343
rect 10805 19309 10811 19343
rect 10765 19271 10811 19309
rect 10765 19237 10771 19271
rect 10805 19237 10811 19271
rect 10765 19199 10811 19237
rect 10765 19165 10771 19199
rect 10805 19165 10811 19199
rect 10765 19127 10811 19165
rect 10765 19093 10771 19127
rect 10805 19093 10811 19127
rect 10765 19055 10811 19093
rect 10765 19021 10771 19055
rect 10805 19021 10811 19055
rect 10765 18983 10811 19021
rect 10765 18949 10771 18983
rect 10805 18949 10811 18983
rect 10765 18911 10811 18949
rect 10765 18877 10771 18911
rect 10805 18877 10811 18911
rect 10765 18839 10811 18877
rect 10765 18805 10771 18839
rect 10805 18805 10811 18839
rect 10765 18767 10811 18805
rect 10765 18733 10771 18767
rect 10805 18733 10811 18767
rect 10765 18695 10811 18733
rect 10765 18661 10771 18695
rect 10805 18661 10811 18695
rect 10765 18623 10811 18661
rect 10765 18589 10771 18623
rect 10805 18589 10811 18623
rect 10765 18551 10811 18589
rect 10765 18517 10771 18551
rect 10805 18517 10811 18551
rect 10765 18479 10811 18517
rect 10765 18445 10771 18479
rect 10805 18445 10811 18479
rect 10765 18407 10811 18445
rect 10765 18373 10771 18407
rect 10805 18373 10811 18407
rect 10765 18335 10811 18373
rect 10765 18301 10771 18335
rect 10805 18301 10811 18335
rect 10765 18263 10811 18301
rect 10765 18229 10771 18263
rect 10805 18229 10811 18263
rect 10765 18191 10811 18229
rect 10765 18157 10771 18191
rect 10805 18157 10811 18191
rect 10765 18119 10811 18157
rect 10765 18085 10771 18119
rect 10805 18085 10811 18119
rect 10765 18047 10811 18085
rect 10765 18013 10771 18047
rect 10805 18013 10811 18047
rect 10765 17975 10811 18013
rect 10765 17941 10771 17975
rect 10805 17941 10811 17975
rect 10765 17903 10811 17941
rect 10765 17869 10771 17903
rect 10805 17869 10811 17903
rect 10765 17831 10811 17869
rect 10765 17797 10771 17831
rect 10805 17797 10811 17831
rect 10765 17759 10811 17797
rect 10765 17725 10771 17759
rect 10805 17725 10811 17759
rect 10765 17687 10811 17725
rect 10765 17653 10771 17687
rect 10805 17653 10811 17687
rect 10765 17615 10811 17653
rect 10765 17581 10771 17615
rect 10805 17581 10811 17615
rect 10765 17543 10811 17581
rect 10765 17509 10771 17543
rect 10805 17509 10811 17543
rect 10765 17471 10811 17509
rect 10765 17437 10771 17471
rect 10805 17437 10811 17471
rect 10765 17399 10811 17437
rect 10765 17365 10771 17399
rect 10805 17365 10811 17399
rect 10765 17327 10811 17365
rect 10765 17293 10771 17327
rect 10805 17293 10811 17327
rect 10765 17255 10811 17293
rect 10765 17221 10771 17255
rect 10805 17221 10811 17255
rect 10765 17183 10811 17221
rect 10765 17149 10771 17183
rect 10805 17149 10811 17183
rect 10765 17111 10811 17149
rect 10765 17077 10771 17111
rect 10805 17077 10811 17111
rect 10765 17039 10811 17077
rect 10765 17005 10771 17039
rect 10805 17005 10811 17039
rect 10765 16967 10811 17005
rect 10765 16933 10771 16967
rect 10805 16933 10811 16967
rect 10765 16895 10811 16933
rect 10765 16861 10771 16895
rect 10805 16861 10811 16895
rect 10765 16823 10811 16861
rect 10765 16789 10771 16823
rect 10805 16789 10811 16823
rect 10765 16751 10811 16789
rect 10765 16717 10771 16751
rect 10805 16717 10811 16751
rect 10765 16679 10811 16717
rect 10765 16645 10771 16679
rect 10805 16645 10811 16679
rect 10765 16607 10811 16645
rect 10765 16573 10771 16607
rect 10805 16573 10811 16607
rect 10765 16535 10811 16573
rect 10765 16501 10771 16535
rect 10805 16501 10811 16535
rect 10765 16463 10811 16501
rect 10765 16429 10771 16463
rect 10805 16429 10811 16463
rect 10765 16391 10811 16429
rect 10765 16357 10771 16391
rect 10805 16357 10811 16391
rect 10765 16319 10811 16357
rect 10765 16285 10771 16319
rect 10805 16285 10811 16319
rect 10765 16247 10811 16285
rect 10765 16213 10771 16247
rect 10805 16213 10811 16247
rect 10765 16175 10811 16213
rect 10765 16141 10771 16175
rect 10805 16141 10811 16175
rect 10765 16103 10811 16141
rect 10765 16069 10771 16103
rect 10805 16069 10811 16103
rect 10765 16031 10811 16069
rect 10765 15997 10771 16031
rect 10805 15997 10811 16031
rect 10765 15959 10811 15997
rect 10765 15925 10771 15959
rect 10805 15925 10811 15959
rect 10765 15887 10811 15925
rect 10765 15853 10771 15887
rect 10805 15853 10811 15887
rect 10765 15815 10811 15853
rect 10765 15781 10771 15815
rect 10805 15781 10811 15815
rect 10765 15743 10811 15781
rect 10765 15709 10771 15743
rect 10805 15709 10811 15743
rect 10765 15671 10811 15709
rect 10765 15637 10771 15671
rect 10805 15637 10811 15671
rect 10765 15599 10811 15637
rect 10765 15565 10771 15599
rect 10805 15565 10811 15599
rect 10765 15527 10811 15565
rect 10765 15493 10771 15527
rect 10805 15493 10811 15527
rect 10765 15455 10811 15493
rect 10765 15421 10771 15455
rect 10805 15421 10811 15455
rect 10765 15383 10811 15421
rect 10765 15349 10771 15383
rect 10805 15349 10811 15383
rect 10765 15311 10811 15349
rect 10765 15277 10771 15311
rect 10805 15277 10811 15311
rect 10765 15239 10811 15277
rect 10765 15205 10771 15239
rect 10805 15205 10811 15239
rect 10765 15167 10811 15205
rect 10765 15133 10771 15167
rect 10805 15133 10811 15167
rect 10765 15095 10811 15133
rect 10765 15061 10771 15095
rect 10805 15061 10811 15095
rect 10765 15023 10811 15061
rect 10765 14989 10771 15023
rect 10805 14989 10811 15023
rect 10765 14951 10811 14989
rect 10765 14917 10771 14951
rect 10805 14917 10811 14951
rect 10765 14879 10811 14917
rect 10765 14845 10771 14879
rect 10805 14845 10811 14879
rect 10765 14807 10811 14845
rect 10765 14773 10771 14807
rect 10805 14773 10811 14807
rect 10765 14735 10811 14773
rect 10765 14701 10771 14735
rect 10805 14701 10811 14735
rect 10765 14663 10811 14701
rect 10765 14629 10771 14663
rect 10805 14629 10811 14663
rect 10765 14591 10811 14629
rect 10765 14557 10771 14591
rect 10805 14557 10811 14591
rect 10765 14519 10811 14557
rect 10765 14485 10771 14519
rect 10805 14485 10811 14519
rect 10765 14447 10811 14485
rect 10765 14413 10771 14447
rect 10805 14413 10811 14447
rect 10765 14375 10811 14413
rect 10765 14341 10771 14375
rect 10805 14341 10811 14375
rect 10765 14303 10811 14341
rect 10765 14269 10771 14303
rect 10805 14269 10811 14303
rect 10765 14231 10811 14269
rect 10765 14197 10771 14231
rect 10805 14197 10811 14231
rect 10765 14159 10811 14197
rect 10765 14125 10771 14159
rect 10805 14125 10811 14159
rect 10765 14087 10811 14125
rect 10765 14053 10771 14087
rect 10805 14053 10811 14087
rect 10765 14015 10811 14053
rect 10765 13981 10771 14015
rect 10805 13981 10811 14015
rect 10765 13943 10811 13981
rect 10765 13909 10771 13943
rect 10805 13909 10811 13943
rect 10765 13871 10811 13909
rect 10765 13837 10771 13871
rect 10805 13837 10811 13871
rect 10765 13799 10811 13837
rect 10765 13765 10771 13799
rect 10805 13765 10811 13799
rect 10765 13727 10811 13765
rect 10765 13693 10771 13727
rect 10805 13693 10811 13727
rect 10765 13655 10811 13693
rect 10765 13621 10771 13655
rect 10805 13621 10811 13655
rect 10765 13583 10811 13621
rect 10765 13549 10771 13583
rect 10805 13549 10811 13583
rect 10765 13511 10811 13549
rect 10765 13477 10771 13511
rect 10805 13477 10811 13511
rect 10765 13439 10811 13477
rect 10765 13405 10771 13439
rect 10805 13405 10811 13439
rect 10765 13367 10811 13405
rect 10765 13333 10771 13367
rect 10805 13333 10811 13367
rect 10765 13295 10811 13333
rect 10765 13261 10771 13295
rect 10805 13261 10811 13295
rect 10765 13223 10811 13261
rect 10765 13189 10771 13223
rect 10805 13189 10811 13223
rect 10765 13151 10811 13189
rect 10765 13117 10771 13151
rect 10805 13117 10811 13151
rect 10765 13079 10811 13117
rect 10765 13045 10771 13079
rect 10805 13045 10811 13079
rect 10765 13007 10811 13045
rect 10765 12973 10771 13007
rect 10805 12973 10811 13007
rect 10765 12935 10811 12973
rect 10765 12901 10771 12935
rect 10805 12901 10811 12935
rect 10765 12863 10811 12901
rect 10765 12829 10771 12863
rect 10805 12829 10811 12863
tri 9945 12791 9959 12805 sw
rect 10765 12791 10811 12829
rect 9893 12757 9959 12791
tri 9959 12757 9993 12791 sw
rect 10765 12757 10771 12791
rect 10805 12757 10811 12791
rect 9893 12754 9993 12757
tri 9993 12754 9996 12757 sw
rect 9893 12741 10265 12754
tri 10265 12741 10278 12754 sw
rect 9893 12719 10278 12741
tri 10278 12719 10300 12741 sw
rect 10765 12719 10811 12757
rect 9893 12708 10300 12719
tri 10300 12708 10311 12719 sw
rect 9893 12685 9973 12708
tri 9973 12685 9996 12708 nw
tri 10245 12685 10268 12708 ne
rect 10268 12695 10311 12708
tri 10311 12695 10324 12708 sw
rect 10268 12685 10324 12695
rect 9893 -1080 9945 12685
tri 9945 12657 9973 12685 nw
tri 10268 12675 10278 12685 ne
rect 10278 12627 10324 12685
rect 10278 12593 10284 12627
rect 10318 12593 10324 12627
rect 10278 12555 10324 12593
rect 10278 12521 10284 12555
rect 10318 12521 10324 12555
rect 10278 12509 10324 12521
rect 10765 12685 10771 12719
rect 10805 12685 10811 12719
rect 10765 12647 10811 12685
rect 10765 12613 10771 12647
rect 10805 12613 10811 12647
rect 10765 12575 10811 12613
rect 10765 12541 10771 12575
rect 10805 12541 10811 12575
rect 10765 12503 10811 12541
rect 10765 12469 10771 12503
rect 10805 12469 10811 12503
rect 10765 12431 10811 12469
rect 10765 12397 10771 12431
rect 10805 12397 10811 12431
rect 10765 12359 10811 12397
rect 10765 12325 10771 12359
rect 10805 12325 10811 12359
rect 10765 12287 10811 12325
rect 10765 12253 10771 12287
rect 10805 12253 10811 12287
rect 10765 12215 10811 12253
rect 10765 12181 10771 12215
rect 10805 12181 10811 12215
rect 10765 12143 10811 12181
rect 10765 12109 10771 12143
rect 10805 12109 10811 12143
rect 10765 12071 10811 12109
rect 10765 12037 10771 12071
rect 10805 12037 10811 12071
rect 10765 11999 10811 12037
rect 10765 11965 10771 11999
rect 10805 11965 10811 11999
rect 10765 11927 10811 11965
rect 10765 11893 10771 11927
rect 10805 11893 10811 11927
rect 10765 11855 10811 11893
rect 10765 11821 10771 11855
rect 10805 11821 10811 11855
rect 10765 11783 10811 11821
rect 10765 11749 10771 11783
rect 10805 11749 10811 11783
rect 10765 11711 10811 11749
rect 10765 11677 10771 11711
rect 10805 11677 10811 11711
rect 10765 11639 10811 11677
rect 10765 11605 10771 11639
rect 10805 11605 10811 11639
rect 10765 11567 10811 11605
rect 10765 11533 10771 11567
rect 10805 11533 10811 11567
rect 10765 11495 10811 11533
rect 10765 11461 10771 11495
rect 10805 11461 10811 11495
rect 10765 11423 10811 11461
rect 10765 11389 10771 11423
rect 10805 11389 10811 11423
rect 10765 11351 10811 11389
rect 10765 11317 10771 11351
rect 10805 11317 10811 11351
rect 10765 11279 10811 11317
rect 10765 11245 10771 11279
rect 10805 11245 10811 11279
rect 10765 11207 10811 11245
rect 10765 11173 10771 11207
rect 10805 11173 10811 11207
rect 10765 11135 10811 11173
rect 10765 11101 10771 11135
rect 10805 11101 10811 11135
rect 10765 11063 10811 11101
rect 10765 11029 10771 11063
rect 10805 11029 10811 11063
rect 10765 10991 10811 11029
rect 10765 10957 10771 10991
rect 10805 10957 10811 10991
rect 10765 10919 10811 10957
rect 10765 10885 10771 10919
rect 10805 10885 10811 10919
rect 10765 10847 10811 10885
rect 10765 10813 10771 10847
rect 10805 10813 10811 10847
rect 10765 10775 10811 10813
rect 10765 10741 10771 10775
rect 10805 10741 10811 10775
rect 10765 10703 10811 10741
rect 10765 10669 10771 10703
rect 10805 10669 10811 10703
rect 10765 10631 10811 10669
rect 10765 10597 10771 10631
rect 10805 10597 10811 10631
rect 10765 10559 10811 10597
rect 10765 10525 10771 10559
rect 10805 10525 10811 10559
rect 10765 10487 10811 10525
rect 10765 10453 10771 10487
rect 10805 10453 10811 10487
rect 10765 10415 10811 10453
rect 10765 10381 10771 10415
rect 10805 10381 10811 10415
rect 10765 10343 10811 10381
rect 10765 10309 10771 10343
rect 10805 10309 10811 10343
rect 10765 10271 10811 10309
rect 10765 10237 10771 10271
rect 10805 10237 10811 10271
rect 10765 10199 10811 10237
rect 10765 10165 10771 10199
rect 10805 10165 10811 10199
rect 10765 10127 10811 10165
rect 10765 10093 10771 10127
rect 10805 10093 10811 10127
rect 10765 10055 10811 10093
rect 10765 10021 10771 10055
rect 10805 10021 10811 10055
rect 10765 9983 10811 10021
rect 10765 9949 10771 9983
rect 10805 9949 10811 9983
rect 10765 9911 10811 9949
rect 10765 9877 10771 9911
rect 10805 9877 10811 9911
rect 10765 9839 10811 9877
rect 10765 9805 10771 9839
rect 10805 9805 10811 9839
rect 10765 9767 10811 9805
rect 10765 9733 10771 9767
rect 10805 9733 10811 9767
rect 10765 9695 10811 9733
rect 10765 9661 10771 9695
rect 10805 9661 10811 9695
rect 10765 9623 10811 9661
rect 10765 9589 10771 9623
rect 10805 9589 10811 9623
rect 10765 9551 10811 9589
rect 10765 9517 10771 9551
rect 10805 9517 10811 9551
rect 10765 9479 10811 9517
rect 10765 9445 10771 9479
rect 10805 9445 10811 9479
rect 10765 9407 10811 9445
rect 10765 9373 10771 9407
rect 10805 9373 10811 9407
rect 10765 9335 10811 9373
rect 10765 9301 10771 9335
rect 10805 9301 10811 9335
rect 10765 9263 10811 9301
rect 10765 9229 10771 9263
rect 10805 9229 10811 9263
rect 10765 9191 10811 9229
rect 10765 9157 10771 9191
rect 10805 9157 10811 9191
rect 10765 9119 10811 9157
rect 10765 9085 10771 9119
rect 10805 9085 10811 9119
rect 10765 9047 10811 9085
rect 10765 9013 10771 9047
rect 10805 9013 10811 9047
rect 10765 8975 10811 9013
rect 10765 8941 10771 8975
rect 10805 8941 10811 8975
rect 10765 8903 10811 8941
rect 10765 8869 10771 8903
rect 10805 8869 10811 8903
rect 10765 8831 10811 8869
rect 10765 8797 10771 8831
rect 10805 8797 10811 8831
rect 10765 8759 10811 8797
rect 10765 8725 10771 8759
rect 10805 8725 10811 8759
rect 10765 8687 10811 8725
rect 10765 8653 10771 8687
rect 10805 8653 10811 8687
rect 10765 8615 10811 8653
rect 10765 8581 10771 8615
rect 10805 8581 10811 8615
rect 10765 8543 10811 8581
rect 10765 8509 10771 8543
rect 10805 8509 10811 8543
rect 10765 8471 10811 8509
rect 10765 8437 10771 8471
rect 10805 8437 10811 8471
rect 10765 8399 10811 8437
rect 10765 8365 10771 8399
rect 10805 8365 10811 8399
rect 10765 8327 10811 8365
rect 10765 8293 10771 8327
rect 10805 8293 10811 8327
rect 10765 8255 10811 8293
rect 10765 8221 10771 8255
rect 10805 8221 10811 8255
rect 10765 8183 10811 8221
rect 10765 8149 10771 8183
rect 10805 8149 10811 8183
rect 10765 8111 10811 8149
rect 10765 8077 10771 8111
rect 10805 8077 10811 8111
rect 10765 8039 10811 8077
rect 10765 8005 10771 8039
rect 10805 8005 10811 8039
rect 10765 7967 10811 8005
rect 10765 7933 10771 7967
rect 10805 7933 10811 7967
rect 10765 7895 10811 7933
rect 10765 7861 10771 7895
rect 10805 7861 10811 7895
rect 10765 7823 10811 7861
rect 10765 7789 10771 7823
rect 10805 7789 10811 7823
rect 10765 7751 10811 7789
rect 10765 7717 10771 7751
rect 10805 7717 10811 7751
rect 10765 7679 10811 7717
rect 10765 7645 10771 7679
rect 10805 7645 10811 7679
rect 10765 7607 10811 7645
rect 10765 7573 10771 7607
rect 10805 7573 10811 7607
rect 10765 7535 10811 7573
rect 10765 7501 10771 7535
rect 10805 7501 10811 7535
rect 10765 7463 10811 7501
rect 10765 7429 10771 7463
rect 10805 7429 10811 7463
rect 10765 7391 10811 7429
rect 10765 7357 10771 7391
rect 10805 7357 10811 7391
rect 10765 7319 10811 7357
rect 10765 7285 10771 7319
rect 10805 7285 10811 7319
rect 10765 7247 10811 7285
rect 10765 7213 10771 7247
rect 10805 7213 10811 7247
rect 10765 7175 10811 7213
rect 10765 7141 10771 7175
rect 10805 7141 10811 7175
rect 10765 7103 10811 7141
rect 10765 7069 10771 7103
rect 10805 7069 10811 7103
rect 10765 7031 10811 7069
rect 10765 6997 10771 7031
rect 10805 6997 10811 7031
rect 10765 6959 10811 6997
rect 10765 6925 10771 6959
rect 10805 6925 10811 6959
rect 10765 6887 10811 6925
rect 10765 6853 10771 6887
rect 10805 6853 10811 6887
rect 10765 6815 10811 6853
rect 10765 6781 10771 6815
rect 10805 6781 10811 6815
rect 10765 6743 10811 6781
rect 10765 6709 10771 6743
rect 10805 6709 10811 6743
rect 10765 6671 10811 6709
rect 10765 6637 10771 6671
rect 10805 6637 10811 6671
rect 10765 6599 10811 6637
rect 10765 6565 10771 6599
rect 10805 6565 10811 6599
rect 10765 6527 10811 6565
rect 10765 6493 10771 6527
rect 10805 6493 10811 6527
rect 10765 6455 10811 6493
rect 10765 6421 10771 6455
rect 10805 6421 10811 6455
rect 10765 6383 10811 6421
rect 10765 6349 10771 6383
rect 10805 6349 10811 6383
rect 10765 6311 10811 6349
rect 10765 6277 10771 6311
rect 10805 6277 10811 6311
rect 10765 6239 10811 6277
rect 10765 6205 10771 6239
rect 10805 6205 10811 6239
rect 10765 6167 10811 6205
rect 10765 6133 10771 6167
rect 10805 6133 10811 6167
rect 10765 6095 10811 6133
rect 10765 6061 10771 6095
rect 10805 6061 10811 6095
rect 10765 6023 10811 6061
rect 10765 5989 10771 6023
rect 10805 5989 10811 6023
rect 10765 5951 10811 5989
rect 10765 5917 10771 5951
rect 10805 5917 10811 5951
rect 10765 5879 10811 5917
rect 10765 5845 10771 5879
rect 10805 5845 10811 5879
rect 10765 5807 10811 5845
rect 10765 5773 10771 5807
rect 10805 5773 10811 5807
rect 10765 5735 10811 5773
rect 10765 5701 10771 5735
rect 10805 5701 10811 5735
rect 10765 5663 10811 5701
rect 10765 5629 10771 5663
rect 10805 5629 10811 5663
rect 10765 5591 10811 5629
rect 10765 5557 10771 5591
rect 10805 5557 10811 5591
rect 10765 5519 10811 5557
rect 10765 5485 10771 5519
rect 10805 5485 10811 5519
rect 10765 5447 10811 5485
rect 10765 5413 10771 5447
rect 10805 5413 10811 5447
rect 10765 5375 10811 5413
rect 10765 5341 10771 5375
rect 10805 5341 10811 5375
rect 10765 5303 10811 5341
rect 10765 5269 10771 5303
rect 10805 5269 10811 5303
rect 10765 5231 10811 5269
rect 10765 5197 10771 5231
rect 10805 5197 10811 5231
rect 10765 5159 10811 5197
rect 10765 5125 10771 5159
rect 10805 5125 10811 5159
rect 10765 5087 10811 5125
rect 10765 5053 10771 5087
rect 10805 5053 10811 5087
rect 10765 5015 10811 5053
rect 10765 4981 10771 5015
rect 10805 4981 10811 5015
rect 10765 4943 10811 4981
rect 10765 4909 10771 4943
rect 10805 4909 10811 4943
rect 10765 4871 10811 4909
rect 10765 4837 10771 4871
rect 10805 4837 10811 4871
rect 10765 4799 10811 4837
rect 10765 4765 10771 4799
rect 10805 4765 10811 4799
rect 10765 4727 10811 4765
rect 10765 4693 10771 4727
rect 10805 4693 10811 4727
rect 10765 4655 10811 4693
rect 10765 4621 10771 4655
rect 10805 4621 10811 4655
rect 10765 4583 10811 4621
rect 10765 4549 10771 4583
rect 10805 4549 10811 4583
rect 10765 4511 10811 4549
rect 10765 4477 10771 4511
rect 10805 4477 10811 4511
rect 10765 4439 10811 4477
rect 10765 4405 10771 4439
rect 10805 4405 10811 4439
rect 10765 4367 10811 4405
rect 10765 4333 10771 4367
rect 10805 4333 10811 4367
rect 10765 4295 10811 4333
rect 10765 4261 10771 4295
rect 10805 4261 10811 4295
rect 10765 4223 10811 4261
rect 10765 4189 10771 4223
rect 10805 4189 10811 4223
rect 10765 4151 10811 4189
rect 10765 4117 10771 4151
rect 10805 4117 10811 4151
rect 10765 4079 10811 4117
rect 10765 4045 10771 4079
rect 10805 4045 10811 4079
rect 10765 4007 10811 4045
rect 10765 3973 10771 4007
rect 10805 3973 10811 4007
rect 10765 3935 10811 3973
rect 10765 3901 10771 3935
rect 10805 3901 10811 3935
rect 10765 3863 10811 3901
rect 10765 3829 10771 3863
rect 10805 3829 10811 3863
rect 10765 3791 10811 3829
rect 10765 3757 10771 3791
rect 10805 3757 10811 3791
rect 10765 3719 10811 3757
rect 10765 3685 10771 3719
rect 10805 3685 10811 3719
rect 10765 3647 10811 3685
rect 10765 3613 10771 3647
rect 10805 3613 10811 3647
rect 10765 3575 10811 3613
rect 10765 3541 10771 3575
rect 10805 3541 10811 3575
rect 10765 3503 10811 3541
rect 10765 3469 10771 3503
rect 10805 3469 10811 3503
rect 10765 3431 10811 3469
rect 10765 3397 10771 3431
rect 10805 3397 10811 3431
rect 10765 3359 10811 3397
rect 10765 3325 10771 3359
rect 10805 3325 10811 3359
rect 10765 3287 10811 3325
rect 10765 3253 10771 3287
rect 10805 3253 10811 3287
rect 10765 3215 10811 3253
rect 10765 3181 10771 3215
rect 10805 3181 10811 3215
rect 10765 3143 10811 3181
rect 10765 3109 10771 3143
rect 10805 3109 10811 3143
rect 10765 3071 10811 3109
rect 10765 3037 10771 3071
rect 10805 3037 10811 3071
rect 10765 2999 10811 3037
rect 10765 2965 10771 2999
rect 10805 2965 10811 2999
rect 10765 2927 10811 2965
rect 10765 2893 10771 2927
rect 10805 2893 10811 2927
rect 10765 2855 10811 2893
rect 10765 2821 10771 2855
rect 10805 2821 10811 2855
rect 10765 2783 10811 2821
rect 10765 2749 10771 2783
rect 10805 2749 10811 2783
rect 10765 2711 10811 2749
rect 10765 2677 10771 2711
rect 10805 2677 10811 2711
rect 10765 2639 10811 2677
rect 10765 2605 10771 2639
rect 10805 2605 10811 2639
rect 10765 2567 10811 2605
rect 10765 2533 10771 2567
rect 10805 2533 10811 2567
rect 10765 2495 10811 2533
rect 10765 2461 10771 2495
rect 10805 2461 10811 2495
rect 10765 2423 10811 2461
rect 10765 2389 10771 2423
rect 10805 2389 10811 2423
rect 10765 2351 10811 2389
rect 10765 2317 10771 2351
rect 10805 2317 10811 2351
rect 10765 2279 10811 2317
rect 10765 2245 10771 2279
rect 10805 2245 10811 2279
rect 10765 2207 10811 2245
rect 10765 2173 10771 2207
rect 10805 2173 10811 2207
rect 10765 2135 10811 2173
rect 10765 2101 10771 2135
rect 10805 2101 10811 2135
rect 10765 2063 10811 2101
rect 10765 2029 10771 2063
rect 10805 2029 10811 2063
rect 10765 1991 10811 2029
rect 10765 1957 10771 1991
rect 10805 1957 10811 1991
rect 10765 1919 10811 1957
rect 10765 1885 10771 1919
rect 10805 1885 10811 1919
rect 10765 1847 10811 1885
rect 10765 1813 10771 1847
rect 10805 1813 10811 1847
rect 10765 1775 10811 1813
rect 10765 1741 10771 1775
rect 10805 1741 10811 1775
rect 10765 1703 10811 1741
rect 10765 1669 10771 1703
rect 10805 1669 10811 1703
rect 9986 1644 10038 1650
rect 9986 1580 10038 1592
rect 9986 -702 10038 1528
rect 10765 1631 10811 1669
rect 10765 1597 10771 1631
rect 10805 1597 10811 1631
rect 10765 1559 10811 1597
rect 10765 1525 10771 1559
rect 10805 1525 10811 1559
rect 10765 1487 10811 1525
rect 10765 1453 10771 1487
rect 10805 1453 10811 1487
rect 10765 1415 10811 1453
rect 10765 1381 10771 1415
rect 10805 1381 10811 1415
rect 10765 1343 10811 1381
rect 10765 1309 10771 1343
rect 10805 1309 10811 1343
rect 10765 1271 10811 1309
rect 10765 1237 10771 1271
rect 10805 1237 10811 1271
rect 10765 1199 10811 1237
rect 10765 1165 10771 1199
rect 10805 1165 10811 1199
rect 10765 1127 10811 1165
rect 10765 1093 10771 1127
rect 10805 1093 10811 1127
rect 10765 1055 10811 1093
rect 10765 1021 10771 1055
rect 10805 1021 10811 1055
rect 10765 983 10811 1021
rect 10765 949 10771 983
rect 10805 949 10811 983
rect 10765 911 10811 949
rect 10765 877 10771 911
rect 10805 877 10811 911
rect 10765 839 10811 877
rect 10765 805 10771 839
rect 10805 805 10811 839
rect 10765 767 10811 805
rect 10765 733 10771 767
rect 10805 733 10811 767
rect 10765 695 10811 733
rect 10765 661 10771 695
rect 10805 661 10811 695
rect 10765 623 10811 661
rect 10765 589 10771 623
rect 10805 589 10811 623
rect 10765 551 10811 589
rect 10765 517 10771 551
rect 10805 517 10811 551
rect 10765 479 10811 517
rect 10765 445 10771 479
rect 10805 445 10811 479
rect 10765 407 10811 445
rect 10765 373 10771 407
rect 10805 373 10811 407
rect 10765 335 10811 373
rect 10765 301 10771 335
rect 10805 301 10811 335
rect 10765 263 10811 301
rect 10765 229 10771 263
rect 10805 229 10811 263
rect 10765 191 10811 229
rect 10765 157 10771 191
rect 10805 157 10811 191
rect 10765 119 10811 157
rect 10765 85 10771 119
rect 10805 85 10811 119
rect 10765 47 10811 85
rect 10765 13 10771 47
rect 10805 13 10811 47
rect 10765 -25 10811 13
rect 10765 -59 10771 -25
rect 10805 -59 10811 -25
rect 10765 -97 10811 -59
rect 10765 -131 10771 -97
rect 10805 -131 10811 -97
rect 10765 -169 10811 -131
rect 10765 -203 10771 -169
rect 10805 -203 10811 -169
rect 10765 -241 10811 -203
rect 10765 -275 10771 -241
rect 10805 -275 10811 -241
rect 10765 -313 10811 -275
rect 10765 -347 10771 -313
rect 10805 -347 10811 -313
rect 10765 -385 10811 -347
rect 10765 -419 10771 -385
rect 10805 -419 10811 -385
rect 10765 -457 10811 -419
rect 10765 -491 10771 -457
rect 10805 -491 10811 -457
rect 10765 -529 10811 -491
rect 10765 -563 10771 -529
rect 10805 -563 10811 -529
rect 10765 -601 10811 -563
rect 10765 -635 10771 -601
rect 10805 -635 10811 -601
rect 10765 -673 10811 -635
tri 9986 -707 9991 -702 ne
rect 9991 -707 10038 -702
tri 10038 -707 10065 -680 sw
rect 10765 -707 10771 -673
rect 10805 -707 10811 -673
tri 9991 -738 10022 -707 ne
rect 10022 -738 10065 -707
tri 10065 -738 10096 -707 sw
tri 10022 -745 10029 -738 ne
rect 10029 -745 10096 -738
tri 10096 -745 10103 -738 sw
rect 10765 -745 10811 -707
tri 10029 -754 10038 -745 ne
rect 10038 -754 10103 -745
tri 10038 -779 10063 -754 ne
rect 10063 -779 10103 -754
tri 10103 -779 10137 -745 sw
rect 10765 -779 10771 -745
rect 10805 -779 10811 -745
tri 10063 -812 10096 -779 ne
rect 10096 -812 10137 -779
tri 10137 -812 10170 -779 sw
tri 10096 -817 10101 -812 ne
rect 10101 -817 10170 -812
tri 10170 -817 10175 -812 sw
rect 10765 -817 10811 -779
tri 10101 -851 10135 -817 ne
rect 10135 -851 10175 -817
tri 10175 -851 10209 -817 sw
rect 10765 -851 10771 -817
rect 10805 -851 10811 -817
tri 10135 -886 10170 -851 ne
rect 10170 -886 10209 -851
tri 10209 -886 10244 -851 sw
tri 10170 -889 10173 -886 ne
rect 10173 -889 10244 -886
tri 10244 -889 10247 -886 sw
rect 10765 -889 10811 -851
tri 10173 -923 10207 -889 ne
rect 10207 -923 10247 -889
tri 10247 -923 10281 -889 sw
rect 10765 -923 10771 -889
rect 10805 -923 10811 -889
tri 10207 -960 10244 -923 ne
rect 10244 -960 10281 -923
tri 10281 -960 10318 -923 sw
tri 10244 -961 10245 -960 ne
rect 10245 -961 10318 -960
tri 10318 -961 10319 -960 sw
rect 10765 -961 10811 -923
tri 10245 -995 10279 -961 ne
rect 10279 -995 10319 -961
tri 10319 -995 10353 -961 sw
rect 10765 -995 10771 -961
rect 10805 -995 10811 -961
tri 10279 -1033 10317 -995 ne
rect 10317 -1033 10353 -995
tri 10353 -1033 10391 -995 sw
rect 10765 -1033 10811 -995
tri 10317 -1034 10318 -1033 ne
rect 10318 -1034 10391 -1033
tri 10391 -1034 10392 -1033 sw
tri 10318 -1067 10351 -1034 ne
rect 10351 -1067 10392 -1034
tri 10392 -1067 10425 -1034 sw
rect 10765 -1067 10771 -1033
rect 10805 -1067 10811 -1033
tri 10351 -1071 10355 -1067 ne
rect 10355 -1071 10425 -1067
tri 9945 -1080 9954 -1071 sw
tri 10355 -1080 10364 -1071 ne
rect 10364 -1080 10425 -1071
rect 9893 -1093 9954 -1080
tri 9893 -1105 9905 -1093 ne
rect 9905 -1105 9954 -1093
tri 9954 -1105 9979 -1080 sw
tri 10364 -1105 10389 -1080 ne
rect 10389 -1105 10425 -1080
tri 10425 -1105 10463 -1067 sw
rect 10765 -1105 10811 -1067
tri 9905 -1139 9939 -1105 ne
rect 9939 -1108 9979 -1105
tri 9979 -1108 9982 -1105 sw
tri 10389 -1108 10392 -1105 ne
rect 10392 -1108 10463 -1105
tri 10463 -1108 10466 -1105 sw
rect 9939 -1139 9982 -1108
tri 9982 -1139 10013 -1108 sw
tri 10392 -1139 10423 -1108 ne
rect 10423 -1139 10466 -1108
tri 10466 -1139 10497 -1108 sw
rect 10765 -1139 10771 -1105
rect 10805 -1139 10811 -1105
tri 9939 -1154 9954 -1139 ne
rect 9954 -1154 10013 -1139
tri 10013 -1154 10028 -1139 sw
tri 10423 -1154 10438 -1139 ne
rect 10438 -1154 10497 -1139
tri 9954 -1177 9977 -1154 ne
rect 9977 -1177 10028 -1154
tri 10028 -1177 10051 -1154 sw
tri 10438 -1177 10461 -1154 ne
rect 10461 -1177 10497 -1154
tri 10497 -1177 10535 -1139 sw
rect 10765 -1177 10811 -1139
tri 9977 -1211 10011 -1177 ne
rect 10011 -1182 10051 -1177
tri 10051 -1182 10056 -1177 sw
tri 10461 -1182 10466 -1177 ne
rect 10466 -1182 10535 -1177
tri 10535 -1182 10540 -1177 sw
rect 10011 -1211 10056 -1182
tri 10056 -1211 10085 -1182 sw
tri 10466 -1211 10495 -1182 ne
rect 10495 -1211 10540 -1182
tri 10540 -1211 10569 -1182 sw
rect 10765 -1211 10771 -1177
rect 10805 -1211 10811 -1177
tri 10011 -1228 10028 -1211 ne
rect 10028 -1228 10085 -1211
tri 10085 -1228 10102 -1211 sw
tri 10495 -1228 10512 -1211 ne
rect 10512 -1228 10569 -1211
tri 10028 -1249 10049 -1228 ne
rect 10049 -1249 10102 -1228
tri 10102 -1249 10123 -1228 sw
tri 10512 -1249 10533 -1228 ne
rect 10533 -1249 10569 -1228
tri 10569 -1249 10607 -1211 sw
rect 10765 -1249 10811 -1211
tri 10049 -1283 10083 -1249 ne
rect 10083 -1256 10123 -1249
tri 10123 -1256 10130 -1249 sw
tri 10533 -1256 10540 -1249 ne
rect 10540 -1256 10607 -1249
tri 10607 -1256 10614 -1249 sw
rect 10083 -1283 10130 -1256
tri 10130 -1283 10157 -1256 sw
tri 10540 -1283 10567 -1256 ne
rect 10567 -1283 10614 -1256
tri 10614 -1283 10641 -1256 sw
rect 10765 -1283 10771 -1249
rect 10805 -1283 10811 -1249
tri 10083 -1302 10102 -1283 ne
rect 10102 -1302 10157 -1283
tri 10157 -1302 10176 -1283 sw
tri 10567 -1302 10586 -1283 ne
rect 10586 -1302 10641 -1283
tri 10102 -1321 10121 -1302 ne
rect 10121 -1321 10176 -1302
tri 10176 -1321 10195 -1302 sw
tri 10586 -1321 10605 -1302 ne
rect 10605 -1321 10641 -1302
tri 10641 -1321 10679 -1283 sw
rect 10765 -1321 10811 -1283
tri 10121 -1355 10155 -1321 ne
rect 10155 -1330 10195 -1321
tri 10195 -1330 10204 -1321 sw
tri 10605 -1330 10614 -1321 ne
rect 10614 -1330 10679 -1321
tri 10679 -1330 10688 -1321 sw
rect 10155 -1352 10204 -1330
tri 10204 -1352 10226 -1330 sw
tri 10614 -1352 10636 -1330 ne
rect 10155 -1355 10226 -1352
tri 10226 -1355 10229 -1352 sw
tri 10155 -1376 10176 -1355 ne
rect 10176 -1376 10229 -1355
tri 10229 -1376 10250 -1355 sw
tri 10176 -1393 10193 -1376 ne
rect 10193 -1393 10250 -1376
tri 10250 -1393 10267 -1376 sw
tri 10193 -1427 10227 -1393 ne
rect 10227 -1427 10267 -1393
tri 10267 -1427 10301 -1393 sw
tri 10227 -1450 10250 -1427 ne
rect 10250 -1450 10301 -1427
tri 10301 -1450 10324 -1427 sw
tri 10250 -1465 10265 -1450 ne
rect 10265 -1465 10324 -1450
tri 10265 -1472 10272 -1465 ne
rect 10272 -1589 10324 -1465
rect 10431 -1555 10497 -1536
tri 10324 -1589 10327 -1586 sw
rect 10431 -1589 10446 -1555
rect 10480 -1589 10497 -1555
rect 10272 -1590 10327 -1589
tri 10327 -1590 10328 -1589 sw
rect 10272 -1597 10328 -1590
tri 10328 -1597 10335 -1590 sw
rect 10272 -1609 10335 -1597
tri 10335 -1609 10347 -1597 sw
tri 10419 -1609 10431 -1597 se
rect 10431 -1600 10497 -1589
rect 10636 -1556 10688 -1330
rect 10636 -1590 10642 -1556
rect 10676 -1590 10688 -1556
tri 10497 -1600 10500 -1597 sw
rect 10431 -1609 10500 -1600
tri 10500 -1609 10509 -1600 sw
tri 10627 -1609 10636 -1600 se
rect 10636 -1609 10688 -1590
rect 10272 -1622 10347 -1609
tri 10347 -1622 10360 -1609 sw
tri 10406 -1622 10419 -1609 se
rect 10419 -1622 10509 -1609
tri 10509 -1622 10522 -1609 sw
tri 10614 -1622 10627 -1609 se
rect 10627 -1622 10688 -1609
rect 10272 -1627 10573 -1622
rect 10272 -1661 10446 -1627
rect 10480 -1661 10573 -1627
rect 10272 -1674 10573 -1661
rect 10574 -1673 10575 -1623
rect 10611 -1673 10612 -1623
rect 10613 -1628 10688 -1622
rect 10613 -1662 10642 -1628
rect 10676 -1662 10688 -1628
rect 10613 -1674 10688 -1662
rect 10765 -1355 10771 -1321
rect 10805 -1355 10811 -1321
rect 10765 -1393 10811 -1355
rect 10765 -1427 10771 -1393
rect 10805 -1427 10811 -1393
rect 10765 -1465 10811 -1427
rect 10765 -1499 10771 -1465
rect 10805 -1499 10811 -1465
rect 10765 -1537 10811 -1499
rect 10765 -1571 10771 -1537
rect 10805 -1571 10811 -1537
rect 10765 -1609 10811 -1571
rect 10765 -1643 10771 -1609
rect 10805 -1643 10811 -1609
rect 9121 -3093 9194 -3076
rect 9069 -3128 9194 -3093
rect 9195 -3127 9196 -3077
rect 9232 -3127 9233 -3077
rect 9234 -3109 9367 -3076
rect 9234 -3128 9277 -3109
rect 9069 -3131 9156 -3128
rect 9069 -3165 9087 -3131
rect 9121 -3143 9156 -3131
tri 9156 -3143 9171 -3128 nw
tri 9238 -3143 9253 -3128 ne
rect 9253 -3143 9277 -3128
rect 9311 -3128 9367 -3109
rect 9368 -3127 9369 -3077
rect 9405 -3127 9406 -3077
rect 9407 -3128 9546 -3076
rect 10765 -1681 10811 -1643
rect 10765 -1715 10771 -1681
rect 10805 -1715 10811 -1681
rect 10765 -1753 10811 -1715
rect 10765 -1787 10771 -1753
rect 10805 -1787 10811 -1753
rect 10765 -1825 10811 -1787
rect 10765 -1859 10771 -1825
rect 10805 -1859 10811 -1825
rect 10765 -1897 10811 -1859
rect 10765 -1931 10771 -1897
rect 10805 -1931 10811 -1897
rect 10765 -1969 10811 -1931
rect 10765 -2003 10771 -1969
rect 10805 -2003 10811 -1969
rect 10765 -2041 10811 -2003
rect 10765 -2075 10771 -2041
rect 10805 -2075 10811 -2041
rect 10765 -2113 10811 -2075
rect 10765 -2147 10771 -2113
rect 10805 -2147 10811 -2113
rect 10765 -2185 10811 -2147
rect 10765 -2219 10771 -2185
rect 10805 -2219 10811 -2185
rect 10765 -2257 10811 -2219
rect 10765 -2291 10771 -2257
rect 10805 -2291 10811 -2257
rect 10765 -2329 10811 -2291
rect 10765 -2363 10771 -2329
rect 10805 -2363 10811 -2329
rect 10765 -2401 10811 -2363
rect 10765 -2435 10771 -2401
rect 10805 -2435 10811 -2401
rect 10765 -2473 10811 -2435
rect 10765 -2507 10771 -2473
rect 10805 -2507 10811 -2473
rect 10765 -2545 10811 -2507
rect 10765 -2579 10771 -2545
rect 10805 -2579 10811 -2545
rect 10765 -2617 10811 -2579
rect 10765 -2651 10771 -2617
rect 10805 -2651 10811 -2617
rect 10765 -2689 10811 -2651
rect 10765 -2723 10771 -2689
rect 10805 -2723 10811 -2689
rect 10765 -2761 10811 -2723
rect 10765 -2795 10771 -2761
rect 10805 -2795 10811 -2761
rect 10765 -2833 10811 -2795
rect 10765 -2867 10771 -2833
rect 10805 -2867 10811 -2833
rect 10765 -2905 10811 -2867
rect 10765 -2939 10771 -2905
rect 10805 -2939 10811 -2905
rect 10765 -2977 10811 -2939
rect 10765 -3011 10771 -2977
rect 10805 -3011 10811 -2977
rect 10765 -3049 10811 -3011
rect 10765 -3083 10771 -3049
rect 10805 -3083 10811 -3049
rect 10765 -3121 10811 -3083
rect 9311 -3143 9321 -3128
rect 9121 -3155 9144 -3143
tri 9144 -3155 9156 -3143 nw
tri 9253 -3155 9265 -3143 ne
rect 9265 -3155 9321 -3143
tri 9321 -3155 9348 -3128 nw
rect 10765 -3155 10771 -3121
rect 10805 -3155 10811 -3121
rect 9121 -3165 9142 -3155
tri 9142 -3157 9144 -3155 nw
tri 9265 -3157 9267 -3155 ne
rect 9267 -3157 9317 -3155
tri 9267 -3159 9269 -3157 ne
rect 9269 -3159 9317 -3157
tri 9317 -3159 9321 -3155 nw
tri 9269 -3161 9271 -3159 ne
rect 9069 -3177 9142 -3165
rect 9271 -3181 9317 -3159
rect 9271 -3215 9277 -3181
rect 9311 -3215 9317 -3181
rect 9271 -3227 9317 -3215
rect 10765 -3193 10811 -3155
rect 10765 -3227 10771 -3193
rect 10805 -3227 10811 -3193
rect 10765 -3265 10811 -3227
rect 10765 -3299 10771 -3265
rect 10805 -3299 10811 -3265
rect 10765 -3337 10811 -3299
rect 10765 -3371 10771 -3337
rect 10805 -3371 10811 -3337
rect 10765 -3409 10811 -3371
rect 10765 -3443 10771 -3409
rect 10805 -3443 10811 -3409
rect 10765 -3481 10811 -3443
rect 10765 -3515 10771 -3481
rect 10805 -3515 10811 -3481
rect 10765 -3553 10811 -3515
rect 10765 -3587 10771 -3553
rect 10805 -3587 10811 -3553
rect 10765 -3625 10811 -3587
rect 10765 -3659 10771 -3625
rect 10805 -3659 10811 -3625
rect 10765 -3697 10811 -3659
rect 10765 -3731 10771 -3697
rect 10805 -3731 10811 -3697
rect 10765 -3769 10811 -3731
rect 10765 -3803 10771 -3769
rect 10805 -3803 10811 -3769
rect 9169 -3835 9339 -3818
rect 9169 -3869 9221 -3835
rect 9255 -3869 9293 -3835
rect 9327 -3869 9339 -3835
rect 9169 -3886 9339 -3869
tri 9169 -3913 9196 -3886 ne
rect 9196 -3913 9312 -3886
tri 9312 -3913 9339 -3886 nw
rect 10765 -3841 10811 -3803
rect 10765 -3875 10771 -3841
rect 10805 -3875 10811 -3841
rect 10765 -3913 10811 -3875
tri 9196 -3947 9230 -3913 ne
rect 9230 -3947 9299 -3913
tri 9299 -3926 9312 -3913 nw
tri 9230 -3948 9231 -3947 ne
rect 9231 -5857 9299 -3947
rect 10765 -3947 10771 -3913
rect 10805 -3947 10811 -3913
rect 10765 -3985 10811 -3947
rect 10765 -4019 10771 -3985
rect 10805 -4019 10811 -3985
rect 10765 -4057 10811 -4019
rect 10765 -4091 10771 -4057
rect 10805 -4091 10811 -4057
rect 10765 -4129 10811 -4091
rect 10765 -4163 10771 -4129
rect 10805 -4163 10811 -4129
rect 10765 -4201 10811 -4163
rect 10765 -4235 10771 -4201
rect 10805 -4235 10811 -4201
rect 10765 -4273 10811 -4235
rect 10765 -4307 10771 -4273
rect 10805 -4307 10811 -4273
rect 10765 -4345 10811 -4307
rect 10765 -4379 10771 -4345
rect 10805 -4379 10811 -4345
rect 10765 -4417 10811 -4379
rect 10765 -4451 10771 -4417
rect 10805 -4451 10811 -4417
rect 10765 -4489 10811 -4451
rect 10765 -4523 10771 -4489
rect 10805 -4523 10811 -4489
rect 10765 -4561 10811 -4523
rect 10765 -4595 10771 -4561
rect 10805 -4595 10811 -4561
rect 10765 -4633 10811 -4595
rect 10765 -4667 10771 -4633
rect 10805 -4667 10811 -4633
rect 10765 -4705 10811 -4667
rect 10765 -4739 10771 -4705
rect 10805 -4739 10811 -4705
rect 10765 -4777 10811 -4739
rect 10765 -4811 10771 -4777
rect 10805 -4811 10811 -4777
rect 10765 -4849 10811 -4811
rect 10765 -4883 10771 -4849
rect 10805 -4883 10811 -4849
rect 10765 -4921 10811 -4883
rect 10765 -4955 10771 -4921
rect 10805 -4955 10811 -4921
rect 10765 -4993 10811 -4955
rect 10765 -5027 10771 -4993
rect 10805 -5027 10811 -4993
rect 10765 -5065 10811 -5027
rect 10765 -5099 10771 -5065
rect 10805 -5099 10811 -5065
rect 10765 -5137 10811 -5099
rect 10765 -5171 10771 -5137
rect 10805 -5171 10811 -5137
rect 10765 -5209 10811 -5171
rect 10765 -5243 10771 -5209
rect 10805 -5243 10811 -5209
rect 10765 -5281 10811 -5243
rect 10765 -5315 10771 -5281
rect 10805 -5315 10811 -5281
rect 10765 -5353 10811 -5315
rect 10765 -5387 10771 -5353
rect 10805 -5387 10811 -5353
rect 10765 -5425 10811 -5387
rect 10765 -5459 10771 -5425
rect 10805 -5459 10811 -5425
rect 10765 -5497 10811 -5459
rect 10765 -5531 10771 -5497
rect 10805 -5531 10811 -5497
rect 10765 -5569 10811 -5531
rect 10765 -5603 10771 -5569
rect 10805 -5603 10811 -5569
rect 10765 -5641 10811 -5603
rect 10765 -5675 10771 -5641
rect 10805 -5675 10811 -5641
rect 10765 -5713 10811 -5675
rect 10765 -5747 10771 -5713
rect 10805 -5747 10811 -5713
rect 10765 -5785 10811 -5747
rect 10765 -5819 10771 -5785
rect 10805 -5819 10811 -5785
tri 9299 -5857 9321 -5835 sw
rect 10765 -5857 10811 -5819
rect 9231 -5891 9321 -5857
tri 9321 -5891 9355 -5857 sw
rect 10765 -5891 10771 -5857
rect 10805 -5891 10811 -5857
rect 9231 -5904 9355 -5891
tri 9355 -5904 9368 -5891 sw
rect 9231 -5916 9525 -5904
rect 9231 -5950 9477 -5916
rect 9511 -5950 9525 -5916
rect 9231 -5988 9525 -5950
rect 9231 -6022 9477 -5988
rect 9511 -6022 9525 -5988
rect 9231 -6034 9525 -6022
rect 10765 -5929 10811 -5891
rect 10765 -5963 10771 -5929
rect 10805 -5963 10811 -5929
rect 10765 -6001 10811 -5963
rect 10765 -6035 10771 -6001
rect 10805 -6035 10811 -6001
rect 10765 -6073 10811 -6035
rect 10765 -6107 10771 -6073
rect 10805 -6107 10811 -6073
rect 10765 -6145 10811 -6107
rect 10765 -6179 10771 -6145
rect 10805 -6179 10811 -6145
rect 10765 -6217 10811 -6179
rect 10765 -6251 10771 -6217
rect 10805 -6251 10811 -6217
tri 10714 -6334 10765 -6283 se
rect 10765 -6334 10811 -6251
rect 10031 -6340 10811 -6334
rect 10031 -6374 10045 -6340
rect 10079 -6374 10117 -6340
rect 10151 -6374 10189 -6340
rect 10223 -6374 10261 -6340
rect 10295 -6374 10333 -6340
rect 10367 -6374 10405 -6340
rect 10439 -6374 10477 -6340
rect 10511 -6374 10549 -6340
rect 10583 -6374 10621 -6340
rect 10655 -6374 10693 -6340
rect 10727 -6374 10765 -6340
rect 10799 -6374 10811 -6340
rect 10031 -6380 10811 -6374
<< rmetal1 >>
rect 9719 21949 9721 21950
rect 9719 21899 9720 21949
rect 9719 21898 9721 21899
rect 9757 21949 9759 21950
rect 9758 21899 9759 21949
rect 10033 21949 10035 21950
rect 9757 21898 9759 21899
rect 10033 21899 10034 21949
rect 10033 21898 10035 21899
rect 10071 21949 10073 21950
rect 10072 21899 10073 21949
rect 10071 21898 10073 21899
rect 10272 21815 10274 21816
rect 10273 21765 10274 21815
rect 10272 21764 10274 21765
rect 10322 21815 10324 21816
rect 10322 21765 10323 21815
rect 10322 21764 10324 21765
rect 10573 -1623 10575 -1622
rect 10573 -1673 10574 -1623
rect 10573 -1674 10575 -1673
rect 10611 -1623 10613 -1622
rect 10612 -1673 10613 -1623
rect 10611 -1674 10613 -1673
rect 9194 -3077 9196 -3076
rect 9194 -3127 9195 -3077
rect 9194 -3128 9196 -3127
rect 9232 -3077 9234 -3076
rect 9233 -3127 9234 -3077
rect 9367 -3077 9369 -3076
rect 9232 -3128 9234 -3127
rect 9367 -3127 9368 -3077
rect 9367 -3128 9369 -3127
rect 9405 -3077 9407 -3076
rect 9406 -3127 9407 -3077
rect 9405 -3128 9407 -3127
<< via1 >>
rect 3987 2025 4103 2093
rect 3987 1991 4000 2025
rect 4000 1991 4034 2025
rect 4034 1991 4074 2025
rect 4074 1991 4103 2025
rect 3987 1953 4103 1991
rect 3987 1919 4000 1953
rect 4000 1919 4034 1953
rect 4034 1919 4074 1953
rect 4074 1919 4103 1953
rect 3987 1913 4103 1919
rect 3755 1719 3807 1725
rect 3755 1685 3759 1719
rect 3759 1685 3793 1719
rect 3793 1685 3807 1719
rect 3755 1673 3807 1685
rect 3819 1673 3871 1725
rect 9061 1598 9113 1650
rect 9125 1598 9177 1650
rect 7335 1445 7387 1497
rect 7399 1445 7451 1497
rect 3981 1399 4033 1405
rect 3981 1365 3986 1399
rect 3986 1365 4020 1399
rect 4020 1365 4033 1399
rect 3981 1353 4033 1365
rect 4045 1399 4097 1405
rect 4045 1365 4058 1399
rect 4058 1365 4092 1399
rect 4092 1365 4097 1399
rect 4045 1353 4097 1365
rect 3981 1324 4033 1340
rect 3981 1290 3986 1324
rect 3986 1290 4020 1324
rect 4020 1290 4033 1324
rect 3981 1288 4033 1290
rect 4045 1324 4097 1340
rect 4045 1290 4058 1324
rect 4058 1290 4092 1324
rect 4092 1290 4097 1324
rect 4045 1288 4097 1290
rect 8302 1313 8335 1347
rect 8335 1313 8418 1347
rect 3981 1249 4033 1275
rect 3981 1223 3986 1249
rect 3986 1223 4020 1249
rect 4020 1223 4033 1249
rect 4045 1249 4097 1275
rect 4045 1223 4058 1249
rect 4058 1223 4092 1249
rect 4092 1223 4097 1249
rect 3981 1174 4033 1210
rect 3981 1158 3986 1174
rect 3986 1158 4020 1174
rect 4020 1158 4033 1174
rect 4045 1174 4097 1210
rect 4045 1158 4058 1174
rect 4058 1158 4092 1174
rect 4092 1158 4097 1174
rect 3981 1140 3986 1145
rect 3986 1140 4020 1145
rect 4020 1140 4033 1145
rect 3981 1099 4033 1140
rect 3981 1093 3986 1099
rect 3986 1093 4020 1099
rect 4020 1093 4033 1099
rect 4045 1140 4058 1145
rect 4058 1140 4092 1145
rect 4092 1140 4097 1145
rect 4045 1099 4097 1140
rect 4045 1093 4058 1099
rect 4058 1093 4092 1099
rect 4092 1093 4097 1099
rect 3981 1065 3986 1080
rect 3986 1065 4020 1080
rect 4020 1065 4033 1080
rect 3981 1028 4033 1065
rect 4045 1065 4058 1080
rect 4058 1065 4092 1080
rect 4092 1065 4097 1080
rect 4045 1028 4097 1065
rect 3981 990 3986 1015
rect 3986 990 4020 1015
rect 4020 990 4033 1015
rect 3981 963 4033 990
rect 4045 990 4058 1015
rect 4058 990 4092 1015
rect 4092 990 4097 1015
rect 4045 963 4097 990
rect 3981 949 4033 950
rect 3981 915 3986 949
rect 3986 915 4020 949
rect 4020 915 4033 949
rect 3981 898 4033 915
rect 4045 949 4097 950
rect 4045 915 4058 949
rect 4058 915 4092 949
rect 4092 915 4097 949
rect 4045 898 4097 915
rect 3981 874 4033 885
rect 3981 840 3986 874
rect 3986 840 4020 874
rect 4020 840 4033 874
rect 3981 833 4033 840
rect 4045 874 4097 885
rect 4045 840 4058 874
rect 4058 840 4092 874
rect 4092 840 4097 874
rect 4045 833 4097 840
rect 6281 870 6461 986
rect 3981 799 4033 820
rect 3981 768 3986 799
rect 3986 768 4020 799
rect 4020 768 4033 799
rect 4045 799 4097 820
rect 4045 768 4058 799
rect 4058 768 4092 799
rect 4092 768 4097 799
rect 3981 724 4033 754
rect 3981 702 3986 724
rect 3986 702 4020 724
rect 4020 702 4033 724
rect 4045 724 4097 754
rect 4045 702 4058 724
rect 4058 702 4092 724
rect 4092 702 4097 724
rect 3593 531 3709 647
rect 3755 491 3871 631
rect 3755 457 3780 491
rect 3780 457 3871 491
rect 3755 451 3871 457
rect 3981 649 4033 688
rect 3981 636 3986 649
rect 3986 636 4020 649
rect 4020 636 4033 649
rect 4045 649 4097 688
rect 4045 636 4058 649
rect 4058 636 4092 649
rect 4092 636 4097 649
rect 7329 755 7381 807
rect 7329 691 7381 743
rect 3981 615 3986 622
rect 3986 615 4020 622
rect 4020 615 4033 622
rect 3981 574 4033 615
rect 3981 570 3986 574
rect 3986 570 4020 574
rect 4020 570 4033 574
rect 4045 615 4058 622
rect 4058 615 4092 622
rect 4092 615 4097 622
rect 4045 574 4097 615
rect 4045 570 4058 574
rect 4058 570 4092 574
rect 4092 570 4097 574
rect 3981 540 3986 556
rect 3986 540 4020 556
rect 4020 540 4033 556
rect 3981 504 4033 540
rect 4045 540 4058 556
rect 4058 540 4092 556
rect 4092 540 4097 556
rect 4045 504 4097 540
rect 3981 466 3986 490
rect 3986 466 4020 490
rect 4020 466 4033 490
rect 3981 438 4033 466
rect 4045 466 4058 490
rect 4058 466 4092 490
rect 4092 466 4097 490
rect 4045 438 4097 466
rect 3981 392 3986 424
rect 3986 392 4020 424
rect 4020 392 4033 424
rect 3981 372 4033 392
rect 4045 392 4058 424
rect 4058 392 4092 424
rect 4092 392 4097 424
rect 4045 372 4097 392
rect 3981 352 4033 358
rect 3981 318 3986 352
rect 3986 318 4020 352
rect 4020 318 4033 352
rect 3981 306 4033 318
rect 4045 352 4097 358
rect 4045 318 4058 352
rect 4058 318 4092 352
rect 4092 318 4097 352
rect 4045 306 4097 318
rect 3981 280 4033 292
rect 3981 246 4013 280
rect 4013 246 4033 280
rect 3981 240 4033 246
rect 4045 280 4097 292
rect 4045 246 4052 280
rect 4052 246 4086 280
rect 4086 246 4097 280
rect 4045 240 4097 246
rect 3981 208 4033 226
rect 3981 174 4013 208
rect 4013 174 4033 208
rect 4045 208 4097 226
rect 4045 174 4052 208
rect 4052 174 4086 208
rect 4086 174 4097 208
rect 3415 57 3467 109
rect 3481 57 3533 109
rect 6748 -35 6800 17
rect 6814 -35 6866 17
rect 5026 -169 5078 -117
rect 5092 -169 5144 -117
rect 8302 1275 8418 1313
rect 8302 1241 8307 1275
rect 8307 1241 8341 1275
rect 8341 1241 8418 1275
rect 8302 1201 8418 1241
rect 8302 1167 8307 1201
rect 8307 1167 8341 1201
rect 8341 1167 8418 1201
rect 8302 1127 8418 1167
rect 8302 1103 8307 1127
rect 8307 1103 8341 1127
rect 8341 1103 8418 1127
rect 8302 1053 8354 1090
rect 8302 1038 8307 1053
rect 8307 1038 8341 1053
rect 8341 1038 8354 1053
rect 8366 1038 8418 1090
rect 8302 1019 8307 1025
rect 8307 1019 8341 1025
rect 8341 1019 8354 1025
rect 8302 979 8354 1019
rect 8302 973 8307 979
rect 8307 973 8341 979
rect 8341 973 8354 979
rect 8366 973 8418 1025
rect 8302 945 8307 960
rect 8307 945 8341 960
rect 8341 945 8354 960
rect 8302 908 8354 945
rect 8366 908 8418 960
rect 8302 872 8307 895
rect 8307 872 8341 895
rect 8341 872 8354 895
rect 8302 843 8354 872
rect 8366 843 8418 895
rect 8302 799 8307 830
rect 8307 799 8341 830
rect 8341 799 8354 830
rect 8302 778 8354 799
rect 8366 778 8418 830
rect 8302 760 8354 765
rect 8302 726 8307 760
rect 8307 726 8341 760
rect 8341 726 8354 760
rect 8302 713 8354 726
rect 8366 713 8418 765
rect 8302 687 8354 700
rect 8302 653 8307 687
rect 8307 653 8341 687
rect 8341 653 8354 687
rect 8302 648 8354 653
rect 8366 648 8418 700
rect 8302 614 8354 635
rect 8302 583 8307 614
rect 8307 583 8341 614
rect 8341 583 8354 614
rect 8366 583 8418 635
rect 8302 541 8354 570
rect 8302 518 8307 541
rect 8307 518 8341 541
rect 8341 518 8354 541
rect 8366 518 8418 570
rect 8302 468 8354 505
rect 8302 453 8307 468
rect 8307 453 8341 468
rect 8341 453 8354 468
rect 8366 453 8418 505
rect 8302 434 8307 440
rect 8307 434 8341 440
rect 8341 434 8354 440
rect 8302 395 8354 434
rect 8302 388 8307 395
rect 8307 388 8341 395
rect 8341 388 8354 395
rect 8366 388 8418 440
rect 8302 361 8307 375
rect 8307 361 8341 375
rect 8341 361 8354 375
rect 8302 323 8354 361
rect 8366 323 8418 375
rect 8302 288 8307 310
rect 8307 288 8341 310
rect 8341 288 8354 310
rect 8302 258 8354 288
rect 8366 258 8418 310
rect 8302 215 8307 245
rect 8307 215 8341 245
rect 8341 215 8354 245
rect 8302 193 8354 215
rect 8366 193 8418 245
rect 8302 176 8354 180
rect 8302 142 8307 176
rect 8307 142 8341 176
rect 8341 142 8354 176
rect 8302 128 8354 142
rect 8366 128 8418 180
rect 8302 103 8354 115
rect 8302 69 8307 103
rect 8307 69 8341 103
rect 8341 69 8354 103
rect 8302 63 8354 69
rect 8366 63 8418 115
rect 7111 -249 7163 -197
rect 7177 -249 7229 -197
rect 3599 -367 3651 -315
rect 3663 -367 3715 -315
rect 3755 -367 3807 -315
rect 3819 -367 3871 -315
rect 9986 1592 10038 1644
rect 9986 1528 10038 1580
<< metal2 >>
rect -5926 -3990 -5606 -12
rect -4390 -35 -3565 -12
tri -3565 -35 -3542 -12 sw
rect -4390 -117 -3542 -35
tri -3542 -117 -3460 -35 sw
rect -4390 -169 -3460 -117
tri -3460 -169 -3408 -117 sw
rect -4390 -197 -3408 -169
tri -3408 -197 -3380 -169 sw
rect -4390 -222 -3380 -197
tri -3380 -222 -3355 -197 sw
rect -4390 -249 -3355 -222
tri -3355 -249 -3328 -222 sw
tri -898 -249 -881 -232 se
rect -881 -249 -751 -232
rect -4390 -315 -3328 -249
tri -3328 -315 -3262 -249 sw
tri -957 -308 -898 -249 se
rect -898 -308 -751 -249
tri 2309 -308 2322 -295 se
rect 2322 -308 2515 2076
rect -4390 -354 -3262 -315
tri -4390 -367 -4377 -354 ne
rect -4377 -367 -3262 -354
tri -3262 -367 -3210 -315 sw
tri -4377 -418 -4326 -367 ne
rect -4326 -418 -3210 -367
tri -3210 -418 -3159 -367 sw
rect -5224 -3614 -4414 -418
tri -4326 -1389 -3355 -418 ne
rect -3355 -1389 -3159 -418
tri -3159 -1389 -2188 -418 sw
tri -3355 -1731 -3013 -1389 ne
rect -3917 -3614 -3069 -1755
rect -3013 -3614 -2188 -1389
tri -2132 -1213 -2130 -1211 se
rect -2132 -1256 -1816 -1213
rect -2132 -3614 -1830 -1256
tri -1830 -1270 -1816 -1256 nw
rect -1620 -3210 -1428 -308
tri -964 -315 -957 -308 se
rect -957 -315 -751 -308
tri -1016 -367 -964 -315 se
rect -964 -367 -751 -315
tri -1067 -418 -1016 -367 se
rect -1016 -418 -751 -367
rect -1067 -1228 -751 -418
rect -734 -3614 -323 -1776
rect -185 -3614 7 -308
rect 303 -3614 355 -308
rect 395 -511 447 -308
rect 455 -3614 906 -1776
rect 996 -3614 1188 -308
rect 1518 -2984 1710 -308
tri 2302 -315 2309 -308 se
rect 2309 -315 2515 -308
tri 2250 -367 2302 -315 se
rect 2302 -367 2515 -315
tri 2199 -418 2250 -367 se
rect 2250 -418 2515 -367
rect 2199 -1228 2515 -418
rect 2643 -1605 2909 2076
tri 3481 128 3487 134 se
rect 3487 128 3539 2161
tri 3468 115 3481 128 se
rect 3481 115 3539 128
tri 3462 109 3468 115 se
rect 3468 109 3539 115
rect 3409 57 3415 109
rect 3467 57 3481 109
rect 3533 57 3539 109
rect 3593 647 3721 2104
rect 3709 531 3721 647
rect 2643 -1677 2837 -1605
tri 2837 -1677 2909 -1605 nw
rect 3593 -315 3721 531
rect 3593 -367 3599 -315
rect 3651 -367 3663 -315
rect 3715 -367 3721 -315
rect 3593 -1324 3721 -367
rect 3749 1725 3877 2104
rect 3749 1673 3755 1725
rect 3807 1673 3819 1725
rect 3871 1673 3877 1725
rect 3749 631 3877 1673
rect 3749 451 3755 631
rect 3871 451 3877 631
rect 3749 -315 3877 451
rect 3981 2093 4109 2104
rect 3981 1913 3987 2093
rect 4103 1913 4109 2093
rect 3981 1405 4109 1913
rect 4033 1353 4045 1405
rect 4097 1353 4109 1405
rect 3981 1340 4109 1353
rect 4033 1288 4045 1340
rect 4097 1288 4109 1340
rect 3981 1275 4109 1288
rect 4033 1223 4045 1275
rect 4097 1223 4109 1275
rect 3981 1210 4109 1223
rect 4033 1158 4045 1210
rect 4097 1158 4109 1210
rect 3981 1145 4109 1158
rect 4033 1093 4045 1145
rect 4097 1093 4109 1145
rect 3981 1080 4109 1093
rect 4033 1028 4045 1080
rect 4097 1028 4109 1080
rect 3981 1015 4109 1028
rect 4033 963 4045 1015
rect 4097 963 4109 1015
rect 3981 950 4109 963
rect 4033 898 4045 950
rect 4097 898 4109 950
rect 3981 885 4109 898
rect 4033 833 4045 885
rect 4097 833 4109 885
rect 3981 820 4109 833
rect 4033 768 4045 820
rect 4097 768 4109 820
rect 3981 754 4109 768
rect 4033 702 4045 754
rect 4097 702 4109 754
rect 3981 688 4109 702
rect 4033 636 4045 688
rect 4097 636 4109 688
rect 3981 622 4109 636
rect 4033 570 4045 622
rect 4097 570 4109 622
rect 3981 556 4109 570
rect 4033 504 4045 556
rect 4097 504 4109 556
rect 3981 490 4109 504
rect 4033 438 4045 490
rect 4097 438 4109 490
rect 3981 424 4109 438
rect 4033 372 4045 424
rect 4097 372 4109 424
rect 3981 358 4109 372
rect 4033 306 4045 358
rect 4097 306 4109 358
rect 3981 292 4109 306
rect 4033 240 4045 292
rect 4097 240 4109 292
rect 3981 226 4109 240
rect 4033 174 4045 226
rect 4097 174 4109 226
rect 3981 168 4109 174
tri 4399 -315 4419 -295 se
rect 4419 -315 4612 2076
tri 5073 -117 5098 -92 se
rect 5098 -117 5150 2161
tri 5772 2135 5797 2160 sw
rect 5020 -169 5026 -117
rect 5078 -169 5092 -117
rect 5144 -169 5150 -117
tri 5644 -169 5772 -41 se
rect 5772 -169 6205 2135
rect 6261 1027 6483 2161
tri 6993 1362 7068 1437 se
rect 7068 1414 7120 2161
tri 7068 1362 7120 1414 nw
tri 6978 1347 6993 1362 se
rect 6993 1347 7053 1362
tri 7053 1347 7068 1362 nw
tri 6918 1287 6978 1347 se
rect 6978 1287 6993 1347
tri 6993 1287 7053 1347 nw
tri 6843 1212 6918 1287 se
tri 6918 1212 6993 1287 nw
tri 6820 1189 6843 1212 se
rect 6843 1189 6895 1212
tri 6895 1189 6918 1212 nw
rect 6275 870 6281 986
rect 6461 870 6467 986
tri 5616 -197 5644 -169 se
rect 5644 -197 6205 -169
tri 5564 -249 5616 -197 se
rect 5616 -249 6205 -197
rect 3749 -367 3755 -315
rect 3807 -367 3819 -315
rect 3871 -367 3877 -315
tri 4347 -367 4399 -315 se
rect 4399 -367 4612 -315
rect 3749 -1324 3877 -367
tri 4296 -418 4347 -367 se
rect 4347 -418 4612 -367
rect 4296 -1228 4612 -418
tri 5395 -418 5564 -249 se
rect 5564 -418 6205 -249
rect 5395 -1238 6205 -418
tri 5395 -1296 5453 -1238 ne
rect 3593 -1424 3877 -1324
tri 3877 -1424 3977 -1324 sw
rect 5453 -1330 6205 -1238
rect 5453 -1424 6111 -1330
tri 6111 -1424 6205 -1330 nw
rect 6261 -1424 6483 57
tri 6795 17 6820 42 se
rect 6820 17 6872 1189
tri 6872 1166 6895 1189 nw
rect 6742 -35 6748 17
rect 6800 -35 6814 17
rect 6866 -35 6872 17
tri 7158 -197 7183 -172 se
rect 7183 -197 7235 2161
rect 7329 1445 7335 1497
rect 7387 1445 7399 1497
rect 7451 1445 7457 1497
rect 7329 807 7381 1445
tri 7381 1369 7457 1445 nw
tri 8318 1369 8352 1403 se
rect 8352 1369 8890 2161
rect 9055 1598 9061 1650
rect 9113 1598 9125 1650
rect 9177 1644 10038 1650
rect 9177 1598 9986 1644
tri 9959 1592 9965 1598 ne
rect 9965 1592 9986 1598
tri 9965 1580 9977 1592 ne
rect 9977 1580 10038 1592
tri 9977 1571 9986 1580 ne
rect 9986 1522 10038 1528
rect 7329 743 7381 755
rect 7329 685 7381 691
tri 8302 1353 8318 1369 se
rect 8318 1353 8890 1369
rect 8302 1347 8890 1353
rect 8418 1103 8890 1347
rect 8302 1090 8890 1103
rect 8354 1038 8366 1090
rect 8418 1038 8890 1090
rect 8302 1025 8890 1038
rect 8354 973 8366 1025
rect 8418 973 8890 1025
rect 8302 960 8890 973
rect 8354 908 8366 960
rect 8418 908 8890 960
rect 8302 895 8890 908
rect 8354 843 8366 895
rect 8418 843 8890 895
rect 8302 830 8890 843
rect 8354 778 8366 830
rect 8418 778 8890 830
rect 8302 765 8890 778
rect 8354 713 8366 765
rect 8418 713 8890 765
rect 8302 700 8890 713
rect 8354 648 8366 700
rect 8418 648 8890 700
rect 8302 635 8890 648
rect 8354 583 8366 635
rect 8418 583 8890 635
rect 8302 570 8890 583
rect 8354 518 8366 570
rect 8418 518 8890 570
rect 8302 505 8890 518
rect 8354 453 8366 505
rect 8418 453 8890 505
rect 8302 440 8890 453
rect 8354 388 8366 440
rect 8418 388 8890 440
rect 8302 375 8890 388
rect 8354 323 8366 375
rect 8418 323 8890 375
rect 8302 310 8890 323
rect 8354 258 8366 310
rect 8418 258 8890 310
rect 8302 245 8890 258
rect 8354 193 8366 245
rect 8418 193 8890 245
rect 8302 180 8890 193
rect 8354 128 8366 180
rect 8418 128 8890 180
rect 8302 115 8890 128
rect 8354 63 8366 115
rect 8418 63 8890 115
rect 8302 57 8890 63
tri 8302 -180 8539 57 ne
rect 7105 -249 7111 -197
rect 7163 -249 7177 -197
rect 7229 -249 7235 -197
tri 6483 -1424 6502 -1405 sw
tri 2582 -1738 2643 -1677 se
rect 2643 -1738 2776 -1677
tri 2776 -1738 2837 -1677 nw
rect 2582 -1776 2738 -1738
tri 2738 -1776 2776 -1738 nw
rect 3593 -1776 3977 -1424
tri 3977 -1776 4329 -1424 sw
tri 1710 -2984 1760 -2934 sw
rect 1518 -3012 1760 -2984
tri 1518 -3072 1578 -3012 ne
rect 1578 -3614 1760 -3012
rect 1816 -3614 2523 -1776
rect 2582 -3438 2720 -1776
tri 2720 -1794 2738 -1776 nw
rect 2581 -3614 2720 -3438
rect 3009 -3614 3422 -1776
rect 3593 -2582 4329 -1776
tri 3593 -2869 3880 -2582 ne
rect 3880 -3614 4329 -2582
rect 5453 -1457 6078 -1424
tri 6078 -1457 6111 -1424 nw
rect 5453 -1495 6040 -1457
tri 6040 -1495 6078 -1457 nw
tri 6223 -1495 6261 -1457 se
rect 6261 -1495 6502 -1424
rect 5453 -3632 5927 -1495
tri 5927 -1608 6040 -1495 nw
tri 6110 -1608 6223 -1495 se
rect 6223 -1608 6502 -1495
tri 6502 -1608 6686 -1424 sw
tri 6040 -1678 6110 -1608 se
rect 6110 -1678 6686 -1608
rect 6040 -1776 6686 -1678
tri 6686 -1776 6854 -1608 sw
rect 6040 -2586 6854 -1776
rect 6040 -3632 6360 -2586
tri 6360 -3080 6854 -2586 nw
rect 8062 -2586 8378 -1761
rect 8062 -3632 8261 -2586
tri 8261 -2703 8378 -2586 nw
rect 8539 -3632 8890 57
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 1 0 3563 0 1 1457
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 1 0 7931 0 1 1219
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 1 0 6275 0 1 870
box 0 0 1 1
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_0
timestamp 1707688321
transform 1 0 -2505 0 1 -2580
box -5 0 301 794
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_1
timestamp 1707688321
transform 1 0 -2985 0 1 -2580
box -5 0 301 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_0
timestamp 1707688321
transform 1 0 -1592 0 1 -2580
box -5 0 141 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_1
timestamp 1707688321
transform 1 0 -158 0 1 -2580
box -5 0 141 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_2
timestamp 1707688321
transform 1 0 1023 0 1 -2580
box -5 0 141 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_3
timestamp 1707688321
transform 1 0 1542 0 1 -2580
box -5 0 141 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_4
timestamp 1707688321
transform 1 0 2582 0 1 -2580
box -5 0 141 794
use M2M3_CDNS_524688791851606  M2M3_CDNS_524688791851606_0
timestamp 1707688321
transform 1 0 3629 0 1 -2580
box -5 0 221 794
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_0
timestamp 1707688321
transform 1 0 3020 0 1 565
box -79 -26 535 1026
use nfet_CDNS_524688791851608  nfet_CDNS_524688791851608_1
timestamp 1707688321
transform 1 0 2508 0 1 565
box -79 -26 535 1026
use nfet_CDNS_524688791851609  nfet_CDNS_524688791851609_0
timestamp 1707688321
transform -1 0 2452 0 1 565
box -79 -26 179 1026
use nfet_CDNS_524688791851609  nfet_CDNS_524688791851609_1
timestamp 1707688321
transform 1 0 3532 0 1 565
box -79 -26 179 1026
use pfet_CDNS_524688791851610  pfet_CDNS_524688791851610_0
timestamp 1707688321
transform -1 0 8180 0 -1 1171
box -89 -36 245 1036
use PYbentRes_CDNS_524688791851611  PYbentRes_CDNS_524688791851611_0
timestamp 1707688321
transform 0 -1 9137 1 0 -3340
box -50 -162 25348 66
use PYbentRes_CDNS_524688791851612  PYbentRes_CDNS_524688791851612_0
timestamp 1707688321
transform 0 -1 10497 1 0 -1630
box -50 -162 23637 66
use PYbentRes_CDNS_524688791851613  PYbentRes_CDNS_524688791851613_0
timestamp 1707688321
transform 0 -1 10335 1 0 12543
box -50 0 9462 66
use PYbentRes_CDNS_524688791851614  PYbentRes_CDNS_524688791851614_0
timestamp 1707688321
transform 0 -1 10011 -1 0 21957
box -50 -162 24463 66
use PYbentRes_CDNS_524688791851615  PYbentRes_CDNS_524688791851615_0
timestamp 1707688321
transform 0 -1 9687 -1 0 21957
box -50 -162 28185 66
use PYbentRes_CDNS_524688791851616  PYbentRes_CDNS_524688791851616_0
timestamp 1707688321
transform 0 -1 9525 1 0 -6000
box -50 0 28008 66
use sky130_fd_io__sio_tk_em1c_CDNS_524688791851607  sky130_fd_io__sio_tk_em1c_CDNS_524688791851607_0
timestamp 1707688321
transform 0 1 10272 1 0 21718
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1707688321
transform -1 0 9286 0 1 -3128
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1707688321
transform -1 0 10665 0 1 -1674
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_2
timestamp 1707688321
transform -1 0 10125 0 1 21898
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_3
timestamp 1707688321
transform -1 0 9459 0 1 -3128
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_4
timestamp 1707688321
transform -1 0 9811 0 1 21898
box 0 0 1 1
<< labels >>
flabel comment s 5121 -3597 5121 -3597 3 FreeSans 200 90 0 0 vnb
flabel comment s 4404 -3597 4404 -3597 3 FreeSans 200 90 0 0 vnb
flabel comment s 3235 -3604 3235 -3604 3 FreeSans 200 90 0 0 vnb
flabel comment s 2152 -3616 2152 -3616 3 FreeSans 200 90 0 0 vnb
flabel comment s 654 -3579 654 -3579 3 FreeSans 200 90 0 0 vnb
flabel comment s -530 -3560 -530 -3560 3 FreeSans 200 90 0 0 vnb
flabel comment s -5761 -36 -5761 -36 3 FreeSans 200 270 0 0 pad
flabel comment s -5997 -1299 -5997 -1299 3 FreeSans 200 0 0 0 oe_hs_h
flabel comment s 328 -3535 328 -3535 3 FreeSans 200 90 0 0 od_h
flabel comment s 328 -374 328 -374 3 FreeSans 200 270 0 0 od_h
flabel comment s 418 -374 418 -374 3 FreeSans 200 270 0 0 oe_hs_h
flabel comment s 2284 -229 2284 -229 3 FreeSans 200 0 0 0 drvhi_h
flabel comment s 2284 -156 2284 -156 3 FreeSans 200 0 0 0 puen_reg_h
flabel comment s 2284 -16 2284 -16 3 FreeSans 200 0 0 0 vreg_en_h
flabel comment s 2284 75 2284 75 3 FreeSans 200 0 0 0 slow_h_n
flabel comment s 1610 -3536 1610 -3536 3 FreeSans 200 90 0 0 vgnd
flabel comment s 1090 -3536 1090 -3536 3 FreeSans 200 90 0 0 vgnd
flabel comment s -89 -3536 -89 -3536 3 FreeSans 200 90 0 0 vgnd
flabel comment s -819 -1150 -819 -1150 3 FreeSans 200 90 0 0 vcc_io
flabel comment s -1519 -3536 -1519 -3536 3 FreeSans 200 90 0 0 vgnd
flabel comment s -5761 -3536 -5761 -3536 3 FreeSans 200 90 0 0 pad
flabel comment s -3972 -378 -3972 -378 3 FreeSans 200 270 0 0 vgnd
flabel comment s -1519 -378 -1519 -378 3 FreeSans 200 270 0 0 vgnd
flabel comment s -819 -378 -819 -378 3 FreeSans 200 270 0 0 vcc_io
flabel comment s -89 -378 -89 -378 3 FreeSans 200 270 0 0 vgnd
flabel comment s 1090 -378 1090 -378 3 FreeSans 200 270 0 0 vgnd
flabel comment s 1610 -378 1610 -378 3 FreeSans 200 270 0 0 vgnd
flabel comment s 2775 -3522 2775 -3522 3 FreeSans 200 90 0 0 vgnd
flabel comment s 2409 -416 2409 -416 3 FreeSans 200 90 0 0 vcc_io
flabel comment s 3506 2051 3506 2051 3 FreeSans 200 270 0 0 slow_h_n
flabel comment s 2775 2051 2775 2051 3 FreeSans 200 270 0 0 vgnd
flabel comment s 2409 2051 2409 2051 3 FreeSans 200 270 0 0 vcc_io
flabel comment s 6082 -3509 6082 -3509 3 FreeSans 200 90 0 0 vcc_io
flabel comment s 8445 -3588 8445 -3588 3 FreeSans 200 90 0 0 vpwr_ka
flabel comment s 8445 2051 8445 2051 3 FreeSans 200 270 0 0 vpwr_ka
flabel comment s 7085 2051 7085 2051 3 FreeSans 200 270 0 0 vreg_en_h
flabel comment s 6424 2051 6424 2051 3 FreeSans 200 270 0 0 vnb
flabel comment s 6082 2051 6082 2051 3 FreeSans 200 270 0 0 vcc_io
flabel comment s 5115 2051 5115 2051 3 FreeSans 200 270 0 0 puen_reg_h
flabel comment s 4520 2051 4520 2051 3 FreeSans 200 270 0 0 vcc_io
flabel comment s 7208 2128 7208 2128 3 FreeSans 200 270 0 0 drvhi_h
flabel metal1 s 2269 1505 2323 1557 0 FreeSans 600 0 0 0 ngate
port 2 nsew
flabel metal2 s 3593 2076 3721 2104 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 7329 1369 7381 1414 0 FreeSans 200 0 0 0 vreg_en_n
port 4 nsew
<< properties >>
string GDS_END 98190060
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98012502
string path 55.350 4.775 101.475 4.775 101.475 46.800 
<< end >>
