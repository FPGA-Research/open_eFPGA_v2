magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 129 226
<< nmos >>
rect 0 0 50 200
<< ndiff >>
rect -50 0 0 200
rect 50 182 103 200
rect 50 148 61 182
rect 95 148 103 182
rect 50 114 103 148
rect 50 80 61 114
rect 95 80 103 114
rect 50 46 103 80
rect 50 12 61 46
rect 95 12 103 46
rect 50 0 103 12
<< ndiffc >>
rect 61 148 95 182
rect 61 80 95 114
rect 61 12 95 46
<< poly >>
rect 0 200 50 226
rect 0 -26 50 0
<< locali >>
rect 61 182 95 198
rect 61 114 95 148
rect 61 46 95 80
rect 61 -4 95 12
<< metal1 >>
rect -51 -16 -5 186
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_0
timestamp 1707688321
transform 1 0 50 0 1 0
box 0 0 1 1
use DFM1sd_CDNS_52468879185186  DFM1sd_CDNS_52468879185186_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 78 97 78 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85976448
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85975626
<< end >>
