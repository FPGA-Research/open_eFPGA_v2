magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 151 47 181 177
rect 254 47 284 177
rect 349 47 379 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 254 297 284 497
rect 349 297 379 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 47 151 177
rect 181 47 254 177
rect 284 161 349 177
rect 284 127 294 161
rect 328 127 349 161
rect 284 93 349 127
rect 284 59 294 93
rect 328 59 349 93
rect 284 47 349 59
rect 379 97 433 177
rect 379 63 391 97
rect 425 63 433 97
rect 379 47 433 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 467 163 497
rect 109 433 119 467
rect 153 433 163 467
rect 109 297 163 433
rect 193 485 254 497
rect 193 451 203 485
rect 237 451 254 485
rect 193 297 254 451
rect 284 467 349 497
rect 284 433 294 467
rect 328 433 349 467
rect 284 297 349 433
rect 379 485 433 497
rect 379 451 391 485
rect 425 451 433 485
rect 379 417 433 451
rect 379 383 391 417
rect 425 383 433 417
rect 379 349 433 383
rect 379 315 391 349
rect 425 315 433 349
rect 379 297 433 315
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 294 127 328 161
rect 294 59 328 93
rect 391 63 425 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 433 153 467
rect 203 451 237 485
rect 294 433 328 467
rect 391 451 425 485
rect 391 383 425 417
rect 391 315 425 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 254 497 284 523
rect 349 497 379 523
rect 79 265 109 297
rect 163 265 193 297
rect 254 265 284 297
rect 349 265 379 297
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 79 177 109 199
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 301 265
rect 247 215 257 249
rect 291 215 301 249
rect 247 199 301 215
rect 349 249 439 265
rect 349 215 395 249
rect 429 215 439 249
rect 349 199 439 215
rect 151 177 181 199
rect 254 177 284 199
rect 349 177 379 199
rect 79 21 109 47
rect 151 21 181 47
rect 254 21 284 47
rect 349 21 379 47
<< polycont >>
rect 31 215 65 249
rect 161 215 195 249
rect 257 215 291 249
rect 395 215 429 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 18 485 84 527
rect 18 451 35 485
rect 69 451 84 485
rect 187 485 253 527
rect 18 417 84 451
rect 18 383 35 417
rect 69 383 84 417
rect 18 349 84 383
rect 118 467 153 483
rect 118 433 119 467
rect 187 451 203 485
rect 237 451 253 485
rect 375 485 442 489
rect 187 435 253 451
rect 294 467 339 483
rect 118 401 153 433
rect 328 433 339 467
rect 294 401 339 433
rect 118 367 339 401
rect 375 451 391 485
rect 425 451 442 485
rect 375 417 442 451
rect 375 383 391 417
rect 425 383 442 417
rect 18 315 35 349
rect 69 315 84 349
rect 375 349 442 383
rect 375 333 391 349
rect 18 299 84 315
rect 214 289 291 333
rect 17 249 73 265
rect 17 215 31 249
rect 65 215 73 249
rect 17 199 73 215
rect 122 249 211 255
rect 122 215 161 249
rect 195 215 211 249
rect 18 129 35 163
rect 69 129 86 163
rect 18 95 86 129
rect 18 61 35 95
rect 69 61 86 95
rect 122 67 211 215
rect 254 249 291 289
rect 254 215 257 249
rect 254 199 291 215
rect 325 315 391 333
rect 425 315 442 349
rect 325 299 442 315
rect 325 165 359 299
rect 393 249 443 265
rect 393 215 395 249
rect 429 215 443 249
rect 393 199 443 215
rect 276 161 359 165
rect 276 127 294 161
rect 328 143 359 161
rect 328 127 357 143
rect 276 93 357 127
rect 18 17 86 61
rect 276 59 294 93
rect 328 59 357 93
rect 391 97 443 113
rect 425 63 443 97
rect 391 17 443 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 396 425 430 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 396 357 430 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 85 156 119 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a31oi_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 4127366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4122120
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
