magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -66 377 4098 897
<< pwell >>
rect 1330 226 1890 230
rect 1064 217 1890 226
rect 2215 217 4028 283
rect 9 43 4028 217
rect -26 -43 4058 43
<< locali >>
rect 121 333 359 433
rect 395 369 461 471
rect 536 333 591 353
rect 121 299 591 333
rect 536 219 591 299
rect 697 162 738 430
rect 876 236 942 430
rect 2041 242 2471 276
rect 2437 87 2471 242
rect 2800 285 2969 329
rect 2800 87 2834 285
rect 2437 53 2834 87
rect 3481 99 3557 747
rect 3940 471 4007 687
rect 3961 265 4007 471
rect 3940 99 4007 265
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 128 735 318 741
rect 128 701 134 735
rect 168 701 206 735
rect 240 701 278 735
rect 312 701 318 735
rect 26 541 92 661
rect 128 577 318 701
rect 683 735 861 741
rect 717 701 755 735
rect 789 701 827 735
rect 480 611 546 661
rect 480 577 647 611
rect 26 507 577 541
rect 26 263 60 507
rect 527 403 577 507
rect 613 525 647 577
rect 683 561 861 701
rect 897 727 1103 761
rect 897 525 931 727
rect 967 561 1033 691
rect 613 491 931 525
rect 26 219 460 263
rect 26 99 97 219
rect 627 183 661 491
rect 133 113 323 183
rect 133 79 139 113
rect 173 79 211 113
rect 245 79 283 113
rect 317 79 323 113
rect 485 149 661 183
rect 988 374 1033 561
rect 1069 444 1103 727
rect 1139 735 1173 741
rect 1723 735 1913 741
rect 1139 480 1173 701
rect 1209 678 1459 712
rect 1209 444 1243 678
rect 1069 410 1243 444
rect 1279 458 1329 642
rect 1368 548 1459 678
rect 1723 701 1729 735
rect 1763 701 1801 735
rect 1835 701 1873 735
rect 1907 701 1913 735
rect 988 340 1213 374
rect 485 99 551 149
rect 774 113 952 199
rect 133 73 323 79
rect 808 79 846 113
rect 880 79 918 113
rect 988 103 1038 340
rect 1147 240 1213 340
rect 1279 204 1313 458
rect 1368 212 1402 548
rect 1074 113 1192 204
rect 774 73 952 79
rect 1074 79 1080 113
rect 1114 79 1152 113
rect 1186 79 1192 113
rect 1074 73 1192 79
rect 1238 87 1313 204
rect 1352 123 1402 212
rect 1438 458 1504 512
rect 1438 87 1472 458
rect 1540 416 1599 648
rect 1723 592 1913 701
rect 2191 735 2381 751
rect 2191 701 2197 735
rect 2231 701 2269 735
rect 2303 701 2341 735
rect 2375 701 2381 735
rect 2191 670 2381 701
rect 1949 634 2155 668
rect 1949 556 1983 634
rect 2121 600 2467 634
rect 1640 522 1983 556
rect 1640 458 1706 522
rect 2019 486 2085 598
rect 1782 452 2085 486
rect 2263 416 2329 511
rect 2405 459 2467 600
rect 2503 539 2569 751
rect 2700 735 2890 741
rect 2700 701 2706 735
rect 2740 701 2778 735
rect 2812 701 2850 735
rect 2884 701 2890 735
rect 2700 575 2890 701
rect 3248 735 3438 747
rect 3248 701 3254 735
rect 3288 701 3326 735
rect 3360 701 3398 735
rect 3432 701 3438 735
rect 2994 539 3060 635
rect 2503 505 3060 539
rect 2405 425 2681 459
rect 1540 382 2329 416
rect 1540 212 1574 382
rect 2440 346 2506 375
rect 1508 128 1574 212
rect 1610 312 2506 346
rect 1610 230 1665 312
rect 2633 283 2681 425
rect 2717 399 2751 505
rect 3137 469 3212 535
rect 2787 435 3212 469
rect 3248 439 3438 701
rect 2717 365 3109 399
rect 1610 87 1644 230
rect 1782 228 1982 276
rect 1238 53 1644 87
rect 1682 113 1872 192
rect 1682 79 1688 113
rect 1722 79 1760 113
rect 1794 79 1832 113
rect 1866 79 1872 113
rect 1916 103 1982 228
rect 2109 113 2299 206
rect 1682 73 1872 79
rect 2109 79 2115 113
rect 2149 79 2187 113
rect 2221 79 2259 113
rect 2293 79 2299 113
rect 2109 73 2299 79
rect 2531 157 2597 265
rect 2717 157 2751 365
rect 2531 123 2751 157
rect 3043 285 3109 365
rect 2870 113 3060 249
rect 3146 165 3212 435
rect 2870 79 2876 113
rect 2910 79 2948 113
rect 2982 79 3020 113
rect 3054 79 3060 113
rect 2870 73 3060 79
rect 3248 113 3438 265
rect 3248 79 3254 113
rect 3288 79 3326 113
rect 3360 79 3398 113
rect 3432 79 3438 113
rect 3707 735 3897 741
rect 3707 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 3897 735
rect 3605 335 3671 637
rect 3707 471 3897 701
rect 3849 335 3915 435
rect 3605 301 3915 335
rect 3605 165 3671 301
rect 3707 113 3897 265
rect 3248 73 3438 79
rect 3707 79 3713 113
rect 3747 79 3785 113
rect 3819 79 3857 113
rect 3891 79 3897 113
rect 3707 73 3897 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 3391 797 3425 831
rect 3487 797 3521 831
rect 3583 797 3617 831
rect 3679 797 3713 831
rect 3775 797 3809 831
rect 3871 797 3905 831
rect 3967 797 4001 831
rect 134 701 168 735
rect 206 701 240 735
rect 278 701 312 735
rect 683 701 717 735
rect 755 701 789 735
rect 827 701 861 735
rect 139 79 173 113
rect 211 79 245 113
rect 283 79 317 113
rect 1139 701 1173 735
rect 1729 701 1763 735
rect 1801 701 1835 735
rect 1873 701 1907 735
rect 774 79 808 113
rect 846 79 880 113
rect 918 79 952 113
rect 1080 79 1114 113
rect 1152 79 1186 113
rect 2197 701 2231 735
rect 2269 701 2303 735
rect 2341 701 2375 735
rect 2706 701 2740 735
rect 2778 701 2812 735
rect 2850 701 2884 735
rect 3254 701 3288 735
rect 3326 701 3360 735
rect 3398 701 3432 735
rect 1688 79 1722 113
rect 1760 79 1794 113
rect 1832 79 1866 113
rect 2115 79 2149 113
rect 2187 79 2221 113
rect 2259 79 2293 113
rect 2876 79 2910 113
rect 2948 79 2982 113
rect 3020 79 3054 113
rect 3254 79 3288 113
rect 3326 79 3360 113
rect 3398 79 3432 113
rect 3713 701 3747 735
rect 3785 701 3819 735
rect 3857 701 3891 735
rect 3713 79 3747 113
rect 3785 79 3819 113
rect 3857 79 3891 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
<< metal1 >>
rect 0 831 4032 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3391 831
rect 3425 797 3487 831
rect 3521 797 3583 831
rect 3617 797 3679 831
rect 3713 797 3775 831
rect 3809 797 3871 831
rect 3905 797 3967 831
rect 4001 797 4032 831
rect 0 791 4032 797
rect 0 735 4032 763
rect 0 701 134 735
rect 168 701 206 735
rect 240 701 278 735
rect 312 701 683 735
rect 717 701 755 735
rect 789 701 827 735
rect 861 701 1139 735
rect 1173 701 1729 735
rect 1763 701 1801 735
rect 1835 701 1873 735
rect 1907 701 2197 735
rect 2231 701 2269 735
rect 2303 701 2341 735
rect 2375 701 2706 735
rect 2740 701 2778 735
rect 2812 701 2850 735
rect 2884 701 3254 735
rect 3288 701 3326 735
rect 3360 701 3398 735
rect 3432 701 3713 735
rect 3747 701 3785 735
rect 3819 701 3857 735
rect 3891 701 4032 735
rect 0 689 4032 701
rect 0 113 4032 125
rect 0 79 139 113
rect 173 79 211 113
rect 245 79 283 113
rect 317 79 774 113
rect 808 79 846 113
rect 880 79 918 113
rect 952 79 1080 113
rect 1114 79 1152 113
rect 1186 79 1688 113
rect 1722 79 1760 113
rect 1794 79 1832 113
rect 1866 79 2115 113
rect 2149 79 2187 113
rect 2221 79 2259 113
rect 2293 79 2876 113
rect 2910 79 2948 113
rect 2982 79 3020 113
rect 3054 79 3254 113
rect 3288 79 3326 113
rect 3360 79 3398 113
rect 3432 79 3713 113
rect 3747 79 3785 113
rect 3819 79 3857 113
rect 3891 79 4032 113
rect 0 51 4032 79
rect 0 17 4032 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4032 17
rect 0 -23 4032 -17
<< labels >>
rlabel locali s 876 236 942 430 6 CLK
port 1 nsew clock input
rlabel locali s 395 369 461 471 6 D
port 2 nsew signal input
rlabel locali s 697 162 738 430 6 SCD
port 3 nsew signal input
rlabel locali s 536 219 591 299 6 SCE
port 4 nsew signal input
rlabel locali s 121 299 591 333 6 SCE
port 4 nsew signal input
rlabel locali s 536 333 591 353 6 SCE
port 4 nsew signal input
rlabel locali s 121 333 359 433 6 SCE
port 4 nsew signal input
rlabel locali s 2437 53 2834 87 6 SET_B
port 5 nsew signal input
rlabel locali s 2800 87 2834 285 6 SET_B
port 5 nsew signal input
rlabel locali s 2437 87 2471 242 6 SET_B
port 5 nsew signal input
rlabel locali s 2041 242 2471 276 6 SET_B
port 5 nsew signal input
rlabel locali s 2800 285 2969 329 6 SET_B
port 5 nsew signal input
rlabel metal1 s 0 51 4032 125 6 VGND
port 6 nsew ground bidirectional
rlabel metal1 s 0 -23 4032 23 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s -26 -43 4058 43 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 9 43 4028 217 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2215 217 4028 283 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1064 217 1890 226 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1330 226 1890 230 6 VNB
port 7 nsew ground bidirectional
rlabel metal1 s 0 791 4032 837 6 VPB
port 8 nsew power bidirectional
rlabel nwell s -66 377 4098 897 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 689 4032 763 6 VPWR
port 9 nsew power bidirectional
rlabel locali s 3940 99 4007 265 6 Q
port 10 nsew signal output
rlabel locali s 3961 265 4007 471 6 Q
port 10 nsew signal output
rlabel locali s 3940 471 4007 687 6 Q
port 10 nsew signal output
rlabel locali s 3481 99 3557 747 6 Q_N
port 11 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 4032 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 570340
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 531624
<< end >>
