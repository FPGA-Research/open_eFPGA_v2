magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1563 203
rect 30 -17 64 21
<< locali >>
rect 1215 383 1449 417
rect 24 199 347 265
rect 387 199 710 265
rect 765 199 1084 265
rect 1134 199 1371 326
rect 1409 161 1449 383
rect 795 127 1517 161
rect 1315 51 1349 127
rect 1483 51 1517 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 35 333 69 493
rect 103 383 169 527
rect 203 333 237 493
rect 271 383 337 527
rect 371 333 405 493
rect 439 383 505 527
rect 539 333 573 493
rect 607 383 673 527
rect 707 333 741 493
rect 779 383 845 527
rect 879 333 913 493
rect 947 451 1013 527
rect 1047 485 1081 493
rect 1047 451 1533 485
rect 1047 333 1081 451
rect 35 299 1081 333
rect 1483 299 1533 451
rect 35 127 757 161
rect 35 51 69 127
rect 103 17 169 93
rect 203 51 237 127
rect 271 17 337 93
rect 371 51 405 127
rect 439 59 1113 93
rect 1215 17 1281 93
rect 1383 17 1449 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 765 199 1084 265 6 A1
port 1 nsew signal input
rlabel locali s 387 199 710 265 6 A2
port 2 nsew signal input
rlabel locali s 24 199 347 265 6 A3
port 3 nsew signal input
rlabel locali s 1134 199 1371 326 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1563 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1483 51 1517 127 6 Y
port 9 nsew signal output
rlabel locali s 1315 51 1349 127 6 Y
port 9 nsew signal output
rlabel locali s 795 127 1517 161 6 Y
port 9 nsew signal output
rlabel locali s 1409 161 1449 383 6 Y
port 9 nsew signal output
rlabel locali s 1215 383 1449 417 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4149346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4136480
<< end >>
