magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 876 1026
<< nmos >>
rect 0 0 800 1000
<< ndiff >>
rect -50 0 0 1000
rect 800 0 850 1000
<< poly >>
rect 0 1000 800 1032
rect 0 -32 800 0
<< locali >>
rect -45 -4 -11 946
rect 811 -4 845 946
use hvDFL1sd_CDNS_5595914180851  hvDFL1sd_CDNS_5595914180851_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 1026
use hvDFL1sd_CDNS_5595914180851  hvDFL1sd_CDNS_5595914180851_1
timestamp 1707688321
transform 1 0 800 0 1 0
box -26 -26 79 1026
<< labels >>
flabel comment s 828 471 828 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 43011900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43011074
<< end >>
