magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect 3644 -1467 3778 -1451
rect 3644 -1501 3660 -1467
rect 3694 -1501 3728 -1467
rect 3762 -1501 3778 -1467
rect 3644 -1517 3778 -1501
<< polycont >>
rect 3660 -1501 3694 -1467
rect 3728 -1501 3762 -1467
<< locali >>
rect 2919 7276 3388 7282
rect 2919 7242 2931 7276
rect 2965 7242 3021 7276
rect 3055 7272 3388 7276
rect 3055 7242 3193 7272
rect 2919 7238 3193 7242
rect 3227 7238 3268 7272
rect 3302 7238 3342 7272
rect 3376 7238 3388 7272
rect 2919 7180 3388 7238
rect 2919 7146 2931 7180
rect 2965 7146 3021 7180
rect 3055 7176 3388 7180
rect 3055 7146 3193 7176
rect 2919 7142 3193 7146
rect 3227 7142 3268 7176
rect 3302 7142 3342 7176
rect 3376 7142 3388 7176
rect 2919 7133 3388 7142
rect 3644 -1501 3654 -1467
rect 3694 -1501 3726 -1467
rect 3762 -1501 3778 -1467
<< viali >>
rect 2931 7242 2965 7276
rect 3021 7242 3055 7276
rect 3193 7238 3227 7272
rect 3268 7238 3302 7272
rect 3342 7238 3376 7272
rect 2931 7146 2965 7180
rect 3021 7146 3055 7180
rect 3193 7142 3227 7176
rect 3268 7142 3302 7176
rect 3342 7142 3376 7176
rect 3654 -1501 3660 -1467
rect 3660 -1501 3688 -1467
rect 3726 -1501 3728 -1467
rect 3728 -1501 3760 -1467
<< metal1 >>
tri 4502 8653 4531 8682 ne
tri 4500 7282 4531 7313 se
rect 4531 7282 4577 8682
tri 4577 8653 4606 8682 nw
tri 2902 7276 2908 7282 se
rect 2908 7276 3067 7282
tri 4496 7278 4500 7282 se
rect 4500 7278 4577 7282
tri 2868 7242 2902 7276 se
rect 2902 7242 2931 7276
rect 2965 7242 3021 7276
rect 3055 7242 3067 7276
tri 2864 7238 2868 7242 se
rect 2868 7238 3067 7242
tri 2817 7191 2864 7238 se
rect 2864 7191 3067 7238
rect 2817 7180 3067 7191
rect 2817 7146 2931 7180
rect 2965 7146 3021 7180
rect 3055 7146 3067 7180
rect 2817 7140 3067 7146
rect 3181 7272 4577 7278
rect 3181 7238 3193 7272
rect 3227 7238 3268 7272
rect 3302 7238 3342 7272
rect 3376 7238 4577 7272
rect 3181 7226 4577 7238
rect 3181 7176 4487 7226
rect 3181 7142 3193 7176
rect 3227 7142 3268 7176
rect 3302 7142 3342 7176
rect 3376 7142 4487 7176
rect 2817 7136 2897 7140
tri 2897 7136 2901 7140 nw
rect 3181 7136 4487 7142
tri 4487 7136 4577 7226 nw
rect 2817 -997 2863 7136
tri 2863 7102 2897 7136 nw
tri 2817 -1039 2859 -997 ne
rect 2859 -1039 2863 -997
tri 2863 -1039 2925 -977 sw
tri 2859 -1043 2863 -1039 ne
rect 2863 -1043 3617 -1039
tri 2863 -1085 2905 -1043 ne
rect 2905 -1085 3617 -1043
tri 3597 -1095 3607 -1085 ne
rect 3607 -1095 3617 -1085
tri 3617 -1095 3673 -1039 sw
tri 3607 -1105 3617 -1095 ne
rect 3617 -1105 3673 -1095
tri 3617 -1115 3627 -1105 ne
rect 3627 -1239 3673 -1105
rect 3783 -1209 3835 -1203
rect 3783 -1281 3835 -1261
rect 3783 -1353 3835 -1333
rect 3783 -1411 3835 -1405
tri 3571 -1461 3598 -1434 sw
rect 3571 -1467 3772 -1461
rect 3571 -1501 3654 -1467
rect 3688 -1501 3726 -1467
rect 3760 -1501 3772 -1467
rect 3571 -1507 3772 -1501
tri 3571 -1534 3598 -1507 nw
<< via1 >>
rect 3783 -1261 3835 -1209
rect 3783 -1333 3835 -1281
rect 3783 -1405 3835 -1353
<< metal2 >>
rect 3783 -1209 3835 -1203
rect 3783 -1281 3835 -1261
rect 3783 -1353 3835 -1333
rect 3783 -1411 3835 -1405
use nfet_CDNS_524688791851003  nfet_CDNS_524688791851003_0
timestamp 1707688321
transform 1 0 3678 0 -1 -1219
box -79 -32 179 232
use sky130_fd_io__opamp_biasgen_1  sky130_fd_io__opamp_biasgen_1_0
timestamp 1707688321
transform 1 0 2747 0 1 -1600
box -570 0 4434 12782
use sky130_fd_io__opamp_stage  sky130_fd_io__opamp_stage_0
timestamp 1707688321
transform 1 0 0 0 1 0
box -59 -46 2937 8816
<< properties >>
string GDS_END 80489548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80487222
string path 95.225 -35.275 95.225 -30.075 
<< end >>
