magic
tech sky130B
magscale 1 2
timestamp 1707688321
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_0
timestamp 1707688321
transform -1 0 14983 0 1 494
box 0 0 1 1
use sky130_fd_io__gpiov2_amux_ctl_inv_1  sky130_fd_io__gpiov2_amux_ctl_inv_1_1
timestamp 1707688321
transform -1 0 15292 0 1 494
box 0 0 1 1
use sky130_fd_io__gpiov2_amux_ctl_ls  sky130_fd_io__gpiov2_amux_ctl_ls_0
timestamp 1707688321
transform 1 0 14705 0 1 1344
box 174 163 2111 1297
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv2  sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0
timestamp 1707688321
transform 1 0 748 0 1 13628
box 290 665 1777 3319
use sky130_fd_io__gpiov2_amux_ctl_lshv2hv  sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0
timestamp 1707688321
transform -1 0 8787 0 1 10523
box 3564 882 6767 1251
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1707688321
transform -1 0 14675 0 1 494
box -38 -49 134 715
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808586  sky130_fd_pr__model__nfet_highvoltage__example_55959141808586_0
timestamp 1707688321
transform -1 0 1459 0 -1 11410
box -1 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808421  sky130_fd_pr__model__pfet_highvoltage__example_55959141808421_0
timestamp 1707688321
transform 1 0 1286 0 -1 10835
box -1 0 297 1
<< properties >>
string GDS_END 22069112
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22043456
<< end >>
