magic
tech sky130A
timestamp 1707688321
<< properties >>
string GDS_END 94744154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94743386
<< end >>
