magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -266 -66 239 666
<< mvpmos >>
rect 0 0 120 600
<< mvpdiff >>
rect -50 0 0 600
rect 120 0 170 600
<< poly >>
rect 0 600 120 632
rect 0 -32 120 0
<< locali >>
rect -113 -4 -11 550
rect 131 -4 165 538
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_0
timestamp 1707688321
transform 1 0 120 0 1 0
box -36 -36 89 636
use hvDFTPL1s_CDNS_52468879185914  hvDFTPL1s_CDNS_52468879185914_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 236 636
<< labels >>
flabel comment s -62 273 -62 273 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80652720
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80651702
<< end >>
