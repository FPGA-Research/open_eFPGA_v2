magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 458 2540 899
<< pwell >>
rect 43 0 2421 86
<< mvpsubdiff >>
rect 69 26 93 60
rect 127 26 161 60
rect 195 26 229 60
rect 263 26 297 60
rect 331 26 365 60
rect 399 26 433 60
rect 467 26 501 60
rect 535 26 569 60
rect 603 26 637 60
rect 671 26 705 60
rect 739 26 773 60
rect 807 26 841 60
rect 875 26 909 60
rect 943 26 977 60
rect 1011 26 1045 60
rect 1079 26 1113 60
rect 1147 26 1181 60
rect 1215 26 1249 60
rect 1283 26 1317 60
rect 1351 26 1385 60
rect 1419 26 1453 60
rect 1487 26 1521 60
rect 1555 26 1589 60
rect 1623 26 1657 60
rect 1691 26 1725 60
rect 1759 26 1793 60
rect 1827 26 1861 60
rect 1895 26 1929 60
rect 1963 26 1997 60
rect 2031 26 2065 60
rect 2099 26 2133 60
rect 2167 26 2201 60
rect 2235 26 2269 60
rect 2303 26 2337 60
rect 2371 26 2395 60
<< mvnsubdiff >>
rect 67 798 101 832
rect 135 798 169 832
rect 203 798 237 832
rect 271 798 305 832
rect 339 798 373 832
rect 407 798 441 832
rect 475 798 509 832
rect 543 798 577 832
rect 611 798 645 832
rect 679 798 713 832
rect 747 798 781 832
rect 815 798 849 832
rect 883 798 917 832
rect 951 798 985 832
rect 1019 798 1053 832
rect 1087 798 1121 832
rect 1155 798 1189 832
rect 1223 798 1257 832
rect 1291 798 1325 832
rect 1359 798 1393 832
rect 1427 798 1461 832
rect 1495 798 1529 832
rect 1563 798 1597 832
rect 1631 798 1665 832
rect 1699 798 1733 832
rect 1767 798 1801 832
rect 1835 798 1869 832
rect 1903 798 1937 832
rect 1971 798 2005 832
rect 2039 798 2073 832
rect 2107 798 2141 832
rect 2175 798 2209 832
rect 2243 798 2277 832
rect 2311 798 2403 832
<< mvpsubdiffcont >>
rect 93 26 127 60
rect 161 26 195 60
rect 229 26 263 60
rect 297 26 331 60
rect 365 26 399 60
rect 433 26 467 60
rect 501 26 535 60
rect 569 26 603 60
rect 637 26 671 60
rect 705 26 739 60
rect 773 26 807 60
rect 841 26 875 60
rect 909 26 943 60
rect 977 26 1011 60
rect 1045 26 1079 60
rect 1113 26 1147 60
rect 1181 26 1215 60
rect 1249 26 1283 60
rect 1317 26 1351 60
rect 1385 26 1419 60
rect 1453 26 1487 60
rect 1521 26 1555 60
rect 1589 26 1623 60
rect 1657 26 1691 60
rect 1725 26 1759 60
rect 1793 26 1827 60
rect 1861 26 1895 60
rect 1929 26 1963 60
rect 1997 26 2031 60
rect 2065 26 2099 60
rect 2133 26 2167 60
rect 2201 26 2235 60
rect 2269 26 2303 60
rect 2337 26 2371 60
<< mvnsubdiffcont >>
rect 101 798 135 832
rect 169 798 203 832
rect 237 798 271 832
rect 305 798 339 832
rect 373 798 407 832
rect 441 798 475 832
rect 509 798 543 832
rect 577 798 611 832
rect 645 798 679 832
rect 713 798 747 832
rect 781 798 815 832
rect 849 798 883 832
rect 917 798 951 832
rect 985 798 1019 832
rect 1053 798 1087 832
rect 1121 798 1155 832
rect 1189 798 1223 832
rect 1257 798 1291 832
rect 1325 798 1359 832
rect 1393 798 1427 832
rect 1461 798 1495 832
rect 1529 798 1563 832
rect 1597 798 1631 832
rect 1665 798 1699 832
rect 1733 798 1767 832
rect 1801 798 1835 832
rect 1869 798 1903 832
rect 1937 798 1971 832
rect 2005 798 2039 832
rect 2073 798 2107 832
rect 2141 798 2175 832
rect 2209 798 2243 832
rect 2277 798 2311 832
<< poly >>
rect 2009 476 2421 492
rect 2009 442 2025 476
rect 2059 442 2095 476
rect 2129 442 2164 476
rect 2198 442 2233 476
rect 2267 442 2302 476
rect 2336 442 2371 476
rect 2405 442 2421 476
rect 2009 426 2421 442
rect 1853 368 2421 384
rect 1853 334 1869 368
rect 1903 334 1941 368
rect 1975 334 2013 368
rect 2047 334 2085 368
rect 2119 334 2157 368
rect 2191 334 2229 368
rect 2263 334 2300 368
rect 2334 334 2371 368
rect 2405 334 2421 368
rect 1853 318 2421 334
<< polycont >>
rect 2025 442 2059 476
rect 2095 442 2129 476
rect 2164 442 2198 476
rect 2233 442 2267 476
rect 2302 442 2336 476
rect 2371 442 2405 476
rect 1869 334 1903 368
rect 1941 334 1975 368
rect 2013 334 2047 368
rect 2085 334 2119 368
rect 2157 334 2191 368
rect 2229 334 2263 368
rect 2300 334 2334 368
rect 2371 334 2405 368
<< locali >>
rect 135 798 141 832
rect 203 798 215 832
rect 271 798 289 832
rect 339 798 363 832
rect 407 798 437 832
rect 475 798 509 832
rect 545 798 577 832
rect 619 798 645 832
rect 693 798 713 832
rect 767 798 781 832
rect 841 798 849 832
rect 915 798 917 832
rect 951 798 955 832
rect 1019 798 1029 832
rect 1087 798 1103 832
rect 1155 798 1177 832
rect 1223 798 1251 832
rect 1291 798 1325 832
rect 1359 798 1393 832
rect 1433 798 1461 832
rect 1507 798 1529 832
rect 1581 798 1597 832
rect 1655 798 1665 832
rect 1729 798 1733 832
rect 1767 798 1769 832
rect 1835 798 1843 832
rect 1903 798 1917 832
rect 1971 798 1991 832
rect 2039 798 2065 832
rect 2107 798 2138 832
rect 2175 798 2209 832
rect 2245 798 2277 832
rect 2318 798 2357 832
rect 2391 798 2403 832
rect 1963 694 2001 728
rect 2283 694 2321 728
rect 2118 532 2156 566
rect 2430 535 2468 569
rect 2009 442 2025 476
rect 2059 442 2095 476
rect 2145 442 2164 476
rect 2231 442 2233 476
rect 2267 442 2283 476
rect 2336 442 2368 476
rect 2405 442 2421 476
rect 1853 334 1869 368
rect 1903 334 1941 368
rect 1975 334 2013 368
rect 2060 334 2085 368
rect 2145 334 2157 368
rect 2191 334 2195 368
rect 2263 334 2279 368
rect 2334 334 2363 368
rect 2405 334 2421 368
rect 1962 232 2000 266
rect 2274 232 2312 266
rect 1806 132 1844 166
rect 2118 132 2156 166
rect 2430 132 2468 166
rect 69 26 81 60
rect 127 26 155 60
rect 195 26 229 60
rect 263 26 297 60
rect 337 26 365 60
rect 411 26 433 60
rect 485 26 501 60
rect 558 26 569 60
rect 631 26 637 60
rect 704 26 705 60
rect 739 26 743 60
rect 807 26 816 60
rect 875 26 889 60
rect 943 26 962 60
rect 1011 26 1035 60
rect 1079 26 1108 60
rect 1147 26 1181 60
rect 1215 26 1249 60
rect 1288 26 1317 60
rect 1361 26 1385 60
rect 1434 26 1453 60
rect 1507 26 1521 60
rect 1580 26 1589 60
rect 1653 26 1657 60
rect 1691 26 1692 60
rect 1759 26 1765 60
rect 1827 26 1838 60
rect 1895 26 1911 60
rect 1963 26 1984 60
rect 2031 26 2057 60
rect 2099 26 2130 60
rect 2167 26 2201 60
rect 2237 26 2269 60
rect 2310 26 2337 60
rect 2383 26 2395 60
<< viali >>
rect 67 798 101 832
rect 141 798 169 832
rect 169 798 175 832
rect 215 798 237 832
rect 237 798 249 832
rect 289 798 305 832
rect 305 798 323 832
rect 363 798 373 832
rect 373 798 397 832
rect 437 798 441 832
rect 441 798 471 832
rect 511 798 543 832
rect 543 798 545 832
rect 585 798 611 832
rect 611 798 619 832
rect 659 798 679 832
rect 679 798 693 832
rect 733 798 747 832
rect 747 798 767 832
rect 807 798 815 832
rect 815 798 841 832
rect 881 798 883 832
rect 883 798 915 832
rect 955 798 985 832
rect 985 798 989 832
rect 1029 798 1053 832
rect 1053 798 1063 832
rect 1103 798 1121 832
rect 1121 798 1137 832
rect 1177 798 1189 832
rect 1189 798 1211 832
rect 1251 798 1257 832
rect 1257 798 1285 832
rect 1325 798 1359 832
rect 1399 798 1427 832
rect 1427 798 1433 832
rect 1473 798 1495 832
rect 1495 798 1507 832
rect 1547 798 1563 832
rect 1563 798 1581 832
rect 1621 798 1631 832
rect 1631 798 1655 832
rect 1695 798 1699 832
rect 1699 798 1729 832
rect 1769 798 1801 832
rect 1801 798 1803 832
rect 1843 798 1869 832
rect 1869 798 1877 832
rect 1917 798 1937 832
rect 1937 798 1951 832
rect 1991 798 2005 832
rect 2005 798 2025 832
rect 2065 798 2073 832
rect 2073 798 2099 832
rect 2138 798 2141 832
rect 2141 798 2172 832
rect 2211 798 2243 832
rect 2243 798 2245 832
rect 2284 798 2311 832
rect 2311 798 2318 832
rect 2357 798 2391 832
rect 1929 694 1963 728
rect 2001 694 2035 728
rect 2249 694 2283 728
rect 2321 694 2355 728
rect 2084 532 2118 566
rect 2156 532 2190 566
rect 2396 535 2430 569
rect 2468 535 2502 569
rect 2025 442 2059 476
rect 2111 442 2129 476
rect 2129 442 2145 476
rect 2197 442 2198 476
rect 2198 442 2231 476
rect 2283 442 2302 476
rect 2302 442 2317 476
rect 2368 442 2371 476
rect 2371 442 2402 476
rect 1941 334 1975 368
rect 2026 334 2047 368
rect 2047 334 2060 368
rect 2111 334 2119 368
rect 2119 334 2145 368
rect 2195 334 2229 368
rect 2279 334 2300 368
rect 2300 334 2313 368
rect 2363 334 2371 368
rect 2371 334 2397 368
rect 1928 232 1962 266
rect 2000 232 2034 266
rect 2240 232 2274 266
rect 2312 232 2346 266
rect 1772 132 1806 166
rect 1844 132 1878 166
rect 2084 132 2118 166
rect 2156 132 2190 166
rect 2396 132 2430 166
rect 2468 132 2502 166
rect 81 26 93 60
rect 93 26 115 60
rect 155 26 161 60
rect 161 26 189 60
rect 229 26 263 60
rect 303 26 331 60
rect 331 26 337 60
rect 377 26 399 60
rect 399 26 411 60
rect 451 26 467 60
rect 467 26 485 60
rect 524 26 535 60
rect 535 26 558 60
rect 597 26 603 60
rect 603 26 631 60
rect 670 26 671 60
rect 671 26 704 60
rect 743 26 773 60
rect 773 26 777 60
rect 816 26 841 60
rect 841 26 850 60
rect 889 26 909 60
rect 909 26 923 60
rect 962 26 977 60
rect 977 26 996 60
rect 1035 26 1045 60
rect 1045 26 1069 60
rect 1108 26 1113 60
rect 1113 26 1142 60
rect 1181 26 1215 60
rect 1254 26 1283 60
rect 1283 26 1288 60
rect 1327 26 1351 60
rect 1351 26 1361 60
rect 1400 26 1419 60
rect 1419 26 1434 60
rect 1473 26 1487 60
rect 1487 26 1507 60
rect 1546 26 1555 60
rect 1555 26 1580 60
rect 1619 26 1623 60
rect 1623 26 1653 60
rect 1692 26 1725 60
rect 1725 26 1726 60
rect 1765 26 1793 60
rect 1793 26 1799 60
rect 1838 26 1861 60
rect 1861 26 1872 60
rect 1911 26 1929 60
rect 1929 26 1945 60
rect 1984 26 1997 60
rect 1997 26 2018 60
rect 2057 26 2065 60
rect 2065 26 2091 60
rect 2130 26 2133 60
rect 2133 26 2164 60
rect 2203 26 2235 60
rect 2235 26 2237 60
rect 2276 26 2303 60
rect 2303 26 2310 60
rect 2349 26 2371 60
rect 2371 26 2383 60
<< metal1 >>
rect 0 832 2540 838
rect 0 798 67 832
rect 101 798 141 832
rect 175 798 215 832
rect 249 798 289 832
rect 323 798 363 832
rect 397 798 437 832
rect 471 798 511 832
rect 545 798 585 832
rect 619 798 659 832
rect 693 798 733 832
rect 767 798 807 832
rect 841 798 881 832
rect 915 798 955 832
rect 989 798 1029 832
rect 1063 798 1103 832
rect 1137 798 1177 832
rect 1211 798 1251 832
rect 1285 798 1325 832
rect 1359 798 1399 832
rect 1433 798 1473 832
rect 1507 798 1547 832
rect 1581 798 1621 832
rect 1655 798 1695 832
rect 1729 798 1769 832
rect 1803 798 1843 832
rect 1877 798 1917 832
rect 1951 798 1991 832
rect 2025 798 2065 832
rect 2099 798 2138 832
rect 2172 798 2211 832
rect 2245 798 2284 832
rect 2318 798 2357 832
rect 2391 798 2540 832
rect 0 792 2540 798
rect 0 690 1738 792
tri 1738 758 1772 792 nw
rect 1917 728 1945 740
rect 1997 728 2009 740
rect 2061 728 2367 740
rect 1917 694 1929 728
rect 1997 694 2001 728
rect 2061 694 2249 728
rect 2283 694 2321 728
rect 2355 694 2367 728
tri 190 688 192 690 ne
rect 192 688 224 690
tri 192 656 224 688 ne
rect 894 688 926 690
tri 926 688 928 690 nw
rect 1917 688 1945 694
rect 1997 688 2009 694
rect 2061 688 2367 694
tri 894 656 926 688 nw
rect 2072 566 2248 578
rect 1845 482 1897 537
rect 2072 532 2084 566
rect 2118 532 2156 566
rect 2190 532 2248 566
rect 2072 526 2248 532
rect 2300 526 2312 578
rect 2364 569 2514 578
rect 2364 535 2396 569
rect 2430 535 2468 569
rect 2502 535 2514 569
rect 2364 526 2514 535
tri 1897 482 1931 516 sw
tri 894 476 898 480 sw
tri 1005 476 1009 480 se
rect 894 447 898 476
tri 898 447 927 476 sw
tri 976 447 1005 476 se
rect 1005 447 1009 476
rect 154 365 179 439
rect 310 361 339 437
rect 465 364 493 444
rect 625 358 648 425
rect 780 358 806 447
rect 894 446 927 447
tri 927 446 928 447 sw
tri 975 446 976 447 se
rect 976 446 1009 447
rect 1845 476 2414 482
rect 882 405 1026 446
rect 1845 442 2025 476
rect 2059 442 2111 476
rect 2145 442 2197 476
rect 2231 442 2283 476
rect 2317 442 2368 476
rect 2402 442 2414 476
rect 1845 436 2414 442
rect 879 394 1026 405
tri 1813 394 1827 408 sw
rect 879 354 1014 394
rect 1813 374 1827 394
tri 1827 374 1847 394 sw
tri 1221 372 1223 374 se
rect 1223 372 1247 374
tri 1217 368 1221 372 se
rect 1221 368 1247 372
rect 877 338 1014 354
tri 1187 338 1217 368 se
rect 1217 338 1247 368
rect 877 334 966 338
tri 966 334 970 338 nw
tri 1183 334 1187 338 se
rect 1187 334 1247 338
rect 877 328 960 334
tri 960 328 966 334 nw
tri 1177 328 1183 334 se
rect 1183 328 1247 334
tri 1564 328 1570 334 se
rect 1570 328 1622 372
rect 1688 368 2409 374
rect 1688 334 1941 368
rect 1975 334 2026 368
rect 2060 334 2111 368
rect 2145 334 2195 368
rect 2229 334 2279 368
rect 2313 334 2363 368
rect 2397 334 2409 368
rect 1688 328 2409 334
rect 877 310 942 328
tri 942 310 960 328 nw
tri 1159 310 1177 328 se
rect 1177 310 1229 328
tri 1229 310 1247 328 nw
tri 1546 310 1564 328 se
rect 1564 310 1628 328
rect 877 290 936 310
tri 936 304 942 310 nw
tri 1035 304 1041 310 se
rect 1041 304 1219 310
tri 1031 300 1035 304 se
rect 1035 300 1219 304
tri 1219 300 1229 310 nw
tri 1536 300 1546 310 se
rect 1546 300 1628 310
tri 1628 300 1656 328 nw
tri 1021 290 1031 300 se
rect 1031 290 1198 300
tri 997 266 1021 290 se
rect 1021 279 1198 290
tri 1198 279 1219 300 nw
rect 1466 290 1622 300
tri 1622 294 1628 300 nw
rect 1021 266 1075 279
tri 1075 266 1088 279 nw
rect 1466 275 1607 290
tri 1607 275 1622 290 nw
rect 1466 266 1598 275
tri 1598 266 1607 275 nw
rect 1916 266 1945 275
rect 1997 266 2009 275
rect 2061 266 2358 275
tri 985 254 997 266 se
rect 997 254 1057 266
tri 114 248 120 254 sw
tri 979 248 985 254 se
rect 985 248 1057 254
tri 1057 248 1075 266 nw
rect 1466 248 1580 266
tri 1580 248 1598 266 nw
rect 114 232 120 248
tri 120 232 136 248 sw
tri 963 232 979 248 se
rect 979 232 1041 248
tri 1041 232 1057 248 nw
rect 1916 232 1928 266
rect 1997 232 2000 266
rect 2061 232 2240 266
rect 2274 232 2312 266
rect 2346 232 2358 266
rect 114 223 136 232
tri 136 223 145 232 sw
tri 954 223 963 232 se
rect 963 223 1032 232
tri 1032 223 1041 232 nw
rect 1916 223 1945 232
rect 1997 223 2009 232
rect 2061 223 2358 232
rect 114 220 145 223
tri 145 220 148 223 sw
tri 951 220 954 223 se
rect 954 220 1029 223
tri 1029 220 1032 223 nw
rect 114 192 1001 220
tri 1001 192 1029 220 nw
rect 1760 166 2249 176
rect 0 66 1603 164
rect 1760 132 1772 166
rect 1806 132 1844 166
rect 1878 132 2084 166
rect 2118 132 2156 166
rect 2190 132 2249 166
rect 1760 124 2249 132
rect 2301 124 2313 176
rect 2365 166 2514 176
rect 2365 132 2396 166
rect 2430 132 2468 166
rect 2502 132 2514 166
rect 2365 124 2514 132
tri 1603 66 1637 100 sw
rect 0 60 2540 66
rect 0 26 81 60
rect 115 26 155 60
rect 189 26 229 60
rect 263 26 303 60
rect 337 26 377 60
rect 411 26 451 60
rect 485 26 524 60
rect 558 26 597 60
rect 631 26 670 60
rect 704 26 743 60
rect 777 26 816 60
rect 850 26 889 60
rect 923 26 962 60
rect 996 26 1035 60
rect 1069 26 1108 60
rect 1142 26 1181 60
rect 1215 26 1254 60
rect 1288 26 1327 60
rect 1361 26 1400 60
rect 1434 26 1473 60
rect 1507 26 1546 60
rect 1580 26 1619 60
rect 1653 26 1692 60
rect 1726 26 1765 60
rect 1799 26 1838 60
rect 1872 26 1911 60
rect 1945 26 1984 60
rect 2018 26 2057 60
rect 2091 26 2130 60
rect 2164 26 2203 60
rect 2237 26 2276 60
rect 2310 26 2349 60
rect 2383 26 2540 60
rect 0 0 2540 26
<< via1 >>
rect 1945 728 1997 740
rect 2009 728 2061 740
rect 1945 694 1963 728
rect 1963 694 1997 728
rect 2009 694 2035 728
rect 2035 694 2061 728
rect 1945 688 1997 694
rect 2009 688 2061 694
rect 2248 526 2300 578
rect 2312 526 2364 578
rect 1945 266 1997 275
rect 2009 266 2061 275
rect 1945 232 1962 266
rect 1962 232 1997 266
rect 2009 232 2034 266
rect 2034 232 2061 266
rect 1945 223 1997 232
rect 2009 223 2061 232
rect 2249 124 2301 176
rect 2313 124 2365 176
<< metal2 >>
rect 1939 688 1945 740
rect 1997 688 2009 740
rect 2061 688 2067 740
tri 1389 578 1392 581 ne
rect 1392 578 1423 581
tri 1392 547 1423 578 ne
rect 1475 578 1506 581
tri 1506 578 1509 581 nw
tri 1475 547 1506 578 nw
tri 1389 300 1423 334 se
rect 1939 275 1991 688
tri 1991 654 2025 688 nw
rect 2242 526 2248 578
rect 2300 526 2312 578
rect 2364 526 2371 578
tri 2285 492 2319 526 ne
tri 1991 275 2025 309 sw
rect 1939 223 1945 275
rect 1997 223 2009 275
rect 2061 223 2067 275
tri 2285 176 2319 210 se
rect 2319 176 2371 526
rect 2243 124 2249 176
rect 2301 124 2313 176
rect 2365 124 2371 176
use nfet_CDNS_52468879185815  nfet_CDNS_52468879185815_0
timestamp 1707688321
transform 1 0 1853 0 1 136
box -82 -32 650 182
use pfet_CDNS_52468879185816  pfet_CDNS_52468879185816_0
timestamp 1707688321
transform 1 0 2009 0 -1 724
box -119 -66 531 266
use sky130_fd_io__gpiovrefv2_hv_inv  sky130_fd_io__gpiovrefv2_hv_inv_0
timestamp 1707688321
transform 1 0 1624 0 1 100
box -244 0 338 690
use sky130_fd_io__gpiovrefv2_hv_nand2  sky130_fd_io__gpiovrefv2_hv_nand2_0
timestamp 1707688321
transform 1 0 468 0 1 100
box 0 0 494 690
use sky130_fd_io__gpiovrefv2_hv_nand3  sky130_fd_io__gpiovrefv2_hv_nand3_0
timestamp 1707688321
transform -1 0 650 0 1 100
box 0 0 650 690
use sky130_fd_io__gpiovrefv2_hv_nor2  sky130_fd_io__gpiovrefv2_hv_nor2_0
timestamp 1707688321
transform 1 0 890 0 1 100
box 0 0 806 690
<< labels >>
flabel metal1 s 2357 132 2463 163 3 FreeSans 200 0 0 0 vrefout
port 1 nsew
flabel metal1 s 74 10 418 124 3 FreeSans 200 0 0 0 vssd
port 2 nsew
flabel metal1 s 2009 698 2128 735 3 FreeSans 200 0 0 0 vrefin
port 3 nsew
flabel metal1 s 153 728 385 818 3 FreeSans 200 0 0 0 vddio_q
port 4 nsew
flabel metal1 s 780 358 806 447 3 FreeSans 200 0 0 0 in3
port 5 nsew
flabel metal1 s 625 358 648 425 3 FreeSans 200 0 0 0 in4
port 6 nsew
flabel metal1 s 465 364 493 444 3 FreeSans 200 0 0 0 in2
port 7 nsew
flabel metal1 s 310 361 339 437 3 FreeSans 200 0 0 0 in1
port 8 nsew
flabel metal1 s 154 365 179 439 3 FreeSans 200 0 0 0 in0
port 9 nsew
<< properties >>
string GDS_END 25758212
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25740504
string path 48.475 17.850 51.675 17.850 
<< end >>
