##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 18:03:01 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO W_IO
  CLASS BLOCK ;
  SIZE 69.9200 BY 219.6400 ;
  FOREIGN W_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2207 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5676 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.72 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 84.7600 69.9200 84.9000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8301 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.53 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 83.4000 69.9200 83.5400 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.32 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 81.7000 69.9200 81.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.968 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 80.3400 69.9200 80.4800 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4713 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.252 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 96.6600 69.9200 96.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.24 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 94.9600 69.9200 95.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.6001 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.896 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 93.6000 69.9200 93.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.36 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 92.2400 69.9200 92.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.0011 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.901 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 90.5400 69.9200 90.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2809 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.6628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.672 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 89.1800 69.9200 89.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9421 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 87.8200 69.9200 87.9600 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 86.1200 69.9200 86.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4881 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 108.2200 69.9200 108.3600 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.2848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.656 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 106.8600 69.9200 107.0000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.5049 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.42 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 105.5000 69.9200 105.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.7128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.272 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 103.8000 69.9200 103.9400 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3897 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.332 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 102.4400 69.9200 102.5800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.7658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.888 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 101.0800 69.9200 101.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2451 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.24 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 99.3800 69.9200 99.5200 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4313 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 98.0200 69.9200 98.1600 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2073 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.959 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.356 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 132.0200 69.9200 132.1600 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5893 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.288 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 130.3200 69.9200 130.4600 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2683 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.7748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 128.9600 69.9200 129.1000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.2288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.024 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 127.6000 69.9200 127.7400 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.12 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.482 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 125.9000 69.9200 126.0400 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9861 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 124.5400 69.9200 124.6800 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4237 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.48 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 123.1800 69.9200 123.3200 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 121.4800 69.9200 121.6200 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.698 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 120.1200 69.9200 120.2600 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.198 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 118.7600 69.9200 118.9000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.373 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 117.0600 69.9200 117.2000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.96 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.564 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 115.7000 69.9200 115.8400 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.296 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 114.3400 69.9200 114.4800 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.72 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 112.6400 69.9200 112.7800 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.32 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 111.2800 69.9200 111.4200 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0201 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.0068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.84 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 109.9200 69.9200 110.0600 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4405 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.098 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 149.7000 69.9200 149.8400 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.3208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.848 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 148.0000 69.9200 148.1400 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.4696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.112 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 146.6400 69.9200 146.7800 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7457 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.9868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.4 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 145.2800 69.9200 145.4200 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0709 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 143.5800 69.9200 143.7200 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.3438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.304 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 142.2200 69.9200 142.3600 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.3117 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.454 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 140.8600 69.9200 141.0000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.048 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 139.1600 69.9200 139.3000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0541 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5185 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.7408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.088 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 137.8000 69.9200 137.9400 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.5698 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 62.176 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 136.4400 69.9200 136.5800 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0065 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 134.4000 69.9200 134.5400 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5081 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 133.3800 69.9200 133.5200 ;
    END
  END E6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3155 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4695 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met2  ;
    ANTENNAMAXAREACAR 38.5257 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 186.373 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.104472 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 14.0400 69.9200 14.1800 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.4348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.712 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 89.8814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 429.686 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 12.6800 69.9200 12.8200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.416 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 49.8946 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 260.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.267073 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 11.3200 69.9200 11.4600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7149 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.47 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 175.967 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 918.893 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 9.9600 69.9200 10.1000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.4275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.491 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3284 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.488 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 25.9400 69.9200 26.0800 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2851 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 24.5800 69.9200 24.7200 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.805 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.0526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.408 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 22.8800 69.9200 23.0200 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5145 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.8685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.0933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.3547 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.024 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 21.5200 69.9200 21.6600 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2269 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.0181 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.9195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8732 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 20.1600 69.9200 20.3000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3249 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.228 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 18.4600 69.9200 18.6000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5731 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.7443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.5505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9432 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 17.1000 69.9200 17.2400 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9081 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.3599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.6285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.936 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 15.7400 69.9200 15.8800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4275 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.1418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7596 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.192 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 37.8400 69.9200 37.9800 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4505 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.192 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 36.1400 69.9200 36.2800 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4605 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2547 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8981 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 34.7800 69.9200 34.9200 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.2758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 33.4200 69.9200 33.5600 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.8 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 31.7200 69.9200 31.8600 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.1245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9432 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7062 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.509 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 30.3600 69.9200 30.5000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.8259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 29.0000 69.9200 29.1400 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8705 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1268 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 27.3000 69.9200 27.4400 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6845 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.1401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.5295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.242 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 61.3000 69.9200 61.4400 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9421 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.137 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.272 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 59.9400 69.9200 60.0800 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.403 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.6018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.68 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 58.2400 69.9200 58.3800 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.424 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 56.8800 69.9200 57.0200 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.3896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 55.1800 69.9200 55.3200 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0369 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 53.8200 69.9200 53.9600 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5028 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.152 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 52.4600 69.9200 52.6000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8405 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.31 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.098 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 51.1000 69.9200 51.2400 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6501 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.4648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 49.4000 69.9200 49.5400 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1269 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.389 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.4905 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.552 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 48.0400 69.9200 48.1800 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.592 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 46.6800 69.9200 46.8200 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.608 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 44.9800 69.9200 45.1200 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.8468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.32 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 43.6200 69.9200 43.7600 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3117 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.6395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 42.2600 69.9200 42.4000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2061 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.9225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.808 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 40.5600 69.9200 40.7000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1657 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 64.554 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 39.2000 69.9200 39.3400 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9113 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7685 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.368 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 78.9800 69.9200 79.1200 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 77.6200 69.9200 77.7600 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1661 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.2627 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.6805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.768 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 75.9200 69.9200 76.0600 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5049 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.488 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 74.5600 69.9200 74.7000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.134 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.6484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.318 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 73.2000 69.9200 73.3400 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.6214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.392 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 71.5000 69.9200 71.6400 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0777 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.2805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.7254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.296 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 70.1400 69.9200 70.2800 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6545 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.1015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.7558 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.168 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 68.7800 69.9200 68.9200 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8777 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.1412 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.8243 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.656 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 66.7400 69.9200 66.8800 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.1983 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.464 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 65.7200 69.9200 65.8600 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.931 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.288 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 64.3600 69.9200 64.5000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5841 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 69.3250 62.6600 69.9200 62.8000 ;
    END
  END W6END[0]
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2851 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8938 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.904 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 100.4000 0.5950 100.5400 ;
    END
  END A_I_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.0395 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.056 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 98.3600 0.5950 98.5000 ;
    END
  END A_T_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.243 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.854 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0675 LAYER via  ;
    ANTENNADIFFAREA 0.954 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.9652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.922 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met2  ;
    ANTENNAMAXAREACAR 26.8269 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 95.9800 0.5950 96.1200 ;
    END
  END A_O_top
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.8566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 12.2191 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.4966 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END UserCLK
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1337 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5235 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.4200 0.5950 84.5600 ;
    END
  END B_I_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.4083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.8705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.7798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.296 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 82.0400 0.5950 82.1800 ;
    END
  END B_T_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.08 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.618 LAYER met4  ;
    ANTENNAMAXAREACAR 47.053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 232.736 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.780683 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 80.0000 0.5950 80.1400 ;
    END
  END B_O_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7131 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.461 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 102.7800 0.5950 102.9200 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.4583 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.187 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.1600 0.5950 105.3000 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1493 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.1739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.5805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.1918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.16 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 107.5400 0.5950 107.6800 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1353 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.4008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.608 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.9200 0.5950 110.0600 ;
    END
  END A_config_C_bit3
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.5017 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.404 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 86.8000 0.5950 86.9400 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.9661 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.726 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 89.1800 0.5950 89.3200 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8269 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.7199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.496 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 91.2200 0.5950 91.3600 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.6000 0.5950 93.7400 ;
    END
  END B_config_C_bit3
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 25.3686 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.019 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.60386 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 209.3500 0.8000 209.6500 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 17.5691 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 84.0652 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 207.5200 0.8000 207.8200 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.4672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.624 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 31.0245 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.185 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6900 0.8000 205.9900 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.7392 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 29.1645 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.286 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 203.8600 0.8000 204.1600 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 21.3368 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.027 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 202.0300 0.8000 202.3300 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.4578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1498 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.661 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 200.2000 0.8000 200.5000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.9164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 39.2231 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 194.22 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.635306 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 198.3700 0.8000 198.6700 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0001 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.128 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 20.7784 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 104.08 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5400 0.8000 196.8400 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4756 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.6558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 35.6897 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 183.024 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 195.3200 0.8000 195.6200 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.9978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 34.0864 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.953 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.381305 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4900 0.8000 193.7900 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 35.4696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 53.6849 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 274.945 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 191.6600 0.8000 191.9600 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.5596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.5448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 33.1422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.863 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 189.8300 0.8000 190.1300 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.9596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 44.6664 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 231.502 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 188.0000 0.8000 188.3000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7446 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.5648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met4  ;
    ANTENNAMAXAREACAR 37.4718 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.225 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.522814 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 186.1700 0.8000 186.4700 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.1404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.744 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 25.95 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.837 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.493797 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3400 0.8000 184.6400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9112 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.992 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 22.5585 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 112.231 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.412011 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 182.5100 0.8000 182.8100 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 14.3145 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 68.7143 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2900 0.8000 181.5900 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 20.1747 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.9812 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.352288 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 179.4600 0.8000 179.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.256 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 16.0333 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 77.5575 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 177.6300 0.8000 177.9300 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.696 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 10.458 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.5965 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.8000 0.8000 176.1000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 12.1528 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 58.4534 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 173.9700 0.8000 174.2700 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 9.07778 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 42.4673 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.356071 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1400 0.8000 172.4400 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 27.434 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.678 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 170.3100 0.8000 170.6100 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.567 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 73.0792 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 364.962 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 168.4800 0.8000 168.7800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.632 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 18.9304 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 91.9638 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 167.2600 0.8000 167.5600 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 22.4922 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 108.486 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 165.4300 0.8000 165.7300 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9996 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.5656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 38.5837 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 200.396 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 163.6000 0.8000 163.9000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.4708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 44.3882 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.571 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 161.7700 0.8000 162.0700 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.0528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 96.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 30.4886 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 154.665 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.388871 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9400 0.8000 160.2400 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.7998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4159 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.638 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.530381 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 158.1100 0.8000 158.4100 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 29.8418 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 149.424 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.2800 0.8000 156.5800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.328 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2195 LAYER met3  ;
    ANTENNAMAXAREACAR 17.7175 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 87.5456 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.49758 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 155.0600 0.8000 155.3600 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.9414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 209.3500 69.9200 209.6500 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.4484 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 207.5200 69.9200 207.8200 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.6304 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.024 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 205.6900 69.9200 205.9900 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.48 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 203.8600 69.9200 204.1600 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.9328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 202.0300 69.9200 202.3300 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.944 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 200.2000 69.9200 200.5000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5846 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.4228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.392 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 198.3700 69.9200 198.6700 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 196.5400 69.9200 196.8400 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2089 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.4508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.208 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 195.3200 69.9200 195.6200 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1066 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.4528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.552 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 193.4900 69.9200 193.7900 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 191.6600 69.9200 191.9600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.1718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.72 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 189.8300 69.9200 190.1300 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.7746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.072 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 188.0000 69.9200 188.3000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.4946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.272 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 186.1700 69.9200 186.4700 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 184.3400 69.9200 184.6400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 182.5100 69.9200 182.8100 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 181.2900 69.9200 181.5900 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.5584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 179.4600 69.9200 179.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.7224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 177.6300 69.9200 177.9300 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 175.8000 69.9200 176.1000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.016 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 173.9700 69.9200 174.2700 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.7904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 172.1400 69.9200 172.4400 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.9438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.504 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 170.3100 69.9200 170.6100 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9244 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 168.4800 69.9200 168.7800 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.7698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.576 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 167.2600 69.9200 167.5600 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.3714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 165.4300 69.9200 165.7300 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.8628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.072 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 163.6000 69.9200 163.9000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.304 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 161.1600 69.9200 161.4600 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 159.9400 69.9200 160.2400 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8326 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.264 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 158.1100 69.9200 158.4100 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 156.2800 69.9200 156.5800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 69.1200 155.0600 69.9200 155.3600 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.22155 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.7131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 0.0000 59.6550 0.3300 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.87465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.029 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.678 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.35798 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.3953 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.7250 0.0000 56.8950 0.3300 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.3176 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.514 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 8.80485 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 42.7933 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 53.9650 0.0000 54.1350 0.3300 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.02236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.71717 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 51.2050 0.0000 51.3750 0.3300 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.55 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.39569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 10.5838 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 48.4450 0.0000 48.6150 0.3300 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.8428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.632 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.493 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.7208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.648 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 64.7162 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.071 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 40.1650 0.0000 40.3350 0.3300 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.7818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 64.2063 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 340.094 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 37.4050 0.0000 37.5750 0.3300 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 30.5924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 152.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 41.816 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 207.527 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 34.6450 0.0000 34.8150 0.3300 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.40013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.60606 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 0.0000 32.0550 0.3300 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.4832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 137.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 38.3696 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 190.453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 29.5850 0.0000 29.7550 0.3300 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.988 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.9802 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.5064 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.99596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.58519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.0650 0.0000 24.2350 0.3300 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.0576 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.17 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 38.9635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 193.423 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 21.3050 0.0000 21.4750 0.3300 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.1444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.648 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 7.22478 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 34.8929 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 18.5450 0.0000 18.7150 0.3300 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.37993 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.5051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.7850 0.0000 15.9550 0.3300 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2972 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 24.5885 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 121.062 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.4225 LAYER met2  ;
    ANTENNAMAXAREACAR 22.3045 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.923 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.569907 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.3747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.464 LAYER met3  ;
    ANTENNAGATEAREA 3.0585 LAYER met3  ;
    ANTENNAMAXAREACAR 25.3696 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.423 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 13.0250 0.0000 13.1950 0.3300 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.9619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 78.5505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2464 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 95.9309 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.12 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.414908 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.6614 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.592 LAYER met3  ;
    ANTENNAGATEAREA 3.0585 LAYER met3  ;
    ANTENNAMAXAREACAR 25.04 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 121.954 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.587921 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 25.6858 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.608535 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.6035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.4745 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.908 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0265 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 101.687 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.6991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.792 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 32.785 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 113.758 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 7.5050 0.0000 7.6750 0.3300 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 30.6122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 149.884 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.4895 LAYER met2  ;
    ANTENNAMAXAREACAR 29.7067 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 142.162 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.655451 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.44 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 30.9474 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 148.869 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.655451 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 0.0000 5.3750 0.3300 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.6228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 219.3100 59.6550 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.9055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 219.3100 56.4350 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 219.3100 53.6750 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3763 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.6228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 219.3100 50.9150 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2162 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0035 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.2459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.3878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 219.3100 48.1550 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 44.7650 219.3100 44.9350 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.0050 219.3100 42.1750 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.782 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.942 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.2450 219.3100 39.4150 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.466 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 219.3100 36.6550 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.7250 219.3100 33.8950 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.25 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 219.3100 30.6750 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.5795 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.7265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.2548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 219.3100 27.9150 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.7427 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 219.3100 25.1550 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 219.3100 22.3950 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 219.3100 19.6350 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.7727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.6298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.2450 219.3100 16.4150 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.4036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.9 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 219.3100 13.6550 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.2032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 100.898 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.7250 219.3100 10.8950 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.9548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 7.9650 219.3100 8.1350 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.8348 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.688 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.588 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 219.3100 5.3750 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 3.3900 5.3300 66.5300 6.3300 ;
        RECT 3.3900 212.6300 66.5300 213.6300 ;
        RECT 3.3900 12.3400 4.3900 12.8200 ;
        RECT 3.3900 23.2200 4.3900 23.7000 ;
        RECT 3.3900 17.7800 4.3900 18.2600 ;
        RECT 3.3900 39.5400 4.3900 40.0200 ;
        RECT 3.3900 34.1000 4.3900 34.5800 ;
        RECT 3.3900 28.6600 4.3900 29.1400 ;
        RECT 3.3900 50.4200 4.3900 50.9000 ;
        RECT 3.3900 44.9800 4.3900 45.4600 ;
        RECT 3.3900 66.7400 4.3900 67.2200 ;
        RECT 3.3900 61.3000 4.3900 61.7800 ;
        RECT 3.3900 55.8600 4.3900 56.3400 ;
        RECT 3.3900 77.6200 4.3900 78.1000 ;
        RECT 3.3900 72.1800 4.3900 72.6600 ;
        RECT 3.3900 93.9400 4.3900 94.4200 ;
        RECT 3.3900 88.5000 4.3900 88.9800 ;
        RECT 3.3900 83.0600 4.3900 83.5400 ;
        RECT 3.3900 104.8200 4.3900 105.3000 ;
        RECT 3.3900 99.3800 4.3900 99.8600 ;
        RECT 65.5300 12.3400 66.5300 12.8200 ;
        RECT 65.5300 23.2200 66.5300 23.7000 ;
        RECT 65.5300 17.7800 66.5300 18.2600 ;
        RECT 65.5300 39.5400 66.5300 40.0200 ;
        RECT 65.5300 34.1000 66.5300 34.5800 ;
        RECT 65.5300 28.6600 66.5300 29.1400 ;
        RECT 65.5300 50.4200 66.5300 50.9000 ;
        RECT 65.5300 44.9800 66.5300 45.4600 ;
        RECT 65.5300 66.7400 66.5300 67.2200 ;
        RECT 65.5300 61.3000 66.5300 61.7800 ;
        RECT 65.5300 55.8600 66.5300 56.3400 ;
        RECT 65.5300 77.6200 66.5300 78.1000 ;
        RECT 65.5300 72.1800 66.5300 72.6600 ;
        RECT 65.5300 93.9400 66.5300 94.4200 ;
        RECT 65.5300 88.5000 66.5300 88.9800 ;
        RECT 65.5300 83.0600 66.5300 83.5400 ;
        RECT 65.5300 104.8200 66.5300 105.3000 ;
        RECT 65.5300 99.3800 66.5300 99.8600 ;
        RECT 3.3900 164.6600 4.3900 165.1400 ;
        RECT 3.3900 121.1400 4.3900 121.6200 ;
        RECT 3.3900 115.7000 4.3900 116.1800 ;
        RECT 3.3900 110.2600 4.3900 110.7400 ;
        RECT 3.3900 132.0200 4.3900 132.5000 ;
        RECT 3.3900 126.5800 4.3900 127.0600 ;
        RECT 3.3900 148.3400 4.3900 148.8200 ;
        RECT 3.3900 142.9000 4.3900 143.3800 ;
        RECT 3.3900 137.4600 4.3900 137.9400 ;
        RECT 3.3900 159.2200 4.3900 159.7000 ;
        RECT 3.3900 153.7800 4.3900 154.2600 ;
        RECT 3.3900 191.8600 4.3900 192.3400 ;
        RECT 3.3900 175.5400 4.3900 176.0200 ;
        RECT 3.3900 170.1000 4.3900 170.5800 ;
        RECT 3.3900 186.4200 4.3900 186.9000 ;
        RECT 3.3900 180.9800 4.3900 181.4600 ;
        RECT 3.3900 202.7400 4.3900 203.2200 ;
        RECT 3.3900 197.3000 4.3900 197.7800 ;
        RECT 3.3900 208.1800 4.3900 208.6600 ;
        RECT 65.5300 164.6600 66.5300 165.1400 ;
        RECT 65.5300 121.1400 66.5300 121.6200 ;
        RECT 65.5300 115.7000 66.5300 116.1800 ;
        RECT 65.5300 110.2600 66.5300 110.7400 ;
        RECT 65.5300 132.0200 66.5300 132.5000 ;
        RECT 65.5300 126.5800 66.5300 127.0600 ;
        RECT 65.5300 148.3400 66.5300 148.8200 ;
        RECT 65.5300 142.9000 66.5300 143.3800 ;
        RECT 65.5300 137.4600 66.5300 137.9400 ;
        RECT 65.5300 159.2200 66.5300 159.7000 ;
        RECT 65.5300 153.7800 66.5300 154.2600 ;
        RECT 65.5300 191.8600 66.5300 192.3400 ;
        RECT 65.5300 175.5400 66.5300 176.0200 ;
        RECT 65.5300 170.1000 66.5300 170.5800 ;
        RECT 65.5300 186.4200 66.5300 186.9000 ;
        RECT 65.5300 180.9800 66.5300 181.4600 ;
        RECT 65.5300 202.7400 66.5300 203.2200 ;
        RECT 65.5300 197.3000 66.5300 197.7800 ;
        RECT 65.5300 208.1800 66.5300 208.6600 ;
      LAYER met4 ;
        RECT 3.3900 5.3300 4.3900 213.6300 ;
        RECT 65.5300 5.3300 66.5300 213.6300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5900 3.5300 68.3300 4.5300 ;
        RECT 1.5900 214.4300 68.3300 215.4300 ;
        RECT 1.5900 9.6200 2.5900 10.1000 ;
        RECT 1.5900 25.9400 2.5900 26.4200 ;
        RECT 1.5900 20.5000 2.5900 20.9800 ;
        RECT 1.5900 15.0600 2.5900 15.5400 ;
        RECT 1.5900 36.8200 2.5900 37.3000 ;
        RECT 1.5900 31.3800 2.5900 31.8600 ;
        RECT 1.5900 53.1400 2.5900 53.6200 ;
        RECT 1.5900 47.7000 2.5900 48.1800 ;
        RECT 1.5900 42.2600 2.5900 42.7400 ;
        RECT 1.5900 64.0200 2.5900 64.5000 ;
        RECT 1.5900 58.5800 2.5900 59.0600 ;
        RECT 1.5900 80.3400 2.5900 80.8200 ;
        RECT 1.5900 74.9000 2.5900 75.3800 ;
        RECT 1.5900 69.4600 2.5900 69.9400 ;
        RECT 1.5900 91.2200 2.5900 91.7000 ;
        RECT 1.5900 85.7800 2.5900 86.2600 ;
        RECT 1.5900 107.5400 2.5900 108.0200 ;
        RECT 1.5900 102.1000 2.5900 102.5800 ;
        RECT 1.5900 96.6600 2.5900 97.1400 ;
        RECT 67.3300 9.6200 68.3300 10.1000 ;
        RECT 67.3300 25.9400 68.3300 26.4200 ;
        RECT 67.3300 20.5000 68.3300 20.9800 ;
        RECT 67.3300 15.0600 68.3300 15.5400 ;
        RECT 67.3300 36.8200 68.3300 37.3000 ;
        RECT 67.3300 31.3800 68.3300 31.8600 ;
        RECT 67.3300 53.1400 68.3300 53.6200 ;
        RECT 67.3300 47.7000 68.3300 48.1800 ;
        RECT 67.3300 42.2600 68.3300 42.7400 ;
        RECT 67.3300 64.0200 68.3300 64.5000 ;
        RECT 67.3300 58.5800 68.3300 59.0600 ;
        RECT 67.3300 80.3400 68.3300 80.8200 ;
        RECT 67.3300 74.9000 68.3300 75.3800 ;
        RECT 67.3300 69.4600 68.3300 69.9400 ;
        RECT 67.3300 91.2200 68.3300 91.7000 ;
        RECT 67.3300 85.7800 68.3300 86.2600 ;
        RECT 67.3300 107.5400 68.3300 108.0200 ;
        RECT 67.3300 102.1000 68.3300 102.5800 ;
        RECT 67.3300 96.6600 68.3300 97.1400 ;
        RECT 1.5900 118.4200 2.5900 118.9000 ;
        RECT 1.5900 112.9800 2.5900 113.4600 ;
        RECT 1.5900 134.7400 2.5900 135.2200 ;
        RECT 1.5900 129.3000 2.5900 129.7800 ;
        RECT 1.5900 123.8600 2.5900 124.3400 ;
        RECT 1.5900 145.6200 2.5900 146.1000 ;
        RECT 1.5900 140.1800 2.5900 140.6600 ;
        RECT 1.5900 161.9400 2.5900 162.4200 ;
        RECT 1.5900 156.5000 2.5900 156.9800 ;
        RECT 1.5900 151.0600 2.5900 151.5400 ;
        RECT 1.5900 178.2600 2.5900 178.7400 ;
        RECT 1.5900 172.8200 2.5900 173.3000 ;
        RECT 1.5900 167.3800 2.5900 167.8600 ;
        RECT 1.5900 189.1400 2.5900 189.6200 ;
        RECT 1.5900 183.7000 2.5900 184.1800 ;
        RECT 1.5900 205.4600 2.5900 205.9400 ;
        RECT 1.5900 200.0200 2.5900 200.5000 ;
        RECT 1.5900 194.5800 2.5900 195.0600 ;
        RECT 67.3300 118.4200 68.3300 118.9000 ;
        RECT 67.3300 112.9800 68.3300 113.4600 ;
        RECT 67.3300 134.7400 68.3300 135.2200 ;
        RECT 67.3300 129.3000 68.3300 129.7800 ;
        RECT 67.3300 123.8600 68.3300 124.3400 ;
        RECT 67.3300 145.6200 68.3300 146.1000 ;
        RECT 67.3300 140.1800 68.3300 140.6600 ;
        RECT 67.3300 161.9400 68.3300 162.4200 ;
        RECT 67.3300 156.5000 68.3300 156.9800 ;
        RECT 67.3300 151.0600 68.3300 151.5400 ;
        RECT 67.3300 178.2600 68.3300 178.7400 ;
        RECT 67.3300 172.8200 68.3300 173.3000 ;
        RECT 67.3300 167.3800 68.3300 167.8600 ;
        RECT 67.3300 189.1400 68.3300 189.6200 ;
        RECT 67.3300 183.7000 68.3300 184.1800 ;
        RECT 67.3300 205.4600 68.3300 205.9400 ;
        RECT 67.3300 200.0200 68.3300 200.5000 ;
        RECT 67.3300 194.5800 68.3300 195.0600 ;
      LAYER met4 ;
        RECT 1.5900 3.5300 2.5900 215.4300 ;
        RECT 67.3300 3.5300 68.3300 215.4300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 59.8250 219.1400 69.9200 219.6400 ;
      RECT 56.6050 219.1400 59.3150 219.6400 ;
      RECT 53.8450 219.1400 56.0950 219.6400 ;
      RECT 51.0850 219.1400 53.3350 219.6400 ;
      RECT 48.3250 219.1400 50.5750 219.6400 ;
      RECT 45.1050 219.1400 47.8150 219.6400 ;
      RECT 42.3450 219.1400 44.5950 219.6400 ;
      RECT 39.5850 219.1400 41.8350 219.6400 ;
      RECT 36.8250 219.1400 39.0750 219.6400 ;
      RECT 34.0650 219.1400 36.3150 219.6400 ;
      RECT 30.8450 219.1400 33.5550 219.6400 ;
      RECT 28.0850 219.1400 30.3350 219.6400 ;
      RECT 25.3250 219.1400 27.5750 219.6400 ;
      RECT 22.5650 219.1400 24.8150 219.6400 ;
      RECT 19.8050 219.1400 22.0550 219.6400 ;
      RECT 16.5850 219.1400 19.2950 219.6400 ;
      RECT 13.8250 219.1400 16.0750 219.6400 ;
      RECT 11.0650 219.1400 13.3150 219.6400 ;
      RECT 8.3050 219.1400 10.5550 219.6400 ;
      RECT 5.5450 219.1400 7.7950 219.6400 ;
      RECT 0.0000 219.1400 5.0350 219.6400 ;
      RECT 0.0000 0.5000 69.9200 219.1400 ;
      RECT 59.8250 0.0000 69.9200 0.5000 ;
      RECT 57.0650 0.0000 59.3150 0.5000 ;
      RECT 54.3050 0.0000 56.5550 0.5000 ;
      RECT 51.5450 0.0000 53.7950 0.5000 ;
      RECT 48.7850 0.0000 51.0350 0.5000 ;
      RECT 46.0250 0.0000 48.2750 0.5000 ;
      RECT 43.2650 0.0000 45.5150 0.5000 ;
      RECT 40.5050 0.0000 42.7550 0.5000 ;
      RECT 37.7450 0.0000 39.9950 0.5000 ;
      RECT 34.9850 0.0000 37.2350 0.5000 ;
      RECT 32.2250 0.0000 34.4750 0.5000 ;
      RECT 29.9250 0.0000 31.7150 0.5000 ;
      RECT 27.1650 0.0000 29.4150 0.5000 ;
      RECT 24.4050 0.0000 26.6550 0.5000 ;
      RECT 21.6450 0.0000 23.8950 0.5000 ;
      RECT 18.8850 0.0000 21.1350 0.5000 ;
      RECT 16.1250 0.0000 18.3750 0.5000 ;
      RECT 13.3650 0.0000 15.6150 0.5000 ;
      RECT 10.6050 0.0000 12.8550 0.5000 ;
      RECT 7.8450 0.0000 10.0950 0.5000 ;
      RECT 5.5450 0.0000 7.3350 0.5000 ;
      RECT 0.0000 0.0000 5.0350 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 149.9800 69.9200 219.6400 ;
      RECT 0.0000 149.5600 69.1850 149.9800 ;
      RECT 0.0000 148.2800 69.9200 149.5600 ;
      RECT 0.0000 147.8600 69.1850 148.2800 ;
      RECT 0.0000 146.9200 69.9200 147.8600 ;
      RECT 0.0000 146.5000 69.1850 146.9200 ;
      RECT 0.0000 145.5600 69.9200 146.5000 ;
      RECT 0.0000 145.1400 69.1850 145.5600 ;
      RECT 0.0000 143.8600 69.9200 145.1400 ;
      RECT 0.0000 143.4400 69.1850 143.8600 ;
      RECT 0.0000 142.5000 69.9200 143.4400 ;
      RECT 0.0000 142.0800 69.1850 142.5000 ;
      RECT 0.0000 141.1400 69.9200 142.0800 ;
      RECT 0.0000 140.7200 69.1850 141.1400 ;
      RECT 0.0000 139.4400 69.9200 140.7200 ;
      RECT 0.0000 139.0200 69.1850 139.4400 ;
      RECT 0.0000 138.0800 69.9200 139.0200 ;
      RECT 0.0000 137.6600 69.1850 138.0800 ;
      RECT 0.0000 136.7200 69.9200 137.6600 ;
      RECT 0.0000 136.3000 69.1850 136.7200 ;
      RECT 0.0000 134.6800 69.9200 136.3000 ;
      RECT 0.0000 134.2600 69.1850 134.6800 ;
      RECT 0.0000 133.6600 69.9200 134.2600 ;
      RECT 0.0000 133.2400 69.1850 133.6600 ;
      RECT 0.0000 132.3000 69.9200 133.2400 ;
      RECT 0.0000 131.8800 69.1850 132.3000 ;
      RECT 0.0000 130.6000 69.9200 131.8800 ;
      RECT 0.0000 130.1800 69.1850 130.6000 ;
      RECT 0.0000 129.2400 69.9200 130.1800 ;
      RECT 0.0000 128.8200 69.1850 129.2400 ;
      RECT 0.0000 127.8800 69.9200 128.8200 ;
      RECT 0.0000 127.4600 69.1850 127.8800 ;
      RECT 0.0000 126.1800 69.9200 127.4600 ;
      RECT 0.0000 125.7600 69.1850 126.1800 ;
      RECT 0.0000 124.8200 69.9200 125.7600 ;
      RECT 0.0000 124.4000 69.1850 124.8200 ;
      RECT 0.0000 123.4600 69.9200 124.4000 ;
      RECT 0.0000 123.0400 69.1850 123.4600 ;
      RECT 0.0000 121.7600 69.9200 123.0400 ;
      RECT 0.0000 121.3400 69.1850 121.7600 ;
      RECT 0.0000 120.4000 69.9200 121.3400 ;
      RECT 0.0000 119.9800 69.1850 120.4000 ;
      RECT 0.0000 119.0400 69.9200 119.9800 ;
      RECT 0.0000 118.6200 69.1850 119.0400 ;
      RECT 0.0000 117.3400 69.9200 118.6200 ;
      RECT 0.0000 116.9200 69.1850 117.3400 ;
      RECT 0.0000 115.9800 69.9200 116.9200 ;
      RECT 0.0000 115.5600 69.1850 115.9800 ;
      RECT 0.0000 114.6200 69.9200 115.5600 ;
      RECT 0.0000 114.2000 69.1850 114.6200 ;
      RECT 0.0000 112.9200 69.9200 114.2000 ;
      RECT 0.0000 112.5000 69.1850 112.9200 ;
      RECT 0.0000 111.5600 69.9200 112.5000 ;
      RECT 0.0000 111.1400 69.1850 111.5600 ;
      RECT 0.0000 110.2000 69.9200 111.1400 ;
      RECT 0.7350 109.7800 69.1850 110.2000 ;
      RECT 0.0000 108.5000 69.9200 109.7800 ;
      RECT 0.0000 108.0800 69.1850 108.5000 ;
      RECT 0.0000 107.8200 69.9200 108.0800 ;
      RECT 0.7350 107.4000 69.9200 107.8200 ;
      RECT 0.0000 107.1400 69.9200 107.4000 ;
      RECT 0.0000 106.7200 69.1850 107.1400 ;
      RECT 0.0000 105.7800 69.9200 106.7200 ;
      RECT 0.0000 105.4400 69.1850 105.7800 ;
      RECT 0.7350 105.3600 69.1850 105.4400 ;
      RECT 0.7350 105.0200 69.9200 105.3600 ;
      RECT 0.0000 104.0800 69.9200 105.0200 ;
      RECT 0.0000 103.6600 69.1850 104.0800 ;
      RECT 0.0000 103.0600 69.9200 103.6600 ;
      RECT 0.7350 102.7200 69.9200 103.0600 ;
      RECT 0.7350 102.6400 69.1850 102.7200 ;
      RECT 0.0000 102.3000 69.1850 102.6400 ;
      RECT 0.0000 101.3600 69.9200 102.3000 ;
      RECT 0.0000 100.9400 69.1850 101.3600 ;
      RECT 0.0000 100.6800 69.9200 100.9400 ;
      RECT 0.7350 100.2600 69.9200 100.6800 ;
      RECT 0.0000 99.6600 69.9200 100.2600 ;
      RECT 0.0000 99.2400 69.1850 99.6600 ;
      RECT 0.0000 98.6400 69.9200 99.2400 ;
      RECT 0.7350 98.3000 69.9200 98.6400 ;
      RECT 0.7350 98.2200 69.1850 98.3000 ;
      RECT 0.0000 97.8800 69.1850 98.2200 ;
      RECT 0.0000 96.9400 69.9200 97.8800 ;
      RECT 0.0000 96.5200 69.1850 96.9400 ;
      RECT 0.0000 96.2600 69.9200 96.5200 ;
      RECT 0.7350 95.8400 69.9200 96.2600 ;
      RECT 0.0000 95.2400 69.9200 95.8400 ;
      RECT 0.0000 94.8200 69.1850 95.2400 ;
      RECT 0.0000 93.8800 69.9200 94.8200 ;
      RECT 0.7350 93.4600 69.1850 93.8800 ;
      RECT 0.0000 92.5200 69.9200 93.4600 ;
      RECT 0.0000 92.1000 69.1850 92.5200 ;
      RECT 0.0000 91.5000 69.9200 92.1000 ;
      RECT 0.7350 91.0800 69.9200 91.5000 ;
      RECT 0.0000 90.8200 69.9200 91.0800 ;
      RECT 0.0000 90.4000 69.1850 90.8200 ;
      RECT 0.0000 89.4600 69.9200 90.4000 ;
      RECT 0.7350 89.0400 69.1850 89.4600 ;
      RECT 0.0000 88.1000 69.9200 89.0400 ;
      RECT 0.0000 87.6800 69.1850 88.1000 ;
      RECT 0.0000 87.0800 69.9200 87.6800 ;
      RECT 0.7350 86.6600 69.9200 87.0800 ;
      RECT 0.0000 86.4000 69.9200 86.6600 ;
      RECT 0.0000 85.9800 69.1850 86.4000 ;
      RECT 0.0000 85.0400 69.9200 85.9800 ;
      RECT 0.0000 84.7000 69.1850 85.0400 ;
      RECT 0.7350 84.6200 69.1850 84.7000 ;
      RECT 0.7350 84.2800 69.9200 84.6200 ;
      RECT 0.0000 83.6800 69.9200 84.2800 ;
      RECT 0.0000 83.2600 69.1850 83.6800 ;
      RECT 0.0000 82.3200 69.9200 83.2600 ;
      RECT 0.7350 81.9800 69.9200 82.3200 ;
      RECT 0.7350 81.9000 69.1850 81.9800 ;
      RECT 0.0000 81.5600 69.1850 81.9000 ;
      RECT 0.0000 80.6200 69.9200 81.5600 ;
      RECT 0.0000 80.2800 69.1850 80.6200 ;
      RECT 0.7350 80.2000 69.1850 80.2800 ;
      RECT 0.7350 79.8600 69.9200 80.2000 ;
      RECT 0.0000 79.2600 69.9200 79.8600 ;
      RECT 0.0000 78.8400 69.1850 79.2600 ;
      RECT 0.0000 77.9000 69.9200 78.8400 ;
      RECT 0.0000 77.4800 69.1850 77.9000 ;
      RECT 0.0000 76.2000 69.9200 77.4800 ;
      RECT 0.0000 75.7800 69.1850 76.2000 ;
      RECT 0.0000 74.8400 69.9200 75.7800 ;
      RECT 0.0000 74.4200 69.1850 74.8400 ;
      RECT 0.0000 73.4800 69.9200 74.4200 ;
      RECT 0.0000 73.0600 69.1850 73.4800 ;
      RECT 0.0000 71.7800 69.9200 73.0600 ;
      RECT 0.0000 71.3600 69.1850 71.7800 ;
      RECT 0.0000 70.4200 69.9200 71.3600 ;
      RECT 0.0000 70.0000 69.1850 70.4200 ;
      RECT 0.0000 69.0600 69.9200 70.0000 ;
      RECT 0.0000 68.6400 69.1850 69.0600 ;
      RECT 0.0000 67.0200 69.9200 68.6400 ;
      RECT 0.0000 66.6000 69.1850 67.0200 ;
      RECT 0.0000 66.0000 69.9200 66.6000 ;
      RECT 0.0000 65.5800 69.1850 66.0000 ;
      RECT 0.0000 64.6400 69.9200 65.5800 ;
      RECT 0.0000 64.2200 69.1850 64.6400 ;
      RECT 0.0000 62.9400 69.9200 64.2200 ;
      RECT 0.0000 62.5200 69.1850 62.9400 ;
      RECT 0.0000 61.5800 69.9200 62.5200 ;
      RECT 0.0000 61.1600 69.1850 61.5800 ;
      RECT 0.0000 60.2200 69.9200 61.1600 ;
      RECT 0.0000 59.8000 69.1850 60.2200 ;
      RECT 0.0000 58.5200 69.9200 59.8000 ;
      RECT 0.0000 58.1000 69.1850 58.5200 ;
      RECT 0.0000 57.1600 69.9200 58.1000 ;
      RECT 0.0000 56.7400 69.1850 57.1600 ;
      RECT 0.0000 55.4600 69.9200 56.7400 ;
      RECT 0.0000 55.0400 69.1850 55.4600 ;
      RECT 0.0000 54.1000 69.9200 55.0400 ;
      RECT 0.0000 53.6800 69.1850 54.1000 ;
      RECT 0.0000 52.7400 69.9200 53.6800 ;
      RECT 0.0000 52.3200 69.1850 52.7400 ;
      RECT 0.0000 51.3800 69.9200 52.3200 ;
      RECT 0.0000 50.9600 69.1850 51.3800 ;
      RECT 0.0000 49.6800 69.9200 50.9600 ;
      RECT 0.0000 49.2600 69.1850 49.6800 ;
      RECT 0.0000 48.3200 69.9200 49.2600 ;
      RECT 0.0000 47.9000 69.1850 48.3200 ;
      RECT 0.0000 46.9600 69.9200 47.9000 ;
      RECT 0.0000 46.5400 69.1850 46.9600 ;
      RECT 0.0000 45.2600 69.9200 46.5400 ;
      RECT 0.0000 44.8400 69.1850 45.2600 ;
      RECT 0.0000 43.9000 69.9200 44.8400 ;
      RECT 0.0000 43.4800 69.1850 43.9000 ;
      RECT 0.0000 42.5400 69.9200 43.4800 ;
      RECT 0.0000 42.1200 69.1850 42.5400 ;
      RECT 0.0000 40.8400 69.9200 42.1200 ;
      RECT 0.0000 40.4200 69.1850 40.8400 ;
      RECT 0.0000 39.4800 69.9200 40.4200 ;
      RECT 0.0000 39.0600 69.1850 39.4800 ;
      RECT 0.0000 38.1200 69.9200 39.0600 ;
      RECT 0.0000 37.7000 69.1850 38.1200 ;
      RECT 0.0000 36.4200 69.9200 37.7000 ;
      RECT 0.0000 36.0000 69.1850 36.4200 ;
      RECT 0.0000 35.0600 69.9200 36.0000 ;
      RECT 0.0000 34.6400 69.1850 35.0600 ;
      RECT 0.0000 33.7000 69.9200 34.6400 ;
      RECT 0.0000 33.2800 69.1850 33.7000 ;
      RECT 0.0000 32.0000 69.9200 33.2800 ;
      RECT 0.0000 31.5800 69.1850 32.0000 ;
      RECT 0.0000 30.6400 69.9200 31.5800 ;
      RECT 0.0000 30.2200 69.1850 30.6400 ;
      RECT 0.0000 29.2800 69.9200 30.2200 ;
      RECT 0.0000 28.8600 69.1850 29.2800 ;
      RECT 0.0000 27.5800 69.9200 28.8600 ;
      RECT 0.0000 27.1600 69.1850 27.5800 ;
      RECT 0.0000 26.2200 69.9200 27.1600 ;
      RECT 0.0000 25.8000 69.1850 26.2200 ;
      RECT 0.0000 24.8600 69.9200 25.8000 ;
      RECT 0.0000 24.4400 69.1850 24.8600 ;
      RECT 0.0000 23.1600 69.9200 24.4400 ;
      RECT 0.0000 22.7400 69.1850 23.1600 ;
      RECT 0.0000 21.8000 69.9200 22.7400 ;
      RECT 0.0000 21.3800 69.1850 21.8000 ;
      RECT 0.0000 20.4400 69.9200 21.3800 ;
      RECT 0.0000 20.0200 69.1850 20.4400 ;
      RECT 0.0000 18.7400 69.9200 20.0200 ;
      RECT 0.0000 18.3200 69.1850 18.7400 ;
      RECT 0.0000 17.3800 69.9200 18.3200 ;
      RECT 0.0000 16.9600 69.1850 17.3800 ;
      RECT 0.0000 16.0200 69.9200 16.9600 ;
      RECT 0.0000 15.6000 69.1850 16.0200 ;
      RECT 0.0000 14.3200 69.9200 15.6000 ;
      RECT 0.0000 13.9000 69.1850 14.3200 ;
      RECT 0.0000 12.9600 69.9200 13.9000 ;
      RECT 0.0000 12.5400 69.1850 12.9600 ;
      RECT 0.0000 11.6000 69.9200 12.5400 ;
      RECT 0.0000 11.1800 69.1850 11.6000 ;
      RECT 0.0000 10.2400 69.9200 11.1800 ;
      RECT 0.0000 9.8200 69.1850 10.2400 ;
      RECT 0.0000 0.0000 69.9200 9.8200 ;
    LAYER met2 ;
      RECT 0.0000 0.0000 69.9200 219.6400 ;
    LAYER met3 ;
      RECT 0.0000 215.7300 69.9200 219.6400 ;
      RECT 68.6300 214.1300 69.9200 215.7300 ;
      RECT 0.0000 214.1300 1.2900 215.7300 ;
      RECT 0.0000 213.9300 69.9200 214.1300 ;
      RECT 66.8300 212.3300 69.9200 213.9300 ;
      RECT 0.0000 212.3300 3.0900 213.9300 ;
      RECT 0.0000 209.9500 69.9200 212.3300 ;
      RECT 1.1000 209.0500 68.8200 209.9500 ;
      RECT 0.0000 208.9600 69.9200 209.0500 ;
      RECT 66.8300 208.1200 69.9200 208.9600 ;
      RECT 0.0000 208.1200 3.0900 208.9600 ;
      RECT 66.8300 207.8800 68.8200 208.1200 ;
      RECT 4.6900 207.8800 65.2300 208.9600 ;
      RECT 1.1000 207.8800 3.0900 208.1200 ;
      RECT 1.1000 207.2200 68.8200 207.8800 ;
      RECT 0.0000 206.2900 69.9200 207.2200 ;
      RECT 1.1000 206.2400 68.8200 206.2900 ;
      RECT 68.6300 205.3900 68.8200 206.2400 ;
      RECT 1.1000 205.3900 1.2900 206.2400 ;
      RECT 68.6300 205.1600 69.9200 205.3900 ;
      RECT 2.8900 205.1600 67.0300 206.2400 ;
      RECT 0.0000 205.1600 1.2900 205.3900 ;
      RECT 0.0000 204.4600 69.9200 205.1600 ;
      RECT 1.1000 203.5600 68.8200 204.4600 ;
      RECT 0.0000 203.5200 69.9200 203.5600 ;
      RECT 66.8300 202.6300 69.9200 203.5200 ;
      RECT 0.0000 202.6300 3.0900 203.5200 ;
      RECT 66.8300 202.4400 68.8200 202.6300 ;
      RECT 4.6900 202.4400 65.2300 203.5200 ;
      RECT 1.1000 202.4400 3.0900 202.6300 ;
      RECT 1.1000 201.7300 68.8200 202.4400 ;
      RECT 0.0000 200.8000 69.9200 201.7300 ;
      RECT 68.6300 199.9000 68.8200 200.8000 ;
      RECT 1.1000 199.9000 1.2900 200.8000 ;
      RECT 68.6300 199.7200 69.9200 199.9000 ;
      RECT 2.8900 199.7200 67.0300 200.8000 ;
      RECT 0.0000 199.7200 1.2900 199.9000 ;
      RECT 0.0000 198.9700 69.9200 199.7200 ;
      RECT 1.1000 198.0800 68.8200 198.9700 ;
      RECT 66.8300 198.0700 68.8200 198.0800 ;
      RECT 1.1000 198.0700 3.0900 198.0800 ;
      RECT 66.8300 197.1400 69.9200 198.0700 ;
      RECT 0.0000 197.1400 3.0900 198.0700 ;
      RECT 66.8300 197.0000 68.8200 197.1400 ;
      RECT 4.6900 197.0000 65.2300 198.0800 ;
      RECT 1.1000 197.0000 3.0900 197.1400 ;
      RECT 1.1000 196.2400 68.8200 197.0000 ;
      RECT 0.0000 195.9200 69.9200 196.2400 ;
      RECT 1.1000 195.3600 68.8200 195.9200 ;
      RECT 68.6300 195.0200 68.8200 195.3600 ;
      RECT 1.1000 195.0200 1.2900 195.3600 ;
      RECT 68.6300 194.2800 69.9200 195.0200 ;
      RECT 2.8900 194.2800 67.0300 195.3600 ;
      RECT 0.0000 194.2800 1.2900 195.0200 ;
      RECT 0.0000 194.0900 69.9200 194.2800 ;
      RECT 1.1000 193.1900 68.8200 194.0900 ;
      RECT 0.0000 192.6400 69.9200 193.1900 ;
      RECT 66.8300 192.2600 69.9200 192.6400 ;
      RECT 0.0000 192.2600 3.0900 192.6400 ;
      RECT 66.8300 191.5600 68.8200 192.2600 ;
      RECT 4.6900 191.5600 65.2300 192.6400 ;
      RECT 1.1000 191.5600 3.0900 192.2600 ;
      RECT 1.1000 191.3600 68.8200 191.5600 ;
      RECT 0.0000 190.4300 69.9200 191.3600 ;
      RECT 1.1000 189.9200 68.8200 190.4300 ;
      RECT 68.6300 189.5300 68.8200 189.9200 ;
      RECT 1.1000 189.5300 1.2900 189.9200 ;
      RECT 68.6300 188.8400 69.9200 189.5300 ;
      RECT 2.8900 188.8400 67.0300 189.9200 ;
      RECT 0.0000 188.8400 1.2900 189.5300 ;
      RECT 0.0000 188.6000 69.9200 188.8400 ;
      RECT 1.1000 187.7000 68.8200 188.6000 ;
      RECT 0.0000 187.2000 69.9200 187.7000 ;
      RECT 66.8300 186.7700 69.9200 187.2000 ;
      RECT 0.0000 186.7700 3.0900 187.2000 ;
      RECT 66.8300 186.1200 68.8200 186.7700 ;
      RECT 4.6900 186.1200 65.2300 187.2000 ;
      RECT 1.1000 186.1200 3.0900 186.7700 ;
      RECT 1.1000 185.8700 68.8200 186.1200 ;
      RECT 0.0000 184.9400 69.9200 185.8700 ;
      RECT 1.1000 184.4800 68.8200 184.9400 ;
      RECT 68.6300 184.0400 68.8200 184.4800 ;
      RECT 1.1000 184.0400 1.2900 184.4800 ;
      RECT 68.6300 183.4000 69.9200 184.0400 ;
      RECT 2.8900 183.4000 67.0300 184.4800 ;
      RECT 0.0000 183.4000 1.2900 184.0400 ;
      RECT 0.0000 183.1100 69.9200 183.4000 ;
      RECT 1.1000 182.2100 68.8200 183.1100 ;
      RECT 0.0000 181.8900 69.9200 182.2100 ;
      RECT 1.1000 181.7600 68.8200 181.8900 ;
      RECT 66.8300 180.9900 68.8200 181.7600 ;
      RECT 1.1000 180.9900 3.0900 181.7600 ;
      RECT 66.8300 180.6800 69.9200 180.9900 ;
      RECT 4.6900 180.6800 65.2300 181.7600 ;
      RECT 0.0000 180.6800 3.0900 180.9900 ;
      RECT 0.0000 180.0600 69.9200 180.6800 ;
      RECT 1.1000 179.1600 68.8200 180.0600 ;
      RECT 0.0000 179.0400 69.9200 179.1600 ;
      RECT 68.6300 178.2300 69.9200 179.0400 ;
      RECT 0.0000 178.2300 1.2900 179.0400 ;
      RECT 68.6300 177.9600 68.8200 178.2300 ;
      RECT 2.8900 177.9600 67.0300 179.0400 ;
      RECT 1.1000 177.9600 1.2900 178.2300 ;
      RECT 1.1000 177.3300 68.8200 177.9600 ;
      RECT 0.0000 176.4000 69.9200 177.3300 ;
      RECT 1.1000 176.3200 68.8200 176.4000 ;
      RECT 66.8300 175.5000 68.8200 176.3200 ;
      RECT 1.1000 175.5000 3.0900 176.3200 ;
      RECT 66.8300 175.2400 69.9200 175.5000 ;
      RECT 4.6900 175.2400 65.2300 176.3200 ;
      RECT 0.0000 175.2400 3.0900 175.5000 ;
      RECT 0.0000 174.5700 69.9200 175.2400 ;
      RECT 1.1000 173.6700 68.8200 174.5700 ;
      RECT 0.0000 173.6000 69.9200 173.6700 ;
      RECT 68.6300 172.7400 69.9200 173.6000 ;
      RECT 0.0000 172.7400 1.2900 173.6000 ;
      RECT 68.6300 172.5200 68.8200 172.7400 ;
      RECT 2.8900 172.5200 67.0300 173.6000 ;
      RECT 1.1000 172.5200 1.2900 172.7400 ;
      RECT 1.1000 171.8400 68.8200 172.5200 ;
      RECT 0.0000 170.9100 69.9200 171.8400 ;
      RECT 1.1000 170.8800 68.8200 170.9100 ;
      RECT 66.8300 170.0100 68.8200 170.8800 ;
      RECT 1.1000 170.0100 3.0900 170.8800 ;
      RECT 66.8300 169.8000 69.9200 170.0100 ;
      RECT 4.6900 169.8000 65.2300 170.8800 ;
      RECT 0.0000 169.8000 3.0900 170.0100 ;
      RECT 0.0000 169.0800 69.9200 169.8000 ;
      RECT 1.1000 168.1800 68.8200 169.0800 ;
      RECT 0.0000 168.1600 69.9200 168.1800 ;
      RECT 68.6300 167.8600 69.9200 168.1600 ;
      RECT 0.0000 167.8600 1.2900 168.1600 ;
      RECT 68.6300 167.0800 68.8200 167.8600 ;
      RECT 2.8900 167.0800 67.0300 168.1600 ;
      RECT 1.1000 167.0800 1.2900 167.8600 ;
      RECT 1.1000 166.9600 68.8200 167.0800 ;
      RECT 0.0000 166.0300 69.9200 166.9600 ;
      RECT 1.1000 165.4400 68.8200 166.0300 ;
      RECT 66.8300 165.1300 68.8200 165.4400 ;
      RECT 1.1000 165.1300 3.0900 165.4400 ;
      RECT 66.8300 164.3600 69.9200 165.1300 ;
      RECT 4.6900 164.3600 65.2300 165.4400 ;
      RECT 0.0000 164.3600 3.0900 165.1300 ;
      RECT 0.0000 164.2000 69.9200 164.3600 ;
      RECT 1.1000 163.3000 68.8200 164.2000 ;
      RECT 0.0000 162.7200 69.9200 163.3000 ;
      RECT 0.0000 162.3700 1.2900 162.7200 ;
      RECT 68.6300 161.7600 69.9200 162.7200 ;
      RECT 68.6300 161.6400 68.8200 161.7600 ;
      RECT 2.8900 161.6400 67.0300 162.7200 ;
      RECT 1.1000 161.6400 1.2900 162.3700 ;
      RECT 1.1000 161.4700 68.8200 161.6400 ;
      RECT 0.0000 160.8600 68.8200 161.4700 ;
      RECT 0.0000 160.5400 69.9200 160.8600 ;
      RECT 1.1000 160.0000 68.8200 160.5400 ;
      RECT 66.8300 159.6400 68.8200 160.0000 ;
      RECT 1.1000 159.6400 3.0900 160.0000 ;
      RECT 66.8300 158.9200 69.9200 159.6400 ;
      RECT 4.6900 158.9200 65.2300 160.0000 ;
      RECT 0.0000 158.9200 3.0900 159.6400 ;
      RECT 0.0000 158.7100 69.9200 158.9200 ;
      RECT 1.1000 157.8100 68.8200 158.7100 ;
      RECT 0.0000 157.2800 69.9200 157.8100 ;
      RECT 68.6300 156.8800 69.9200 157.2800 ;
      RECT 0.0000 156.8800 1.2900 157.2800 ;
      RECT 68.6300 156.2000 68.8200 156.8800 ;
      RECT 2.8900 156.2000 67.0300 157.2800 ;
      RECT 1.1000 156.2000 1.2900 156.8800 ;
      RECT 1.1000 155.9800 68.8200 156.2000 ;
      RECT 0.0000 155.6600 69.9200 155.9800 ;
      RECT 1.1000 154.7600 68.8200 155.6600 ;
      RECT 0.0000 154.5600 69.9200 154.7600 ;
      RECT 66.8300 153.4800 69.9200 154.5600 ;
      RECT 4.6900 153.4800 65.2300 154.5600 ;
      RECT 0.0000 153.4800 3.0900 154.5600 ;
      RECT 0.0000 151.8400 69.9200 153.4800 ;
      RECT 68.6300 150.7600 69.9200 151.8400 ;
      RECT 2.8900 150.7600 67.0300 151.8400 ;
      RECT 0.0000 150.7600 1.2900 151.8400 ;
      RECT 0.0000 149.1200 69.9200 150.7600 ;
      RECT 66.8300 148.0400 69.9200 149.1200 ;
      RECT 4.6900 148.0400 65.2300 149.1200 ;
      RECT 0.0000 148.0400 3.0900 149.1200 ;
      RECT 0.0000 146.4000 69.9200 148.0400 ;
      RECT 68.6300 145.3200 69.9200 146.4000 ;
      RECT 2.8900 145.3200 67.0300 146.4000 ;
      RECT 0.0000 145.3200 1.2900 146.4000 ;
      RECT 0.0000 143.6800 69.9200 145.3200 ;
      RECT 66.8300 142.6000 69.9200 143.6800 ;
      RECT 4.6900 142.6000 65.2300 143.6800 ;
      RECT 0.0000 142.6000 3.0900 143.6800 ;
      RECT 0.0000 140.9600 69.9200 142.6000 ;
      RECT 68.6300 139.8800 69.9200 140.9600 ;
      RECT 2.8900 139.8800 67.0300 140.9600 ;
      RECT 0.0000 139.8800 1.2900 140.9600 ;
      RECT 0.0000 138.2400 69.9200 139.8800 ;
      RECT 66.8300 137.1600 69.9200 138.2400 ;
      RECT 4.6900 137.1600 65.2300 138.2400 ;
      RECT 0.0000 137.1600 3.0900 138.2400 ;
      RECT 0.0000 135.5200 69.9200 137.1600 ;
      RECT 68.6300 134.4400 69.9200 135.5200 ;
      RECT 2.8900 134.4400 67.0300 135.5200 ;
      RECT 0.0000 134.4400 1.2900 135.5200 ;
      RECT 0.0000 132.8000 69.9200 134.4400 ;
      RECT 66.8300 131.7200 69.9200 132.8000 ;
      RECT 4.6900 131.7200 65.2300 132.8000 ;
      RECT 0.0000 131.7200 3.0900 132.8000 ;
      RECT 0.0000 130.0800 69.9200 131.7200 ;
      RECT 68.6300 129.0000 69.9200 130.0800 ;
      RECT 2.8900 129.0000 67.0300 130.0800 ;
      RECT 0.0000 129.0000 1.2900 130.0800 ;
      RECT 0.0000 127.3600 69.9200 129.0000 ;
      RECT 66.8300 126.2800 69.9200 127.3600 ;
      RECT 4.6900 126.2800 65.2300 127.3600 ;
      RECT 0.0000 126.2800 3.0900 127.3600 ;
      RECT 0.0000 124.6400 69.9200 126.2800 ;
      RECT 68.6300 123.5600 69.9200 124.6400 ;
      RECT 2.8900 123.5600 67.0300 124.6400 ;
      RECT 0.0000 123.5600 1.2900 124.6400 ;
      RECT 0.0000 121.9200 69.9200 123.5600 ;
      RECT 66.8300 120.8400 69.9200 121.9200 ;
      RECT 4.6900 120.8400 65.2300 121.9200 ;
      RECT 0.0000 120.8400 3.0900 121.9200 ;
      RECT 0.0000 119.2000 69.9200 120.8400 ;
      RECT 68.6300 118.1200 69.9200 119.2000 ;
      RECT 2.8900 118.1200 67.0300 119.2000 ;
      RECT 0.0000 118.1200 1.2900 119.2000 ;
      RECT 0.0000 116.4800 69.9200 118.1200 ;
      RECT 66.8300 115.4000 69.9200 116.4800 ;
      RECT 4.6900 115.4000 65.2300 116.4800 ;
      RECT 0.0000 115.4000 3.0900 116.4800 ;
      RECT 0.0000 113.7600 69.9200 115.4000 ;
      RECT 68.6300 112.6800 69.9200 113.7600 ;
      RECT 2.8900 112.6800 67.0300 113.7600 ;
      RECT 0.0000 112.6800 1.2900 113.7600 ;
      RECT 0.0000 111.0400 69.9200 112.6800 ;
      RECT 66.8300 109.9600 69.9200 111.0400 ;
      RECT 4.6900 109.9600 65.2300 111.0400 ;
      RECT 0.0000 109.9600 3.0900 111.0400 ;
      RECT 0.0000 108.3200 69.9200 109.9600 ;
      RECT 68.6300 107.2400 69.9200 108.3200 ;
      RECT 2.8900 107.2400 67.0300 108.3200 ;
      RECT 0.0000 107.2400 1.2900 108.3200 ;
      RECT 0.0000 105.6000 69.9200 107.2400 ;
      RECT 66.8300 104.5200 69.9200 105.6000 ;
      RECT 4.6900 104.5200 65.2300 105.6000 ;
      RECT 0.0000 104.5200 3.0900 105.6000 ;
      RECT 0.0000 102.8800 69.9200 104.5200 ;
      RECT 68.6300 101.8000 69.9200 102.8800 ;
      RECT 2.8900 101.8000 67.0300 102.8800 ;
      RECT 0.0000 101.8000 1.2900 102.8800 ;
      RECT 0.0000 100.1600 69.9200 101.8000 ;
      RECT 66.8300 99.0800 69.9200 100.1600 ;
      RECT 4.6900 99.0800 65.2300 100.1600 ;
      RECT 0.0000 99.0800 3.0900 100.1600 ;
      RECT 0.0000 97.4400 69.9200 99.0800 ;
      RECT 68.6300 96.3600 69.9200 97.4400 ;
      RECT 2.8900 96.3600 67.0300 97.4400 ;
      RECT 0.0000 96.3600 1.2900 97.4400 ;
      RECT 0.0000 94.7200 69.9200 96.3600 ;
      RECT 66.8300 93.6400 69.9200 94.7200 ;
      RECT 4.6900 93.6400 65.2300 94.7200 ;
      RECT 0.0000 93.6400 3.0900 94.7200 ;
      RECT 0.0000 92.0000 69.9200 93.6400 ;
      RECT 68.6300 90.9200 69.9200 92.0000 ;
      RECT 2.8900 90.9200 67.0300 92.0000 ;
      RECT 0.0000 90.9200 1.2900 92.0000 ;
      RECT 0.0000 89.2800 69.9200 90.9200 ;
      RECT 66.8300 88.2000 69.9200 89.2800 ;
      RECT 4.6900 88.2000 65.2300 89.2800 ;
      RECT 0.0000 88.2000 3.0900 89.2800 ;
      RECT 0.0000 86.5600 69.9200 88.2000 ;
      RECT 68.6300 85.4800 69.9200 86.5600 ;
      RECT 2.8900 85.4800 67.0300 86.5600 ;
      RECT 0.0000 85.4800 1.2900 86.5600 ;
      RECT 0.0000 83.8400 69.9200 85.4800 ;
      RECT 66.8300 82.7600 69.9200 83.8400 ;
      RECT 4.6900 82.7600 65.2300 83.8400 ;
      RECT 0.0000 82.7600 3.0900 83.8400 ;
      RECT 0.0000 81.1200 69.9200 82.7600 ;
      RECT 68.6300 80.0400 69.9200 81.1200 ;
      RECT 2.8900 80.0400 67.0300 81.1200 ;
      RECT 0.0000 80.0400 1.2900 81.1200 ;
      RECT 0.0000 78.4000 69.9200 80.0400 ;
      RECT 66.8300 77.3200 69.9200 78.4000 ;
      RECT 4.6900 77.3200 65.2300 78.4000 ;
      RECT 0.0000 77.3200 3.0900 78.4000 ;
      RECT 0.0000 75.6800 69.9200 77.3200 ;
      RECT 68.6300 74.6000 69.9200 75.6800 ;
      RECT 2.8900 74.6000 67.0300 75.6800 ;
      RECT 0.0000 74.6000 1.2900 75.6800 ;
      RECT 0.0000 72.9600 69.9200 74.6000 ;
      RECT 66.8300 71.8800 69.9200 72.9600 ;
      RECT 4.6900 71.8800 65.2300 72.9600 ;
      RECT 0.0000 71.8800 3.0900 72.9600 ;
      RECT 0.0000 70.2400 69.9200 71.8800 ;
      RECT 68.6300 69.1600 69.9200 70.2400 ;
      RECT 2.8900 69.1600 67.0300 70.2400 ;
      RECT 0.0000 69.1600 1.2900 70.2400 ;
      RECT 0.0000 67.5200 69.9200 69.1600 ;
      RECT 66.8300 66.4400 69.9200 67.5200 ;
      RECT 4.6900 66.4400 65.2300 67.5200 ;
      RECT 0.0000 66.4400 3.0900 67.5200 ;
      RECT 0.0000 64.8000 69.9200 66.4400 ;
      RECT 68.6300 63.7200 69.9200 64.8000 ;
      RECT 2.8900 63.7200 67.0300 64.8000 ;
      RECT 0.0000 63.7200 1.2900 64.8000 ;
      RECT 0.0000 62.0800 69.9200 63.7200 ;
      RECT 66.8300 61.0000 69.9200 62.0800 ;
      RECT 4.6900 61.0000 65.2300 62.0800 ;
      RECT 0.0000 61.0000 3.0900 62.0800 ;
      RECT 0.0000 59.3600 69.9200 61.0000 ;
      RECT 68.6300 58.2800 69.9200 59.3600 ;
      RECT 2.8900 58.2800 67.0300 59.3600 ;
      RECT 0.0000 58.2800 1.2900 59.3600 ;
      RECT 0.0000 56.6400 69.9200 58.2800 ;
      RECT 66.8300 55.5600 69.9200 56.6400 ;
      RECT 4.6900 55.5600 65.2300 56.6400 ;
      RECT 0.0000 55.5600 3.0900 56.6400 ;
      RECT 0.0000 53.9200 69.9200 55.5600 ;
      RECT 68.6300 52.8400 69.9200 53.9200 ;
      RECT 2.8900 52.8400 67.0300 53.9200 ;
      RECT 0.0000 52.8400 1.2900 53.9200 ;
      RECT 0.0000 51.2000 69.9200 52.8400 ;
      RECT 66.8300 50.1200 69.9200 51.2000 ;
      RECT 4.6900 50.1200 65.2300 51.2000 ;
      RECT 0.0000 50.1200 3.0900 51.2000 ;
      RECT 0.0000 48.4800 69.9200 50.1200 ;
      RECT 68.6300 47.4000 69.9200 48.4800 ;
      RECT 2.8900 47.4000 67.0300 48.4800 ;
      RECT 0.0000 47.4000 1.2900 48.4800 ;
      RECT 0.0000 45.7600 69.9200 47.4000 ;
      RECT 66.8300 44.6800 69.9200 45.7600 ;
      RECT 4.6900 44.6800 65.2300 45.7600 ;
      RECT 0.0000 44.6800 3.0900 45.7600 ;
      RECT 0.0000 43.0400 69.9200 44.6800 ;
      RECT 68.6300 41.9600 69.9200 43.0400 ;
      RECT 2.8900 41.9600 67.0300 43.0400 ;
      RECT 0.0000 41.9600 1.2900 43.0400 ;
      RECT 0.0000 40.3200 69.9200 41.9600 ;
      RECT 66.8300 39.2400 69.9200 40.3200 ;
      RECT 4.6900 39.2400 65.2300 40.3200 ;
      RECT 0.0000 39.2400 3.0900 40.3200 ;
      RECT 0.0000 37.6000 69.9200 39.2400 ;
      RECT 68.6300 36.5200 69.9200 37.6000 ;
      RECT 2.8900 36.5200 67.0300 37.6000 ;
      RECT 0.0000 36.5200 1.2900 37.6000 ;
      RECT 0.0000 34.8800 69.9200 36.5200 ;
      RECT 66.8300 33.8000 69.9200 34.8800 ;
      RECT 4.6900 33.8000 65.2300 34.8800 ;
      RECT 0.0000 33.8000 3.0900 34.8800 ;
      RECT 0.0000 32.1600 69.9200 33.8000 ;
      RECT 68.6300 31.0800 69.9200 32.1600 ;
      RECT 2.8900 31.0800 67.0300 32.1600 ;
      RECT 0.0000 31.0800 1.2900 32.1600 ;
      RECT 0.0000 29.4400 69.9200 31.0800 ;
      RECT 66.8300 28.3600 69.9200 29.4400 ;
      RECT 4.6900 28.3600 65.2300 29.4400 ;
      RECT 0.0000 28.3600 3.0900 29.4400 ;
      RECT 0.0000 26.7200 69.9200 28.3600 ;
      RECT 68.6300 25.6400 69.9200 26.7200 ;
      RECT 2.8900 25.6400 67.0300 26.7200 ;
      RECT 0.0000 25.6400 1.2900 26.7200 ;
      RECT 0.0000 24.0000 69.9200 25.6400 ;
      RECT 66.8300 22.9200 69.9200 24.0000 ;
      RECT 4.6900 22.9200 65.2300 24.0000 ;
      RECT 0.0000 22.9200 3.0900 24.0000 ;
      RECT 0.0000 21.2800 69.9200 22.9200 ;
      RECT 68.6300 20.2000 69.9200 21.2800 ;
      RECT 2.8900 20.2000 67.0300 21.2800 ;
      RECT 0.0000 20.2000 1.2900 21.2800 ;
      RECT 0.0000 18.5600 69.9200 20.2000 ;
      RECT 66.8300 17.4800 69.9200 18.5600 ;
      RECT 4.6900 17.4800 65.2300 18.5600 ;
      RECT 0.0000 17.4800 3.0900 18.5600 ;
      RECT 0.0000 15.8400 69.9200 17.4800 ;
      RECT 68.6300 14.7600 69.9200 15.8400 ;
      RECT 2.8900 14.7600 67.0300 15.8400 ;
      RECT 0.0000 14.7600 1.2900 15.8400 ;
      RECT 0.0000 13.1200 69.9200 14.7600 ;
      RECT 66.8300 12.0400 69.9200 13.1200 ;
      RECT 4.6900 12.0400 65.2300 13.1200 ;
      RECT 0.0000 12.0400 3.0900 13.1200 ;
      RECT 0.0000 10.4000 69.9200 12.0400 ;
      RECT 68.6300 9.3200 69.9200 10.4000 ;
      RECT 2.8900 9.3200 67.0300 10.4000 ;
      RECT 0.0000 9.3200 1.2900 10.4000 ;
      RECT 0.0000 6.6300 69.9200 9.3200 ;
      RECT 66.8300 5.0300 69.9200 6.6300 ;
      RECT 0.0000 5.0300 3.0900 6.6300 ;
      RECT 0.0000 4.8300 69.9200 5.0300 ;
      RECT 68.6300 3.2300 69.9200 4.8300 ;
      RECT 0.0000 3.2300 1.2900 4.8300 ;
      RECT 0.0000 0.0000 69.9200 3.2300 ;
    LAYER met4 ;
      RECT 0.0000 215.7300 69.9200 219.6400 ;
      RECT 2.8900 213.9300 67.0300 215.7300 ;
      RECT 66.8300 5.0300 67.0300 213.9300 ;
      RECT 4.6900 5.0300 65.2300 213.9300 ;
      RECT 2.8900 5.0300 3.0900 213.9300 ;
      RECT 68.6300 3.2300 69.9200 215.7300 ;
      RECT 2.8900 3.2300 67.0300 5.0300 ;
      RECT 0.0000 3.2300 1.2900 215.7300 ;
      RECT 0.0000 0.0000 69.9200 3.2300 ;
  END
END W_IO

END LIBRARY
