magic
tech sky130A
timestamp 1707688321
<< pwell >>
rect -13 -13 1924 54
<< psubdiff >>
rect 0 29 1911 41
rect 0 12 12 29
rect 29 12 46 29
rect 63 12 80 29
rect 97 12 114 29
rect 131 12 148 29
rect 165 12 182 29
rect 199 12 216 29
rect 233 12 250 29
rect 267 12 284 29
rect 301 12 318 29
rect 335 12 352 29
rect 369 12 386 29
rect 403 12 420 29
rect 437 12 454 29
rect 471 12 488 29
rect 505 12 522 29
rect 539 12 556 29
rect 573 12 590 29
rect 607 12 624 29
rect 641 12 658 29
rect 675 12 692 29
rect 709 12 726 29
rect 743 12 760 29
rect 777 12 794 29
rect 811 12 828 29
rect 845 12 862 29
rect 879 12 896 29
rect 913 12 930 29
rect 947 12 964 29
rect 981 12 998 29
rect 1015 12 1032 29
rect 1049 12 1066 29
rect 1083 12 1100 29
rect 1117 12 1134 29
rect 1151 12 1168 29
rect 1185 12 1202 29
rect 1219 12 1236 29
rect 1253 12 1270 29
rect 1287 12 1304 29
rect 1321 12 1338 29
rect 1355 12 1372 29
rect 1389 12 1406 29
rect 1423 12 1440 29
rect 1457 12 1474 29
rect 1491 12 1508 29
rect 1525 12 1542 29
rect 1559 12 1576 29
rect 1593 12 1610 29
rect 1627 12 1644 29
rect 1661 12 1678 29
rect 1695 12 1712 29
rect 1729 12 1746 29
rect 1763 12 1780 29
rect 1797 12 1814 29
rect 1831 12 1848 29
rect 1865 12 1882 29
rect 1899 12 1911 29
rect 0 0 1911 12
<< psubdiffcont >>
rect 12 12 29 29
rect 46 12 63 29
rect 80 12 97 29
rect 114 12 131 29
rect 148 12 165 29
rect 182 12 199 29
rect 216 12 233 29
rect 250 12 267 29
rect 284 12 301 29
rect 318 12 335 29
rect 352 12 369 29
rect 386 12 403 29
rect 420 12 437 29
rect 454 12 471 29
rect 488 12 505 29
rect 522 12 539 29
rect 556 12 573 29
rect 590 12 607 29
rect 624 12 641 29
rect 658 12 675 29
rect 692 12 709 29
rect 726 12 743 29
rect 760 12 777 29
rect 794 12 811 29
rect 828 12 845 29
rect 862 12 879 29
rect 896 12 913 29
rect 930 12 947 29
rect 964 12 981 29
rect 998 12 1015 29
rect 1032 12 1049 29
rect 1066 12 1083 29
rect 1100 12 1117 29
rect 1134 12 1151 29
rect 1168 12 1185 29
rect 1202 12 1219 29
rect 1236 12 1253 29
rect 1270 12 1287 29
rect 1304 12 1321 29
rect 1338 12 1355 29
rect 1372 12 1389 29
rect 1406 12 1423 29
rect 1440 12 1457 29
rect 1474 12 1491 29
rect 1508 12 1525 29
rect 1542 12 1559 29
rect 1576 12 1593 29
rect 1610 12 1627 29
rect 1644 12 1661 29
rect 1678 12 1695 29
rect 1712 12 1729 29
rect 1746 12 1763 29
rect 1780 12 1797 29
rect 1814 12 1831 29
rect 1848 12 1865 29
rect 1882 12 1899 29
<< locali >>
rect 12 29 1899 37
rect 29 12 46 29
rect 63 12 80 29
rect 97 12 114 29
rect 131 12 148 29
rect 165 12 182 29
rect 199 12 216 29
rect 233 12 250 29
rect 267 12 284 29
rect 301 12 318 29
rect 335 12 352 29
rect 369 12 386 29
rect 403 12 420 29
rect 437 12 454 29
rect 471 12 488 29
rect 505 12 522 29
rect 539 12 556 29
rect 573 12 590 29
rect 607 12 624 29
rect 641 12 658 29
rect 675 12 692 29
rect 709 12 726 29
rect 743 12 760 29
rect 777 12 794 29
rect 811 12 828 29
rect 845 12 862 29
rect 879 12 896 29
rect 913 12 930 29
rect 947 12 964 29
rect 981 12 998 29
rect 1015 12 1032 29
rect 1049 12 1066 29
rect 1083 12 1100 29
rect 1117 12 1134 29
rect 1151 12 1168 29
rect 1185 12 1202 29
rect 1219 12 1236 29
rect 1253 12 1270 29
rect 1287 12 1304 29
rect 1321 12 1338 29
rect 1355 12 1372 29
rect 1389 12 1406 29
rect 1423 12 1440 29
rect 1457 12 1474 29
rect 1491 12 1508 29
rect 1525 12 1542 29
rect 1559 12 1576 29
rect 1593 12 1610 29
rect 1627 12 1644 29
rect 1661 12 1678 29
rect 1695 12 1712 29
rect 1729 12 1746 29
rect 1763 12 1780 29
rect 1797 12 1814 29
rect 1831 12 1848 29
rect 1865 12 1882 29
rect 12 4 1899 12
<< properties >>
string GDS_END 42946140
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42942360
<< end >>
