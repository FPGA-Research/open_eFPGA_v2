magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 145 157 415 203
rect 48 21 415 157
rect 48 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 126 47 156 131
rect 223 47 253 177
rect 307 47 337 177
<< scpmoshvt >>
rect 127 297 157 381
rect 235 297 265 497
rect 307 297 337 497
<< ndiff >>
rect 171 163 223 177
rect 171 131 179 163
rect 74 108 126 131
rect 74 74 82 108
rect 116 74 126 108
rect 74 47 126 74
rect 156 129 179 131
rect 213 129 223 163
rect 156 95 223 129
rect 156 61 179 95
rect 213 61 223 95
rect 156 47 223 61
rect 253 163 307 177
rect 253 129 263 163
rect 297 129 307 163
rect 253 95 307 129
rect 253 61 263 95
rect 297 61 307 95
rect 253 47 307 61
rect 337 95 389 177
rect 337 61 347 95
rect 381 61 389 95
rect 337 47 389 61
<< pdiff >>
rect 183 485 235 497
rect 183 451 191 485
rect 225 451 235 485
rect 183 417 235 451
rect 183 383 191 417
rect 225 383 235 417
rect 183 381 235 383
rect 75 363 127 381
rect 75 329 83 363
rect 117 329 127 363
rect 75 297 127 329
rect 157 297 235 381
rect 265 297 307 497
rect 337 485 389 497
rect 337 451 347 485
rect 381 451 389 485
rect 337 417 389 451
rect 337 383 347 417
rect 381 383 389 417
rect 337 297 389 383
<< ndiffc >>
rect 82 74 116 108
rect 179 129 213 163
rect 179 61 213 95
rect 263 129 297 163
rect 263 61 297 95
rect 347 61 381 95
<< pdiffc >>
rect 191 451 225 485
rect 191 383 225 417
rect 83 329 117 363
rect 347 451 381 485
rect 347 383 381 417
<< poly >>
rect 235 497 265 523
rect 307 497 337 523
rect 127 381 157 407
rect 127 265 157 297
rect 235 265 265 297
rect 21 249 157 265
rect 21 215 31 249
rect 65 215 157 249
rect 21 199 157 215
rect 199 249 265 265
rect 199 215 215 249
rect 249 215 265 249
rect 199 199 265 215
rect 307 265 337 297
rect 307 249 373 265
rect 307 215 323 249
rect 357 215 373 249
rect 307 199 373 215
rect 126 131 156 199
rect 223 177 253 199
rect 307 177 337 199
rect 126 21 156 47
rect 223 21 253 47
rect 307 21 337 47
<< polycont >>
rect 31 215 65 249
rect 215 215 249 249
rect 323 215 357 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 175 485 241 527
rect 175 451 191 485
rect 225 451 241 485
rect 175 417 241 451
rect 175 383 191 417
rect 225 383 241 417
rect 83 363 135 381
rect 175 371 241 383
rect 331 485 443 493
rect 331 451 347 485
rect 381 451 443 485
rect 331 417 443 451
rect 331 383 347 417
rect 381 383 443 417
rect 331 370 443 383
rect 117 336 135 363
rect 117 329 341 336
rect 83 302 341 329
rect 20 249 65 265
rect 20 215 31 249
rect 20 145 65 215
rect 99 109 135 302
rect 192 249 265 265
rect 192 215 215 249
rect 249 215 265 249
rect 307 249 341 302
rect 307 215 323 249
rect 357 215 373 249
rect 192 213 265 215
rect 407 179 443 370
rect 66 108 135 109
rect 66 74 82 108
rect 116 74 135 108
rect 171 163 213 179
rect 171 129 179 163
rect 171 95 213 129
rect 171 61 179 95
rect 171 17 213 61
rect 247 163 443 179
rect 247 129 263 163
rect 297 145 443 163
rect 297 129 313 145
rect 247 95 313 129
rect 247 61 263 95
rect 297 61 313 95
rect 247 51 313 61
rect 347 95 424 111
rect 381 61 424 95
rect 347 17 424 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 400 180 0 0 B_N
port 2 nsew signal input
flabel locali s 397 425 431 459 0 FreeSans 400 180 0 0 Y
port 7 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 400 180 0 0 A
port 1 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nor2b_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1980508
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1976254
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
