magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 378
rect 93 0 96 378
<< via1 >>
rect 3 0 93 378
<< metal2 >>
rect 0 0 3 378
rect 93 0 96 378
<< properties >>
string GDS_END 87632188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87629752
<< end >>
