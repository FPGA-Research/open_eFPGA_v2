magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 1719 266
<< mvpmos >>
rect 0 0 1600 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 1600 182 1653 200
rect 1600 148 1611 182
rect 1645 148 1653 182
rect 1600 114 1653 148
rect 1600 80 1611 114
rect 1645 80 1653 114
rect 1600 46 1653 80
rect 1600 12 1611 46
rect 1645 12 1653 46
rect 1600 0 1653 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 1611 148 1645 182
rect 1611 80 1645 114
rect 1611 12 1645 46
<< poly >>
rect 0 200 1600 232
rect 0 -32 1600 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 1611 182 1645 198
rect 1611 114 1645 148
rect 1611 46 1645 80
rect 1611 -4 1645 12
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_1
timestamp 1707688321
transform 1 0 1600 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 1628 97 1628 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6680826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6679812
<< end >>
