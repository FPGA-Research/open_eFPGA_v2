magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 531 666
<< mvpmos >>
rect 0 0 100 600
rect 156 0 256 600
rect 312 0 412 600
<< mvpdiff >>
rect -50 0 0 600
rect 412 0 462 600
<< poly >>
rect 0 600 100 626
rect 0 -26 100 0
rect 156 600 256 626
rect 156 -26 256 0
rect 312 600 412 626
rect 312 -26 412 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
rect 267 -4 301 538
rect 423 -4 457 538
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_0
timestamp 1707688321
transform 1 0 256 0 1 0
box -36 -36 92 636
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_1
timestamp 1707688321
transform 1 0 100 0 1 0
box -36 -36 92 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_1
timestamp 1707688321
transform 1 0 412 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 440 267 440 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87980864
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87978846
<< end >>
