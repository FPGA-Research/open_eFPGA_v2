magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 665 136 674
rect 56 609 80 665
rect 0 465 136 609
rect 56 409 80 465
rect 0 265 136 409
rect 56 209 80 265
rect 0 65 136 209
rect 56 9 80 65
rect 0 0 136 9
<< via2 >>
rect 0 609 56 665
rect 80 609 136 665
rect 0 409 56 465
rect 80 409 136 465
rect 0 209 56 265
rect 80 209 136 265
rect 0 9 56 65
rect 80 9 136 65
<< metal3 >>
rect -5 665 141 670
rect -5 609 0 665
rect 56 609 80 665
rect 136 609 141 665
rect -5 465 141 609
rect -5 409 0 465
rect 56 409 80 465
rect 136 409 141 465
rect -5 265 141 409
rect -5 209 0 265
rect 56 209 80 265
rect 136 209 141 265
rect -5 65 141 209
rect -5 9 0 65
rect 56 9 80 65
rect 136 9 141 65
rect -5 4 141 9
<< properties >>
string GDS_END 78395850
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78395206
<< end >>
