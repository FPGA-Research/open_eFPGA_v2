magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 80 80 3376 39920
<< nwell >>
rect 0 39714 3456 40000
rect 0 286 286 39714
rect 3170 286 3456 39714
rect 0 0 3456 286
<< pwell >>
rect 347 39105 3109 39217
rect 347 606 459 39105
rect 2997 606 3109 39105
rect 347 494 3109 606
<< mvpsubdiff >>
rect 373 39178 3083 39191
rect 373 39144 465 39178
rect 499 39144 533 39178
rect 567 39144 601 39178
rect 635 39144 669 39178
rect 703 39144 737 39178
rect 771 39144 805 39178
rect 839 39144 873 39178
rect 907 39144 941 39178
rect 975 39144 1009 39178
rect 1043 39144 1077 39178
rect 1111 39144 1145 39178
rect 1179 39144 1213 39178
rect 1247 39144 1281 39178
rect 1315 39144 1349 39178
rect 1383 39144 1417 39178
rect 1451 39144 1485 39178
rect 1519 39144 1553 39178
rect 1587 39144 1621 39178
rect 1655 39144 1689 39178
rect 1723 39144 1757 39178
rect 1791 39144 1825 39178
rect 1859 39144 1893 39178
rect 1927 39144 1961 39178
rect 1995 39144 2029 39178
rect 2063 39144 2097 39178
rect 2131 39144 2165 39178
rect 2199 39144 2233 39178
rect 2267 39144 2301 39178
rect 2335 39144 2369 39178
rect 2403 39144 2437 39178
rect 2471 39144 2505 39178
rect 2539 39144 2573 39178
rect 2607 39144 2641 39178
rect 2675 39144 2709 39178
rect 2743 39144 2777 39178
rect 2811 39144 2845 39178
rect 2879 39144 2913 39178
rect 2947 39144 2981 39178
rect 3015 39144 3083 39178
rect 373 39131 3083 39144
rect 373 39123 433 39131
rect 373 39089 386 39123
rect 420 39089 433 39123
rect 373 39055 433 39089
rect 3023 39110 3083 39131
rect 3023 39076 3036 39110
rect 3070 39076 3083 39110
rect 373 39021 386 39055
rect 420 39021 433 39055
rect 373 38987 433 39021
rect 3023 39042 3083 39076
rect 3023 39008 3036 39042
rect 3070 39008 3083 39042
rect 373 38953 386 38987
rect 420 38953 433 38987
rect 373 38919 433 38953
rect 373 38885 386 38919
rect 420 38885 433 38919
rect 373 38851 433 38885
rect 373 38817 386 38851
rect 420 38817 433 38851
rect 373 38783 433 38817
rect 373 38749 386 38783
rect 420 38749 433 38783
rect 373 38715 433 38749
rect 373 38681 386 38715
rect 420 38681 433 38715
rect 373 38647 433 38681
rect 373 38613 386 38647
rect 420 38613 433 38647
rect 373 38579 433 38613
rect 373 38545 386 38579
rect 420 38545 433 38579
rect 373 38511 433 38545
rect 373 38477 386 38511
rect 420 38477 433 38511
rect 373 38443 433 38477
rect 373 38409 386 38443
rect 420 38409 433 38443
rect 373 38375 433 38409
rect 373 38341 386 38375
rect 420 38341 433 38375
rect 373 38307 433 38341
rect 373 38273 386 38307
rect 420 38273 433 38307
rect 373 38239 433 38273
rect 373 38205 386 38239
rect 420 38205 433 38239
rect 373 38171 433 38205
rect 373 38137 386 38171
rect 420 38137 433 38171
rect 373 38103 433 38137
rect 373 38069 386 38103
rect 420 38069 433 38103
rect 373 38035 433 38069
rect 373 38001 386 38035
rect 420 38001 433 38035
rect 373 37967 433 38001
rect 373 37933 386 37967
rect 420 37933 433 37967
rect 373 37899 433 37933
rect 373 37865 386 37899
rect 420 37865 433 37899
rect 373 37831 433 37865
rect 373 37797 386 37831
rect 420 37797 433 37831
rect 373 37763 433 37797
rect 373 37729 386 37763
rect 420 37729 433 37763
rect 373 37695 433 37729
rect 373 37661 386 37695
rect 420 37661 433 37695
rect 373 37627 433 37661
rect 373 37593 386 37627
rect 420 37593 433 37627
rect 373 37559 433 37593
rect 373 37525 386 37559
rect 420 37525 433 37559
rect 373 37491 433 37525
rect 373 37457 386 37491
rect 420 37457 433 37491
rect 373 37423 433 37457
rect 373 37389 386 37423
rect 420 37389 433 37423
rect 373 37355 433 37389
rect 373 37321 386 37355
rect 420 37321 433 37355
rect 373 37287 433 37321
rect 373 37253 386 37287
rect 420 37253 433 37287
rect 373 37219 433 37253
rect 373 37185 386 37219
rect 420 37185 433 37219
rect 373 37151 433 37185
rect 373 37117 386 37151
rect 420 37117 433 37151
rect 373 37083 433 37117
rect 373 37049 386 37083
rect 420 37049 433 37083
rect 373 37015 433 37049
rect 373 36981 386 37015
rect 420 36981 433 37015
rect 373 36947 433 36981
rect 373 36913 386 36947
rect 420 36913 433 36947
rect 3023 38974 3083 39008
rect 3023 38940 3036 38974
rect 3070 38940 3083 38974
rect 3023 38906 3083 38940
rect 3023 38872 3036 38906
rect 3070 38872 3083 38906
rect 3023 38838 3083 38872
rect 3023 38804 3036 38838
rect 3070 38804 3083 38838
rect 3023 38770 3083 38804
rect 3023 38736 3036 38770
rect 3070 38736 3083 38770
rect 3023 38702 3083 38736
rect 3023 38668 3036 38702
rect 3070 38668 3083 38702
rect 3023 38634 3083 38668
rect 3023 38600 3036 38634
rect 3070 38600 3083 38634
rect 3023 38566 3083 38600
rect 3023 38532 3036 38566
rect 3070 38532 3083 38566
rect 3023 38498 3083 38532
rect 3023 38464 3036 38498
rect 3070 38464 3083 38498
rect 3023 38430 3083 38464
rect 3023 38396 3036 38430
rect 3070 38396 3083 38430
rect 3023 38362 3083 38396
rect 3023 38328 3036 38362
rect 3070 38328 3083 38362
rect 3023 38294 3083 38328
rect 3023 38260 3036 38294
rect 3070 38260 3083 38294
rect 3023 38226 3083 38260
rect 3023 38192 3036 38226
rect 3070 38192 3083 38226
rect 3023 38158 3083 38192
rect 3023 38124 3036 38158
rect 3070 38124 3083 38158
rect 3023 38090 3083 38124
rect 3023 38056 3036 38090
rect 3070 38056 3083 38090
rect 3023 38022 3083 38056
rect 3023 37988 3036 38022
rect 3070 37988 3083 38022
rect 3023 37954 3083 37988
rect 3023 37920 3036 37954
rect 3070 37920 3083 37954
rect 3023 37886 3083 37920
rect 3023 37852 3036 37886
rect 3070 37852 3083 37886
rect 3023 37818 3083 37852
rect 3023 37784 3036 37818
rect 3070 37784 3083 37818
rect 3023 37750 3083 37784
rect 3023 37716 3036 37750
rect 3070 37716 3083 37750
rect 3023 37682 3083 37716
rect 3023 37648 3036 37682
rect 3070 37648 3083 37682
rect 3023 37614 3083 37648
rect 3023 37580 3036 37614
rect 3070 37580 3083 37614
rect 3023 37546 3083 37580
rect 3023 37512 3036 37546
rect 3070 37512 3083 37546
rect 3023 37478 3083 37512
rect 3023 37444 3036 37478
rect 3070 37444 3083 37478
rect 3023 37410 3083 37444
rect 3023 37376 3036 37410
rect 3070 37376 3083 37410
rect 3023 37342 3083 37376
rect 3023 37308 3036 37342
rect 3070 37308 3083 37342
rect 3023 37274 3083 37308
rect 3023 37240 3036 37274
rect 3070 37240 3083 37274
rect 3023 37206 3083 37240
rect 3023 37172 3036 37206
rect 3070 37172 3083 37206
rect 3023 37138 3083 37172
rect 3023 37104 3036 37138
rect 3070 37104 3083 37138
rect 3023 37070 3083 37104
rect 3023 37036 3036 37070
rect 3070 37036 3083 37070
rect 3023 37002 3083 37036
rect 3023 36968 3036 37002
rect 3070 36968 3083 37002
rect 373 36879 433 36913
rect 373 36845 386 36879
rect 420 36845 433 36879
rect 3023 36934 3083 36968
rect 3023 36900 3036 36934
rect 3070 36900 3083 36934
rect 373 36811 433 36845
rect 373 36777 386 36811
rect 420 36777 433 36811
rect 373 36743 433 36777
rect 373 36709 386 36743
rect 420 36709 433 36743
rect 373 36675 433 36709
rect 373 36641 386 36675
rect 420 36641 433 36675
rect 373 36607 433 36641
rect 373 36573 386 36607
rect 420 36573 433 36607
rect 373 36539 433 36573
rect 373 36505 386 36539
rect 420 36505 433 36539
rect 373 36471 433 36505
rect 373 36437 386 36471
rect 420 36437 433 36471
rect 373 36403 433 36437
rect 373 36369 386 36403
rect 420 36369 433 36403
rect 373 36335 433 36369
rect 373 36301 386 36335
rect 420 36301 433 36335
rect 373 36267 433 36301
rect 373 36233 386 36267
rect 420 36233 433 36267
rect 373 36199 433 36233
rect 373 36165 386 36199
rect 420 36165 433 36199
rect 373 36131 433 36165
rect 373 36097 386 36131
rect 420 36097 433 36131
rect 373 36063 433 36097
rect 373 36029 386 36063
rect 420 36029 433 36063
rect 373 35995 433 36029
rect 373 35961 386 35995
rect 420 35961 433 35995
rect 373 35927 433 35961
rect 373 35893 386 35927
rect 420 35893 433 35927
rect 373 35859 433 35893
rect 373 35825 386 35859
rect 420 35825 433 35859
rect 373 35791 433 35825
rect 373 35757 386 35791
rect 420 35757 433 35791
rect 373 35723 433 35757
rect 373 35689 386 35723
rect 420 35689 433 35723
rect 373 35655 433 35689
rect 373 35621 386 35655
rect 420 35621 433 35655
rect 373 35587 433 35621
rect 373 35553 386 35587
rect 420 35553 433 35587
rect 373 35519 433 35553
rect 373 35485 386 35519
rect 420 35485 433 35519
rect 373 35451 433 35485
rect 373 35417 386 35451
rect 420 35417 433 35451
rect 373 35383 433 35417
rect 373 35349 386 35383
rect 420 35349 433 35383
rect 373 35315 433 35349
rect 373 35281 386 35315
rect 420 35281 433 35315
rect 373 35247 433 35281
rect 373 35213 386 35247
rect 420 35213 433 35247
rect 373 35179 433 35213
rect 373 35145 386 35179
rect 420 35145 433 35179
rect 373 35111 433 35145
rect 373 35077 386 35111
rect 420 35077 433 35111
rect 373 35043 433 35077
rect 373 35009 386 35043
rect 420 35009 433 35043
rect 373 34975 433 35009
rect 373 34941 386 34975
rect 420 34941 433 34975
rect 373 34907 433 34941
rect 373 34873 386 34907
rect 420 34873 433 34907
rect 373 34839 433 34873
rect 373 34805 386 34839
rect 420 34805 433 34839
rect 3023 36866 3083 36900
rect 3023 36832 3036 36866
rect 3070 36832 3083 36866
rect 3023 36798 3083 36832
rect 3023 36764 3036 36798
rect 3070 36764 3083 36798
rect 3023 36730 3083 36764
rect 3023 36696 3036 36730
rect 3070 36696 3083 36730
rect 3023 36662 3083 36696
rect 3023 36628 3036 36662
rect 3070 36628 3083 36662
rect 3023 36594 3083 36628
rect 3023 36560 3036 36594
rect 3070 36560 3083 36594
rect 3023 36526 3083 36560
rect 3023 36492 3036 36526
rect 3070 36492 3083 36526
rect 3023 36458 3083 36492
rect 3023 36424 3036 36458
rect 3070 36424 3083 36458
rect 3023 36390 3083 36424
rect 3023 36356 3036 36390
rect 3070 36356 3083 36390
rect 3023 36322 3083 36356
rect 3023 36288 3036 36322
rect 3070 36288 3083 36322
rect 3023 36254 3083 36288
rect 3023 36220 3036 36254
rect 3070 36220 3083 36254
rect 3023 36186 3083 36220
rect 3023 36152 3036 36186
rect 3070 36152 3083 36186
rect 3023 36118 3083 36152
rect 3023 36084 3036 36118
rect 3070 36084 3083 36118
rect 3023 36050 3083 36084
rect 3023 36016 3036 36050
rect 3070 36016 3083 36050
rect 3023 35982 3083 36016
rect 3023 35948 3036 35982
rect 3070 35948 3083 35982
rect 3023 35914 3083 35948
rect 3023 35880 3036 35914
rect 3070 35880 3083 35914
rect 3023 35846 3083 35880
rect 3023 35812 3036 35846
rect 3070 35812 3083 35846
rect 3023 35778 3083 35812
rect 3023 35744 3036 35778
rect 3070 35744 3083 35778
rect 3023 35710 3083 35744
rect 3023 35676 3036 35710
rect 3070 35676 3083 35710
rect 3023 35642 3083 35676
rect 3023 35608 3036 35642
rect 3070 35608 3083 35642
rect 3023 35574 3083 35608
rect 3023 35540 3036 35574
rect 3070 35540 3083 35574
rect 3023 35506 3083 35540
rect 3023 35472 3036 35506
rect 3070 35472 3083 35506
rect 3023 35438 3083 35472
rect 3023 35404 3036 35438
rect 3070 35404 3083 35438
rect 3023 35370 3083 35404
rect 3023 35336 3036 35370
rect 3070 35336 3083 35370
rect 3023 35302 3083 35336
rect 3023 35268 3036 35302
rect 3070 35268 3083 35302
rect 3023 35234 3083 35268
rect 3023 35200 3036 35234
rect 3070 35200 3083 35234
rect 3023 35166 3083 35200
rect 3023 35132 3036 35166
rect 3070 35132 3083 35166
rect 3023 35098 3083 35132
rect 3023 35064 3036 35098
rect 3070 35064 3083 35098
rect 3023 35030 3083 35064
rect 3023 34996 3036 35030
rect 3070 34996 3083 35030
rect 3023 34962 3083 34996
rect 3023 34928 3036 34962
rect 3070 34928 3083 34962
rect 3023 34894 3083 34928
rect 3023 34860 3036 34894
rect 3070 34860 3083 34894
rect 3023 34826 3083 34860
rect 373 34771 433 34805
rect 373 34737 386 34771
rect 420 34737 433 34771
rect 3023 34792 3036 34826
rect 3070 34792 3083 34826
rect 3023 34758 3083 34792
rect 373 34703 433 34737
rect 373 34669 386 34703
rect 420 34669 433 34703
rect 373 34635 433 34669
rect 373 34601 386 34635
rect 420 34601 433 34635
rect 373 34567 433 34601
rect 373 34533 386 34567
rect 420 34533 433 34567
rect 373 34499 433 34533
rect 373 34465 386 34499
rect 420 34465 433 34499
rect 373 34431 433 34465
rect 373 34397 386 34431
rect 420 34397 433 34431
rect 373 34363 433 34397
rect 373 34329 386 34363
rect 420 34329 433 34363
rect 373 34295 433 34329
rect 373 34261 386 34295
rect 420 34261 433 34295
rect 373 34227 433 34261
rect 373 34193 386 34227
rect 420 34193 433 34227
rect 373 34159 433 34193
rect 373 34125 386 34159
rect 420 34125 433 34159
rect 373 34091 433 34125
rect 373 34057 386 34091
rect 420 34057 433 34091
rect 373 34023 433 34057
rect 373 33989 386 34023
rect 420 33989 433 34023
rect 373 33955 433 33989
rect 373 33921 386 33955
rect 420 33921 433 33955
rect 373 33887 433 33921
rect 373 33853 386 33887
rect 420 33853 433 33887
rect 373 33819 433 33853
rect 373 33785 386 33819
rect 420 33785 433 33819
rect 373 33751 433 33785
rect 373 33717 386 33751
rect 420 33717 433 33751
rect 373 33683 433 33717
rect 373 33649 386 33683
rect 420 33649 433 33683
rect 373 33615 433 33649
rect 373 33581 386 33615
rect 420 33581 433 33615
rect 373 33547 433 33581
rect 373 33513 386 33547
rect 420 33513 433 33547
rect 373 33479 433 33513
rect 373 33445 386 33479
rect 420 33445 433 33479
rect 373 33411 433 33445
rect 373 33377 386 33411
rect 420 33377 433 33411
rect 373 33343 433 33377
rect 373 33309 386 33343
rect 420 33309 433 33343
rect 373 33275 433 33309
rect 373 33241 386 33275
rect 420 33241 433 33275
rect 373 33207 433 33241
rect 373 33173 386 33207
rect 420 33173 433 33207
rect 373 33139 433 33173
rect 373 33105 386 33139
rect 420 33105 433 33139
rect 373 33071 433 33105
rect 373 33037 386 33071
rect 420 33037 433 33071
rect 373 33003 433 33037
rect 373 32969 386 33003
rect 420 32969 433 33003
rect 373 32935 433 32969
rect 373 32901 386 32935
rect 420 32901 433 32935
rect 373 32867 433 32901
rect 373 32833 386 32867
rect 420 32833 433 32867
rect 373 32799 433 32833
rect 373 32765 386 32799
rect 420 32765 433 32799
rect 373 32731 433 32765
rect 373 32697 386 32731
rect 420 32697 433 32731
rect 373 32663 433 32697
rect 3023 34724 3036 34758
rect 3070 34724 3083 34758
rect 3023 34690 3083 34724
rect 3023 34656 3036 34690
rect 3070 34656 3083 34690
rect 3023 34622 3083 34656
rect 3023 34588 3036 34622
rect 3070 34588 3083 34622
rect 3023 34554 3083 34588
rect 3023 34520 3036 34554
rect 3070 34520 3083 34554
rect 3023 34486 3083 34520
rect 3023 34452 3036 34486
rect 3070 34452 3083 34486
rect 3023 34418 3083 34452
rect 3023 34384 3036 34418
rect 3070 34384 3083 34418
rect 3023 34350 3083 34384
rect 3023 34316 3036 34350
rect 3070 34316 3083 34350
rect 3023 34282 3083 34316
rect 3023 34248 3036 34282
rect 3070 34248 3083 34282
rect 3023 34214 3083 34248
rect 3023 34180 3036 34214
rect 3070 34180 3083 34214
rect 3023 34146 3083 34180
rect 3023 34112 3036 34146
rect 3070 34112 3083 34146
rect 3023 34078 3083 34112
rect 3023 34044 3036 34078
rect 3070 34044 3083 34078
rect 3023 34010 3083 34044
rect 3023 33976 3036 34010
rect 3070 33976 3083 34010
rect 3023 33942 3083 33976
rect 3023 33908 3036 33942
rect 3070 33908 3083 33942
rect 3023 33874 3083 33908
rect 3023 33840 3036 33874
rect 3070 33840 3083 33874
rect 3023 33806 3083 33840
rect 3023 33772 3036 33806
rect 3070 33772 3083 33806
rect 3023 33738 3083 33772
rect 3023 33704 3036 33738
rect 3070 33704 3083 33738
rect 3023 33670 3083 33704
rect 3023 33636 3036 33670
rect 3070 33636 3083 33670
rect 3023 33602 3083 33636
rect 3023 33568 3036 33602
rect 3070 33568 3083 33602
rect 3023 33534 3083 33568
rect 3023 33500 3036 33534
rect 3070 33500 3083 33534
rect 3023 33466 3083 33500
rect 3023 33432 3036 33466
rect 3070 33432 3083 33466
rect 3023 33398 3083 33432
rect 3023 33364 3036 33398
rect 3070 33364 3083 33398
rect 3023 33330 3083 33364
rect 3023 33296 3036 33330
rect 3070 33296 3083 33330
rect 3023 33262 3083 33296
rect 3023 33228 3036 33262
rect 3070 33228 3083 33262
rect 3023 33194 3083 33228
rect 3023 33160 3036 33194
rect 3070 33160 3083 33194
rect 3023 33126 3083 33160
rect 3023 33092 3036 33126
rect 3070 33092 3083 33126
rect 3023 33058 3083 33092
rect 3023 33024 3036 33058
rect 3070 33024 3083 33058
rect 3023 32990 3083 33024
rect 3023 32956 3036 32990
rect 3070 32956 3083 32990
rect 3023 32922 3083 32956
rect 3023 32888 3036 32922
rect 3070 32888 3083 32922
rect 3023 32854 3083 32888
rect 3023 32820 3036 32854
rect 3070 32820 3083 32854
rect 3023 32786 3083 32820
rect 3023 32752 3036 32786
rect 3070 32752 3083 32786
rect 3023 32718 3083 32752
rect 3023 32684 3036 32718
rect 3070 32684 3083 32718
rect 373 32629 386 32663
rect 420 32629 433 32663
rect 373 32595 433 32629
rect 3023 32650 3083 32684
rect 3023 32616 3036 32650
rect 3070 32616 3083 32650
rect 373 32561 386 32595
rect 420 32561 433 32595
rect 373 32527 433 32561
rect 373 32493 386 32527
rect 420 32493 433 32527
rect 373 32459 433 32493
rect 373 32425 386 32459
rect 420 32425 433 32459
rect 373 32391 433 32425
rect 373 32357 386 32391
rect 420 32357 433 32391
rect 373 32323 433 32357
rect 373 32289 386 32323
rect 420 32289 433 32323
rect 373 32255 433 32289
rect 373 32221 386 32255
rect 420 32221 433 32255
rect 373 32187 433 32221
rect 373 32153 386 32187
rect 420 32153 433 32187
rect 373 32119 433 32153
rect 373 32085 386 32119
rect 420 32085 433 32119
rect 373 32051 433 32085
rect 373 32017 386 32051
rect 420 32017 433 32051
rect 373 31983 433 32017
rect 373 31949 386 31983
rect 420 31949 433 31983
rect 373 31915 433 31949
rect 373 31881 386 31915
rect 420 31881 433 31915
rect 373 31847 433 31881
rect 373 31813 386 31847
rect 420 31813 433 31847
rect 373 31779 433 31813
rect 373 31745 386 31779
rect 420 31745 433 31779
rect 373 31711 433 31745
rect 373 31677 386 31711
rect 420 31677 433 31711
rect 373 31643 433 31677
rect 373 31609 386 31643
rect 420 31609 433 31643
rect 373 31575 433 31609
rect 373 31541 386 31575
rect 420 31541 433 31575
rect 373 31507 433 31541
rect 373 31473 386 31507
rect 420 31473 433 31507
rect 373 31439 433 31473
rect 373 31405 386 31439
rect 420 31405 433 31439
rect 373 31371 433 31405
rect 373 31337 386 31371
rect 420 31337 433 31371
rect 373 31303 433 31337
rect 373 31269 386 31303
rect 420 31269 433 31303
rect 373 31235 433 31269
rect 373 31201 386 31235
rect 420 31201 433 31235
rect 373 31167 433 31201
rect 373 31133 386 31167
rect 420 31133 433 31167
rect 373 31099 433 31133
rect 373 31065 386 31099
rect 420 31065 433 31099
rect 373 31031 433 31065
rect 373 30997 386 31031
rect 420 30997 433 31031
rect 373 30963 433 30997
rect 373 30929 386 30963
rect 420 30929 433 30963
rect 373 30895 433 30929
rect 373 30861 386 30895
rect 420 30861 433 30895
rect 373 30827 433 30861
rect 373 30793 386 30827
rect 420 30793 433 30827
rect 373 30759 433 30793
rect 373 30725 386 30759
rect 420 30725 433 30759
rect 373 30691 433 30725
rect 373 30657 386 30691
rect 420 30657 433 30691
rect 373 30623 433 30657
rect 373 30589 386 30623
rect 420 30589 433 30623
rect 373 30555 433 30589
rect 373 30521 386 30555
rect 420 30521 433 30555
rect 3023 32582 3083 32616
rect 3023 32548 3036 32582
rect 3070 32548 3083 32582
rect 3023 32514 3083 32548
rect 3023 32480 3036 32514
rect 3070 32480 3083 32514
rect 3023 32446 3083 32480
rect 3023 32412 3036 32446
rect 3070 32412 3083 32446
rect 3023 32378 3083 32412
rect 3023 32344 3036 32378
rect 3070 32344 3083 32378
rect 3023 32310 3083 32344
rect 3023 32276 3036 32310
rect 3070 32276 3083 32310
rect 3023 32242 3083 32276
rect 3023 32208 3036 32242
rect 3070 32208 3083 32242
rect 3023 32174 3083 32208
rect 3023 32140 3036 32174
rect 3070 32140 3083 32174
rect 3023 32106 3083 32140
rect 3023 32072 3036 32106
rect 3070 32072 3083 32106
rect 3023 32038 3083 32072
rect 3023 32004 3036 32038
rect 3070 32004 3083 32038
rect 3023 31970 3083 32004
rect 3023 31936 3036 31970
rect 3070 31936 3083 31970
rect 3023 31902 3083 31936
rect 3023 31868 3036 31902
rect 3070 31868 3083 31902
rect 3023 31834 3083 31868
rect 3023 31800 3036 31834
rect 3070 31800 3083 31834
rect 3023 31766 3083 31800
rect 3023 31732 3036 31766
rect 3070 31732 3083 31766
rect 3023 31698 3083 31732
rect 3023 31664 3036 31698
rect 3070 31664 3083 31698
rect 3023 31630 3083 31664
rect 3023 31596 3036 31630
rect 3070 31596 3083 31630
rect 3023 31562 3083 31596
rect 3023 31528 3036 31562
rect 3070 31528 3083 31562
rect 3023 31494 3083 31528
rect 3023 31460 3036 31494
rect 3070 31460 3083 31494
rect 3023 31426 3083 31460
rect 3023 31392 3036 31426
rect 3070 31392 3083 31426
rect 3023 31358 3083 31392
rect 3023 31324 3036 31358
rect 3070 31324 3083 31358
rect 3023 31290 3083 31324
rect 3023 31256 3036 31290
rect 3070 31256 3083 31290
rect 3023 31222 3083 31256
rect 3023 31188 3036 31222
rect 3070 31188 3083 31222
rect 3023 31154 3083 31188
rect 3023 31120 3036 31154
rect 3070 31120 3083 31154
rect 3023 31086 3083 31120
rect 3023 31052 3036 31086
rect 3070 31052 3083 31086
rect 3023 31018 3083 31052
rect 3023 30984 3036 31018
rect 3070 30984 3083 31018
rect 3023 30950 3083 30984
rect 3023 30916 3036 30950
rect 3070 30916 3083 30950
rect 3023 30882 3083 30916
rect 3023 30848 3036 30882
rect 3070 30848 3083 30882
rect 3023 30814 3083 30848
rect 3023 30780 3036 30814
rect 3070 30780 3083 30814
rect 3023 30746 3083 30780
rect 3023 30712 3036 30746
rect 3070 30712 3083 30746
rect 3023 30678 3083 30712
rect 3023 30644 3036 30678
rect 3070 30644 3083 30678
rect 3023 30610 3083 30644
rect 3023 30576 3036 30610
rect 3070 30576 3083 30610
rect 373 30487 433 30521
rect 373 30453 386 30487
rect 420 30453 433 30487
rect 3023 30542 3083 30576
rect 3023 30508 3036 30542
rect 3070 30508 3083 30542
rect 373 30419 433 30453
rect 373 30385 386 30419
rect 420 30385 433 30419
rect 373 30351 433 30385
rect 373 30317 386 30351
rect 420 30317 433 30351
rect 373 30283 433 30317
rect 373 30249 386 30283
rect 420 30249 433 30283
rect 373 30215 433 30249
rect 373 30181 386 30215
rect 420 30181 433 30215
rect 373 30147 433 30181
rect 373 30113 386 30147
rect 420 30113 433 30147
rect 373 30079 433 30113
rect 373 30045 386 30079
rect 420 30045 433 30079
rect 373 30011 433 30045
rect 373 29977 386 30011
rect 420 29977 433 30011
rect 373 29943 433 29977
rect 373 29909 386 29943
rect 420 29909 433 29943
rect 373 29875 433 29909
rect 373 29841 386 29875
rect 420 29841 433 29875
rect 373 29807 433 29841
rect 373 29773 386 29807
rect 420 29773 433 29807
rect 373 29739 433 29773
rect 373 29705 386 29739
rect 420 29705 433 29739
rect 373 29671 433 29705
rect 373 29637 386 29671
rect 420 29637 433 29671
rect 373 29603 433 29637
rect 373 29569 386 29603
rect 420 29569 433 29603
rect 373 29535 433 29569
rect 373 29501 386 29535
rect 420 29501 433 29535
rect 373 29467 433 29501
rect 373 29433 386 29467
rect 420 29433 433 29467
rect 373 29399 433 29433
rect 373 29365 386 29399
rect 420 29365 433 29399
rect 373 29331 433 29365
rect 373 29297 386 29331
rect 420 29297 433 29331
rect 373 29263 433 29297
rect 373 29229 386 29263
rect 420 29229 433 29263
rect 373 29195 433 29229
rect 373 29161 386 29195
rect 420 29161 433 29195
rect 373 29127 433 29161
rect 373 29093 386 29127
rect 420 29093 433 29127
rect 373 29059 433 29093
rect 373 29025 386 29059
rect 420 29025 433 29059
rect 373 28991 433 29025
rect 373 28957 386 28991
rect 420 28957 433 28991
rect 373 28923 433 28957
rect 373 28889 386 28923
rect 420 28889 433 28923
rect 373 28855 433 28889
rect 373 28821 386 28855
rect 420 28821 433 28855
rect 373 28787 433 28821
rect 373 28753 386 28787
rect 420 28753 433 28787
rect 373 28719 433 28753
rect 373 28685 386 28719
rect 420 28685 433 28719
rect 373 28651 433 28685
rect 373 28617 386 28651
rect 420 28617 433 28651
rect 373 28583 433 28617
rect 373 28549 386 28583
rect 420 28549 433 28583
rect 373 28515 433 28549
rect 373 28481 386 28515
rect 420 28481 433 28515
rect 373 28447 433 28481
rect 373 28413 386 28447
rect 420 28413 433 28447
rect 3023 30474 3083 30508
rect 3023 30440 3036 30474
rect 3070 30440 3083 30474
rect 3023 30406 3083 30440
rect 3023 30372 3036 30406
rect 3070 30372 3083 30406
rect 3023 30338 3083 30372
rect 3023 30304 3036 30338
rect 3070 30304 3083 30338
rect 3023 30270 3083 30304
rect 3023 30236 3036 30270
rect 3070 30236 3083 30270
rect 3023 30202 3083 30236
rect 3023 30168 3036 30202
rect 3070 30168 3083 30202
rect 3023 30134 3083 30168
rect 3023 30100 3036 30134
rect 3070 30100 3083 30134
rect 3023 30066 3083 30100
rect 3023 30032 3036 30066
rect 3070 30032 3083 30066
rect 3023 29998 3083 30032
rect 3023 29964 3036 29998
rect 3070 29964 3083 29998
rect 3023 29930 3083 29964
rect 3023 29896 3036 29930
rect 3070 29896 3083 29930
rect 3023 29862 3083 29896
rect 3023 29828 3036 29862
rect 3070 29828 3083 29862
rect 3023 29794 3083 29828
rect 3023 29760 3036 29794
rect 3070 29760 3083 29794
rect 3023 29726 3083 29760
rect 3023 29692 3036 29726
rect 3070 29692 3083 29726
rect 3023 29658 3083 29692
rect 3023 29624 3036 29658
rect 3070 29624 3083 29658
rect 3023 29590 3083 29624
rect 3023 29556 3036 29590
rect 3070 29556 3083 29590
rect 3023 29522 3083 29556
rect 3023 29488 3036 29522
rect 3070 29488 3083 29522
rect 3023 29454 3083 29488
rect 3023 29420 3036 29454
rect 3070 29420 3083 29454
rect 3023 29386 3083 29420
rect 3023 29352 3036 29386
rect 3070 29352 3083 29386
rect 3023 29318 3083 29352
rect 3023 29284 3036 29318
rect 3070 29284 3083 29318
rect 3023 29250 3083 29284
rect 3023 29216 3036 29250
rect 3070 29216 3083 29250
rect 3023 29182 3083 29216
rect 3023 29148 3036 29182
rect 3070 29148 3083 29182
rect 3023 29114 3083 29148
rect 3023 29080 3036 29114
rect 3070 29080 3083 29114
rect 3023 29046 3083 29080
rect 3023 29012 3036 29046
rect 3070 29012 3083 29046
rect 3023 28978 3083 29012
rect 3023 28944 3036 28978
rect 3070 28944 3083 28978
rect 3023 28910 3083 28944
rect 3023 28876 3036 28910
rect 3070 28876 3083 28910
rect 3023 28842 3083 28876
rect 3023 28808 3036 28842
rect 3070 28808 3083 28842
rect 3023 28774 3083 28808
rect 3023 28740 3036 28774
rect 3070 28740 3083 28774
rect 3023 28706 3083 28740
rect 3023 28672 3036 28706
rect 3070 28672 3083 28706
rect 3023 28638 3083 28672
rect 3023 28604 3036 28638
rect 3070 28604 3083 28638
rect 3023 28570 3083 28604
rect 3023 28536 3036 28570
rect 3070 28536 3083 28570
rect 3023 28502 3083 28536
rect 3023 28468 3036 28502
rect 3070 28468 3083 28502
rect 3023 28434 3083 28468
rect 373 28379 433 28413
rect 373 28345 386 28379
rect 420 28345 433 28379
rect 3023 28400 3036 28434
rect 3070 28400 3083 28434
rect 3023 28366 3083 28400
rect 373 28311 433 28345
rect 373 28277 386 28311
rect 420 28277 433 28311
rect 373 28243 433 28277
rect 373 28209 386 28243
rect 420 28209 433 28243
rect 373 28175 433 28209
rect 373 28141 386 28175
rect 420 28141 433 28175
rect 373 28107 433 28141
rect 373 28073 386 28107
rect 420 28073 433 28107
rect 373 28039 433 28073
rect 373 28005 386 28039
rect 420 28005 433 28039
rect 373 27971 433 28005
rect 373 27937 386 27971
rect 420 27937 433 27971
rect 373 27903 433 27937
rect 373 27869 386 27903
rect 420 27869 433 27903
rect 373 27835 433 27869
rect 373 27801 386 27835
rect 420 27801 433 27835
rect 373 27767 433 27801
rect 373 27733 386 27767
rect 420 27733 433 27767
rect 373 27699 433 27733
rect 373 27665 386 27699
rect 420 27665 433 27699
rect 373 27631 433 27665
rect 373 27597 386 27631
rect 420 27597 433 27631
rect 373 27563 433 27597
rect 373 27529 386 27563
rect 420 27529 433 27563
rect 373 27495 433 27529
rect 373 27461 386 27495
rect 420 27461 433 27495
rect 373 27427 433 27461
rect 373 27393 386 27427
rect 420 27393 433 27427
rect 373 27359 433 27393
rect 373 27325 386 27359
rect 420 27325 433 27359
rect 373 27291 433 27325
rect 373 27257 386 27291
rect 420 27257 433 27291
rect 373 27223 433 27257
rect 373 27189 386 27223
rect 420 27189 433 27223
rect 373 27155 433 27189
rect 373 27121 386 27155
rect 420 27121 433 27155
rect 373 27087 433 27121
rect 373 27053 386 27087
rect 420 27053 433 27087
rect 373 27019 433 27053
rect 373 26985 386 27019
rect 420 26985 433 27019
rect 373 26951 433 26985
rect 373 26917 386 26951
rect 420 26917 433 26951
rect 373 26883 433 26917
rect 373 26849 386 26883
rect 420 26849 433 26883
rect 373 26815 433 26849
rect 373 26781 386 26815
rect 420 26781 433 26815
rect 373 26747 433 26781
rect 373 26713 386 26747
rect 420 26713 433 26747
rect 373 26679 433 26713
rect 373 26645 386 26679
rect 420 26645 433 26679
rect 373 26611 433 26645
rect 373 26577 386 26611
rect 420 26577 433 26611
rect 373 26543 433 26577
rect 373 26509 386 26543
rect 420 26509 433 26543
rect 373 26475 433 26509
rect 373 26441 386 26475
rect 420 26441 433 26475
rect 373 26407 433 26441
rect 373 26373 386 26407
rect 420 26373 433 26407
rect 373 26339 433 26373
rect 373 26305 386 26339
rect 420 26305 433 26339
rect 373 26271 433 26305
rect 3023 28332 3036 28366
rect 3070 28332 3083 28366
rect 3023 28298 3083 28332
rect 3023 28264 3036 28298
rect 3070 28264 3083 28298
rect 3023 28230 3083 28264
rect 3023 28196 3036 28230
rect 3070 28196 3083 28230
rect 3023 28162 3083 28196
rect 3023 28128 3036 28162
rect 3070 28128 3083 28162
rect 3023 28094 3083 28128
rect 3023 28060 3036 28094
rect 3070 28060 3083 28094
rect 3023 28026 3083 28060
rect 3023 27992 3036 28026
rect 3070 27992 3083 28026
rect 3023 27958 3083 27992
rect 3023 27924 3036 27958
rect 3070 27924 3083 27958
rect 3023 27890 3083 27924
rect 3023 27856 3036 27890
rect 3070 27856 3083 27890
rect 3023 27822 3083 27856
rect 3023 27788 3036 27822
rect 3070 27788 3083 27822
rect 3023 27754 3083 27788
rect 3023 27720 3036 27754
rect 3070 27720 3083 27754
rect 3023 27686 3083 27720
rect 3023 27652 3036 27686
rect 3070 27652 3083 27686
rect 3023 27618 3083 27652
rect 3023 27584 3036 27618
rect 3070 27584 3083 27618
rect 3023 27550 3083 27584
rect 3023 27516 3036 27550
rect 3070 27516 3083 27550
rect 3023 27482 3083 27516
rect 3023 27448 3036 27482
rect 3070 27448 3083 27482
rect 3023 27414 3083 27448
rect 3023 27380 3036 27414
rect 3070 27380 3083 27414
rect 3023 27346 3083 27380
rect 3023 27312 3036 27346
rect 3070 27312 3083 27346
rect 3023 27278 3083 27312
rect 3023 27244 3036 27278
rect 3070 27244 3083 27278
rect 3023 27210 3083 27244
rect 3023 27176 3036 27210
rect 3070 27176 3083 27210
rect 3023 27142 3083 27176
rect 3023 27108 3036 27142
rect 3070 27108 3083 27142
rect 3023 27074 3083 27108
rect 3023 27040 3036 27074
rect 3070 27040 3083 27074
rect 3023 27006 3083 27040
rect 3023 26972 3036 27006
rect 3070 26972 3083 27006
rect 3023 26938 3083 26972
rect 3023 26904 3036 26938
rect 3070 26904 3083 26938
rect 3023 26870 3083 26904
rect 3023 26836 3036 26870
rect 3070 26836 3083 26870
rect 3023 26802 3083 26836
rect 3023 26768 3036 26802
rect 3070 26768 3083 26802
rect 3023 26734 3083 26768
rect 3023 26700 3036 26734
rect 3070 26700 3083 26734
rect 3023 26666 3083 26700
rect 3023 26632 3036 26666
rect 3070 26632 3083 26666
rect 3023 26598 3083 26632
rect 3023 26564 3036 26598
rect 3070 26564 3083 26598
rect 3023 26530 3083 26564
rect 3023 26496 3036 26530
rect 3070 26496 3083 26530
rect 3023 26462 3083 26496
rect 3023 26428 3036 26462
rect 3070 26428 3083 26462
rect 3023 26394 3083 26428
rect 3023 26360 3036 26394
rect 3070 26360 3083 26394
rect 3023 26326 3083 26360
rect 3023 26292 3036 26326
rect 3070 26292 3083 26326
rect 373 26237 386 26271
rect 420 26237 433 26271
rect 373 26203 433 26237
rect 3023 26258 3083 26292
rect 3023 26224 3036 26258
rect 3070 26224 3083 26258
rect 373 26169 386 26203
rect 420 26169 433 26203
rect 373 26135 433 26169
rect 373 26101 386 26135
rect 420 26101 433 26135
rect 373 26067 433 26101
rect 373 26033 386 26067
rect 420 26033 433 26067
rect 373 25999 433 26033
rect 373 25965 386 25999
rect 420 25965 433 25999
rect 373 25931 433 25965
rect 373 25897 386 25931
rect 420 25897 433 25931
rect 373 25863 433 25897
rect 373 25829 386 25863
rect 420 25829 433 25863
rect 373 25795 433 25829
rect 373 25761 386 25795
rect 420 25761 433 25795
rect 373 25727 433 25761
rect 373 25693 386 25727
rect 420 25693 433 25727
rect 373 25659 433 25693
rect 373 25625 386 25659
rect 420 25625 433 25659
rect 373 25591 433 25625
rect 373 25557 386 25591
rect 420 25557 433 25591
rect 373 25523 433 25557
rect 373 25489 386 25523
rect 420 25489 433 25523
rect 373 25455 433 25489
rect 373 25421 386 25455
rect 420 25421 433 25455
rect 373 25387 433 25421
rect 373 25353 386 25387
rect 420 25353 433 25387
rect 373 25319 433 25353
rect 373 25285 386 25319
rect 420 25285 433 25319
rect 373 25251 433 25285
rect 373 25217 386 25251
rect 420 25217 433 25251
rect 373 25183 433 25217
rect 373 25149 386 25183
rect 420 25149 433 25183
rect 373 25115 433 25149
rect 373 25081 386 25115
rect 420 25081 433 25115
rect 373 25047 433 25081
rect 373 25013 386 25047
rect 420 25013 433 25047
rect 373 24979 433 25013
rect 373 24945 386 24979
rect 420 24945 433 24979
rect 373 24911 433 24945
rect 373 24877 386 24911
rect 420 24877 433 24911
rect 373 24843 433 24877
rect 373 24809 386 24843
rect 420 24809 433 24843
rect 373 24775 433 24809
rect 373 24741 386 24775
rect 420 24741 433 24775
rect 373 24707 433 24741
rect 373 24673 386 24707
rect 420 24673 433 24707
rect 373 24639 433 24673
rect 373 24605 386 24639
rect 420 24605 433 24639
rect 373 24571 433 24605
rect 373 24537 386 24571
rect 420 24537 433 24571
rect 373 24503 433 24537
rect 373 24469 386 24503
rect 420 24469 433 24503
rect 373 24435 433 24469
rect 373 24401 386 24435
rect 420 24401 433 24435
rect 373 24367 433 24401
rect 373 24333 386 24367
rect 420 24333 433 24367
rect 373 24299 433 24333
rect 373 24265 386 24299
rect 420 24265 433 24299
rect 373 24231 433 24265
rect 373 24197 386 24231
rect 420 24197 433 24231
rect 373 24163 433 24197
rect 373 24129 386 24163
rect 420 24129 433 24163
rect 3023 26190 3083 26224
rect 3023 26156 3036 26190
rect 3070 26156 3083 26190
rect 3023 26122 3083 26156
rect 3023 26088 3036 26122
rect 3070 26088 3083 26122
rect 3023 26054 3083 26088
rect 3023 26020 3036 26054
rect 3070 26020 3083 26054
rect 3023 25986 3083 26020
rect 3023 25952 3036 25986
rect 3070 25952 3083 25986
rect 3023 25918 3083 25952
rect 3023 25884 3036 25918
rect 3070 25884 3083 25918
rect 3023 25850 3083 25884
rect 3023 25816 3036 25850
rect 3070 25816 3083 25850
rect 3023 25782 3083 25816
rect 3023 25748 3036 25782
rect 3070 25748 3083 25782
rect 3023 25714 3083 25748
rect 3023 25680 3036 25714
rect 3070 25680 3083 25714
rect 3023 25646 3083 25680
rect 3023 25612 3036 25646
rect 3070 25612 3083 25646
rect 3023 25578 3083 25612
rect 3023 25544 3036 25578
rect 3070 25544 3083 25578
rect 3023 25510 3083 25544
rect 3023 25476 3036 25510
rect 3070 25476 3083 25510
rect 3023 25442 3083 25476
rect 3023 25408 3036 25442
rect 3070 25408 3083 25442
rect 3023 25374 3083 25408
rect 3023 25340 3036 25374
rect 3070 25340 3083 25374
rect 3023 25306 3083 25340
rect 3023 25272 3036 25306
rect 3070 25272 3083 25306
rect 3023 25238 3083 25272
rect 3023 25204 3036 25238
rect 3070 25204 3083 25238
rect 3023 25170 3083 25204
rect 3023 25136 3036 25170
rect 3070 25136 3083 25170
rect 3023 25102 3083 25136
rect 3023 25068 3036 25102
rect 3070 25068 3083 25102
rect 3023 25034 3083 25068
rect 3023 25000 3036 25034
rect 3070 25000 3083 25034
rect 3023 24966 3083 25000
rect 3023 24932 3036 24966
rect 3070 24932 3083 24966
rect 3023 24898 3083 24932
rect 3023 24864 3036 24898
rect 3070 24864 3083 24898
rect 3023 24830 3083 24864
rect 3023 24796 3036 24830
rect 3070 24796 3083 24830
rect 3023 24762 3083 24796
rect 3023 24728 3036 24762
rect 3070 24728 3083 24762
rect 3023 24694 3083 24728
rect 3023 24660 3036 24694
rect 3070 24660 3083 24694
rect 3023 24626 3083 24660
rect 3023 24592 3036 24626
rect 3070 24592 3083 24626
rect 3023 24558 3083 24592
rect 3023 24524 3036 24558
rect 3070 24524 3083 24558
rect 3023 24490 3083 24524
rect 3023 24456 3036 24490
rect 3070 24456 3083 24490
rect 3023 24422 3083 24456
rect 3023 24388 3036 24422
rect 3070 24388 3083 24422
rect 3023 24354 3083 24388
rect 3023 24320 3036 24354
rect 3070 24320 3083 24354
rect 3023 24286 3083 24320
rect 3023 24252 3036 24286
rect 3070 24252 3083 24286
rect 3023 24218 3083 24252
rect 3023 24184 3036 24218
rect 3070 24184 3083 24218
rect 373 24095 433 24129
rect 373 24061 386 24095
rect 420 24061 433 24095
rect 3023 24150 3083 24184
rect 3023 24116 3036 24150
rect 3070 24116 3083 24150
rect 373 24027 433 24061
rect 373 23993 386 24027
rect 420 23993 433 24027
rect 373 23959 433 23993
rect 373 23925 386 23959
rect 420 23925 433 23959
rect 373 23891 433 23925
rect 373 23857 386 23891
rect 420 23857 433 23891
rect 373 23823 433 23857
rect 373 23789 386 23823
rect 420 23789 433 23823
rect 373 23755 433 23789
rect 373 23721 386 23755
rect 420 23721 433 23755
rect 373 23687 433 23721
rect 373 23653 386 23687
rect 420 23653 433 23687
rect 373 23619 433 23653
rect 373 23585 386 23619
rect 420 23585 433 23619
rect 373 23551 433 23585
rect 373 23517 386 23551
rect 420 23517 433 23551
rect 373 23483 433 23517
rect 373 23449 386 23483
rect 420 23449 433 23483
rect 373 23415 433 23449
rect 373 23381 386 23415
rect 420 23381 433 23415
rect 373 23347 433 23381
rect 373 23313 386 23347
rect 420 23313 433 23347
rect 373 23279 433 23313
rect 373 23245 386 23279
rect 420 23245 433 23279
rect 373 23211 433 23245
rect 373 23177 386 23211
rect 420 23177 433 23211
rect 373 23143 433 23177
rect 373 23109 386 23143
rect 420 23109 433 23143
rect 373 23075 433 23109
rect 373 23041 386 23075
rect 420 23041 433 23075
rect 373 23007 433 23041
rect 373 22973 386 23007
rect 420 22973 433 23007
rect 373 22939 433 22973
rect 373 22905 386 22939
rect 420 22905 433 22939
rect 373 22871 433 22905
rect 373 22837 386 22871
rect 420 22837 433 22871
rect 373 22803 433 22837
rect 373 22769 386 22803
rect 420 22769 433 22803
rect 373 22735 433 22769
rect 373 22701 386 22735
rect 420 22701 433 22735
rect 373 22667 433 22701
rect 373 22633 386 22667
rect 420 22633 433 22667
rect 373 22599 433 22633
rect 373 22565 386 22599
rect 420 22565 433 22599
rect 373 22531 433 22565
rect 373 22497 386 22531
rect 420 22497 433 22531
rect 373 22463 433 22497
rect 373 22429 386 22463
rect 420 22429 433 22463
rect 373 22395 433 22429
rect 373 22361 386 22395
rect 420 22361 433 22395
rect 373 22327 433 22361
rect 373 22293 386 22327
rect 420 22293 433 22327
rect 373 22259 433 22293
rect 373 22225 386 22259
rect 420 22225 433 22259
rect 373 22191 433 22225
rect 373 22157 386 22191
rect 420 22157 433 22191
rect 373 22123 433 22157
rect 373 22089 386 22123
rect 420 22089 433 22123
rect 373 22055 433 22089
rect 373 22021 386 22055
rect 420 22021 433 22055
rect 3023 24082 3083 24116
rect 3023 24048 3036 24082
rect 3070 24048 3083 24082
rect 3023 24014 3083 24048
rect 3023 23980 3036 24014
rect 3070 23980 3083 24014
rect 3023 23946 3083 23980
rect 3023 23912 3036 23946
rect 3070 23912 3083 23946
rect 3023 23878 3083 23912
rect 3023 23844 3036 23878
rect 3070 23844 3083 23878
rect 3023 23810 3083 23844
rect 3023 23776 3036 23810
rect 3070 23776 3083 23810
rect 3023 23742 3083 23776
rect 3023 23708 3036 23742
rect 3070 23708 3083 23742
rect 3023 23674 3083 23708
rect 3023 23640 3036 23674
rect 3070 23640 3083 23674
rect 3023 23606 3083 23640
rect 3023 23572 3036 23606
rect 3070 23572 3083 23606
rect 3023 23538 3083 23572
rect 3023 23504 3036 23538
rect 3070 23504 3083 23538
rect 3023 23470 3083 23504
rect 3023 23436 3036 23470
rect 3070 23436 3083 23470
rect 3023 23402 3083 23436
rect 3023 23368 3036 23402
rect 3070 23368 3083 23402
rect 3023 23334 3083 23368
rect 3023 23300 3036 23334
rect 3070 23300 3083 23334
rect 3023 23266 3083 23300
rect 3023 23232 3036 23266
rect 3070 23232 3083 23266
rect 3023 23198 3083 23232
rect 3023 23164 3036 23198
rect 3070 23164 3083 23198
rect 3023 23130 3083 23164
rect 3023 23096 3036 23130
rect 3070 23096 3083 23130
rect 3023 23062 3083 23096
rect 3023 23028 3036 23062
rect 3070 23028 3083 23062
rect 3023 22994 3083 23028
rect 3023 22960 3036 22994
rect 3070 22960 3083 22994
rect 3023 22926 3083 22960
rect 3023 22892 3036 22926
rect 3070 22892 3083 22926
rect 3023 22858 3083 22892
rect 3023 22824 3036 22858
rect 3070 22824 3083 22858
rect 3023 22790 3083 22824
rect 3023 22756 3036 22790
rect 3070 22756 3083 22790
rect 3023 22722 3083 22756
rect 3023 22688 3036 22722
rect 3070 22688 3083 22722
rect 3023 22654 3083 22688
rect 3023 22620 3036 22654
rect 3070 22620 3083 22654
rect 3023 22586 3083 22620
rect 3023 22552 3036 22586
rect 3070 22552 3083 22586
rect 3023 22518 3083 22552
rect 3023 22484 3036 22518
rect 3070 22484 3083 22518
rect 3023 22450 3083 22484
rect 3023 22416 3036 22450
rect 3070 22416 3083 22450
rect 3023 22382 3083 22416
rect 3023 22348 3036 22382
rect 3070 22348 3083 22382
rect 3023 22314 3083 22348
rect 3023 22280 3036 22314
rect 3070 22280 3083 22314
rect 3023 22246 3083 22280
rect 3023 22212 3036 22246
rect 3070 22212 3083 22246
rect 3023 22178 3083 22212
rect 3023 22144 3036 22178
rect 3070 22144 3083 22178
rect 3023 22110 3083 22144
rect 3023 22076 3036 22110
rect 3070 22076 3083 22110
rect 3023 22042 3083 22076
rect 373 21987 433 22021
rect 373 21953 386 21987
rect 420 21953 433 21987
rect 3023 22008 3036 22042
rect 3070 22008 3083 22042
rect 3023 21974 3083 22008
rect 373 21919 433 21953
rect 373 21885 386 21919
rect 420 21885 433 21919
rect 373 21851 433 21885
rect 373 21817 386 21851
rect 420 21817 433 21851
rect 373 21783 433 21817
rect 373 21749 386 21783
rect 420 21749 433 21783
rect 373 21715 433 21749
rect 373 21681 386 21715
rect 420 21681 433 21715
rect 373 21647 433 21681
rect 373 21613 386 21647
rect 420 21613 433 21647
rect 373 21579 433 21613
rect 373 21545 386 21579
rect 420 21545 433 21579
rect 373 21511 433 21545
rect 373 21477 386 21511
rect 420 21477 433 21511
rect 373 21443 433 21477
rect 373 21409 386 21443
rect 420 21409 433 21443
rect 373 21375 433 21409
rect 373 21341 386 21375
rect 420 21341 433 21375
rect 373 21307 433 21341
rect 373 21273 386 21307
rect 420 21273 433 21307
rect 373 21239 433 21273
rect 373 21205 386 21239
rect 420 21205 433 21239
rect 373 21171 433 21205
rect 373 21137 386 21171
rect 420 21137 433 21171
rect 373 21103 433 21137
rect 373 21069 386 21103
rect 420 21069 433 21103
rect 373 21035 433 21069
rect 373 21001 386 21035
rect 420 21001 433 21035
rect 373 20967 433 21001
rect 373 20933 386 20967
rect 420 20933 433 20967
rect 373 20899 433 20933
rect 373 20865 386 20899
rect 420 20865 433 20899
rect 373 20831 433 20865
rect 373 20797 386 20831
rect 420 20797 433 20831
rect 373 20763 433 20797
rect 373 20729 386 20763
rect 420 20729 433 20763
rect 373 20695 433 20729
rect 373 20661 386 20695
rect 420 20661 433 20695
rect 373 20627 433 20661
rect 373 20593 386 20627
rect 420 20593 433 20627
rect 373 20559 433 20593
rect 373 20525 386 20559
rect 420 20525 433 20559
rect 373 20491 433 20525
rect 373 20457 386 20491
rect 420 20457 433 20491
rect 373 20423 433 20457
rect 373 20389 386 20423
rect 420 20389 433 20423
rect 373 20355 433 20389
rect 373 20321 386 20355
rect 420 20321 433 20355
rect 373 20287 433 20321
rect 373 20253 386 20287
rect 420 20253 433 20287
rect 373 20219 433 20253
rect 373 20185 386 20219
rect 420 20185 433 20219
rect 373 20151 433 20185
rect 373 20117 386 20151
rect 420 20117 433 20151
rect 373 20083 433 20117
rect 373 20049 386 20083
rect 420 20049 433 20083
rect 373 20015 433 20049
rect 373 19981 386 20015
rect 420 19981 433 20015
rect 373 19947 433 19981
rect 373 19913 386 19947
rect 420 19913 433 19947
rect 373 19879 433 19913
rect 3023 21940 3036 21974
rect 3070 21940 3083 21974
rect 3023 21906 3083 21940
rect 3023 21872 3036 21906
rect 3070 21872 3083 21906
rect 3023 21838 3083 21872
rect 3023 21804 3036 21838
rect 3070 21804 3083 21838
rect 3023 21770 3083 21804
rect 3023 21736 3036 21770
rect 3070 21736 3083 21770
rect 3023 21702 3083 21736
rect 3023 21668 3036 21702
rect 3070 21668 3083 21702
rect 3023 21634 3083 21668
rect 3023 21600 3036 21634
rect 3070 21600 3083 21634
rect 3023 21566 3083 21600
rect 3023 21532 3036 21566
rect 3070 21532 3083 21566
rect 3023 21498 3083 21532
rect 3023 21464 3036 21498
rect 3070 21464 3083 21498
rect 3023 21430 3083 21464
rect 3023 21396 3036 21430
rect 3070 21396 3083 21430
rect 3023 21362 3083 21396
rect 3023 21328 3036 21362
rect 3070 21328 3083 21362
rect 3023 21294 3083 21328
rect 3023 21260 3036 21294
rect 3070 21260 3083 21294
rect 3023 21226 3083 21260
rect 3023 21192 3036 21226
rect 3070 21192 3083 21226
rect 3023 21158 3083 21192
rect 3023 21124 3036 21158
rect 3070 21124 3083 21158
rect 3023 21090 3083 21124
rect 3023 21056 3036 21090
rect 3070 21056 3083 21090
rect 3023 21022 3083 21056
rect 3023 20988 3036 21022
rect 3070 20988 3083 21022
rect 3023 20954 3083 20988
rect 3023 20920 3036 20954
rect 3070 20920 3083 20954
rect 3023 20886 3083 20920
rect 3023 20852 3036 20886
rect 3070 20852 3083 20886
rect 3023 20818 3083 20852
rect 3023 20784 3036 20818
rect 3070 20784 3083 20818
rect 3023 20750 3083 20784
rect 3023 20716 3036 20750
rect 3070 20716 3083 20750
rect 3023 20682 3083 20716
rect 3023 20648 3036 20682
rect 3070 20648 3083 20682
rect 3023 20614 3083 20648
rect 3023 20580 3036 20614
rect 3070 20580 3083 20614
rect 3023 20546 3083 20580
rect 3023 20512 3036 20546
rect 3070 20512 3083 20546
rect 3023 20478 3083 20512
rect 3023 20444 3036 20478
rect 3070 20444 3083 20478
rect 3023 20410 3083 20444
rect 3023 20376 3036 20410
rect 3070 20376 3083 20410
rect 3023 20342 3083 20376
rect 3023 20308 3036 20342
rect 3070 20308 3083 20342
rect 3023 20274 3083 20308
rect 3023 20240 3036 20274
rect 3070 20240 3083 20274
rect 3023 20206 3083 20240
rect 3023 20172 3036 20206
rect 3070 20172 3083 20206
rect 3023 20138 3083 20172
rect 3023 20104 3036 20138
rect 3070 20104 3083 20138
rect 3023 20070 3083 20104
rect 3023 20036 3036 20070
rect 3070 20036 3083 20070
rect 3023 20002 3083 20036
rect 3023 19968 3036 20002
rect 3070 19968 3083 20002
rect 3023 19934 3083 19968
rect 3023 19900 3036 19934
rect 3070 19900 3083 19934
rect 373 19845 386 19879
rect 420 19845 433 19879
rect 373 19811 433 19845
rect 3023 19866 3083 19900
rect 373 19777 386 19811
rect 420 19777 433 19811
rect 373 19743 433 19777
rect 373 19709 386 19743
rect 420 19709 433 19743
rect 373 19675 433 19709
rect 373 19641 386 19675
rect 420 19641 433 19675
rect 373 19607 433 19641
rect 373 19573 386 19607
rect 420 19573 433 19607
rect 373 19539 433 19573
rect 373 19505 386 19539
rect 420 19505 433 19539
rect 373 19471 433 19505
rect 373 19437 386 19471
rect 420 19437 433 19471
rect 373 19403 433 19437
rect 373 19369 386 19403
rect 420 19369 433 19403
rect 373 19335 433 19369
rect 373 19301 386 19335
rect 420 19301 433 19335
rect 373 19267 433 19301
rect 373 19233 386 19267
rect 420 19233 433 19267
rect 373 19199 433 19233
rect 373 19165 386 19199
rect 420 19165 433 19199
rect 373 19131 433 19165
rect 373 19097 386 19131
rect 420 19097 433 19131
rect 373 19063 433 19097
rect 373 19029 386 19063
rect 420 19029 433 19063
rect 373 18995 433 19029
rect 373 18961 386 18995
rect 420 18961 433 18995
rect 373 18927 433 18961
rect 373 18893 386 18927
rect 420 18893 433 18927
rect 373 18859 433 18893
rect 373 18825 386 18859
rect 420 18825 433 18859
rect 373 18791 433 18825
rect 373 18757 386 18791
rect 420 18757 433 18791
rect 373 18723 433 18757
rect 373 18689 386 18723
rect 420 18689 433 18723
rect 373 18655 433 18689
rect 373 18621 386 18655
rect 420 18621 433 18655
rect 373 18587 433 18621
rect 373 18553 386 18587
rect 420 18553 433 18587
rect 373 18519 433 18553
rect 373 18485 386 18519
rect 420 18485 433 18519
rect 373 18451 433 18485
rect 373 18417 386 18451
rect 420 18417 433 18451
rect 373 18383 433 18417
rect 373 18349 386 18383
rect 420 18349 433 18383
rect 373 18315 433 18349
rect 373 18281 386 18315
rect 420 18281 433 18315
rect 373 18247 433 18281
rect 373 18213 386 18247
rect 420 18213 433 18247
rect 373 18179 433 18213
rect 373 18145 386 18179
rect 420 18145 433 18179
rect 373 18111 433 18145
rect 373 18077 386 18111
rect 420 18077 433 18111
rect 373 18043 433 18077
rect 373 18009 386 18043
rect 420 18009 433 18043
rect 373 17975 433 18009
rect 373 17941 386 17975
rect 420 17941 433 17975
rect 373 17907 433 17941
rect 373 17873 386 17907
rect 420 17873 433 17907
rect 373 17839 433 17873
rect 373 17805 386 17839
rect 420 17805 433 17839
rect 373 17771 433 17805
rect 373 17737 386 17771
rect 420 17737 433 17771
rect 3023 19832 3036 19866
rect 3070 19832 3083 19866
rect 3023 19798 3083 19832
rect 3023 19764 3036 19798
rect 3070 19764 3083 19798
rect 3023 19730 3083 19764
rect 3023 19696 3036 19730
rect 3070 19696 3083 19730
rect 3023 19662 3083 19696
rect 3023 19628 3036 19662
rect 3070 19628 3083 19662
rect 3023 19594 3083 19628
rect 3023 19560 3036 19594
rect 3070 19560 3083 19594
rect 3023 19526 3083 19560
rect 3023 19492 3036 19526
rect 3070 19492 3083 19526
rect 3023 19458 3083 19492
rect 3023 19424 3036 19458
rect 3070 19424 3083 19458
rect 3023 19390 3083 19424
rect 3023 19356 3036 19390
rect 3070 19356 3083 19390
rect 3023 19322 3083 19356
rect 3023 19288 3036 19322
rect 3070 19288 3083 19322
rect 3023 19254 3083 19288
rect 3023 19220 3036 19254
rect 3070 19220 3083 19254
rect 3023 19186 3083 19220
rect 3023 19152 3036 19186
rect 3070 19152 3083 19186
rect 3023 19118 3083 19152
rect 3023 19084 3036 19118
rect 3070 19084 3083 19118
rect 3023 19050 3083 19084
rect 3023 19016 3036 19050
rect 3070 19016 3083 19050
rect 3023 18982 3083 19016
rect 3023 18948 3036 18982
rect 3070 18948 3083 18982
rect 3023 18914 3083 18948
rect 3023 18880 3036 18914
rect 3070 18880 3083 18914
rect 3023 18846 3083 18880
rect 3023 18812 3036 18846
rect 3070 18812 3083 18846
rect 3023 18778 3083 18812
rect 3023 18744 3036 18778
rect 3070 18744 3083 18778
rect 3023 18710 3083 18744
rect 3023 18676 3036 18710
rect 3070 18676 3083 18710
rect 3023 18642 3083 18676
rect 3023 18608 3036 18642
rect 3070 18608 3083 18642
rect 3023 18574 3083 18608
rect 3023 18540 3036 18574
rect 3070 18540 3083 18574
rect 3023 18506 3083 18540
rect 3023 18472 3036 18506
rect 3070 18472 3083 18506
rect 3023 18438 3083 18472
rect 3023 18404 3036 18438
rect 3070 18404 3083 18438
rect 3023 18370 3083 18404
rect 3023 18336 3036 18370
rect 3070 18336 3083 18370
rect 3023 18302 3083 18336
rect 3023 18268 3036 18302
rect 3070 18268 3083 18302
rect 3023 18234 3083 18268
rect 3023 18200 3036 18234
rect 3070 18200 3083 18234
rect 3023 18166 3083 18200
rect 3023 18132 3036 18166
rect 3070 18132 3083 18166
rect 3023 18098 3083 18132
rect 3023 18064 3036 18098
rect 3070 18064 3083 18098
rect 3023 18030 3083 18064
rect 3023 17996 3036 18030
rect 3070 17996 3083 18030
rect 3023 17962 3083 17996
rect 3023 17928 3036 17962
rect 3070 17928 3083 17962
rect 3023 17894 3083 17928
rect 3023 17860 3036 17894
rect 3070 17860 3083 17894
rect 3023 17826 3083 17860
rect 3023 17792 3036 17826
rect 3070 17792 3083 17826
rect 373 17703 433 17737
rect 3023 17758 3083 17792
rect 3023 17724 3036 17758
rect 3070 17724 3083 17758
rect 373 17669 386 17703
rect 420 17669 433 17703
rect 373 17635 433 17669
rect 373 17601 386 17635
rect 420 17601 433 17635
rect 373 17567 433 17601
rect 373 17533 386 17567
rect 420 17533 433 17567
rect 373 17499 433 17533
rect 373 17465 386 17499
rect 420 17465 433 17499
rect 373 17431 433 17465
rect 373 17397 386 17431
rect 420 17397 433 17431
rect 373 17363 433 17397
rect 373 17329 386 17363
rect 420 17329 433 17363
rect 373 17295 433 17329
rect 373 17261 386 17295
rect 420 17261 433 17295
rect 373 17227 433 17261
rect 373 17193 386 17227
rect 420 17193 433 17227
rect 373 17159 433 17193
rect 373 17125 386 17159
rect 420 17125 433 17159
rect 373 17091 433 17125
rect 373 17057 386 17091
rect 420 17057 433 17091
rect 373 17023 433 17057
rect 373 16989 386 17023
rect 420 16989 433 17023
rect 373 16955 433 16989
rect 373 16921 386 16955
rect 420 16921 433 16955
rect 373 16887 433 16921
rect 373 16853 386 16887
rect 420 16853 433 16887
rect 373 16819 433 16853
rect 373 16785 386 16819
rect 420 16785 433 16819
rect 373 16751 433 16785
rect 373 16717 386 16751
rect 420 16717 433 16751
rect 373 16683 433 16717
rect 373 16649 386 16683
rect 420 16649 433 16683
rect 373 16615 433 16649
rect 373 16581 386 16615
rect 420 16581 433 16615
rect 373 16547 433 16581
rect 373 16513 386 16547
rect 420 16513 433 16547
rect 373 16479 433 16513
rect 373 16445 386 16479
rect 420 16445 433 16479
rect 373 16411 433 16445
rect 373 16377 386 16411
rect 420 16377 433 16411
rect 373 16343 433 16377
rect 373 16309 386 16343
rect 420 16309 433 16343
rect 373 16275 433 16309
rect 373 16241 386 16275
rect 420 16241 433 16275
rect 373 16207 433 16241
rect 373 16173 386 16207
rect 420 16173 433 16207
rect 373 16139 433 16173
rect 373 16105 386 16139
rect 420 16105 433 16139
rect 373 16071 433 16105
rect 373 16037 386 16071
rect 420 16037 433 16071
rect 373 16003 433 16037
rect 373 15969 386 16003
rect 420 15969 433 16003
rect 373 15935 433 15969
rect 373 15901 386 15935
rect 420 15901 433 15935
rect 373 15867 433 15901
rect 373 15833 386 15867
rect 420 15833 433 15867
rect 373 15799 433 15833
rect 373 15765 386 15799
rect 420 15765 433 15799
rect 373 15731 433 15765
rect 373 15697 386 15731
rect 420 15697 433 15731
rect 373 15663 433 15697
rect 373 15629 386 15663
rect 420 15629 433 15663
rect 3023 17690 3083 17724
rect 3023 17656 3036 17690
rect 3070 17656 3083 17690
rect 3023 17622 3083 17656
rect 3023 17588 3036 17622
rect 3070 17588 3083 17622
rect 3023 17554 3083 17588
rect 3023 17520 3036 17554
rect 3070 17520 3083 17554
rect 3023 17486 3083 17520
rect 3023 17452 3036 17486
rect 3070 17452 3083 17486
rect 3023 17418 3083 17452
rect 3023 17384 3036 17418
rect 3070 17384 3083 17418
rect 3023 17350 3083 17384
rect 3023 17316 3036 17350
rect 3070 17316 3083 17350
rect 3023 17282 3083 17316
rect 3023 17248 3036 17282
rect 3070 17248 3083 17282
rect 3023 17214 3083 17248
rect 3023 17180 3036 17214
rect 3070 17180 3083 17214
rect 3023 17146 3083 17180
rect 3023 17112 3036 17146
rect 3070 17112 3083 17146
rect 3023 17078 3083 17112
rect 3023 17044 3036 17078
rect 3070 17044 3083 17078
rect 3023 17010 3083 17044
rect 3023 16976 3036 17010
rect 3070 16976 3083 17010
rect 3023 16942 3083 16976
rect 3023 16908 3036 16942
rect 3070 16908 3083 16942
rect 3023 16874 3083 16908
rect 3023 16840 3036 16874
rect 3070 16840 3083 16874
rect 3023 16806 3083 16840
rect 3023 16772 3036 16806
rect 3070 16772 3083 16806
rect 3023 16738 3083 16772
rect 3023 16704 3036 16738
rect 3070 16704 3083 16738
rect 3023 16670 3083 16704
rect 3023 16636 3036 16670
rect 3070 16636 3083 16670
rect 3023 16602 3083 16636
rect 3023 16568 3036 16602
rect 3070 16568 3083 16602
rect 3023 16534 3083 16568
rect 3023 16500 3036 16534
rect 3070 16500 3083 16534
rect 3023 16466 3083 16500
rect 3023 16432 3036 16466
rect 3070 16432 3083 16466
rect 3023 16398 3083 16432
rect 3023 16364 3036 16398
rect 3070 16364 3083 16398
rect 3023 16330 3083 16364
rect 3023 16296 3036 16330
rect 3070 16296 3083 16330
rect 3023 16262 3083 16296
rect 3023 16228 3036 16262
rect 3070 16228 3083 16262
rect 3023 16194 3083 16228
rect 3023 16160 3036 16194
rect 3070 16160 3083 16194
rect 3023 16126 3083 16160
rect 3023 16092 3036 16126
rect 3070 16092 3083 16126
rect 3023 16058 3083 16092
rect 3023 16024 3036 16058
rect 3070 16024 3083 16058
rect 3023 15990 3083 16024
rect 3023 15956 3036 15990
rect 3070 15956 3083 15990
rect 3023 15922 3083 15956
rect 3023 15888 3036 15922
rect 3070 15888 3083 15922
rect 3023 15854 3083 15888
rect 3023 15820 3036 15854
rect 3070 15820 3083 15854
rect 3023 15786 3083 15820
rect 3023 15752 3036 15786
rect 3070 15752 3083 15786
rect 3023 15718 3083 15752
rect 3023 15684 3036 15718
rect 3070 15684 3083 15718
rect 3023 15650 3083 15684
rect 373 15595 433 15629
rect 373 15561 386 15595
rect 420 15561 433 15595
rect 3023 15616 3036 15650
rect 3070 15616 3083 15650
rect 3023 15582 3083 15616
rect 373 15527 433 15561
rect 373 15493 386 15527
rect 420 15493 433 15527
rect 373 15459 433 15493
rect 373 15425 386 15459
rect 420 15425 433 15459
rect 373 15391 433 15425
rect 373 15357 386 15391
rect 420 15357 433 15391
rect 373 15323 433 15357
rect 373 15289 386 15323
rect 420 15289 433 15323
rect 373 15255 433 15289
rect 373 15221 386 15255
rect 420 15221 433 15255
rect 373 15187 433 15221
rect 373 15153 386 15187
rect 420 15153 433 15187
rect 373 15119 433 15153
rect 373 15085 386 15119
rect 420 15085 433 15119
rect 373 15051 433 15085
rect 373 15017 386 15051
rect 420 15017 433 15051
rect 373 14983 433 15017
rect 373 14949 386 14983
rect 420 14949 433 14983
rect 373 14915 433 14949
rect 373 14881 386 14915
rect 420 14881 433 14915
rect 373 14847 433 14881
rect 373 14813 386 14847
rect 420 14813 433 14847
rect 373 14779 433 14813
rect 373 14745 386 14779
rect 420 14745 433 14779
rect 373 14711 433 14745
rect 373 14677 386 14711
rect 420 14677 433 14711
rect 373 14643 433 14677
rect 373 14609 386 14643
rect 420 14609 433 14643
rect 373 14575 433 14609
rect 373 14541 386 14575
rect 420 14541 433 14575
rect 373 14507 433 14541
rect 373 14473 386 14507
rect 420 14473 433 14507
rect 373 14439 433 14473
rect 373 14405 386 14439
rect 420 14405 433 14439
rect 373 14371 433 14405
rect 373 14337 386 14371
rect 420 14337 433 14371
rect 373 14303 433 14337
rect 373 14269 386 14303
rect 420 14269 433 14303
rect 373 14235 433 14269
rect 373 14201 386 14235
rect 420 14201 433 14235
rect 373 14167 433 14201
rect 373 14133 386 14167
rect 420 14133 433 14167
rect 373 14099 433 14133
rect 373 14065 386 14099
rect 420 14065 433 14099
rect 373 14031 433 14065
rect 373 13997 386 14031
rect 420 13997 433 14031
rect 373 13963 433 13997
rect 373 13929 386 13963
rect 420 13929 433 13963
rect 373 13895 433 13929
rect 373 13861 386 13895
rect 420 13861 433 13895
rect 373 13827 433 13861
rect 373 13793 386 13827
rect 420 13793 433 13827
rect 373 13759 433 13793
rect 373 13725 386 13759
rect 420 13725 433 13759
rect 373 13691 433 13725
rect 373 13657 386 13691
rect 420 13657 433 13691
rect 373 13623 433 13657
rect 373 13589 386 13623
rect 420 13589 433 13623
rect 373 13555 433 13589
rect 373 13521 386 13555
rect 420 13521 433 13555
rect 373 13487 433 13521
rect 3023 15548 3036 15582
rect 3070 15548 3083 15582
rect 3023 15514 3083 15548
rect 3023 15480 3036 15514
rect 3070 15480 3083 15514
rect 3023 15446 3083 15480
rect 3023 15412 3036 15446
rect 3070 15412 3083 15446
rect 3023 15378 3083 15412
rect 3023 15344 3036 15378
rect 3070 15344 3083 15378
rect 3023 15310 3083 15344
rect 3023 15276 3036 15310
rect 3070 15276 3083 15310
rect 3023 15242 3083 15276
rect 3023 15208 3036 15242
rect 3070 15208 3083 15242
rect 3023 15174 3083 15208
rect 3023 15140 3036 15174
rect 3070 15140 3083 15174
rect 3023 15106 3083 15140
rect 3023 15072 3036 15106
rect 3070 15072 3083 15106
rect 3023 15038 3083 15072
rect 3023 15004 3036 15038
rect 3070 15004 3083 15038
rect 3023 14970 3083 15004
rect 3023 14936 3036 14970
rect 3070 14936 3083 14970
rect 3023 14902 3083 14936
rect 3023 14868 3036 14902
rect 3070 14868 3083 14902
rect 3023 14834 3083 14868
rect 3023 14800 3036 14834
rect 3070 14800 3083 14834
rect 3023 14766 3083 14800
rect 3023 14732 3036 14766
rect 3070 14732 3083 14766
rect 3023 14698 3083 14732
rect 3023 14664 3036 14698
rect 3070 14664 3083 14698
rect 3023 14630 3083 14664
rect 3023 14596 3036 14630
rect 3070 14596 3083 14630
rect 3023 14562 3083 14596
rect 3023 14528 3036 14562
rect 3070 14528 3083 14562
rect 3023 14494 3083 14528
rect 3023 14460 3036 14494
rect 3070 14460 3083 14494
rect 3023 14426 3083 14460
rect 3023 14392 3036 14426
rect 3070 14392 3083 14426
rect 3023 14358 3083 14392
rect 3023 14324 3036 14358
rect 3070 14324 3083 14358
rect 3023 14290 3083 14324
rect 3023 14256 3036 14290
rect 3070 14256 3083 14290
rect 3023 14222 3083 14256
rect 3023 14188 3036 14222
rect 3070 14188 3083 14222
rect 3023 14154 3083 14188
rect 3023 14120 3036 14154
rect 3070 14120 3083 14154
rect 3023 14086 3083 14120
rect 3023 14052 3036 14086
rect 3070 14052 3083 14086
rect 3023 14018 3083 14052
rect 3023 13984 3036 14018
rect 3070 13984 3083 14018
rect 3023 13950 3083 13984
rect 3023 13916 3036 13950
rect 3070 13916 3083 13950
rect 3023 13882 3083 13916
rect 3023 13848 3036 13882
rect 3070 13848 3083 13882
rect 3023 13814 3083 13848
rect 3023 13780 3036 13814
rect 3070 13780 3083 13814
rect 3023 13746 3083 13780
rect 3023 13712 3036 13746
rect 3070 13712 3083 13746
rect 3023 13678 3083 13712
rect 3023 13644 3036 13678
rect 3070 13644 3083 13678
rect 3023 13610 3083 13644
rect 3023 13576 3036 13610
rect 3070 13576 3083 13610
rect 3023 13542 3083 13576
rect 373 13453 386 13487
rect 420 13453 433 13487
rect 373 13419 433 13453
rect 3023 13508 3036 13542
rect 3070 13508 3083 13542
rect 3023 13474 3083 13508
rect 373 13385 386 13419
rect 420 13385 433 13419
rect 373 13351 433 13385
rect 373 13317 386 13351
rect 420 13317 433 13351
rect 373 13283 433 13317
rect 373 13249 386 13283
rect 420 13249 433 13283
rect 373 13215 433 13249
rect 373 13181 386 13215
rect 420 13181 433 13215
rect 373 13147 433 13181
rect 373 13113 386 13147
rect 420 13113 433 13147
rect 373 13079 433 13113
rect 373 13045 386 13079
rect 420 13045 433 13079
rect 373 13011 433 13045
rect 373 12977 386 13011
rect 420 12977 433 13011
rect 373 12943 433 12977
rect 373 12909 386 12943
rect 420 12909 433 12943
rect 373 12875 433 12909
rect 373 12841 386 12875
rect 420 12841 433 12875
rect 373 12807 433 12841
rect 373 12773 386 12807
rect 420 12773 433 12807
rect 373 12739 433 12773
rect 373 12705 386 12739
rect 420 12705 433 12739
rect 373 12671 433 12705
rect 373 12637 386 12671
rect 420 12637 433 12671
rect 373 12603 433 12637
rect 373 12569 386 12603
rect 420 12569 433 12603
rect 373 12535 433 12569
rect 373 12501 386 12535
rect 420 12501 433 12535
rect 373 12467 433 12501
rect 373 12433 386 12467
rect 420 12433 433 12467
rect 373 12399 433 12433
rect 373 12365 386 12399
rect 420 12365 433 12399
rect 373 12331 433 12365
rect 373 12297 386 12331
rect 420 12297 433 12331
rect 373 12263 433 12297
rect 373 12229 386 12263
rect 420 12229 433 12263
rect 373 12195 433 12229
rect 373 12161 386 12195
rect 420 12161 433 12195
rect 373 12127 433 12161
rect 373 12093 386 12127
rect 420 12093 433 12127
rect 373 12059 433 12093
rect 373 12025 386 12059
rect 420 12025 433 12059
rect 373 11991 433 12025
rect 373 11957 386 11991
rect 420 11957 433 11991
rect 373 11923 433 11957
rect 373 11889 386 11923
rect 420 11889 433 11923
rect 373 11855 433 11889
rect 373 11821 386 11855
rect 420 11821 433 11855
rect 373 11787 433 11821
rect 373 11753 386 11787
rect 420 11753 433 11787
rect 373 11719 433 11753
rect 373 11685 386 11719
rect 420 11685 433 11719
rect 373 11651 433 11685
rect 373 11617 386 11651
rect 420 11617 433 11651
rect 373 11583 433 11617
rect 373 11549 386 11583
rect 420 11549 433 11583
rect 373 11515 433 11549
rect 373 11481 386 11515
rect 420 11481 433 11515
rect 373 11447 433 11481
rect 373 11413 386 11447
rect 420 11413 433 11447
rect 373 11379 433 11413
rect 3023 13440 3036 13474
rect 3070 13440 3083 13474
rect 3023 13406 3083 13440
rect 3023 13372 3036 13406
rect 3070 13372 3083 13406
rect 3023 13338 3083 13372
rect 3023 13304 3036 13338
rect 3070 13304 3083 13338
rect 3023 13270 3083 13304
rect 3023 13236 3036 13270
rect 3070 13236 3083 13270
rect 3023 13202 3083 13236
rect 3023 13168 3036 13202
rect 3070 13168 3083 13202
rect 3023 13134 3083 13168
rect 3023 13100 3036 13134
rect 3070 13100 3083 13134
rect 3023 13066 3083 13100
rect 3023 13032 3036 13066
rect 3070 13032 3083 13066
rect 3023 12998 3083 13032
rect 3023 12964 3036 12998
rect 3070 12964 3083 12998
rect 3023 12930 3083 12964
rect 3023 12896 3036 12930
rect 3070 12896 3083 12930
rect 3023 12862 3083 12896
rect 3023 12828 3036 12862
rect 3070 12828 3083 12862
rect 3023 12794 3083 12828
rect 3023 12760 3036 12794
rect 3070 12760 3083 12794
rect 3023 12726 3083 12760
rect 3023 12692 3036 12726
rect 3070 12692 3083 12726
rect 3023 12658 3083 12692
rect 3023 12624 3036 12658
rect 3070 12624 3083 12658
rect 3023 12590 3083 12624
rect 3023 12556 3036 12590
rect 3070 12556 3083 12590
rect 3023 12522 3083 12556
rect 3023 12488 3036 12522
rect 3070 12488 3083 12522
rect 3023 12454 3083 12488
rect 3023 12420 3036 12454
rect 3070 12420 3083 12454
rect 3023 12386 3083 12420
rect 3023 12352 3036 12386
rect 3070 12352 3083 12386
rect 3023 12318 3083 12352
rect 3023 12284 3036 12318
rect 3070 12284 3083 12318
rect 3023 12250 3083 12284
rect 3023 12216 3036 12250
rect 3070 12216 3083 12250
rect 3023 12182 3083 12216
rect 3023 12148 3036 12182
rect 3070 12148 3083 12182
rect 3023 12114 3083 12148
rect 3023 12080 3036 12114
rect 3070 12080 3083 12114
rect 3023 12046 3083 12080
rect 3023 12012 3036 12046
rect 3070 12012 3083 12046
rect 3023 11978 3083 12012
rect 3023 11944 3036 11978
rect 3070 11944 3083 11978
rect 3023 11910 3083 11944
rect 3023 11876 3036 11910
rect 3070 11876 3083 11910
rect 3023 11842 3083 11876
rect 3023 11808 3036 11842
rect 3070 11808 3083 11842
rect 3023 11774 3083 11808
rect 3023 11740 3036 11774
rect 3070 11740 3083 11774
rect 3023 11706 3083 11740
rect 3023 11672 3036 11706
rect 3070 11672 3083 11706
rect 3023 11638 3083 11672
rect 3023 11604 3036 11638
rect 3070 11604 3083 11638
rect 3023 11570 3083 11604
rect 3023 11536 3036 11570
rect 3070 11536 3083 11570
rect 3023 11502 3083 11536
rect 3023 11468 3036 11502
rect 3070 11468 3083 11502
rect 3023 11434 3083 11468
rect 3023 11400 3036 11434
rect 3070 11400 3083 11434
rect 373 11345 386 11379
rect 420 11345 433 11379
rect 373 11311 433 11345
rect 3023 11366 3083 11400
rect 3023 11332 3036 11366
rect 3070 11332 3083 11366
rect 373 11277 386 11311
rect 420 11277 433 11311
rect 373 11243 433 11277
rect 373 11209 386 11243
rect 420 11209 433 11243
rect 373 11175 433 11209
rect 373 11141 386 11175
rect 420 11141 433 11175
rect 373 11107 433 11141
rect 373 11073 386 11107
rect 420 11073 433 11107
rect 373 11039 433 11073
rect 373 11005 386 11039
rect 420 11005 433 11039
rect 373 10971 433 11005
rect 373 10937 386 10971
rect 420 10937 433 10971
rect 373 10903 433 10937
rect 373 10869 386 10903
rect 420 10869 433 10903
rect 373 10835 433 10869
rect 373 10801 386 10835
rect 420 10801 433 10835
rect 373 10767 433 10801
rect 373 10733 386 10767
rect 420 10733 433 10767
rect 373 10699 433 10733
rect 373 10665 386 10699
rect 420 10665 433 10699
rect 373 10631 433 10665
rect 373 10597 386 10631
rect 420 10597 433 10631
rect 373 10563 433 10597
rect 373 10529 386 10563
rect 420 10529 433 10563
rect 373 10495 433 10529
rect 373 10461 386 10495
rect 420 10461 433 10495
rect 373 10427 433 10461
rect 373 10393 386 10427
rect 420 10393 433 10427
rect 373 10359 433 10393
rect 373 10325 386 10359
rect 420 10325 433 10359
rect 373 10291 433 10325
rect 373 10257 386 10291
rect 420 10257 433 10291
rect 373 10223 433 10257
rect 373 10189 386 10223
rect 420 10189 433 10223
rect 373 10155 433 10189
rect 373 10121 386 10155
rect 420 10121 433 10155
rect 373 10087 433 10121
rect 373 10053 386 10087
rect 420 10053 433 10087
rect 373 10019 433 10053
rect 373 9985 386 10019
rect 420 9985 433 10019
rect 373 9951 433 9985
rect 373 9917 386 9951
rect 420 9917 433 9951
rect 373 9883 433 9917
rect 373 9849 386 9883
rect 420 9849 433 9883
rect 373 9815 433 9849
rect 373 9781 386 9815
rect 420 9781 433 9815
rect 373 9747 433 9781
rect 373 9713 386 9747
rect 420 9713 433 9747
rect 373 9679 433 9713
rect 373 9645 386 9679
rect 420 9645 433 9679
rect 373 9611 433 9645
rect 373 9577 386 9611
rect 420 9577 433 9611
rect 373 9543 433 9577
rect 373 9509 386 9543
rect 420 9509 433 9543
rect 373 9475 433 9509
rect 373 9441 386 9475
rect 420 9441 433 9475
rect 373 9407 433 9441
rect 373 9373 386 9407
rect 420 9373 433 9407
rect 373 9339 433 9373
rect 373 9305 386 9339
rect 420 9305 433 9339
rect 373 9271 433 9305
rect 373 9237 386 9271
rect 420 9237 433 9271
rect 3023 11298 3083 11332
rect 3023 11264 3036 11298
rect 3070 11264 3083 11298
rect 3023 11230 3083 11264
rect 3023 11196 3036 11230
rect 3070 11196 3083 11230
rect 3023 11162 3083 11196
rect 3023 11128 3036 11162
rect 3070 11128 3083 11162
rect 3023 11094 3083 11128
rect 3023 11060 3036 11094
rect 3070 11060 3083 11094
rect 3023 11026 3083 11060
rect 3023 10992 3036 11026
rect 3070 10992 3083 11026
rect 3023 10958 3083 10992
rect 3023 10924 3036 10958
rect 3070 10924 3083 10958
rect 3023 10890 3083 10924
rect 3023 10856 3036 10890
rect 3070 10856 3083 10890
rect 3023 10822 3083 10856
rect 3023 10788 3036 10822
rect 3070 10788 3083 10822
rect 3023 10754 3083 10788
rect 3023 10720 3036 10754
rect 3070 10720 3083 10754
rect 3023 10686 3083 10720
rect 3023 10652 3036 10686
rect 3070 10652 3083 10686
rect 3023 10618 3083 10652
rect 3023 10584 3036 10618
rect 3070 10584 3083 10618
rect 3023 10550 3083 10584
rect 3023 10516 3036 10550
rect 3070 10516 3083 10550
rect 3023 10482 3083 10516
rect 3023 10448 3036 10482
rect 3070 10448 3083 10482
rect 3023 10414 3083 10448
rect 3023 10380 3036 10414
rect 3070 10380 3083 10414
rect 3023 10346 3083 10380
rect 3023 10312 3036 10346
rect 3070 10312 3083 10346
rect 3023 10278 3083 10312
rect 3023 10244 3036 10278
rect 3070 10244 3083 10278
rect 3023 10210 3083 10244
rect 3023 10176 3036 10210
rect 3070 10176 3083 10210
rect 3023 10142 3083 10176
rect 3023 10108 3036 10142
rect 3070 10108 3083 10142
rect 3023 10074 3083 10108
rect 3023 10040 3036 10074
rect 3070 10040 3083 10074
rect 3023 10006 3083 10040
rect 3023 9972 3036 10006
rect 3070 9972 3083 10006
rect 3023 9938 3083 9972
rect 3023 9904 3036 9938
rect 3070 9904 3083 9938
rect 3023 9870 3083 9904
rect 3023 9836 3036 9870
rect 3070 9836 3083 9870
rect 3023 9802 3083 9836
rect 3023 9768 3036 9802
rect 3070 9768 3083 9802
rect 3023 9734 3083 9768
rect 3023 9700 3036 9734
rect 3070 9700 3083 9734
rect 3023 9666 3083 9700
rect 3023 9632 3036 9666
rect 3070 9632 3083 9666
rect 3023 9598 3083 9632
rect 3023 9564 3036 9598
rect 3070 9564 3083 9598
rect 3023 9530 3083 9564
rect 3023 9496 3036 9530
rect 3070 9496 3083 9530
rect 3023 9462 3083 9496
rect 3023 9428 3036 9462
rect 3070 9428 3083 9462
rect 3023 9394 3083 9428
rect 3023 9360 3036 9394
rect 3070 9360 3083 9394
rect 3023 9326 3083 9360
rect 3023 9292 3036 9326
rect 3070 9292 3083 9326
rect 3023 9258 3083 9292
rect 373 9203 433 9237
rect 373 9169 386 9203
rect 420 9169 433 9203
rect 3023 9224 3036 9258
rect 3070 9224 3083 9258
rect 3023 9190 3083 9224
rect 373 9135 433 9169
rect 373 9101 386 9135
rect 420 9101 433 9135
rect 373 9067 433 9101
rect 373 9033 386 9067
rect 420 9033 433 9067
rect 373 8999 433 9033
rect 373 8965 386 8999
rect 420 8965 433 8999
rect 373 8931 433 8965
rect 373 8897 386 8931
rect 420 8897 433 8931
rect 373 8863 433 8897
rect 373 8829 386 8863
rect 420 8829 433 8863
rect 373 8795 433 8829
rect 373 8761 386 8795
rect 420 8761 433 8795
rect 373 8727 433 8761
rect 373 8693 386 8727
rect 420 8693 433 8727
rect 373 8659 433 8693
rect 373 8625 386 8659
rect 420 8625 433 8659
rect 373 8591 433 8625
rect 373 8557 386 8591
rect 420 8557 433 8591
rect 373 8523 433 8557
rect 373 8489 386 8523
rect 420 8489 433 8523
rect 373 8455 433 8489
rect 373 8421 386 8455
rect 420 8421 433 8455
rect 373 8387 433 8421
rect 373 8353 386 8387
rect 420 8353 433 8387
rect 373 8319 433 8353
rect 373 8285 386 8319
rect 420 8285 433 8319
rect 373 8251 433 8285
rect 373 8217 386 8251
rect 420 8217 433 8251
rect 373 8183 433 8217
rect 373 8149 386 8183
rect 420 8149 433 8183
rect 373 8115 433 8149
rect 373 8081 386 8115
rect 420 8081 433 8115
rect 373 8047 433 8081
rect 373 8013 386 8047
rect 420 8013 433 8047
rect 373 7979 433 8013
rect 373 7945 386 7979
rect 420 7945 433 7979
rect 373 7911 433 7945
rect 373 7877 386 7911
rect 420 7877 433 7911
rect 373 7843 433 7877
rect 373 7809 386 7843
rect 420 7809 433 7843
rect 373 7775 433 7809
rect 373 7741 386 7775
rect 420 7741 433 7775
rect 373 7707 433 7741
rect 373 7673 386 7707
rect 420 7673 433 7707
rect 373 7639 433 7673
rect 373 7605 386 7639
rect 420 7605 433 7639
rect 373 7571 433 7605
rect 373 7537 386 7571
rect 420 7537 433 7571
rect 373 7503 433 7537
rect 373 7469 386 7503
rect 420 7469 433 7503
rect 373 7435 433 7469
rect 373 7401 386 7435
rect 420 7401 433 7435
rect 373 7367 433 7401
rect 373 7333 386 7367
rect 420 7333 433 7367
rect 373 7299 433 7333
rect 373 7265 386 7299
rect 420 7265 433 7299
rect 373 7231 433 7265
rect 373 7197 386 7231
rect 420 7197 433 7231
rect 373 7163 433 7197
rect 373 7129 386 7163
rect 420 7129 433 7163
rect 373 7095 433 7129
rect 3023 9156 3036 9190
rect 3070 9156 3083 9190
rect 3023 9122 3083 9156
rect 3023 9088 3036 9122
rect 3070 9088 3083 9122
rect 3023 9054 3083 9088
rect 3023 9020 3036 9054
rect 3070 9020 3083 9054
rect 3023 8986 3083 9020
rect 3023 8952 3036 8986
rect 3070 8952 3083 8986
rect 3023 8918 3083 8952
rect 3023 8884 3036 8918
rect 3070 8884 3083 8918
rect 3023 8850 3083 8884
rect 3023 8816 3036 8850
rect 3070 8816 3083 8850
rect 3023 8782 3083 8816
rect 3023 8748 3036 8782
rect 3070 8748 3083 8782
rect 3023 8714 3083 8748
rect 3023 8680 3036 8714
rect 3070 8680 3083 8714
rect 3023 8646 3083 8680
rect 3023 8612 3036 8646
rect 3070 8612 3083 8646
rect 3023 8578 3083 8612
rect 3023 8544 3036 8578
rect 3070 8544 3083 8578
rect 3023 8510 3083 8544
rect 3023 8476 3036 8510
rect 3070 8476 3083 8510
rect 3023 8442 3083 8476
rect 3023 8408 3036 8442
rect 3070 8408 3083 8442
rect 3023 8374 3083 8408
rect 3023 8340 3036 8374
rect 3070 8340 3083 8374
rect 3023 8306 3083 8340
rect 3023 8272 3036 8306
rect 3070 8272 3083 8306
rect 3023 8238 3083 8272
rect 3023 8204 3036 8238
rect 3070 8204 3083 8238
rect 3023 8170 3083 8204
rect 3023 8136 3036 8170
rect 3070 8136 3083 8170
rect 3023 8102 3083 8136
rect 3023 8068 3036 8102
rect 3070 8068 3083 8102
rect 3023 8034 3083 8068
rect 3023 8000 3036 8034
rect 3070 8000 3083 8034
rect 3023 7966 3083 8000
rect 3023 7932 3036 7966
rect 3070 7932 3083 7966
rect 3023 7898 3083 7932
rect 3023 7864 3036 7898
rect 3070 7864 3083 7898
rect 3023 7830 3083 7864
rect 3023 7796 3036 7830
rect 3070 7796 3083 7830
rect 3023 7762 3083 7796
rect 3023 7728 3036 7762
rect 3070 7728 3083 7762
rect 3023 7694 3083 7728
rect 3023 7660 3036 7694
rect 3070 7660 3083 7694
rect 3023 7626 3083 7660
rect 3023 7592 3036 7626
rect 3070 7592 3083 7626
rect 3023 7558 3083 7592
rect 3023 7524 3036 7558
rect 3070 7524 3083 7558
rect 3023 7490 3083 7524
rect 3023 7456 3036 7490
rect 3070 7456 3083 7490
rect 3023 7422 3083 7456
rect 3023 7388 3036 7422
rect 3070 7388 3083 7422
rect 3023 7354 3083 7388
rect 3023 7320 3036 7354
rect 3070 7320 3083 7354
rect 3023 7286 3083 7320
rect 3023 7252 3036 7286
rect 3070 7252 3083 7286
rect 3023 7218 3083 7252
rect 3023 7184 3036 7218
rect 3070 7184 3083 7218
rect 3023 7150 3083 7184
rect 373 7061 386 7095
rect 420 7061 433 7095
rect 373 7027 433 7061
rect 3023 7116 3036 7150
rect 3070 7116 3083 7150
rect 3023 7082 3083 7116
rect 373 6993 386 7027
rect 420 6993 433 7027
rect 373 6959 433 6993
rect 373 6925 386 6959
rect 420 6925 433 6959
rect 373 6891 433 6925
rect 373 6857 386 6891
rect 420 6857 433 6891
rect 373 6823 433 6857
rect 373 6789 386 6823
rect 420 6789 433 6823
rect 373 6755 433 6789
rect 373 6721 386 6755
rect 420 6721 433 6755
rect 373 6687 433 6721
rect 373 6653 386 6687
rect 420 6653 433 6687
rect 373 6619 433 6653
rect 373 6585 386 6619
rect 420 6585 433 6619
rect 373 6551 433 6585
rect 373 6517 386 6551
rect 420 6517 433 6551
rect 373 6483 433 6517
rect 373 6449 386 6483
rect 420 6449 433 6483
rect 373 6415 433 6449
rect 373 6381 386 6415
rect 420 6381 433 6415
rect 373 6347 433 6381
rect 373 6313 386 6347
rect 420 6313 433 6347
rect 373 6279 433 6313
rect 373 6245 386 6279
rect 420 6245 433 6279
rect 373 6211 433 6245
rect 373 6177 386 6211
rect 420 6177 433 6211
rect 373 6143 433 6177
rect 373 6109 386 6143
rect 420 6109 433 6143
rect 373 6075 433 6109
rect 373 6041 386 6075
rect 420 6041 433 6075
rect 373 6007 433 6041
rect 373 5973 386 6007
rect 420 5973 433 6007
rect 373 5939 433 5973
rect 373 5905 386 5939
rect 420 5905 433 5939
rect 373 5871 433 5905
rect 373 5837 386 5871
rect 420 5837 433 5871
rect 373 5803 433 5837
rect 373 5769 386 5803
rect 420 5769 433 5803
rect 373 5735 433 5769
rect 373 5701 386 5735
rect 420 5701 433 5735
rect 373 5667 433 5701
rect 373 5633 386 5667
rect 420 5633 433 5667
rect 373 5599 433 5633
rect 373 5565 386 5599
rect 420 5565 433 5599
rect 373 5531 433 5565
rect 373 5497 386 5531
rect 420 5497 433 5531
rect 373 5463 433 5497
rect 373 5429 386 5463
rect 420 5429 433 5463
rect 373 5395 433 5429
rect 373 5361 386 5395
rect 420 5361 433 5395
rect 373 5327 433 5361
rect 373 5293 386 5327
rect 420 5293 433 5327
rect 373 5259 433 5293
rect 373 5225 386 5259
rect 420 5225 433 5259
rect 373 5191 433 5225
rect 373 5157 386 5191
rect 420 5157 433 5191
rect 373 5123 433 5157
rect 373 5089 386 5123
rect 420 5089 433 5123
rect 373 5055 433 5089
rect 373 5021 386 5055
rect 420 5021 433 5055
rect 373 4987 433 5021
rect 3023 7048 3036 7082
rect 3070 7048 3083 7082
rect 3023 7014 3083 7048
rect 3023 6980 3036 7014
rect 3070 6980 3083 7014
rect 3023 6946 3083 6980
rect 3023 6912 3036 6946
rect 3070 6912 3083 6946
rect 3023 6878 3083 6912
rect 3023 6844 3036 6878
rect 3070 6844 3083 6878
rect 3023 6810 3083 6844
rect 3023 6776 3036 6810
rect 3070 6776 3083 6810
rect 3023 6742 3083 6776
rect 3023 6708 3036 6742
rect 3070 6708 3083 6742
rect 3023 6674 3083 6708
rect 3023 6640 3036 6674
rect 3070 6640 3083 6674
rect 3023 6606 3083 6640
rect 3023 6572 3036 6606
rect 3070 6572 3083 6606
rect 3023 6538 3083 6572
rect 3023 6504 3036 6538
rect 3070 6504 3083 6538
rect 3023 6470 3083 6504
rect 3023 6436 3036 6470
rect 3070 6436 3083 6470
rect 3023 6402 3083 6436
rect 3023 6368 3036 6402
rect 3070 6368 3083 6402
rect 3023 6334 3083 6368
rect 3023 6300 3036 6334
rect 3070 6300 3083 6334
rect 3023 6266 3083 6300
rect 3023 6232 3036 6266
rect 3070 6232 3083 6266
rect 3023 6198 3083 6232
rect 3023 6164 3036 6198
rect 3070 6164 3083 6198
rect 3023 6130 3083 6164
rect 3023 6096 3036 6130
rect 3070 6096 3083 6130
rect 3023 6062 3083 6096
rect 3023 6028 3036 6062
rect 3070 6028 3083 6062
rect 3023 5994 3083 6028
rect 3023 5960 3036 5994
rect 3070 5960 3083 5994
rect 3023 5926 3083 5960
rect 3023 5892 3036 5926
rect 3070 5892 3083 5926
rect 3023 5858 3083 5892
rect 3023 5824 3036 5858
rect 3070 5824 3083 5858
rect 3023 5790 3083 5824
rect 3023 5756 3036 5790
rect 3070 5756 3083 5790
rect 3023 5722 3083 5756
rect 3023 5688 3036 5722
rect 3070 5688 3083 5722
rect 3023 5654 3083 5688
rect 3023 5620 3036 5654
rect 3070 5620 3083 5654
rect 3023 5586 3083 5620
rect 3023 5552 3036 5586
rect 3070 5552 3083 5586
rect 3023 5518 3083 5552
rect 3023 5484 3036 5518
rect 3070 5484 3083 5518
rect 3023 5450 3083 5484
rect 3023 5416 3036 5450
rect 3070 5416 3083 5450
rect 3023 5382 3083 5416
rect 3023 5348 3036 5382
rect 3070 5348 3083 5382
rect 3023 5314 3083 5348
rect 3023 5280 3036 5314
rect 3070 5280 3083 5314
rect 3023 5246 3083 5280
rect 3023 5212 3036 5246
rect 3070 5212 3083 5246
rect 3023 5178 3083 5212
rect 3023 5144 3036 5178
rect 3070 5144 3083 5178
rect 3023 5110 3083 5144
rect 3023 5076 3036 5110
rect 3070 5076 3083 5110
rect 3023 5042 3083 5076
rect 3023 5008 3036 5042
rect 3070 5008 3083 5042
rect 373 4953 386 4987
rect 420 4953 433 4987
rect 373 4919 433 4953
rect 3023 4974 3083 5008
rect 3023 4940 3036 4974
rect 3070 4940 3083 4974
rect 373 4885 386 4919
rect 420 4885 433 4919
rect 373 4851 433 4885
rect 373 4817 386 4851
rect 420 4817 433 4851
rect 373 4783 433 4817
rect 373 4749 386 4783
rect 420 4749 433 4783
rect 373 4715 433 4749
rect 373 4681 386 4715
rect 420 4681 433 4715
rect 373 4647 433 4681
rect 373 4613 386 4647
rect 420 4613 433 4647
rect 373 4579 433 4613
rect 373 4545 386 4579
rect 420 4545 433 4579
rect 373 4511 433 4545
rect 373 4477 386 4511
rect 420 4477 433 4511
rect 373 4443 433 4477
rect 373 4409 386 4443
rect 420 4409 433 4443
rect 373 4375 433 4409
rect 373 4341 386 4375
rect 420 4341 433 4375
rect 373 4307 433 4341
rect 373 4273 386 4307
rect 420 4273 433 4307
rect 373 4239 433 4273
rect 373 4205 386 4239
rect 420 4205 433 4239
rect 373 4171 433 4205
rect 373 4137 386 4171
rect 420 4137 433 4171
rect 373 4103 433 4137
rect 373 4069 386 4103
rect 420 4069 433 4103
rect 373 4035 433 4069
rect 373 4001 386 4035
rect 420 4001 433 4035
rect 373 3967 433 4001
rect 373 3933 386 3967
rect 420 3933 433 3967
rect 373 3899 433 3933
rect 373 3865 386 3899
rect 420 3865 433 3899
rect 373 3831 433 3865
rect 373 3797 386 3831
rect 420 3797 433 3831
rect 373 3763 433 3797
rect 373 3729 386 3763
rect 420 3729 433 3763
rect 373 3695 433 3729
rect 373 3661 386 3695
rect 420 3661 433 3695
rect 373 3627 433 3661
rect 373 3593 386 3627
rect 420 3593 433 3627
rect 373 3559 433 3593
rect 373 3525 386 3559
rect 420 3525 433 3559
rect 373 3491 433 3525
rect 373 3457 386 3491
rect 420 3457 433 3491
rect 373 3423 433 3457
rect 373 3389 386 3423
rect 420 3389 433 3423
rect 373 3355 433 3389
rect 373 3321 386 3355
rect 420 3321 433 3355
rect 373 3287 433 3321
rect 373 3253 386 3287
rect 420 3253 433 3287
rect 373 3219 433 3253
rect 373 3185 386 3219
rect 420 3185 433 3219
rect 373 3151 433 3185
rect 373 3117 386 3151
rect 420 3117 433 3151
rect 373 3083 433 3117
rect 373 3049 386 3083
rect 420 3049 433 3083
rect 373 3015 433 3049
rect 373 2981 386 3015
rect 420 2981 433 3015
rect 373 2947 433 2981
rect 373 2913 386 2947
rect 420 2913 433 2947
rect 373 2879 433 2913
rect 373 2845 386 2879
rect 420 2845 433 2879
rect 3023 4906 3083 4940
rect 3023 4872 3036 4906
rect 3070 4872 3083 4906
rect 3023 4838 3083 4872
rect 3023 4804 3036 4838
rect 3070 4804 3083 4838
rect 3023 4770 3083 4804
rect 3023 4736 3036 4770
rect 3070 4736 3083 4770
rect 3023 4702 3083 4736
rect 3023 4668 3036 4702
rect 3070 4668 3083 4702
rect 3023 4634 3083 4668
rect 3023 4600 3036 4634
rect 3070 4600 3083 4634
rect 3023 4566 3083 4600
rect 3023 4532 3036 4566
rect 3070 4532 3083 4566
rect 3023 4498 3083 4532
rect 3023 4464 3036 4498
rect 3070 4464 3083 4498
rect 3023 4430 3083 4464
rect 3023 4396 3036 4430
rect 3070 4396 3083 4430
rect 3023 4362 3083 4396
rect 3023 4328 3036 4362
rect 3070 4328 3083 4362
rect 3023 4294 3083 4328
rect 3023 4260 3036 4294
rect 3070 4260 3083 4294
rect 3023 4226 3083 4260
rect 3023 4192 3036 4226
rect 3070 4192 3083 4226
rect 3023 4158 3083 4192
rect 3023 4124 3036 4158
rect 3070 4124 3083 4158
rect 3023 4090 3083 4124
rect 3023 4056 3036 4090
rect 3070 4056 3083 4090
rect 3023 4022 3083 4056
rect 3023 3988 3036 4022
rect 3070 3988 3083 4022
rect 3023 3954 3083 3988
rect 3023 3920 3036 3954
rect 3070 3920 3083 3954
rect 3023 3886 3083 3920
rect 3023 3852 3036 3886
rect 3070 3852 3083 3886
rect 3023 3818 3083 3852
rect 3023 3784 3036 3818
rect 3070 3784 3083 3818
rect 3023 3750 3083 3784
rect 3023 3716 3036 3750
rect 3070 3716 3083 3750
rect 3023 3682 3083 3716
rect 3023 3648 3036 3682
rect 3070 3648 3083 3682
rect 3023 3614 3083 3648
rect 3023 3580 3036 3614
rect 3070 3580 3083 3614
rect 3023 3546 3083 3580
rect 3023 3512 3036 3546
rect 3070 3512 3083 3546
rect 3023 3478 3083 3512
rect 3023 3444 3036 3478
rect 3070 3444 3083 3478
rect 3023 3410 3083 3444
rect 3023 3376 3036 3410
rect 3070 3376 3083 3410
rect 3023 3342 3083 3376
rect 3023 3308 3036 3342
rect 3070 3308 3083 3342
rect 3023 3274 3083 3308
rect 3023 3240 3036 3274
rect 3070 3240 3083 3274
rect 3023 3206 3083 3240
rect 3023 3172 3036 3206
rect 3070 3172 3083 3206
rect 3023 3138 3083 3172
rect 3023 3104 3036 3138
rect 3070 3104 3083 3138
rect 3023 3070 3083 3104
rect 3023 3036 3036 3070
rect 3070 3036 3083 3070
rect 3023 3002 3083 3036
rect 3023 2968 3036 3002
rect 3070 2968 3083 3002
rect 3023 2934 3083 2968
rect 3023 2900 3036 2934
rect 3070 2900 3083 2934
rect 3023 2866 3083 2900
rect 373 2811 433 2845
rect 373 2777 386 2811
rect 420 2777 433 2811
rect 3023 2832 3036 2866
rect 3070 2832 3083 2866
rect 3023 2798 3083 2832
rect 373 2743 433 2777
rect 373 2709 386 2743
rect 420 2709 433 2743
rect 373 2675 433 2709
rect 373 2641 386 2675
rect 420 2641 433 2675
rect 373 2607 433 2641
rect 373 2573 386 2607
rect 420 2573 433 2607
rect 373 2539 433 2573
rect 373 2505 386 2539
rect 420 2505 433 2539
rect 373 2471 433 2505
rect 373 2437 386 2471
rect 420 2437 433 2471
rect 373 2403 433 2437
rect 373 2369 386 2403
rect 420 2369 433 2403
rect 373 2335 433 2369
rect 373 2301 386 2335
rect 420 2301 433 2335
rect 373 2267 433 2301
rect 373 2233 386 2267
rect 420 2233 433 2267
rect 373 2199 433 2233
rect 373 2165 386 2199
rect 420 2165 433 2199
rect 373 2131 433 2165
rect 373 2097 386 2131
rect 420 2097 433 2131
rect 373 2063 433 2097
rect 373 2029 386 2063
rect 420 2029 433 2063
rect 373 1995 433 2029
rect 373 1961 386 1995
rect 420 1961 433 1995
rect 373 1927 433 1961
rect 373 1893 386 1927
rect 420 1893 433 1927
rect 373 1859 433 1893
rect 373 1825 386 1859
rect 420 1825 433 1859
rect 373 1791 433 1825
rect 373 1757 386 1791
rect 420 1757 433 1791
rect 373 1723 433 1757
rect 373 1689 386 1723
rect 420 1689 433 1723
rect 373 1655 433 1689
rect 373 1621 386 1655
rect 420 1621 433 1655
rect 373 1587 433 1621
rect 373 1553 386 1587
rect 420 1553 433 1587
rect 373 1519 433 1553
rect 373 1485 386 1519
rect 420 1485 433 1519
rect 373 1451 433 1485
rect 373 1417 386 1451
rect 420 1417 433 1451
rect 373 1383 433 1417
rect 373 1349 386 1383
rect 420 1349 433 1383
rect 373 1315 433 1349
rect 373 1281 386 1315
rect 420 1281 433 1315
rect 373 1247 433 1281
rect 373 1213 386 1247
rect 420 1213 433 1247
rect 373 1179 433 1213
rect 373 1145 386 1179
rect 420 1145 433 1179
rect 373 1111 433 1145
rect 373 1077 386 1111
rect 420 1077 433 1111
rect 373 1043 433 1077
rect 373 1009 386 1043
rect 420 1009 433 1043
rect 373 975 433 1009
rect 373 941 386 975
rect 420 941 433 975
rect 373 907 433 941
rect 373 873 386 907
rect 420 873 433 907
rect 373 839 433 873
rect 373 805 386 839
rect 420 805 433 839
rect 373 771 433 805
rect 373 737 386 771
rect 420 737 433 771
rect 373 703 433 737
rect 3023 2764 3036 2798
rect 3070 2764 3083 2798
rect 3023 2730 3083 2764
rect 3023 2696 3036 2730
rect 3070 2696 3083 2730
rect 3023 2662 3083 2696
rect 3023 2628 3036 2662
rect 3070 2628 3083 2662
rect 3023 2594 3083 2628
rect 3023 2560 3036 2594
rect 3070 2560 3083 2594
rect 3023 2526 3083 2560
rect 3023 2492 3036 2526
rect 3070 2492 3083 2526
rect 3023 2458 3083 2492
rect 3023 2424 3036 2458
rect 3070 2424 3083 2458
rect 3023 2390 3083 2424
rect 3023 2356 3036 2390
rect 3070 2356 3083 2390
rect 3023 2322 3083 2356
rect 3023 2288 3036 2322
rect 3070 2288 3083 2322
rect 3023 2254 3083 2288
rect 3023 2220 3036 2254
rect 3070 2220 3083 2254
rect 3023 2186 3083 2220
rect 3023 2152 3036 2186
rect 3070 2152 3083 2186
rect 3023 2118 3083 2152
rect 3023 2084 3036 2118
rect 3070 2084 3083 2118
rect 3023 2050 3083 2084
rect 3023 2016 3036 2050
rect 3070 2016 3083 2050
rect 3023 1982 3083 2016
rect 3023 1948 3036 1982
rect 3070 1948 3083 1982
rect 3023 1914 3083 1948
rect 3023 1880 3036 1914
rect 3070 1880 3083 1914
rect 3023 1846 3083 1880
rect 3023 1812 3036 1846
rect 3070 1812 3083 1846
rect 3023 1778 3083 1812
rect 3023 1744 3036 1778
rect 3070 1744 3083 1778
rect 3023 1710 3083 1744
rect 3023 1676 3036 1710
rect 3070 1676 3083 1710
rect 3023 1642 3083 1676
rect 3023 1608 3036 1642
rect 3070 1608 3083 1642
rect 3023 1574 3083 1608
rect 3023 1540 3036 1574
rect 3070 1540 3083 1574
rect 3023 1506 3083 1540
rect 3023 1472 3036 1506
rect 3070 1472 3083 1506
rect 3023 1438 3083 1472
rect 3023 1404 3036 1438
rect 3070 1404 3083 1438
rect 3023 1370 3083 1404
rect 3023 1336 3036 1370
rect 3070 1336 3083 1370
rect 3023 1302 3083 1336
rect 3023 1268 3036 1302
rect 3070 1268 3083 1302
rect 3023 1234 3083 1268
rect 3023 1200 3036 1234
rect 3070 1200 3083 1234
rect 3023 1166 3083 1200
rect 3023 1132 3036 1166
rect 3070 1132 3083 1166
rect 3023 1098 3083 1132
rect 3023 1064 3036 1098
rect 3070 1064 3083 1098
rect 3023 1030 3083 1064
rect 3023 996 3036 1030
rect 3070 996 3083 1030
rect 3023 962 3083 996
rect 3023 928 3036 962
rect 3070 928 3083 962
rect 3023 894 3083 928
rect 3023 860 3036 894
rect 3070 860 3083 894
rect 3023 826 3083 860
rect 3023 792 3036 826
rect 3070 792 3083 826
rect 3023 758 3083 792
rect 373 669 386 703
rect 420 669 433 703
rect 373 580 433 669
rect 3023 724 3036 758
rect 3070 724 3083 758
rect 3023 690 3083 724
rect 3023 656 3036 690
rect 3070 656 3083 690
rect 3023 622 3083 656
rect 3023 588 3036 622
rect 3070 588 3083 622
rect 3023 580 3083 588
rect 373 567 3083 580
rect 373 533 441 567
rect 475 533 509 567
rect 543 533 577 567
rect 611 533 645 567
rect 679 533 713 567
rect 747 533 781 567
rect 815 533 849 567
rect 883 533 917 567
rect 951 533 985 567
rect 1019 533 1053 567
rect 1087 533 1121 567
rect 1155 533 1189 567
rect 1223 533 1257 567
rect 1291 533 1325 567
rect 1359 533 1393 567
rect 1427 533 1461 567
rect 1495 533 1529 567
rect 1563 533 1597 567
rect 1631 533 1665 567
rect 1699 533 1733 567
rect 1767 533 1801 567
rect 1835 533 1869 567
rect 1903 533 1937 567
rect 1971 533 2005 567
rect 2039 533 2073 567
rect 2107 533 2141 567
rect 2175 533 2209 567
rect 2243 533 2277 567
rect 2311 533 2345 567
rect 2379 533 2413 567
rect 2447 533 2481 567
rect 2515 533 2549 567
rect 2583 533 2617 567
rect 2651 533 2685 567
rect 2719 533 2753 567
rect 2787 533 2821 567
rect 2855 533 2889 567
rect 2923 533 2957 567
rect 2991 533 3083 567
rect 373 520 3083 533
<< mvnsubdiff >>
rect 126 39840 236 39874
rect 270 39840 304 39874
rect 338 39840 372 39874
rect 406 39840 440 39874
rect 474 39840 508 39874
rect 542 39840 576 39874
rect 610 39840 644 39874
rect 678 39840 712 39874
rect 746 39840 780 39874
rect 814 39840 848 39874
rect 882 39840 916 39874
rect 950 39840 984 39874
rect 1018 39840 1052 39874
rect 1086 39840 1120 39874
rect 1154 39840 1188 39874
rect 1222 39840 1256 39874
rect 1290 39840 1324 39874
rect 1358 39840 1392 39874
rect 1426 39840 1460 39874
rect 1494 39840 1528 39874
rect 1562 39840 1596 39874
rect 1630 39840 1664 39874
rect 1698 39840 1732 39874
rect 1766 39840 1800 39874
rect 1834 39840 1868 39874
rect 1902 39840 1936 39874
rect 1970 39840 2004 39874
rect 2038 39840 2072 39874
rect 2106 39840 2140 39874
rect 2174 39840 2208 39874
rect 2242 39840 2276 39874
rect 2310 39840 2344 39874
rect 2378 39840 2412 39874
rect 2446 39840 2480 39874
rect 2514 39840 2548 39874
rect 2582 39840 2616 39874
rect 2650 39840 2684 39874
rect 2718 39840 2752 39874
rect 2786 39840 2820 39874
rect 2854 39840 2888 39874
rect 2922 39840 2956 39874
rect 2990 39840 3024 39874
rect 3058 39840 3092 39874
rect 3126 39840 3160 39874
rect 3194 39840 3228 39874
rect 3262 39840 3330 39874
rect 126 39806 160 39840
rect 126 39738 160 39772
rect 126 39670 160 39704
rect 126 39602 160 39636
rect 126 39534 160 39568
rect 126 39466 160 39500
rect 126 39398 160 39432
rect 126 39330 160 39364
rect 126 39262 160 39296
rect 126 39194 160 39228
rect 3296 39804 3330 39840
rect 3296 39736 3330 39770
rect 3296 39668 3330 39702
rect 3296 39600 3330 39634
rect 3296 39532 3330 39566
rect 3296 39464 3330 39498
rect 3296 39396 3330 39430
rect 3296 39328 3330 39362
rect 3296 39260 3330 39294
rect 3296 39192 3330 39226
rect 126 39126 160 39160
rect 126 39058 160 39092
rect 126 38990 160 39024
rect 126 38922 160 38956
rect 126 38854 160 38888
rect 126 38786 160 38820
rect 126 38718 160 38752
rect 126 38650 160 38684
rect 126 38582 160 38616
rect 126 38514 160 38548
rect 126 38446 160 38480
rect 126 38378 160 38412
rect 126 38310 160 38344
rect 126 38242 160 38276
rect 126 38174 160 38208
rect 126 38106 160 38140
rect 126 38038 160 38072
rect 126 37970 160 38004
rect 126 37902 160 37936
rect 126 37834 160 37868
rect 126 37766 160 37800
rect 126 37698 160 37732
rect 126 37630 160 37664
rect 126 37562 160 37596
rect 126 37494 160 37528
rect 126 37426 160 37460
rect 126 37358 160 37392
rect 126 37290 160 37324
rect 126 37222 160 37256
rect 126 37154 160 37188
rect 126 37086 160 37120
rect 126 37018 160 37052
rect 126 36950 160 36984
rect 126 36882 160 36916
rect 126 36814 160 36848
rect 126 36746 160 36780
rect 126 36678 160 36712
rect 126 36610 160 36644
rect 126 36542 160 36576
rect 126 36474 160 36508
rect 126 36406 160 36440
rect 126 36338 160 36372
rect 126 36270 160 36304
rect 126 36202 160 36236
rect 126 36134 160 36168
rect 126 36066 160 36100
rect 126 35998 160 36032
rect 126 35930 160 35964
rect 126 35862 160 35896
rect 126 35794 160 35828
rect 126 35726 160 35760
rect 126 35658 160 35692
rect 126 35590 160 35624
rect 126 35522 160 35556
rect 126 35454 160 35488
rect 126 35386 160 35420
rect 126 35318 160 35352
rect 126 35250 160 35284
rect 126 35182 160 35216
rect 126 35114 160 35148
rect 126 35046 160 35080
rect 126 34978 160 35012
rect 126 34910 160 34944
rect 126 34842 160 34876
rect 126 34774 160 34808
rect 126 34706 160 34740
rect 126 34638 160 34672
rect 126 34570 160 34604
rect 126 34502 160 34536
rect 126 34434 160 34468
rect 126 34366 160 34400
rect 126 34298 160 34332
rect 126 34230 160 34264
rect 126 34162 160 34196
rect 126 34094 160 34128
rect 126 34026 160 34060
rect 126 33958 160 33992
rect 126 33890 160 33924
rect 126 33822 160 33856
rect 126 33754 160 33788
rect 126 33686 160 33720
rect 126 33618 160 33652
rect 126 33550 160 33584
rect 126 33482 160 33516
rect 126 33414 160 33448
rect 126 33346 160 33380
rect 126 33278 160 33312
rect 126 33210 160 33244
rect 126 33142 160 33176
rect 126 33074 160 33108
rect 126 33006 160 33040
rect 126 32938 160 32972
rect 126 32870 160 32904
rect 126 32802 160 32836
rect 126 32734 160 32768
rect 126 32666 160 32700
rect 126 32598 160 32632
rect 126 32530 160 32564
rect 126 32462 160 32496
rect 126 32394 160 32428
rect 126 32326 160 32360
rect 126 32258 160 32292
rect 126 32190 160 32224
rect 126 32122 160 32156
rect 126 32054 160 32088
rect 126 31986 160 32020
rect 126 31918 160 31952
rect 126 31850 160 31884
rect 126 31782 160 31816
rect 126 31714 160 31748
rect 126 31646 160 31680
rect 126 31578 160 31612
rect 126 31510 160 31544
rect 126 31442 160 31476
rect 126 31374 160 31408
rect 126 31306 160 31340
rect 126 31238 160 31272
rect 126 31170 160 31204
rect 126 31102 160 31136
rect 126 31034 160 31068
rect 126 30966 160 31000
rect 126 30898 160 30932
rect 126 30830 160 30864
rect 126 30762 160 30796
rect 126 30694 160 30728
rect 126 30626 160 30660
rect 126 30558 160 30592
rect 126 30490 160 30524
rect 126 30422 160 30456
rect 126 30354 160 30388
rect 126 30286 160 30320
rect 126 30218 160 30252
rect 126 30150 160 30184
rect 126 30082 160 30116
rect 126 30014 160 30048
rect 126 29946 160 29980
rect 126 29878 160 29912
rect 126 29810 160 29844
rect 126 29742 160 29776
rect 126 29674 160 29708
rect 126 29606 160 29640
rect 126 29538 160 29572
rect 126 29470 160 29504
rect 126 29402 160 29436
rect 126 29334 160 29368
rect 126 29266 160 29300
rect 126 29198 160 29232
rect 126 29130 160 29164
rect 126 29062 160 29096
rect 126 28994 160 29028
rect 126 28926 160 28960
rect 126 28858 160 28892
rect 126 28790 160 28824
rect 126 28722 160 28756
rect 126 28654 160 28688
rect 126 28586 160 28620
rect 126 28518 160 28552
rect 126 28450 160 28484
rect 126 28382 160 28416
rect 126 28314 160 28348
rect 126 28246 160 28280
rect 126 28178 160 28212
rect 126 28110 160 28144
rect 126 28042 160 28076
rect 126 27974 160 28008
rect 126 27906 160 27940
rect 126 27838 160 27872
rect 126 27770 160 27804
rect 126 27702 160 27736
rect 126 27634 160 27668
rect 126 27566 160 27600
rect 126 27498 160 27532
rect 126 27430 160 27464
rect 126 27362 160 27396
rect 126 27294 160 27328
rect 126 27226 160 27260
rect 126 27158 160 27192
rect 126 27090 160 27124
rect 126 27022 160 27056
rect 126 26954 160 26988
rect 126 26886 160 26920
rect 126 26818 160 26852
rect 126 26750 160 26784
rect 126 26682 160 26716
rect 126 26614 160 26648
rect 126 26546 160 26580
rect 126 26478 160 26512
rect 126 26410 160 26444
rect 126 26342 160 26376
rect 126 26274 160 26308
rect 126 26206 160 26240
rect 126 26138 160 26172
rect 126 26070 160 26104
rect 126 26002 160 26036
rect 126 25934 160 25968
rect 126 25866 160 25900
rect 126 25798 160 25832
rect 126 25730 160 25764
rect 126 25662 160 25696
rect 126 25594 160 25628
rect 126 25526 160 25560
rect 126 25458 160 25492
rect 126 25390 160 25424
rect 126 25322 160 25356
rect 126 25254 160 25288
rect 126 25186 160 25220
rect 126 25118 160 25152
rect 126 25050 160 25084
rect 126 24982 160 25016
rect 126 24914 160 24948
rect 126 24846 160 24880
rect 126 24778 160 24812
rect 126 24710 160 24744
rect 126 24642 160 24676
rect 126 24574 160 24608
rect 126 24506 160 24540
rect 126 24438 160 24472
rect 126 24370 160 24404
rect 126 24302 160 24336
rect 126 24234 160 24268
rect 126 24166 160 24200
rect 126 24098 160 24132
rect 126 24030 160 24064
rect 126 23962 160 23996
rect 126 23894 160 23928
rect 126 23826 160 23860
rect 126 23758 160 23792
rect 126 23690 160 23724
rect 126 23622 160 23656
rect 126 23554 160 23588
rect 126 23486 160 23520
rect 126 23418 160 23452
rect 126 23350 160 23384
rect 126 23282 160 23316
rect 126 23214 160 23248
rect 126 23146 160 23180
rect 126 23078 160 23112
rect 126 23010 160 23044
rect 126 22942 160 22976
rect 126 22874 160 22908
rect 126 22806 160 22840
rect 126 22738 160 22772
rect 126 22670 160 22704
rect 126 22602 160 22636
rect 126 22534 160 22568
rect 126 22466 160 22500
rect 126 22398 160 22432
rect 126 22330 160 22364
rect 126 22262 160 22296
rect 126 22194 160 22228
rect 126 22126 160 22160
rect 126 22058 160 22092
rect 126 21990 160 22024
rect 126 21922 160 21956
rect 126 21854 160 21888
rect 126 21786 160 21820
rect 126 21718 160 21752
rect 126 21650 160 21684
rect 126 21582 160 21616
rect 126 21514 160 21548
rect 126 21446 160 21480
rect 126 21378 160 21412
rect 126 21310 160 21344
rect 126 21242 160 21276
rect 126 21174 160 21208
rect 126 21106 160 21140
rect 126 21038 160 21072
rect 126 20970 160 21004
rect 126 20902 160 20936
rect 126 20834 160 20868
rect 126 20766 160 20800
rect 126 20698 160 20732
rect 126 20630 160 20664
rect 126 20562 160 20596
rect 126 20494 160 20528
rect 126 20426 160 20460
rect 126 20358 160 20392
rect 126 20290 160 20324
rect 126 20222 160 20256
rect 126 20154 160 20188
rect 126 20086 160 20120
rect 126 20018 160 20052
rect 126 19950 160 19984
rect 126 19882 160 19916
rect 126 19814 160 19848
rect 126 19746 160 19780
rect 126 19678 160 19712
rect 126 19610 160 19644
rect 126 19542 160 19576
rect 126 19474 160 19508
rect 126 19406 160 19440
rect 126 19338 160 19372
rect 126 19270 160 19304
rect 126 19202 160 19236
rect 126 19134 160 19168
rect 126 19066 160 19100
rect 126 18998 160 19032
rect 126 18930 160 18964
rect 126 18862 160 18896
rect 126 18794 160 18828
rect 126 18726 160 18760
rect 126 18658 160 18692
rect 126 18590 160 18624
rect 126 18522 160 18556
rect 126 18454 160 18488
rect 126 18386 160 18420
rect 126 18318 160 18352
rect 126 18250 160 18284
rect 126 18182 160 18216
rect 126 18114 160 18148
rect 126 18046 160 18080
rect 126 17978 160 18012
rect 126 17910 160 17944
rect 126 17842 160 17876
rect 126 17774 160 17808
rect 126 17706 160 17740
rect 126 17638 160 17672
rect 126 17570 160 17604
rect 126 17502 160 17536
rect 126 17434 160 17468
rect 126 17366 160 17400
rect 126 17298 160 17332
rect 126 17230 160 17264
rect 126 17162 160 17196
rect 126 17094 160 17128
rect 126 17026 160 17060
rect 126 16958 160 16992
rect 126 16890 160 16924
rect 126 16822 160 16856
rect 126 16754 160 16788
rect 126 16686 160 16720
rect 126 16618 160 16652
rect 126 16550 160 16584
rect 126 16482 160 16516
rect 126 16414 160 16448
rect 126 16346 160 16380
rect 126 16278 160 16312
rect 126 16210 160 16244
rect 126 16142 160 16176
rect 126 16074 160 16108
rect 126 16006 160 16040
rect 126 15938 160 15972
rect 126 15870 160 15904
rect 126 15802 160 15836
rect 126 15734 160 15768
rect 126 15666 160 15700
rect 126 15598 160 15632
rect 126 15530 160 15564
rect 126 15462 160 15496
rect 126 15394 160 15428
rect 126 15326 160 15360
rect 126 15258 160 15292
rect 126 15190 160 15224
rect 126 15122 160 15156
rect 126 15054 160 15088
rect 126 14986 160 15020
rect 126 14918 160 14952
rect 126 14850 160 14884
rect 126 14782 160 14816
rect 126 14714 160 14748
rect 126 14646 160 14680
rect 126 14578 160 14612
rect 126 14510 160 14544
rect 126 14442 160 14476
rect 126 14374 160 14408
rect 126 14306 160 14340
rect 126 14238 160 14272
rect 126 14170 160 14204
rect 126 14102 160 14136
rect 126 14034 160 14068
rect 126 13966 160 14000
rect 126 13898 160 13932
rect 126 13830 160 13864
rect 126 13762 160 13796
rect 126 13694 160 13728
rect 126 13626 160 13660
rect 126 13558 160 13592
rect 126 13490 160 13524
rect 126 13422 160 13456
rect 126 13354 160 13388
rect 126 13286 160 13320
rect 126 13218 160 13252
rect 126 13150 160 13184
rect 126 13082 160 13116
rect 126 13014 160 13048
rect 126 12946 160 12980
rect 126 12878 160 12912
rect 126 12810 160 12844
rect 126 12742 160 12776
rect 126 12674 160 12708
rect 126 12606 160 12640
rect 126 12538 160 12572
rect 126 12470 160 12504
rect 126 12402 160 12436
rect 126 12334 160 12368
rect 126 12266 160 12300
rect 126 12198 160 12232
rect 126 12130 160 12164
rect 126 12062 160 12096
rect 126 11994 160 12028
rect 126 11926 160 11960
rect 126 11858 160 11892
rect 126 11790 160 11824
rect 126 11722 160 11756
rect 126 11654 160 11688
rect 126 11586 160 11620
rect 126 11518 160 11552
rect 126 11450 160 11484
rect 126 11382 160 11416
rect 126 11314 160 11348
rect 126 11246 160 11280
rect 126 11178 160 11212
rect 126 11110 160 11144
rect 126 11042 160 11076
rect 126 10974 160 11008
rect 126 10906 160 10940
rect 126 10838 160 10872
rect 126 10770 160 10804
rect 126 10702 160 10736
rect 126 10634 160 10668
rect 126 10566 160 10600
rect 126 10498 160 10532
rect 126 10430 160 10464
rect 126 10362 160 10396
rect 126 10294 160 10328
rect 126 10226 160 10260
rect 126 10158 160 10192
rect 126 10090 160 10124
rect 126 10022 160 10056
rect 126 9954 160 9988
rect 126 9886 160 9920
rect 126 9818 160 9852
rect 126 9750 160 9784
rect 126 9682 160 9716
rect 126 9614 160 9648
rect 126 9546 160 9580
rect 126 9478 160 9512
rect 126 9410 160 9444
rect 126 9342 160 9376
rect 126 9274 160 9308
rect 126 9206 160 9240
rect 126 9138 160 9172
rect 126 9070 160 9104
rect 126 9002 160 9036
rect 126 8934 160 8968
rect 126 8866 160 8900
rect 126 8798 160 8832
rect 126 8730 160 8764
rect 126 8662 160 8696
rect 126 8594 160 8628
rect 126 8526 160 8560
rect 126 8458 160 8492
rect 126 8390 160 8424
rect 126 8322 160 8356
rect 126 8254 160 8288
rect 126 8186 160 8220
rect 126 8118 160 8152
rect 126 8050 160 8084
rect 126 7982 160 8016
rect 126 7914 160 7948
rect 126 7846 160 7880
rect 126 7778 160 7812
rect 126 7710 160 7744
rect 126 7642 160 7676
rect 126 7574 160 7608
rect 126 7506 160 7540
rect 126 7438 160 7472
rect 126 7370 160 7404
rect 126 7302 160 7336
rect 126 7234 160 7268
rect 126 7166 160 7200
rect 126 7098 160 7132
rect 126 7030 160 7064
rect 126 6962 160 6996
rect 126 6894 160 6928
rect 126 6826 160 6860
rect 126 6758 160 6792
rect 126 6690 160 6724
rect 126 6622 160 6656
rect 126 6554 160 6588
rect 126 6486 160 6520
rect 126 6418 160 6452
rect 126 6350 160 6384
rect 126 6282 160 6316
rect 126 6214 160 6248
rect 126 6146 160 6180
rect 126 6078 160 6112
rect 126 6010 160 6044
rect 126 5942 160 5976
rect 126 5874 160 5908
rect 126 5806 160 5840
rect 126 5738 160 5772
rect 126 5670 160 5704
rect 126 5602 160 5636
rect 126 5534 160 5568
rect 126 5466 160 5500
rect 126 5398 160 5432
rect 126 5330 160 5364
rect 126 5262 160 5296
rect 126 5194 160 5228
rect 126 5126 160 5160
rect 126 5058 160 5092
rect 126 4990 160 5024
rect 126 4922 160 4956
rect 126 4854 160 4888
rect 126 4786 160 4820
rect 126 4718 160 4752
rect 126 4650 160 4684
rect 126 4582 160 4616
rect 126 4514 160 4548
rect 126 4446 160 4480
rect 126 4378 160 4412
rect 126 4310 160 4344
rect 126 4242 160 4276
rect 126 4174 160 4208
rect 126 4106 160 4140
rect 126 4038 160 4072
rect 126 3970 160 4004
rect 126 3902 160 3936
rect 126 3834 160 3868
rect 126 3766 160 3800
rect 126 3698 160 3732
rect 126 3630 160 3664
rect 126 3562 160 3596
rect 126 3494 160 3528
rect 126 3426 160 3460
rect 126 3358 160 3392
rect 126 3290 160 3324
rect 126 3222 160 3256
rect 126 3154 160 3188
rect 126 3086 160 3120
rect 126 3018 160 3052
rect 126 2950 160 2984
rect 126 2882 160 2916
rect 126 2814 160 2848
rect 126 2746 160 2780
rect 126 2678 160 2712
rect 126 2610 160 2644
rect 126 2542 160 2576
rect 126 2474 160 2508
rect 126 2406 160 2440
rect 126 2338 160 2372
rect 126 2270 160 2304
rect 126 2202 160 2236
rect 126 2134 160 2168
rect 126 2066 160 2100
rect 126 1998 160 2032
rect 126 1930 160 1964
rect 126 1862 160 1896
rect 126 1794 160 1828
rect 126 1726 160 1760
rect 126 1658 160 1692
rect 126 1590 160 1624
rect 126 1522 160 1556
rect 126 1454 160 1488
rect 126 1386 160 1420
rect 126 1318 160 1352
rect 126 1250 160 1284
rect 126 1182 160 1216
rect 126 1114 160 1148
rect 126 1046 160 1080
rect 126 978 160 1012
rect 126 910 160 944
rect 126 842 160 876
rect 126 774 160 808
rect 126 706 160 740
rect 126 638 160 672
rect 126 570 160 604
rect 126 502 160 536
rect 3296 39124 3330 39158
rect 3296 39056 3330 39090
rect 3296 38988 3330 39022
rect 3296 38920 3330 38954
rect 3296 38852 3330 38886
rect 3296 38784 3330 38818
rect 3296 38716 3330 38750
rect 3296 38648 3330 38682
rect 3296 38580 3330 38614
rect 3296 38512 3330 38546
rect 3296 38444 3330 38478
rect 3296 38376 3330 38410
rect 3296 38308 3330 38342
rect 3296 38240 3330 38274
rect 3296 38172 3330 38206
rect 3296 38104 3330 38138
rect 3296 38036 3330 38070
rect 3296 37968 3330 38002
rect 3296 37900 3330 37934
rect 3296 37832 3330 37866
rect 3296 37764 3330 37798
rect 3296 37696 3330 37730
rect 3296 37628 3330 37662
rect 3296 37560 3330 37594
rect 3296 37492 3330 37526
rect 3296 37424 3330 37458
rect 3296 37356 3330 37390
rect 3296 37288 3330 37322
rect 3296 37220 3330 37254
rect 3296 37152 3330 37186
rect 3296 37084 3330 37118
rect 3296 37016 3330 37050
rect 3296 36948 3330 36982
rect 3296 36880 3330 36914
rect 3296 36812 3330 36846
rect 3296 36744 3330 36778
rect 3296 36676 3330 36710
rect 3296 36608 3330 36642
rect 3296 36540 3330 36574
rect 3296 36472 3330 36506
rect 3296 36404 3330 36438
rect 3296 36336 3330 36370
rect 3296 36268 3330 36302
rect 3296 36200 3330 36234
rect 3296 36132 3330 36166
rect 3296 36064 3330 36098
rect 3296 35996 3330 36030
rect 3296 35928 3330 35962
rect 3296 35860 3330 35894
rect 3296 35792 3330 35826
rect 3296 35724 3330 35758
rect 3296 35656 3330 35690
rect 3296 35588 3330 35622
rect 3296 35520 3330 35554
rect 3296 35452 3330 35486
rect 3296 35384 3330 35418
rect 3296 35316 3330 35350
rect 3296 35248 3330 35282
rect 3296 35180 3330 35214
rect 3296 35112 3330 35146
rect 3296 35044 3330 35078
rect 3296 34976 3330 35010
rect 3296 34908 3330 34942
rect 3296 34840 3330 34874
rect 3296 34772 3330 34806
rect 3296 34704 3330 34738
rect 3296 34636 3330 34670
rect 3296 34568 3330 34602
rect 3296 34500 3330 34534
rect 3296 34432 3330 34466
rect 3296 34364 3330 34398
rect 3296 34296 3330 34330
rect 3296 34228 3330 34262
rect 3296 34160 3330 34194
rect 3296 34092 3330 34126
rect 3296 34024 3330 34058
rect 3296 33956 3330 33990
rect 3296 33888 3330 33922
rect 3296 33820 3330 33854
rect 3296 33752 3330 33786
rect 3296 33684 3330 33718
rect 3296 33616 3330 33650
rect 3296 33548 3330 33582
rect 3296 33480 3330 33514
rect 3296 33412 3330 33446
rect 3296 33344 3330 33378
rect 3296 33276 3330 33310
rect 3296 33208 3330 33242
rect 3296 33140 3330 33174
rect 3296 33072 3330 33106
rect 3296 33004 3330 33038
rect 3296 32936 3330 32970
rect 3296 32868 3330 32902
rect 3296 32800 3330 32834
rect 3296 32732 3330 32766
rect 3296 32664 3330 32698
rect 3296 32596 3330 32630
rect 3296 32528 3330 32562
rect 3296 32460 3330 32494
rect 3296 32392 3330 32426
rect 3296 32324 3330 32358
rect 3296 32256 3330 32290
rect 3296 32188 3330 32222
rect 3296 32120 3330 32154
rect 3296 32052 3330 32086
rect 3296 31984 3330 32018
rect 3296 31916 3330 31950
rect 3296 31848 3330 31882
rect 3296 31780 3330 31814
rect 3296 31712 3330 31746
rect 3296 31644 3330 31678
rect 3296 31576 3330 31610
rect 3296 31508 3330 31542
rect 3296 31440 3330 31474
rect 3296 31372 3330 31406
rect 3296 31304 3330 31338
rect 3296 31236 3330 31270
rect 3296 31168 3330 31202
rect 3296 31100 3330 31134
rect 3296 31032 3330 31066
rect 3296 30964 3330 30998
rect 3296 30896 3330 30930
rect 3296 30828 3330 30862
rect 3296 30760 3330 30794
rect 3296 30692 3330 30726
rect 3296 30624 3330 30658
rect 3296 30556 3330 30590
rect 3296 30488 3330 30522
rect 3296 30420 3330 30454
rect 3296 30352 3330 30386
rect 3296 30284 3330 30318
rect 3296 30216 3330 30250
rect 3296 30148 3330 30182
rect 3296 30080 3330 30114
rect 3296 30012 3330 30046
rect 3296 29944 3330 29978
rect 3296 29876 3330 29910
rect 3296 29808 3330 29842
rect 3296 29740 3330 29774
rect 3296 29672 3330 29706
rect 3296 29604 3330 29638
rect 3296 29536 3330 29570
rect 3296 29468 3330 29502
rect 3296 29400 3330 29434
rect 3296 29332 3330 29366
rect 3296 29264 3330 29298
rect 3296 29196 3330 29230
rect 3296 29128 3330 29162
rect 3296 29060 3330 29094
rect 3296 28992 3330 29026
rect 3296 28924 3330 28958
rect 3296 28856 3330 28890
rect 3296 28788 3330 28822
rect 3296 28720 3330 28754
rect 3296 28652 3330 28686
rect 3296 28584 3330 28618
rect 3296 28516 3330 28550
rect 3296 28448 3330 28482
rect 3296 28380 3330 28414
rect 3296 28312 3330 28346
rect 3296 28244 3330 28278
rect 3296 28176 3330 28210
rect 3296 28108 3330 28142
rect 3296 28040 3330 28074
rect 3296 27972 3330 28006
rect 3296 27904 3330 27938
rect 3296 27836 3330 27870
rect 3296 27768 3330 27802
rect 3296 27700 3330 27734
rect 3296 27632 3330 27666
rect 3296 27564 3330 27598
rect 3296 27496 3330 27530
rect 3296 27428 3330 27462
rect 3296 27360 3330 27394
rect 3296 27292 3330 27326
rect 3296 27224 3330 27258
rect 3296 27156 3330 27190
rect 3296 27088 3330 27122
rect 3296 27020 3330 27054
rect 3296 26952 3330 26986
rect 3296 26884 3330 26918
rect 3296 26816 3330 26850
rect 3296 26748 3330 26782
rect 3296 26680 3330 26714
rect 3296 26612 3330 26646
rect 3296 26544 3330 26578
rect 3296 26476 3330 26510
rect 3296 26408 3330 26442
rect 3296 26340 3330 26374
rect 3296 26272 3330 26306
rect 3296 26204 3330 26238
rect 3296 26136 3330 26170
rect 3296 26068 3330 26102
rect 3296 26000 3330 26034
rect 3296 25932 3330 25966
rect 3296 25864 3330 25898
rect 3296 25796 3330 25830
rect 3296 25728 3330 25762
rect 3296 25660 3330 25694
rect 3296 25592 3330 25626
rect 3296 25524 3330 25558
rect 3296 25456 3330 25490
rect 3296 25388 3330 25422
rect 3296 25320 3330 25354
rect 3296 25252 3330 25286
rect 3296 25184 3330 25218
rect 3296 25116 3330 25150
rect 3296 25048 3330 25082
rect 3296 24980 3330 25014
rect 3296 24912 3330 24946
rect 3296 24844 3330 24878
rect 3296 24776 3330 24810
rect 3296 24708 3330 24742
rect 3296 24640 3330 24674
rect 3296 24572 3330 24606
rect 3296 24504 3330 24538
rect 3296 24436 3330 24470
rect 3296 24368 3330 24402
rect 3296 24300 3330 24334
rect 3296 24232 3330 24266
rect 3296 24164 3330 24198
rect 3296 24096 3330 24130
rect 3296 24028 3330 24062
rect 3296 23960 3330 23994
rect 3296 23892 3330 23926
rect 3296 23824 3330 23858
rect 3296 23756 3330 23790
rect 3296 23688 3330 23722
rect 3296 23620 3330 23654
rect 3296 23552 3330 23586
rect 3296 23484 3330 23518
rect 3296 23416 3330 23450
rect 3296 23348 3330 23382
rect 3296 23280 3330 23314
rect 3296 23212 3330 23246
rect 3296 23144 3330 23178
rect 3296 23076 3330 23110
rect 3296 23008 3330 23042
rect 3296 22940 3330 22974
rect 3296 22872 3330 22906
rect 3296 22804 3330 22838
rect 3296 22736 3330 22770
rect 3296 22668 3330 22702
rect 3296 22600 3330 22634
rect 3296 22532 3330 22566
rect 3296 22464 3330 22498
rect 3296 22396 3330 22430
rect 3296 22328 3330 22362
rect 3296 22260 3330 22294
rect 3296 22192 3330 22226
rect 3296 22124 3330 22158
rect 3296 22056 3330 22090
rect 3296 21988 3330 22022
rect 3296 21920 3330 21954
rect 3296 21852 3330 21886
rect 3296 21784 3330 21818
rect 3296 21716 3330 21750
rect 3296 21648 3330 21682
rect 3296 21580 3330 21614
rect 3296 21512 3330 21546
rect 3296 21444 3330 21478
rect 3296 21376 3330 21410
rect 3296 21308 3330 21342
rect 3296 21240 3330 21274
rect 3296 21172 3330 21206
rect 3296 21104 3330 21138
rect 3296 21036 3330 21070
rect 3296 20968 3330 21002
rect 3296 20900 3330 20934
rect 3296 20832 3330 20866
rect 3296 20764 3330 20798
rect 3296 20696 3330 20730
rect 3296 20628 3330 20662
rect 3296 20560 3330 20594
rect 3296 20492 3330 20526
rect 3296 20424 3330 20458
rect 3296 20356 3330 20390
rect 3296 20288 3330 20322
rect 3296 20220 3330 20254
rect 3296 20152 3330 20186
rect 3296 20084 3330 20118
rect 3296 20016 3330 20050
rect 3296 19948 3330 19982
rect 3296 19880 3330 19914
rect 3296 19812 3330 19846
rect 3296 19744 3330 19778
rect 3296 19676 3330 19710
rect 3296 19608 3330 19642
rect 3296 19540 3330 19574
rect 3296 19472 3330 19506
rect 3296 19404 3330 19438
rect 3296 19336 3330 19370
rect 3296 19268 3330 19302
rect 3296 19200 3330 19234
rect 3296 19132 3330 19166
rect 3296 19064 3330 19098
rect 3296 18996 3330 19030
rect 3296 18928 3330 18962
rect 3296 18860 3330 18894
rect 3296 18792 3330 18826
rect 3296 18724 3330 18758
rect 3296 18656 3330 18690
rect 3296 18588 3330 18622
rect 3296 18520 3330 18554
rect 3296 18452 3330 18486
rect 3296 18384 3330 18418
rect 3296 18316 3330 18350
rect 3296 18248 3330 18282
rect 3296 18180 3330 18214
rect 3296 18112 3330 18146
rect 3296 18044 3330 18078
rect 3296 17976 3330 18010
rect 3296 17908 3330 17942
rect 3296 17840 3330 17874
rect 3296 17772 3330 17806
rect 3296 17704 3330 17738
rect 3296 17636 3330 17670
rect 3296 17568 3330 17602
rect 3296 17500 3330 17534
rect 3296 17432 3330 17466
rect 3296 17364 3330 17398
rect 3296 17296 3330 17330
rect 3296 17228 3330 17262
rect 3296 17160 3330 17194
rect 3296 17092 3330 17126
rect 3296 17024 3330 17058
rect 3296 16956 3330 16990
rect 3296 16888 3330 16922
rect 3296 16820 3330 16854
rect 3296 16752 3330 16786
rect 3296 16684 3330 16718
rect 3296 16616 3330 16650
rect 3296 16548 3330 16582
rect 3296 16480 3330 16514
rect 3296 16412 3330 16446
rect 3296 16344 3330 16378
rect 3296 16276 3330 16310
rect 3296 16208 3330 16242
rect 3296 16140 3330 16174
rect 3296 16072 3330 16106
rect 3296 16004 3330 16038
rect 3296 15936 3330 15970
rect 3296 15868 3330 15902
rect 3296 15800 3330 15834
rect 3296 15732 3330 15766
rect 3296 15664 3330 15698
rect 3296 15596 3330 15630
rect 3296 15528 3330 15562
rect 3296 15460 3330 15494
rect 3296 15392 3330 15426
rect 3296 15324 3330 15358
rect 3296 15256 3330 15290
rect 3296 15188 3330 15222
rect 3296 15120 3330 15154
rect 3296 15052 3330 15086
rect 3296 14984 3330 15018
rect 3296 14916 3330 14950
rect 3296 14848 3330 14882
rect 3296 14780 3330 14814
rect 3296 14712 3330 14746
rect 3296 14644 3330 14678
rect 3296 14576 3330 14610
rect 3296 14508 3330 14542
rect 3296 14440 3330 14474
rect 3296 14372 3330 14406
rect 3296 14304 3330 14338
rect 3296 14236 3330 14270
rect 3296 14168 3330 14202
rect 3296 14100 3330 14134
rect 3296 14032 3330 14066
rect 3296 13964 3330 13998
rect 3296 13896 3330 13930
rect 3296 13828 3330 13862
rect 3296 13760 3330 13794
rect 3296 13692 3330 13726
rect 3296 13624 3330 13658
rect 3296 13556 3330 13590
rect 3296 13488 3330 13522
rect 3296 13420 3330 13454
rect 3296 13352 3330 13386
rect 3296 13284 3330 13318
rect 3296 13216 3330 13250
rect 3296 13148 3330 13182
rect 3296 13080 3330 13114
rect 3296 13012 3330 13046
rect 3296 12944 3330 12978
rect 3296 12876 3330 12910
rect 3296 12808 3330 12842
rect 3296 12740 3330 12774
rect 3296 12672 3330 12706
rect 3296 12604 3330 12638
rect 3296 12536 3330 12570
rect 3296 12468 3330 12502
rect 3296 12400 3330 12434
rect 3296 12332 3330 12366
rect 3296 12264 3330 12298
rect 3296 12196 3330 12230
rect 3296 12128 3330 12162
rect 3296 12060 3330 12094
rect 3296 11992 3330 12026
rect 3296 11924 3330 11958
rect 3296 11856 3330 11890
rect 3296 11788 3330 11822
rect 3296 11720 3330 11754
rect 3296 11652 3330 11686
rect 3296 11584 3330 11618
rect 3296 11516 3330 11550
rect 3296 11448 3330 11482
rect 3296 11380 3330 11414
rect 3296 11312 3330 11346
rect 3296 11244 3330 11278
rect 3296 11176 3330 11210
rect 3296 11108 3330 11142
rect 3296 11040 3330 11074
rect 3296 10972 3330 11006
rect 3296 10904 3330 10938
rect 3296 10836 3330 10870
rect 3296 10768 3330 10802
rect 3296 10700 3330 10734
rect 3296 10632 3330 10666
rect 3296 10564 3330 10598
rect 3296 10496 3330 10530
rect 3296 10428 3330 10462
rect 3296 10360 3330 10394
rect 3296 10292 3330 10326
rect 3296 10224 3330 10258
rect 3296 10156 3330 10190
rect 3296 10088 3330 10122
rect 3296 10020 3330 10054
rect 3296 9952 3330 9986
rect 3296 9884 3330 9918
rect 3296 9816 3330 9850
rect 3296 9748 3330 9782
rect 3296 9680 3330 9714
rect 3296 9612 3330 9646
rect 3296 9544 3330 9578
rect 3296 9476 3330 9510
rect 3296 9408 3330 9442
rect 3296 9340 3330 9374
rect 3296 9272 3330 9306
rect 3296 9204 3330 9238
rect 3296 9136 3330 9170
rect 3296 9068 3330 9102
rect 3296 9000 3330 9034
rect 3296 8932 3330 8966
rect 3296 8864 3330 8898
rect 3296 8796 3330 8830
rect 3296 8728 3330 8762
rect 3296 8660 3330 8694
rect 3296 8592 3330 8626
rect 3296 8524 3330 8558
rect 3296 8456 3330 8490
rect 3296 8388 3330 8422
rect 3296 8320 3330 8354
rect 3296 8252 3330 8286
rect 3296 8184 3330 8218
rect 3296 8116 3330 8150
rect 3296 8048 3330 8082
rect 3296 7980 3330 8014
rect 3296 7912 3330 7946
rect 3296 7844 3330 7878
rect 3296 7776 3330 7810
rect 3296 7708 3330 7742
rect 3296 7640 3330 7674
rect 3296 7572 3330 7606
rect 3296 7504 3330 7538
rect 3296 7436 3330 7470
rect 3296 7368 3330 7402
rect 3296 7300 3330 7334
rect 3296 7232 3330 7266
rect 3296 7164 3330 7198
rect 3296 7096 3330 7130
rect 3296 7028 3330 7062
rect 3296 6960 3330 6994
rect 3296 6892 3330 6926
rect 3296 6824 3330 6858
rect 3296 6756 3330 6790
rect 3296 6688 3330 6722
rect 3296 6620 3330 6654
rect 3296 6552 3330 6586
rect 3296 6484 3330 6518
rect 3296 6416 3330 6450
rect 3296 6348 3330 6382
rect 3296 6280 3330 6314
rect 3296 6212 3330 6246
rect 3296 6144 3330 6178
rect 3296 6076 3330 6110
rect 3296 6008 3330 6042
rect 3296 5940 3330 5974
rect 3296 5872 3330 5906
rect 3296 5804 3330 5838
rect 3296 5736 3330 5770
rect 3296 5668 3330 5702
rect 3296 5600 3330 5634
rect 3296 5532 3330 5566
rect 3296 5464 3330 5498
rect 3296 5396 3330 5430
rect 3296 5328 3330 5362
rect 3296 5260 3330 5294
rect 3296 5192 3330 5226
rect 3296 5124 3330 5158
rect 3296 5056 3330 5090
rect 3296 4988 3330 5022
rect 3296 4920 3330 4954
rect 3296 4852 3330 4886
rect 3296 4784 3330 4818
rect 3296 4716 3330 4750
rect 3296 4648 3330 4682
rect 3296 4580 3330 4614
rect 3296 4512 3330 4546
rect 3296 4444 3330 4478
rect 3296 4376 3330 4410
rect 3296 4308 3330 4342
rect 3296 4240 3330 4274
rect 3296 4172 3330 4206
rect 3296 4104 3330 4138
rect 3296 4036 3330 4070
rect 3296 3968 3330 4002
rect 3296 3900 3330 3934
rect 3296 3832 3330 3866
rect 3296 3764 3330 3798
rect 3296 3696 3330 3730
rect 3296 3628 3330 3662
rect 3296 3560 3330 3594
rect 3296 3492 3330 3526
rect 3296 3424 3330 3458
rect 3296 3356 3330 3390
rect 3296 3288 3330 3322
rect 3296 3220 3330 3254
rect 3296 3152 3330 3186
rect 3296 3084 3330 3118
rect 3296 3016 3330 3050
rect 3296 2948 3330 2982
rect 3296 2880 3330 2914
rect 3296 2812 3330 2846
rect 3296 2744 3330 2778
rect 3296 2676 3330 2710
rect 3296 2608 3330 2642
rect 3296 2540 3330 2574
rect 3296 2472 3330 2506
rect 3296 2404 3330 2438
rect 3296 2336 3330 2370
rect 3296 2268 3330 2302
rect 3296 2200 3330 2234
rect 3296 2132 3330 2166
rect 3296 2064 3330 2098
rect 3296 1996 3330 2030
rect 3296 1928 3330 1962
rect 3296 1860 3330 1894
rect 3296 1792 3330 1826
rect 3296 1724 3330 1758
rect 3296 1656 3330 1690
rect 3296 1588 3330 1622
rect 3296 1520 3330 1554
rect 3296 1452 3330 1486
rect 3296 1384 3330 1418
rect 3296 1316 3330 1350
rect 3296 1248 3330 1282
rect 3296 1180 3330 1214
rect 3296 1112 3330 1146
rect 3296 1044 3330 1078
rect 3296 976 3330 1010
rect 3296 908 3330 942
rect 3296 840 3330 874
rect 3296 772 3330 806
rect 3296 704 3330 738
rect 3296 636 3330 670
rect 3296 568 3330 602
rect 126 434 160 468
rect 126 366 160 400
rect 126 252 160 332
rect 126 160 160 218
rect 3296 500 3330 534
rect 3296 432 3330 466
rect 3296 364 3330 398
rect 3296 296 3330 330
rect 3296 228 3330 262
rect 3296 160 3330 194
rect 126 126 194 160
rect 228 126 262 160
rect 296 126 330 160
rect 364 126 398 160
rect 432 126 466 160
rect 500 126 534 160
rect 568 126 602 160
rect 636 126 670 160
rect 704 126 738 160
rect 772 126 806 160
rect 840 126 874 160
rect 908 126 942 160
rect 976 126 1010 160
rect 1044 126 1078 160
rect 1112 126 1146 160
rect 1180 126 1214 160
rect 1248 126 1282 160
rect 1316 126 1350 160
rect 1384 126 1418 160
rect 1452 126 1486 160
rect 1520 126 1554 160
rect 1588 126 1622 160
rect 1656 126 1690 160
rect 1724 126 1758 160
rect 1792 126 1826 160
rect 1860 126 1894 160
rect 1928 126 1962 160
rect 1996 126 2030 160
rect 2064 126 2098 160
rect 2132 126 2166 160
rect 2200 126 2234 160
rect 2268 126 2302 160
rect 2336 126 2370 160
rect 2404 126 2438 160
rect 2472 126 2506 160
rect 2540 126 2574 160
rect 2608 126 2642 160
rect 2676 126 2710 160
rect 2744 126 2778 160
rect 2812 126 2846 160
rect 2880 126 2914 160
rect 2948 126 2982 160
rect 3016 126 3050 160
rect 3084 126 3118 160
rect 3152 126 3186 160
rect 3220 126 3330 160
<< mvpsubdiffcont >>
rect 465 39144 499 39178
rect 533 39144 567 39178
rect 601 39144 635 39178
rect 669 39144 703 39178
rect 737 39144 771 39178
rect 805 39144 839 39178
rect 873 39144 907 39178
rect 941 39144 975 39178
rect 1009 39144 1043 39178
rect 1077 39144 1111 39178
rect 1145 39144 1179 39178
rect 1213 39144 1247 39178
rect 1281 39144 1315 39178
rect 1349 39144 1383 39178
rect 1417 39144 1451 39178
rect 1485 39144 1519 39178
rect 1553 39144 1587 39178
rect 1621 39144 1655 39178
rect 1689 39144 1723 39178
rect 1757 39144 1791 39178
rect 1825 39144 1859 39178
rect 1893 39144 1927 39178
rect 1961 39144 1995 39178
rect 2029 39144 2063 39178
rect 2097 39144 2131 39178
rect 2165 39144 2199 39178
rect 2233 39144 2267 39178
rect 2301 39144 2335 39178
rect 2369 39144 2403 39178
rect 2437 39144 2471 39178
rect 2505 39144 2539 39178
rect 2573 39144 2607 39178
rect 2641 39144 2675 39178
rect 2709 39144 2743 39178
rect 2777 39144 2811 39178
rect 2845 39144 2879 39178
rect 2913 39144 2947 39178
rect 2981 39144 3015 39178
rect 386 39089 420 39123
rect 3036 39076 3070 39110
rect 386 39021 420 39055
rect 3036 39008 3070 39042
rect 386 38953 420 38987
rect 386 38885 420 38919
rect 386 38817 420 38851
rect 386 38749 420 38783
rect 386 38681 420 38715
rect 386 38613 420 38647
rect 386 38545 420 38579
rect 386 38477 420 38511
rect 386 38409 420 38443
rect 386 38341 420 38375
rect 386 38273 420 38307
rect 386 38205 420 38239
rect 386 38137 420 38171
rect 386 38069 420 38103
rect 386 38001 420 38035
rect 386 37933 420 37967
rect 386 37865 420 37899
rect 386 37797 420 37831
rect 386 37729 420 37763
rect 386 37661 420 37695
rect 386 37593 420 37627
rect 386 37525 420 37559
rect 386 37457 420 37491
rect 386 37389 420 37423
rect 386 37321 420 37355
rect 386 37253 420 37287
rect 386 37185 420 37219
rect 386 37117 420 37151
rect 386 37049 420 37083
rect 386 36981 420 37015
rect 386 36913 420 36947
rect 3036 38940 3070 38974
rect 3036 38872 3070 38906
rect 3036 38804 3070 38838
rect 3036 38736 3070 38770
rect 3036 38668 3070 38702
rect 3036 38600 3070 38634
rect 3036 38532 3070 38566
rect 3036 38464 3070 38498
rect 3036 38396 3070 38430
rect 3036 38328 3070 38362
rect 3036 38260 3070 38294
rect 3036 38192 3070 38226
rect 3036 38124 3070 38158
rect 3036 38056 3070 38090
rect 3036 37988 3070 38022
rect 3036 37920 3070 37954
rect 3036 37852 3070 37886
rect 3036 37784 3070 37818
rect 3036 37716 3070 37750
rect 3036 37648 3070 37682
rect 3036 37580 3070 37614
rect 3036 37512 3070 37546
rect 3036 37444 3070 37478
rect 3036 37376 3070 37410
rect 3036 37308 3070 37342
rect 3036 37240 3070 37274
rect 3036 37172 3070 37206
rect 3036 37104 3070 37138
rect 3036 37036 3070 37070
rect 3036 36968 3070 37002
rect 386 36845 420 36879
rect 3036 36900 3070 36934
rect 386 36777 420 36811
rect 386 36709 420 36743
rect 386 36641 420 36675
rect 386 36573 420 36607
rect 386 36505 420 36539
rect 386 36437 420 36471
rect 386 36369 420 36403
rect 386 36301 420 36335
rect 386 36233 420 36267
rect 386 36165 420 36199
rect 386 36097 420 36131
rect 386 36029 420 36063
rect 386 35961 420 35995
rect 386 35893 420 35927
rect 386 35825 420 35859
rect 386 35757 420 35791
rect 386 35689 420 35723
rect 386 35621 420 35655
rect 386 35553 420 35587
rect 386 35485 420 35519
rect 386 35417 420 35451
rect 386 35349 420 35383
rect 386 35281 420 35315
rect 386 35213 420 35247
rect 386 35145 420 35179
rect 386 35077 420 35111
rect 386 35009 420 35043
rect 386 34941 420 34975
rect 386 34873 420 34907
rect 386 34805 420 34839
rect 3036 36832 3070 36866
rect 3036 36764 3070 36798
rect 3036 36696 3070 36730
rect 3036 36628 3070 36662
rect 3036 36560 3070 36594
rect 3036 36492 3070 36526
rect 3036 36424 3070 36458
rect 3036 36356 3070 36390
rect 3036 36288 3070 36322
rect 3036 36220 3070 36254
rect 3036 36152 3070 36186
rect 3036 36084 3070 36118
rect 3036 36016 3070 36050
rect 3036 35948 3070 35982
rect 3036 35880 3070 35914
rect 3036 35812 3070 35846
rect 3036 35744 3070 35778
rect 3036 35676 3070 35710
rect 3036 35608 3070 35642
rect 3036 35540 3070 35574
rect 3036 35472 3070 35506
rect 3036 35404 3070 35438
rect 3036 35336 3070 35370
rect 3036 35268 3070 35302
rect 3036 35200 3070 35234
rect 3036 35132 3070 35166
rect 3036 35064 3070 35098
rect 3036 34996 3070 35030
rect 3036 34928 3070 34962
rect 3036 34860 3070 34894
rect 386 34737 420 34771
rect 3036 34792 3070 34826
rect 386 34669 420 34703
rect 386 34601 420 34635
rect 386 34533 420 34567
rect 386 34465 420 34499
rect 386 34397 420 34431
rect 386 34329 420 34363
rect 386 34261 420 34295
rect 386 34193 420 34227
rect 386 34125 420 34159
rect 386 34057 420 34091
rect 386 33989 420 34023
rect 386 33921 420 33955
rect 386 33853 420 33887
rect 386 33785 420 33819
rect 386 33717 420 33751
rect 386 33649 420 33683
rect 386 33581 420 33615
rect 386 33513 420 33547
rect 386 33445 420 33479
rect 386 33377 420 33411
rect 386 33309 420 33343
rect 386 33241 420 33275
rect 386 33173 420 33207
rect 386 33105 420 33139
rect 386 33037 420 33071
rect 386 32969 420 33003
rect 386 32901 420 32935
rect 386 32833 420 32867
rect 386 32765 420 32799
rect 386 32697 420 32731
rect 3036 34724 3070 34758
rect 3036 34656 3070 34690
rect 3036 34588 3070 34622
rect 3036 34520 3070 34554
rect 3036 34452 3070 34486
rect 3036 34384 3070 34418
rect 3036 34316 3070 34350
rect 3036 34248 3070 34282
rect 3036 34180 3070 34214
rect 3036 34112 3070 34146
rect 3036 34044 3070 34078
rect 3036 33976 3070 34010
rect 3036 33908 3070 33942
rect 3036 33840 3070 33874
rect 3036 33772 3070 33806
rect 3036 33704 3070 33738
rect 3036 33636 3070 33670
rect 3036 33568 3070 33602
rect 3036 33500 3070 33534
rect 3036 33432 3070 33466
rect 3036 33364 3070 33398
rect 3036 33296 3070 33330
rect 3036 33228 3070 33262
rect 3036 33160 3070 33194
rect 3036 33092 3070 33126
rect 3036 33024 3070 33058
rect 3036 32956 3070 32990
rect 3036 32888 3070 32922
rect 3036 32820 3070 32854
rect 3036 32752 3070 32786
rect 3036 32684 3070 32718
rect 386 32629 420 32663
rect 3036 32616 3070 32650
rect 386 32561 420 32595
rect 386 32493 420 32527
rect 386 32425 420 32459
rect 386 32357 420 32391
rect 386 32289 420 32323
rect 386 32221 420 32255
rect 386 32153 420 32187
rect 386 32085 420 32119
rect 386 32017 420 32051
rect 386 31949 420 31983
rect 386 31881 420 31915
rect 386 31813 420 31847
rect 386 31745 420 31779
rect 386 31677 420 31711
rect 386 31609 420 31643
rect 386 31541 420 31575
rect 386 31473 420 31507
rect 386 31405 420 31439
rect 386 31337 420 31371
rect 386 31269 420 31303
rect 386 31201 420 31235
rect 386 31133 420 31167
rect 386 31065 420 31099
rect 386 30997 420 31031
rect 386 30929 420 30963
rect 386 30861 420 30895
rect 386 30793 420 30827
rect 386 30725 420 30759
rect 386 30657 420 30691
rect 386 30589 420 30623
rect 386 30521 420 30555
rect 3036 32548 3070 32582
rect 3036 32480 3070 32514
rect 3036 32412 3070 32446
rect 3036 32344 3070 32378
rect 3036 32276 3070 32310
rect 3036 32208 3070 32242
rect 3036 32140 3070 32174
rect 3036 32072 3070 32106
rect 3036 32004 3070 32038
rect 3036 31936 3070 31970
rect 3036 31868 3070 31902
rect 3036 31800 3070 31834
rect 3036 31732 3070 31766
rect 3036 31664 3070 31698
rect 3036 31596 3070 31630
rect 3036 31528 3070 31562
rect 3036 31460 3070 31494
rect 3036 31392 3070 31426
rect 3036 31324 3070 31358
rect 3036 31256 3070 31290
rect 3036 31188 3070 31222
rect 3036 31120 3070 31154
rect 3036 31052 3070 31086
rect 3036 30984 3070 31018
rect 3036 30916 3070 30950
rect 3036 30848 3070 30882
rect 3036 30780 3070 30814
rect 3036 30712 3070 30746
rect 3036 30644 3070 30678
rect 3036 30576 3070 30610
rect 386 30453 420 30487
rect 3036 30508 3070 30542
rect 386 30385 420 30419
rect 386 30317 420 30351
rect 386 30249 420 30283
rect 386 30181 420 30215
rect 386 30113 420 30147
rect 386 30045 420 30079
rect 386 29977 420 30011
rect 386 29909 420 29943
rect 386 29841 420 29875
rect 386 29773 420 29807
rect 386 29705 420 29739
rect 386 29637 420 29671
rect 386 29569 420 29603
rect 386 29501 420 29535
rect 386 29433 420 29467
rect 386 29365 420 29399
rect 386 29297 420 29331
rect 386 29229 420 29263
rect 386 29161 420 29195
rect 386 29093 420 29127
rect 386 29025 420 29059
rect 386 28957 420 28991
rect 386 28889 420 28923
rect 386 28821 420 28855
rect 386 28753 420 28787
rect 386 28685 420 28719
rect 386 28617 420 28651
rect 386 28549 420 28583
rect 386 28481 420 28515
rect 386 28413 420 28447
rect 3036 30440 3070 30474
rect 3036 30372 3070 30406
rect 3036 30304 3070 30338
rect 3036 30236 3070 30270
rect 3036 30168 3070 30202
rect 3036 30100 3070 30134
rect 3036 30032 3070 30066
rect 3036 29964 3070 29998
rect 3036 29896 3070 29930
rect 3036 29828 3070 29862
rect 3036 29760 3070 29794
rect 3036 29692 3070 29726
rect 3036 29624 3070 29658
rect 3036 29556 3070 29590
rect 3036 29488 3070 29522
rect 3036 29420 3070 29454
rect 3036 29352 3070 29386
rect 3036 29284 3070 29318
rect 3036 29216 3070 29250
rect 3036 29148 3070 29182
rect 3036 29080 3070 29114
rect 3036 29012 3070 29046
rect 3036 28944 3070 28978
rect 3036 28876 3070 28910
rect 3036 28808 3070 28842
rect 3036 28740 3070 28774
rect 3036 28672 3070 28706
rect 3036 28604 3070 28638
rect 3036 28536 3070 28570
rect 3036 28468 3070 28502
rect 386 28345 420 28379
rect 3036 28400 3070 28434
rect 386 28277 420 28311
rect 386 28209 420 28243
rect 386 28141 420 28175
rect 386 28073 420 28107
rect 386 28005 420 28039
rect 386 27937 420 27971
rect 386 27869 420 27903
rect 386 27801 420 27835
rect 386 27733 420 27767
rect 386 27665 420 27699
rect 386 27597 420 27631
rect 386 27529 420 27563
rect 386 27461 420 27495
rect 386 27393 420 27427
rect 386 27325 420 27359
rect 386 27257 420 27291
rect 386 27189 420 27223
rect 386 27121 420 27155
rect 386 27053 420 27087
rect 386 26985 420 27019
rect 386 26917 420 26951
rect 386 26849 420 26883
rect 386 26781 420 26815
rect 386 26713 420 26747
rect 386 26645 420 26679
rect 386 26577 420 26611
rect 386 26509 420 26543
rect 386 26441 420 26475
rect 386 26373 420 26407
rect 386 26305 420 26339
rect 3036 28332 3070 28366
rect 3036 28264 3070 28298
rect 3036 28196 3070 28230
rect 3036 28128 3070 28162
rect 3036 28060 3070 28094
rect 3036 27992 3070 28026
rect 3036 27924 3070 27958
rect 3036 27856 3070 27890
rect 3036 27788 3070 27822
rect 3036 27720 3070 27754
rect 3036 27652 3070 27686
rect 3036 27584 3070 27618
rect 3036 27516 3070 27550
rect 3036 27448 3070 27482
rect 3036 27380 3070 27414
rect 3036 27312 3070 27346
rect 3036 27244 3070 27278
rect 3036 27176 3070 27210
rect 3036 27108 3070 27142
rect 3036 27040 3070 27074
rect 3036 26972 3070 27006
rect 3036 26904 3070 26938
rect 3036 26836 3070 26870
rect 3036 26768 3070 26802
rect 3036 26700 3070 26734
rect 3036 26632 3070 26666
rect 3036 26564 3070 26598
rect 3036 26496 3070 26530
rect 3036 26428 3070 26462
rect 3036 26360 3070 26394
rect 3036 26292 3070 26326
rect 386 26237 420 26271
rect 3036 26224 3070 26258
rect 386 26169 420 26203
rect 386 26101 420 26135
rect 386 26033 420 26067
rect 386 25965 420 25999
rect 386 25897 420 25931
rect 386 25829 420 25863
rect 386 25761 420 25795
rect 386 25693 420 25727
rect 386 25625 420 25659
rect 386 25557 420 25591
rect 386 25489 420 25523
rect 386 25421 420 25455
rect 386 25353 420 25387
rect 386 25285 420 25319
rect 386 25217 420 25251
rect 386 25149 420 25183
rect 386 25081 420 25115
rect 386 25013 420 25047
rect 386 24945 420 24979
rect 386 24877 420 24911
rect 386 24809 420 24843
rect 386 24741 420 24775
rect 386 24673 420 24707
rect 386 24605 420 24639
rect 386 24537 420 24571
rect 386 24469 420 24503
rect 386 24401 420 24435
rect 386 24333 420 24367
rect 386 24265 420 24299
rect 386 24197 420 24231
rect 386 24129 420 24163
rect 3036 26156 3070 26190
rect 3036 26088 3070 26122
rect 3036 26020 3070 26054
rect 3036 25952 3070 25986
rect 3036 25884 3070 25918
rect 3036 25816 3070 25850
rect 3036 25748 3070 25782
rect 3036 25680 3070 25714
rect 3036 25612 3070 25646
rect 3036 25544 3070 25578
rect 3036 25476 3070 25510
rect 3036 25408 3070 25442
rect 3036 25340 3070 25374
rect 3036 25272 3070 25306
rect 3036 25204 3070 25238
rect 3036 25136 3070 25170
rect 3036 25068 3070 25102
rect 3036 25000 3070 25034
rect 3036 24932 3070 24966
rect 3036 24864 3070 24898
rect 3036 24796 3070 24830
rect 3036 24728 3070 24762
rect 3036 24660 3070 24694
rect 3036 24592 3070 24626
rect 3036 24524 3070 24558
rect 3036 24456 3070 24490
rect 3036 24388 3070 24422
rect 3036 24320 3070 24354
rect 3036 24252 3070 24286
rect 3036 24184 3070 24218
rect 386 24061 420 24095
rect 3036 24116 3070 24150
rect 386 23993 420 24027
rect 386 23925 420 23959
rect 386 23857 420 23891
rect 386 23789 420 23823
rect 386 23721 420 23755
rect 386 23653 420 23687
rect 386 23585 420 23619
rect 386 23517 420 23551
rect 386 23449 420 23483
rect 386 23381 420 23415
rect 386 23313 420 23347
rect 386 23245 420 23279
rect 386 23177 420 23211
rect 386 23109 420 23143
rect 386 23041 420 23075
rect 386 22973 420 23007
rect 386 22905 420 22939
rect 386 22837 420 22871
rect 386 22769 420 22803
rect 386 22701 420 22735
rect 386 22633 420 22667
rect 386 22565 420 22599
rect 386 22497 420 22531
rect 386 22429 420 22463
rect 386 22361 420 22395
rect 386 22293 420 22327
rect 386 22225 420 22259
rect 386 22157 420 22191
rect 386 22089 420 22123
rect 386 22021 420 22055
rect 3036 24048 3070 24082
rect 3036 23980 3070 24014
rect 3036 23912 3070 23946
rect 3036 23844 3070 23878
rect 3036 23776 3070 23810
rect 3036 23708 3070 23742
rect 3036 23640 3070 23674
rect 3036 23572 3070 23606
rect 3036 23504 3070 23538
rect 3036 23436 3070 23470
rect 3036 23368 3070 23402
rect 3036 23300 3070 23334
rect 3036 23232 3070 23266
rect 3036 23164 3070 23198
rect 3036 23096 3070 23130
rect 3036 23028 3070 23062
rect 3036 22960 3070 22994
rect 3036 22892 3070 22926
rect 3036 22824 3070 22858
rect 3036 22756 3070 22790
rect 3036 22688 3070 22722
rect 3036 22620 3070 22654
rect 3036 22552 3070 22586
rect 3036 22484 3070 22518
rect 3036 22416 3070 22450
rect 3036 22348 3070 22382
rect 3036 22280 3070 22314
rect 3036 22212 3070 22246
rect 3036 22144 3070 22178
rect 3036 22076 3070 22110
rect 386 21953 420 21987
rect 3036 22008 3070 22042
rect 386 21885 420 21919
rect 386 21817 420 21851
rect 386 21749 420 21783
rect 386 21681 420 21715
rect 386 21613 420 21647
rect 386 21545 420 21579
rect 386 21477 420 21511
rect 386 21409 420 21443
rect 386 21341 420 21375
rect 386 21273 420 21307
rect 386 21205 420 21239
rect 386 21137 420 21171
rect 386 21069 420 21103
rect 386 21001 420 21035
rect 386 20933 420 20967
rect 386 20865 420 20899
rect 386 20797 420 20831
rect 386 20729 420 20763
rect 386 20661 420 20695
rect 386 20593 420 20627
rect 386 20525 420 20559
rect 386 20457 420 20491
rect 386 20389 420 20423
rect 386 20321 420 20355
rect 386 20253 420 20287
rect 386 20185 420 20219
rect 386 20117 420 20151
rect 386 20049 420 20083
rect 386 19981 420 20015
rect 386 19913 420 19947
rect 3036 21940 3070 21974
rect 3036 21872 3070 21906
rect 3036 21804 3070 21838
rect 3036 21736 3070 21770
rect 3036 21668 3070 21702
rect 3036 21600 3070 21634
rect 3036 21532 3070 21566
rect 3036 21464 3070 21498
rect 3036 21396 3070 21430
rect 3036 21328 3070 21362
rect 3036 21260 3070 21294
rect 3036 21192 3070 21226
rect 3036 21124 3070 21158
rect 3036 21056 3070 21090
rect 3036 20988 3070 21022
rect 3036 20920 3070 20954
rect 3036 20852 3070 20886
rect 3036 20784 3070 20818
rect 3036 20716 3070 20750
rect 3036 20648 3070 20682
rect 3036 20580 3070 20614
rect 3036 20512 3070 20546
rect 3036 20444 3070 20478
rect 3036 20376 3070 20410
rect 3036 20308 3070 20342
rect 3036 20240 3070 20274
rect 3036 20172 3070 20206
rect 3036 20104 3070 20138
rect 3036 20036 3070 20070
rect 3036 19968 3070 20002
rect 3036 19900 3070 19934
rect 386 19845 420 19879
rect 386 19777 420 19811
rect 386 19709 420 19743
rect 386 19641 420 19675
rect 386 19573 420 19607
rect 386 19505 420 19539
rect 386 19437 420 19471
rect 386 19369 420 19403
rect 386 19301 420 19335
rect 386 19233 420 19267
rect 386 19165 420 19199
rect 386 19097 420 19131
rect 386 19029 420 19063
rect 386 18961 420 18995
rect 386 18893 420 18927
rect 386 18825 420 18859
rect 386 18757 420 18791
rect 386 18689 420 18723
rect 386 18621 420 18655
rect 386 18553 420 18587
rect 386 18485 420 18519
rect 386 18417 420 18451
rect 386 18349 420 18383
rect 386 18281 420 18315
rect 386 18213 420 18247
rect 386 18145 420 18179
rect 386 18077 420 18111
rect 386 18009 420 18043
rect 386 17941 420 17975
rect 386 17873 420 17907
rect 386 17805 420 17839
rect 386 17737 420 17771
rect 3036 19832 3070 19866
rect 3036 19764 3070 19798
rect 3036 19696 3070 19730
rect 3036 19628 3070 19662
rect 3036 19560 3070 19594
rect 3036 19492 3070 19526
rect 3036 19424 3070 19458
rect 3036 19356 3070 19390
rect 3036 19288 3070 19322
rect 3036 19220 3070 19254
rect 3036 19152 3070 19186
rect 3036 19084 3070 19118
rect 3036 19016 3070 19050
rect 3036 18948 3070 18982
rect 3036 18880 3070 18914
rect 3036 18812 3070 18846
rect 3036 18744 3070 18778
rect 3036 18676 3070 18710
rect 3036 18608 3070 18642
rect 3036 18540 3070 18574
rect 3036 18472 3070 18506
rect 3036 18404 3070 18438
rect 3036 18336 3070 18370
rect 3036 18268 3070 18302
rect 3036 18200 3070 18234
rect 3036 18132 3070 18166
rect 3036 18064 3070 18098
rect 3036 17996 3070 18030
rect 3036 17928 3070 17962
rect 3036 17860 3070 17894
rect 3036 17792 3070 17826
rect 3036 17724 3070 17758
rect 386 17669 420 17703
rect 386 17601 420 17635
rect 386 17533 420 17567
rect 386 17465 420 17499
rect 386 17397 420 17431
rect 386 17329 420 17363
rect 386 17261 420 17295
rect 386 17193 420 17227
rect 386 17125 420 17159
rect 386 17057 420 17091
rect 386 16989 420 17023
rect 386 16921 420 16955
rect 386 16853 420 16887
rect 386 16785 420 16819
rect 386 16717 420 16751
rect 386 16649 420 16683
rect 386 16581 420 16615
rect 386 16513 420 16547
rect 386 16445 420 16479
rect 386 16377 420 16411
rect 386 16309 420 16343
rect 386 16241 420 16275
rect 386 16173 420 16207
rect 386 16105 420 16139
rect 386 16037 420 16071
rect 386 15969 420 16003
rect 386 15901 420 15935
rect 386 15833 420 15867
rect 386 15765 420 15799
rect 386 15697 420 15731
rect 386 15629 420 15663
rect 3036 17656 3070 17690
rect 3036 17588 3070 17622
rect 3036 17520 3070 17554
rect 3036 17452 3070 17486
rect 3036 17384 3070 17418
rect 3036 17316 3070 17350
rect 3036 17248 3070 17282
rect 3036 17180 3070 17214
rect 3036 17112 3070 17146
rect 3036 17044 3070 17078
rect 3036 16976 3070 17010
rect 3036 16908 3070 16942
rect 3036 16840 3070 16874
rect 3036 16772 3070 16806
rect 3036 16704 3070 16738
rect 3036 16636 3070 16670
rect 3036 16568 3070 16602
rect 3036 16500 3070 16534
rect 3036 16432 3070 16466
rect 3036 16364 3070 16398
rect 3036 16296 3070 16330
rect 3036 16228 3070 16262
rect 3036 16160 3070 16194
rect 3036 16092 3070 16126
rect 3036 16024 3070 16058
rect 3036 15956 3070 15990
rect 3036 15888 3070 15922
rect 3036 15820 3070 15854
rect 3036 15752 3070 15786
rect 3036 15684 3070 15718
rect 386 15561 420 15595
rect 3036 15616 3070 15650
rect 386 15493 420 15527
rect 386 15425 420 15459
rect 386 15357 420 15391
rect 386 15289 420 15323
rect 386 15221 420 15255
rect 386 15153 420 15187
rect 386 15085 420 15119
rect 386 15017 420 15051
rect 386 14949 420 14983
rect 386 14881 420 14915
rect 386 14813 420 14847
rect 386 14745 420 14779
rect 386 14677 420 14711
rect 386 14609 420 14643
rect 386 14541 420 14575
rect 386 14473 420 14507
rect 386 14405 420 14439
rect 386 14337 420 14371
rect 386 14269 420 14303
rect 386 14201 420 14235
rect 386 14133 420 14167
rect 386 14065 420 14099
rect 386 13997 420 14031
rect 386 13929 420 13963
rect 386 13861 420 13895
rect 386 13793 420 13827
rect 386 13725 420 13759
rect 386 13657 420 13691
rect 386 13589 420 13623
rect 386 13521 420 13555
rect 3036 15548 3070 15582
rect 3036 15480 3070 15514
rect 3036 15412 3070 15446
rect 3036 15344 3070 15378
rect 3036 15276 3070 15310
rect 3036 15208 3070 15242
rect 3036 15140 3070 15174
rect 3036 15072 3070 15106
rect 3036 15004 3070 15038
rect 3036 14936 3070 14970
rect 3036 14868 3070 14902
rect 3036 14800 3070 14834
rect 3036 14732 3070 14766
rect 3036 14664 3070 14698
rect 3036 14596 3070 14630
rect 3036 14528 3070 14562
rect 3036 14460 3070 14494
rect 3036 14392 3070 14426
rect 3036 14324 3070 14358
rect 3036 14256 3070 14290
rect 3036 14188 3070 14222
rect 3036 14120 3070 14154
rect 3036 14052 3070 14086
rect 3036 13984 3070 14018
rect 3036 13916 3070 13950
rect 3036 13848 3070 13882
rect 3036 13780 3070 13814
rect 3036 13712 3070 13746
rect 3036 13644 3070 13678
rect 3036 13576 3070 13610
rect 386 13453 420 13487
rect 3036 13508 3070 13542
rect 386 13385 420 13419
rect 386 13317 420 13351
rect 386 13249 420 13283
rect 386 13181 420 13215
rect 386 13113 420 13147
rect 386 13045 420 13079
rect 386 12977 420 13011
rect 386 12909 420 12943
rect 386 12841 420 12875
rect 386 12773 420 12807
rect 386 12705 420 12739
rect 386 12637 420 12671
rect 386 12569 420 12603
rect 386 12501 420 12535
rect 386 12433 420 12467
rect 386 12365 420 12399
rect 386 12297 420 12331
rect 386 12229 420 12263
rect 386 12161 420 12195
rect 386 12093 420 12127
rect 386 12025 420 12059
rect 386 11957 420 11991
rect 386 11889 420 11923
rect 386 11821 420 11855
rect 386 11753 420 11787
rect 386 11685 420 11719
rect 386 11617 420 11651
rect 386 11549 420 11583
rect 386 11481 420 11515
rect 386 11413 420 11447
rect 3036 13440 3070 13474
rect 3036 13372 3070 13406
rect 3036 13304 3070 13338
rect 3036 13236 3070 13270
rect 3036 13168 3070 13202
rect 3036 13100 3070 13134
rect 3036 13032 3070 13066
rect 3036 12964 3070 12998
rect 3036 12896 3070 12930
rect 3036 12828 3070 12862
rect 3036 12760 3070 12794
rect 3036 12692 3070 12726
rect 3036 12624 3070 12658
rect 3036 12556 3070 12590
rect 3036 12488 3070 12522
rect 3036 12420 3070 12454
rect 3036 12352 3070 12386
rect 3036 12284 3070 12318
rect 3036 12216 3070 12250
rect 3036 12148 3070 12182
rect 3036 12080 3070 12114
rect 3036 12012 3070 12046
rect 3036 11944 3070 11978
rect 3036 11876 3070 11910
rect 3036 11808 3070 11842
rect 3036 11740 3070 11774
rect 3036 11672 3070 11706
rect 3036 11604 3070 11638
rect 3036 11536 3070 11570
rect 3036 11468 3070 11502
rect 3036 11400 3070 11434
rect 386 11345 420 11379
rect 3036 11332 3070 11366
rect 386 11277 420 11311
rect 386 11209 420 11243
rect 386 11141 420 11175
rect 386 11073 420 11107
rect 386 11005 420 11039
rect 386 10937 420 10971
rect 386 10869 420 10903
rect 386 10801 420 10835
rect 386 10733 420 10767
rect 386 10665 420 10699
rect 386 10597 420 10631
rect 386 10529 420 10563
rect 386 10461 420 10495
rect 386 10393 420 10427
rect 386 10325 420 10359
rect 386 10257 420 10291
rect 386 10189 420 10223
rect 386 10121 420 10155
rect 386 10053 420 10087
rect 386 9985 420 10019
rect 386 9917 420 9951
rect 386 9849 420 9883
rect 386 9781 420 9815
rect 386 9713 420 9747
rect 386 9645 420 9679
rect 386 9577 420 9611
rect 386 9509 420 9543
rect 386 9441 420 9475
rect 386 9373 420 9407
rect 386 9305 420 9339
rect 386 9237 420 9271
rect 3036 11264 3070 11298
rect 3036 11196 3070 11230
rect 3036 11128 3070 11162
rect 3036 11060 3070 11094
rect 3036 10992 3070 11026
rect 3036 10924 3070 10958
rect 3036 10856 3070 10890
rect 3036 10788 3070 10822
rect 3036 10720 3070 10754
rect 3036 10652 3070 10686
rect 3036 10584 3070 10618
rect 3036 10516 3070 10550
rect 3036 10448 3070 10482
rect 3036 10380 3070 10414
rect 3036 10312 3070 10346
rect 3036 10244 3070 10278
rect 3036 10176 3070 10210
rect 3036 10108 3070 10142
rect 3036 10040 3070 10074
rect 3036 9972 3070 10006
rect 3036 9904 3070 9938
rect 3036 9836 3070 9870
rect 3036 9768 3070 9802
rect 3036 9700 3070 9734
rect 3036 9632 3070 9666
rect 3036 9564 3070 9598
rect 3036 9496 3070 9530
rect 3036 9428 3070 9462
rect 3036 9360 3070 9394
rect 3036 9292 3070 9326
rect 386 9169 420 9203
rect 3036 9224 3070 9258
rect 386 9101 420 9135
rect 386 9033 420 9067
rect 386 8965 420 8999
rect 386 8897 420 8931
rect 386 8829 420 8863
rect 386 8761 420 8795
rect 386 8693 420 8727
rect 386 8625 420 8659
rect 386 8557 420 8591
rect 386 8489 420 8523
rect 386 8421 420 8455
rect 386 8353 420 8387
rect 386 8285 420 8319
rect 386 8217 420 8251
rect 386 8149 420 8183
rect 386 8081 420 8115
rect 386 8013 420 8047
rect 386 7945 420 7979
rect 386 7877 420 7911
rect 386 7809 420 7843
rect 386 7741 420 7775
rect 386 7673 420 7707
rect 386 7605 420 7639
rect 386 7537 420 7571
rect 386 7469 420 7503
rect 386 7401 420 7435
rect 386 7333 420 7367
rect 386 7265 420 7299
rect 386 7197 420 7231
rect 386 7129 420 7163
rect 3036 9156 3070 9190
rect 3036 9088 3070 9122
rect 3036 9020 3070 9054
rect 3036 8952 3070 8986
rect 3036 8884 3070 8918
rect 3036 8816 3070 8850
rect 3036 8748 3070 8782
rect 3036 8680 3070 8714
rect 3036 8612 3070 8646
rect 3036 8544 3070 8578
rect 3036 8476 3070 8510
rect 3036 8408 3070 8442
rect 3036 8340 3070 8374
rect 3036 8272 3070 8306
rect 3036 8204 3070 8238
rect 3036 8136 3070 8170
rect 3036 8068 3070 8102
rect 3036 8000 3070 8034
rect 3036 7932 3070 7966
rect 3036 7864 3070 7898
rect 3036 7796 3070 7830
rect 3036 7728 3070 7762
rect 3036 7660 3070 7694
rect 3036 7592 3070 7626
rect 3036 7524 3070 7558
rect 3036 7456 3070 7490
rect 3036 7388 3070 7422
rect 3036 7320 3070 7354
rect 3036 7252 3070 7286
rect 3036 7184 3070 7218
rect 386 7061 420 7095
rect 3036 7116 3070 7150
rect 386 6993 420 7027
rect 386 6925 420 6959
rect 386 6857 420 6891
rect 386 6789 420 6823
rect 386 6721 420 6755
rect 386 6653 420 6687
rect 386 6585 420 6619
rect 386 6517 420 6551
rect 386 6449 420 6483
rect 386 6381 420 6415
rect 386 6313 420 6347
rect 386 6245 420 6279
rect 386 6177 420 6211
rect 386 6109 420 6143
rect 386 6041 420 6075
rect 386 5973 420 6007
rect 386 5905 420 5939
rect 386 5837 420 5871
rect 386 5769 420 5803
rect 386 5701 420 5735
rect 386 5633 420 5667
rect 386 5565 420 5599
rect 386 5497 420 5531
rect 386 5429 420 5463
rect 386 5361 420 5395
rect 386 5293 420 5327
rect 386 5225 420 5259
rect 386 5157 420 5191
rect 386 5089 420 5123
rect 386 5021 420 5055
rect 3036 7048 3070 7082
rect 3036 6980 3070 7014
rect 3036 6912 3070 6946
rect 3036 6844 3070 6878
rect 3036 6776 3070 6810
rect 3036 6708 3070 6742
rect 3036 6640 3070 6674
rect 3036 6572 3070 6606
rect 3036 6504 3070 6538
rect 3036 6436 3070 6470
rect 3036 6368 3070 6402
rect 3036 6300 3070 6334
rect 3036 6232 3070 6266
rect 3036 6164 3070 6198
rect 3036 6096 3070 6130
rect 3036 6028 3070 6062
rect 3036 5960 3070 5994
rect 3036 5892 3070 5926
rect 3036 5824 3070 5858
rect 3036 5756 3070 5790
rect 3036 5688 3070 5722
rect 3036 5620 3070 5654
rect 3036 5552 3070 5586
rect 3036 5484 3070 5518
rect 3036 5416 3070 5450
rect 3036 5348 3070 5382
rect 3036 5280 3070 5314
rect 3036 5212 3070 5246
rect 3036 5144 3070 5178
rect 3036 5076 3070 5110
rect 3036 5008 3070 5042
rect 386 4953 420 4987
rect 3036 4940 3070 4974
rect 386 4885 420 4919
rect 386 4817 420 4851
rect 386 4749 420 4783
rect 386 4681 420 4715
rect 386 4613 420 4647
rect 386 4545 420 4579
rect 386 4477 420 4511
rect 386 4409 420 4443
rect 386 4341 420 4375
rect 386 4273 420 4307
rect 386 4205 420 4239
rect 386 4137 420 4171
rect 386 4069 420 4103
rect 386 4001 420 4035
rect 386 3933 420 3967
rect 386 3865 420 3899
rect 386 3797 420 3831
rect 386 3729 420 3763
rect 386 3661 420 3695
rect 386 3593 420 3627
rect 386 3525 420 3559
rect 386 3457 420 3491
rect 386 3389 420 3423
rect 386 3321 420 3355
rect 386 3253 420 3287
rect 386 3185 420 3219
rect 386 3117 420 3151
rect 386 3049 420 3083
rect 386 2981 420 3015
rect 386 2913 420 2947
rect 386 2845 420 2879
rect 3036 4872 3070 4906
rect 3036 4804 3070 4838
rect 3036 4736 3070 4770
rect 3036 4668 3070 4702
rect 3036 4600 3070 4634
rect 3036 4532 3070 4566
rect 3036 4464 3070 4498
rect 3036 4396 3070 4430
rect 3036 4328 3070 4362
rect 3036 4260 3070 4294
rect 3036 4192 3070 4226
rect 3036 4124 3070 4158
rect 3036 4056 3070 4090
rect 3036 3988 3070 4022
rect 3036 3920 3070 3954
rect 3036 3852 3070 3886
rect 3036 3784 3070 3818
rect 3036 3716 3070 3750
rect 3036 3648 3070 3682
rect 3036 3580 3070 3614
rect 3036 3512 3070 3546
rect 3036 3444 3070 3478
rect 3036 3376 3070 3410
rect 3036 3308 3070 3342
rect 3036 3240 3070 3274
rect 3036 3172 3070 3206
rect 3036 3104 3070 3138
rect 3036 3036 3070 3070
rect 3036 2968 3070 3002
rect 3036 2900 3070 2934
rect 386 2777 420 2811
rect 3036 2832 3070 2866
rect 386 2709 420 2743
rect 386 2641 420 2675
rect 386 2573 420 2607
rect 386 2505 420 2539
rect 386 2437 420 2471
rect 386 2369 420 2403
rect 386 2301 420 2335
rect 386 2233 420 2267
rect 386 2165 420 2199
rect 386 2097 420 2131
rect 386 2029 420 2063
rect 386 1961 420 1995
rect 386 1893 420 1927
rect 386 1825 420 1859
rect 386 1757 420 1791
rect 386 1689 420 1723
rect 386 1621 420 1655
rect 386 1553 420 1587
rect 386 1485 420 1519
rect 386 1417 420 1451
rect 386 1349 420 1383
rect 386 1281 420 1315
rect 386 1213 420 1247
rect 386 1145 420 1179
rect 386 1077 420 1111
rect 386 1009 420 1043
rect 386 941 420 975
rect 386 873 420 907
rect 386 805 420 839
rect 386 737 420 771
rect 3036 2764 3070 2798
rect 3036 2696 3070 2730
rect 3036 2628 3070 2662
rect 3036 2560 3070 2594
rect 3036 2492 3070 2526
rect 3036 2424 3070 2458
rect 3036 2356 3070 2390
rect 3036 2288 3070 2322
rect 3036 2220 3070 2254
rect 3036 2152 3070 2186
rect 3036 2084 3070 2118
rect 3036 2016 3070 2050
rect 3036 1948 3070 1982
rect 3036 1880 3070 1914
rect 3036 1812 3070 1846
rect 3036 1744 3070 1778
rect 3036 1676 3070 1710
rect 3036 1608 3070 1642
rect 3036 1540 3070 1574
rect 3036 1472 3070 1506
rect 3036 1404 3070 1438
rect 3036 1336 3070 1370
rect 3036 1268 3070 1302
rect 3036 1200 3070 1234
rect 3036 1132 3070 1166
rect 3036 1064 3070 1098
rect 3036 996 3070 1030
rect 3036 928 3070 962
rect 3036 860 3070 894
rect 3036 792 3070 826
rect 386 669 420 703
rect 3036 724 3070 758
rect 3036 656 3070 690
rect 3036 588 3070 622
rect 441 533 475 567
rect 509 533 543 567
rect 577 533 611 567
rect 645 533 679 567
rect 713 533 747 567
rect 781 533 815 567
rect 849 533 883 567
rect 917 533 951 567
rect 985 533 1019 567
rect 1053 533 1087 567
rect 1121 533 1155 567
rect 1189 533 1223 567
rect 1257 533 1291 567
rect 1325 533 1359 567
rect 1393 533 1427 567
rect 1461 533 1495 567
rect 1529 533 1563 567
rect 1597 533 1631 567
rect 1665 533 1699 567
rect 1733 533 1767 567
rect 1801 533 1835 567
rect 1869 533 1903 567
rect 1937 533 1971 567
rect 2005 533 2039 567
rect 2073 533 2107 567
rect 2141 533 2175 567
rect 2209 533 2243 567
rect 2277 533 2311 567
rect 2345 533 2379 567
rect 2413 533 2447 567
rect 2481 533 2515 567
rect 2549 533 2583 567
rect 2617 533 2651 567
rect 2685 533 2719 567
rect 2753 533 2787 567
rect 2821 533 2855 567
rect 2889 533 2923 567
rect 2957 533 2991 567
<< mvnsubdiffcont >>
rect 236 39840 270 39874
rect 304 39840 338 39874
rect 372 39840 406 39874
rect 440 39840 474 39874
rect 508 39840 542 39874
rect 576 39840 610 39874
rect 644 39840 678 39874
rect 712 39840 746 39874
rect 780 39840 814 39874
rect 848 39840 882 39874
rect 916 39840 950 39874
rect 984 39840 1018 39874
rect 1052 39840 1086 39874
rect 1120 39840 1154 39874
rect 1188 39840 1222 39874
rect 1256 39840 1290 39874
rect 1324 39840 1358 39874
rect 1392 39840 1426 39874
rect 1460 39840 1494 39874
rect 1528 39840 1562 39874
rect 1596 39840 1630 39874
rect 1664 39840 1698 39874
rect 1732 39840 1766 39874
rect 1800 39840 1834 39874
rect 1868 39840 1902 39874
rect 1936 39840 1970 39874
rect 2004 39840 2038 39874
rect 2072 39840 2106 39874
rect 2140 39840 2174 39874
rect 2208 39840 2242 39874
rect 2276 39840 2310 39874
rect 2344 39840 2378 39874
rect 2412 39840 2446 39874
rect 2480 39840 2514 39874
rect 2548 39840 2582 39874
rect 2616 39840 2650 39874
rect 2684 39840 2718 39874
rect 2752 39840 2786 39874
rect 2820 39840 2854 39874
rect 2888 39840 2922 39874
rect 2956 39840 2990 39874
rect 3024 39840 3058 39874
rect 3092 39840 3126 39874
rect 3160 39840 3194 39874
rect 3228 39840 3262 39874
rect 126 39772 160 39806
rect 126 39704 160 39738
rect 126 39636 160 39670
rect 126 39568 160 39602
rect 126 39500 160 39534
rect 126 39432 160 39466
rect 126 39364 160 39398
rect 126 39296 160 39330
rect 126 39228 160 39262
rect 126 39160 160 39194
rect 3296 39770 3330 39804
rect 3296 39702 3330 39736
rect 3296 39634 3330 39668
rect 3296 39566 3330 39600
rect 3296 39498 3330 39532
rect 3296 39430 3330 39464
rect 3296 39362 3330 39396
rect 3296 39294 3330 39328
rect 3296 39226 3330 39260
rect 126 39092 160 39126
rect 126 39024 160 39058
rect 126 38956 160 38990
rect 126 38888 160 38922
rect 126 38820 160 38854
rect 126 38752 160 38786
rect 126 38684 160 38718
rect 126 38616 160 38650
rect 126 38548 160 38582
rect 126 38480 160 38514
rect 126 38412 160 38446
rect 126 38344 160 38378
rect 126 38276 160 38310
rect 126 38208 160 38242
rect 126 38140 160 38174
rect 126 38072 160 38106
rect 126 38004 160 38038
rect 126 37936 160 37970
rect 126 37868 160 37902
rect 126 37800 160 37834
rect 126 37732 160 37766
rect 126 37664 160 37698
rect 126 37596 160 37630
rect 126 37528 160 37562
rect 126 37460 160 37494
rect 126 37392 160 37426
rect 126 37324 160 37358
rect 126 37256 160 37290
rect 126 37188 160 37222
rect 126 37120 160 37154
rect 126 37052 160 37086
rect 126 36984 160 37018
rect 126 36916 160 36950
rect 126 36848 160 36882
rect 126 36780 160 36814
rect 126 36712 160 36746
rect 126 36644 160 36678
rect 126 36576 160 36610
rect 126 36508 160 36542
rect 126 36440 160 36474
rect 126 36372 160 36406
rect 126 36304 160 36338
rect 126 36236 160 36270
rect 126 36168 160 36202
rect 126 36100 160 36134
rect 126 36032 160 36066
rect 126 35964 160 35998
rect 126 35896 160 35930
rect 126 35828 160 35862
rect 126 35760 160 35794
rect 126 35692 160 35726
rect 126 35624 160 35658
rect 126 35556 160 35590
rect 126 35488 160 35522
rect 126 35420 160 35454
rect 126 35352 160 35386
rect 126 35284 160 35318
rect 126 35216 160 35250
rect 126 35148 160 35182
rect 126 35080 160 35114
rect 126 35012 160 35046
rect 126 34944 160 34978
rect 126 34876 160 34910
rect 126 34808 160 34842
rect 126 34740 160 34774
rect 126 34672 160 34706
rect 126 34604 160 34638
rect 126 34536 160 34570
rect 126 34468 160 34502
rect 126 34400 160 34434
rect 126 34332 160 34366
rect 126 34264 160 34298
rect 126 34196 160 34230
rect 126 34128 160 34162
rect 126 34060 160 34094
rect 126 33992 160 34026
rect 126 33924 160 33958
rect 126 33856 160 33890
rect 126 33788 160 33822
rect 126 33720 160 33754
rect 126 33652 160 33686
rect 126 33584 160 33618
rect 126 33516 160 33550
rect 126 33448 160 33482
rect 126 33380 160 33414
rect 126 33312 160 33346
rect 126 33244 160 33278
rect 126 33176 160 33210
rect 126 33108 160 33142
rect 126 33040 160 33074
rect 126 32972 160 33006
rect 126 32904 160 32938
rect 126 32836 160 32870
rect 126 32768 160 32802
rect 126 32700 160 32734
rect 126 32632 160 32666
rect 126 32564 160 32598
rect 126 32496 160 32530
rect 126 32428 160 32462
rect 126 32360 160 32394
rect 126 32292 160 32326
rect 126 32224 160 32258
rect 126 32156 160 32190
rect 126 32088 160 32122
rect 126 32020 160 32054
rect 126 31952 160 31986
rect 126 31884 160 31918
rect 126 31816 160 31850
rect 126 31748 160 31782
rect 126 31680 160 31714
rect 126 31612 160 31646
rect 126 31544 160 31578
rect 126 31476 160 31510
rect 126 31408 160 31442
rect 126 31340 160 31374
rect 126 31272 160 31306
rect 126 31204 160 31238
rect 126 31136 160 31170
rect 126 31068 160 31102
rect 126 31000 160 31034
rect 126 30932 160 30966
rect 126 30864 160 30898
rect 126 30796 160 30830
rect 126 30728 160 30762
rect 126 30660 160 30694
rect 126 30592 160 30626
rect 126 30524 160 30558
rect 126 30456 160 30490
rect 126 30388 160 30422
rect 126 30320 160 30354
rect 126 30252 160 30286
rect 126 30184 160 30218
rect 126 30116 160 30150
rect 126 30048 160 30082
rect 126 29980 160 30014
rect 126 29912 160 29946
rect 126 29844 160 29878
rect 126 29776 160 29810
rect 126 29708 160 29742
rect 126 29640 160 29674
rect 126 29572 160 29606
rect 126 29504 160 29538
rect 126 29436 160 29470
rect 126 29368 160 29402
rect 126 29300 160 29334
rect 126 29232 160 29266
rect 126 29164 160 29198
rect 126 29096 160 29130
rect 126 29028 160 29062
rect 126 28960 160 28994
rect 126 28892 160 28926
rect 126 28824 160 28858
rect 126 28756 160 28790
rect 126 28688 160 28722
rect 126 28620 160 28654
rect 126 28552 160 28586
rect 126 28484 160 28518
rect 126 28416 160 28450
rect 126 28348 160 28382
rect 126 28280 160 28314
rect 126 28212 160 28246
rect 126 28144 160 28178
rect 126 28076 160 28110
rect 126 28008 160 28042
rect 126 27940 160 27974
rect 126 27872 160 27906
rect 126 27804 160 27838
rect 126 27736 160 27770
rect 126 27668 160 27702
rect 126 27600 160 27634
rect 126 27532 160 27566
rect 126 27464 160 27498
rect 126 27396 160 27430
rect 126 27328 160 27362
rect 126 27260 160 27294
rect 126 27192 160 27226
rect 126 27124 160 27158
rect 126 27056 160 27090
rect 126 26988 160 27022
rect 126 26920 160 26954
rect 126 26852 160 26886
rect 126 26784 160 26818
rect 126 26716 160 26750
rect 126 26648 160 26682
rect 126 26580 160 26614
rect 126 26512 160 26546
rect 126 26444 160 26478
rect 126 26376 160 26410
rect 126 26308 160 26342
rect 126 26240 160 26274
rect 126 26172 160 26206
rect 126 26104 160 26138
rect 126 26036 160 26070
rect 126 25968 160 26002
rect 126 25900 160 25934
rect 126 25832 160 25866
rect 126 25764 160 25798
rect 126 25696 160 25730
rect 126 25628 160 25662
rect 126 25560 160 25594
rect 126 25492 160 25526
rect 126 25424 160 25458
rect 126 25356 160 25390
rect 126 25288 160 25322
rect 126 25220 160 25254
rect 126 25152 160 25186
rect 126 25084 160 25118
rect 126 25016 160 25050
rect 126 24948 160 24982
rect 126 24880 160 24914
rect 126 24812 160 24846
rect 126 24744 160 24778
rect 126 24676 160 24710
rect 126 24608 160 24642
rect 126 24540 160 24574
rect 126 24472 160 24506
rect 126 24404 160 24438
rect 126 24336 160 24370
rect 126 24268 160 24302
rect 126 24200 160 24234
rect 126 24132 160 24166
rect 126 24064 160 24098
rect 126 23996 160 24030
rect 126 23928 160 23962
rect 126 23860 160 23894
rect 126 23792 160 23826
rect 126 23724 160 23758
rect 126 23656 160 23690
rect 126 23588 160 23622
rect 126 23520 160 23554
rect 126 23452 160 23486
rect 126 23384 160 23418
rect 126 23316 160 23350
rect 126 23248 160 23282
rect 126 23180 160 23214
rect 126 23112 160 23146
rect 126 23044 160 23078
rect 126 22976 160 23010
rect 126 22908 160 22942
rect 126 22840 160 22874
rect 126 22772 160 22806
rect 126 22704 160 22738
rect 126 22636 160 22670
rect 126 22568 160 22602
rect 126 22500 160 22534
rect 126 22432 160 22466
rect 126 22364 160 22398
rect 126 22296 160 22330
rect 126 22228 160 22262
rect 126 22160 160 22194
rect 126 22092 160 22126
rect 126 22024 160 22058
rect 126 21956 160 21990
rect 126 21888 160 21922
rect 126 21820 160 21854
rect 126 21752 160 21786
rect 126 21684 160 21718
rect 126 21616 160 21650
rect 126 21548 160 21582
rect 126 21480 160 21514
rect 126 21412 160 21446
rect 126 21344 160 21378
rect 126 21276 160 21310
rect 126 21208 160 21242
rect 126 21140 160 21174
rect 126 21072 160 21106
rect 126 21004 160 21038
rect 126 20936 160 20970
rect 126 20868 160 20902
rect 126 20800 160 20834
rect 126 20732 160 20766
rect 126 20664 160 20698
rect 126 20596 160 20630
rect 126 20528 160 20562
rect 126 20460 160 20494
rect 126 20392 160 20426
rect 126 20324 160 20358
rect 126 20256 160 20290
rect 126 20188 160 20222
rect 126 20120 160 20154
rect 126 20052 160 20086
rect 126 19984 160 20018
rect 126 19916 160 19950
rect 126 19848 160 19882
rect 126 19780 160 19814
rect 126 19712 160 19746
rect 126 19644 160 19678
rect 126 19576 160 19610
rect 126 19508 160 19542
rect 126 19440 160 19474
rect 126 19372 160 19406
rect 126 19304 160 19338
rect 126 19236 160 19270
rect 126 19168 160 19202
rect 126 19100 160 19134
rect 126 19032 160 19066
rect 126 18964 160 18998
rect 126 18896 160 18930
rect 126 18828 160 18862
rect 126 18760 160 18794
rect 126 18692 160 18726
rect 126 18624 160 18658
rect 126 18556 160 18590
rect 126 18488 160 18522
rect 126 18420 160 18454
rect 126 18352 160 18386
rect 126 18284 160 18318
rect 126 18216 160 18250
rect 126 18148 160 18182
rect 126 18080 160 18114
rect 126 18012 160 18046
rect 126 17944 160 17978
rect 126 17876 160 17910
rect 126 17808 160 17842
rect 126 17740 160 17774
rect 126 17672 160 17706
rect 126 17604 160 17638
rect 126 17536 160 17570
rect 126 17468 160 17502
rect 126 17400 160 17434
rect 126 17332 160 17366
rect 126 17264 160 17298
rect 126 17196 160 17230
rect 126 17128 160 17162
rect 126 17060 160 17094
rect 126 16992 160 17026
rect 126 16924 160 16958
rect 126 16856 160 16890
rect 126 16788 160 16822
rect 126 16720 160 16754
rect 126 16652 160 16686
rect 126 16584 160 16618
rect 126 16516 160 16550
rect 126 16448 160 16482
rect 126 16380 160 16414
rect 126 16312 160 16346
rect 126 16244 160 16278
rect 126 16176 160 16210
rect 126 16108 160 16142
rect 126 16040 160 16074
rect 126 15972 160 16006
rect 126 15904 160 15938
rect 126 15836 160 15870
rect 126 15768 160 15802
rect 126 15700 160 15734
rect 126 15632 160 15666
rect 126 15564 160 15598
rect 126 15496 160 15530
rect 126 15428 160 15462
rect 126 15360 160 15394
rect 126 15292 160 15326
rect 126 15224 160 15258
rect 126 15156 160 15190
rect 126 15088 160 15122
rect 126 15020 160 15054
rect 126 14952 160 14986
rect 126 14884 160 14918
rect 126 14816 160 14850
rect 126 14748 160 14782
rect 126 14680 160 14714
rect 126 14612 160 14646
rect 126 14544 160 14578
rect 126 14476 160 14510
rect 126 14408 160 14442
rect 126 14340 160 14374
rect 126 14272 160 14306
rect 126 14204 160 14238
rect 126 14136 160 14170
rect 126 14068 160 14102
rect 126 14000 160 14034
rect 126 13932 160 13966
rect 126 13864 160 13898
rect 126 13796 160 13830
rect 126 13728 160 13762
rect 126 13660 160 13694
rect 126 13592 160 13626
rect 126 13524 160 13558
rect 126 13456 160 13490
rect 126 13388 160 13422
rect 126 13320 160 13354
rect 126 13252 160 13286
rect 126 13184 160 13218
rect 126 13116 160 13150
rect 126 13048 160 13082
rect 126 12980 160 13014
rect 126 12912 160 12946
rect 126 12844 160 12878
rect 126 12776 160 12810
rect 126 12708 160 12742
rect 126 12640 160 12674
rect 126 12572 160 12606
rect 126 12504 160 12538
rect 126 12436 160 12470
rect 126 12368 160 12402
rect 126 12300 160 12334
rect 126 12232 160 12266
rect 126 12164 160 12198
rect 126 12096 160 12130
rect 126 12028 160 12062
rect 126 11960 160 11994
rect 126 11892 160 11926
rect 126 11824 160 11858
rect 126 11756 160 11790
rect 126 11688 160 11722
rect 126 11620 160 11654
rect 126 11552 160 11586
rect 126 11484 160 11518
rect 126 11416 160 11450
rect 126 11348 160 11382
rect 126 11280 160 11314
rect 126 11212 160 11246
rect 126 11144 160 11178
rect 126 11076 160 11110
rect 126 11008 160 11042
rect 126 10940 160 10974
rect 126 10872 160 10906
rect 126 10804 160 10838
rect 126 10736 160 10770
rect 126 10668 160 10702
rect 126 10600 160 10634
rect 126 10532 160 10566
rect 126 10464 160 10498
rect 126 10396 160 10430
rect 126 10328 160 10362
rect 126 10260 160 10294
rect 126 10192 160 10226
rect 126 10124 160 10158
rect 126 10056 160 10090
rect 126 9988 160 10022
rect 126 9920 160 9954
rect 126 9852 160 9886
rect 126 9784 160 9818
rect 126 9716 160 9750
rect 126 9648 160 9682
rect 126 9580 160 9614
rect 126 9512 160 9546
rect 126 9444 160 9478
rect 126 9376 160 9410
rect 126 9308 160 9342
rect 126 9240 160 9274
rect 126 9172 160 9206
rect 126 9104 160 9138
rect 126 9036 160 9070
rect 126 8968 160 9002
rect 126 8900 160 8934
rect 126 8832 160 8866
rect 126 8764 160 8798
rect 126 8696 160 8730
rect 126 8628 160 8662
rect 126 8560 160 8594
rect 126 8492 160 8526
rect 126 8424 160 8458
rect 126 8356 160 8390
rect 126 8288 160 8322
rect 126 8220 160 8254
rect 126 8152 160 8186
rect 126 8084 160 8118
rect 126 8016 160 8050
rect 126 7948 160 7982
rect 126 7880 160 7914
rect 126 7812 160 7846
rect 126 7744 160 7778
rect 126 7676 160 7710
rect 126 7608 160 7642
rect 126 7540 160 7574
rect 126 7472 160 7506
rect 126 7404 160 7438
rect 126 7336 160 7370
rect 126 7268 160 7302
rect 126 7200 160 7234
rect 126 7132 160 7166
rect 126 7064 160 7098
rect 126 6996 160 7030
rect 126 6928 160 6962
rect 126 6860 160 6894
rect 126 6792 160 6826
rect 126 6724 160 6758
rect 126 6656 160 6690
rect 126 6588 160 6622
rect 126 6520 160 6554
rect 126 6452 160 6486
rect 126 6384 160 6418
rect 126 6316 160 6350
rect 126 6248 160 6282
rect 126 6180 160 6214
rect 126 6112 160 6146
rect 126 6044 160 6078
rect 126 5976 160 6010
rect 126 5908 160 5942
rect 126 5840 160 5874
rect 126 5772 160 5806
rect 126 5704 160 5738
rect 126 5636 160 5670
rect 126 5568 160 5602
rect 126 5500 160 5534
rect 126 5432 160 5466
rect 126 5364 160 5398
rect 126 5296 160 5330
rect 126 5228 160 5262
rect 126 5160 160 5194
rect 126 5092 160 5126
rect 126 5024 160 5058
rect 126 4956 160 4990
rect 126 4888 160 4922
rect 126 4820 160 4854
rect 126 4752 160 4786
rect 126 4684 160 4718
rect 126 4616 160 4650
rect 126 4548 160 4582
rect 126 4480 160 4514
rect 126 4412 160 4446
rect 126 4344 160 4378
rect 126 4276 160 4310
rect 126 4208 160 4242
rect 126 4140 160 4174
rect 126 4072 160 4106
rect 126 4004 160 4038
rect 126 3936 160 3970
rect 126 3868 160 3902
rect 126 3800 160 3834
rect 126 3732 160 3766
rect 126 3664 160 3698
rect 126 3596 160 3630
rect 126 3528 160 3562
rect 126 3460 160 3494
rect 126 3392 160 3426
rect 126 3324 160 3358
rect 126 3256 160 3290
rect 126 3188 160 3222
rect 126 3120 160 3154
rect 126 3052 160 3086
rect 126 2984 160 3018
rect 126 2916 160 2950
rect 126 2848 160 2882
rect 126 2780 160 2814
rect 126 2712 160 2746
rect 126 2644 160 2678
rect 126 2576 160 2610
rect 126 2508 160 2542
rect 126 2440 160 2474
rect 126 2372 160 2406
rect 126 2304 160 2338
rect 126 2236 160 2270
rect 126 2168 160 2202
rect 126 2100 160 2134
rect 126 2032 160 2066
rect 126 1964 160 1998
rect 126 1896 160 1930
rect 126 1828 160 1862
rect 126 1760 160 1794
rect 126 1692 160 1726
rect 126 1624 160 1658
rect 126 1556 160 1590
rect 126 1488 160 1522
rect 126 1420 160 1454
rect 126 1352 160 1386
rect 126 1284 160 1318
rect 126 1216 160 1250
rect 126 1148 160 1182
rect 126 1080 160 1114
rect 126 1012 160 1046
rect 126 944 160 978
rect 126 876 160 910
rect 126 808 160 842
rect 126 740 160 774
rect 126 672 160 706
rect 126 604 160 638
rect 126 536 160 570
rect 3296 39158 3330 39192
rect 3296 39090 3330 39124
rect 3296 39022 3330 39056
rect 3296 38954 3330 38988
rect 3296 38886 3330 38920
rect 3296 38818 3330 38852
rect 3296 38750 3330 38784
rect 3296 38682 3330 38716
rect 3296 38614 3330 38648
rect 3296 38546 3330 38580
rect 3296 38478 3330 38512
rect 3296 38410 3330 38444
rect 3296 38342 3330 38376
rect 3296 38274 3330 38308
rect 3296 38206 3330 38240
rect 3296 38138 3330 38172
rect 3296 38070 3330 38104
rect 3296 38002 3330 38036
rect 3296 37934 3330 37968
rect 3296 37866 3330 37900
rect 3296 37798 3330 37832
rect 3296 37730 3330 37764
rect 3296 37662 3330 37696
rect 3296 37594 3330 37628
rect 3296 37526 3330 37560
rect 3296 37458 3330 37492
rect 3296 37390 3330 37424
rect 3296 37322 3330 37356
rect 3296 37254 3330 37288
rect 3296 37186 3330 37220
rect 3296 37118 3330 37152
rect 3296 37050 3330 37084
rect 3296 36982 3330 37016
rect 3296 36914 3330 36948
rect 3296 36846 3330 36880
rect 3296 36778 3330 36812
rect 3296 36710 3330 36744
rect 3296 36642 3330 36676
rect 3296 36574 3330 36608
rect 3296 36506 3330 36540
rect 3296 36438 3330 36472
rect 3296 36370 3330 36404
rect 3296 36302 3330 36336
rect 3296 36234 3330 36268
rect 3296 36166 3330 36200
rect 3296 36098 3330 36132
rect 3296 36030 3330 36064
rect 3296 35962 3330 35996
rect 3296 35894 3330 35928
rect 3296 35826 3330 35860
rect 3296 35758 3330 35792
rect 3296 35690 3330 35724
rect 3296 35622 3330 35656
rect 3296 35554 3330 35588
rect 3296 35486 3330 35520
rect 3296 35418 3330 35452
rect 3296 35350 3330 35384
rect 3296 35282 3330 35316
rect 3296 35214 3330 35248
rect 3296 35146 3330 35180
rect 3296 35078 3330 35112
rect 3296 35010 3330 35044
rect 3296 34942 3330 34976
rect 3296 34874 3330 34908
rect 3296 34806 3330 34840
rect 3296 34738 3330 34772
rect 3296 34670 3330 34704
rect 3296 34602 3330 34636
rect 3296 34534 3330 34568
rect 3296 34466 3330 34500
rect 3296 34398 3330 34432
rect 3296 34330 3330 34364
rect 3296 34262 3330 34296
rect 3296 34194 3330 34228
rect 3296 34126 3330 34160
rect 3296 34058 3330 34092
rect 3296 33990 3330 34024
rect 3296 33922 3330 33956
rect 3296 33854 3330 33888
rect 3296 33786 3330 33820
rect 3296 33718 3330 33752
rect 3296 33650 3330 33684
rect 3296 33582 3330 33616
rect 3296 33514 3330 33548
rect 3296 33446 3330 33480
rect 3296 33378 3330 33412
rect 3296 33310 3330 33344
rect 3296 33242 3330 33276
rect 3296 33174 3330 33208
rect 3296 33106 3330 33140
rect 3296 33038 3330 33072
rect 3296 32970 3330 33004
rect 3296 32902 3330 32936
rect 3296 32834 3330 32868
rect 3296 32766 3330 32800
rect 3296 32698 3330 32732
rect 3296 32630 3330 32664
rect 3296 32562 3330 32596
rect 3296 32494 3330 32528
rect 3296 32426 3330 32460
rect 3296 32358 3330 32392
rect 3296 32290 3330 32324
rect 3296 32222 3330 32256
rect 3296 32154 3330 32188
rect 3296 32086 3330 32120
rect 3296 32018 3330 32052
rect 3296 31950 3330 31984
rect 3296 31882 3330 31916
rect 3296 31814 3330 31848
rect 3296 31746 3330 31780
rect 3296 31678 3330 31712
rect 3296 31610 3330 31644
rect 3296 31542 3330 31576
rect 3296 31474 3330 31508
rect 3296 31406 3330 31440
rect 3296 31338 3330 31372
rect 3296 31270 3330 31304
rect 3296 31202 3330 31236
rect 3296 31134 3330 31168
rect 3296 31066 3330 31100
rect 3296 30998 3330 31032
rect 3296 30930 3330 30964
rect 3296 30862 3330 30896
rect 3296 30794 3330 30828
rect 3296 30726 3330 30760
rect 3296 30658 3330 30692
rect 3296 30590 3330 30624
rect 3296 30522 3330 30556
rect 3296 30454 3330 30488
rect 3296 30386 3330 30420
rect 3296 30318 3330 30352
rect 3296 30250 3330 30284
rect 3296 30182 3330 30216
rect 3296 30114 3330 30148
rect 3296 30046 3330 30080
rect 3296 29978 3330 30012
rect 3296 29910 3330 29944
rect 3296 29842 3330 29876
rect 3296 29774 3330 29808
rect 3296 29706 3330 29740
rect 3296 29638 3330 29672
rect 3296 29570 3330 29604
rect 3296 29502 3330 29536
rect 3296 29434 3330 29468
rect 3296 29366 3330 29400
rect 3296 29298 3330 29332
rect 3296 29230 3330 29264
rect 3296 29162 3330 29196
rect 3296 29094 3330 29128
rect 3296 29026 3330 29060
rect 3296 28958 3330 28992
rect 3296 28890 3330 28924
rect 3296 28822 3330 28856
rect 3296 28754 3330 28788
rect 3296 28686 3330 28720
rect 3296 28618 3330 28652
rect 3296 28550 3330 28584
rect 3296 28482 3330 28516
rect 3296 28414 3330 28448
rect 3296 28346 3330 28380
rect 3296 28278 3330 28312
rect 3296 28210 3330 28244
rect 3296 28142 3330 28176
rect 3296 28074 3330 28108
rect 3296 28006 3330 28040
rect 3296 27938 3330 27972
rect 3296 27870 3330 27904
rect 3296 27802 3330 27836
rect 3296 27734 3330 27768
rect 3296 27666 3330 27700
rect 3296 27598 3330 27632
rect 3296 27530 3330 27564
rect 3296 27462 3330 27496
rect 3296 27394 3330 27428
rect 3296 27326 3330 27360
rect 3296 27258 3330 27292
rect 3296 27190 3330 27224
rect 3296 27122 3330 27156
rect 3296 27054 3330 27088
rect 3296 26986 3330 27020
rect 3296 26918 3330 26952
rect 3296 26850 3330 26884
rect 3296 26782 3330 26816
rect 3296 26714 3330 26748
rect 3296 26646 3330 26680
rect 3296 26578 3330 26612
rect 3296 26510 3330 26544
rect 3296 26442 3330 26476
rect 3296 26374 3330 26408
rect 3296 26306 3330 26340
rect 3296 26238 3330 26272
rect 3296 26170 3330 26204
rect 3296 26102 3330 26136
rect 3296 26034 3330 26068
rect 3296 25966 3330 26000
rect 3296 25898 3330 25932
rect 3296 25830 3330 25864
rect 3296 25762 3330 25796
rect 3296 25694 3330 25728
rect 3296 25626 3330 25660
rect 3296 25558 3330 25592
rect 3296 25490 3330 25524
rect 3296 25422 3330 25456
rect 3296 25354 3330 25388
rect 3296 25286 3330 25320
rect 3296 25218 3330 25252
rect 3296 25150 3330 25184
rect 3296 25082 3330 25116
rect 3296 25014 3330 25048
rect 3296 24946 3330 24980
rect 3296 24878 3330 24912
rect 3296 24810 3330 24844
rect 3296 24742 3330 24776
rect 3296 24674 3330 24708
rect 3296 24606 3330 24640
rect 3296 24538 3330 24572
rect 3296 24470 3330 24504
rect 3296 24402 3330 24436
rect 3296 24334 3330 24368
rect 3296 24266 3330 24300
rect 3296 24198 3330 24232
rect 3296 24130 3330 24164
rect 3296 24062 3330 24096
rect 3296 23994 3330 24028
rect 3296 23926 3330 23960
rect 3296 23858 3330 23892
rect 3296 23790 3330 23824
rect 3296 23722 3330 23756
rect 3296 23654 3330 23688
rect 3296 23586 3330 23620
rect 3296 23518 3330 23552
rect 3296 23450 3330 23484
rect 3296 23382 3330 23416
rect 3296 23314 3330 23348
rect 3296 23246 3330 23280
rect 3296 23178 3330 23212
rect 3296 23110 3330 23144
rect 3296 23042 3330 23076
rect 3296 22974 3330 23008
rect 3296 22906 3330 22940
rect 3296 22838 3330 22872
rect 3296 22770 3330 22804
rect 3296 22702 3330 22736
rect 3296 22634 3330 22668
rect 3296 22566 3330 22600
rect 3296 22498 3330 22532
rect 3296 22430 3330 22464
rect 3296 22362 3330 22396
rect 3296 22294 3330 22328
rect 3296 22226 3330 22260
rect 3296 22158 3330 22192
rect 3296 22090 3330 22124
rect 3296 22022 3330 22056
rect 3296 21954 3330 21988
rect 3296 21886 3330 21920
rect 3296 21818 3330 21852
rect 3296 21750 3330 21784
rect 3296 21682 3330 21716
rect 3296 21614 3330 21648
rect 3296 21546 3330 21580
rect 3296 21478 3330 21512
rect 3296 21410 3330 21444
rect 3296 21342 3330 21376
rect 3296 21274 3330 21308
rect 3296 21206 3330 21240
rect 3296 21138 3330 21172
rect 3296 21070 3330 21104
rect 3296 21002 3330 21036
rect 3296 20934 3330 20968
rect 3296 20866 3330 20900
rect 3296 20798 3330 20832
rect 3296 20730 3330 20764
rect 3296 20662 3330 20696
rect 3296 20594 3330 20628
rect 3296 20526 3330 20560
rect 3296 20458 3330 20492
rect 3296 20390 3330 20424
rect 3296 20322 3330 20356
rect 3296 20254 3330 20288
rect 3296 20186 3330 20220
rect 3296 20118 3330 20152
rect 3296 20050 3330 20084
rect 3296 19982 3330 20016
rect 3296 19914 3330 19948
rect 3296 19846 3330 19880
rect 3296 19778 3330 19812
rect 3296 19710 3330 19744
rect 3296 19642 3330 19676
rect 3296 19574 3330 19608
rect 3296 19506 3330 19540
rect 3296 19438 3330 19472
rect 3296 19370 3330 19404
rect 3296 19302 3330 19336
rect 3296 19234 3330 19268
rect 3296 19166 3330 19200
rect 3296 19098 3330 19132
rect 3296 19030 3330 19064
rect 3296 18962 3330 18996
rect 3296 18894 3330 18928
rect 3296 18826 3330 18860
rect 3296 18758 3330 18792
rect 3296 18690 3330 18724
rect 3296 18622 3330 18656
rect 3296 18554 3330 18588
rect 3296 18486 3330 18520
rect 3296 18418 3330 18452
rect 3296 18350 3330 18384
rect 3296 18282 3330 18316
rect 3296 18214 3330 18248
rect 3296 18146 3330 18180
rect 3296 18078 3330 18112
rect 3296 18010 3330 18044
rect 3296 17942 3330 17976
rect 3296 17874 3330 17908
rect 3296 17806 3330 17840
rect 3296 17738 3330 17772
rect 3296 17670 3330 17704
rect 3296 17602 3330 17636
rect 3296 17534 3330 17568
rect 3296 17466 3330 17500
rect 3296 17398 3330 17432
rect 3296 17330 3330 17364
rect 3296 17262 3330 17296
rect 3296 17194 3330 17228
rect 3296 17126 3330 17160
rect 3296 17058 3330 17092
rect 3296 16990 3330 17024
rect 3296 16922 3330 16956
rect 3296 16854 3330 16888
rect 3296 16786 3330 16820
rect 3296 16718 3330 16752
rect 3296 16650 3330 16684
rect 3296 16582 3330 16616
rect 3296 16514 3330 16548
rect 3296 16446 3330 16480
rect 3296 16378 3330 16412
rect 3296 16310 3330 16344
rect 3296 16242 3330 16276
rect 3296 16174 3330 16208
rect 3296 16106 3330 16140
rect 3296 16038 3330 16072
rect 3296 15970 3330 16004
rect 3296 15902 3330 15936
rect 3296 15834 3330 15868
rect 3296 15766 3330 15800
rect 3296 15698 3330 15732
rect 3296 15630 3330 15664
rect 3296 15562 3330 15596
rect 3296 15494 3330 15528
rect 3296 15426 3330 15460
rect 3296 15358 3330 15392
rect 3296 15290 3330 15324
rect 3296 15222 3330 15256
rect 3296 15154 3330 15188
rect 3296 15086 3330 15120
rect 3296 15018 3330 15052
rect 3296 14950 3330 14984
rect 3296 14882 3330 14916
rect 3296 14814 3330 14848
rect 3296 14746 3330 14780
rect 3296 14678 3330 14712
rect 3296 14610 3330 14644
rect 3296 14542 3330 14576
rect 3296 14474 3330 14508
rect 3296 14406 3330 14440
rect 3296 14338 3330 14372
rect 3296 14270 3330 14304
rect 3296 14202 3330 14236
rect 3296 14134 3330 14168
rect 3296 14066 3330 14100
rect 3296 13998 3330 14032
rect 3296 13930 3330 13964
rect 3296 13862 3330 13896
rect 3296 13794 3330 13828
rect 3296 13726 3330 13760
rect 3296 13658 3330 13692
rect 3296 13590 3330 13624
rect 3296 13522 3330 13556
rect 3296 13454 3330 13488
rect 3296 13386 3330 13420
rect 3296 13318 3330 13352
rect 3296 13250 3330 13284
rect 3296 13182 3330 13216
rect 3296 13114 3330 13148
rect 3296 13046 3330 13080
rect 3296 12978 3330 13012
rect 3296 12910 3330 12944
rect 3296 12842 3330 12876
rect 3296 12774 3330 12808
rect 3296 12706 3330 12740
rect 3296 12638 3330 12672
rect 3296 12570 3330 12604
rect 3296 12502 3330 12536
rect 3296 12434 3330 12468
rect 3296 12366 3330 12400
rect 3296 12298 3330 12332
rect 3296 12230 3330 12264
rect 3296 12162 3330 12196
rect 3296 12094 3330 12128
rect 3296 12026 3330 12060
rect 3296 11958 3330 11992
rect 3296 11890 3330 11924
rect 3296 11822 3330 11856
rect 3296 11754 3330 11788
rect 3296 11686 3330 11720
rect 3296 11618 3330 11652
rect 3296 11550 3330 11584
rect 3296 11482 3330 11516
rect 3296 11414 3330 11448
rect 3296 11346 3330 11380
rect 3296 11278 3330 11312
rect 3296 11210 3330 11244
rect 3296 11142 3330 11176
rect 3296 11074 3330 11108
rect 3296 11006 3330 11040
rect 3296 10938 3330 10972
rect 3296 10870 3330 10904
rect 3296 10802 3330 10836
rect 3296 10734 3330 10768
rect 3296 10666 3330 10700
rect 3296 10598 3330 10632
rect 3296 10530 3330 10564
rect 3296 10462 3330 10496
rect 3296 10394 3330 10428
rect 3296 10326 3330 10360
rect 3296 10258 3330 10292
rect 3296 10190 3330 10224
rect 3296 10122 3330 10156
rect 3296 10054 3330 10088
rect 3296 9986 3330 10020
rect 3296 9918 3330 9952
rect 3296 9850 3330 9884
rect 3296 9782 3330 9816
rect 3296 9714 3330 9748
rect 3296 9646 3330 9680
rect 3296 9578 3330 9612
rect 3296 9510 3330 9544
rect 3296 9442 3330 9476
rect 3296 9374 3330 9408
rect 3296 9306 3330 9340
rect 3296 9238 3330 9272
rect 3296 9170 3330 9204
rect 3296 9102 3330 9136
rect 3296 9034 3330 9068
rect 3296 8966 3330 9000
rect 3296 8898 3330 8932
rect 3296 8830 3330 8864
rect 3296 8762 3330 8796
rect 3296 8694 3330 8728
rect 3296 8626 3330 8660
rect 3296 8558 3330 8592
rect 3296 8490 3330 8524
rect 3296 8422 3330 8456
rect 3296 8354 3330 8388
rect 3296 8286 3330 8320
rect 3296 8218 3330 8252
rect 3296 8150 3330 8184
rect 3296 8082 3330 8116
rect 3296 8014 3330 8048
rect 3296 7946 3330 7980
rect 3296 7878 3330 7912
rect 3296 7810 3330 7844
rect 3296 7742 3330 7776
rect 3296 7674 3330 7708
rect 3296 7606 3330 7640
rect 3296 7538 3330 7572
rect 3296 7470 3330 7504
rect 3296 7402 3330 7436
rect 3296 7334 3330 7368
rect 3296 7266 3330 7300
rect 3296 7198 3330 7232
rect 3296 7130 3330 7164
rect 3296 7062 3330 7096
rect 3296 6994 3330 7028
rect 3296 6926 3330 6960
rect 3296 6858 3330 6892
rect 3296 6790 3330 6824
rect 3296 6722 3330 6756
rect 3296 6654 3330 6688
rect 3296 6586 3330 6620
rect 3296 6518 3330 6552
rect 3296 6450 3330 6484
rect 3296 6382 3330 6416
rect 3296 6314 3330 6348
rect 3296 6246 3330 6280
rect 3296 6178 3330 6212
rect 3296 6110 3330 6144
rect 3296 6042 3330 6076
rect 3296 5974 3330 6008
rect 3296 5906 3330 5940
rect 3296 5838 3330 5872
rect 3296 5770 3330 5804
rect 3296 5702 3330 5736
rect 3296 5634 3330 5668
rect 3296 5566 3330 5600
rect 3296 5498 3330 5532
rect 3296 5430 3330 5464
rect 3296 5362 3330 5396
rect 3296 5294 3330 5328
rect 3296 5226 3330 5260
rect 3296 5158 3330 5192
rect 3296 5090 3330 5124
rect 3296 5022 3330 5056
rect 3296 4954 3330 4988
rect 3296 4886 3330 4920
rect 3296 4818 3330 4852
rect 3296 4750 3330 4784
rect 3296 4682 3330 4716
rect 3296 4614 3330 4648
rect 3296 4546 3330 4580
rect 3296 4478 3330 4512
rect 3296 4410 3330 4444
rect 3296 4342 3330 4376
rect 3296 4274 3330 4308
rect 3296 4206 3330 4240
rect 3296 4138 3330 4172
rect 3296 4070 3330 4104
rect 3296 4002 3330 4036
rect 3296 3934 3330 3968
rect 3296 3866 3330 3900
rect 3296 3798 3330 3832
rect 3296 3730 3330 3764
rect 3296 3662 3330 3696
rect 3296 3594 3330 3628
rect 3296 3526 3330 3560
rect 3296 3458 3330 3492
rect 3296 3390 3330 3424
rect 3296 3322 3330 3356
rect 3296 3254 3330 3288
rect 3296 3186 3330 3220
rect 3296 3118 3330 3152
rect 3296 3050 3330 3084
rect 3296 2982 3330 3016
rect 3296 2914 3330 2948
rect 3296 2846 3330 2880
rect 3296 2778 3330 2812
rect 3296 2710 3330 2744
rect 3296 2642 3330 2676
rect 3296 2574 3330 2608
rect 3296 2506 3330 2540
rect 3296 2438 3330 2472
rect 3296 2370 3330 2404
rect 3296 2302 3330 2336
rect 3296 2234 3330 2268
rect 3296 2166 3330 2200
rect 3296 2098 3330 2132
rect 3296 2030 3330 2064
rect 3296 1962 3330 1996
rect 3296 1894 3330 1928
rect 3296 1826 3330 1860
rect 3296 1758 3330 1792
rect 3296 1690 3330 1724
rect 3296 1622 3330 1656
rect 3296 1554 3330 1588
rect 3296 1486 3330 1520
rect 3296 1418 3330 1452
rect 3296 1350 3330 1384
rect 3296 1282 3330 1316
rect 3296 1214 3330 1248
rect 3296 1146 3330 1180
rect 3296 1078 3330 1112
rect 3296 1010 3330 1044
rect 3296 942 3330 976
rect 3296 874 3330 908
rect 3296 806 3330 840
rect 3296 738 3330 772
rect 3296 670 3330 704
rect 3296 602 3330 636
rect 3296 534 3330 568
rect 126 468 160 502
rect 126 400 160 434
rect 126 332 160 366
rect 126 218 160 252
rect 3296 466 3330 500
rect 3296 398 3330 432
rect 3296 330 3330 364
rect 3296 262 3330 296
rect 3296 194 3330 228
rect 194 126 228 160
rect 262 126 296 160
rect 330 126 364 160
rect 398 126 432 160
rect 466 126 500 160
rect 534 126 568 160
rect 602 126 636 160
rect 670 126 704 160
rect 738 126 772 160
rect 806 126 840 160
rect 874 126 908 160
rect 942 126 976 160
rect 1010 126 1044 160
rect 1078 126 1112 160
rect 1146 126 1180 160
rect 1214 126 1248 160
rect 1282 126 1316 160
rect 1350 126 1384 160
rect 1418 126 1452 160
rect 1486 126 1520 160
rect 1554 126 1588 160
rect 1622 126 1656 160
rect 1690 126 1724 160
rect 1758 126 1792 160
rect 1826 126 1860 160
rect 1894 126 1928 160
rect 1962 126 1996 160
rect 2030 126 2064 160
rect 2098 126 2132 160
rect 2166 126 2200 160
rect 2234 126 2268 160
rect 2302 126 2336 160
rect 2370 126 2404 160
rect 2438 126 2472 160
rect 2506 126 2540 160
rect 2574 126 2608 160
rect 2642 126 2676 160
rect 2710 126 2744 160
rect 2778 126 2812 160
rect 2846 126 2880 160
rect 2914 126 2948 160
rect 2982 126 3016 160
rect 3050 126 3084 160
rect 3118 126 3152 160
rect 3186 126 3220 160
<< poly >>
rect 576 39054 2880 39070
rect 576 39020 592 39054
rect 626 39020 662 39054
rect 696 39020 732 39054
rect 766 39020 802 39054
rect 836 39020 872 39054
rect 906 39020 942 39054
rect 976 39020 1012 39054
rect 1046 39020 1082 39054
rect 1116 39020 1152 39054
rect 1186 39020 1222 39054
rect 1256 39020 1292 39054
rect 1326 39020 1362 39054
rect 1396 39020 1432 39054
rect 1466 39020 1502 39054
rect 1536 39020 1572 39054
rect 1606 39020 1642 39054
rect 1676 39020 1712 39054
rect 1746 39020 1782 39054
rect 1816 39020 1852 39054
rect 1886 39020 1922 39054
rect 1956 39020 1992 39054
rect 2026 39020 2062 39054
rect 2096 39020 2132 39054
rect 2166 39020 2202 39054
rect 2236 39020 2272 39054
rect 2306 39020 2342 39054
rect 2376 39020 2412 39054
rect 2446 39020 2482 39054
rect 2516 39020 2552 39054
rect 2586 39020 2622 39054
rect 2656 39020 2692 39054
rect 2726 39020 2761 39054
rect 2795 39020 2830 39054
rect 2864 39020 2880 39054
rect 576 39004 2880 39020
rect 576 36924 2880 36940
rect 576 36890 592 36924
rect 626 36890 662 36924
rect 696 36890 732 36924
rect 766 36890 802 36924
rect 836 36890 872 36924
rect 906 36890 942 36924
rect 976 36890 1012 36924
rect 1046 36890 1082 36924
rect 1116 36890 1152 36924
rect 1186 36890 1222 36924
rect 1256 36890 1292 36924
rect 1326 36890 1362 36924
rect 1396 36890 1432 36924
rect 1466 36890 1502 36924
rect 1536 36890 1572 36924
rect 1606 36890 1642 36924
rect 1676 36890 1712 36924
rect 1746 36890 1782 36924
rect 1816 36890 1852 36924
rect 1886 36890 1922 36924
rect 1956 36890 1992 36924
rect 2026 36890 2062 36924
rect 2096 36890 2132 36924
rect 2166 36890 2202 36924
rect 2236 36890 2272 36924
rect 2306 36890 2342 36924
rect 2376 36890 2412 36924
rect 2446 36890 2482 36924
rect 2516 36890 2552 36924
rect 2586 36890 2622 36924
rect 2656 36890 2692 36924
rect 2726 36890 2761 36924
rect 2795 36890 2830 36924
rect 2864 36890 2880 36924
rect 576 36874 2880 36890
rect 576 34794 2880 34810
rect 576 34760 592 34794
rect 626 34760 662 34794
rect 696 34760 732 34794
rect 766 34760 802 34794
rect 836 34760 872 34794
rect 906 34760 942 34794
rect 976 34760 1012 34794
rect 1046 34760 1082 34794
rect 1116 34760 1152 34794
rect 1186 34760 1222 34794
rect 1256 34760 1292 34794
rect 1326 34760 1362 34794
rect 1396 34760 1432 34794
rect 1466 34760 1502 34794
rect 1536 34760 1572 34794
rect 1606 34760 1642 34794
rect 1676 34760 1712 34794
rect 1746 34760 1782 34794
rect 1816 34760 1852 34794
rect 1886 34760 1922 34794
rect 1956 34760 1992 34794
rect 2026 34760 2062 34794
rect 2096 34760 2132 34794
rect 2166 34760 2202 34794
rect 2236 34760 2272 34794
rect 2306 34760 2342 34794
rect 2376 34760 2412 34794
rect 2446 34760 2482 34794
rect 2516 34760 2552 34794
rect 2586 34760 2622 34794
rect 2656 34760 2692 34794
rect 2726 34760 2761 34794
rect 2795 34760 2830 34794
rect 2864 34760 2880 34794
rect 576 34744 2880 34760
rect 576 32664 2880 32680
rect 576 32630 592 32664
rect 626 32630 662 32664
rect 696 32630 732 32664
rect 766 32630 802 32664
rect 836 32630 872 32664
rect 906 32630 942 32664
rect 976 32630 1012 32664
rect 1046 32630 1082 32664
rect 1116 32630 1152 32664
rect 1186 32630 1222 32664
rect 1256 32630 1292 32664
rect 1326 32630 1362 32664
rect 1396 32630 1432 32664
rect 1466 32630 1502 32664
rect 1536 32630 1572 32664
rect 1606 32630 1642 32664
rect 1676 32630 1712 32664
rect 1746 32630 1782 32664
rect 1816 32630 1852 32664
rect 1886 32630 1922 32664
rect 1956 32630 1992 32664
rect 2026 32630 2062 32664
rect 2096 32630 2132 32664
rect 2166 32630 2202 32664
rect 2236 32630 2272 32664
rect 2306 32630 2342 32664
rect 2376 32630 2412 32664
rect 2446 32630 2482 32664
rect 2516 32630 2552 32664
rect 2586 32630 2622 32664
rect 2656 32630 2692 32664
rect 2726 32630 2761 32664
rect 2795 32630 2830 32664
rect 2864 32630 2880 32664
rect 576 32614 2880 32630
rect 576 30534 2880 30550
rect 576 30500 592 30534
rect 626 30500 662 30534
rect 696 30500 732 30534
rect 766 30500 802 30534
rect 836 30500 872 30534
rect 906 30500 942 30534
rect 976 30500 1012 30534
rect 1046 30500 1082 30534
rect 1116 30500 1152 30534
rect 1186 30500 1222 30534
rect 1256 30500 1292 30534
rect 1326 30500 1362 30534
rect 1396 30500 1432 30534
rect 1466 30500 1502 30534
rect 1536 30500 1572 30534
rect 1606 30500 1642 30534
rect 1676 30500 1712 30534
rect 1746 30500 1782 30534
rect 1816 30500 1852 30534
rect 1886 30500 1922 30534
rect 1956 30500 1992 30534
rect 2026 30500 2062 30534
rect 2096 30500 2132 30534
rect 2166 30500 2202 30534
rect 2236 30500 2272 30534
rect 2306 30500 2342 30534
rect 2376 30500 2412 30534
rect 2446 30500 2482 30534
rect 2516 30500 2552 30534
rect 2586 30500 2622 30534
rect 2656 30500 2692 30534
rect 2726 30500 2761 30534
rect 2795 30500 2830 30534
rect 2864 30500 2880 30534
rect 576 30484 2880 30500
rect 576 28404 2880 28420
rect 576 28370 592 28404
rect 626 28370 662 28404
rect 696 28370 732 28404
rect 766 28370 802 28404
rect 836 28370 872 28404
rect 906 28370 942 28404
rect 976 28370 1012 28404
rect 1046 28370 1082 28404
rect 1116 28370 1152 28404
rect 1186 28370 1222 28404
rect 1256 28370 1292 28404
rect 1326 28370 1362 28404
rect 1396 28370 1432 28404
rect 1466 28370 1502 28404
rect 1536 28370 1572 28404
rect 1606 28370 1642 28404
rect 1676 28370 1712 28404
rect 1746 28370 1782 28404
rect 1816 28370 1852 28404
rect 1886 28370 1922 28404
rect 1956 28370 1992 28404
rect 2026 28370 2062 28404
rect 2096 28370 2132 28404
rect 2166 28370 2202 28404
rect 2236 28370 2272 28404
rect 2306 28370 2342 28404
rect 2376 28370 2412 28404
rect 2446 28370 2482 28404
rect 2516 28370 2552 28404
rect 2586 28370 2622 28404
rect 2656 28370 2692 28404
rect 2726 28370 2761 28404
rect 2795 28370 2830 28404
rect 2864 28370 2880 28404
rect 576 28354 2880 28370
rect 576 26274 2880 26290
rect 576 26240 592 26274
rect 626 26240 662 26274
rect 696 26240 732 26274
rect 766 26240 802 26274
rect 836 26240 872 26274
rect 906 26240 942 26274
rect 976 26240 1012 26274
rect 1046 26240 1082 26274
rect 1116 26240 1152 26274
rect 1186 26240 1222 26274
rect 1256 26240 1292 26274
rect 1326 26240 1362 26274
rect 1396 26240 1432 26274
rect 1466 26240 1502 26274
rect 1536 26240 1572 26274
rect 1606 26240 1642 26274
rect 1676 26240 1712 26274
rect 1746 26240 1782 26274
rect 1816 26240 1852 26274
rect 1886 26240 1922 26274
rect 1956 26240 1992 26274
rect 2026 26240 2062 26274
rect 2096 26240 2132 26274
rect 2166 26240 2202 26274
rect 2236 26240 2272 26274
rect 2306 26240 2342 26274
rect 2376 26240 2412 26274
rect 2446 26240 2482 26274
rect 2516 26240 2552 26274
rect 2586 26240 2622 26274
rect 2656 26240 2692 26274
rect 2726 26240 2761 26274
rect 2795 26240 2830 26274
rect 2864 26240 2880 26274
rect 576 26224 2880 26240
rect 576 24144 2880 24160
rect 576 24110 592 24144
rect 626 24110 662 24144
rect 696 24110 732 24144
rect 766 24110 802 24144
rect 836 24110 872 24144
rect 906 24110 942 24144
rect 976 24110 1012 24144
rect 1046 24110 1082 24144
rect 1116 24110 1152 24144
rect 1186 24110 1222 24144
rect 1256 24110 1292 24144
rect 1326 24110 1362 24144
rect 1396 24110 1432 24144
rect 1466 24110 1502 24144
rect 1536 24110 1572 24144
rect 1606 24110 1642 24144
rect 1676 24110 1712 24144
rect 1746 24110 1782 24144
rect 1816 24110 1852 24144
rect 1886 24110 1922 24144
rect 1956 24110 1992 24144
rect 2026 24110 2062 24144
rect 2096 24110 2132 24144
rect 2166 24110 2202 24144
rect 2236 24110 2272 24144
rect 2306 24110 2342 24144
rect 2376 24110 2412 24144
rect 2446 24110 2482 24144
rect 2516 24110 2552 24144
rect 2586 24110 2622 24144
rect 2656 24110 2692 24144
rect 2726 24110 2761 24144
rect 2795 24110 2830 24144
rect 2864 24110 2880 24144
rect 576 24094 2880 24110
rect 576 22014 2880 22030
rect 576 21980 592 22014
rect 626 21980 662 22014
rect 696 21980 732 22014
rect 766 21980 802 22014
rect 836 21980 872 22014
rect 906 21980 942 22014
rect 976 21980 1012 22014
rect 1046 21980 1082 22014
rect 1116 21980 1152 22014
rect 1186 21980 1222 22014
rect 1256 21980 1292 22014
rect 1326 21980 1362 22014
rect 1396 21980 1432 22014
rect 1466 21980 1502 22014
rect 1536 21980 1572 22014
rect 1606 21980 1642 22014
rect 1676 21980 1712 22014
rect 1746 21980 1782 22014
rect 1816 21980 1852 22014
rect 1886 21980 1922 22014
rect 1956 21980 1992 22014
rect 2026 21980 2062 22014
rect 2096 21980 2132 22014
rect 2166 21980 2202 22014
rect 2236 21980 2272 22014
rect 2306 21980 2342 22014
rect 2376 21980 2412 22014
rect 2446 21980 2482 22014
rect 2516 21980 2552 22014
rect 2586 21980 2622 22014
rect 2656 21980 2692 22014
rect 2726 21980 2761 22014
rect 2795 21980 2830 22014
rect 2864 21980 2880 22014
rect 576 21964 2880 21980
rect 576 19884 2880 19900
rect 576 19850 592 19884
rect 626 19850 662 19884
rect 696 19850 732 19884
rect 766 19850 802 19884
rect 836 19850 872 19884
rect 906 19850 942 19884
rect 976 19850 1012 19884
rect 1046 19850 1082 19884
rect 1116 19850 1152 19884
rect 1186 19850 1222 19884
rect 1256 19850 1292 19884
rect 1326 19850 1362 19884
rect 1396 19850 1432 19884
rect 1466 19850 1502 19884
rect 1536 19850 1572 19884
rect 1606 19850 1642 19884
rect 1676 19850 1712 19884
rect 1746 19850 1782 19884
rect 1816 19850 1852 19884
rect 1886 19850 1922 19884
rect 1956 19850 1992 19884
rect 2026 19850 2062 19884
rect 2096 19850 2132 19884
rect 2166 19850 2202 19884
rect 2236 19850 2272 19884
rect 2306 19850 2342 19884
rect 2376 19850 2412 19884
rect 2446 19850 2482 19884
rect 2516 19850 2552 19884
rect 2586 19850 2622 19884
rect 2656 19850 2692 19884
rect 2726 19850 2761 19884
rect 2795 19850 2830 19884
rect 2864 19850 2880 19884
rect 576 19834 2880 19850
rect 576 17754 2880 17770
rect 576 17720 592 17754
rect 626 17720 662 17754
rect 696 17720 732 17754
rect 766 17720 802 17754
rect 836 17720 872 17754
rect 906 17720 942 17754
rect 976 17720 1012 17754
rect 1046 17720 1082 17754
rect 1116 17720 1152 17754
rect 1186 17720 1222 17754
rect 1256 17720 1292 17754
rect 1326 17720 1362 17754
rect 1396 17720 1432 17754
rect 1466 17720 1502 17754
rect 1536 17720 1572 17754
rect 1606 17720 1642 17754
rect 1676 17720 1712 17754
rect 1746 17720 1782 17754
rect 1816 17720 1852 17754
rect 1886 17720 1922 17754
rect 1956 17720 1992 17754
rect 2026 17720 2062 17754
rect 2096 17720 2132 17754
rect 2166 17720 2202 17754
rect 2236 17720 2272 17754
rect 2306 17720 2342 17754
rect 2376 17720 2412 17754
rect 2446 17720 2482 17754
rect 2516 17720 2552 17754
rect 2586 17720 2622 17754
rect 2656 17720 2692 17754
rect 2726 17720 2761 17754
rect 2795 17720 2830 17754
rect 2864 17720 2880 17754
rect 576 17704 2880 17720
rect 576 15624 2880 15640
rect 576 15590 592 15624
rect 626 15590 662 15624
rect 696 15590 732 15624
rect 766 15590 802 15624
rect 836 15590 872 15624
rect 906 15590 942 15624
rect 976 15590 1012 15624
rect 1046 15590 1082 15624
rect 1116 15590 1152 15624
rect 1186 15590 1222 15624
rect 1256 15590 1292 15624
rect 1326 15590 1362 15624
rect 1396 15590 1432 15624
rect 1466 15590 1502 15624
rect 1536 15590 1572 15624
rect 1606 15590 1642 15624
rect 1676 15590 1712 15624
rect 1746 15590 1782 15624
rect 1816 15590 1852 15624
rect 1886 15590 1922 15624
rect 1956 15590 1992 15624
rect 2026 15590 2062 15624
rect 2096 15590 2132 15624
rect 2166 15590 2202 15624
rect 2236 15590 2272 15624
rect 2306 15590 2342 15624
rect 2376 15590 2412 15624
rect 2446 15590 2482 15624
rect 2516 15590 2552 15624
rect 2586 15590 2622 15624
rect 2656 15590 2692 15624
rect 2726 15590 2761 15624
rect 2795 15590 2830 15624
rect 2864 15590 2880 15624
rect 576 15574 2880 15590
rect 576 13494 2880 13510
rect 576 13460 592 13494
rect 626 13460 662 13494
rect 696 13460 732 13494
rect 766 13460 802 13494
rect 836 13460 872 13494
rect 906 13460 942 13494
rect 976 13460 1012 13494
rect 1046 13460 1082 13494
rect 1116 13460 1152 13494
rect 1186 13460 1222 13494
rect 1256 13460 1292 13494
rect 1326 13460 1362 13494
rect 1396 13460 1432 13494
rect 1466 13460 1502 13494
rect 1536 13460 1572 13494
rect 1606 13460 1642 13494
rect 1676 13460 1712 13494
rect 1746 13460 1782 13494
rect 1816 13460 1852 13494
rect 1886 13460 1922 13494
rect 1956 13460 1992 13494
rect 2026 13460 2062 13494
rect 2096 13460 2132 13494
rect 2166 13460 2202 13494
rect 2236 13460 2272 13494
rect 2306 13460 2342 13494
rect 2376 13460 2412 13494
rect 2446 13460 2482 13494
rect 2516 13460 2552 13494
rect 2586 13460 2622 13494
rect 2656 13460 2692 13494
rect 2726 13460 2761 13494
rect 2795 13460 2830 13494
rect 2864 13460 2880 13494
rect 576 13444 2880 13460
rect 576 11364 2880 11380
rect 576 11330 592 11364
rect 626 11330 662 11364
rect 696 11330 732 11364
rect 766 11330 802 11364
rect 836 11330 872 11364
rect 906 11330 942 11364
rect 976 11330 1012 11364
rect 1046 11330 1082 11364
rect 1116 11330 1152 11364
rect 1186 11330 1222 11364
rect 1256 11330 1292 11364
rect 1326 11330 1362 11364
rect 1396 11330 1432 11364
rect 1466 11330 1502 11364
rect 1536 11330 1572 11364
rect 1606 11330 1642 11364
rect 1676 11330 1712 11364
rect 1746 11330 1782 11364
rect 1816 11330 1852 11364
rect 1886 11330 1922 11364
rect 1956 11330 1992 11364
rect 2026 11330 2062 11364
rect 2096 11330 2132 11364
rect 2166 11330 2202 11364
rect 2236 11330 2272 11364
rect 2306 11330 2342 11364
rect 2376 11330 2412 11364
rect 2446 11330 2482 11364
rect 2516 11330 2552 11364
rect 2586 11330 2622 11364
rect 2656 11330 2692 11364
rect 2726 11330 2761 11364
rect 2795 11330 2830 11364
rect 2864 11330 2880 11364
rect 576 11314 2880 11330
rect 576 9234 2880 9250
rect 576 9200 592 9234
rect 626 9200 662 9234
rect 696 9200 732 9234
rect 766 9200 802 9234
rect 836 9200 872 9234
rect 906 9200 942 9234
rect 976 9200 1012 9234
rect 1046 9200 1082 9234
rect 1116 9200 1152 9234
rect 1186 9200 1222 9234
rect 1256 9200 1292 9234
rect 1326 9200 1362 9234
rect 1396 9200 1432 9234
rect 1466 9200 1502 9234
rect 1536 9200 1572 9234
rect 1606 9200 1642 9234
rect 1676 9200 1712 9234
rect 1746 9200 1782 9234
rect 1816 9200 1852 9234
rect 1886 9200 1922 9234
rect 1956 9200 1992 9234
rect 2026 9200 2062 9234
rect 2096 9200 2132 9234
rect 2166 9200 2202 9234
rect 2236 9200 2272 9234
rect 2306 9200 2342 9234
rect 2376 9200 2412 9234
rect 2446 9200 2482 9234
rect 2516 9200 2552 9234
rect 2586 9200 2622 9234
rect 2656 9200 2692 9234
rect 2726 9200 2761 9234
rect 2795 9200 2830 9234
rect 2864 9200 2880 9234
rect 576 9184 2880 9200
rect 576 7104 2880 7120
rect 576 7070 592 7104
rect 626 7070 662 7104
rect 696 7070 732 7104
rect 766 7070 802 7104
rect 836 7070 872 7104
rect 906 7070 942 7104
rect 976 7070 1012 7104
rect 1046 7070 1082 7104
rect 1116 7070 1152 7104
rect 1186 7070 1222 7104
rect 1256 7070 1292 7104
rect 1326 7070 1362 7104
rect 1396 7070 1432 7104
rect 1466 7070 1502 7104
rect 1536 7070 1572 7104
rect 1606 7070 1642 7104
rect 1676 7070 1712 7104
rect 1746 7070 1782 7104
rect 1816 7070 1852 7104
rect 1886 7070 1922 7104
rect 1956 7070 1992 7104
rect 2026 7070 2062 7104
rect 2096 7070 2132 7104
rect 2166 7070 2202 7104
rect 2236 7070 2272 7104
rect 2306 7070 2342 7104
rect 2376 7070 2412 7104
rect 2446 7070 2482 7104
rect 2516 7070 2552 7104
rect 2586 7070 2622 7104
rect 2656 7070 2692 7104
rect 2726 7070 2761 7104
rect 2795 7070 2830 7104
rect 2864 7070 2880 7104
rect 576 7054 2880 7070
rect 576 4974 2880 4990
rect 576 4940 592 4974
rect 626 4940 662 4974
rect 696 4940 732 4974
rect 766 4940 802 4974
rect 836 4940 872 4974
rect 906 4940 942 4974
rect 976 4940 1012 4974
rect 1046 4940 1082 4974
rect 1116 4940 1152 4974
rect 1186 4940 1222 4974
rect 1256 4940 1292 4974
rect 1326 4940 1362 4974
rect 1396 4940 1432 4974
rect 1466 4940 1502 4974
rect 1536 4940 1572 4974
rect 1606 4940 1642 4974
rect 1676 4940 1712 4974
rect 1746 4940 1782 4974
rect 1816 4940 1852 4974
rect 1886 4940 1922 4974
rect 1956 4940 1992 4974
rect 2026 4940 2062 4974
rect 2096 4940 2132 4974
rect 2166 4940 2202 4974
rect 2236 4940 2272 4974
rect 2306 4940 2342 4974
rect 2376 4940 2412 4974
rect 2446 4940 2482 4974
rect 2516 4940 2552 4974
rect 2586 4940 2622 4974
rect 2656 4940 2692 4974
rect 2726 4940 2761 4974
rect 2795 4940 2830 4974
rect 2864 4940 2880 4974
rect 576 4924 2880 4940
rect 576 2844 2880 2860
rect 576 2810 592 2844
rect 626 2810 662 2844
rect 696 2810 732 2844
rect 766 2810 802 2844
rect 836 2810 872 2844
rect 906 2810 942 2844
rect 976 2810 1012 2844
rect 1046 2810 1082 2844
rect 1116 2810 1152 2844
rect 1186 2810 1222 2844
rect 1256 2810 1292 2844
rect 1326 2810 1362 2844
rect 1396 2810 1432 2844
rect 1466 2810 1502 2844
rect 1536 2810 1572 2844
rect 1606 2810 1642 2844
rect 1676 2810 1712 2844
rect 1746 2810 1782 2844
rect 1816 2810 1852 2844
rect 1886 2810 1922 2844
rect 1956 2810 1992 2844
rect 2026 2810 2062 2844
rect 2096 2810 2132 2844
rect 2166 2810 2202 2844
rect 2236 2810 2272 2844
rect 2306 2810 2342 2844
rect 2376 2810 2412 2844
rect 2446 2810 2482 2844
rect 2516 2810 2552 2844
rect 2586 2810 2622 2844
rect 2656 2810 2692 2844
rect 2726 2810 2761 2844
rect 2795 2810 2830 2844
rect 2864 2810 2880 2844
rect 576 2794 2880 2810
rect 576 714 2880 730
rect 576 680 592 714
rect 626 680 662 714
rect 696 680 732 714
rect 766 680 802 714
rect 836 680 872 714
rect 906 680 942 714
rect 976 680 1012 714
rect 1046 680 1082 714
rect 1116 680 1152 714
rect 1186 680 1222 714
rect 1256 680 1292 714
rect 1326 680 1362 714
rect 1396 680 1432 714
rect 1466 680 1502 714
rect 1536 680 1572 714
rect 1606 680 1642 714
rect 1676 680 1712 714
rect 1746 680 1782 714
rect 1816 680 1852 714
rect 1886 680 1922 714
rect 1956 680 1992 714
rect 2026 680 2062 714
rect 2096 680 2132 714
rect 2166 680 2202 714
rect 2236 680 2272 714
rect 2306 680 2342 714
rect 2376 680 2412 714
rect 2446 680 2482 714
rect 2516 680 2552 714
rect 2586 680 2622 714
rect 2656 680 2692 714
rect 2726 680 2761 714
rect 2795 680 2830 714
rect 2864 680 2880 714
rect 576 664 2880 680
<< polycont >>
rect 592 39020 626 39054
rect 662 39020 696 39054
rect 732 39020 766 39054
rect 802 39020 836 39054
rect 872 39020 906 39054
rect 942 39020 976 39054
rect 1012 39020 1046 39054
rect 1082 39020 1116 39054
rect 1152 39020 1186 39054
rect 1222 39020 1256 39054
rect 1292 39020 1326 39054
rect 1362 39020 1396 39054
rect 1432 39020 1466 39054
rect 1502 39020 1536 39054
rect 1572 39020 1606 39054
rect 1642 39020 1676 39054
rect 1712 39020 1746 39054
rect 1782 39020 1816 39054
rect 1852 39020 1886 39054
rect 1922 39020 1956 39054
rect 1992 39020 2026 39054
rect 2062 39020 2096 39054
rect 2132 39020 2166 39054
rect 2202 39020 2236 39054
rect 2272 39020 2306 39054
rect 2342 39020 2376 39054
rect 2412 39020 2446 39054
rect 2482 39020 2516 39054
rect 2552 39020 2586 39054
rect 2622 39020 2656 39054
rect 2692 39020 2726 39054
rect 2761 39020 2795 39054
rect 2830 39020 2864 39054
rect 592 36890 626 36924
rect 662 36890 696 36924
rect 732 36890 766 36924
rect 802 36890 836 36924
rect 872 36890 906 36924
rect 942 36890 976 36924
rect 1012 36890 1046 36924
rect 1082 36890 1116 36924
rect 1152 36890 1186 36924
rect 1222 36890 1256 36924
rect 1292 36890 1326 36924
rect 1362 36890 1396 36924
rect 1432 36890 1466 36924
rect 1502 36890 1536 36924
rect 1572 36890 1606 36924
rect 1642 36890 1676 36924
rect 1712 36890 1746 36924
rect 1782 36890 1816 36924
rect 1852 36890 1886 36924
rect 1922 36890 1956 36924
rect 1992 36890 2026 36924
rect 2062 36890 2096 36924
rect 2132 36890 2166 36924
rect 2202 36890 2236 36924
rect 2272 36890 2306 36924
rect 2342 36890 2376 36924
rect 2412 36890 2446 36924
rect 2482 36890 2516 36924
rect 2552 36890 2586 36924
rect 2622 36890 2656 36924
rect 2692 36890 2726 36924
rect 2761 36890 2795 36924
rect 2830 36890 2864 36924
rect 592 34760 626 34794
rect 662 34760 696 34794
rect 732 34760 766 34794
rect 802 34760 836 34794
rect 872 34760 906 34794
rect 942 34760 976 34794
rect 1012 34760 1046 34794
rect 1082 34760 1116 34794
rect 1152 34760 1186 34794
rect 1222 34760 1256 34794
rect 1292 34760 1326 34794
rect 1362 34760 1396 34794
rect 1432 34760 1466 34794
rect 1502 34760 1536 34794
rect 1572 34760 1606 34794
rect 1642 34760 1676 34794
rect 1712 34760 1746 34794
rect 1782 34760 1816 34794
rect 1852 34760 1886 34794
rect 1922 34760 1956 34794
rect 1992 34760 2026 34794
rect 2062 34760 2096 34794
rect 2132 34760 2166 34794
rect 2202 34760 2236 34794
rect 2272 34760 2306 34794
rect 2342 34760 2376 34794
rect 2412 34760 2446 34794
rect 2482 34760 2516 34794
rect 2552 34760 2586 34794
rect 2622 34760 2656 34794
rect 2692 34760 2726 34794
rect 2761 34760 2795 34794
rect 2830 34760 2864 34794
rect 592 32630 626 32664
rect 662 32630 696 32664
rect 732 32630 766 32664
rect 802 32630 836 32664
rect 872 32630 906 32664
rect 942 32630 976 32664
rect 1012 32630 1046 32664
rect 1082 32630 1116 32664
rect 1152 32630 1186 32664
rect 1222 32630 1256 32664
rect 1292 32630 1326 32664
rect 1362 32630 1396 32664
rect 1432 32630 1466 32664
rect 1502 32630 1536 32664
rect 1572 32630 1606 32664
rect 1642 32630 1676 32664
rect 1712 32630 1746 32664
rect 1782 32630 1816 32664
rect 1852 32630 1886 32664
rect 1922 32630 1956 32664
rect 1992 32630 2026 32664
rect 2062 32630 2096 32664
rect 2132 32630 2166 32664
rect 2202 32630 2236 32664
rect 2272 32630 2306 32664
rect 2342 32630 2376 32664
rect 2412 32630 2446 32664
rect 2482 32630 2516 32664
rect 2552 32630 2586 32664
rect 2622 32630 2656 32664
rect 2692 32630 2726 32664
rect 2761 32630 2795 32664
rect 2830 32630 2864 32664
rect 592 30500 626 30534
rect 662 30500 696 30534
rect 732 30500 766 30534
rect 802 30500 836 30534
rect 872 30500 906 30534
rect 942 30500 976 30534
rect 1012 30500 1046 30534
rect 1082 30500 1116 30534
rect 1152 30500 1186 30534
rect 1222 30500 1256 30534
rect 1292 30500 1326 30534
rect 1362 30500 1396 30534
rect 1432 30500 1466 30534
rect 1502 30500 1536 30534
rect 1572 30500 1606 30534
rect 1642 30500 1676 30534
rect 1712 30500 1746 30534
rect 1782 30500 1816 30534
rect 1852 30500 1886 30534
rect 1922 30500 1956 30534
rect 1992 30500 2026 30534
rect 2062 30500 2096 30534
rect 2132 30500 2166 30534
rect 2202 30500 2236 30534
rect 2272 30500 2306 30534
rect 2342 30500 2376 30534
rect 2412 30500 2446 30534
rect 2482 30500 2516 30534
rect 2552 30500 2586 30534
rect 2622 30500 2656 30534
rect 2692 30500 2726 30534
rect 2761 30500 2795 30534
rect 2830 30500 2864 30534
rect 592 28370 626 28404
rect 662 28370 696 28404
rect 732 28370 766 28404
rect 802 28370 836 28404
rect 872 28370 906 28404
rect 942 28370 976 28404
rect 1012 28370 1046 28404
rect 1082 28370 1116 28404
rect 1152 28370 1186 28404
rect 1222 28370 1256 28404
rect 1292 28370 1326 28404
rect 1362 28370 1396 28404
rect 1432 28370 1466 28404
rect 1502 28370 1536 28404
rect 1572 28370 1606 28404
rect 1642 28370 1676 28404
rect 1712 28370 1746 28404
rect 1782 28370 1816 28404
rect 1852 28370 1886 28404
rect 1922 28370 1956 28404
rect 1992 28370 2026 28404
rect 2062 28370 2096 28404
rect 2132 28370 2166 28404
rect 2202 28370 2236 28404
rect 2272 28370 2306 28404
rect 2342 28370 2376 28404
rect 2412 28370 2446 28404
rect 2482 28370 2516 28404
rect 2552 28370 2586 28404
rect 2622 28370 2656 28404
rect 2692 28370 2726 28404
rect 2761 28370 2795 28404
rect 2830 28370 2864 28404
rect 592 26240 626 26274
rect 662 26240 696 26274
rect 732 26240 766 26274
rect 802 26240 836 26274
rect 872 26240 906 26274
rect 942 26240 976 26274
rect 1012 26240 1046 26274
rect 1082 26240 1116 26274
rect 1152 26240 1186 26274
rect 1222 26240 1256 26274
rect 1292 26240 1326 26274
rect 1362 26240 1396 26274
rect 1432 26240 1466 26274
rect 1502 26240 1536 26274
rect 1572 26240 1606 26274
rect 1642 26240 1676 26274
rect 1712 26240 1746 26274
rect 1782 26240 1816 26274
rect 1852 26240 1886 26274
rect 1922 26240 1956 26274
rect 1992 26240 2026 26274
rect 2062 26240 2096 26274
rect 2132 26240 2166 26274
rect 2202 26240 2236 26274
rect 2272 26240 2306 26274
rect 2342 26240 2376 26274
rect 2412 26240 2446 26274
rect 2482 26240 2516 26274
rect 2552 26240 2586 26274
rect 2622 26240 2656 26274
rect 2692 26240 2726 26274
rect 2761 26240 2795 26274
rect 2830 26240 2864 26274
rect 592 24110 626 24144
rect 662 24110 696 24144
rect 732 24110 766 24144
rect 802 24110 836 24144
rect 872 24110 906 24144
rect 942 24110 976 24144
rect 1012 24110 1046 24144
rect 1082 24110 1116 24144
rect 1152 24110 1186 24144
rect 1222 24110 1256 24144
rect 1292 24110 1326 24144
rect 1362 24110 1396 24144
rect 1432 24110 1466 24144
rect 1502 24110 1536 24144
rect 1572 24110 1606 24144
rect 1642 24110 1676 24144
rect 1712 24110 1746 24144
rect 1782 24110 1816 24144
rect 1852 24110 1886 24144
rect 1922 24110 1956 24144
rect 1992 24110 2026 24144
rect 2062 24110 2096 24144
rect 2132 24110 2166 24144
rect 2202 24110 2236 24144
rect 2272 24110 2306 24144
rect 2342 24110 2376 24144
rect 2412 24110 2446 24144
rect 2482 24110 2516 24144
rect 2552 24110 2586 24144
rect 2622 24110 2656 24144
rect 2692 24110 2726 24144
rect 2761 24110 2795 24144
rect 2830 24110 2864 24144
rect 592 21980 626 22014
rect 662 21980 696 22014
rect 732 21980 766 22014
rect 802 21980 836 22014
rect 872 21980 906 22014
rect 942 21980 976 22014
rect 1012 21980 1046 22014
rect 1082 21980 1116 22014
rect 1152 21980 1186 22014
rect 1222 21980 1256 22014
rect 1292 21980 1326 22014
rect 1362 21980 1396 22014
rect 1432 21980 1466 22014
rect 1502 21980 1536 22014
rect 1572 21980 1606 22014
rect 1642 21980 1676 22014
rect 1712 21980 1746 22014
rect 1782 21980 1816 22014
rect 1852 21980 1886 22014
rect 1922 21980 1956 22014
rect 1992 21980 2026 22014
rect 2062 21980 2096 22014
rect 2132 21980 2166 22014
rect 2202 21980 2236 22014
rect 2272 21980 2306 22014
rect 2342 21980 2376 22014
rect 2412 21980 2446 22014
rect 2482 21980 2516 22014
rect 2552 21980 2586 22014
rect 2622 21980 2656 22014
rect 2692 21980 2726 22014
rect 2761 21980 2795 22014
rect 2830 21980 2864 22014
rect 592 19850 626 19884
rect 662 19850 696 19884
rect 732 19850 766 19884
rect 802 19850 836 19884
rect 872 19850 906 19884
rect 942 19850 976 19884
rect 1012 19850 1046 19884
rect 1082 19850 1116 19884
rect 1152 19850 1186 19884
rect 1222 19850 1256 19884
rect 1292 19850 1326 19884
rect 1362 19850 1396 19884
rect 1432 19850 1466 19884
rect 1502 19850 1536 19884
rect 1572 19850 1606 19884
rect 1642 19850 1676 19884
rect 1712 19850 1746 19884
rect 1782 19850 1816 19884
rect 1852 19850 1886 19884
rect 1922 19850 1956 19884
rect 1992 19850 2026 19884
rect 2062 19850 2096 19884
rect 2132 19850 2166 19884
rect 2202 19850 2236 19884
rect 2272 19850 2306 19884
rect 2342 19850 2376 19884
rect 2412 19850 2446 19884
rect 2482 19850 2516 19884
rect 2552 19850 2586 19884
rect 2622 19850 2656 19884
rect 2692 19850 2726 19884
rect 2761 19850 2795 19884
rect 2830 19850 2864 19884
rect 592 17720 626 17754
rect 662 17720 696 17754
rect 732 17720 766 17754
rect 802 17720 836 17754
rect 872 17720 906 17754
rect 942 17720 976 17754
rect 1012 17720 1046 17754
rect 1082 17720 1116 17754
rect 1152 17720 1186 17754
rect 1222 17720 1256 17754
rect 1292 17720 1326 17754
rect 1362 17720 1396 17754
rect 1432 17720 1466 17754
rect 1502 17720 1536 17754
rect 1572 17720 1606 17754
rect 1642 17720 1676 17754
rect 1712 17720 1746 17754
rect 1782 17720 1816 17754
rect 1852 17720 1886 17754
rect 1922 17720 1956 17754
rect 1992 17720 2026 17754
rect 2062 17720 2096 17754
rect 2132 17720 2166 17754
rect 2202 17720 2236 17754
rect 2272 17720 2306 17754
rect 2342 17720 2376 17754
rect 2412 17720 2446 17754
rect 2482 17720 2516 17754
rect 2552 17720 2586 17754
rect 2622 17720 2656 17754
rect 2692 17720 2726 17754
rect 2761 17720 2795 17754
rect 2830 17720 2864 17754
rect 592 15590 626 15624
rect 662 15590 696 15624
rect 732 15590 766 15624
rect 802 15590 836 15624
rect 872 15590 906 15624
rect 942 15590 976 15624
rect 1012 15590 1046 15624
rect 1082 15590 1116 15624
rect 1152 15590 1186 15624
rect 1222 15590 1256 15624
rect 1292 15590 1326 15624
rect 1362 15590 1396 15624
rect 1432 15590 1466 15624
rect 1502 15590 1536 15624
rect 1572 15590 1606 15624
rect 1642 15590 1676 15624
rect 1712 15590 1746 15624
rect 1782 15590 1816 15624
rect 1852 15590 1886 15624
rect 1922 15590 1956 15624
rect 1992 15590 2026 15624
rect 2062 15590 2096 15624
rect 2132 15590 2166 15624
rect 2202 15590 2236 15624
rect 2272 15590 2306 15624
rect 2342 15590 2376 15624
rect 2412 15590 2446 15624
rect 2482 15590 2516 15624
rect 2552 15590 2586 15624
rect 2622 15590 2656 15624
rect 2692 15590 2726 15624
rect 2761 15590 2795 15624
rect 2830 15590 2864 15624
rect 592 13460 626 13494
rect 662 13460 696 13494
rect 732 13460 766 13494
rect 802 13460 836 13494
rect 872 13460 906 13494
rect 942 13460 976 13494
rect 1012 13460 1046 13494
rect 1082 13460 1116 13494
rect 1152 13460 1186 13494
rect 1222 13460 1256 13494
rect 1292 13460 1326 13494
rect 1362 13460 1396 13494
rect 1432 13460 1466 13494
rect 1502 13460 1536 13494
rect 1572 13460 1606 13494
rect 1642 13460 1676 13494
rect 1712 13460 1746 13494
rect 1782 13460 1816 13494
rect 1852 13460 1886 13494
rect 1922 13460 1956 13494
rect 1992 13460 2026 13494
rect 2062 13460 2096 13494
rect 2132 13460 2166 13494
rect 2202 13460 2236 13494
rect 2272 13460 2306 13494
rect 2342 13460 2376 13494
rect 2412 13460 2446 13494
rect 2482 13460 2516 13494
rect 2552 13460 2586 13494
rect 2622 13460 2656 13494
rect 2692 13460 2726 13494
rect 2761 13460 2795 13494
rect 2830 13460 2864 13494
rect 592 11330 626 11364
rect 662 11330 696 11364
rect 732 11330 766 11364
rect 802 11330 836 11364
rect 872 11330 906 11364
rect 942 11330 976 11364
rect 1012 11330 1046 11364
rect 1082 11330 1116 11364
rect 1152 11330 1186 11364
rect 1222 11330 1256 11364
rect 1292 11330 1326 11364
rect 1362 11330 1396 11364
rect 1432 11330 1466 11364
rect 1502 11330 1536 11364
rect 1572 11330 1606 11364
rect 1642 11330 1676 11364
rect 1712 11330 1746 11364
rect 1782 11330 1816 11364
rect 1852 11330 1886 11364
rect 1922 11330 1956 11364
rect 1992 11330 2026 11364
rect 2062 11330 2096 11364
rect 2132 11330 2166 11364
rect 2202 11330 2236 11364
rect 2272 11330 2306 11364
rect 2342 11330 2376 11364
rect 2412 11330 2446 11364
rect 2482 11330 2516 11364
rect 2552 11330 2586 11364
rect 2622 11330 2656 11364
rect 2692 11330 2726 11364
rect 2761 11330 2795 11364
rect 2830 11330 2864 11364
rect 592 9200 626 9234
rect 662 9200 696 9234
rect 732 9200 766 9234
rect 802 9200 836 9234
rect 872 9200 906 9234
rect 942 9200 976 9234
rect 1012 9200 1046 9234
rect 1082 9200 1116 9234
rect 1152 9200 1186 9234
rect 1222 9200 1256 9234
rect 1292 9200 1326 9234
rect 1362 9200 1396 9234
rect 1432 9200 1466 9234
rect 1502 9200 1536 9234
rect 1572 9200 1606 9234
rect 1642 9200 1676 9234
rect 1712 9200 1746 9234
rect 1782 9200 1816 9234
rect 1852 9200 1886 9234
rect 1922 9200 1956 9234
rect 1992 9200 2026 9234
rect 2062 9200 2096 9234
rect 2132 9200 2166 9234
rect 2202 9200 2236 9234
rect 2272 9200 2306 9234
rect 2342 9200 2376 9234
rect 2412 9200 2446 9234
rect 2482 9200 2516 9234
rect 2552 9200 2586 9234
rect 2622 9200 2656 9234
rect 2692 9200 2726 9234
rect 2761 9200 2795 9234
rect 2830 9200 2864 9234
rect 592 7070 626 7104
rect 662 7070 696 7104
rect 732 7070 766 7104
rect 802 7070 836 7104
rect 872 7070 906 7104
rect 942 7070 976 7104
rect 1012 7070 1046 7104
rect 1082 7070 1116 7104
rect 1152 7070 1186 7104
rect 1222 7070 1256 7104
rect 1292 7070 1326 7104
rect 1362 7070 1396 7104
rect 1432 7070 1466 7104
rect 1502 7070 1536 7104
rect 1572 7070 1606 7104
rect 1642 7070 1676 7104
rect 1712 7070 1746 7104
rect 1782 7070 1816 7104
rect 1852 7070 1886 7104
rect 1922 7070 1956 7104
rect 1992 7070 2026 7104
rect 2062 7070 2096 7104
rect 2132 7070 2166 7104
rect 2202 7070 2236 7104
rect 2272 7070 2306 7104
rect 2342 7070 2376 7104
rect 2412 7070 2446 7104
rect 2482 7070 2516 7104
rect 2552 7070 2586 7104
rect 2622 7070 2656 7104
rect 2692 7070 2726 7104
rect 2761 7070 2795 7104
rect 2830 7070 2864 7104
rect 592 4940 626 4974
rect 662 4940 696 4974
rect 732 4940 766 4974
rect 802 4940 836 4974
rect 872 4940 906 4974
rect 942 4940 976 4974
rect 1012 4940 1046 4974
rect 1082 4940 1116 4974
rect 1152 4940 1186 4974
rect 1222 4940 1256 4974
rect 1292 4940 1326 4974
rect 1362 4940 1396 4974
rect 1432 4940 1466 4974
rect 1502 4940 1536 4974
rect 1572 4940 1606 4974
rect 1642 4940 1676 4974
rect 1712 4940 1746 4974
rect 1782 4940 1816 4974
rect 1852 4940 1886 4974
rect 1922 4940 1956 4974
rect 1992 4940 2026 4974
rect 2062 4940 2096 4974
rect 2132 4940 2166 4974
rect 2202 4940 2236 4974
rect 2272 4940 2306 4974
rect 2342 4940 2376 4974
rect 2412 4940 2446 4974
rect 2482 4940 2516 4974
rect 2552 4940 2586 4974
rect 2622 4940 2656 4974
rect 2692 4940 2726 4974
rect 2761 4940 2795 4974
rect 2830 4940 2864 4974
rect 592 2810 626 2844
rect 662 2810 696 2844
rect 732 2810 766 2844
rect 802 2810 836 2844
rect 872 2810 906 2844
rect 942 2810 976 2844
rect 1012 2810 1046 2844
rect 1082 2810 1116 2844
rect 1152 2810 1186 2844
rect 1222 2810 1256 2844
rect 1292 2810 1326 2844
rect 1362 2810 1396 2844
rect 1432 2810 1466 2844
rect 1502 2810 1536 2844
rect 1572 2810 1606 2844
rect 1642 2810 1676 2844
rect 1712 2810 1746 2844
rect 1782 2810 1816 2844
rect 1852 2810 1886 2844
rect 1922 2810 1956 2844
rect 1992 2810 2026 2844
rect 2062 2810 2096 2844
rect 2132 2810 2166 2844
rect 2202 2810 2236 2844
rect 2272 2810 2306 2844
rect 2342 2810 2376 2844
rect 2412 2810 2446 2844
rect 2482 2810 2516 2844
rect 2552 2810 2586 2844
rect 2622 2810 2656 2844
rect 2692 2810 2726 2844
rect 2761 2810 2795 2844
rect 2830 2810 2864 2844
rect 592 680 626 714
rect 662 680 696 714
rect 732 680 766 714
rect 802 680 836 714
rect 872 680 906 714
rect 942 680 976 714
rect 1012 680 1046 714
rect 1082 680 1116 714
rect 1152 680 1186 714
rect 1222 680 1256 714
rect 1292 680 1326 714
rect 1362 680 1396 714
rect 1432 680 1466 714
rect 1502 680 1536 714
rect 1572 680 1606 714
rect 1642 680 1676 714
rect 1712 680 1746 714
rect 1782 680 1816 714
rect 1852 680 1886 714
rect 1922 680 1956 714
rect 1992 680 2026 714
rect 2062 680 2096 714
rect 2132 680 2166 714
rect 2202 680 2236 714
rect 2272 680 2306 714
rect 2342 680 2376 714
rect 2412 680 2446 714
rect 2482 680 2516 714
rect 2552 680 2586 714
rect 2622 680 2656 714
rect 2692 680 2726 714
rect 2761 680 2795 714
rect 2830 680 2864 714
<< locali >>
rect 120 39874 3336 39880
rect 120 39840 206 39874
rect 270 39840 286 39874
rect 338 39840 366 39874
rect 406 39840 440 39874
rect 481 39840 508 39874
rect 562 39840 576 39874
rect 643 39840 644 39874
rect 678 39840 690 39874
rect 746 39840 780 39874
rect 834 39840 848 39874
rect 907 39840 916 39874
rect 980 39840 984 39874
rect 1018 39840 1019 39874
rect 1086 39840 1092 39874
rect 1154 39840 1165 39874
rect 1222 39840 1238 39874
rect 1290 39840 1311 39874
rect 1358 39840 1384 39874
rect 1426 39840 1457 39874
rect 1494 39840 1528 39874
rect 1564 39840 1596 39874
rect 1637 39840 1664 39874
rect 1710 39840 1732 39874
rect 1783 39840 1800 39874
rect 1856 39840 1868 39874
rect 1929 39840 1936 39874
rect 2002 39840 2004 39874
rect 2038 39840 2041 39874
rect 2106 39840 2114 39874
rect 2174 39840 2188 39874
rect 2242 39840 2262 39874
rect 2310 39840 2336 39874
rect 2378 39840 2410 39874
rect 2446 39840 2480 39874
rect 2518 39840 2548 39874
rect 2592 39840 2616 39874
rect 2666 39840 2684 39874
rect 2740 39840 2752 39874
rect 2814 39840 2820 39874
rect 2922 39840 2928 39874
rect 2990 39840 3002 39874
rect 3058 39840 3076 39874
rect 3126 39840 3150 39874
rect 3194 39840 3224 39874
rect 3262 39840 3336 39874
rect 120 39834 3336 39840
rect 120 39806 166 39834
rect 120 39768 126 39806
rect 160 39768 166 39806
rect 120 39738 166 39768
rect 120 39695 126 39738
rect 160 39695 166 39738
rect 120 39670 166 39695
rect 120 39622 126 39670
rect 160 39622 166 39670
rect 120 39602 166 39622
rect 120 39549 126 39602
rect 160 39549 166 39602
rect 120 39534 166 39549
rect 120 39476 126 39534
rect 160 39476 166 39534
rect 120 39466 166 39476
rect 120 39403 126 39466
rect 160 39403 166 39466
rect 120 39398 166 39403
rect 120 39296 126 39398
rect 160 39296 166 39398
rect 120 39291 166 39296
rect 120 39228 126 39291
rect 160 39228 166 39291
rect 120 39218 166 39228
rect 120 39160 126 39218
rect 160 39160 166 39218
rect 3290 39804 3336 39834
rect 3290 39768 3296 39804
rect 3330 39768 3336 39804
rect 3290 39736 3336 39768
rect 3290 39696 3296 39736
rect 3330 39696 3336 39736
rect 3290 39668 3336 39696
rect 3290 39624 3296 39668
rect 3330 39624 3336 39668
rect 3290 39600 3336 39624
rect 3290 39552 3296 39600
rect 3330 39552 3336 39600
rect 3290 39532 3336 39552
rect 3290 39480 3296 39532
rect 3330 39480 3336 39532
rect 3290 39464 3336 39480
rect 3290 39408 3296 39464
rect 3330 39408 3336 39464
rect 3290 39396 3336 39408
rect 3290 39336 3296 39396
rect 3330 39336 3336 39396
rect 3290 39328 3336 39336
rect 3290 39264 3296 39328
rect 3330 39264 3336 39328
rect 3290 39260 3336 39264
rect 120 39145 166 39160
rect 120 39092 126 39145
rect 160 39092 166 39145
rect 120 39072 166 39092
rect 120 39024 126 39072
rect 160 39024 166 39072
rect 120 38999 166 39024
rect 120 38956 126 38999
rect 160 38956 166 38999
rect 120 38926 166 38956
rect 120 38888 126 38926
rect 160 38888 166 38926
rect 120 38854 166 38888
rect 120 38819 126 38854
rect 160 38819 166 38854
rect 120 38786 166 38819
rect 120 38746 126 38786
rect 160 38746 166 38786
rect 120 38718 166 38746
rect 120 38673 126 38718
rect 160 38673 166 38718
rect 120 38650 166 38673
rect 120 38600 126 38650
rect 160 38600 166 38650
rect 120 38582 166 38600
rect 120 38527 126 38582
rect 160 38527 166 38582
rect 120 38514 166 38527
rect 120 38454 126 38514
rect 160 38454 166 38514
rect 120 38446 166 38454
rect 120 38381 126 38446
rect 160 38381 166 38446
rect 120 38378 166 38381
rect 120 38344 126 38378
rect 160 38344 166 38378
rect 120 38342 166 38344
rect 120 38276 126 38342
rect 160 38276 166 38342
rect 120 38269 166 38276
rect 120 38208 126 38269
rect 160 38208 166 38269
rect 120 38196 166 38208
rect 120 38140 126 38196
rect 160 38140 166 38196
rect 120 38123 166 38140
rect 120 38072 126 38123
rect 160 38072 166 38123
rect 120 38050 166 38072
rect 120 38004 126 38050
rect 160 38004 166 38050
rect 120 37977 166 38004
rect 120 37936 126 37977
rect 160 37936 166 37977
rect 120 37904 166 37936
rect 120 37868 126 37904
rect 160 37868 166 37904
rect 120 37834 166 37868
rect 120 37797 126 37834
rect 160 37797 166 37834
rect 120 37766 166 37797
rect 120 37724 126 37766
rect 160 37724 166 37766
rect 120 37698 166 37724
rect 120 37651 126 37698
rect 160 37651 166 37698
rect 120 37630 166 37651
rect 120 37578 126 37630
rect 160 37578 166 37630
rect 120 37562 166 37578
rect 120 37505 126 37562
rect 160 37505 166 37562
rect 120 37494 166 37505
rect 120 37432 126 37494
rect 160 37432 166 37494
rect 120 37426 166 37432
rect 120 37359 126 37426
rect 160 37359 166 37426
rect 120 37358 166 37359
rect 120 37324 126 37358
rect 160 37324 166 37358
rect 120 37320 166 37324
rect 120 37256 126 37320
rect 160 37256 166 37320
rect 120 37247 166 37256
rect 120 37188 126 37247
rect 160 37188 166 37247
rect 120 37174 166 37188
rect 120 37120 126 37174
rect 160 37120 166 37174
rect 120 37101 166 37120
rect 120 37052 126 37101
rect 160 37052 166 37101
rect 120 37028 166 37052
rect 120 36984 126 37028
rect 160 36984 166 37028
rect 120 36955 166 36984
rect 120 36916 126 36955
rect 160 36916 166 36955
rect 120 36882 166 36916
rect 120 36848 126 36882
rect 160 36848 166 36882
rect 120 36814 166 36848
rect 120 36775 126 36814
rect 160 36775 166 36814
rect 120 36746 166 36775
rect 120 36702 126 36746
rect 160 36702 166 36746
rect 120 36678 166 36702
rect 120 36630 126 36678
rect 160 36630 166 36678
rect 120 36610 166 36630
rect 120 36558 126 36610
rect 160 36558 166 36610
rect 120 36542 166 36558
rect 120 36486 126 36542
rect 160 36486 166 36542
rect 120 36474 166 36486
rect 120 36414 126 36474
rect 160 36414 166 36474
rect 120 36406 166 36414
rect 120 36342 126 36406
rect 160 36342 166 36406
rect 120 36338 166 36342
rect 120 36236 126 36338
rect 160 36236 166 36338
rect 120 36232 166 36236
rect 120 36168 126 36232
rect 160 36168 166 36232
rect 120 36160 166 36168
rect 120 36100 126 36160
rect 160 36100 166 36160
rect 120 36088 166 36100
rect 120 36032 126 36088
rect 160 36032 166 36088
rect 120 36016 166 36032
rect 120 35964 126 36016
rect 160 35964 166 36016
rect 120 35944 166 35964
rect 120 35896 126 35944
rect 160 35896 166 35944
rect 120 35872 166 35896
rect 120 35828 126 35872
rect 160 35828 166 35872
rect 120 35800 166 35828
rect 120 35760 126 35800
rect 160 35760 166 35800
rect 120 35728 166 35760
rect 120 35692 126 35728
rect 160 35692 166 35728
rect 120 35658 166 35692
rect 120 35622 126 35658
rect 160 35622 166 35658
rect 120 35590 166 35622
rect 120 35550 126 35590
rect 160 35550 166 35590
rect 120 35522 166 35550
rect 120 35478 126 35522
rect 160 35478 166 35522
rect 120 35454 166 35478
rect 120 35406 126 35454
rect 160 35406 166 35454
rect 120 35386 166 35406
rect 120 35334 126 35386
rect 160 35334 166 35386
rect 120 35318 166 35334
rect 120 35262 126 35318
rect 160 35262 166 35318
rect 120 35250 166 35262
rect 120 35190 126 35250
rect 160 35190 166 35250
rect 120 35182 166 35190
rect 120 35118 126 35182
rect 160 35118 166 35182
rect 120 35114 166 35118
rect 120 35012 126 35114
rect 160 35012 166 35114
rect 120 35008 166 35012
rect 120 34944 126 35008
rect 160 34944 166 35008
rect 120 34936 166 34944
rect 120 34876 126 34936
rect 160 34876 166 34936
rect 120 34864 166 34876
rect 120 34808 126 34864
rect 160 34808 166 34864
rect 120 34792 166 34808
rect 120 34740 126 34792
rect 160 34740 166 34792
rect 120 34720 166 34740
rect 120 34672 126 34720
rect 160 34672 166 34720
rect 120 34648 166 34672
rect 120 34604 126 34648
rect 160 34604 166 34648
rect 120 34576 166 34604
rect 120 34536 126 34576
rect 160 34536 166 34576
rect 120 34504 166 34536
rect 120 34468 126 34504
rect 160 34468 166 34504
rect 120 34434 166 34468
rect 120 34398 126 34434
rect 160 34398 166 34434
rect 120 34366 166 34398
rect 120 34326 126 34366
rect 160 34326 166 34366
rect 120 34298 166 34326
rect 120 34254 126 34298
rect 160 34254 166 34298
rect 120 34230 166 34254
rect 120 34182 126 34230
rect 160 34182 166 34230
rect 120 34162 166 34182
rect 120 34110 126 34162
rect 160 34110 166 34162
rect 120 34094 166 34110
rect 120 34038 126 34094
rect 160 34038 166 34094
rect 120 34026 166 34038
rect 120 33966 126 34026
rect 160 33966 166 34026
rect 120 33958 166 33966
rect 120 33894 126 33958
rect 160 33894 166 33958
rect 120 33890 166 33894
rect 120 33788 126 33890
rect 160 33788 166 33890
rect 120 33784 166 33788
rect 120 33720 126 33784
rect 160 33720 166 33784
rect 120 33712 166 33720
rect 120 33652 126 33712
rect 160 33652 166 33712
rect 120 33640 166 33652
rect 120 33584 126 33640
rect 160 33584 166 33640
rect 120 33568 166 33584
rect 120 33516 126 33568
rect 160 33516 166 33568
rect 120 33496 166 33516
rect 120 33448 126 33496
rect 160 33448 166 33496
rect 120 33424 166 33448
rect 120 33380 126 33424
rect 160 33380 166 33424
rect 120 33352 166 33380
rect 120 33312 126 33352
rect 160 33312 166 33352
rect 120 33280 166 33312
rect 120 33244 126 33280
rect 160 33244 166 33280
rect 120 33210 166 33244
rect 120 33174 126 33210
rect 160 33174 166 33210
rect 120 33142 166 33174
rect 120 33102 126 33142
rect 160 33102 166 33142
rect 120 33074 166 33102
rect 120 33030 126 33074
rect 160 33030 166 33074
rect 120 33006 166 33030
rect 120 32958 126 33006
rect 160 32958 166 33006
rect 120 32938 166 32958
rect 120 32886 126 32938
rect 160 32886 166 32938
rect 120 32870 166 32886
rect 120 32814 126 32870
rect 160 32814 166 32870
rect 120 32802 166 32814
rect 120 32742 126 32802
rect 160 32742 166 32802
rect 120 32734 166 32742
rect 120 32670 126 32734
rect 160 32670 166 32734
rect 120 32666 166 32670
rect 120 32564 126 32666
rect 160 32564 166 32666
rect 120 32560 166 32564
rect 120 32496 126 32560
rect 160 32496 166 32560
rect 120 32488 166 32496
rect 120 32428 126 32488
rect 160 32428 166 32488
rect 120 32416 166 32428
rect 120 32360 126 32416
rect 160 32360 166 32416
rect 120 32344 166 32360
rect 120 32292 126 32344
rect 160 32292 166 32344
rect 120 32272 166 32292
rect 120 32224 126 32272
rect 160 32224 166 32272
rect 120 32200 166 32224
rect 120 32156 126 32200
rect 160 32156 166 32200
rect 120 32128 166 32156
rect 120 32088 126 32128
rect 160 32088 166 32128
rect 120 32056 166 32088
rect 120 32020 126 32056
rect 160 32020 166 32056
rect 120 31986 166 32020
rect 120 31950 126 31986
rect 160 31950 166 31986
rect 120 31918 166 31950
rect 120 31878 126 31918
rect 160 31878 166 31918
rect 120 31850 166 31878
rect 120 31806 126 31850
rect 160 31806 166 31850
rect 120 31782 166 31806
rect 120 31734 126 31782
rect 160 31734 166 31782
rect 120 31714 166 31734
rect 120 31662 126 31714
rect 160 31662 166 31714
rect 120 31646 166 31662
rect 120 31590 126 31646
rect 160 31590 166 31646
rect 120 31578 166 31590
rect 120 31518 126 31578
rect 160 31518 166 31578
rect 120 31510 166 31518
rect 120 31446 126 31510
rect 160 31446 166 31510
rect 120 31442 166 31446
rect 120 31340 126 31442
rect 160 31340 166 31442
rect 120 31336 166 31340
rect 120 31272 126 31336
rect 160 31272 166 31336
rect 120 31264 166 31272
rect 120 31204 126 31264
rect 160 31204 166 31264
rect 120 31192 166 31204
rect 120 31136 126 31192
rect 160 31136 166 31192
rect 120 31120 166 31136
rect 120 31068 126 31120
rect 160 31068 166 31120
rect 120 31048 166 31068
rect 120 31000 126 31048
rect 160 31000 166 31048
rect 120 30976 166 31000
rect 120 30932 126 30976
rect 160 30932 166 30976
rect 120 30904 166 30932
rect 120 30864 126 30904
rect 160 30864 166 30904
rect 120 30832 166 30864
rect 120 30796 126 30832
rect 160 30796 166 30832
rect 120 30762 166 30796
rect 120 30726 126 30762
rect 160 30726 166 30762
rect 120 30694 166 30726
rect 120 30654 126 30694
rect 160 30654 166 30694
rect 120 30626 166 30654
rect 120 30582 126 30626
rect 160 30582 166 30626
rect 120 30558 166 30582
rect 120 30510 126 30558
rect 160 30510 166 30558
rect 120 30490 166 30510
rect 120 30438 126 30490
rect 160 30438 166 30490
rect 120 30422 166 30438
rect 120 30366 126 30422
rect 160 30366 166 30422
rect 120 30354 166 30366
rect 120 30294 126 30354
rect 160 30294 166 30354
rect 120 30286 166 30294
rect 120 30222 126 30286
rect 160 30222 166 30286
rect 120 30218 166 30222
rect 120 30116 126 30218
rect 160 30116 166 30218
rect 120 30112 166 30116
rect 120 30048 126 30112
rect 160 30048 166 30112
rect 120 30040 166 30048
rect 120 29980 126 30040
rect 160 29980 166 30040
rect 120 29968 166 29980
rect 120 29912 126 29968
rect 160 29912 166 29968
rect 120 29896 166 29912
rect 120 29844 126 29896
rect 160 29844 166 29896
rect 120 29824 166 29844
rect 120 29776 126 29824
rect 160 29776 166 29824
rect 120 29752 166 29776
rect 120 29708 126 29752
rect 160 29708 166 29752
rect 120 29680 166 29708
rect 120 29640 126 29680
rect 160 29640 166 29680
rect 120 29608 166 29640
rect 120 29572 126 29608
rect 160 29572 166 29608
rect 120 29538 166 29572
rect 120 29502 126 29538
rect 160 29502 166 29538
rect 120 29470 166 29502
rect 120 29430 126 29470
rect 160 29430 166 29470
rect 120 29402 166 29430
rect 120 29358 126 29402
rect 160 29358 166 29402
rect 120 29334 166 29358
rect 120 29286 126 29334
rect 160 29286 166 29334
rect 120 29266 166 29286
rect 120 29214 126 29266
rect 160 29214 166 29266
rect 120 29198 166 29214
rect 120 29142 126 29198
rect 160 29142 166 29198
rect 120 29130 166 29142
rect 120 29070 126 29130
rect 160 29070 166 29130
rect 120 29062 166 29070
rect 120 28998 126 29062
rect 160 28998 166 29062
rect 120 28994 166 28998
rect 120 28892 126 28994
rect 160 28892 166 28994
rect 120 28888 166 28892
rect 120 28824 126 28888
rect 160 28824 166 28888
rect 120 28816 166 28824
rect 120 28756 126 28816
rect 160 28756 166 28816
rect 120 28744 166 28756
rect 120 28688 126 28744
rect 160 28688 166 28744
rect 120 28672 166 28688
rect 120 28620 126 28672
rect 160 28620 166 28672
rect 120 28600 166 28620
rect 120 28552 126 28600
rect 160 28552 166 28600
rect 120 28528 166 28552
rect 120 28484 126 28528
rect 160 28484 166 28528
rect 120 28456 166 28484
rect 120 28416 126 28456
rect 160 28416 166 28456
rect 120 28384 166 28416
rect 120 28348 126 28384
rect 160 28348 166 28384
rect 120 28314 166 28348
rect 120 28278 126 28314
rect 160 28278 166 28314
rect 120 28246 166 28278
rect 120 28206 126 28246
rect 160 28206 166 28246
rect 120 28178 166 28206
rect 120 28134 126 28178
rect 160 28134 166 28178
rect 120 28110 166 28134
rect 120 28062 126 28110
rect 160 28062 166 28110
rect 120 28042 166 28062
rect 120 27990 126 28042
rect 160 27990 166 28042
rect 120 27974 166 27990
rect 120 27918 126 27974
rect 160 27918 166 27974
rect 120 27906 166 27918
rect 120 27846 126 27906
rect 160 27846 166 27906
rect 120 27838 166 27846
rect 120 27774 126 27838
rect 160 27774 166 27838
rect 120 27770 166 27774
rect 120 27668 126 27770
rect 160 27668 166 27770
rect 120 27664 166 27668
rect 120 27600 126 27664
rect 160 27600 166 27664
rect 120 27592 166 27600
rect 120 27532 126 27592
rect 160 27532 166 27592
rect 120 27520 166 27532
rect 120 27464 126 27520
rect 160 27464 166 27520
rect 120 27448 166 27464
rect 120 27396 126 27448
rect 160 27396 166 27448
rect 120 27376 166 27396
rect 120 27328 126 27376
rect 160 27328 166 27376
rect 120 27304 166 27328
rect 120 27260 126 27304
rect 160 27260 166 27304
rect 120 27232 166 27260
rect 120 27192 126 27232
rect 160 27192 166 27232
rect 120 27160 166 27192
rect 120 27124 126 27160
rect 160 27124 166 27160
rect 120 27090 166 27124
rect 120 27054 126 27090
rect 160 27054 166 27090
rect 120 27022 166 27054
rect 120 26982 126 27022
rect 160 26982 166 27022
rect 120 26954 166 26982
rect 120 26910 126 26954
rect 160 26910 166 26954
rect 120 26886 166 26910
rect 120 26838 126 26886
rect 160 26838 166 26886
rect 120 26818 166 26838
rect 120 26766 126 26818
rect 160 26766 166 26818
rect 120 26750 166 26766
rect 120 26694 126 26750
rect 160 26694 166 26750
rect 120 26682 166 26694
rect 120 26622 126 26682
rect 160 26622 166 26682
rect 120 26614 166 26622
rect 120 26550 126 26614
rect 160 26550 166 26614
rect 120 26546 166 26550
rect 120 26444 126 26546
rect 160 26444 166 26546
rect 120 26440 166 26444
rect 120 26376 126 26440
rect 160 26376 166 26440
rect 120 26368 166 26376
rect 120 26308 126 26368
rect 160 26308 166 26368
rect 120 26296 166 26308
rect 120 26240 126 26296
rect 160 26240 166 26296
rect 120 26224 166 26240
rect 120 26172 126 26224
rect 160 26172 166 26224
rect 120 26152 166 26172
rect 120 26104 126 26152
rect 160 26104 166 26152
rect 120 26080 166 26104
rect 120 26036 126 26080
rect 160 26036 166 26080
rect 120 26008 166 26036
rect 120 25968 126 26008
rect 160 25968 166 26008
rect 120 25936 166 25968
rect 120 25900 126 25936
rect 160 25900 166 25936
rect 120 25866 166 25900
rect 120 25830 126 25866
rect 160 25830 166 25866
rect 120 25798 166 25830
rect 120 25758 126 25798
rect 160 25758 166 25798
rect 120 25730 166 25758
rect 120 25686 126 25730
rect 160 25686 166 25730
rect 120 25662 166 25686
rect 120 25614 126 25662
rect 160 25614 166 25662
rect 120 25594 166 25614
rect 120 25542 126 25594
rect 160 25542 166 25594
rect 120 25526 166 25542
rect 120 25470 126 25526
rect 160 25470 166 25526
rect 120 25458 166 25470
rect 120 25398 126 25458
rect 160 25398 166 25458
rect 120 25390 166 25398
rect 120 25326 126 25390
rect 160 25326 166 25390
rect 120 25322 166 25326
rect 120 25220 126 25322
rect 160 25220 166 25322
rect 120 25216 166 25220
rect 120 25152 126 25216
rect 160 25152 166 25216
rect 120 25144 166 25152
rect 120 25084 126 25144
rect 160 25084 166 25144
rect 120 25072 166 25084
rect 120 25016 126 25072
rect 160 25016 166 25072
rect 120 25000 166 25016
rect 120 24948 126 25000
rect 160 24948 166 25000
rect 120 24928 166 24948
rect 120 24880 126 24928
rect 160 24880 166 24928
rect 120 24856 166 24880
rect 120 24812 126 24856
rect 160 24812 166 24856
rect 120 24784 166 24812
rect 120 24744 126 24784
rect 160 24744 166 24784
rect 120 24712 166 24744
rect 120 24676 126 24712
rect 160 24676 166 24712
rect 120 24642 166 24676
rect 120 24606 126 24642
rect 160 24606 166 24642
rect 120 24574 166 24606
rect 120 24534 126 24574
rect 160 24534 166 24574
rect 120 24506 166 24534
rect 120 24462 126 24506
rect 160 24462 166 24506
rect 120 24438 166 24462
rect 120 24390 126 24438
rect 160 24390 166 24438
rect 120 24370 166 24390
rect 120 24318 126 24370
rect 160 24318 166 24370
rect 120 24302 166 24318
rect 120 24246 126 24302
rect 160 24246 166 24302
rect 120 24234 166 24246
rect 120 24174 126 24234
rect 160 24174 166 24234
rect 120 24166 166 24174
rect 120 24102 126 24166
rect 160 24102 166 24166
rect 120 24098 166 24102
rect 120 23996 126 24098
rect 160 23996 166 24098
rect 120 23992 166 23996
rect 120 23928 126 23992
rect 160 23928 166 23992
rect 120 23920 166 23928
rect 120 23860 126 23920
rect 160 23860 166 23920
rect 120 23848 166 23860
rect 120 23792 126 23848
rect 160 23792 166 23848
rect 120 23776 166 23792
rect 120 23724 126 23776
rect 160 23724 166 23776
rect 120 23704 166 23724
rect 120 23656 126 23704
rect 160 23656 166 23704
rect 120 23632 166 23656
rect 120 23588 126 23632
rect 160 23588 166 23632
rect 120 23560 166 23588
rect 120 23520 126 23560
rect 160 23520 166 23560
rect 120 23488 166 23520
rect 120 23452 126 23488
rect 160 23452 166 23488
rect 120 23418 166 23452
rect 120 23382 126 23418
rect 160 23382 166 23418
rect 120 23350 166 23382
rect 120 23310 126 23350
rect 160 23310 166 23350
rect 120 23282 166 23310
rect 120 23238 126 23282
rect 160 23238 166 23282
rect 120 23214 166 23238
rect 120 23166 126 23214
rect 160 23166 166 23214
rect 120 23146 166 23166
rect 120 23094 126 23146
rect 160 23094 166 23146
rect 120 23078 166 23094
rect 120 23022 126 23078
rect 160 23022 166 23078
rect 120 23010 166 23022
rect 120 22950 126 23010
rect 160 22950 166 23010
rect 120 22942 166 22950
rect 120 22878 126 22942
rect 160 22878 166 22942
rect 120 22874 166 22878
rect 120 22772 126 22874
rect 160 22772 166 22874
rect 120 22768 166 22772
rect 120 22704 126 22768
rect 160 22704 166 22768
rect 120 22696 166 22704
rect 120 22636 126 22696
rect 160 22636 166 22696
rect 120 22624 166 22636
rect 120 22568 126 22624
rect 160 22568 166 22624
rect 120 22552 166 22568
rect 120 22500 126 22552
rect 160 22500 166 22552
rect 120 22480 166 22500
rect 120 22432 126 22480
rect 160 22432 166 22480
rect 120 22408 166 22432
rect 120 22364 126 22408
rect 160 22364 166 22408
rect 120 22336 166 22364
rect 120 22296 126 22336
rect 160 22296 166 22336
rect 120 22264 166 22296
rect 120 22228 126 22264
rect 160 22228 166 22264
rect 120 22194 166 22228
rect 120 22158 126 22194
rect 160 22158 166 22194
rect 120 22126 166 22158
rect 120 22086 126 22126
rect 160 22086 166 22126
rect 120 22058 166 22086
rect 120 22014 126 22058
rect 160 22014 166 22058
rect 120 21990 166 22014
rect 120 21942 126 21990
rect 160 21942 166 21990
rect 120 21922 166 21942
rect 120 21870 126 21922
rect 160 21870 166 21922
rect 120 21854 166 21870
rect 120 21798 126 21854
rect 160 21798 166 21854
rect 120 21786 166 21798
rect 120 21726 126 21786
rect 160 21726 166 21786
rect 120 21718 166 21726
rect 120 21654 126 21718
rect 160 21654 166 21718
rect 120 21650 166 21654
rect 120 21548 126 21650
rect 160 21548 166 21650
rect 120 21544 166 21548
rect 120 21480 126 21544
rect 160 21480 166 21544
rect 120 21472 166 21480
rect 120 21412 126 21472
rect 160 21412 166 21472
rect 120 21400 166 21412
rect 120 21344 126 21400
rect 160 21344 166 21400
rect 120 21328 166 21344
rect 120 21276 126 21328
rect 160 21276 166 21328
rect 120 21256 166 21276
rect 120 21208 126 21256
rect 160 21208 166 21256
rect 120 21184 166 21208
rect 120 21140 126 21184
rect 160 21140 166 21184
rect 120 21112 166 21140
rect 120 21072 126 21112
rect 160 21072 166 21112
rect 120 21040 166 21072
rect 120 21004 126 21040
rect 160 21004 166 21040
rect 120 20970 166 21004
rect 120 20934 126 20970
rect 160 20934 166 20970
rect 120 20902 166 20934
rect 120 20862 126 20902
rect 160 20862 166 20902
rect 120 20834 166 20862
rect 120 20790 126 20834
rect 160 20790 166 20834
rect 120 20766 166 20790
rect 120 20718 126 20766
rect 160 20718 166 20766
rect 120 20698 166 20718
rect 120 20646 126 20698
rect 160 20646 166 20698
rect 120 20630 166 20646
rect 120 20574 126 20630
rect 160 20574 166 20630
rect 120 20562 166 20574
rect 120 20502 126 20562
rect 160 20502 166 20562
rect 120 20494 166 20502
rect 120 20430 126 20494
rect 160 20430 166 20494
rect 120 20426 166 20430
rect 120 20324 126 20426
rect 160 20324 166 20426
rect 120 20320 166 20324
rect 120 20256 126 20320
rect 160 20256 166 20320
rect 120 20248 166 20256
rect 120 20188 126 20248
rect 160 20188 166 20248
rect 120 20176 166 20188
rect 120 20120 126 20176
rect 160 20120 166 20176
rect 120 20104 166 20120
rect 120 20052 126 20104
rect 160 20052 166 20104
rect 120 20032 166 20052
rect 120 19984 126 20032
rect 160 19984 166 20032
rect 120 19960 166 19984
rect 120 19916 126 19960
rect 160 19916 166 19960
rect 120 19888 166 19916
rect 120 19848 126 19888
rect 160 19848 166 19888
rect 120 19816 166 19848
rect 120 19780 126 19816
rect 160 19780 166 19816
rect 120 19746 166 19780
rect 120 19710 126 19746
rect 160 19710 166 19746
rect 120 19678 166 19710
rect 120 19638 126 19678
rect 160 19638 166 19678
rect 120 19610 166 19638
rect 120 19566 126 19610
rect 160 19566 166 19610
rect 120 19542 166 19566
rect 120 19494 126 19542
rect 160 19494 166 19542
rect 120 19474 166 19494
rect 120 19422 126 19474
rect 160 19422 166 19474
rect 120 19406 166 19422
rect 120 19350 126 19406
rect 160 19350 166 19406
rect 120 19338 166 19350
rect 120 19278 126 19338
rect 160 19278 166 19338
rect 120 19270 166 19278
rect 120 19206 126 19270
rect 160 19206 166 19270
rect 120 19202 166 19206
rect 120 19100 126 19202
rect 160 19100 166 19202
rect 120 19096 166 19100
rect 120 19032 126 19096
rect 160 19032 166 19096
rect 120 19024 166 19032
rect 120 18964 126 19024
rect 160 18964 166 19024
rect 120 18952 166 18964
rect 120 18896 126 18952
rect 160 18896 166 18952
rect 120 18880 166 18896
rect 120 18828 126 18880
rect 160 18828 166 18880
rect 120 18808 166 18828
rect 120 18760 126 18808
rect 160 18760 166 18808
rect 120 18736 166 18760
rect 120 18692 126 18736
rect 160 18692 166 18736
rect 120 18664 166 18692
rect 120 18624 126 18664
rect 160 18624 166 18664
rect 120 18592 166 18624
rect 120 18556 126 18592
rect 160 18556 166 18592
rect 120 18522 166 18556
rect 120 18486 126 18522
rect 160 18486 166 18522
rect 120 18454 166 18486
rect 120 18414 126 18454
rect 160 18414 166 18454
rect 120 18386 166 18414
rect 120 18342 126 18386
rect 160 18342 166 18386
rect 120 18318 166 18342
rect 120 18270 126 18318
rect 160 18270 166 18318
rect 120 18250 166 18270
rect 120 18198 126 18250
rect 160 18198 166 18250
rect 120 18182 166 18198
rect 120 18126 126 18182
rect 160 18126 166 18182
rect 120 18114 166 18126
rect 120 18054 126 18114
rect 160 18054 166 18114
rect 120 18046 166 18054
rect 120 17982 126 18046
rect 160 17982 166 18046
rect 120 17978 166 17982
rect 120 17876 126 17978
rect 160 17876 166 17978
rect 120 17872 166 17876
rect 120 17808 126 17872
rect 160 17808 166 17872
rect 120 17800 166 17808
rect 120 17740 126 17800
rect 160 17740 166 17800
rect 120 17728 166 17740
rect 120 17672 126 17728
rect 160 17672 166 17728
rect 120 17656 166 17672
rect 120 17604 126 17656
rect 160 17604 166 17656
rect 120 17584 166 17604
rect 120 17536 126 17584
rect 160 17536 166 17584
rect 120 17512 166 17536
rect 120 17468 126 17512
rect 160 17468 166 17512
rect 120 17440 166 17468
rect 120 17400 126 17440
rect 160 17400 166 17440
rect 120 17368 166 17400
rect 120 17332 126 17368
rect 160 17332 166 17368
rect 120 17298 166 17332
rect 120 17262 126 17298
rect 160 17262 166 17298
rect 120 17230 166 17262
rect 120 17190 126 17230
rect 160 17190 166 17230
rect 120 17162 166 17190
rect 120 17118 126 17162
rect 160 17118 166 17162
rect 120 17094 166 17118
rect 120 17046 126 17094
rect 160 17046 166 17094
rect 120 17026 166 17046
rect 120 16974 126 17026
rect 160 16974 166 17026
rect 120 16958 166 16974
rect 120 16902 126 16958
rect 160 16902 166 16958
rect 120 16890 166 16902
rect 120 16830 126 16890
rect 160 16830 166 16890
rect 120 16822 166 16830
rect 120 16758 126 16822
rect 160 16758 166 16822
rect 120 16754 166 16758
rect 120 16652 126 16754
rect 160 16652 166 16754
rect 120 16648 166 16652
rect 120 16584 126 16648
rect 160 16584 166 16648
rect 120 16576 166 16584
rect 120 16516 126 16576
rect 160 16516 166 16576
rect 120 16504 166 16516
rect 120 16448 126 16504
rect 160 16448 166 16504
rect 120 16432 166 16448
rect 120 16380 126 16432
rect 160 16380 166 16432
rect 120 16360 166 16380
rect 120 16312 126 16360
rect 160 16312 166 16360
rect 120 16288 166 16312
rect 120 16244 126 16288
rect 160 16244 166 16288
rect 120 16216 166 16244
rect 120 16176 126 16216
rect 160 16176 166 16216
rect 120 16144 166 16176
rect 120 16108 126 16144
rect 160 16108 166 16144
rect 120 16074 166 16108
rect 120 16038 126 16074
rect 160 16038 166 16074
rect 120 16006 166 16038
rect 120 15966 126 16006
rect 160 15966 166 16006
rect 120 15938 166 15966
rect 120 15894 126 15938
rect 160 15894 166 15938
rect 120 15870 166 15894
rect 120 15822 126 15870
rect 160 15822 166 15870
rect 120 15802 166 15822
rect 120 15750 126 15802
rect 160 15750 166 15802
rect 120 15734 166 15750
rect 120 15678 126 15734
rect 160 15678 166 15734
rect 120 15666 166 15678
rect 120 15606 126 15666
rect 160 15606 166 15666
rect 120 15598 166 15606
rect 120 15534 126 15598
rect 160 15534 166 15598
rect 120 15530 166 15534
rect 120 15428 126 15530
rect 160 15428 166 15530
rect 120 15424 166 15428
rect 120 15360 126 15424
rect 160 15360 166 15424
rect 120 15352 166 15360
rect 120 15292 126 15352
rect 160 15292 166 15352
rect 120 15280 166 15292
rect 120 15224 126 15280
rect 160 15224 166 15280
rect 120 15208 166 15224
rect 120 15156 126 15208
rect 160 15156 166 15208
rect 120 15136 166 15156
rect 120 15088 126 15136
rect 160 15088 166 15136
rect 120 15064 166 15088
rect 120 15020 126 15064
rect 160 15020 166 15064
rect 120 14992 166 15020
rect 120 14952 126 14992
rect 160 14952 166 14992
rect 120 14920 166 14952
rect 120 14884 126 14920
rect 160 14884 166 14920
rect 120 14850 166 14884
rect 120 14814 126 14850
rect 160 14814 166 14850
rect 120 14782 166 14814
rect 120 14742 126 14782
rect 160 14742 166 14782
rect 120 14714 166 14742
rect 120 14670 126 14714
rect 160 14670 166 14714
rect 120 14646 166 14670
rect 120 14598 126 14646
rect 160 14598 166 14646
rect 120 14578 166 14598
rect 120 14526 126 14578
rect 160 14526 166 14578
rect 120 14510 166 14526
rect 120 14454 126 14510
rect 160 14454 166 14510
rect 120 14442 166 14454
rect 120 14382 126 14442
rect 160 14382 166 14442
rect 120 14374 166 14382
rect 120 14310 126 14374
rect 160 14310 166 14374
rect 120 14306 166 14310
rect 120 14204 126 14306
rect 160 14204 166 14306
rect 120 14200 166 14204
rect 120 14136 126 14200
rect 160 14136 166 14200
rect 120 14128 166 14136
rect 120 14068 126 14128
rect 160 14068 166 14128
rect 120 14056 166 14068
rect 120 14000 126 14056
rect 160 14000 166 14056
rect 120 13984 166 14000
rect 120 13932 126 13984
rect 160 13932 166 13984
rect 120 13912 166 13932
rect 120 13864 126 13912
rect 160 13864 166 13912
rect 120 13840 166 13864
rect 120 13796 126 13840
rect 160 13796 166 13840
rect 120 13768 166 13796
rect 120 13728 126 13768
rect 160 13728 166 13768
rect 120 13696 166 13728
rect 120 13660 126 13696
rect 160 13660 166 13696
rect 120 13626 166 13660
rect 120 13590 126 13626
rect 160 13590 166 13626
rect 120 13558 166 13590
rect 120 13518 126 13558
rect 160 13518 166 13558
rect 120 13490 166 13518
rect 120 13446 126 13490
rect 160 13446 166 13490
rect 120 13422 166 13446
rect 120 13374 126 13422
rect 160 13374 166 13422
rect 120 13354 166 13374
rect 120 13302 126 13354
rect 160 13302 166 13354
rect 120 13286 166 13302
rect 120 13230 126 13286
rect 160 13230 166 13286
rect 120 13218 166 13230
rect 120 13158 126 13218
rect 160 13158 166 13218
rect 120 13150 166 13158
rect 120 13086 126 13150
rect 160 13086 166 13150
rect 120 13082 166 13086
rect 120 12980 126 13082
rect 160 12980 166 13082
rect 120 12976 166 12980
rect 120 12912 126 12976
rect 160 12912 166 12976
rect 120 12904 166 12912
rect 120 12844 126 12904
rect 160 12844 166 12904
rect 120 12832 166 12844
rect 120 12776 126 12832
rect 160 12776 166 12832
rect 120 12760 166 12776
rect 120 12708 126 12760
rect 160 12708 166 12760
rect 120 12688 166 12708
rect 120 12640 126 12688
rect 160 12640 166 12688
rect 120 12616 166 12640
rect 120 12572 126 12616
rect 160 12572 166 12616
rect 120 12544 166 12572
rect 120 12504 126 12544
rect 160 12504 166 12544
rect 120 12472 166 12504
rect 120 12436 126 12472
rect 160 12436 166 12472
rect 120 12402 166 12436
rect 120 12366 126 12402
rect 160 12366 166 12402
rect 120 12334 166 12366
rect 120 12294 126 12334
rect 160 12294 166 12334
rect 120 12266 166 12294
rect 120 12222 126 12266
rect 160 12222 166 12266
rect 120 12198 166 12222
rect 120 12150 126 12198
rect 160 12150 166 12198
rect 120 12130 166 12150
rect 120 12078 126 12130
rect 160 12078 166 12130
rect 120 12062 166 12078
rect 120 12006 126 12062
rect 160 12006 166 12062
rect 120 11994 166 12006
rect 120 11934 126 11994
rect 160 11934 166 11994
rect 120 11926 166 11934
rect 120 11862 126 11926
rect 160 11862 166 11926
rect 120 11858 166 11862
rect 120 11756 126 11858
rect 160 11756 166 11858
rect 120 11752 166 11756
rect 120 11688 126 11752
rect 160 11688 166 11752
rect 120 11680 166 11688
rect 120 11620 126 11680
rect 160 11620 166 11680
rect 120 11608 166 11620
rect 120 11552 126 11608
rect 160 11552 166 11608
rect 120 11536 166 11552
rect 120 11484 126 11536
rect 160 11484 166 11536
rect 120 11464 166 11484
rect 120 11416 126 11464
rect 160 11416 166 11464
rect 120 11392 166 11416
rect 120 11348 126 11392
rect 160 11348 166 11392
rect 120 11320 166 11348
rect 120 11280 126 11320
rect 160 11280 166 11320
rect 120 11248 166 11280
rect 120 11212 126 11248
rect 160 11212 166 11248
rect 120 11178 166 11212
rect 120 11142 126 11178
rect 160 11142 166 11178
rect 120 11110 166 11142
rect 120 11070 126 11110
rect 160 11070 166 11110
rect 120 11042 166 11070
rect 120 10998 126 11042
rect 160 10998 166 11042
rect 120 10974 166 10998
rect 120 10926 126 10974
rect 160 10926 166 10974
rect 120 10906 166 10926
rect 120 10854 126 10906
rect 160 10854 166 10906
rect 120 10838 166 10854
rect 120 10782 126 10838
rect 160 10782 166 10838
rect 120 10770 166 10782
rect 120 10710 126 10770
rect 160 10710 166 10770
rect 120 10702 166 10710
rect 120 10638 126 10702
rect 160 10638 166 10702
rect 120 10634 166 10638
rect 120 10532 126 10634
rect 160 10532 166 10634
rect 120 10528 166 10532
rect 120 10464 126 10528
rect 160 10464 166 10528
rect 120 10456 166 10464
rect 120 10396 126 10456
rect 160 10396 166 10456
rect 120 10384 166 10396
rect 120 10328 126 10384
rect 160 10328 166 10384
rect 120 10312 166 10328
rect 120 10260 126 10312
rect 160 10260 166 10312
rect 120 10240 166 10260
rect 120 10192 126 10240
rect 160 10192 166 10240
rect 120 10168 166 10192
rect 120 10124 126 10168
rect 160 10124 166 10168
rect 120 10096 166 10124
rect 120 10056 126 10096
rect 160 10056 166 10096
rect 120 10024 166 10056
rect 120 9988 126 10024
rect 160 9988 166 10024
rect 120 9954 166 9988
rect 120 9918 126 9954
rect 160 9918 166 9954
rect 120 9886 166 9918
rect 120 9846 126 9886
rect 160 9846 166 9886
rect 120 9818 166 9846
rect 120 9774 126 9818
rect 160 9774 166 9818
rect 120 9750 166 9774
rect 120 9702 126 9750
rect 160 9702 166 9750
rect 120 9682 166 9702
rect 120 9630 126 9682
rect 160 9630 166 9682
rect 120 9614 166 9630
rect 120 9558 126 9614
rect 160 9558 166 9614
rect 120 9546 166 9558
rect 120 9486 126 9546
rect 160 9486 166 9546
rect 120 9478 166 9486
rect 120 9414 126 9478
rect 160 9414 166 9478
rect 120 9410 166 9414
rect 120 9308 126 9410
rect 160 9308 166 9410
rect 120 9304 166 9308
rect 120 9240 126 9304
rect 160 9240 166 9304
rect 120 9232 166 9240
rect 120 9172 126 9232
rect 160 9172 166 9232
rect 120 9160 166 9172
rect 120 9104 126 9160
rect 160 9104 166 9160
rect 120 9088 166 9104
rect 120 9036 126 9088
rect 160 9036 166 9088
rect 120 9016 166 9036
rect 120 8968 126 9016
rect 160 8968 166 9016
rect 120 8944 166 8968
rect 120 8900 126 8944
rect 160 8900 166 8944
rect 120 8872 166 8900
rect 120 8832 126 8872
rect 160 8832 166 8872
rect 120 8800 166 8832
rect 120 8764 126 8800
rect 160 8764 166 8800
rect 120 8730 166 8764
rect 120 8694 126 8730
rect 160 8694 166 8730
rect 120 8662 166 8694
rect 120 8622 126 8662
rect 160 8622 166 8662
rect 120 8594 166 8622
rect 120 8550 126 8594
rect 160 8550 166 8594
rect 120 8526 166 8550
rect 120 8478 126 8526
rect 160 8478 166 8526
rect 120 8458 166 8478
rect 120 8406 126 8458
rect 160 8406 166 8458
rect 120 8390 166 8406
rect 120 8334 126 8390
rect 160 8334 166 8390
rect 120 8322 166 8334
rect 120 8262 126 8322
rect 160 8262 166 8322
rect 120 8254 166 8262
rect 120 8190 126 8254
rect 160 8190 166 8254
rect 120 8186 166 8190
rect 120 8084 126 8186
rect 160 8084 166 8186
rect 120 8080 166 8084
rect 120 8016 126 8080
rect 160 8016 166 8080
rect 120 8008 166 8016
rect 120 7948 126 8008
rect 160 7948 166 8008
rect 120 7936 166 7948
rect 120 7880 126 7936
rect 160 7880 166 7936
rect 120 7864 166 7880
rect 120 7812 126 7864
rect 160 7812 166 7864
rect 120 7792 166 7812
rect 120 7744 126 7792
rect 160 7744 166 7792
rect 120 7720 166 7744
rect 120 7676 126 7720
rect 160 7676 166 7720
rect 120 7648 166 7676
rect 120 7608 126 7648
rect 160 7608 166 7648
rect 120 7576 166 7608
rect 120 7540 126 7576
rect 160 7540 166 7576
rect 120 7506 166 7540
rect 120 7470 126 7506
rect 160 7470 166 7506
rect 120 7438 166 7470
rect 120 7398 126 7438
rect 160 7398 166 7438
rect 120 7370 166 7398
rect 120 7326 126 7370
rect 160 7326 166 7370
rect 120 7302 166 7326
rect 120 7254 126 7302
rect 160 7254 166 7302
rect 120 7234 166 7254
rect 120 7182 126 7234
rect 160 7182 166 7234
rect 120 7166 166 7182
rect 120 7110 126 7166
rect 160 7110 166 7166
rect 120 7098 166 7110
rect 120 7038 126 7098
rect 160 7038 166 7098
rect 120 7030 166 7038
rect 120 6966 126 7030
rect 160 6966 166 7030
rect 120 6962 166 6966
rect 120 6860 126 6962
rect 160 6860 166 6962
rect 120 6856 166 6860
rect 120 6792 126 6856
rect 160 6792 166 6856
rect 120 6784 166 6792
rect 120 6724 126 6784
rect 160 6724 166 6784
rect 120 6712 166 6724
rect 120 6656 126 6712
rect 160 6656 166 6712
rect 120 6640 166 6656
rect 120 6588 126 6640
rect 160 6588 166 6640
rect 120 6568 166 6588
rect 120 6520 126 6568
rect 160 6520 166 6568
rect 120 6496 166 6520
rect 120 6452 126 6496
rect 160 6452 166 6496
rect 120 6424 166 6452
rect 120 6384 126 6424
rect 160 6384 166 6424
rect 120 6352 166 6384
rect 120 6316 126 6352
rect 160 6316 166 6352
rect 120 6282 166 6316
rect 120 6246 126 6282
rect 160 6246 166 6282
rect 120 6214 166 6246
rect 120 6174 126 6214
rect 160 6174 166 6214
rect 120 6146 166 6174
rect 120 6102 126 6146
rect 160 6102 166 6146
rect 120 6078 166 6102
rect 120 6030 126 6078
rect 160 6030 166 6078
rect 120 6010 166 6030
rect 120 5958 126 6010
rect 160 5958 166 6010
rect 120 5942 166 5958
rect 120 5886 126 5942
rect 160 5886 166 5942
rect 120 5874 166 5886
rect 120 5814 126 5874
rect 160 5814 166 5874
rect 120 5806 166 5814
rect 120 5742 126 5806
rect 160 5742 166 5806
rect 120 5738 166 5742
rect 120 5636 126 5738
rect 160 5636 166 5738
rect 120 5632 166 5636
rect 120 5568 126 5632
rect 160 5568 166 5632
rect 120 5560 166 5568
rect 120 5500 126 5560
rect 160 5500 166 5560
rect 120 5488 166 5500
rect 120 5432 126 5488
rect 160 5432 166 5488
rect 120 5416 166 5432
rect 120 5364 126 5416
rect 160 5364 166 5416
rect 120 5344 166 5364
rect 120 5296 126 5344
rect 160 5296 166 5344
rect 120 5272 166 5296
rect 120 5228 126 5272
rect 160 5228 166 5272
rect 120 5200 166 5228
rect 120 5160 126 5200
rect 160 5160 166 5200
rect 120 5128 166 5160
rect 120 5092 126 5128
rect 160 5092 166 5128
rect 120 5058 166 5092
rect 120 5022 126 5058
rect 160 5022 166 5058
rect 120 4990 166 5022
rect 120 4950 126 4990
rect 160 4950 166 4990
rect 120 4922 166 4950
rect 120 4878 126 4922
rect 160 4878 166 4922
rect 120 4854 166 4878
rect 120 4806 126 4854
rect 160 4806 166 4854
rect 120 4786 166 4806
rect 120 4734 126 4786
rect 160 4734 166 4786
rect 120 4718 166 4734
rect 120 4662 126 4718
rect 160 4662 166 4718
rect 120 4650 166 4662
rect 120 4590 126 4650
rect 160 4590 166 4650
rect 120 4582 166 4590
rect 120 4518 126 4582
rect 160 4518 166 4582
rect 120 4514 166 4518
rect 120 4412 126 4514
rect 160 4412 166 4514
rect 120 4408 166 4412
rect 120 4344 126 4408
rect 160 4344 166 4408
rect 120 4336 166 4344
rect 120 4276 126 4336
rect 160 4276 166 4336
rect 120 4264 166 4276
rect 120 4208 126 4264
rect 160 4208 166 4264
rect 120 4192 166 4208
rect 120 4140 126 4192
rect 160 4140 166 4192
rect 120 4120 166 4140
rect 120 4072 126 4120
rect 160 4072 166 4120
rect 120 4048 166 4072
rect 120 4004 126 4048
rect 160 4004 166 4048
rect 120 3976 166 4004
rect 120 3936 126 3976
rect 160 3936 166 3976
rect 120 3904 166 3936
rect 120 3868 126 3904
rect 160 3868 166 3904
rect 120 3834 166 3868
rect 120 3798 126 3834
rect 160 3798 166 3834
rect 120 3766 166 3798
rect 120 3726 126 3766
rect 160 3726 166 3766
rect 120 3698 166 3726
rect 120 3654 126 3698
rect 160 3654 166 3698
rect 120 3630 166 3654
rect 120 3582 126 3630
rect 160 3582 166 3630
rect 120 3562 166 3582
rect 120 3510 126 3562
rect 160 3510 166 3562
rect 120 3494 166 3510
rect 120 3438 126 3494
rect 160 3438 166 3494
rect 120 3426 166 3438
rect 120 3366 126 3426
rect 160 3366 166 3426
rect 120 3358 166 3366
rect 120 3294 126 3358
rect 160 3294 166 3358
rect 120 3290 166 3294
rect 120 3188 126 3290
rect 160 3188 166 3290
rect 120 3184 166 3188
rect 120 3120 126 3184
rect 160 3120 166 3184
rect 120 3112 166 3120
rect 120 3052 126 3112
rect 160 3052 166 3112
rect 120 3040 166 3052
rect 120 2984 126 3040
rect 160 2984 166 3040
rect 120 2968 166 2984
rect 120 2916 126 2968
rect 160 2916 166 2968
rect 120 2896 166 2916
rect 120 2848 126 2896
rect 160 2848 166 2896
rect 120 2824 166 2848
rect 120 2780 126 2824
rect 160 2780 166 2824
rect 120 2752 166 2780
rect 120 2712 126 2752
rect 160 2712 166 2752
rect 120 2680 166 2712
rect 120 2644 126 2680
rect 160 2644 166 2680
rect 120 2610 166 2644
rect 120 2574 126 2610
rect 160 2574 166 2610
rect 120 2542 166 2574
rect 120 2502 126 2542
rect 160 2502 166 2542
rect 120 2474 166 2502
rect 120 2430 126 2474
rect 160 2430 166 2474
rect 120 2406 166 2430
rect 120 2358 126 2406
rect 160 2358 166 2406
rect 120 2338 166 2358
rect 120 2286 126 2338
rect 160 2286 166 2338
rect 120 2270 166 2286
rect 120 2214 126 2270
rect 160 2214 166 2270
rect 120 2202 166 2214
rect 120 2142 126 2202
rect 160 2142 166 2202
rect 120 2134 166 2142
rect 120 2070 126 2134
rect 160 2070 166 2134
rect 120 2066 166 2070
rect 120 1964 126 2066
rect 160 1964 166 2066
rect 120 1960 166 1964
rect 120 1896 126 1960
rect 160 1896 166 1960
rect 120 1888 166 1896
rect 120 1828 126 1888
rect 160 1828 166 1888
rect 120 1816 166 1828
rect 120 1760 126 1816
rect 160 1760 166 1816
rect 120 1744 166 1760
rect 120 1692 126 1744
rect 160 1692 166 1744
rect 120 1672 166 1692
rect 120 1624 126 1672
rect 160 1624 166 1672
rect 120 1600 166 1624
rect 120 1556 126 1600
rect 160 1556 166 1600
rect 120 1528 166 1556
rect 120 1488 126 1528
rect 160 1488 166 1528
rect 120 1456 166 1488
rect 120 1420 126 1456
rect 160 1420 166 1456
rect 120 1386 166 1420
rect 120 1350 126 1386
rect 160 1350 166 1386
rect 120 1318 166 1350
rect 120 1278 126 1318
rect 160 1278 166 1318
rect 120 1250 166 1278
rect 120 1206 126 1250
rect 160 1206 166 1250
rect 120 1182 166 1206
rect 120 1134 126 1182
rect 160 1134 166 1182
rect 120 1114 166 1134
rect 120 1062 126 1114
rect 160 1062 166 1114
rect 120 1046 166 1062
rect 120 990 126 1046
rect 160 990 166 1046
rect 120 978 166 990
rect 120 918 126 978
rect 160 918 166 978
rect 120 910 166 918
rect 120 846 126 910
rect 160 846 166 910
rect 120 842 166 846
rect 120 740 126 842
rect 160 740 166 842
rect 120 736 166 740
rect 120 672 126 736
rect 160 672 166 736
rect 120 664 166 672
rect 120 604 126 664
rect 160 604 166 664
rect 120 592 166 604
rect 120 536 126 592
rect 160 536 166 592
rect 120 520 166 536
rect 373 39178 3083 39191
rect 373 39144 462 39178
rect 499 39144 533 39178
rect 572 39144 601 39178
rect 635 39144 648 39178
rect 703 39144 720 39178
rect 771 39144 792 39178
rect 839 39144 864 39178
rect 907 39144 936 39178
rect 975 39144 1008 39178
rect 1043 39144 1077 39178
rect 1114 39144 1145 39178
rect 1186 39144 1213 39178
rect 1258 39144 1281 39178
rect 1330 39144 1349 39178
rect 1402 39144 1417 39178
rect 1474 39144 1485 39178
rect 1546 39144 1553 39178
rect 1618 39144 1621 39178
rect 1655 39144 1656 39178
rect 1723 39144 1728 39178
rect 1791 39144 1800 39178
rect 1859 39144 1872 39178
rect 1927 39144 1944 39178
rect 1995 39144 2016 39178
rect 2063 39144 2088 39178
rect 2131 39144 2161 39178
rect 2199 39144 2233 39178
rect 2268 39144 2301 39178
rect 2341 39144 2369 39178
rect 2414 39144 2437 39178
rect 2487 39144 2505 39178
rect 2560 39144 2573 39178
rect 2633 39144 2641 39178
rect 2706 39144 2709 39178
rect 2743 39144 2745 39178
rect 2811 39144 2818 39178
rect 2879 39144 2891 39178
rect 2947 39144 2964 39178
rect 3015 39144 3083 39178
rect 373 39131 3083 39144
rect 373 39123 433 39131
rect 373 39072 386 39123
rect 420 39072 433 39123
rect 373 39055 433 39072
rect 373 38999 386 39055
rect 420 38999 433 39055
rect 3023 39110 3083 39131
rect 3023 39072 3036 39110
rect 3070 39072 3083 39110
rect 576 39020 592 39054
rect 626 39020 662 39054
rect 696 39020 732 39054
rect 766 39020 802 39054
rect 836 39020 872 39054
rect 906 39020 942 39054
rect 976 39020 1012 39054
rect 1046 39020 1082 39054
rect 1116 39020 1152 39054
rect 1186 39020 1222 39054
rect 1256 39020 1292 39054
rect 1326 39020 1362 39054
rect 1396 39020 1432 39054
rect 1466 39020 1502 39054
rect 1536 39020 1572 39054
rect 1606 39020 1642 39054
rect 1676 39020 1712 39054
rect 1746 39020 1782 39054
rect 1816 39020 1852 39054
rect 1886 39020 1922 39054
rect 1956 39020 1992 39054
rect 2026 39020 2062 39054
rect 2096 39020 2132 39054
rect 2166 39020 2202 39054
rect 2236 39020 2272 39054
rect 2306 39020 2342 39054
rect 2376 39020 2412 39054
rect 2446 39020 2482 39054
rect 2516 39020 2552 39054
rect 2586 39020 2622 39054
rect 2656 39020 2692 39054
rect 2726 39020 2761 39054
rect 2795 39020 2830 39054
rect 2864 39020 2880 39054
rect 3023 39042 3083 39072
rect 373 38987 433 38999
rect 373 38926 386 38987
rect 420 38926 433 38987
rect 3023 39000 3036 39042
rect 3070 39000 3083 39042
rect 3023 38974 3083 39000
rect 373 38919 433 38926
rect 373 38853 386 38919
rect 420 38853 433 38919
rect 373 38851 433 38853
rect 373 38817 386 38851
rect 420 38817 433 38851
rect 373 38814 433 38817
rect 373 38749 386 38814
rect 420 38749 433 38814
rect 373 38741 433 38749
rect 373 38681 386 38741
rect 420 38681 433 38741
rect 373 38668 433 38681
rect 373 38613 386 38668
rect 420 38613 433 38668
rect 373 38595 433 38613
rect 373 38545 386 38595
rect 420 38545 433 38595
rect 373 38522 433 38545
rect 373 38477 386 38522
rect 420 38477 433 38522
rect 373 38449 433 38477
rect 373 38409 386 38449
rect 420 38409 433 38449
rect 373 38376 433 38409
rect 373 38341 386 38376
rect 420 38341 433 38376
rect 373 38307 433 38341
rect 373 38269 386 38307
rect 420 38269 433 38307
rect 373 38239 433 38269
rect 373 38196 386 38239
rect 420 38196 433 38239
rect 373 38171 433 38196
rect 373 38123 386 38171
rect 420 38123 433 38171
rect 373 38103 433 38123
rect 373 38050 386 38103
rect 420 38050 433 38103
rect 373 38035 433 38050
rect 373 37977 386 38035
rect 420 37977 433 38035
rect 373 37967 433 37977
rect 373 37904 386 37967
rect 420 37904 433 37967
rect 373 37899 433 37904
rect 373 37797 386 37899
rect 420 37797 433 37899
rect 373 37792 433 37797
rect 373 37729 386 37792
rect 420 37729 433 37792
rect 373 37719 433 37729
rect 373 37661 386 37719
rect 420 37661 433 37719
rect 373 37647 433 37661
rect 373 37593 386 37647
rect 420 37593 433 37647
rect 373 37575 433 37593
rect 373 37525 386 37575
rect 420 37525 433 37575
rect 373 37503 433 37525
rect 373 37457 386 37503
rect 420 37457 433 37503
rect 373 37431 433 37457
rect 373 37389 386 37431
rect 420 37389 433 37431
rect 373 37359 433 37389
rect 373 37321 386 37359
rect 420 37321 433 37359
rect 373 37287 433 37321
rect 373 37253 386 37287
rect 420 37253 433 37287
rect 373 37219 433 37253
rect 373 37181 386 37219
rect 420 37181 433 37219
rect 373 37151 433 37181
rect 373 37109 386 37151
rect 420 37109 433 37151
rect 373 37083 433 37109
rect 373 37037 386 37083
rect 420 37037 433 37083
rect 373 37015 433 37037
rect 531 38891 565 38930
rect 531 38818 565 38857
rect 531 38745 565 38784
rect 531 38672 565 38711
rect 531 38599 565 38638
rect 531 38526 565 38565
rect 531 38453 565 38492
rect 531 38380 565 38419
rect 531 38307 565 38346
rect 531 38234 565 38273
rect 531 38161 565 38200
rect 531 38088 565 38127
rect 531 38014 565 38054
rect 531 37940 565 37980
rect 531 37866 565 37906
rect 531 37792 565 37832
rect 531 37718 565 37758
rect 531 37644 565 37684
rect 531 37570 565 37610
rect 531 37496 565 37536
rect 531 37422 565 37462
rect 531 37348 565 37388
rect 531 37274 565 37314
rect 531 37200 565 37240
rect 531 37126 565 37166
rect 531 37052 565 37092
rect 767 38891 801 38930
rect 767 38818 801 38857
rect 767 38745 801 38784
rect 767 38672 801 38711
rect 767 38599 801 38638
rect 767 38526 801 38565
rect 767 38453 801 38492
rect 767 38380 801 38419
rect 767 38307 801 38346
rect 767 38234 801 38273
rect 767 38161 801 38200
rect 767 38088 801 38127
rect 767 38014 801 38054
rect 767 37940 801 37980
rect 767 37866 801 37906
rect 767 37792 801 37832
rect 767 37718 801 37758
rect 767 37644 801 37684
rect 767 37570 801 37610
rect 767 37496 801 37536
rect 767 37422 801 37462
rect 767 37348 801 37388
rect 767 37274 801 37314
rect 767 37200 801 37240
rect 767 37126 801 37166
rect 767 37052 801 37092
rect 1003 38891 1037 38930
rect 1003 38818 1037 38857
rect 1003 38745 1037 38784
rect 1003 38672 1037 38711
rect 1003 38599 1037 38638
rect 1003 38526 1037 38565
rect 1003 38453 1037 38492
rect 1003 38380 1037 38419
rect 1003 38307 1037 38346
rect 1003 38234 1037 38273
rect 1003 38161 1037 38200
rect 1003 38088 1037 38127
rect 1003 38014 1037 38054
rect 1003 37940 1037 37980
rect 1003 37866 1037 37906
rect 1003 37792 1037 37832
rect 1003 37718 1037 37758
rect 1003 37644 1037 37684
rect 1003 37570 1037 37610
rect 1003 37496 1037 37536
rect 1003 37422 1037 37462
rect 1003 37348 1037 37388
rect 1003 37274 1037 37314
rect 1003 37200 1037 37240
rect 1003 37126 1037 37166
rect 1003 37052 1037 37092
rect 1239 38891 1273 38930
rect 1239 38818 1273 38857
rect 1239 38745 1273 38784
rect 1239 38672 1273 38711
rect 1239 38599 1273 38638
rect 1239 38526 1273 38565
rect 1239 38453 1273 38492
rect 1239 38380 1273 38419
rect 1239 38307 1273 38346
rect 1239 38234 1273 38273
rect 1239 38161 1273 38200
rect 1239 38088 1273 38127
rect 1239 38014 1273 38054
rect 1239 37940 1273 37980
rect 1239 37866 1273 37906
rect 1239 37792 1273 37832
rect 1239 37718 1273 37758
rect 1239 37644 1273 37684
rect 1239 37570 1273 37610
rect 1239 37496 1273 37536
rect 1239 37422 1273 37462
rect 1239 37348 1273 37388
rect 1239 37274 1273 37314
rect 1239 37200 1273 37240
rect 1239 37126 1273 37166
rect 1239 37052 1273 37092
rect 1475 38891 1509 38930
rect 1475 38818 1509 38857
rect 1475 38745 1509 38784
rect 1475 38672 1509 38711
rect 1475 38599 1509 38638
rect 1475 38526 1509 38565
rect 1475 38453 1509 38492
rect 1475 38380 1509 38419
rect 1475 38307 1509 38346
rect 1475 38234 1509 38273
rect 1475 38161 1509 38200
rect 1475 38088 1509 38127
rect 1475 38014 1509 38054
rect 1475 37940 1509 37980
rect 1475 37866 1509 37906
rect 1475 37792 1509 37832
rect 1475 37718 1509 37758
rect 1475 37644 1509 37684
rect 1475 37570 1509 37610
rect 1475 37496 1509 37536
rect 1475 37422 1509 37462
rect 1475 37348 1509 37388
rect 1475 37274 1509 37314
rect 1475 37200 1509 37240
rect 1475 37126 1509 37166
rect 1475 37052 1509 37092
rect 1711 38891 1745 38930
rect 1711 38818 1745 38857
rect 1711 38745 1745 38784
rect 1711 38672 1745 38711
rect 1711 38599 1745 38638
rect 1711 38526 1745 38565
rect 1711 38453 1745 38492
rect 1711 38380 1745 38419
rect 1711 38307 1745 38346
rect 1711 38234 1745 38273
rect 1711 38161 1745 38200
rect 1711 38088 1745 38127
rect 1711 38014 1745 38054
rect 1711 37940 1745 37980
rect 1711 37866 1745 37906
rect 1711 37792 1745 37832
rect 1711 37718 1745 37758
rect 1711 37644 1745 37684
rect 1711 37570 1745 37610
rect 1711 37496 1745 37536
rect 1711 37422 1745 37462
rect 1711 37348 1745 37388
rect 1711 37274 1745 37314
rect 1711 37200 1745 37240
rect 1711 37126 1745 37166
rect 1711 37052 1745 37092
rect 1947 38891 1981 38930
rect 1947 38818 1981 38857
rect 1947 38745 1981 38784
rect 1947 38672 1981 38711
rect 1947 38599 1981 38638
rect 1947 38526 1981 38565
rect 1947 38453 1981 38492
rect 1947 38380 1981 38419
rect 1947 38307 1981 38346
rect 1947 38234 1981 38273
rect 1947 38161 1981 38200
rect 1947 38088 1981 38127
rect 1947 38014 1981 38054
rect 1947 37940 1981 37980
rect 1947 37866 1981 37906
rect 1947 37792 1981 37832
rect 1947 37718 1981 37758
rect 1947 37644 1981 37684
rect 1947 37570 1981 37610
rect 1947 37496 1981 37536
rect 1947 37422 1981 37462
rect 1947 37348 1981 37388
rect 1947 37274 1981 37314
rect 1947 37200 1981 37240
rect 1947 37126 1981 37166
rect 1947 37052 1981 37092
rect 2183 38891 2217 38930
rect 2183 38818 2217 38857
rect 2183 38745 2217 38784
rect 2183 38672 2217 38711
rect 2183 38599 2217 38638
rect 2183 38526 2217 38565
rect 2183 38453 2217 38492
rect 2183 38380 2217 38419
rect 2183 38307 2217 38346
rect 2183 38234 2217 38273
rect 2183 38161 2217 38200
rect 2183 38088 2217 38127
rect 2183 38014 2217 38054
rect 2183 37940 2217 37980
rect 2183 37866 2217 37906
rect 2183 37792 2217 37832
rect 2183 37718 2217 37758
rect 2183 37644 2217 37684
rect 2183 37570 2217 37610
rect 2183 37496 2217 37536
rect 2183 37422 2217 37462
rect 2183 37348 2217 37388
rect 2183 37274 2217 37314
rect 2183 37200 2217 37240
rect 2183 37126 2217 37166
rect 2183 37052 2217 37092
rect 2419 38891 2453 38930
rect 2419 38818 2453 38857
rect 2419 38745 2453 38784
rect 2419 38672 2453 38711
rect 2419 38599 2453 38638
rect 2419 38526 2453 38565
rect 2419 38453 2453 38492
rect 2419 38380 2453 38419
rect 2419 38307 2453 38346
rect 2419 38234 2453 38273
rect 2419 38161 2453 38200
rect 2419 38088 2453 38127
rect 2419 38014 2453 38054
rect 2419 37940 2453 37980
rect 2419 37866 2453 37906
rect 2419 37792 2453 37832
rect 2419 37718 2453 37758
rect 2419 37644 2453 37684
rect 2419 37570 2453 37610
rect 2419 37496 2453 37536
rect 2419 37422 2453 37462
rect 2419 37348 2453 37388
rect 2419 37274 2453 37314
rect 2419 37200 2453 37240
rect 2419 37126 2453 37166
rect 2419 37052 2453 37092
rect 2655 38891 2689 38930
rect 2655 38818 2689 38857
rect 2655 38745 2689 38784
rect 2655 38672 2689 38711
rect 2655 38599 2689 38638
rect 2655 38526 2689 38565
rect 2655 38453 2689 38492
rect 2655 38380 2689 38419
rect 2655 38307 2689 38346
rect 2655 38234 2689 38273
rect 2655 38161 2689 38200
rect 2655 38088 2689 38127
rect 2655 38014 2689 38054
rect 2655 37940 2689 37980
rect 2655 37866 2689 37906
rect 2655 37792 2689 37832
rect 2655 37718 2689 37758
rect 2655 37644 2689 37684
rect 2655 37570 2689 37610
rect 2655 37496 2689 37536
rect 2655 37422 2689 37462
rect 2655 37348 2689 37388
rect 2655 37274 2689 37314
rect 2655 37200 2689 37240
rect 2655 37126 2689 37166
rect 2655 37052 2689 37092
rect 2891 38891 2925 38930
rect 2891 38818 2925 38857
rect 2891 38745 2925 38784
rect 2891 38672 2925 38711
rect 2891 38599 2925 38638
rect 2891 38526 2925 38565
rect 2891 38453 2925 38492
rect 2891 38380 2925 38419
rect 2891 38307 2925 38346
rect 2891 38234 2925 38273
rect 2891 38161 2925 38200
rect 2891 38088 2925 38127
rect 2891 38014 2925 38054
rect 2891 37940 2925 37980
rect 2891 37866 2925 37906
rect 2891 37792 2925 37832
rect 2891 37718 2925 37758
rect 2891 37644 2925 37684
rect 2891 37570 2925 37610
rect 2891 37496 2925 37536
rect 2891 37422 2925 37462
rect 2891 37348 2925 37388
rect 2891 37274 2925 37314
rect 2891 37200 2925 37240
rect 2891 37126 2925 37166
rect 2891 37052 2925 37092
rect 3023 38928 3036 38974
rect 3070 38928 3083 38974
rect 3023 38906 3083 38928
rect 3023 38856 3036 38906
rect 3070 38856 3083 38906
rect 3023 38838 3083 38856
rect 3023 38784 3036 38838
rect 3070 38784 3083 38838
rect 3023 38770 3083 38784
rect 3023 38712 3036 38770
rect 3070 38712 3083 38770
rect 3023 38702 3083 38712
rect 3023 38640 3036 38702
rect 3070 38640 3083 38702
rect 3023 38634 3083 38640
rect 3023 38568 3036 38634
rect 3070 38568 3083 38634
rect 3023 38566 3083 38568
rect 3023 38532 3036 38566
rect 3070 38532 3083 38566
rect 3023 38530 3083 38532
rect 3023 38464 3036 38530
rect 3070 38464 3083 38530
rect 3023 38458 3083 38464
rect 3023 38396 3036 38458
rect 3070 38396 3083 38458
rect 3023 38386 3083 38396
rect 3023 38328 3036 38386
rect 3070 38328 3083 38386
rect 3023 38314 3083 38328
rect 3023 38260 3036 38314
rect 3070 38260 3083 38314
rect 3023 38242 3083 38260
rect 3023 38192 3036 38242
rect 3070 38192 3083 38242
rect 3023 38170 3083 38192
rect 3023 38124 3036 38170
rect 3070 38124 3083 38170
rect 3023 38098 3083 38124
rect 3023 38056 3036 38098
rect 3070 38056 3083 38098
rect 3023 38026 3083 38056
rect 3023 37988 3036 38026
rect 3070 37988 3083 38026
rect 3023 37954 3083 37988
rect 3023 37920 3036 37954
rect 3070 37920 3083 37954
rect 3023 37886 3083 37920
rect 3023 37848 3036 37886
rect 3070 37848 3083 37886
rect 3023 37818 3083 37848
rect 3023 37776 3036 37818
rect 3070 37776 3083 37818
rect 3023 37750 3083 37776
rect 3023 37704 3036 37750
rect 3070 37704 3083 37750
rect 3023 37682 3083 37704
rect 3023 37632 3036 37682
rect 3070 37632 3083 37682
rect 3023 37614 3083 37632
rect 3023 37560 3036 37614
rect 3070 37560 3083 37614
rect 3023 37546 3083 37560
rect 3023 37488 3036 37546
rect 3070 37488 3083 37546
rect 3023 37478 3083 37488
rect 3023 37416 3036 37478
rect 3070 37416 3083 37478
rect 3023 37410 3083 37416
rect 3023 37344 3036 37410
rect 3070 37344 3083 37410
rect 3023 37342 3083 37344
rect 3023 37308 3036 37342
rect 3070 37308 3083 37342
rect 3023 37306 3083 37308
rect 3023 37240 3036 37306
rect 3070 37240 3083 37306
rect 3023 37234 3083 37240
rect 3023 37172 3036 37234
rect 3070 37172 3083 37234
rect 3023 37162 3083 37172
rect 3023 37104 3036 37162
rect 3070 37104 3083 37162
rect 3023 37090 3083 37104
rect 3023 37036 3036 37090
rect 3070 37036 3083 37090
rect 3023 37018 3083 37036
rect 373 36965 386 37015
rect 420 36965 433 37015
rect 373 36947 433 36965
rect 373 36893 386 36947
rect 420 36893 433 36947
rect 3023 36968 3036 37018
rect 3070 36968 3083 37018
rect 3023 36946 3083 36968
rect 373 36879 433 36893
rect 576 36890 592 36924
rect 659 36890 662 36924
rect 696 36890 700 36924
rect 766 36890 775 36924
rect 836 36890 850 36924
rect 906 36890 925 36924
rect 976 36890 1000 36924
rect 1046 36890 1075 36924
rect 1116 36890 1150 36924
rect 1186 36890 1222 36924
rect 1259 36890 1292 36924
rect 1334 36890 1362 36924
rect 1409 36890 1432 36924
rect 1484 36890 1502 36924
rect 1559 36890 1572 36924
rect 1634 36890 1642 36924
rect 1708 36890 1712 36924
rect 1746 36890 1748 36924
rect 1816 36890 1822 36924
rect 1886 36890 1896 36924
rect 1956 36890 1970 36924
rect 2026 36890 2044 36924
rect 2096 36890 2118 36924
rect 2166 36890 2192 36924
rect 2236 36890 2266 36924
rect 2306 36890 2340 36924
rect 2376 36890 2412 36924
rect 2448 36890 2482 36924
rect 2522 36890 2552 36924
rect 2596 36890 2622 36924
rect 2670 36890 2692 36924
rect 2744 36890 2761 36924
rect 2818 36890 2830 36924
rect 2864 36890 2880 36924
rect 3023 36900 3036 36946
rect 3070 36900 3083 36946
rect 373 36821 386 36879
rect 420 36821 433 36879
rect 3023 36874 3083 36900
rect 3023 36832 3036 36874
rect 3070 36832 3083 36874
rect 373 36811 433 36821
rect 373 36749 386 36811
rect 420 36749 433 36811
rect 373 36743 433 36749
rect 373 36677 386 36743
rect 420 36677 433 36743
rect 373 36675 433 36677
rect 373 36641 386 36675
rect 420 36641 433 36675
rect 373 36639 433 36641
rect 373 36573 386 36639
rect 420 36573 433 36639
rect 373 36567 433 36573
rect 373 36505 386 36567
rect 420 36505 433 36567
rect 373 36495 433 36505
rect 373 36437 386 36495
rect 420 36437 433 36495
rect 373 36423 433 36437
rect 373 36369 386 36423
rect 420 36369 433 36423
rect 373 36351 433 36369
rect 373 36301 386 36351
rect 420 36301 433 36351
rect 373 36279 433 36301
rect 373 36233 386 36279
rect 420 36233 433 36279
rect 373 36207 433 36233
rect 373 36165 386 36207
rect 420 36165 433 36207
rect 373 36135 433 36165
rect 373 36097 386 36135
rect 420 36097 433 36135
rect 373 36063 433 36097
rect 373 36029 386 36063
rect 420 36029 433 36063
rect 373 35995 433 36029
rect 373 35957 386 35995
rect 420 35957 433 35995
rect 373 35927 433 35957
rect 373 35885 386 35927
rect 420 35885 433 35927
rect 373 35859 433 35885
rect 373 35813 386 35859
rect 420 35813 433 35859
rect 373 35791 433 35813
rect 373 35741 386 35791
rect 420 35741 433 35791
rect 373 35723 433 35741
rect 373 35669 386 35723
rect 420 35669 433 35723
rect 373 35655 433 35669
rect 373 35597 386 35655
rect 420 35597 433 35655
rect 373 35587 433 35597
rect 373 35525 386 35587
rect 420 35525 433 35587
rect 373 35519 433 35525
rect 373 35453 386 35519
rect 420 35453 433 35519
rect 373 35451 433 35453
rect 373 35417 386 35451
rect 420 35417 433 35451
rect 373 35415 433 35417
rect 373 35349 386 35415
rect 420 35349 433 35415
rect 373 35343 433 35349
rect 373 35281 386 35343
rect 420 35281 433 35343
rect 373 35271 433 35281
rect 373 35213 386 35271
rect 420 35213 433 35271
rect 373 35199 433 35213
rect 373 35145 386 35199
rect 420 35145 433 35199
rect 373 35127 433 35145
rect 373 35077 386 35127
rect 420 35077 433 35127
rect 373 35055 433 35077
rect 373 35009 386 35055
rect 420 35009 433 35055
rect 373 34983 433 35009
rect 373 34941 386 34983
rect 420 34941 433 34983
rect 373 34911 433 34941
rect 373 34873 386 34911
rect 420 34873 433 34911
rect 531 36749 565 36788
rect 531 36676 565 36715
rect 531 36603 565 36642
rect 531 36530 565 36569
rect 531 36457 565 36496
rect 531 36384 565 36423
rect 531 36311 565 36350
rect 531 36238 565 36277
rect 531 36165 565 36204
rect 531 36092 565 36131
rect 531 36019 565 36058
rect 531 35946 565 35985
rect 531 35872 565 35912
rect 531 35798 565 35838
rect 531 35724 565 35764
rect 531 35650 565 35690
rect 531 35576 565 35616
rect 531 35502 565 35542
rect 531 35428 565 35468
rect 531 35354 565 35394
rect 531 35280 565 35320
rect 531 35206 565 35246
rect 531 35132 565 35172
rect 531 35058 565 35098
rect 531 34984 565 35024
rect 531 34910 565 34950
rect 767 36749 801 36788
rect 767 36676 801 36715
rect 767 36603 801 36642
rect 767 36530 801 36569
rect 767 36457 801 36496
rect 767 36384 801 36423
rect 767 36311 801 36350
rect 767 36238 801 36277
rect 767 36165 801 36204
rect 767 36092 801 36131
rect 767 36019 801 36058
rect 767 35946 801 35985
rect 767 35872 801 35912
rect 767 35798 801 35838
rect 767 35724 801 35764
rect 767 35650 801 35690
rect 767 35576 801 35616
rect 767 35502 801 35542
rect 767 35428 801 35468
rect 767 35354 801 35394
rect 767 35280 801 35320
rect 767 35206 801 35246
rect 767 35132 801 35172
rect 767 35058 801 35098
rect 767 34984 801 35024
rect 767 34910 801 34950
rect 1003 36749 1037 36788
rect 1003 36676 1037 36715
rect 1003 36603 1037 36642
rect 1003 36530 1037 36569
rect 1003 36457 1037 36496
rect 1003 36384 1037 36423
rect 1003 36311 1037 36350
rect 1003 36238 1037 36277
rect 1003 36165 1037 36204
rect 1003 36092 1037 36131
rect 1003 36019 1037 36058
rect 1003 35946 1037 35985
rect 1003 35872 1037 35912
rect 1003 35798 1037 35838
rect 1003 35724 1037 35764
rect 1003 35650 1037 35690
rect 1003 35576 1037 35616
rect 1003 35502 1037 35542
rect 1003 35428 1037 35468
rect 1003 35354 1037 35394
rect 1003 35280 1037 35320
rect 1003 35206 1037 35246
rect 1003 35132 1037 35172
rect 1003 35058 1037 35098
rect 1003 34984 1037 35024
rect 1003 34910 1037 34950
rect 1239 36749 1273 36788
rect 1239 36676 1273 36715
rect 1239 36603 1273 36642
rect 1239 36530 1273 36569
rect 1239 36457 1273 36496
rect 1239 36384 1273 36423
rect 1239 36311 1273 36350
rect 1239 36238 1273 36277
rect 1239 36165 1273 36204
rect 1239 36092 1273 36131
rect 1239 36019 1273 36058
rect 1239 35946 1273 35985
rect 1239 35872 1273 35912
rect 1239 35798 1273 35838
rect 1239 35724 1273 35764
rect 1239 35650 1273 35690
rect 1239 35576 1273 35616
rect 1239 35502 1273 35542
rect 1239 35428 1273 35468
rect 1239 35354 1273 35394
rect 1239 35280 1273 35320
rect 1239 35206 1273 35246
rect 1239 35132 1273 35172
rect 1239 35058 1273 35098
rect 1239 34984 1273 35024
rect 1239 34910 1273 34950
rect 1475 36749 1509 36788
rect 1475 36676 1509 36715
rect 1475 36603 1509 36642
rect 1475 36530 1509 36569
rect 1475 36457 1509 36496
rect 1475 36384 1509 36423
rect 1475 36311 1509 36350
rect 1475 36238 1509 36277
rect 1475 36165 1509 36204
rect 1475 36092 1509 36131
rect 1475 36019 1509 36058
rect 1475 35946 1509 35985
rect 1475 35872 1509 35912
rect 1475 35798 1509 35838
rect 1475 35724 1509 35764
rect 1475 35650 1509 35690
rect 1475 35576 1509 35616
rect 1475 35502 1509 35542
rect 1475 35428 1509 35468
rect 1475 35354 1509 35394
rect 1475 35280 1509 35320
rect 1475 35206 1509 35246
rect 1475 35132 1509 35172
rect 1475 35058 1509 35098
rect 1475 34984 1509 35024
rect 1475 34910 1509 34950
rect 1711 36749 1745 36788
rect 1711 36676 1745 36715
rect 1711 36603 1745 36642
rect 1711 36530 1745 36569
rect 1711 36457 1745 36496
rect 1711 36384 1745 36423
rect 1711 36311 1745 36350
rect 1711 36238 1745 36277
rect 1711 36165 1745 36204
rect 1711 36092 1745 36131
rect 1711 36019 1745 36058
rect 1711 35946 1745 35985
rect 1711 35872 1745 35912
rect 1711 35798 1745 35838
rect 1711 35724 1745 35764
rect 1711 35650 1745 35690
rect 1711 35576 1745 35616
rect 1711 35502 1745 35542
rect 1711 35428 1745 35468
rect 1711 35354 1745 35394
rect 1711 35280 1745 35320
rect 1711 35206 1745 35246
rect 1711 35132 1745 35172
rect 1711 35058 1745 35098
rect 1711 34984 1745 35024
rect 1711 34910 1745 34950
rect 1947 36749 1981 36788
rect 1947 36676 1981 36715
rect 1947 36603 1981 36642
rect 1947 36530 1981 36569
rect 1947 36457 1981 36496
rect 1947 36384 1981 36423
rect 1947 36311 1981 36350
rect 1947 36238 1981 36277
rect 1947 36165 1981 36204
rect 1947 36092 1981 36131
rect 1947 36019 1981 36058
rect 1947 35946 1981 35985
rect 1947 35872 1981 35912
rect 1947 35798 1981 35838
rect 1947 35724 1981 35764
rect 1947 35650 1981 35690
rect 1947 35576 1981 35616
rect 1947 35502 1981 35542
rect 1947 35428 1981 35468
rect 1947 35354 1981 35394
rect 1947 35280 1981 35320
rect 1947 35206 1981 35246
rect 1947 35132 1981 35172
rect 1947 35058 1981 35098
rect 1947 34984 1981 35024
rect 1947 34910 1981 34950
rect 2183 36749 2217 36788
rect 2183 36676 2217 36715
rect 2183 36603 2217 36642
rect 2183 36530 2217 36569
rect 2183 36457 2217 36496
rect 2183 36384 2217 36423
rect 2183 36311 2217 36350
rect 2183 36238 2217 36277
rect 2183 36165 2217 36204
rect 2183 36092 2217 36131
rect 2183 36019 2217 36058
rect 2183 35946 2217 35985
rect 2183 35872 2217 35912
rect 2183 35798 2217 35838
rect 2183 35724 2217 35764
rect 2183 35650 2217 35690
rect 2183 35576 2217 35616
rect 2183 35502 2217 35542
rect 2183 35428 2217 35468
rect 2183 35354 2217 35394
rect 2183 35280 2217 35320
rect 2183 35206 2217 35246
rect 2183 35132 2217 35172
rect 2183 35058 2217 35098
rect 2183 34984 2217 35024
rect 2183 34910 2217 34950
rect 2419 36749 2453 36788
rect 2419 36676 2453 36715
rect 2419 36603 2453 36642
rect 2419 36530 2453 36569
rect 2419 36457 2453 36496
rect 2419 36384 2453 36423
rect 2419 36311 2453 36350
rect 2419 36238 2453 36277
rect 2419 36165 2453 36204
rect 2419 36092 2453 36131
rect 2419 36019 2453 36058
rect 2419 35946 2453 35985
rect 2419 35872 2453 35912
rect 2419 35798 2453 35838
rect 2419 35724 2453 35764
rect 2419 35650 2453 35690
rect 2419 35576 2453 35616
rect 2419 35502 2453 35542
rect 2419 35428 2453 35468
rect 2419 35354 2453 35394
rect 2419 35280 2453 35320
rect 2419 35206 2453 35246
rect 2419 35132 2453 35172
rect 2419 35058 2453 35098
rect 2419 34984 2453 35024
rect 2419 34910 2453 34950
rect 2655 36749 2689 36788
rect 2655 36676 2689 36715
rect 2655 36603 2689 36642
rect 2655 36530 2689 36569
rect 2655 36457 2689 36496
rect 2655 36384 2689 36423
rect 2655 36311 2689 36350
rect 2655 36238 2689 36277
rect 2655 36165 2689 36204
rect 2655 36092 2689 36131
rect 2655 36019 2689 36058
rect 2655 35946 2689 35985
rect 2655 35872 2689 35912
rect 2655 35798 2689 35838
rect 2655 35724 2689 35764
rect 2655 35650 2689 35690
rect 2655 35576 2689 35616
rect 2655 35502 2689 35542
rect 2655 35428 2689 35468
rect 2655 35354 2689 35394
rect 2655 35280 2689 35320
rect 2655 35206 2689 35246
rect 2655 35132 2689 35172
rect 2655 35058 2689 35098
rect 2655 34984 2689 35024
rect 2655 34910 2689 34950
rect 2891 36749 2925 36788
rect 2891 36676 2925 36715
rect 2891 36603 2925 36642
rect 2891 36530 2925 36569
rect 2891 36457 2925 36496
rect 2891 36384 2925 36423
rect 2891 36311 2925 36350
rect 2891 36238 2925 36277
rect 2891 36165 2925 36204
rect 2891 36092 2925 36131
rect 2891 36019 2925 36058
rect 2891 35946 2925 35985
rect 2891 35872 2925 35912
rect 2891 35798 2925 35838
rect 2891 35724 2925 35764
rect 2891 35650 2925 35690
rect 2891 35576 2925 35616
rect 2891 35502 2925 35542
rect 2891 35428 2925 35468
rect 2891 35354 2925 35394
rect 2891 35280 2925 35320
rect 2891 35206 2925 35246
rect 2891 35132 2925 35172
rect 2891 35058 2925 35098
rect 2891 34984 2925 35024
rect 2891 34910 2925 34950
rect 3023 36802 3083 36832
rect 3023 36764 3036 36802
rect 3070 36764 3083 36802
rect 3023 36730 3083 36764
rect 3023 36696 3036 36730
rect 3070 36696 3083 36730
rect 3023 36662 3083 36696
rect 3023 36624 3036 36662
rect 3070 36624 3083 36662
rect 3023 36594 3083 36624
rect 3023 36552 3036 36594
rect 3070 36552 3083 36594
rect 3023 36526 3083 36552
rect 3023 36480 3036 36526
rect 3070 36480 3083 36526
rect 3023 36458 3083 36480
rect 3023 36408 3036 36458
rect 3070 36408 3083 36458
rect 3023 36390 3083 36408
rect 3023 36336 3036 36390
rect 3070 36336 3083 36390
rect 3023 36322 3083 36336
rect 3023 36264 3036 36322
rect 3070 36264 3083 36322
rect 3023 36254 3083 36264
rect 3023 36192 3036 36254
rect 3070 36192 3083 36254
rect 3023 36186 3083 36192
rect 3023 36120 3036 36186
rect 3070 36120 3083 36186
rect 3023 36118 3083 36120
rect 3023 36084 3036 36118
rect 3070 36084 3083 36118
rect 3023 36082 3083 36084
rect 3023 36016 3036 36082
rect 3070 36016 3083 36082
rect 3023 36010 3083 36016
rect 3023 35948 3036 36010
rect 3070 35948 3083 36010
rect 3023 35938 3083 35948
rect 3023 35880 3036 35938
rect 3070 35880 3083 35938
rect 3023 35866 3083 35880
rect 3023 35812 3036 35866
rect 3070 35812 3083 35866
rect 3023 35794 3083 35812
rect 3023 35744 3036 35794
rect 3070 35744 3083 35794
rect 3023 35722 3083 35744
rect 3023 35676 3036 35722
rect 3070 35676 3083 35722
rect 3023 35650 3083 35676
rect 3023 35608 3036 35650
rect 3070 35608 3083 35650
rect 3023 35578 3083 35608
rect 3023 35540 3036 35578
rect 3070 35540 3083 35578
rect 3023 35506 3083 35540
rect 3023 35472 3036 35506
rect 3070 35472 3083 35506
rect 3023 35438 3083 35472
rect 3023 35400 3036 35438
rect 3070 35400 3083 35438
rect 3023 35370 3083 35400
rect 3023 35328 3036 35370
rect 3070 35328 3083 35370
rect 3023 35302 3083 35328
rect 3023 35256 3036 35302
rect 3070 35256 3083 35302
rect 3023 35234 3083 35256
rect 3023 35184 3036 35234
rect 3070 35184 3083 35234
rect 3023 35166 3083 35184
rect 3023 35112 3036 35166
rect 3070 35112 3083 35166
rect 3023 35098 3083 35112
rect 3023 35040 3036 35098
rect 3070 35040 3083 35098
rect 3023 35030 3083 35040
rect 3023 34968 3036 35030
rect 3070 34968 3083 35030
rect 3023 34962 3083 34968
rect 3023 34896 3036 34962
rect 3070 34896 3083 34962
rect 3023 34894 3083 34896
rect 373 34839 433 34873
rect 373 34805 386 34839
rect 420 34805 433 34839
rect 373 34771 433 34805
rect 3023 34860 3036 34894
rect 3070 34860 3083 34894
rect 3023 34858 3083 34860
rect 373 34733 386 34771
rect 420 34733 433 34771
rect 576 34760 592 34794
rect 659 34760 662 34794
rect 696 34760 700 34794
rect 766 34760 775 34794
rect 836 34760 850 34794
rect 906 34760 925 34794
rect 976 34760 1000 34794
rect 1046 34760 1075 34794
rect 1116 34760 1150 34794
rect 1186 34760 1222 34794
rect 1259 34760 1292 34794
rect 1334 34760 1362 34794
rect 1409 34760 1432 34794
rect 1484 34760 1502 34794
rect 1559 34760 1572 34794
rect 1634 34760 1642 34794
rect 1708 34760 1712 34794
rect 1746 34760 1748 34794
rect 1816 34760 1822 34794
rect 1886 34760 1896 34794
rect 1956 34760 1970 34794
rect 2026 34760 2044 34794
rect 2096 34760 2118 34794
rect 2166 34760 2192 34794
rect 2236 34760 2266 34794
rect 2306 34760 2340 34794
rect 2376 34760 2412 34794
rect 2448 34760 2482 34794
rect 2522 34760 2552 34794
rect 2596 34760 2622 34794
rect 2670 34760 2692 34794
rect 2744 34760 2761 34794
rect 2818 34760 2830 34794
rect 2864 34760 2880 34794
rect 3023 34792 3036 34858
rect 3070 34792 3083 34858
rect 3023 34786 3083 34792
rect 373 34703 433 34733
rect 373 34661 386 34703
rect 420 34661 433 34703
rect 3023 34724 3036 34786
rect 3070 34724 3083 34786
rect 3023 34714 3083 34724
rect 373 34635 433 34661
rect 373 34589 386 34635
rect 420 34589 433 34635
rect 373 34567 433 34589
rect 373 34517 386 34567
rect 420 34517 433 34567
rect 373 34499 433 34517
rect 373 34445 386 34499
rect 420 34445 433 34499
rect 373 34431 433 34445
rect 373 34373 386 34431
rect 420 34373 433 34431
rect 373 34363 433 34373
rect 373 34301 386 34363
rect 420 34301 433 34363
rect 373 34295 433 34301
rect 373 34229 386 34295
rect 420 34229 433 34295
rect 373 34227 433 34229
rect 373 34193 386 34227
rect 420 34193 433 34227
rect 373 34191 433 34193
rect 373 34125 386 34191
rect 420 34125 433 34191
rect 373 34119 433 34125
rect 373 34057 386 34119
rect 420 34057 433 34119
rect 373 34047 433 34057
rect 373 33989 386 34047
rect 420 33989 433 34047
rect 373 33975 433 33989
rect 373 33921 386 33975
rect 420 33921 433 33975
rect 373 33903 433 33921
rect 373 33853 386 33903
rect 420 33853 433 33903
rect 373 33831 433 33853
rect 373 33785 386 33831
rect 420 33785 433 33831
rect 373 33759 433 33785
rect 373 33717 386 33759
rect 420 33717 433 33759
rect 373 33687 433 33717
rect 373 33649 386 33687
rect 420 33649 433 33687
rect 373 33615 433 33649
rect 373 33581 386 33615
rect 420 33581 433 33615
rect 373 33547 433 33581
rect 373 33509 386 33547
rect 420 33509 433 33547
rect 373 33479 433 33509
rect 373 33437 386 33479
rect 420 33437 433 33479
rect 373 33411 433 33437
rect 373 33365 386 33411
rect 420 33365 433 33411
rect 373 33343 433 33365
rect 373 33293 386 33343
rect 420 33293 433 33343
rect 373 33275 433 33293
rect 373 33221 386 33275
rect 420 33221 433 33275
rect 373 33207 433 33221
rect 373 33149 386 33207
rect 420 33149 433 33207
rect 373 33139 433 33149
rect 373 33077 386 33139
rect 420 33077 433 33139
rect 373 33071 433 33077
rect 373 33005 386 33071
rect 420 33005 433 33071
rect 373 33003 433 33005
rect 373 32969 386 33003
rect 420 32969 433 33003
rect 373 32967 433 32969
rect 373 32901 386 32967
rect 420 32901 433 32967
rect 373 32895 433 32901
rect 373 32833 386 32895
rect 420 32833 433 32895
rect 373 32823 433 32833
rect 373 32765 386 32823
rect 420 32765 433 32823
rect 373 32751 433 32765
rect 373 32697 386 32751
rect 420 32697 433 32751
rect 531 34619 565 34658
rect 531 34546 565 34585
rect 531 34473 565 34512
rect 531 34400 565 34439
rect 531 34327 565 34366
rect 531 34254 565 34293
rect 531 34181 565 34220
rect 531 34108 565 34147
rect 531 34035 565 34074
rect 531 33962 565 34001
rect 531 33889 565 33928
rect 531 33816 565 33855
rect 531 33742 565 33782
rect 531 33668 565 33708
rect 531 33594 565 33634
rect 531 33520 565 33560
rect 531 33446 565 33486
rect 531 33372 565 33412
rect 531 33298 565 33338
rect 531 33224 565 33264
rect 531 33150 565 33190
rect 531 33076 565 33116
rect 531 33002 565 33042
rect 531 32928 565 32968
rect 531 32854 565 32894
rect 531 32780 565 32820
rect 767 34619 801 34658
rect 767 34546 801 34585
rect 767 34473 801 34512
rect 767 34400 801 34439
rect 767 34327 801 34366
rect 767 34254 801 34293
rect 767 34181 801 34220
rect 767 34108 801 34147
rect 767 34035 801 34074
rect 767 33962 801 34001
rect 767 33889 801 33928
rect 767 33816 801 33855
rect 767 33742 801 33782
rect 767 33668 801 33708
rect 767 33594 801 33634
rect 767 33520 801 33560
rect 767 33446 801 33486
rect 767 33372 801 33412
rect 767 33298 801 33338
rect 767 33224 801 33264
rect 767 33150 801 33190
rect 767 33076 801 33116
rect 767 33002 801 33042
rect 767 32928 801 32968
rect 767 32854 801 32894
rect 767 32780 801 32820
rect 1003 34619 1037 34658
rect 1003 34546 1037 34585
rect 1003 34473 1037 34512
rect 1003 34400 1037 34439
rect 1003 34327 1037 34366
rect 1003 34254 1037 34293
rect 1003 34181 1037 34220
rect 1003 34108 1037 34147
rect 1003 34035 1037 34074
rect 1003 33962 1037 34001
rect 1003 33889 1037 33928
rect 1003 33816 1037 33855
rect 1003 33742 1037 33782
rect 1003 33668 1037 33708
rect 1003 33594 1037 33634
rect 1003 33520 1037 33560
rect 1003 33446 1037 33486
rect 1003 33372 1037 33412
rect 1003 33298 1037 33338
rect 1003 33224 1037 33264
rect 1003 33150 1037 33190
rect 1003 33076 1037 33116
rect 1003 33002 1037 33042
rect 1003 32928 1037 32968
rect 1003 32854 1037 32894
rect 1003 32780 1037 32820
rect 1239 34619 1273 34658
rect 1239 34546 1273 34585
rect 1239 34473 1273 34512
rect 1239 34400 1273 34439
rect 1239 34327 1273 34366
rect 1239 34254 1273 34293
rect 1239 34181 1273 34220
rect 1239 34108 1273 34147
rect 1239 34035 1273 34074
rect 1239 33962 1273 34001
rect 1239 33889 1273 33928
rect 1239 33816 1273 33855
rect 1239 33742 1273 33782
rect 1239 33668 1273 33708
rect 1239 33594 1273 33634
rect 1239 33520 1273 33560
rect 1239 33446 1273 33486
rect 1239 33372 1273 33412
rect 1239 33298 1273 33338
rect 1239 33224 1273 33264
rect 1239 33150 1273 33190
rect 1239 33076 1273 33116
rect 1239 33002 1273 33042
rect 1239 32928 1273 32968
rect 1239 32854 1273 32894
rect 1239 32780 1273 32820
rect 1475 34619 1509 34658
rect 1475 34546 1509 34585
rect 1475 34473 1509 34512
rect 1475 34400 1509 34439
rect 1475 34327 1509 34366
rect 1475 34254 1509 34293
rect 1475 34181 1509 34220
rect 1475 34108 1509 34147
rect 1475 34035 1509 34074
rect 1475 33962 1509 34001
rect 1475 33889 1509 33928
rect 1475 33816 1509 33855
rect 1475 33742 1509 33782
rect 1475 33668 1509 33708
rect 1475 33594 1509 33634
rect 1475 33520 1509 33560
rect 1475 33446 1509 33486
rect 1475 33372 1509 33412
rect 1475 33298 1509 33338
rect 1475 33224 1509 33264
rect 1475 33150 1509 33190
rect 1475 33076 1509 33116
rect 1475 33002 1509 33042
rect 1475 32928 1509 32968
rect 1475 32854 1509 32894
rect 1475 32780 1509 32820
rect 1711 34619 1745 34658
rect 1711 34546 1745 34585
rect 1711 34473 1745 34512
rect 1711 34400 1745 34439
rect 1711 34327 1745 34366
rect 1711 34254 1745 34293
rect 1711 34181 1745 34220
rect 1711 34108 1745 34147
rect 1711 34035 1745 34074
rect 1711 33962 1745 34001
rect 1711 33889 1745 33928
rect 1711 33816 1745 33855
rect 1711 33742 1745 33782
rect 1711 33668 1745 33708
rect 1711 33594 1745 33634
rect 1711 33520 1745 33560
rect 1711 33446 1745 33486
rect 1711 33372 1745 33412
rect 1711 33298 1745 33338
rect 1711 33224 1745 33264
rect 1711 33150 1745 33190
rect 1711 33076 1745 33116
rect 1711 33002 1745 33042
rect 1711 32928 1745 32968
rect 1711 32854 1745 32894
rect 1711 32780 1745 32820
rect 1947 34619 1981 34658
rect 1947 34546 1981 34585
rect 1947 34473 1981 34512
rect 1947 34400 1981 34439
rect 1947 34327 1981 34366
rect 1947 34254 1981 34293
rect 1947 34181 1981 34220
rect 1947 34108 1981 34147
rect 1947 34035 1981 34074
rect 1947 33962 1981 34001
rect 1947 33889 1981 33928
rect 1947 33816 1981 33855
rect 1947 33742 1981 33782
rect 1947 33668 1981 33708
rect 1947 33594 1981 33634
rect 1947 33520 1981 33560
rect 1947 33446 1981 33486
rect 1947 33372 1981 33412
rect 1947 33298 1981 33338
rect 1947 33224 1981 33264
rect 1947 33150 1981 33190
rect 1947 33076 1981 33116
rect 1947 33002 1981 33042
rect 1947 32928 1981 32968
rect 1947 32854 1981 32894
rect 1947 32780 1981 32820
rect 2183 34619 2217 34658
rect 2183 34546 2217 34585
rect 2183 34473 2217 34512
rect 2183 34400 2217 34439
rect 2183 34327 2217 34366
rect 2183 34254 2217 34293
rect 2183 34181 2217 34220
rect 2183 34108 2217 34147
rect 2183 34035 2217 34074
rect 2183 33962 2217 34001
rect 2183 33889 2217 33928
rect 2183 33816 2217 33855
rect 2183 33742 2217 33782
rect 2183 33668 2217 33708
rect 2183 33594 2217 33634
rect 2183 33520 2217 33560
rect 2183 33446 2217 33486
rect 2183 33372 2217 33412
rect 2183 33298 2217 33338
rect 2183 33224 2217 33264
rect 2183 33150 2217 33190
rect 2183 33076 2217 33116
rect 2183 33002 2217 33042
rect 2183 32928 2217 32968
rect 2183 32854 2217 32894
rect 2183 32780 2217 32820
rect 2419 34619 2453 34658
rect 2419 34546 2453 34585
rect 2419 34473 2453 34512
rect 2419 34400 2453 34439
rect 2419 34327 2453 34366
rect 2419 34254 2453 34293
rect 2419 34181 2453 34220
rect 2419 34108 2453 34147
rect 2419 34035 2453 34074
rect 2419 33962 2453 34001
rect 2419 33889 2453 33928
rect 2419 33816 2453 33855
rect 2419 33742 2453 33782
rect 2419 33668 2453 33708
rect 2419 33594 2453 33634
rect 2419 33520 2453 33560
rect 2419 33446 2453 33486
rect 2419 33372 2453 33412
rect 2419 33298 2453 33338
rect 2419 33224 2453 33264
rect 2419 33150 2453 33190
rect 2419 33076 2453 33116
rect 2419 33002 2453 33042
rect 2419 32928 2453 32968
rect 2419 32854 2453 32894
rect 2419 32780 2453 32820
rect 2655 34619 2689 34658
rect 2655 34546 2689 34585
rect 2655 34473 2689 34512
rect 2655 34400 2689 34439
rect 2655 34327 2689 34366
rect 2655 34254 2689 34293
rect 2655 34181 2689 34220
rect 2655 34108 2689 34147
rect 2655 34035 2689 34074
rect 2655 33962 2689 34001
rect 2655 33889 2689 33928
rect 2655 33816 2689 33855
rect 2655 33742 2689 33782
rect 2655 33668 2689 33708
rect 2655 33594 2689 33634
rect 2655 33520 2689 33560
rect 2655 33446 2689 33486
rect 2655 33372 2689 33412
rect 2655 33298 2689 33338
rect 2655 33224 2689 33264
rect 2655 33150 2689 33190
rect 2655 33076 2689 33116
rect 2655 33002 2689 33042
rect 2655 32928 2689 32968
rect 2655 32854 2689 32894
rect 2655 32780 2689 32820
rect 2891 34619 2925 34658
rect 2891 34546 2925 34585
rect 2891 34473 2925 34512
rect 2891 34400 2925 34439
rect 2891 34327 2925 34366
rect 2891 34254 2925 34293
rect 2891 34181 2925 34220
rect 2891 34108 2925 34147
rect 2891 34035 2925 34074
rect 2891 33962 2925 34001
rect 2891 33889 2925 33928
rect 2891 33816 2925 33855
rect 2891 33742 2925 33782
rect 2891 33668 2925 33708
rect 2891 33594 2925 33634
rect 2891 33520 2925 33560
rect 2891 33446 2925 33486
rect 2891 33372 2925 33412
rect 2891 33298 2925 33338
rect 2891 33224 2925 33264
rect 2891 33150 2925 33190
rect 2891 33076 2925 33116
rect 2891 33002 2925 33042
rect 2891 32928 2925 32968
rect 2891 32854 2925 32894
rect 2891 32780 2925 32820
rect 3023 34656 3036 34714
rect 3070 34656 3083 34714
rect 3023 34642 3083 34656
rect 3023 34588 3036 34642
rect 3070 34588 3083 34642
rect 3023 34570 3083 34588
rect 3023 34520 3036 34570
rect 3070 34520 3083 34570
rect 3023 34498 3083 34520
rect 3023 34452 3036 34498
rect 3070 34452 3083 34498
rect 3023 34426 3083 34452
rect 3023 34384 3036 34426
rect 3070 34384 3083 34426
rect 3023 34354 3083 34384
rect 3023 34316 3036 34354
rect 3070 34316 3083 34354
rect 3023 34282 3083 34316
rect 3023 34248 3036 34282
rect 3070 34248 3083 34282
rect 3023 34214 3083 34248
rect 3023 34176 3036 34214
rect 3070 34176 3083 34214
rect 3023 34146 3083 34176
rect 3023 34104 3036 34146
rect 3070 34104 3083 34146
rect 3023 34078 3083 34104
rect 3023 34032 3036 34078
rect 3070 34032 3083 34078
rect 3023 34010 3083 34032
rect 3023 33960 3036 34010
rect 3070 33960 3083 34010
rect 3023 33942 3083 33960
rect 3023 33888 3036 33942
rect 3070 33888 3083 33942
rect 3023 33874 3083 33888
rect 3023 33816 3036 33874
rect 3070 33816 3083 33874
rect 3023 33806 3083 33816
rect 3023 33744 3036 33806
rect 3070 33744 3083 33806
rect 3023 33738 3083 33744
rect 3023 33672 3036 33738
rect 3070 33672 3083 33738
rect 3023 33670 3083 33672
rect 3023 33636 3036 33670
rect 3070 33636 3083 33670
rect 3023 33634 3083 33636
rect 3023 33568 3036 33634
rect 3070 33568 3083 33634
rect 3023 33562 3083 33568
rect 3023 33500 3036 33562
rect 3070 33500 3083 33562
rect 3023 33490 3083 33500
rect 3023 33432 3036 33490
rect 3070 33432 3083 33490
rect 3023 33418 3083 33432
rect 3023 33364 3036 33418
rect 3070 33364 3083 33418
rect 3023 33346 3083 33364
rect 3023 33296 3036 33346
rect 3070 33296 3083 33346
rect 3023 33274 3083 33296
rect 3023 33228 3036 33274
rect 3070 33228 3083 33274
rect 3023 33202 3083 33228
rect 3023 33160 3036 33202
rect 3070 33160 3083 33202
rect 3023 33130 3083 33160
rect 3023 33092 3036 33130
rect 3070 33092 3083 33130
rect 3023 33058 3083 33092
rect 3023 33024 3036 33058
rect 3070 33024 3083 33058
rect 3023 32990 3083 33024
rect 3023 32952 3036 32990
rect 3070 32952 3083 32990
rect 3023 32922 3083 32952
rect 3023 32880 3036 32922
rect 3070 32880 3083 32922
rect 3023 32854 3083 32880
rect 3023 32808 3036 32854
rect 3070 32808 3083 32854
rect 3023 32786 3083 32808
rect 373 32679 433 32697
rect 373 32629 386 32679
rect 420 32629 433 32679
rect 3023 32736 3036 32786
rect 3070 32736 3083 32786
rect 3023 32718 3083 32736
rect 3023 32664 3036 32718
rect 3070 32664 3083 32718
rect 576 32630 592 32664
rect 659 32630 662 32664
rect 696 32630 700 32664
rect 766 32630 775 32664
rect 836 32630 850 32664
rect 906 32630 925 32664
rect 976 32630 1000 32664
rect 1046 32630 1075 32664
rect 1116 32630 1150 32664
rect 1186 32630 1222 32664
rect 1259 32630 1292 32664
rect 1334 32630 1362 32664
rect 1409 32630 1432 32664
rect 1484 32630 1502 32664
rect 1559 32630 1572 32664
rect 1634 32630 1642 32664
rect 1708 32630 1712 32664
rect 1746 32630 1748 32664
rect 1816 32630 1822 32664
rect 1886 32630 1896 32664
rect 1956 32630 1970 32664
rect 2026 32630 2044 32664
rect 2096 32630 2118 32664
rect 2166 32630 2192 32664
rect 2236 32630 2266 32664
rect 2306 32630 2340 32664
rect 2376 32630 2412 32664
rect 2448 32630 2482 32664
rect 2522 32630 2552 32664
rect 2596 32630 2622 32664
rect 2670 32630 2692 32664
rect 2744 32630 2761 32664
rect 2818 32630 2830 32664
rect 2864 32630 2880 32664
rect 3023 32650 3083 32664
rect 373 32607 433 32629
rect 373 32561 386 32607
rect 420 32561 433 32607
rect 373 32535 433 32561
rect 3023 32592 3036 32650
rect 3070 32592 3083 32650
rect 3023 32582 3083 32592
rect 373 32493 386 32535
rect 420 32493 433 32535
rect 373 32463 433 32493
rect 373 32425 386 32463
rect 420 32425 433 32463
rect 373 32391 433 32425
rect 373 32357 386 32391
rect 420 32357 433 32391
rect 373 32323 433 32357
rect 373 32285 386 32323
rect 420 32285 433 32323
rect 373 32255 433 32285
rect 373 32213 386 32255
rect 420 32213 433 32255
rect 373 32187 433 32213
rect 373 32141 386 32187
rect 420 32141 433 32187
rect 373 32119 433 32141
rect 373 32069 386 32119
rect 420 32069 433 32119
rect 373 32051 433 32069
rect 373 31997 386 32051
rect 420 31997 433 32051
rect 373 31983 433 31997
rect 373 31925 386 31983
rect 420 31925 433 31983
rect 373 31915 433 31925
rect 373 31853 386 31915
rect 420 31853 433 31915
rect 373 31847 433 31853
rect 373 31781 386 31847
rect 420 31781 433 31847
rect 373 31779 433 31781
rect 373 31745 386 31779
rect 420 31745 433 31779
rect 373 31743 433 31745
rect 373 31677 386 31743
rect 420 31677 433 31743
rect 373 31671 433 31677
rect 373 31609 386 31671
rect 420 31609 433 31671
rect 373 31599 433 31609
rect 373 31541 386 31599
rect 420 31541 433 31599
rect 373 31527 433 31541
rect 373 31473 386 31527
rect 420 31473 433 31527
rect 373 31455 433 31473
rect 373 31405 386 31455
rect 420 31405 433 31455
rect 373 31383 433 31405
rect 373 31337 386 31383
rect 420 31337 433 31383
rect 373 31311 433 31337
rect 373 31269 386 31311
rect 420 31269 433 31311
rect 373 31239 433 31269
rect 373 31201 386 31239
rect 420 31201 433 31239
rect 373 31167 433 31201
rect 373 31133 386 31167
rect 420 31133 433 31167
rect 373 31099 433 31133
rect 373 31061 386 31099
rect 420 31061 433 31099
rect 373 31031 433 31061
rect 373 30989 386 31031
rect 420 30989 433 31031
rect 373 30963 433 30989
rect 373 30917 386 30963
rect 420 30917 433 30963
rect 373 30895 433 30917
rect 373 30845 386 30895
rect 420 30845 433 30895
rect 373 30827 433 30845
rect 373 30773 386 30827
rect 420 30773 433 30827
rect 373 30759 433 30773
rect 373 30701 386 30759
rect 420 30701 433 30759
rect 373 30691 433 30701
rect 373 30629 386 30691
rect 420 30629 433 30691
rect 373 30623 433 30629
rect 373 30557 386 30623
rect 420 30557 433 30623
rect 531 32475 565 32514
rect 531 32402 565 32441
rect 531 32329 565 32368
rect 531 32256 565 32295
rect 531 32183 565 32222
rect 531 32110 565 32149
rect 531 32037 565 32076
rect 531 31964 565 32003
rect 531 31891 565 31930
rect 531 31818 565 31857
rect 531 31745 565 31784
rect 531 31672 565 31711
rect 531 31598 565 31638
rect 531 31524 565 31564
rect 531 31450 565 31490
rect 531 31376 565 31416
rect 531 31302 565 31342
rect 531 31228 565 31268
rect 531 31154 565 31194
rect 531 31080 565 31120
rect 531 31006 565 31046
rect 531 30932 565 30972
rect 531 30858 565 30898
rect 531 30784 565 30824
rect 531 30710 565 30750
rect 531 30636 565 30676
rect 767 32475 801 32514
rect 767 32402 801 32441
rect 767 32329 801 32368
rect 767 32256 801 32295
rect 767 32183 801 32222
rect 767 32110 801 32149
rect 767 32037 801 32076
rect 767 31964 801 32003
rect 767 31891 801 31930
rect 767 31818 801 31857
rect 767 31745 801 31784
rect 767 31672 801 31711
rect 767 31598 801 31638
rect 767 31524 801 31564
rect 767 31450 801 31490
rect 767 31376 801 31416
rect 767 31302 801 31342
rect 767 31228 801 31268
rect 767 31154 801 31194
rect 767 31080 801 31120
rect 767 31006 801 31046
rect 767 30932 801 30972
rect 767 30858 801 30898
rect 767 30784 801 30824
rect 767 30710 801 30750
rect 767 30636 801 30676
rect 1003 32475 1037 32514
rect 1003 32402 1037 32441
rect 1003 32329 1037 32368
rect 1003 32256 1037 32295
rect 1003 32183 1037 32222
rect 1003 32110 1037 32149
rect 1003 32037 1037 32076
rect 1003 31964 1037 32003
rect 1003 31891 1037 31930
rect 1003 31818 1037 31857
rect 1003 31745 1037 31784
rect 1003 31672 1037 31711
rect 1003 31598 1037 31638
rect 1003 31524 1037 31564
rect 1003 31450 1037 31490
rect 1003 31376 1037 31416
rect 1003 31302 1037 31342
rect 1003 31228 1037 31268
rect 1003 31154 1037 31194
rect 1003 31080 1037 31120
rect 1003 31006 1037 31046
rect 1003 30932 1037 30972
rect 1003 30858 1037 30898
rect 1003 30784 1037 30824
rect 1003 30710 1037 30750
rect 1003 30636 1037 30676
rect 1239 32475 1273 32514
rect 1239 32402 1273 32441
rect 1239 32329 1273 32368
rect 1239 32256 1273 32295
rect 1239 32183 1273 32222
rect 1239 32110 1273 32149
rect 1239 32037 1273 32076
rect 1239 31964 1273 32003
rect 1239 31891 1273 31930
rect 1239 31818 1273 31857
rect 1239 31745 1273 31784
rect 1239 31672 1273 31711
rect 1239 31598 1273 31638
rect 1239 31524 1273 31564
rect 1239 31450 1273 31490
rect 1239 31376 1273 31416
rect 1239 31302 1273 31342
rect 1239 31228 1273 31268
rect 1239 31154 1273 31194
rect 1239 31080 1273 31120
rect 1239 31006 1273 31046
rect 1239 30932 1273 30972
rect 1239 30858 1273 30898
rect 1239 30784 1273 30824
rect 1239 30710 1273 30750
rect 1239 30636 1273 30676
rect 1475 32475 1509 32514
rect 1475 32402 1509 32441
rect 1475 32329 1509 32368
rect 1475 32256 1509 32295
rect 1475 32183 1509 32222
rect 1475 32110 1509 32149
rect 1475 32037 1509 32076
rect 1475 31964 1509 32003
rect 1475 31891 1509 31930
rect 1475 31818 1509 31857
rect 1475 31745 1509 31784
rect 1475 31672 1509 31711
rect 1475 31598 1509 31638
rect 1475 31524 1509 31564
rect 1475 31450 1509 31490
rect 1475 31376 1509 31416
rect 1475 31302 1509 31342
rect 1475 31228 1509 31268
rect 1475 31154 1509 31194
rect 1475 31080 1509 31120
rect 1475 31006 1509 31046
rect 1475 30932 1509 30972
rect 1475 30858 1509 30898
rect 1475 30784 1509 30824
rect 1475 30710 1509 30750
rect 1475 30636 1509 30676
rect 1711 32475 1745 32514
rect 1711 32402 1745 32441
rect 1711 32329 1745 32368
rect 1711 32256 1745 32295
rect 1711 32183 1745 32222
rect 1711 32110 1745 32149
rect 1711 32037 1745 32076
rect 1711 31964 1745 32003
rect 1711 31891 1745 31930
rect 1711 31818 1745 31857
rect 1711 31745 1745 31784
rect 1711 31672 1745 31711
rect 1711 31598 1745 31638
rect 1711 31524 1745 31564
rect 1711 31450 1745 31490
rect 1711 31376 1745 31416
rect 1711 31302 1745 31342
rect 1711 31228 1745 31268
rect 1711 31154 1745 31194
rect 1711 31080 1745 31120
rect 1711 31006 1745 31046
rect 1711 30932 1745 30972
rect 1711 30858 1745 30898
rect 1711 30784 1745 30824
rect 1711 30710 1745 30750
rect 1711 30636 1745 30676
rect 1947 32475 1981 32514
rect 1947 32402 1981 32441
rect 1947 32329 1981 32368
rect 1947 32256 1981 32295
rect 1947 32183 1981 32222
rect 1947 32110 1981 32149
rect 1947 32037 1981 32076
rect 1947 31964 1981 32003
rect 1947 31891 1981 31930
rect 1947 31818 1981 31857
rect 1947 31745 1981 31784
rect 1947 31672 1981 31711
rect 1947 31598 1981 31638
rect 1947 31524 1981 31564
rect 1947 31450 1981 31490
rect 1947 31376 1981 31416
rect 1947 31302 1981 31342
rect 1947 31228 1981 31268
rect 1947 31154 1981 31194
rect 1947 31080 1981 31120
rect 1947 31006 1981 31046
rect 1947 30932 1981 30972
rect 1947 30858 1981 30898
rect 1947 30784 1981 30824
rect 1947 30710 1981 30750
rect 1947 30636 1981 30676
rect 2183 32475 2217 32514
rect 2183 32402 2217 32441
rect 2183 32329 2217 32368
rect 2183 32256 2217 32295
rect 2183 32183 2217 32222
rect 2183 32110 2217 32149
rect 2183 32037 2217 32076
rect 2183 31964 2217 32003
rect 2183 31891 2217 31930
rect 2183 31818 2217 31857
rect 2183 31745 2217 31784
rect 2183 31672 2217 31711
rect 2183 31598 2217 31638
rect 2183 31524 2217 31564
rect 2183 31450 2217 31490
rect 2183 31376 2217 31416
rect 2183 31302 2217 31342
rect 2183 31228 2217 31268
rect 2183 31154 2217 31194
rect 2183 31080 2217 31120
rect 2183 31006 2217 31046
rect 2183 30932 2217 30972
rect 2183 30858 2217 30898
rect 2183 30784 2217 30824
rect 2183 30710 2217 30750
rect 2183 30636 2217 30676
rect 2419 32475 2453 32514
rect 2419 32402 2453 32441
rect 2419 32329 2453 32368
rect 2419 32256 2453 32295
rect 2419 32183 2453 32222
rect 2419 32110 2453 32149
rect 2419 32037 2453 32076
rect 2419 31964 2453 32003
rect 2419 31891 2453 31930
rect 2419 31818 2453 31857
rect 2419 31745 2453 31784
rect 2419 31672 2453 31711
rect 2419 31598 2453 31638
rect 2419 31524 2453 31564
rect 2419 31450 2453 31490
rect 2419 31376 2453 31416
rect 2419 31302 2453 31342
rect 2419 31228 2453 31268
rect 2419 31154 2453 31194
rect 2419 31080 2453 31120
rect 2419 31006 2453 31046
rect 2419 30932 2453 30972
rect 2419 30858 2453 30898
rect 2419 30784 2453 30824
rect 2419 30710 2453 30750
rect 2419 30636 2453 30676
rect 2655 32475 2689 32514
rect 2655 32402 2689 32441
rect 2655 32329 2689 32368
rect 2655 32256 2689 32295
rect 2655 32183 2689 32222
rect 2655 32110 2689 32149
rect 2655 32037 2689 32076
rect 2655 31964 2689 32003
rect 2655 31891 2689 31930
rect 2655 31818 2689 31857
rect 2655 31745 2689 31784
rect 2655 31672 2689 31711
rect 2655 31598 2689 31638
rect 2655 31524 2689 31564
rect 2655 31450 2689 31490
rect 2655 31376 2689 31416
rect 2655 31302 2689 31342
rect 2655 31228 2689 31268
rect 2655 31154 2689 31194
rect 2655 31080 2689 31120
rect 2655 31006 2689 31046
rect 2655 30932 2689 30972
rect 2655 30858 2689 30898
rect 2655 30784 2689 30824
rect 2655 30710 2689 30750
rect 2655 30636 2689 30676
rect 2891 32475 2925 32514
rect 2891 32402 2925 32441
rect 2891 32329 2925 32368
rect 2891 32256 2925 32295
rect 2891 32183 2925 32222
rect 2891 32110 2925 32149
rect 2891 32037 2925 32076
rect 2891 31964 2925 32003
rect 2891 31891 2925 31930
rect 2891 31818 2925 31857
rect 2891 31745 2925 31784
rect 2891 31672 2925 31711
rect 2891 31598 2925 31638
rect 2891 31524 2925 31564
rect 2891 31450 2925 31490
rect 2891 31376 2925 31416
rect 2891 31302 2925 31342
rect 2891 31228 2925 31268
rect 2891 31154 2925 31194
rect 2891 31080 2925 31120
rect 2891 31006 2925 31046
rect 2891 30932 2925 30972
rect 2891 30858 2925 30898
rect 2891 30784 2925 30824
rect 2891 30710 2925 30750
rect 2891 30636 2925 30676
rect 3023 32520 3036 32582
rect 3070 32520 3083 32582
rect 3023 32514 3083 32520
rect 3023 32448 3036 32514
rect 3070 32448 3083 32514
rect 3023 32446 3083 32448
rect 3023 32412 3036 32446
rect 3070 32412 3083 32446
rect 3023 32410 3083 32412
rect 3023 32344 3036 32410
rect 3070 32344 3083 32410
rect 3023 32338 3083 32344
rect 3023 32276 3036 32338
rect 3070 32276 3083 32338
rect 3023 32266 3083 32276
rect 3023 32208 3036 32266
rect 3070 32208 3083 32266
rect 3023 32194 3083 32208
rect 3023 32140 3036 32194
rect 3070 32140 3083 32194
rect 3023 32122 3083 32140
rect 3023 32072 3036 32122
rect 3070 32072 3083 32122
rect 3023 32050 3083 32072
rect 3023 32004 3036 32050
rect 3070 32004 3083 32050
rect 3023 31978 3083 32004
rect 3023 31936 3036 31978
rect 3070 31936 3083 31978
rect 3023 31906 3083 31936
rect 3023 31868 3036 31906
rect 3070 31868 3083 31906
rect 3023 31834 3083 31868
rect 3023 31800 3036 31834
rect 3070 31800 3083 31834
rect 3023 31766 3083 31800
rect 3023 31728 3036 31766
rect 3070 31728 3083 31766
rect 3023 31698 3083 31728
rect 3023 31656 3036 31698
rect 3070 31656 3083 31698
rect 3023 31630 3083 31656
rect 3023 31584 3036 31630
rect 3070 31584 3083 31630
rect 3023 31562 3083 31584
rect 3023 31512 3036 31562
rect 3070 31512 3083 31562
rect 3023 31494 3083 31512
rect 3023 31440 3036 31494
rect 3070 31440 3083 31494
rect 3023 31426 3083 31440
rect 3023 31368 3036 31426
rect 3070 31368 3083 31426
rect 3023 31358 3083 31368
rect 3023 31296 3036 31358
rect 3070 31296 3083 31358
rect 3023 31290 3083 31296
rect 3023 31224 3036 31290
rect 3070 31224 3083 31290
rect 3023 31222 3083 31224
rect 3023 31188 3036 31222
rect 3070 31188 3083 31222
rect 3023 31186 3083 31188
rect 3023 31120 3036 31186
rect 3070 31120 3083 31186
rect 3023 31114 3083 31120
rect 3023 31052 3036 31114
rect 3070 31052 3083 31114
rect 3023 31042 3083 31052
rect 3023 30984 3036 31042
rect 3070 30984 3083 31042
rect 3023 30970 3083 30984
rect 3023 30916 3036 30970
rect 3070 30916 3083 30970
rect 3023 30898 3083 30916
rect 3023 30848 3036 30898
rect 3070 30848 3083 30898
rect 3023 30826 3083 30848
rect 3023 30780 3036 30826
rect 3070 30780 3083 30826
rect 3023 30754 3083 30780
rect 3023 30712 3036 30754
rect 3070 30712 3083 30754
rect 3023 30682 3083 30712
rect 3023 30644 3036 30682
rect 3070 30644 3083 30682
rect 3023 30610 3083 30644
rect 373 30555 433 30557
rect 373 30521 386 30555
rect 420 30521 433 30555
rect 3023 30576 3036 30610
rect 3070 30576 3083 30610
rect 3023 30542 3083 30576
rect 373 30519 433 30521
rect 373 30453 386 30519
rect 420 30453 433 30519
rect 576 30500 592 30534
rect 659 30500 662 30534
rect 696 30500 700 30534
rect 766 30500 775 30534
rect 836 30500 850 30534
rect 906 30500 925 30534
rect 976 30500 1000 30534
rect 1046 30500 1075 30534
rect 1116 30500 1150 30534
rect 1186 30500 1222 30534
rect 1259 30500 1292 30534
rect 1334 30500 1362 30534
rect 1409 30500 1432 30534
rect 1484 30500 1502 30534
rect 1559 30500 1572 30534
rect 1634 30500 1642 30534
rect 1708 30500 1712 30534
rect 1746 30500 1748 30534
rect 1816 30500 1822 30534
rect 1886 30500 1896 30534
rect 1956 30500 1970 30534
rect 2026 30500 2044 30534
rect 2096 30500 2118 30534
rect 2166 30500 2192 30534
rect 2236 30500 2266 30534
rect 2306 30500 2340 30534
rect 2376 30500 2412 30534
rect 2448 30500 2482 30534
rect 2522 30500 2552 30534
rect 2596 30500 2622 30534
rect 2670 30500 2692 30534
rect 2744 30500 2761 30534
rect 2818 30500 2830 30534
rect 2864 30500 2880 30534
rect 3023 30504 3036 30542
rect 3070 30504 3083 30542
rect 373 30447 433 30453
rect 373 30385 386 30447
rect 420 30385 433 30447
rect 3023 30474 3083 30504
rect 3023 30432 3036 30474
rect 3070 30432 3083 30474
rect 373 30375 433 30385
rect 373 30317 386 30375
rect 420 30317 433 30375
rect 373 30303 433 30317
rect 373 30249 386 30303
rect 420 30249 433 30303
rect 373 30231 433 30249
rect 373 30181 386 30231
rect 420 30181 433 30231
rect 373 30159 433 30181
rect 373 30113 386 30159
rect 420 30113 433 30159
rect 373 30087 433 30113
rect 373 30045 386 30087
rect 420 30045 433 30087
rect 373 30015 433 30045
rect 373 29977 386 30015
rect 420 29977 433 30015
rect 373 29943 433 29977
rect 373 29909 386 29943
rect 420 29909 433 29943
rect 373 29875 433 29909
rect 373 29837 386 29875
rect 420 29837 433 29875
rect 373 29807 433 29837
rect 373 29765 386 29807
rect 420 29765 433 29807
rect 373 29739 433 29765
rect 373 29693 386 29739
rect 420 29693 433 29739
rect 373 29671 433 29693
rect 373 29621 386 29671
rect 420 29621 433 29671
rect 373 29603 433 29621
rect 373 29549 386 29603
rect 420 29549 433 29603
rect 373 29535 433 29549
rect 373 29477 386 29535
rect 420 29477 433 29535
rect 373 29467 433 29477
rect 373 29405 386 29467
rect 420 29405 433 29467
rect 373 29399 433 29405
rect 373 29333 386 29399
rect 420 29333 433 29399
rect 373 29331 433 29333
rect 373 29297 386 29331
rect 420 29297 433 29331
rect 373 29295 433 29297
rect 373 29229 386 29295
rect 420 29229 433 29295
rect 373 29223 433 29229
rect 373 29161 386 29223
rect 420 29161 433 29223
rect 373 29151 433 29161
rect 373 29093 386 29151
rect 420 29093 433 29151
rect 373 29079 433 29093
rect 373 29025 386 29079
rect 420 29025 433 29079
rect 373 29007 433 29025
rect 373 28957 386 29007
rect 420 28957 433 29007
rect 373 28935 433 28957
rect 373 28889 386 28935
rect 420 28889 433 28935
rect 373 28863 433 28889
rect 373 28821 386 28863
rect 420 28821 433 28863
rect 373 28791 433 28821
rect 373 28753 386 28791
rect 420 28753 433 28791
rect 373 28719 433 28753
rect 373 28685 386 28719
rect 420 28685 433 28719
rect 373 28651 433 28685
rect 373 28613 386 28651
rect 420 28613 433 28651
rect 373 28583 433 28613
rect 373 28541 386 28583
rect 420 28541 433 28583
rect 373 28515 433 28541
rect 373 28469 386 28515
rect 420 28469 433 28515
rect 531 30359 565 30398
rect 531 30286 565 30325
rect 531 30213 565 30252
rect 531 30140 565 30179
rect 531 30067 565 30106
rect 531 29994 565 30033
rect 531 29921 565 29960
rect 531 29848 565 29887
rect 531 29775 565 29814
rect 531 29702 565 29741
rect 531 29629 565 29668
rect 531 29556 565 29595
rect 531 29482 565 29522
rect 531 29408 565 29448
rect 531 29334 565 29374
rect 531 29260 565 29300
rect 531 29186 565 29226
rect 531 29112 565 29152
rect 531 29038 565 29078
rect 531 28964 565 29004
rect 531 28890 565 28930
rect 531 28816 565 28856
rect 531 28742 565 28782
rect 531 28668 565 28708
rect 531 28594 565 28634
rect 531 28520 565 28560
rect 767 30359 801 30398
rect 767 30286 801 30325
rect 767 30213 801 30252
rect 767 30140 801 30179
rect 767 30067 801 30106
rect 767 29994 801 30033
rect 767 29921 801 29960
rect 767 29848 801 29887
rect 767 29775 801 29814
rect 767 29702 801 29741
rect 767 29629 801 29668
rect 767 29556 801 29595
rect 767 29482 801 29522
rect 767 29408 801 29448
rect 767 29334 801 29374
rect 767 29260 801 29300
rect 767 29186 801 29226
rect 767 29112 801 29152
rect 767 29038 801 29078
rect 767 28964 801 29004
rect 767 28890 801 28930
rect 767 28816 801 28856
rect 767 28742 801 28782
rect 767 28668 801 28708
rect 767 28594 801 28634
rect 767 28520 801 28560
rect 1003 30359 1037 30398
rect 1003 30286 1037 30325
rect 1003 30213 1037 30252
rect 1003 30140 1037 30179
rect 1003 30067 1037 30106
rect 1003 29994 1037 30033
rect 1003 29921 1037 29960
rect 1003 29848 1037 29887
rect 1003 29775 1037 29814
rect 1003 29702 1037 29741
rect 1003 29629 1037 29668
rect 1003 29556 1037 29595
rect 1003 29482 1037 29522
rect 1003 29408 1037 29448
rect 1003 29334 1037 29374
rect 1003 29260 1037 29300
rect 1003 29186 1037 29226
rect 1003 29112 1037 29152
rect 1003 29038 1037 29078
rect 1003 28964 1037 29004
rect 1003 28890 1037 28930
rect 1003 28816 1037 28856
rect 1003 28742 1037 28782
rect 1003 28668 1037 28708
rect 1003 28594 1037 28634
rect 1003 28520 1037 28560
rect 1239 30359 1273 30398
rect 1239 30286 1273 30325
rect 1239 30213 1273 30252
rect 1239 30140 1273 30179
rect 1239 30067 1273 30106
rect 1239 29994 1273 30033
rect 1239 29921 1273 29960
rect 1239 29848 1273 29887
rect 1239 29775 1273 29814
rect 1239 29702 1273 29741
rect 1239 29629 1273 29668
rect 1239 29556 1273 29595
rect 1239 29482 1273 29522
rect 1239 29408 1273 29448
rect 1239 29334 1273 29374
rect 1239 29260 1273 29300
rect 1239 29186 1273 29226
rect 1239 29112 1273 29152
rect 1239 29038 1273 29078
rect 1239 28964 1273 29004
rect 1239 28890 1273 28930
rect 1239 28816 1273 28856
rect 1239 28742 1273 28782
rect 1239 28668 1273 28708
rect 1239 28594 1273 28634
rect 1239 28520 1273 28560
rect 1475 30359 1509 30398
rect 1475 30286 1509 30325
rect 1475 30213 1509 30252
rect 1475 30140 1509 30179
rect 1475 30067 1509 30106
rect 1475 29994 1509 30033
rect 1475 29921 1509 29960
rect 1475 29848 1509 29887
rect 1475 29775 1509 29814
rect 1475 29702 1509 29741
rect 1475 29629 1509 29668
rect 1475 29556 1509 29595
rect 1475 29482 1509 29522
rect 1475 29408 1509 29448
rect 1475 29334 1509 29374
rect 1475 29260 1509 29300
rect 1475 29186 1509 29226
rect 1475 29112 1509 29152
rect 1475 29038 1509 29078
rect 1475 28964 1509 29004
rect 1475 28890 1509 28930
rect 1475 28816 1509 28856
rect 1475 28742 1509 28782
rect 1475 28668 1509 28708
rect 1475 28594 1509 28634
rect 1475 28520 1509 28560
rect 1711 30359 1745 30398
rect 1711 30286 1745 30325
rect 1711 30213 1745 30252
rect 1711 30140 1745 30179
rect 1711 30067 1745 30106
rect 1711 29994 1745 30033
rect 1711 29921 1745 29960
rect 1711 29848 1745 29887
rect 1711 29775 1745 29814
rect 1711 29702 1745 29741
rect 1711 29629 1745 29668
rect 1711 29556 1745 29595
rect 1711 29482 1745 29522
rect 1711 29408 1745 29448
rect 1711 29334 1745 29374
rect 1711 29260 1745 29300
rect 1711 29186 1745 29226
rect 1711 29112 1745 29152
rect 1711 29038 1745 29078
rect 1711 28964 1745 29004
rect 1711 28890 1745 28930
rect 1711 28816 1745 28856
rect 1711 28742 1745 28782
rect 1711 28668 1745 28708
rect 1711 28594 1745 28634
rect 1711 28520 1745 28560
rect 1947 30359 1981 30398
rect 1947 30286 1981 30325
rect 1947 30213 1981 30252
rect 1947 30140 1981 30179
rect 1947 30067 1981 30106
rect 1947 29994 1981 30033
rect 1947 29921 1981 29960
rect 1947 29848 1981 29887
rect 1947 29775 1981 29814
rect 1947 29702 1981 29741
rect 1947 29629 1981 29668
rect 1947 29556 1981 29595
rect 1947 29482 1981 29522
rect 1947 29408 1981 29448
rect 1947 29334 1981 29374
rect 1947 29260 1981 29300
rect 1947 29186 1981 29226
rect 1947 29112 1981 29152
rect 1947 29038 1981 29078
rect 1947 28964 1981 29004
rect 1947 28890 1981 28930
rect 1947 28816 1981 28856
rect 1947 28742 1981 28782
rect 1947 28668 1981 28708
rect 1947 28594 1981 28634
rect 1947 28520 1981 28560
rect 2183 30359 2217 30398
rect 2183 30286 2217 30325
rect 2183 30213 2217 30252
rect 2183 30140 2217 30179
rect 2183 30067 2217 30106
rect 2183 29994 2217 30033
rect 2183 29921 2217 29960
rect 2183 29848 2217 29887
rect 2183 29775 2217 29814
rect 2183 29702 2217 29741
rect 2183 29629 2217 29668
rect 2183 29556 2217 29595
rect 2183 29482 2217 29522
rect 2183 29408 2217 29448
rect 2183 29334 2217 29374
rect 2183 29260 2217 29300
rect 2183 29186 2217 29226
rect 2183 29112 2217 29152
rect 2183 29038 2217 29078
rect 2183 28964 2217 29004
rect 2183 28890 2217 28930
rect 2183 28816 2217 28856
rect 2183 28742 2217 28782
rect 2183 28668 2217 28708
rect 2183 28594 2217 28634
rect 2183 28520 2217 28560
rect 2419 30359 2453 30398
rect 2419 30286 2453 30325
rect 2419 30213 2453 30252
rect 2419 30140 2453 30179
rect 2419 30067 2453 30106
rect 2419 29994 2453 30033
rect 2419 29921 2453 29960
rect 2419 29848 2453 29887
rect 2419 29775 2453 29814
rect 2419 29702 2453 29741
rect 2419 29629 2453 29668
rect 2419 29556 2453 29595
rect 2419 29482 2453 29522
rect 2419 29408 2453 29448
rect 2419 29334 2453 29374
rect 2419 29260 2453 29300
rect 2419 29186 2453 29226
rect 2419 29112 2453 29152
rect 2419 29038 2453 29078
rect 2419 28964 2453 29004
rect 2419 28890 2453 28930
rect 2419 28816 2453 28856
rect 2419 28742 2453 28782
rect 2419 28668 2453 28708
rect 2419 28594 2453 28634
rect 2419 28520 2453 28560
rect 2655 30359 2689 30398
rect 2655 30286 2689 30325
rect 2655 30213 2689 30252
rect 2655 30140 2689 30179
rect 2655 30067 2689 30106
rect 2655 29994 2689 30033
rect 2655 29921 2689 29960
rect 2655 29848 2689 29887
rect 2655 29775 2689 29814
rect 2655 29702 2689 29741
rect 2655 29629 2689 29668
rect 2655 29556 2689 29595
rect 2655 29482 2689 29522
rect 2655 29408 2689 29448
rect 2655 29334 2689 29374
rect 2655 29260 2689 29300
rect 2655 29186 2689 29226
rect 2655 29112 2689 29152
rect 2655 29038 2689 29078
rect 2655 28964 2689 29004
rect 2655 28890 2689 28930
rect 2655 28816 2689 28856
rect 2655 28742 2689 28782
rect 2655 28668 2689 28708
rect 2655 28594 2689 28634
rect 2655 28520 2689 28560
rect 2891 30359 2925 30398
rect 2891 30286 2925 30325
rect 2891 30213 2925 30252
rect 2891 30140 2925 30179
rect 2891 30067 2925 30106
rect 2891 29994 2925 30033
rect 2891 29921 2925 29960
rect 2891 29848 2925 29887
rect 2891 29775 2925 29814
rect 2891 29702 2925 29741
rect 2891 29629 2925 29668
rect 2891 29556 2925 29595
rect 2891 29482 2925 29522
rect 2891 29408 2925 29448
rect 2891 29334 2925 29374
rect 2891 29260 2925 29300
rect 2891 29186 2925 29226
rect 2891 29112 2925 29152
rect 2891 29038 2925 29078
rect 2891 28964 2925 29004
rect 2891 28890 2925 28930
rect 2891 28816 2925 28856
rect 2891 28742 2925 28782
rect 2891 28668 2925 28708
rect 2891 28594 2925 28634
rect 2891 28520 2925 28560
rect 3023 30406 3083 30432
rect 3023 30360 3036 30406
rect 3070 30360 3083 30406
rect 3023 30338 3083 30360
rect 3023 30288 3036 30338
rect 3070 30288 3083 30338
rect 3023 30270 3083 30288
rect 3023 30216 3036 30270
rect 3070 30216 3083 30270
rect 3023 30202 3083 30216
rect 3023 30144 3036 30202
rect 3070 30144 3083 30202
rect 3023 30134 3083 30144
rect 3023 30072 3036 30134
rect 3070 30072 3083 30134
rect 3023 30066 3083 30072
rect 3023 30000 3036 30066
rect 3070 30000 3083 30066
rect 3023 29998 3083 30000
rect 3023 29964 3036 29998
rect 3070 29964 3083 29998
rect 3023 29962 3083 29964
rect 3023 29896 3036 29962
rect 3070 29896 3083 29962
rect 3023 29890 3083 29896
rect 3023 29828 3036 29890
rect 3070 29828 3083 29890
rect 3023 29818 3083 29828
rect 3023 29760 3036 29818
rect 3070 29760 3083 29818
rect 3023 29746 3083 29760
rect 3023 29692 3036 29746
rect 3070 29692 3083 29746
rect 3023 29674 3083 29692
rect 3023 29624 3036 29674
rect 3070 29624 3083 29674
rect 3023 29602 3083 29624
rect 3023 29556 3036 29602
rect 3070 29556 3083 29602
rect 3023 29530 3083 29556
rect 3023 29488 3036 29530
rect 3070 29488 3083 29530
rect 3023 29458 3083 29488
rect 3023 29420 3036 29458
rect 3070 29420 3083 29458
rect 3023 29386 3083 29420
rect 3023 29352 3036 29386
rect 3070 29352 3083 29386
rect 3023 29318 3083 29352
rect 3023 29280 3036 29318
rect 3070 29280 3083 29318
rect 3023 29250 3083 29280
rect 3023 29208 3036 29250
rect 3070 29208 3083 29250
rect 3023 29182 3083 29208
rect 3023 29136 3036 29182
rect 3070 29136 3083 29182
rect 3023 29114 3083 29136
rect 3023 29064 3036 29114
rect 3070 29064 3083 29114
rect 3023 29046 3083 29064
rect 3023 28992 3036 29046
rect 3070 28992 3083 29046
rect 3023 28978 3083 28992
rect 3023 28920 3036 28978
rect 3070 28920 3083 28978
rect 3023 28910 3083 28920
rect 3023 28848 3036 28910
rect 3070 28848 3083 28910
rect 3023 28842 3083 28848
rect 3023 28776 3036 28842
rect 3070 28776 3083 28842
rect 3023 28774 3083 28776
rect 3023 28740 3036 28774
rect 3070 28740 3083 28774
rect 3023 28738 3083 28740
rect 3023 28672 3036 28738
rect 3070 28672 3083 28738
rect 3023 28666 3083 28672
rect 3023 28604 3036 28666
rect 3070 28604 3083 28666
rect 3023 28594 3083 28604
rect 3023 28536 3036 28594
rect 3070 28536 3083 28594
rect 3023 28522 3083 28536
rect 373 28447 433 28469
rect 373 28397 386 28447
rect 420 28397 433 28447
rect 3023 28468 3036 28522
rect 3070 28468 3083 28522
rect 3023 28450 3083 28468
rect 373 28379 433 28397
rect 373 28325 386 28379
rect 420 28325 433 28379
rect 576 28370 592 28404
rect 659 28370 662 28404
rect 696 28370 700 28404
rect 766 28370 775 28404
rect 836 28370 850 28404
rect 906 28370 925 28404
rect 976 28370 1000 28404
rect 1046 28370 1075 28404
rect 1116 28370 1150 28404
rect 1186 28370 1222 28404
rect 1259 28370 1292 28404
rect 1334 28370 1362 28404
rect 1409 28370 1432 28404
rect 1484 28370 1502 28404
rect 1559 28370 1572 28404
rect 1634 28370 1642 28404
rect 1708 28370 1712 28404
rect 1746 28370 1748 28404
rect 1816 28370 1822 28404
rect 1886 28370 1896 28404
rect 1956 28370 1970 28404
rect 2026 28370 2044 28404
rect 2096 28370 2118 28404
rect 2166 28370 2192 28404
rect 2236 28370 2266 28404
rect 2306 28370 2340 28404
rect 2376 28370 2412 28404
rect 2448 28370 2482 28404
rect 2522 28370 2552 28404
rect 2596 28370 2622 28404
rect 2670 28370 2692 28404
rect 2744 28370 2761 28404
rect 2818 28370 2830 28404
rect 2864 28370 2880 28404
rect 3023 28400 3036 28450
rect 3070 28400 3083 28450
rect 3023 28378 3083 28400
rect 373 28311 433 28325
rect 373 28253 386 28311
rect 420 28253 433 28311
rect 3023 28332 3036 28378
rect 3070 28332 3083 28378
rect 3023 28306 3083 28332
rect 373 28243 433 28253
rect 373 28181 386 28243
rect 420 28181 433 28243
rect 373 28175 433 28181
rect 373 28109 386 28175
rect 420 28109 433 28175
rect 373 28107 433 28109
rect 373 28073 386 28107
rect 420 28073 433 28107
rect 373 28071 433 28073
rect 373 28005 386 28071
rect 420 28005 433 28071
rect 373 27999 433 28005
rect 373 27937 386 27999
rect 420 27937 433 27999
rect 373 27927 433 27937
rect 373 27869 386 27927
rect 420 27869 433 27927
rect 373 27855 433 27869
rect 373 27801 386 27855
rect 420 27801 433 27855
rect 373 27783 433 27801
rect 373 27733 386 27783
rect 420 27733 433 27783
rect 373 27711 433 27733
rect 373 27665 386 27711
rect 420 27665 433 27711
rect 373 27639 433 27665
rect 373 27597 386 27639
rect 420 27597 433 27639
rect 373 27567 433 27597
rect 373 27529 386 27567
rect 420 27529 433 27567
rect 373 27495 433 27529
rect 373 27461 386 27495
rect 420 27461 433 27495
rect 373 27427 433 27461
rect 373 27389 386 27427
rect 420 27389 433 27427
rect 373 27359 433 27389
rect 373 27317 386 27359
rect 420 27317 433 27359
rect 373 27291 433 27317
rect 373 27245 386 27291
rect 420 27245 433 27291
rect 373 27223 433 27245
rect 373 27173 386 27223
rect 420 27173 433 27223
rect 373 27155 433 27173
rect 373 27101 386 27155
rect 420 27101 433 27155
rect 373 27087 433 27101
rect 373 27029 386 27087
rect 420 27029 433 27087
rect 373 27019 433 27029
rect 373 26957 386 27019
rect 420 26957 433 27019
rect 373 26951 433 26957
rect 373 26885 386 26951
rect 420 26885 433 26951
rect 373 26883 433 26885
rect 373 26849 386 26883
rect 420 26849 433 26883
rect 373 26847 433 26849
rect 373 26781 386 26847
rect 420 26781 433 26847
rect 373 26775 433 26781
rect 373 26713 386 26775
rect 420 26713 433 26775
rect 373 26703 433 26713
rect 373 26645 386 26703
rect 420 26645 433 26703
rect 373 26631 433 26645
rect 373 26577 386 26631
rect 420 26577 433 26631
rect 373 26559 433 26577
rect 373 26509 386 26559
rect 420 26509 433 26559
rect 373 26487 433 26509
rect 373 26441 386 26487
rect 420 26441 433 26487
rect 373 26415 433 26441
rect 373 26373 386 26415
rect 420 26373 433 26415
rect 373 26343 433 26373
rect 373 26305 386 26343
rect 420 26305 433 26343
rect 531 28215 565 28254
rect 531 28142 565 28181
rect 531 28069 565 28108
rect 531 27996 565 28035
rect 531 27923 565 27962
rect 531 27850 565 27889
rect 531 27777 565 27816
rect 531 27704 565 27743
rect 531 27631 565 27670
rect 531 27558 565 27597
rect 531 27485 565 27524
rect 531 27412 565 27451
rect 531 27338 565 27378
rect 531 27264 565 27304
rect 531 27190 565 27230
rect 531 27116 565 27156
rect 531 27042 565 27082
rect 531 26968 565 27008
rect 531 26894 565 26934
rect 531 26820 565 26860
rect 531 26746 565 26786
rect 531 26672 565 26712
rect 531 26598 565 26638
rect 531 26524 565 26564
rect 531 26450 565 26490
rect 531 26376 565 26416
rect 767 28215 801 28254
rect 767 28142 801 28181
rect 767 28069 801 28108
rect 767 27996 801 28035
rect 767 27923 801 27962
rect 767 27850 801 27889
rect 767 27777 801 27816
rect 767 27704 801 27743
rect 767 27631 801 27670
rect 767 27558 801 27597
rect 767 27485 801 27524
rect 767 27412 801 27451
rect 767 27338 801 27378
rect 767 27264 801 27304
rect 767 27190 801 27230
rect 767 27116 801 27156
rect 767 27042 801 27082
rect 767 26968 801 27008
rect 767 26894 801 26934
rect 767 26820 801 26860
rect 767 26746 801 26786
rect 767 26672 801 26712
rect 767 26598 801 26638
rect 767 26524 801 26564
rect 767 26450 801 26490
rect 767 26376 801 26416
rect 1003 28215 1037 28254
rect 1003 28142 1037 28181
rect 1003 28069 1037 28108
rect 1003 27996 1037 28035
rect 1003 27923 1037 27962
rect 1003 27850 1037 27889
rect 1003 27777 1037 27816
rect 1003 27704 1037 27743
rect 1003 27631 1037 27670
rect 1003 27558 1037 27597
rect 1003 27485 1037 27524
rect 1003 27412 1037 27451
rect 1003 27338 1037 27378
rect 1003 27264 1037 27304
rect 1003 27190 1037 27230
rect 1003 27116 1037 27156
rect 1003 27042 1037 27082
rect 1003 26968 1037 27008
rect 1003 26894 1037 26934
rect 1003 26820 1037 26860
rect 1003 26746 1037 26786
rect 1003 26672 1037 26712
rect 1003 26598 1037 26638
rect 1003 26524 1037 26564
rect 1003 26450 1037 26490
rect 1003 26376 1037 26416
rect 1239 28215 1273 28254
rect 1239 28142 1273 28181
rect 1239 28069 1273 28108
rect 1239 27996 1273 28035
rect 1239 27923 1273 27962
rect 1239 27850 1273 27889
rect 1239 27777 1273 27816
rect 1239 27704 1273 27743
rect 1239 27631 1273 27670
rect 1239 27558 1273 27597
rect 1239 27485 1273 27524
rect 1239 27412 1273 27451
rect 1239 27338 1273 27378
rect 1239 27264 1273 27304
rect 1239 27190 1273 27230
rect 1239 27116 1273 27156
rect 1239 27042 1273 27082
rect 1239 26968 1273 27008
rect 1239 26894 1273 26934
rect 1239 26820 1273 26860
rect 1239 26746 1273 26786
rect 1239 26672 1273 26712
rect 1239 26598 1273 26638
rect 1239 26524 1273 26564
rect 1239 26450 1273 26490
rect 1239 26376 1273 26416
rect 1475 28215 1509 28254
rect 1475 28142 1509 28181
rect 1475 28069 1509 28108
rect 1475 27996 1509 28035
rect 1475 27923 1509 27962
rect 1475 27850 1509 27889
rect 1475 27777 1509 27816
rect 1475 27704 1509 27743
rect 1475 27631 1509 27670
rect 1475 27558 1509 27597
rect 1475 27485 1509 27524
rect 1475 27412 1509 27451
rect 1475 27338 1509 27378
rect 1475 27264 1509 27304
rect 1475 27190 1509 27230
rect 1475 27116 1509 27156
rect 1475 27042 1509 27082
rect 1475 26968 1509 27008
rect 1475 26894 1509 26934
rect 1475 26820 1509 26860
rect 1475 26746 1509 26786
rect 1475 26672 1509 26712
rect 1475 26598 1509 26638
rect 1475 26524 1509 26564
rect 1475 26450 1509 26490
rect 1475 26376 1509 26416
rect 1711 28215 1745 28254
rect 1711 28142 1745 28181
rect 1711 28069 1745 28108
rect 1711 27996 1745 28035
rect 1711 27923 1745 27962
rect 1711 27850 1745 27889
rect 1711 27777 1745 27816
rect 1711 27704 1745 27743
rect 1711 27631 1745 27670
rect 1711 27558 1745 27597
rect 1711 27485 1745 27524
rect 1711 27412 1745 27451
rect 1711 27338 1745 27378
rect 1711 27264 1745 27304
rect 1711 27190 1745 27230
rect 1711 27116 1745 27156
rect 1711 27042 1745 27082
rect 1711 26968 1745 27008
rect 1711 26894 1745 26934
rect 1711 26820 1745 26860
rect 1711 26746 1745 26786
rect 1711 26672 1745 26712
rect 1711 26598 1745 26638
rect 1711 26524 1745 26564
rect 1711 26450 1745 26490
rect 1711 26376 1745 26416
rect 1947 28215 1981 28254
rect 1947 28142 1981 28181
rect 1947 28069 1981 28108
rect 1947 27996 1981 28035
rect 1947 27923 1981 27962
rect 1947 27850 1981 27889
rect 1947 27777 1981 27816
rect 1947 27704 1981 27743
rect 1947 27631 1981 27670
rect 1947 27558 1981 27597
rect 1947 27485 1981 27524
rect 1947 27412 1981 27451
rect 1947 27338 1981 27378
rect 1947 27264 1981 27304
rect 1947 27190 1981 27230
rect 1947 27116 1981 27156
rect 1947 27042 1981 27082
rect 1947 26968 1981 27008
rect 1947 26894 1981 26934
rect 1947 26820 1981 26860
rect 1947 26746 1981 26786
rect 1947 26672 1981 26712
rect 1947 26598 1981 26638
rect 1947 26524 1981 26564
rect 1947 26450 1981 26490
rect 1947 26376 1981 26416
rect 2183 28215 2217 28254
rect 2183 28142 2217 28181
rect 2183 28069 2217 28108
rect 2183 27996 2217 28035
rect 2183 27923 2217 27962
rect 2183 27850 2217 27889
rect 2183 27777 2217 27816
rect 2183 27704 2217 27743
rect 2183 27631 2217 27670
rect 2183 27558 2217 27597
rect 2183 27485 2217 27524
rect 2183 27412 2217 27451
rect 2183 27338 2217 27378
rect 2183 27264 2217 27304
rect 2183 27190 2217 27230
rect 2183 27116 2217 27156
rect 2183 27042 2217 27082
rect 2183 26968 2217 27008
rect 2183 26894 2217 26934
rect 2183 26820 2217 26860
rect 2183 26746 2217 26786
rect 2183 26672 2217 26712
rect 2183 26598 2217 26638
rect 2183 26524 2217 26564
rect 2183 26450 2217 26490
rect 2183 26376 2217 26416
rect 2419 28215 2453 28254
rect 2419 28142 2453 28181
rect 2419 28069 2453 28108
rect 2419 27996 2453 28035
rect 2419 27923 2453 27962
rect 2419 27850 2453 27889
rect 2419 27777 2453 27816
rect 2419 27704 2453 27743
rect 2419 27631 2453 27670
rect 2419 27558 2453 27597
rect 2419 27485 2453 27524
rect 2419 27412 2453 27451
rect 2419 27338 2453 27378
rect 2419 27264 2453 27304
rect 2419 27190 2453 27230
rect 2419 27116 2453 27156
rect 2419 27042 2453 27082
rect 2419 26968 2453 27008
rect 2419 26894 2453 26934
rect 2419 26820 2453 26860
rect 2419 26746 2453 26786
rect 2419 26672 2453 26712
rect 2419 26598 2453 26638
rect 2419 26524 2453 26564
rect 2419 26450 2453 26490
rect 2419 26376 2453 26416
rect 2655 28215 2689 28254
rect 2655 28142 2689 28181
rect 2655 28069 2689 28108
rect 2655 27996 2689 28035
rect 2655 27923 2689 27962
rect 2655 27850 2689 27889
rect 2655 27777 2689 27816
rect 2655 27704 2689 27743
rect 2655 27631 2689 27670
rect 2655 27558 2689 27597
rect 2655 27485 2689 27524
rect 2655 27412 2689 27451
rect 2655 27338 2689 27378
rect 2655 27264 2689 27304
rect 2655 27190 2689 27230
rect 2655 27116 2689 27156
rect 2655 27042 2689 27082
rect 2655 26968 2689 27008
rect 2655 26894 2689 26934
rect 2655 26820 2689 26860
rect 2655 26746 2689 26786
rect 2655 26672 2689 26712
rect 2655 26598 2689 26638
rect 2655 26524 2689 26564
rect 2655 26450 2689 26490
rect 2655 26376 2689 26416
rect 2891 28215 2925 28254
rect 2891 28142 2925 28181
rect 2891 28069 2925 28108
rect 2891 27996 2925 28035
rect 2891 27923 2925 27962
rect 2891 27850 2925 27889
rect 2891 27777 2925 27816
rect 2891 27704 2925 27743
rect 2891 27631 2925 27670
rect 2891 27558 2925 27597
rect 2891 27485 2925 27524
rect 2891 27412 2925 27451
rect 2891 27338 2925 27378
rect 2891 27264 2925 27304
rect 2891 27190 2925 27230
rect 2891 27116 2925 27156
rect 2891 27042 2925 27082
rect 2891 26968 2925 27008
rect 2891 26894 2925 26934
rect 2891 26820 2925 26860
rect 2891 26746 2925 26786
rect 2891 26672 2925 26712
rect 2891 26598 2925 26638
rect 2891 26524 2925 26564
rect 2891 26450 2925 26490
rect 2891 26376 2925 26416
rect 3023 28264 3036 28306
rect 3070 28264 3083 28306
rect 3023 28234 3083 28264
rect 3023 28196 3036 28234
rect 3070 28196 3083 28234
rect 3023 28162 3083 28196
rect 3023 28128 3036 28162
rect 3070 28128 3083 28162
rect 3023 28094 3083 28128
rect 3023 28056 3036 28094
rect 3070 28056 3083 28094
rect 3023 28026 3083 28056
rect 3023 27984 3036 28026
rect 3070 27984 3083 28026
rect 3023 27958 3083 27984
rect 3023 27912 3036 27958
rect 3070 27912 3083 27958
rect 3023 27890 3083 27912
rect 3023 27840 3036 27890
rect 3070 27840 3083 27890
rect 3023 27822 3083 27840
rect 3023 27768 3036 27822
rect 3070 27768 3083 27822
rect 3023 27754 3083 27768
rect 3023 27696 3036 27754
rect 3070 27696 3083 27754
rect 3023 27686 3083 27696
rect 3023 27624 3036 27686
rect 3070 27624 3083 27686
rect 3023 27618 3083 27624
rect 3023 27552 3036 27618
rect 3070 27552 3083 27618
rect 3023 27550 3083 27552
rect 3023 27516 3036 27550
rect 3070 27516 3083 27550
rect 3023 27514 3083 27516
rect 3023 27448 3036 27514
rect 3070 27448 3083 27514
rect 3023 27442 3083 27448
rect 3023 27380 3036 27442
rect 3070 27380 3083 27442
rect 3023 27370 3083 27380
rect 3023 27312 3036 27370
rect 3070 27312 3083 27370
rect 3023 27298 3083 27312
rect 3023 27244 3036 27298
rect 3070 27244 3083 27298
rect 3023 27226 3083 27244
rect 3023 27176 3036 27226
rect 3070 27176 3083 27226
rect 3023 27154 3083 27176
rect 3023 27108 3036 27154
rect 3070 27108 3083 27154
rect 3023 27082 3083 27108
rect 3023 27040 3036 27082
rect 3070 27040 3083 27082
rect 3023 27010 3083 27040
rect 3023 26972 3036 27010
rect 3070 26972 3083 27010
rect 3023 26938 3083 26972
rect 3023 26904 3036 26938
rect 3070 26904 3083 26938
rect 3023 26870 3083 26904
rect 3023 26832 3036 26870
rect 3070 26832 3083 26870
rect 3023 26802 3083 26832
rect 3023 26760 3036 26802
rect 3070 26760 3083 26802
rect 3023 26734 3083 26760
rect 3023 26688 3036 26734
rect 3070 26688 3083 26734
rect 3023 26666 3083 26688
rect 3023 26616 3036 26666
rect 3070 26616 3083 26666
rect 3023 26598 3083 26616
rect 3023 26544 3036 26598
rect 3070 26544 3083 26598
rect 3023 26530 3083 26544
rect 3023 26472 3036 26530
rect 3070 26472 3083 26530
rect 3023 26462 3083 26472
rect 3023 26400 3036 26462
rect 3070 26400 3083 26462
rect 3023 26394 3083 26400
rect 373 26271 433 26305
rect 3023 26328 3036 26394
rect 3070 26328 3083 26394
rect 3023 26326 3083 26328
rect 3023 26292 3036 26326
rect 3070 26292 3083 26326
rect 3023 26290 3083 26292
rect 373 26237 386 26271
rect 420 26237 433 26271
rect 576 26240 592 26274
rect 659 26240 662 26274
rect 696 26240 700 26274
rect 766 26240 775 26274
rect 836 26240 850 26274
rect 906 26240 925 26274
rect 976 26240 1000 26274
rect 1046 26240 1075 26274
rect 1116 26240 1150 26274
rect 1186 26240 1222 26274
rect 1259 26240 1292 26274
rect 1334 26240 1362 26274
rect 1409 26240 1432 26274
rect 1484 26240 1502 26274
rect 1559 26240 1572 26274
rect 1634 26240 1642 26274
rect 1708 26240 1712 26274
rect 1746 26240 1748 26274
rect 1816 26240 1822 26274
rect 1886 26240 1896 26274
rect 1956 26240 1970 26274
rect 2026 26240 2044 26274
rect 2096 26240 2118 26274
rect 2166 26240 2192 26274
rect 2236 26240 2266 26274
rect 2306 26240 2340 26274
rect 2376 26240 2412 26274
rect 2448 26240 2482 26274
rect 2522 26240 2552 26274
rect 2596 26240 2622 26274
rect 2670 26240 2692 26274
rect 2744 26240 2761 26274
rect 2818 26240 2830 26274
rect 2864 26240 2880 26274
rect 373 26203 433 26237
rect 373 26165 386 26203
rect 420 26165 433 26203
rect 3023 26224 3036 26290
rect 3070 26224 3083 26290
rect 3023 26218 3083 26224
rect 373 26135 433 26165
rect 373 26093 386 26135
rect 420 26093 433 26135
rect 373 26067 433 26093
rect 373 26021 386 26067
rect 420 26021 433 26067
rect 373 25999 433 26021
rect 373 25949 386 25999
rect 420 25949 433 25999
rect 373 25931 433 25949
rect 373 25877 386 25931
rect 420 25877 433 25931
rect 373 25863 433 25877
rect 373 25805 386 25863
rect 420 25805 433 25863
rect 373 25795 433 25805
rect 373 25733 386 25795
rect 420 25733 433 25795
rect 373 25727 433 25733
rect 373 25661 386 25727
rect 420 25661 433 25727
rect 373 25659 433 25661
rect 373 25625 386 25659
rect 420 25625 433 25659
rect 373 25623 433 25625
rect 373 25557 386 25623
rect 420 25557 433 25623
rect 373 25551 433 25557
rect 373 25489 386 25551
rect 420 25489 433 25551
rect 373 25479 433 25489
rect 373 25421 386 25479
rect 420 25421 433 25479
rect 373 25407 433 25421
rect 373 25353 386 25407
rect 420 25353 433 25407
rect 373 25335 433 25353
rect 373 25285 386 25335
rect 420 25285 433 25335
rect 373 25263 433 25285
rect 373 25217 386 25263
rect 420 25217 433 25263
rect 373 25191 433 25217
rect 373 25149 386 25191
rect 420 25149 433 25191
rect 373 25119 433 25149
rect 373 25081 386 25119
rect 420 25081 433 25119
rect 373 25047 433 25081
rect 373 25013 386 25047
rect 420 25013 433 25047
rect 373 24979 433 25013
rect 373 24941 386 24979
rect 420 24941 433 24979
rect 373 24911 433 24941
rect 373 24869 386 24911
rect 420 24869 433 24911
rect 373 24843 433 24869
rect 373 24797 386 24843
rect 420 24797 433 24843
rect 373 24775 433 24797
rect 373 24725 386 24775
rect 420 24725 433 24775
rect 373 24707 433 24725
rect 373 24653 386 24707
rect 420 24653 433 24707
rect 373 24639 433 24653
rect 373 24581 386 24639
rect 420 24581 433 24639
rect 373 24571 433 24581
rect 373 24509 386 24571
rect 420 24509 433 24571
rect 373 24503 433 24509
rect 373 24437 386 24503
rect 420 24437 433 24503
rect 373 24435 433 24437
rect 373 24401 386 24435
rect 420 24401 433 24435
rect 373 24399 433 24401
rect 373 24333 386 24399
rect 420 24333 433 24399
rect 373 24327 433 24333
rect 373 24265 386 24327
rect 420 24265 433 24327
rect 373 24255 433 24265
rect 373 24197 386 24255
rect 420 24197 433 24255
rect 531 26099 565 26138
rect 531 26026 565 26065
rect 531 25953 565 25992
rect 531 25880 565 25919
rect 531 25807 565 25846
rect 531 25734 565 25773
rect 531 25661 565 25700
rect 531 25588 565 25627
rect 531 25515 565 25554
rect 531 25442 565 25481
rect 531 25369 565 25408
rect 531 25296 565 25335
rect 531 25222 565 25262
rect 531 25148 565 25188
rect 531 25074 565 25114
rect 531 25000 565 25040
rect 531 24926 565 24966
rect 531 24852 565 24892
rect 531 24778 565 24818
rect 531 24704 565 24744
rect 531 24630 565 24670
rect 531 24556 565 24596
rect 531 24482 565 24522
rect 531 24408 565 24448
rect 531 24334 565 24374
rect 531 24260 565 24300
rect 767 26099 801 26138
rect 767 26026 801 26065
rect 767 25953 801 25992
rect 767 25880 801 25919
rect 767 25807 801 25846
rect 767 25734 801 25773
rect 767 25661 801 25700
rect 767 25588 801 25627
rect 767 25515 801 25554
rect 767 25442 801 25481
rect 767 25369 801 25408
rect 767 25296 801 25335
rect 767 25222 801 25262
rect 767 25148 801 25188
rect 767 25074 801 25114
rect 767 25000 801 25040
rect 767 24926 801 24966
rect 767 24852 801 24892
rect 767 24778 801 24818
rect 767 24704 801 24744
rect 767 24630 801 24670
rect 767 24556 801 24596
rect 767 24482 801 24522
rect 767 24408 801 24448
rect 767 24334 801 24374
rect 767 24260 801 24300
rect 1003 26099 1037 26138
rect 1003 26026 1037 26065
rect 1003 25953 1037 25992
rect 1003 25880 1037 25919
rect 1003 25807 1037 25846
rect 1003 25734 1037 25773
rect 1003 25661 1037 25700
rect 1003 25588 1037 25627
rect 1003 25515 1037 25554
rect 1003 25442 1037 25481
rect 1003 25369 1037 25408
rect 1003 25296 1037 25335
rect 1003 25222 1037 25262
rect 1003 25148 1037 25188
rect 1003 25074 1037 25114
rect 1003 25000 1037 25040
rect 1003 24926 1037 24966
rect 1003 24852 1037 24892
rect 1003 24778 1037 24818
rect 1003 24704 1037 24744
rect 1003 24630 1037 24670
rect 1003 24556 1037 24596
rect 1003 24482 1037 24522
rect 1003 24408 1037 24448
rect 1003 24334 1037 24374
rect 1003 24260 1037 24300
rect 1239 26099 1273 26138
rect 1239 26026 1273 26065
rect 1239 25953 1273 25992
rect 1239 25880 1273 25919
rect 1239 25807 1273 25846
rect 1239 25734 1273 25773
rect 1239 25661 1273 25700
rect 1239 25588 1273 25627
rect 1239 25515 1273 25554
rect 1239 25442 1273 25481
rect 1239 25369 1273 25408
rect 1239 25296 1273 25335
rect 1239 25222 1273 25262
rect 1239 25148 1273 25188
rect 1239 25074 1273 25114
rect 1239 25000 1273 25040
rect 1239 24926 1273 24966
rect 1239 24852 1273 24892
rect 1239 24778 1273 24818
rect 1239 24704 1273 24744
rect 1239 24630 1273 24670
rect 1239 24556 1273 24596
rect 1239 24482 1273 24522
rect 1239 24408 1273 24448
rect 1239 24334 1273 24374
rect 1239 24260 1273 24300
rect 1475 26099 1509 26138
rect 1475 26026 1509 26065
rect 1475 25953 1509 25992
rect 1475 25880 1509 25919
rect 1475 25807 1509 25846
rect 1475 25734 1509 25773
rect 1475 25661 1509 25700
rect 1475 25588 1509 25627
rect 1475 25515 1509 25554
rect 1475 25442 1509 25481
rect 1475 25369 1509 25408
rect 1475 25296 1509 25335
rect 1475 25222 1509 25262
rect 1475 25148 1509 25188
rect 1475 25074 1509 25114
rect 1475 25000 1509 25040
rect 1475 24926 1509 24966
rect 1475 24852 1509 24892
rect 1475 24778 1509 24818
rect 1475 24704 1509 24744
rect 1475 24630 1509 24670
rect 1475 24556 1509 24596
rect 1475 24482 1509 24522
rect 1475 24408 1509 24448
rect 1475 24334 1509 24374
rect 1475 24260 1509 24300
rect 1711 26099 1745 26138
rect 1711 26026 1745 26065
rect 1711 25953 1745 25992
rect 1711 25880 1745 25919
rect 1711 25807 1745 25846
rect 1711 25734 1745 25773
rect 1711 25661 1745 25700
rect 1711 25588 1745 25627
rect 1711 25515 1745 25554
rect 1711 25442 1745 25481
rect 1711 25369 1745 25408
rect 1711 25296 1745 25335
rect 1711 25222 1745 25262
rect 1711 25148 1745 25188
rect 1711 25074 1745 25114
rect 1711 25000 1745 25040
rect 1711 24926 1745 24966
rect 1711 24852 1745 24892
rect 1711 24778 1745 24818
rect 1711 24704 1745 24744
rect 1711 24630 1745 24670
rect 1711 24556 1745 24596
rect 1711 24482 1745 24522
rect 1711 24408 1745 24448
rect 1711 24334 1745 24374
rect 1711 24260 1745 24300
rect 1947 26099 1981 26138
rect 1947 26026 1981 26065
rect 1947 25953 1981 25992
rect 1947 25880 1981 25919
rect 1947 25807 1981 25846
rect 1947 25734 1981 25773
rect 1947 25661 1981 25700
rect 1947 25588 1981 25627
rect 1947 25515 1981 25554
rect 1947 25442 1981 25481
rect 1947 25369 1981 25408
rect 1947 25296 1981 25335
rect 1947 25222 1981 25262
rect 1947 25148 1981 25188
rect 1947 25074 1981 25114
rect 1947 25000 1981 25040
rect 1947 24926 1981 24966
rect 1947 24852 1981 24892
rect 1947 24778 1981 24818
rect 1947 24704 1981 24744
rect 1947 24630 1981 24670
rect 1947 24556 1981 24596
rect 1947 24482 1981 24522
rect 1947 24408 1981 24448
rect 1947 24334 1981 24374
rect 1947 24260 1981 24300
rect 2183 26099 2217 26138
rect 2183 26026 2217 26065
rect 2183 25953 2217 25992
rect 2183 25880 2217 25919
rect 2183 25807 2217 25846
rect 2183 25734 2217 25773
rect 2183 25661 2217 25700
rect 2183 25588 2217 25627
rect 2183 25515 2217 25554
rect 2183 25442 2217 25481
rect 2183 25369 2217 25408
rect 2183 25296 2217 25335
rect 2183 25222 2217 25262
rect 2183 25148 2217 25188
rect 2183 25074 2217 25114
rect 2183 25000 2217 25040
rect 2183 24926 2217 24966
rect 2183 24852 2217 24892
rect 2183 24778 2217 24818
rect 2183 24704 2217 24744
rect 2183 24630 2217 24670
rect 2183 24556 2217 24596
rect 2183 24482 2217 24522
rect 2183 24408 2217 24448
rect 2183 24334 2217 24374
rect 2183 24260 2217 24300
rect 2419 26099 2453 26138
rect 2419 26026 2453 26065
rect 2419 25953 2453 25992
rect 2419 25880 2453 25919
rect 2419 25807 2453 25846
rect 2419 25734 2453 25773
rect 2419 25661 2453 25700
rect 2419 25588 2453 25627
rect 2419 25515 2453 25554
rect 2419 25442 2453 25481
rect 2419 25369 2453 25408
rect 2419 25296 2453 25335
rect 2419 25222 2453 25262
rect 2419 25148 2453 25188
rect 2419 25074 2453 25114
rect 2419 25000 2453 25040
rect 2419 24926 2453 24966
rect 2419 24852 2453 24892
rect 2419 24778 2453 24818
rect 2419 24704 2453 24744
rect 2419 24630 2453 24670
rect 2419 24556 2453 24596
rect 2419 24482 2453 24522
rect 2419 24408 2453 24448
rect 2419 24334 2453 24374
rect 2419 24260 2453 24300
rect 2655 26099 2689 26138
rect 2655 26026 2689 26065
rect 2655 25953 2689 25992
rect 2655 25880 2689 25919
rect 2655 25807 2689 25846
rect 2655 25734 2689 25773
rect 2655 25661 2689 25700
rect 2655 25588 2689 25627
rect 2655 25515 2689 25554
rect 2655 25442 2689 25481
rect 2655 25369 2689 25408
rect 2655 25296 2689 25335
rect 2655 25222 2689 25262
rect 2655 25148 2689 25188
rect 2655 25074 2689 25114
rect 2655 25000 2689 25040
rect 2655 24926 2689 24966
rect 2655 24852 2689 24892
rect 2655 24778 2689 24818
rect 2655 24704 2689 24744
rect 2655 24630 2689 24670
rect 2655 24556 2689 24596
rect 2655 24482 2689 24522
rect 2655 24408 2689 24448
rect 2655 24334 2689 24374
rect 2655 24260 2689 24300
rect 2891 26099 2925 26138
rect 2891 26026 2925 26065
rect 2891 25953 2925 25992
rect 2891 25880 2925 25919
rect 2891 25807 2925 25846
rect 2891 25734 2925 25773
rect 2891 25661 2925 25700
rect 2891 25588 2925 25627
rect 2891 25515 2925 25554
rect 2891 25442 2925 25481
rect 2891 25369 2925 25408
rect 2891 25296 2925 25335
rect 2891 25222 2925 25262
rect 2891 25148 2925 25188
rect 2891 25074 2925 25114
rect 2891 25000 2925 25040
rect 2891 24926 2925 24966
rect 2891 24852 2925 24892
rect 2891 24778 2925 24818
rect 2891 24704 2925 24744
rect 2891 24630 2925 24670
rect 2891 24556 2925 24596
rect 2891 24482 2925 24522
rect 2891 24408 2925 24448
rect 2891 24334 2925 24374
rect 2891 24260 2925 24300
rect 3023 26156 3036 26218
rect 3070 26156 3083 26218
rect 3023 26146 3083 26156
rect 3023 26088 3036 26146
rect 3070 26088 3083 26146
rect 3023 26074 3083 26088
rect 3023 26020 3036 26074
rect 3070 26020 3083 26074
rect 3023 26002 3083 26020
rect 3023 25952 3036 26002
rect 3070 25952 3083 26002
rect 3023 25930 3083 25952
rect 3023 25884 3036 25930
rect 3070 25884 3083 25930
rect 3023 25858 3083 25884
rect 3023 25816 3036 25858
rect 3070 25816 3083 25858
rect 3023 25786 3083 25816
rect 3023 25748 3036 25786
rect 3070 25748 3083 25786
rect 3023 25714 3083 25748
rect 3023 25680 3036 25714
rect 3070 25680 3083 25714
rect 3023 25646 3083 25680
rect 3023 25608 3036 25646
rect 3070 25608 3083 25646
rect 3023 25578 3083 25608
rect 3023 25536 3036 25578
rect 3070 25536 3083 25578
rect 3023 25510 3083 25536
rect 3023 25464 3036 25510
rect 3070 25464 3083 25510
rect 3023 25442 3083 25464
rect 3023 25392 3036 25442
rect 3070 25392 3083 25442
rect 3023 25374 3083 25392
rect 3023 25320 3036 25374
rect 3070 25320 3083 25374
rect 3023 25306 3083 25320
rect 3023 25248 3036 25306
rect 3070 25248 3083 25306
rect 3023 25238 3083 25248
rect 3023 25176 3036 25238
rect 3070 25176 3083 25238
rect 3023 25170 3083 25176
rect 3023 25104 3036 25170
rect 3070 25104 3083 25170
rect 3023 25102 3083 25104
rect 3023 25068 3036 25102
rect 3070 25068 3083 25102
rect 3023 25066 3083 25068
rect 3023 25000 3036 25066
rect 3070 25000 3083 25066
rect 3023 24994 3083 25000
rect 3023 24932 3036 24994
rect 3070 24932 3083 24994
rect 3023 24922 3083 24932
rect 3023 24864 3036 24922
rect 3070 24864 3083 24922
rect 3023 24850 3083 24864
rect 3023 24796 3036 24850
rect 3070 24796 3083 24850
rect 3023 24778 3083 24796
rect 3023 24728 3036 24778
rect 3070 24728 3083 24778
rect 3023 24706 3083 24728
rect 3023 24660 3036 24706
rect 3070 24660 3083 24706
rect 3023 24634 3083 24660
rect 3023 24592 3036 24634
rect 3070 24592 3083 24634
rect 3023 24562 3083 24592
rect 3023 24524 3036 24562
rect 3070 24524 3083 24562
rect 3023 24490 3083 24524
rect 3023 24456 3036 24490
rect 3070 24456 3083 24490
rect 3023 24422 3083 24456
rect 3023 24384 3036 24422
rect 3070 24384 3083 24422
rect 3023 24354 3083 24384
rect 3023 24312 3036 24354
rect 3070 24312 3083 24354
rect 3023 24286 3083 24312
rect 3023 24240 3036 24286
rect 3070 24240 3083 24286
rect 373 24183 433 24197
rect 373 24129 386 24183
rect 420 24129 433 24183
rect 3023 24218 3083 24240
rect 3023 24168 3036 24218
rect 3070 24168 3083 24218
rect 3023 24150 3083 24168
rect 373 24111 433 24129
rect 373 24061 386 24111
rect 420 24061 433 24111
rect 576 24110 592 24144
rect 659 24110 662 24144
rect 696 24110 700 24144
rect 766 24110 775 24144
rect 836 24110 850 24144
rect 906 24110 925 24144
rect 976 24110 1000 24144
rect 1046 24110 1075 24144
rect 1116 24110 1150 24144
rect 1186 24110 1222 24144
rect 1259 24110 1292 24144
rect 1334 24110 1362 24144
rect 1409 24110 1432 24144
rect 1484 24110 1502 24144
rect 1559 24110 1572 24144
rect 1634 24110 1642 24144
rect 1708 24110 1712 24144
rect 1746 24110 1748 24144
rect 1816 24110 1822 24144
rect 1886 24110 1896 24144
rect 1956 24110 1970 24144
rect 2026 24110 2044 24144
rect 2096 24110 2118 24144
rect 2166 24110 2192 24144
rect 2236 24110 2266 24144
rect 2306 24110 2340 24144
rect 2376 24110 2412 24144
rect 2448 24110 2482 24144
rect 2522 24110 2552 24144
rect 2596 24110 2622 24144
rect 2670 24110 2692 24144
rect 2744 24110 2761 24144
rect 2818 24110 2830 24144
rect 2864 24110 2880 24144
rect 373 24039 433 24061
rect 373 23993 386 24039
rect 420 23993 433 24039
rect 3023 24096 3036 24150
rect 3070 24096 3083 24150
rect 3023 24082 3083 24096
rect 373 23967 433 23993
rect 373 23925 386 23967
rect 420 23925 433 23967
rect 373 23895 433 23925
rect 373 23857 386 23895
rect 420 23857 433 23895
rect 373 23823 433 23857
rect 373 23789 386 23823
rect 420 23789 433 23823
rect 373 23755 433 23789
rect 373 23717 386 23755
rect 420 23717 433 23755
rect 373 23687 433 23717
rect 373 23645 386 23687
rect 420 23645 433 23687
rect 373 23619 433 23645
rect 373 23573 386 23619
rect 420 23573 433 23619
rect 373 23551 433 23573
rect 373 23501 386 23551
rect 420 23501 433 23551
rect 373 23483 433 23501
rect 373 23429 386 23483
rect 420 23429 433 23483
rect 373 23415 433 23429
rect 373 23357 386 23415
rect 420 23357 433 23415
rect 373 23347 433 23357
rect 373 23285 386 23347
rect 420 23285 433 23347
rect 373 23279 433 23285
rect 373 23213 386 23279
rect 420 23213 433 23279
rect 373 23211 433 23213
rect 373 23177 386 23211
rect 420 23177 433 23211
rect 373 23175 433 23177
rect 373 23109 386 23175
rect 420 23109 433 23175
rect 373 23103 433 23109
rect 373 23041 386 23103
rect 420 23041 433 23103
rect 373 23031 433 23041
rect 373 22973 386 23031
rect 420 22973 433 23031
rect 373 22959 433 22973
rect 373 22905 386 22959
rect 420 22905 433 22959
rect 373 22887 433 22905
rect 373 22837 386 22887
rect 420 22837 433 22887
rect 373 22815 433 22837
rect 373 22769 386 22815
rect 420 22769 433 22815
rect 373 22743 433 22769
rect 373 22701 386 22743
rect 420 22701 433 22743
rect 373 22671 433 22701
rect 373 22633 386 22671
rect 420 22633 433 22671
rect 373 22599 433 22633
rect 373 22565 386 22599
rect 420 22565 433 22599
rect 373 22531 433 22565
rect 373 22493 386 22531
rect 420 22493 433 22531
rect 373 22463 433 22493
rect 373 22421 386 22463
rect 420 22421 433 22463
rect 373 22395 433 22421
rect 373 22349 386 22395
rect 420 22349 433 22395
rect 373 22327 433 22349
rect 373 22277 386 22327
rect 420 22277 433 22327
rect 373 22259 433 22277
rect 373 22205 386 22259
rect 420 22205 433 22259
rect 373 22191 433 22205
rect 373 22133 386 22191
rect 420 22133 433 22191
rect 373 22123 433 22133
rect 373 22061 386 22123
rect 420 22061 433 22123
rect 531 23955 565 23994
rect 531 23882 565 23921
rect 531 23809 565 23848
rect 531 23736 565 23775
rect 531 23663 565 23702
rect 531 23590 565 23629
rect 531 23517 565 23556
rect 531 23444 565 23483
rect 531 23371 565 23410
rect 531 23298 565 23337
rect 531 23225 565 23264
rect 531 23152 565 23191
rect 531 23078 565 23118
rect 531 23004 565 23044
rect 531 22930 565 22970
rect 531 22856 565 22896
rect 531 22782 565 22822
rect 531 22708 565 22748
rect 531 22634 565 22674
rect 531 22560 565 22600
rect 531 22486 565 22526
rect 531 22412 565 22452
rect 531 22338 565 22378
rect 531 22264 565 22304
rect 531 22190 565 22230
rect 531 22116 565 22156
rect 767 23955 801 23994
rect 767 23882 801 23921
rect 767 23809 801 23848
rect 767 23736 801 23775
rect 767 23663 801 23702
rect 767 23590 801 23629
rect 767 23517 801 23556
rect 767 23444 801 23483
rect 767 23371 801 23410
rect 767 23298 801 23337
rect 767 23225 801 23264
rect 767 23152 801 23191
rect 767 23078 801 23118
rect 767 23004 801 23044
rect 767 22930 801 22970
rect 767 22856 801 22896
rect 767 22782 801 22822
rect 767 22708 801 22748
rect 767 22634 801 22674
rect 767 22560 801 22600
rect 767 22486 801 22526
rect 767 22412 801 22452
rect 767 22338 801 22378
rect 767 22264 801 22304
rect 767 22190 801 22230
rect 767 22116 801 22156
rect 1003 23955 1037 23994
rect 1003 23882 1037 23921
rect 1003 23809 1037 23848
rect 1003 23736 1037 23775
rect 1003 23663 1037 23702
rect 1003 23590 1037 23629
rect 1003 23517 1037 23556
rect 1003 23444 1037 23483
rect 1003 23371 1037 23410
rect 1003 23298 1037 23337
rect 1003 23225 1037 23264
rect 1003 23152 1037 23191
rect 1003 23078 1037 23118
rect 1003 23004 1037 23044
rect 1003 22930 1037 22970
rect 1003 22856 1037 22896
rect 1003 22782 1037 22822
rect 1003 22708 1037 22748
rect 1003 22634 1037 22674
rect 1003 22560 1037 22600
rect 1003 22486 1037 22526
rect 1003 22412 1037 22452
rect 1003 22338 1037 22378
rect 1003 22264 1037 22304
rect 1003 22190 1037 22230
rect 1003 22116 1037 22156
rect 1239 23955 1273 23994
rect 1239 23882 1273 23921
rect 1239 23809 1273 23848
rect 1239 23736 1273 23775
rect 1239 23663 1273 23702
rect 1239 23590 1273 23629
rect 1239 23517 1273 23556
rect 1239 23444 1273 23483
rect 1239 23371 1273 23410
rect 1239 23298 1273 23337
rect 1239 23225 1273 23264
rect 1239 23152 1273 23191
rect 1239 23078 1273 23118
rect 1239 23004 1273 23044
rect 1239 22930 1273 22970
rect 1239 22856 1273 22896
rect 1239 22782 1273 22822
rect 1239 22708 1273 22748
rect 1239 22634 1273 22674
rect 1239 22560 1273 22600
rect 1239 22486 1273 22526
rect 1239 22412 1273 22452
rect 1239 22338 1273 22378
rect 1239 22264 1273 22304
rect 1239 22190 1273 22230
rect 1239 22116 1273 22156
rect 1475 23955 1509 23994
rect 1475 23882 1509 23921
rect 1475 23809 1509 23848
rect 1475 23736 1509 23775
rect 1475 23663 1509 23702
rect 1475 23590 1509 23629
rect 1475 23517 1509 23556
rect 1475 23444 1509 23483
rect 1475 23371 1509 23410
rect 1475 23298 1509 23337
rect 1475 23225 1509 23264
rect 1475 23152 1509 23191
rect 1475 23078 1509 23118
rect 1475 23004 1509 23044
rect 1475 22930 1509 22970
rect 1475 22856 1509 22896
rect 1475 22782 1509 22822
rect 1475 22708 1509 22748
rect 1475 22634 1509 22674
rect 1475 22560 1509 22600
rect 1475 22486 1509 22526
rect 1475 22412 1509 22452
rect 1475 22338 1509 22378
rect 1475 22264 1509 22304
rect 1475 22190 1509 22230
rect 1475 22116 1509 22156
rect 1711 23955 1745 23994
rect 1711 23882 1745 23921
rect 1711 23809 1745 23848
rect 1711 23736 1745 23775
rect 1711 23663 1745 23702
rect 1711 23590 1745 23629
rect 1711 23517 1745 23556
rect 1711 23444 1745 23483
rect 1711 23371 1745 23410
rect 1711 23298 1745 23337
rect 1711 23225 1745 23264
rect 1711 23152 1745 23191
rect 1711 23078 1745 23118
rect 1711 23004 1745 23044
rect 1711 22930 1745 22970
rect 1711 22856 1745 22896
rect 1711 22782 1745 22822
rect 1711 22708 1745 22748
rect 1711 22634 1745 22674
rect 1711 22560 1745 22600
rect 1711 22486 1745 22526
rect 1711 22412 1745 22452
rect 1711 22338 1745 22378
rect 1711 22264 1745 22304
rect 1711 22190 1745 22230
rect 1711 22116 1745 22156
rect 1947 23955 1981 23994
rect 1947 23882 1981 23921
rect 1947 23809 1981 23848
rect 1947 23736 1981 23775
rect 1947 23663 1981 23702
rect 1947 23590 1981 23629
rect 1947 23517 1981 23556
rect 1947 23444 1981 23483
rect 1947 23371 1981 23410
rect 1947 23298 1981 23337
rect 1947 23225 1981 23264
rect 1947 23152 1981 23191
rect 1947 23078 1981 23118
rect 1947 23004 1981 23044
rect 1947 22930 1981 22970
rect 1947 22856 1981 22896
rect 1947 22782 1981 22822
rect 1947 22708 1981 22748
rect 1947 22634 1981 22674
rect 1947 22560 1981 22600
rect 1947 22486 1981 22526
rect 1947 22412 1981 22452
rect 1947 22338 1981 22378
rect 1947 22264 1981 22304
rect 1947 22190 1981 22230
rect 1947 22116 1981 22156
rect 2183 23955 2217 23994
rect 2183 23882 2217 23921
rect 2183 23809 2217 23848
rect 2183 23736 2217 23775
rect 2183 23663 2217 23702
rect 2183 23590 2217 23629
rect 2183 23517 2217 23556
rect 2183 23444 2217 23483
rect 2183 23371 2217 23410
rect 2183 23298 2217 23337
rect 2183 23225 2217 23264
rect 2183 23152 2217 23191
rect 2183 23078 2217 23118
rect 2183 23004 2217 23044
rect 2183 22930 2217 22970
rect 2183 22856 2217 22896
rect 2183 22782 2217 22822
rect 2183 22708 2217 22748
rect 2183 22634 2217 22674
rect 2183 22560 2217 22600
rect 2183 22486 2217 22526
rect 2183 22412 2217 22452
rect 2183 22338 2217 22378
rect 2183 22264 2217 22304
rect 2183 22190 2217 22230
rect 2183 22116 2217 22156
rect 2419 23955 2453 23994
rect 2419 23882 2453 23921
rect 2419 23809 2453 23848
rect 2419 23736 2453 23775
rect 2419 23663 2453 23702
rect 2419 23590 2453 23629
rect 2419 23517 2453 23556
rect 2419 23444 2453 23483
rect 2419 23371 2453 23410
rect 2419 23298 2453 23337
rect 2419 23225 2453 23264
rect 2419 23152 2453 23191
rect 2419 23078 2453 23118
rect 2419 23004 2453 23044
rect 2419 22930 2453 22970
rect 2419 22856 2453 22896
rect 2419 22782 2453 22822
rect 2419 22708 2453 22748
rect 2419 22634 2453 22674
rect 2419 22560 2453 22600
rect 2419 22486 2453 22526
rect 2419 22412 2453 22452
rect 2419 22338 2453 22378
rect 2419 22264 2453 22304
rect 2419 22190 2453 22230
rect 2419 22116 2453 22156
rect 2655 23955 2689 23994
rect 2655 23882 2689 23921
rect 2655 23809 2689 23848
rect 2655 23736 2689 23775
rect 2655 23663 2689 23702
rect 2655 23590 2689 23629
rect 2655 23517 2689 23556
rect 2655 23444 2689 23483
rect 2655 23371 2689 23410
rect 2655 23298 2689 23337
rect 2655 23225 2689 23264
rect 2655 23152 2689 23191
rect 2655 23078 2689 23118
rect 2655 23004 2689 23044
rect 2655 22930 2689 22970
rect 2655 22856 2689 22896
rect 2655 22782 2689 22822
rect 2655 22708 2689 22748
rect 2655 22634 2689 22674
rect 2655 22560 2689 22600
rect 2655 22486 2689 22526
rect 2655 22412 2689 22452
rect 2655 22338 2689 22378
rect 2655 22264 2689 22304
rect 2655 22190 2689 22230
rect 2655 22116 2689 22156
rect 2891 23955 2925 23994
rect 2891 23882 2925 23921
rect 2891 23809 2925 23848
rect 2891 23736 2925 23775
rect 2891 23663 2925 23702
rect 2891 23590 2925 23629
rect 2891 23517 2925 23556
rect 2891 23444 2925 23483
rect 2891 23371 2925 23410
rect 2891 23298 2925 23337
rect 2891 23225 2925 23264
rect 2891 23152 2925 23191
rect 2891 23078 2925 23118
rect 2891 23004 2925 23044
rect 2891 22930 2925 22970
rect 2891 22856 2925 22896
rect 2891 22782 2925 22822
rect 2891 22708 2925 22748
rect 2891 22634 2925 22674
rect 2891 22560 2925 22600
rect 2891 22486 2925 22526
rect 2891 22412 2925 22452
rect 2891 22338 2925 22378
rect 2891 22264 2925 22304
rect 2891 22190 2925 22230
rect 2891 22116 2925 22156
rect 3023 24024 3036 24082
rect 3070 24024 3083 24082
rect 3023 24014 3083 24024
rect 3023 23952 3036 24014
rect 3070 23952 3083 24014
rect 3023 23946 3083 23952
rect 3023 23880 3036 23946
rect 3070 23880 3083 23946
rect 3023 23878 3083 23880
rect 3023 23844 3036 23878
rect 3070 23844 3083 23878
rect 3023 23842 3083 23844
rect 3023 23776 3036 23842
rect 3070 23776 3083 23842
rect 3023 23770 3083 23776
rect 3023 23708 3036 23770
rect 3070 23708 3083 23770
rect 3023 23698 3083 23708
rect 3023 23640 3036 23698
rect 3070 23640 3083 23698
rect 3023 23626 3083 23640
rect 3023 23572 3036 23626
rect 3070 23572 3083 23626
rect 3023 23554 3083 23572
rect 3023 23504 3036 23554
rect 3070 23504 3083 23554
rect 3023 23482 3083 23504
rect 3023 23436 3036 23482
rect 3070 23436 3083 23482
rect 3023 23410 3083 23436
rect 3023 23368 3036 23410
rect 3070 23368 3083 23410
rect 3023 23338 3083 23368
rect 3023 23300 3036 23338
rect 3070 23300 3083 23338
rect 3023 23266 3083 23300
rect 3023 23232 3036 23266
rect 3070 23232 3083 23266
rect 3023 23198 3083 23232
rect 3023 23160 3036 23198
rect 3070 23160 3083 23198
rect 3023 23130 3083 23160
rect 3023 23088 3036 23130
rect 3070 23088 3083 23130
rect 3023 23062 3083 23088
rect 3023 23016 3036 23062
rect 3070 23016 3083 23062
rect 3023 22994 3083 23016
rect 3023 22944 3036 22994
rect 3070 22944 3083 22994
rect 3023 22926 3083 22944
rect 3023 22872 3036 22926
rect 3070 22872 3083 22926
rect 3023 22858 3083 22872
rect 3023 22800 3036 22858
rect 3070 22800 3083 22858
rect 3023 22790 3083 22800
rect 3023 22728 3036 22790
rect 3070 22728 3083 22790
rect 3023 22722 3083 22728
rect 3023 22656 3036 22722
rect 3070 22656 3083 22722
rect 3023 22654 3083 22656
rect 3023 22620 3036 22654
rect 3070 22620 3083 22654
rect 3023 22618 3083 22620
rect 3023 22552 3036 22618
rect 3070 22552 3083 22618
rect 3023 22546 3083 22552
rect 3023 22484 3036 22546
rect 3070 22484 3083 22546
rect 3023 22474 3083 22484
rect 3023 22416 3036 22474
rect 3070 22416 3083 22474
rect 3023 22402 3083 22416
rect 3023 22348 3036 22402
rect 3070 22348 3083 22402
rect 3023 22330 3083 22348
rect 3023 22280 3036 22330
rect 3070 22280 3083 22330
rect 3023 22258 3083 22280
rect 3023 22212 3036 22258
rect 3070 22212 3083 22258
rect 3023 22186 3083 22212
rect 3023 22144 3036 22186
rect 3070 22144 3083 22186
rect 3023 22114 3083 22144
rect 373 22055 433 22061
rect 373 21989 386 22055
rect 420 21989 433 22055
rect 3023 22076 3036 22114
rect 3070 22076 3083 22114
rect 3023 22042 3083 22076
rect 373 21987 433 21989
rect 373 21953 386 21987
rect 420 21953 433 21987
rect 576 21980 592 22014
rect 659 21980 662 22014
rect 696 21980 700 22014
rect 766 21980 775 22014
rect 836 21980 850 22014
rect 906 21980 925 22014
rect 976 21980 1000 22014
rect 1046 21980 1075 22014
rect 1116 21980 1150 22014
rect 1186 21980 1222 22014
rect 1259 21980 1292 22014
rect 1334 21980 1362 22014
rect 1409 21980 1432 22014
rect 1484 21980 1502 22014
rect 1559 21980 1572 22014
rect 1634 21980 1642 22014
rect 1708 21980 1712 22014
rect 1746 21980 1748 22014
rect 1816 21980 1822 22014
rect 1886 21980 1896 22014
rect 1956 21980 1970 22014
rect 2026 21980 2044 22014
rect 2096 21980 2118 22014
rect 2166 21980 2192 22014
rect 2236 21980 2266 22014
rect 2306 21980 2340 22014
rect 2376 21980 2412 22014
rect 2448 21980 2482 22014
rect 2522 21980 2552 22014
rect 2596 21980 2622 22014
rect 2670 21980 2692 22014
rect 2744 21980 2761 22014
rect 2818 21980 2830 22014
rect 2864 21980 2880 22014
rect 3023 22008 3036 22042
rect 3070 22008 3083 22042
rect 373 21951 433 21953
rect 373 21885 386 21951
rect 420 21885 433 21951
rect 3023 21974 3083 22008
rect 3023 21936 3036 21974
rect 3070 21936 3083 21974
rect 373 21879 433 21885
rect 373 21817 386 21879
rect 420 21817 433 21879
rect 373 21807 433 21817
rect 373 21749 386 21807
rect 420 21749 433 21807
rect 373 21735 433 21749
rect 373 21681 386 21735
rect 420 21681 433 21735
rect 373 21663 433 21681
rect 373 21613 386 21663
rect 420 21613 433 21663
rect 373 21591 433 21613
rect 373 21545 386 21591
rect 420 21545 433 21591
rect 373 21519 433 21545
rect 373 21477 386 21519
rect 420 21477 433 21519
rect 373 21447 433 21477
rect 373 21409 386 21447
rect 420 21409 433 21447
rect 373 21375 433 21409
rect 373 21341 386 21375
rect 420 21341 433 21375
rect 373 21307 433 21341
rect 373 21269 386 21307
rect 420 21269 433 21307
rect 373 21239 433 21269
rect 373 21197 386 21239
rect 420 21197 433 21239
rect 373 21171 433 21197
rect 373 21125 386 21171
rect 420 21125 433 21171
rect 373 21103 433 21125
rect 373 21053 386 21103
rect 420 21053 433 21103
rect 373 21035 433 21053
rect 373 20981 386 21035
rect 420 20981 433 21035
rect 373 20967 433 20981
rect 373 20909 386 20967
rect 420 20909 433 20967
rect 373 20899 433 20909
rect 373 20837 386 20899
rect 420 20837 433 20899
rect 373 20831 433 20837
rect 373 20765 386 20831
rect 420 20765 433 20831
rect 373 20763 433 20765
rect 373 20729 386 20763
rect 420 20729 433 20763
rect 373 20727 433 20729
rect 373 20661 386 20727
rect 420 20661 433 20727
rect 373 20655 433 20661
rect 373 20593 386 20655
rect 420 20593 433 20655
rect 373 20583 433 20593
rect 373 20525 386 20583
rect 420 20525 433 20583
rect 373 20511 433 20525
rect 373 20457 386 20511
rect 420 20457 433 20511
rect 373 20439 433 20457
rect 373 20389 386 20439
rect 420 20389 433 20439
rect 373 20367 433 20389
rect 373 20321 386 20367
rect 420 20321 433 20367
rect 373 20295 433 20321
rect 373 20253 386 20295
rect 420 20253 433 20295
rect 373 20223 433 20253
rect 373 20185 386 20223
rect 420 20185 433 20223
rect 373 20151 433 20185
rect 373 20117 386 20151
rect 420 20117 433 20151
rect 373 20083 433 20117
rect 373 20045 386 20083
rect 420 20045 433 20083
rect 373 20015 433 20045
rect 373 19973 386 20015
rect 420 19973 433 20015
rect 373 19947 433 19973
rect 531 21839 565 21878
rect 531 21766 565 21805
rect 531 21693 565 21732
rect 531 21620 565 21659
rect 531 21547 565 21586
rect 531 21474 565 21513
rect 531 21401 565 21440
rect 531 21328 565 21367
rect 531 21255 565 21294
rect 531 21182 565 21221
rect 531 21109 565 21148
rect 531 21036 565 21075
rect 531 20962 565 21002
rect 531 20888 565 20928
rect 531 20814 565 20854
rect 531 20740 565 20780
rect 531 20666 565 20706
rect 531 20592 565 20632
rect 531 20518 565 20558
rect 531 20444 565 20484
rect 531 20370 565 20410
rect 531 20296 565 20336
rect 531 20222 565 20262
rect 531 20148 565 20188
rect 531 20074 565 20114
rect 531 20000 565 20040
rect 767 21839 801 21878
rect 767 21766 801 21805
rect 767 21693 801 21732
rect 767 21620 801 21659
rect 767 21547 801 21586
rect 767 21474 801 21513
rect 767 21401 801 21440
rect 767 21328 801 21367
rect 767 21255 801 21294
rect 767 21182 801 21221
rect 767 21109 801 21148
rect 767 21036 801 21075
rect 767 20962 801 21002
rect 767 20888 801 20928
rect 767 20814 801 20854
rect 767 20740 801 20780
rect 767 20666 801 20706
rect 767 20592 801 20632
rect 767 20518 801 20558
rect 767 20444 801 20484
rect 767 20370 801 20410
rect 767 20296 801 20336
rect 767 20222 801 20262
rect 767 20148 801 20188
rect 767 20074 801 20114
rect 767 20000 801 20040
rect 1003 21839 1037 21878
rect 1003 21766 1037 21805
rect 1003 21693 1037 21732
rect 1003 21620 1037 21659
rect 1003 21547 1037 21586
rect 1003 21474 1037 21513
rect 1003 21401 1037 21440
rect 1003 21328 1037 21367
rect 1003 21255 1037 21294
rect 1003 21182 1037 21221
rect 1003 21109 1037 21148
rect 1003 21036 1037 21075
rect 1003 20962 1037 21002
rect 1003 20888 1037 20928
rect 1003 20814 1037 20854
rect 1003 20740 1037 20780
rect 1003 20666 1037 20706
rect 1003 20592 1037 20632
rect 1003 20518 1037 20558
rect 1003 20444 1037 20484
rect 1003 20370 1037 20410
rect 1003 20296 1037 20336
rect 1003 20222 1037 20262
rect 1003 20148 1037 20188
rect 1003 20074 1037 20114
rect 1003 20000 1037 20040
rect 1239 21839 1273 21878
rect 1239 21766 1273 21805
rect 1239 21693 1273 21732
rect 1239 21620 1273 21659
rect 1239 21547 1273 21586
rect 1239 21474 1273 21513
rect 1239 21401 1273 21440
rect 1239 21328 1273 21367
rect 1239 21255 1273 21294
rect 1239 21182 1273 21221
rect 1239 21109 1273 21148
rect 1239 21036 1273 21075
rect 1239 20962 1273 21002
rect 1239 20888 1273 20928
rect 1239 20814 1273 20854
rect 1239 20740 1273 20780
rect 1239 20666 1273 20706
rect 1239 20592 1273 20632
rect 1239 20518 1273 20558
rect 1239 20444 1273 20484
rect 1239 20370 1273 20410
rect 1239 20296 1273 20336
rect 1239 20222 1273 20262
rect 1239 20148 1273 20188
rect 1239 20074 1273 20114
rect 1239 20000 1273 20040
rect 1475 21839 1509 21878
rect 1475 21766 1509 21805
rect 1475 21693 1509 21732
rect 1475 21620 1509 21659
rect 1475 21547 1509 21586
rect 1475 21474 1509 21513
rect 1475 21401 1509 21440
rect 1475 21328 1509 21367
rect 1475 21255 1509 21294
rect 1475 21182 1509 21221
rect 1475 21109 1509 21148
rect 1475 21036 1509 21075
rect 1475 20962 1509 21002
rect 1475 20888 1509 20928
rect 1475 20814 1509 20854
rect 1475 20740 1509 20780
rect 1475 20666 1509 20706
rect 1475 20592 1509 20632
rect 1475 20518 1509 20558
rect 1475 20444 1509 20484
rect 1475 20370 1509 20410
rect 1475 20296 1509 20336
rect 1475 20222 1509 20262
rect 1475 20148 1509 20188
rect 1475 20074 1509 20114
rect 1475 20000 1509 20040
rect 1711 21839 1745 21878
rect 1711 21766 1745 21805
rect 1711 21693 1745 21732
rect 1711 21620 1745 21659
rect 1711 21547 1745 21586
rect 1711 21474 1745 21513
rect 1711 21401 1745 21440
rect 1711 21328 1745 21367
rect 1711 21255 1745 21294
rect 1711 21182 1745 21221
rect 1711 21109 1745 21148
rect 1711 21036 1745 21075
rect 1711 20962 1745 21002
rect 1711 20888 1745 20928
rect 1711 20814 1745 20854
rect 1711 20740 1745 20780
rect 1711 20666 1745 20706
rect 1711 20592 1745 20632
rect 1711 20518 1745 20558
rect 1711 20444 1745 20484
rect 1711 20370 1745 20410
rect 1711 20296 1745 20336
rect 1711 20222 1745 20262
rect 1711 20148 1745 20188
rect 1711 20074 1745 20114
rect 1711 20000 1745 20040
rect 1947 21839 1981 21878
rect 1947 21766 1981 21805
rect 1947 21693 1981 21732
rect 1947 21620 1981 21659
rect 1947 21547 1981 21586
rect 1947 21474 1981 21513
rect 1947 21401 1981 21440
rect 1947 21328 1981 21367
rect 1947 21255 1981 21294
rect 1947 21182 1981 21221
rect 1947 21109 1981 21148
rect 1947 21036 1981 21075
rect 1947 20962 1981 21002
rect 1947 20888 1981 20928
rect 1947 20814 1981 20854
rect 1947 20740 1981 20780
rect 1947 20666 1981 20706
rect 1947 20592 1981 20632
rect 1947 20518 1981 20558
rect 1947 20444 1981 20484
rect 1947 20370 1981 20410
rect 1947 20296 1981 20336
rect 1947 20222 1981 20262
rect 1947 20148 1981 20188
rect 1947 20074 1981 20114
rect 1947 20000 1981 20040
rect 2183 21839 2217 21878
rect 2183 21766 2217 21805
rect 2183 21693 2217 21732
rect 2183 21620 2217 21659
rect 2183 21547 2217 21586
rect 2183 21474 2217 21513
rect 2183 21401 2217 21440
rect 2183 21328 2217 21367
rect 2183 21255 2217 21294
rect 2183 21182 2217 21221
rect 2183 21109 2217 21148
rect 2183 21036 2217 21075
rect 2183 20962 2217 21002
rect 2183 20888 2217 20928
rect 2183 20814 2217 20854
rect 2183 20740 2217 20780
rect 2183 20666 2217 20706
rect 2183 20592 2217 20632
rect 2183 20518 2217 20558
rect 2183 20444 2217 20484
rect 2183 20370 2217 20410
rect 2183 20296 2217 20336
rect 2183 20222 2217 20262
rect 2183 20148 2217 20188
rect 2183 20074 2217 20114
rect 2183 20000 2217 20040
rect 2419 21839 2453 21878
rect 2419 21766 2453 21805
rect 2419 21693 2453 21732
rect 2419 21620 2453 21659
rect 2419 21547 2453 21586
rect 2419 21474 2453 21513
rect 2419 21401 2453 21440
rect 2419 21328 2453 21367
rect 2419 21255 2453 21294
rect 2419 21182 2453 21221
rect 2419 21109 2453 21148
rect 2419 21036 2453 21075
rect 2419 20962 2453 21002
rect 2419 20888 2453 20928
rect 2419 20814 2453 20854
rect 2419 20740 2453 20780
rect 2419 20666 2453 20706
rect 2419 20592 2453 20632
rect 2419 20518 2453 20558
rect 2419 20444 2453 20484
rect 2419 20370 2453 20410
rect 2419 20296 2453 20336
rect 2419 20222 2453 20262
rect 2419 20148 2453 20188
rect 2419 20074 2453 20114
rect 2419 20000 2453 20040
rect 2655 21839 2689 21878
rect 2655 21766 2689 21805
rect 2655 21693 2689 21732
rect 2655 21620 2689 21659
rect 2655 21547 2689 21586
rect 2655 21474 2689 21513
rect 2655 21401 2689 21440
rect 2655 21328 2689 21367
rect 2655 21255 2689 21294
rect 2655 21182 2689 21221
rect 2655 21109 2689 21148
rect 2655 21036 2689 21075
rect 2655 20962 2689 21002
rect 2655 20888 2689 20928
rect 2655 20814 2689 20854
rect 2655 20740 2689 20780
rect 2655 20666 2689 20706
rect 2655 20592 2689 20632
rect 2655 20518 2689 20558
rect 2655 20444 2689 20484
rect 2655 20370 2689 20410
rect 2655 20296 2689 20336
rect 2655 20222 2689 20262
rect 2655 20148 2689 20188
rect 2655 20074 2689 20114
rect 2655 20000 2689 20040
rect 2891 21839 2925 21878
rect 2891 21766 2925 21805
rect 2891 21693 2925 21732
rect 2891 21620 2925 21659
rect 2891 21547 2925 21586
rect 2891 21474 2925 21513
rect 2891 21401 2925 21440
rect 2891 21328 2925 21367
rect 2891 21255 2925 21294
rect 2891 21182 2925 21221
rect 2891 21109 2925 21148
rect 2891 21036 2925 21075
rect 2891 20962 2925 21002
rect 2891 20888 2925 20928
rect 2891 20814 2925 20854
rect 2891 20740 2925 20780
rect 2891 20666 2925 20706
rect 2891 20592 2925 20632
rect 2891 20518 2925 20558
rect 2891 20444 2925 20484
rect 2891 20370 2925 20410
rect 2891 20296 2925 20336
rect 2891 20222 2925 20262
rect 2891 20148 2925 20188
rect 2891 20074 2925 20114
rect 2891 20000 2925 20040
rect 3023 21906 3083 21936
rect 3023 21864 3036 21906
rect 3070 21864 3083 21906
rect 3023 21838 3083 21864
rect 3023 21792 3036 21838
rect 3070 21792 3083 21838
rect 3023 21770 3083 21792
rect 3023 21720 3036 21770
rect 3070 21720 3083 21770
rect 3023 21702 3083 21720
rect 3023 21648 3036 21702
rect 3070 21648 3083 21702
rect 3023 21634 3083 21648
rect 3023 21576 3036 21634
rect 3070 21576 3083 21634
rect 3023 21566 3083 21576
rect 3023 21504 3036 21566
rect 3070 21504 3083 21566
rect 3023 21498 3083 21504
rect 3023 21432 3036 21498
rect 3070 21432 3083 21498
rect 3023 21430 3083 21432
rect 3023 21396 3036 21430
rect 3070 21396 3083 21430
rect 3023 21394 3083 21396
rect 3023 21328 3036 21394
rect 3070 21328 3083 21394
rect 3023 21322 3083 21328
rect 3023 21260 3036 21322
rect 3070 21260 3083 21322
rect 3023 21250 3083 21260
rect 3023 21192 3036 21250
rect 3070 21192 3083 21250
rect 3023 21178 3083 21192
rect 3023 21124 3036 21178
rect 3070 21124 3083 21178
rect 3023 21106 3083 21124
rect 3023 21056 3036 21106
rect 3070 21056 3083 21106
rect 3023 21034 3083 21056
rect 3023 20988 3036 21034
rect 3070 20988 3083 21034
rect 3023 20962 3083 20988
rect 3023 20920 3036 20962
rect 3070 20920 3083 20962
rect 3023 20890 3083 20920
rect 3023 20852 3036 20890
rect 3070 20852 3083 20890
rect 3023 20818 3083 20852
rect 3023 20784 3036 20818
rect 3070 20784 3083 20818
rect 3023 20750 3083 20784
rect 3023 20712 3036 20750
rect 3070 20712 3083 20750
rect 3023 20682 3083 20712
rect 3023 20640 3036 20682
rect 3070 20640 3083 20682
rect 3023 20614 3083 20640
rect 3023 20568 3036 20614
rect 3070 20568 3083 20614
rect 3023 20546 3083 20568
rect 3023 20496 3036 20546
rect 3070 20496 3083 20546
rect 3023 20478 3083 20496
rect 3023 20424 3036 20478
rect 3070 20424 3083 20478
rect 3023 20410 3083 20424
rect 3023 20352 3036 20410
rect 3070 20352 3083 20410
rect 3023 20342 3083 20352
rect 3023 20280 3036 20342
rect 3070 20280 3083 20342
rect 3023 20274 3083 20280
rect 3023 20208 3036 20274
rect 3070 20208 3083 20274
rect 3023 20206 3083 20208
rect 3023 20172 3036 20206
rect 3070 20172 3083 20206
rect 3023 20170 3083 20172
rect 3023 20104 3036 20170
rect 3070 20104 3083 20170
rect 3023 20098 3083 20104
rect 3023 20036 3036 20098
rect 3070 20036 3083 20098
rect 3023 20026 3083 20036
rect 3023 19968 3036 20026
rect 3070 19968 3083 20026
rect 373 19901 386 19947
rect 420 19901 433 19947
rect 373 19879 433 19901
rect 3023 19954 3083 19968
rect 3023 19900 3036 19954
rect 3070 19900 3083 19954
rect 373 19829 386 19879
rect 420 19829 433 19879
rect 576 19850 592 19884
rect 659 19850 662 19884
rect 696 19850 700 19884
rect 766 19850 775 19884
rect 836 19850 850 19884
rect 906 19850 925 19884
rect 976 19850 1000 19884
rect 1046 19850 1075 19884
rect 1116 19850 1150 19884
rect 1186 19850 1222 19884
rect 1259 19850 1292 19884
rect 1334 19850 1362 19884
rect 1409 19850 1432 19884
rect 1484 19850 1502 19884
rect 1559 19850 1572 19884
rect 1634 19850 1642 19884
rect 1708 19850 1712 19884
rect 1746 19850 1748 19884
rect 1816 19850 1822 19884
rect 1886 19850 1896 19884
rect 1956 19850 1970 19884
rect 2026 19850 2044 19884
rect 2096 19850 2118 19884
rect 2166 19850 2192 19884
rect 2236 19850 2266 19884
rect 2306 19850 2340 19884
rect 2376 19850 2412 19884
rect 2448 19850 2482 19884
rect 2522 19850 2552 19884
rect 2596 19850 2622 19884
rect 2670 19850 2692 19884
rect 2744 19850 2761 19884
rect 2818 19850 2830 19884
rect 2864 19850 2880 19884
rect 3023 19882 3083 19900
rect 373 19811 433 19829
rect 373 19757 386 19811
rect 420 19757 433 19811
rect 3023 19832 3036 19882
rect 3070 19832 3083 19882
rect 3023 19810 3083 19832
rect 373 19743 433 19757
rect 373 19685 386 19743
rect 420 19685 433 19743
rect 373 19675 433 19685
rect 373 19613 386 19675
rect 420 19613 433 19675
rect 373 19607 433 19613
rect 373 19541 386 19607
rect 420 19541 433 19607
rect 373 19539 433 19541
rect 373 19505 386 19539
rect 420 19505 433 19539
rect 373 19503 433 19505
rect 373 19437 386 19503
rect 420 19437 433 19503
rect 373 19431 433 19437
rect 373 19369 386 19431
rect 420 19369 433 19431
rect 373 19359 433 19369
rect 373 19301 386 19359
rect 420 19301 433 19359
rect 373 19287 433 19301
rect 373 19233 386 19287
rect 420 19233 433 19287
rect 373 19215 433 19233
rect 373 19165 386 19215
rect 420 19165 433 19215
rect 373 19143 433 19165
rect 373 19097 386 19143
rect 420 19097 433 19143
rect 373 19071 433 19097
rect 373 19029 386 19071
rect 420 19029 433 19071
rect 373 18999 433 19029
rect 373 18961 386 18999
rect 420 18961 433 18999
rect 373 18927 433 18961
rect 373 18893 386 18927
rect 420 18893 433 18927
rect 373 18859 433 18893
rect 373 18821 386 18859
rect 420 18821 433 18859
rect 373 18791 433 18821
rect 373 18749 386 18791
rect 420 18749 433 18791
rect 373 18723 433 18749
rect 373 18677 386 18723
rect 420 18677 433 18723
rect 373 18655 433 18677
rect 373 18605 386 18655
rect 420 18605 433 18655
rect 373 18587 433 18605
rect 373 18533 386 18587
rect 420 18533 433 18587
rect 373 18519 433 18533
rect 373 18461 386 18519
rect 420 18461 433 18519
rect 373 18451 433 18461
rect 373 18389 386 18451
rect 420 18389 433 18451
rect 373 18383 433 18389
rect 373 18317 386 18383
rect 420 18317 433 18383
rect 373 18315 433 18317
rect 373 18281 386 18315
rect 420 18281 433 18315
rect 373 18279 433 18281
rect 373 18213 386 18279
rect 420 18213 433 18279
rect 373 18207 433 18213
rect 373 18145 386 18207
rect 420 18145 433 18207
rect 373 18135 433 18145
rect 373 18077 386 18135
rect 420 18077 433 18135
rect 373 18063 433 18077
rect 373 18009 386 18063
rect 420 18009 433 18063
rect 373 17991 433 18009
rect 373 17941 386 17991
rect 420 17941 433 17991
rect 373 17919 433 17941
rect 373 17873 386 17919
rect 420 17873 433 17919
rect 373 17847 433 17873
rect 373 17805 386 17847
rect 420 17805 433 17847
rect 531 19695 565 19734
rect 531 19622 565 19661
rect 531 19549 565 19588
rect 531 19476 565 19515
rect 531 19403 565 19442
rect 531 19330 565 19369
rect 531 19257 565 19296
rect 531 19184 565 19223
rect 531 19111 565 19150
rect 531 19038 565 19077
rect 531 18965 565 19004
rect 531 18892 565 18931
rect 531 18818 565 18858
rect 531 18744 565 18784
rect 531 18670 565 18710
rect 531 18596 565 18636
rect 531 18522 565 18562
rect 531 18448 565 18488
rect 531 18374 565 18414
rect 531 18300 565 18340
rect 531 18226 565 18266
rect 531 18152 565 18192
rect 531 18078 565 18118
rect 531 18004 565 18044
rect 531 17930 565 17970
rect 531 17856 565 17896
rect 767 19695 801 19734
rect 767 19622 801 19661
rect 767 19549 801 19588
rect 767 19476 801 19515
rect 767 19403 801 19442
rect 767 19330 801 19369
rect 767 19257 801 19296
rect 767 19184 801 19223
rect 767 19111 801 19150
rect 767 19038 801 19077
rect 767 18965 801 19004
rect 767 18892 801 18931
rect 767 18818 801 18858
rect 767 18744 801 18784
rect 767 18670 801 18710
rect 767 18596 801 18636
rect 767 18522 801 18562
rect 767 18448 801 18488
rect 767 18374 801 18414
rect 767 18300 801 18340
rect 767 18226 801 18266
rect 767 18152 801 18192
rect 767 18078 801 18118
rect 767 18004 801 18044
rect 767 17930 801 17970
rect 767 17856 801 17896
rect 1003 19695 1037 19734
rect 1003 19622 1037 19661
rect 1003 19549 1037 19588
rect 1003 19476 1037 19515
rect 1003 19403 1037 19442
rect 1003 19330 1037 19369
rect 1003 19257 1037 19296
rect 1003 19184 1037 19223
rect 1003 19111 1037 19150
rect 1003 19038 1037 19077
rect 1003 18965 1037 19004
rect 1003 18892 1037 18931
rect 1003 18818 1037 18858
rect 1003 18744 1037 18784
rect 1003 18670 1037 18710
rect 1003 18596 1037 18636
rect 1003 18522 1037 18562
rect 1003 18448 1037 18488
rect 1003 18374 1037 18414
rect 1003 18300 1037 18340
rect 1003 18226 1037 18266
rect 1003 18152 1037 18192
rect 1003 18078 1037 18118
rect 1003 18004 1037 18044
rect 1003 17930 1037 17970
rect 1003 17856 1037 17896
rect 1239 19695 1273 19734
rect 1239 19622 1273 19661
rect 1239 19549 1273 19588
rect 1239 19476 1273 19515
rect 1239 19403 1273 19442
rect 1239 19330 1273 19369
rect 1239 19257 1273 19296
rect 1239 19184 1273 19223
rect 1239 19111 1273 19150
rect 1239 19038 1273 19077
rect 1239 18965 1273 19004
rect 1239 18892 1273 18931
rect 1239 18818 1273 18858
rect 1239 18744 1273 18784
rect 1239 18670 1273 18710
rect 1239 18596 1273 18636
rect 1239 18522 1273 18562
rect 1239 18448 1273 18488
rect 1239 18374 1273 18414
rect 1239 18300 1273 18340
rect 1239 18226 1273 18266
rect 1239 18152 1273 18192
rect 1239 18078 1273 18118
rect 1239 18004 1273 18044
rect 1239 17930 1273 17970
rect 1239 17856 1273 17896
rect 1475 19695 1509 19734
rect 1475 19622 1509 19661
rect 1475 19549 1509 19588
rect 1475 19476 1509 19515
rect 1475 19403 1509 19442
rect 1475 19330 1509 19369
rect 1475 19257 1509 19296
rect 1475 19184 1509 19223
rect 1475 19111 1509 19150
rect 1475 19038 1509 19077
rect 1475 18965 1509 19004
rect 1475 18892 1509 18931
rect 1475 18818 1509 18858
rect 1475 18744 1509 18784
rect 1475 18670 1509 18710
rect 1475 18596 1509 18636
rect 1475 18522 1509 18562
rect 1475 18448 1509 18488
rect 1475 18374 1509 18414
rect 1475 18300 1509 18340
rect 1475 18226 1509 18266
rect 1475 18152 1509 18192
rect 1475 18078 1509 18118
rect 1475 18004 1509 18044
rect 1475 17930 1509 17970
rect 1475 17856 1509 17896
rect 1711 19695 1745 19734
rect 1711 19622 1745 19661
rect 1711 19549 1745 19588
rect 1711 19476 1745 19515
rect 1711 19403 1745 19442
rect 1711 19330 1745 19369
rect 1711 19257 1745 19296
rect 1711 19184 1745 19223
rect 1711 19111 1745 19150
rect 1711 19038 1745 19077
rect 1711 18965 1745 19004
rect 1711 18892 1745 18931
rect 1711 18818 1745 18858
rect 1711 18744 1745 18784
rect 1711 18670 1745 18710
rect 1711 18596 1745 18636
rect 1711 18522 1745 18562
rect 1711 18448 1745 18488
rect 1711 18374 1745 18414
rect 1711 18300 1745 18340
rect 1711 18226 1745 18266
rect 1711 18152 1745 18192
rect 1711 18078 1745 18118
rect 1711 18004 1745 18044
rect 1711 17930 1745 17970
rect 1711 17856 1745 17896
rect 1947 19695 1981 19734
rect 1947 19622 1981 19661
rect 1947 19549 1981 19588
rect 1947 19476 1981 19515
rect 1947 19403 1981 19442
rect 1947 19330 1981 19369
rect 1947 19257 1981 19296
rect 1947 19184 1981 19223
rect 1947 19111 1981 19150
rect 1947 19038 1981 19077
rect 1947 18965 1981 19004
rect 1947 18892 1981 18931
rect 1947 18818 1981 18858
rect 1947 18744 1981 18784
rect 1947 18670 1981 18710
rect 1947 18596 1981 18636
rect 1947 18522 1981 18562
rect 1947 18448 1981 18488
rect 1947 18374 1981 18414
rect 1947 18300 1981 18340
rect 1947 18226 1981 18266
rect 1947 18152 1981 18192
rect 1947 18078 1981 18118
rect 1947 18004 1981 18044
rect 1947 17930 1981 17970
rect 1947 17856 1981 17896
rect 2183 19695 2217 19734
rect 2183 19622 2217 19661
rect 2183 19549 2217 19588
rect 2183 19476 2217 19515
rect 2183 19403 2217 19442
rect 2183 19330 2217 19369
rect 2183 19257 2217 19296
rect 2183 19184 2217 19223
rect 2183 19111 2217 19150
rect 2183 19038 2217 19077
rect 2183 18965 2217 19004
rect 2183 18892 2217 18931
rect 2183 18818 2217 18858
rect 2183 18744 2217 18784
rect 2183 18670 2217 18710
rect 2183 18596 2217 18636
rect 2183 18522 2217 18562
rect 2183 18448 2217 18488
rect 2183 18374 2217 18414
rect 2183 18300 2217 18340
rect 2183 18226 2217 18266
rect 2183 18152 2217 18192
rect 2183 18078 2217 18118
rect 2183 18004 2217 18044
rect 2183 17930 2217 17970
rect 2183 17856 2217 17896
rect 2419 19695 2453 19734
rect 2419 19622 2453 19661
rect 2419 19549 2453 19588
rect 2419 19476 2453 19515
rect 2419 19403 2453 19442
rect 2419 19330 2453 19369
rect 2419 19257 2453 19296
rect 2419 19184 2453 19223
rect 2419 19111 2453 19150
rect 2419 19038 2453 19077
rect 2419 18965 2453 19004
rect 2419 18892 2453 18931
rect 2419 18818 2453 18858
rect 2419 18744 2453 18784
rect 2419 18670 2453 18710
rect 2419 18596 2453 18636
rect 2419 18522 2453 18562
rect 2419 18448 2453 18488
rect 2419 18374 2453 18414
rect 2419 18300 2453 18340
rect 2419 18226 2453 18266
rect 2419 18152 2453 18192
rect 2419 18078 2453 18118
rect 2419 18004 2453 18044
rect 2419 17930 2453 17970
rect 2419 17856 2453 17896
rect 2655 19695 2689 19734
rect 2655 19622 2689 19661
rect 2655 19549 2689 19588
rect 2655 19476 2689 19515
rect 2655 19403 2689 19442
rect 2655 19330 2689 19369
rect 2655 19257 2689 19296
rect 2655 19184 2689 19223
rect 2655 19111 2689 19150
rect 2655 19038 2689 19077
rect 2655 18965 2689 19004
rect 2655 18892 2689 18931
rect 2655 18818 2689 18858
rect 2655 18744 2689 18784
rect 2655 18670 2689 18710
rect 2655 18596 2689 18636
rect 2655 18522 2689 18562
rect 2655 18448 2689 18488
rect 2655 18374 2689 18414
rect 2655 18300 2689 18340
rect 2655 18226 2689 18266
rect 2655 18152 2689 18192
rect 2655 18078 2689 18118
rect 2655 18004 2689 18044
rect 2655 17930 2689 17970
rect 2655 17856 2689 17896
rect 2891 19695 2925 19734
rect 2891 19622 2925 19661
rect 2891 19549 2925 19588
rect 2891 19476 2925 19515
rect 2891 19403 2925 19442
rect 2891 19330 2925 19369
rect 2891 19257 2925 19296
rect 2891 19184 2925 19223
rect 2891 19111 2925 19150
rect 2891 19038 2925 19077
rect 2891 18965 2925 19004
rect 2891 18892 2925 18931
rect 2891 18818 2925 18858
rect 2891 18744 2925 18784
rect 2891 18670 2925 18710
rect 2891 18596 2925 18636
rect 2891 18522 2925 18562
rect 2891 18448 2925 18488
rect 2891 18374 2925 18414
rect 2891 18300 2925 18340
rect 2891 18226 2925 18266
rect 2891 18152 2925 18192
rect 2891 18078 2925 18118
rect 2891 18004 2925 18044
rect 2891 17930 2925 17970
rect 2891 17856 2925 17896
rect 3023 19764 3036 19810
rect 3070 19764 3083 19810
rect 3023 19738 3083 19764
rect 3023 19696 3036 19738
rect 3070 19696 3083 19738
rect 3023 19666 3083 19696
rect 3023 19628 3036 19666
rect 3070 19628 3083 19666
rect 3023 19594 3083 19628
rect 3023 19560 3036 19594
rect 3070 19560 3083 19594
rect 3023 19526 3083 19560
rect 3023 19488 3036 19526
rect 3070 19488 3083 19526
rect 3023 19458 3083 19488
rect 3023 19416 3036 19458
rect 3070 19416 3083 19458
rect 3023 19390 3083 19416
rect 3023 19344 3036 19390
rect 3070 19344 3083 19390
rect 3023 19322 3083 19344
rect 3023 19272 3036 19322
rect 3070 19272 3083 19322
rect 3023 19254 3083 19272
rect 3023 19200 3036 19254
rect 3070 19200 3083 19254
rect 3023 19186 3083 19200
rect 3023 19128 3036 19186
rect 3070 19128 3083 19186
rect 3023 19118 3083 19128
rect 3023 19056 3036 19118
rect 3070 19056 3083 19118
rect 3023 19050 3083 19056
rect 3023 18984 3036 19050
rect 3070 18984 3083 19050
rect 3023 18982 3083 18984
rect 3023 18948 3036 18982
rect 3070 18948 3083 18982
rect 3023 18946 3083 18948
rect 3023 18880 3036 18946
rect 3070 18880 3083 18946
rect 3023 18874 3083 18880
rect 3023 18812 3036 18874
rect 3070 18812 3083 18874
rect 3023 18802 3083 18812
rect 3023 18744 3036 18802
rect 3070 18744 3083 18802
rect 3023 18730 3083 18744
rect 3023 18676 3036 18730
rect 3070 18676 3083 18730
rect 3023 18658 3083 18676
rect 3023 18608 3036 18658
rect 3070 18608 3083 18658
rect 3023 18586 3083 18608
rect 3023 18540 3036 18586
rect 3070 18540 3083 18586
rect 3023 18514 3083 18540
rect 3023 18472 3036 18514
rect 3070 18472 3083 18514
rect 3023 18442 3083 18472
rect 3023 18404 3036 18442
rect 3070 18404 3083 18442
rect 3023 18370 3083 18404
rect 3023 18336 3036 18370
rect 3070 18336 3083 18370
rect 3023 18302 3083 18336
rect 3023 18264 3036 18302
rect 3070 18264 3083 18302
rect 3023 18234 3083 18264
rect 3023 18192 3036 18234
rect 3070 18192 3083 18234
rect 3023 18166 3083 18192
rect 3023 18120 3036 18166
rect 3070 18120 3083 18166
rect 3023 18098 3083 18120
rect 3023 18048 3036 18098
rect 3070 18048 3083 18098
rect 3023 18030 3083 18048
rect 3023 17976 3036 18030
rect 3070 17976 3083 18030
rect 3023 17962 3083 17976
rect 3023 17904 3036 17962
rect 3070 17904 3083 17962
rect 3023 17894 3083 17904
rect 3023 17832 3036 17894
rect 3070 17832 3083 17894
rect 3023 17826 3083 17832
rect 373 17775 433 17805
rect 373 17737 386 17775
rect 420 17737 433 17775
rect 3023 17760 3036 17826
rect 3070 17760 3083 17826
rect 3023 17758 3083 17760
rect 373 17703 433 17737
rect 576 17720 592 17754
rect 659 17720 662 17754
rect 696 17720 700 17754
rect 766 17720 775 17754
rect 836 17720 850 17754
rect 906 17720 925 17754
rect 976 17720 1000 17754
rect 1046 17720 1075 17754
rect 1116 17720 1150 17754
rect 1186 17720 1222 17754
rect 1259 17720 1292 17754
rect 1334 17720 1362 17754
rect 1409 17720 1432 17754
rect 1484 17720 1502 17754
rect 1559 17720 1572 17754
rect 1634 17720 1642 17754
rect 1708 17720 1712 17754
rect 1746 17720 1748 17754
rect 1816 17720 1822 17754
rect 1886 17720 1896 17754
rect 1956 17720 1970 17754
rect 2026 17720 2044 17754
rect 2096 17720 2118 17754
rect 2166 17720 2192 17754
rect 2236 17720 2266 17754
rect 2306 17720 2340 17754
rect 2376 17720 2412 17754
rect 2448 17720 2482 17754
rect 2522 17720 2552 17754
rect 2596 17720 2622 17754
rect 2670 17720 2692 17754
rect 2744 17720 2761 17754
rect 2818 17720 2830 17754
rect 2864 17720 2880 17754
rect 3023 17724 3036 17758
rect 3070 17724 3083 17758
rect 3023 17722 3083 17724
rect 373 17669 386 17703
rect 420 17669 433 17703
rect 373 17635 433 17669
rect 3023 17656 3036 17722
rect 3070 17656 3083 17722
rect 373 17597 386 17635
rect 420 17597 433 17635
rect 373 17567 433 17597
rect 373 17525 386 17567
rect 420 17525 433 17567
rect 373 17499 433 17525
rect 373 17453 386 17499
rect 420 17453 433 17499
rect 373 17431 433 17453
rect 373 17381 386 17431
rect 420 17381 433 17431
rect 373 17363 433 17381
rect 373 17309 386 17363
rect 420 17309 433 17363
rect 373 17295 433 17309
rect 373 17237 386 17295
rect 420 17237 433 17295
rect 373 17227 433 17237
rect 373 17165 386 17227
rect 420 17165 433 17227
rect 373 17159 433 17165
rect 373 17093 386 17159
rect 420 17093 433 17159
rect 373 17091 433 17093
rect 373 17057 386 17091
rect 420 17057 433 17091
rect 373 17055 433 17057
rect 373 16989 386 17055
rect 420 16989 433 17055
rect 373 16983 433 16989
rect 373 16921 386 16983
rect 420 16921 433 16983
rect 373 16911 433 16921
rect 373 16853 386 16911
rect 420 16853 433 16911
rect 373 16839 433 16853
rect 373 16785 386 16839
rect 420 16785 433 16839
rect 373 16767 433 16785
rect 373 16717 386 16767
rect 420 16717 433 16767
rect 373 16695 433 16717
rect 373 16649 386 16695
rect 420 16649 433 16695
rect 373 16623 433 16649
rect 373 16581 386 16623
rect 420 16581 433 16623
rect 373 16551 433 16581
rect 373 16513 386 16551
rect 420 16513 433 16551
rect 373 16479 433 16513
rect 373 16445 386 16479
rect 420 16445 433 16479
rect 373 16411 433 16445
rect 373 16373 386 16411
rect 420 16373 433 16411
rect 373 16343 433 16373
rect 373 16301 386 16343
rect 420 16301 433 16343
rect 373 16275 433 16301
rect 373 16229 386 16275
rect 420 16229 433 16275
rect 373 16207 433 16229
rect 373 16157 386 16207
rect 420 16157 433 16207
rect 373 16139 433 16157
rect 373 16085 386 16139
rect 420 16085 433 16139
rect 373 16071 433 16085
rect 373 16013 386 16071
rect 420 16013 433 16071
rect 373 16003 433 16013
rect 373 15941 386 16003
rect 420 15941 433 16003
rect 373 15935 433 15941
rect 373 15869 386 15935
rect 420 15869 433 15935
rect 373 15867 433 15869
rect 373 15833 386 15867
rect 420 15833 433 15867
rect 373 15831 433 15833
rect 373 15765 386 15831
rect 420 15765 433 15831
rect 373 15759 433 15765
rect 373 15697 386 15759
rect 420 15697 433 15759
rect 531 17579 565 17618
rect 531 17506 565 17545
rect 531 17433 565 17472
rect 531 17360 565 17399
rect 531 17287 565 17326
rect 531 17214 565 17253
rect 531 17141 565 17180
rect 531 17068 565 17107
rect 531 16995 565 17034
rect 531 16922 565 16961
rect 531 16849 565 16888
rect 531 16776 565 16815
rect 531 16702 565 16742
rect 531 16628 565 16668
rect 531 16554 565 16594
rect 531 16480 565 16520
rect 531 16406 565 16446
rect 531 16332 565 16372
rect 531 16258 565 16298
rect 531 16184 565 16224
rect 531 16110 565 16150
rect 531 16036 565 16076
rect 531 15962 565 16002
rect 531 15888 565 15928
rect 531 15814 565 15854
rect 531 15740 565 15780
rect 767 17579 801 17618
rect 767 17506 801 17545
rect 767 17433 801 17472
rect 767 17360 801 17399
rect 767 17287 801 17326
rect 767 17214 801 17253
rect 767 17141 801 17180
rect 767 17068 801 17107
rect 767 16995 801 17034
rect 767 16922 801 16961
rect 767 16849 801 16888
rect 767 16776 801 16815
rect 767 16702 801 16742
rect 767 16628 801 16668
rect 767 16554 801 16594
rect 767 16480 801 16520
rect 767 16406 801 16446
rect 767 16332 801 16372
rect 767 16258 801 16298
rect 767 16184 801 16224
rect 767 16110 801 16150
rect 767 16036 801 16076
rect 767 15962 801 16002
rect 767 15888 801 15928
rect 767 15814 801 15854
rect 767 15740 801 15780
rect 1003 17579 1037 17618
rect 1003 17506 1037 17545
rect 1003 17433 1037 17472
rect 1003 17360 1037 17399
rect 1003 17287 1037 17326
rect 1003 17214 1037 17253
rect 1003 17141 1037 17180
rect 1003 17068 1037 17107
rect 1003 16995 1037 17034
rect 1003 16922 1037 16961
rect 1003 16849 1037 16888
rect 1003 16776 1037 16815
rect 1003 16702 1037 16742
rect 1003 16628 1037 16668
rect 1003 16554 1037 16594
rect 1003 16480 1037 16520
rect 1003 16406 1037 16446
rect 1003 16332 1037 16372
rect 1003 16258 1037 16298
rect 1003 16184 1037 16224
rect 1003 16110 1037 16150
rect 1003 16036 1037 16076
rect 1003 15962 1037 16002
rect 1003 15888 1037 15928
rect 1003 15814 1037 15854
rect 1003 15740 1037 15780
rect 1239 17579 1273 17618
rect 1239 17506 1273 17545
rect 1239 17433 1273 17472
rect 1239 17360 1273 17399
rect 1239 17287 1273 17326
rect 1239 17214 1273 17253
rect 1239 17141 1273 17180
rect 1239 17068 1273 17107
rect 1239 16995 1273 17034
rect 1239 16922 1273 16961
rect 1239 16849 1273 16888
rect 1239 16776 1273 16815
rect 1239 16702 1273 16742
rect 1239 16628 1273 16668
rect 1239 16554 1273 16594
rect 1239 16480 1273 16520
rect 1239 16406 1273 16446
rect 1239 16332 1273 16372
rect 1239 16258 1273 16298
rect 1239 16184 1273 16224
rect 1239 16110 1273 16150
rect 1239 16036 1273 16076
rect 1239 15962 1273 16002
rect 1239 15888 1273 15928
rect 1239 15814 1273 15854
rect 1239 15740 1273 15780
rect 1475 17579 1509 17618
rect 1475 17506 1509 17545
rect 1475 17433 1509 17472
rect 1475 17360 1509 17399
rect 1475 17287 1509 17326
rect 1475 17214 1509 17253
rect 1475 17141 1509 17180
rect 1475 17068 1509 17107
rect 1475 16995 1509 17034
rect 1475 16922 1509 16961
rect 1475 16849 1509 16888
rect 1475 16776 1509 16815
rect 1475 16702 1509 16742
rect 1475 16628 1509 16668
rect 1475 16554 1509 16594
rect 1475 16480 1509 16520
rect 1475 16406 1509 16446
rect 1475 16332 1509 16372
rect 1475 16258 1509 16298
rect 1475 16184 1509 16224
rect 1475 16110 1509 16150
rect 1475 16036 1509 16076
rect 1475 15962 1509 16002
rect 1475 15888 1509 15928
rect 1475 15814 1509 15854
rect 1475 15740 1509 15780
rect 1711 17579 1745 17618
rect 1711 17506 1745 17545
rect 1711 17433 1745 17472
rect 1711 17360 1745 17399
rect 1711 17287 1745 17326
rect 1711 17214 1745 17253
rect 1711 17141 1745 17180
rect 1711 17068 1745 17107
rect 1711 16995 1745 17034
rect 1711 16922 1745 16961
rect 1711 16849 1745 16888
rect 1711 16776 1745 16815
rect 1711 16702 1745 16742
rect 1711 16628 1745 16668
rect 1711 16554 1745 16594
rect 1711 16480 1745 16520
rect 1711 16406 1745 16446
rect 1711 16332 1745 16372
rect 1711 16258 1745 16298
rect 1711 16184 1745 16224
rect 1711 16110 1745 16150
rect 1711 16036 1745 16076
rect 1711 15962 1745 16002
rect 1711 15888 1745 15928
rect 1711 15814 1745 15854
rect 1711 15740 1745 15780
rect 1947 17579 1981 17618
rect 1947 17506 1981 17545
rect 1947 17433 1981 17472
rect 1947 17360 1981 17399
rect 1947 17287 1981 17326
rect 1947 17214 1981 17253
rect 1947 17141 1981 17180
rect 1947 17068 1981 17107
rect 1947 16995 1981 17034
rect 1947 16922 1981 16961
rect 1947 16849 1981 16888
rect 1947 16776 1981 16815
rect 1947 16702 1981 16742
rect 1947 16628 1981 16668
rect 1947 16554 1981 16594
rect 1947 16480 1981 16520
rect 1947 16406 1981 16446
rect 1947 16332 1981 16372
rect 1947 16258 1981 16298
rect 1947 16184 1981 16224
rect 1947 16110 1981 16150
rect 1947 16036 1981 16076
rect 1947 15962 1981 16002
rect 1947 15888 1981 15928
rect 1947 15814 1981 15854
rect 1947 15740 1981 15780
rect 2183 17579 2217 17618
rect 2183 17506 2217 17545
rect 2183 17433 2217 17472
rect 2183 17360 2217 17399
rect 2183 17287 2217 17326
rect 2183 17214 2217 17253
rect 2183 17141 2217 17180
rect 2183 17068 2217 17107
rect 2183 16995 2217 17034
rect 2183 16922 2217 16961
rect 2183 16849 2217 16888
rect 2183 16776 2217 16815
rect 2183 16702 2217 16742
rect 2183 16628 2217 16668
rect 2183 16554 2217 16594
rect 2183 16480 2217 16520
rect 2183 16406 2217 16446
rect 2183 16332 2217 16372
rect 2183 16258 2217 16298
rect 2183 16184 2217 16224
rect 2183 16110 2217 16150
rect 2183 16036 2217 16076
rect 2183 15962 2217 16002
rect 2183 15888 2217 15928
rect 2183 15814 2217 15854
rect 2183 15740 2217 15780
rect 2419 17579 2453 17618
rect 2419 17506 2453 17545
rect 2419 17433 2453 17472
rect 2419 17360 2453 17399
rect 2419 17287 2453 17326
rect 2419 17214 2453 17253
rect 2419 17141 2453 17180
rect 2419 17068 2453 17107
rect 2419 16995 2453 17034
rect 2419 16922 2453 16961
rect 2419 16849 2453 16888
rect 2419 16776 2453 16815
rect 2419 16702 2453 16742
rect 2419 16628 2453 16668
rect 2419 16554 2453 16594
rect 2419 16480 2453 16520
rect 2419 16406 2453 16446
rect 2419 16332 2453 16372
rect 2419 16258 2453 16298
rect 2419 16184 2453 16224
rect 2419 16110 2453 16150
rect 2419 16036 2453 16076
rect 2419 15962 2453 16002
rect 2419 15888 2453 15928
rect 2419 15814 2453 15854
rect 2419 15740 2453 15780
rect 2655 17579 2689 17618
rect 2655 17506 2689 17545
rect 2655 17433 2689 17472
rect 2655 17360 2689 17399
rect 2655 17287 2689 17326
rect 2655 17214 2689 17253
rect 2655 17141 2689 17180
rect 2655 17068 2689 17107
rect 2655 16995 2689 17034
rect 2655 16922 2689 16961
rect 2655 16849 2689 16888
rect 2655 16776 2689 16815
rect 2655 16702 2689 16742
rect 2655 16628 2689 16668
rect 2655 16554 2689 16594
rect 2655 16480 2689 16520
rect 2655 16406 2689 16446
rect 2655 16332 2689 16372
rect 2655 16258 2689 16298
rect 2655 16184 2689 16224
rect 2655 16110 2689 16150
rect 2655 16036 2689 16076
rect 2655 15962 2689 16002
rect 2655 15888 2689 15928
rect 2655 15814 2689 15854
rect 2655 15740 2689 15780
rect 2891 17579 2925 17618
rect 2891 17506 2925 17545
rect 2891 17433 2925 17472
rect 2891 17360 2925 17399
rect 2891 17287 2925 17326
rect 2891 17214 2925 17253
rect 2891 17141 2925 17180
rect 2891 17068 2925 17107
rect 2891 16995 2925 17034
rect 2891 16922 2925 16961
rect 2891 16849 2925 16888
rect 2891 16776 2925 16815
rect 2891 16702 2925 16742
rect 2891 16628 2925 16668
rect 2891 16554 2925 16594
rect 2891 16480 2925 16520
rect 2891 16406 2925 16446
rect 2891 16332 2925 16372
rect 2891 16258 2925 16298
rect 2891 16184 2925 16224
rect 2891 16110 2925 16150
rect 2891 16036 2925 16076
rect 2891 15962 2925 16002
rect 2891 15888 2925 15928
rect 2891 15814 2925 15854
rect 2891 15740 2925 15780
rect 3023 17650 3083 17656
rect 3023 17588 3036 17650
rect 3070 17588 3083 17650
rect 3023 17578 3083 17588
rect 3023 17520 3036 17578
rect 3070 17520 3083 17578
rect 3023 17506 3083 17520
rect 3023 17452 3036 17506
rect 3070 17452 3083 17506
rect 3023 17434 3083 17452
rect 3023 17384 3036 17434
rect 3070 17384 3083 17434
rect 3023 17362 3083 17384
rect 3023 17316 3036 17362
rect 3070 17316 3083 17362
rect 3023 17290 3083 17316
rect 3023 17248 3036 17290
rect 3070 17248 3083 17290
rect 3023 17218 3083 17248
rect 3023 17180 3036 17218
rect 3070 17180 3083 17218
rect 3023 17146 3083 17180
rect 3023 17112 3036 17146
rect 3070 17112 3083 17146
rect 3023 17078 3083 17112
rect 3023 17040 3036 17078
rect 3070 17040 3083 17078
rect 3023 17010 3083 17040
rect 3023 16968 3036 17010
rect 3070 16968 3083 17010
rect 3023 16942 3083 16968
rect 3023 16896 3036 16942
rect 3070 16896 3083 16942
rect 3023 16874 3083 16896
rect 3023 16824 3036 16874
rect 3070 16824 3083 16874
rect 3023 16806 3083 16824
rect 3023 16752 3036 16806
rect 3070 16752 3083 16806
rect 3023 16738 3083 16752
rect 3023 16680 3036 16738
rect 3070 16680 3083 16738
rect 3023 16670 3083 16680
rect 3023 16608 3036 16670
rect 3070 16608 3083 16670
rect 3023 16602 3083 16608
rect 3023 16536 3036 16602
rect 3070 16536 3083 16602
rect 3023 16534 3083 16536
rect 3023 16500 3036 16534
rect 3070 16500 3083 16534
rect 3023 16498 3083 16500
rect 3023 16432 3036 16498
rect 3070 16432 3083 16498
rect 3023 16426 3083 16432
rect 3023 16364 3036 16426
rect 3070 16364 3083 16426
rect 3023 16354 3083 16364
rect 3023 16296 3036 16354
rect 3070 16296 3083 16354
rect 3023 16282 3083 16296
rect 3023 16228 3036 16282
rect 3070 16228 3083 16282
rect 3023 16210 3083 16228
rect 3023 16160 3036 16210
rect 3070 16160 3083 16210
rect 3023 16138 3083 16160
rect 3023 16092 3036 16138
rect 3070 16092 3083 16138
rect 3023 16066 3083 16092
rect 3023 16024 3036 16066
rect 3070 16024 3083 16066
rect 3023 15994 3083 16024
rect 3023 15956 3036 15994
rect 3070 15956 3083 15994
rect 3023 15922 3083 15956
rect 3023 15888 3036 15922
rect 3070 15888 3083 15922
rect 3023 15854 3083 15888
rect 3023 15816 3036 15854
rect 3070 15816 3083 15854
rect 3023 15786 3083 15816
rect 3023 15744 3036 15786
rect 3070 15744 3083 15786
rect 3023 15718 3083 15744
rect 373 15687 433 15697
rect 373 15629 386 15687
rect 420 15629 433 15687
rect 373 15615 433 15629
rect 3023 15672 3036 15718
rect 3070 15672 3083 15718
rect 3023 15650 3083 15672
rect 373 15561 386 15615
rect 420 15561 433 15615
rect 576 15590 592 15624
rect 659 15590 662 15624
rect 696 15590 700 15624
rect 766 15590 775 15624
rect 836 15590 850 15624
rect 906 15590 925 15624
rect 976 15590 1000 15624
rect 1046 15590 1075 15624
rect 1116 15590 1150 15624
rect 1186 15590 1222 15624
rect 1259 15590 1292 15624
rect 1334 15590 1362 15624
rect 1409 15590 1432 15624
rect 1484 15590 1502 15624
rect 1559 15590 1572 15624
rect 1634 15590 1642 15624
rect 1708 15590 1712 15624
rect 1746 15590 1748 15624
rect 1816 15590 1822 15624
rect 1886 15590 1896 15624
rect 1956 15590 1970 15624
rect 2026 15590 2044 15624
rect 2096 15590 2118 15624
rect 2166 15590 2192 15624
rect 2236 15590 2266 15624
rect 2306 15590 2340 15624
rect 2376 15590 2412 15624
rect 2448 15590 2482 15624
rect 2522 15590 2552 15624
rect 2596 15590 2622 15624
rect 2670 15590 2692 15624
rect 2744 15590 2761 15624
rect 2818 15590 2830 15624
rect 2864 15590 2880 15624
rect 3023 15600 3036 15650
rect 3070 15600 3083 15650
rect 373 15543 433 15561
rect 373 15493 386 15543
rect 420 15493 433 15543
rect 3023 15582 3083 15600
rect 3023 15528 3036 15582
rect 3070 15528 3083 15582
rect 3023 15514 3083 15528
rect 373 15471 433 15493
rect 373 15425 386 15471
rect 420 15425 433 15471
rect 373 15399 433 15425
rect 373 15357 386 15399
rect 420 15357 433 15399
rect 373 15327 433 15357
rect 373 15289 386 15327
rect 420 15289 433 15327
rect 373 15255 433 15289
rect 373 15221 386 15255
rect 420 15221 433 15255
rect 373 15187 433 15221
rect 373 15149 386 15187
rect 420 15149 433 15187
rect 373 15119 433 15149
rect 373 15077 386 15119
rect 420 15077 433 15119
rect 373 15051 433 15077
rect 373 15005 386 15051
rect 420 15005 433 15051
rect 373 14983 433 15005
rect 373 14933 386 14983
rect 420 14933 433 14983
rect 373 14915 433 14933
rect 373 14861 386 14915
rect 420 14861 433 14915
rect 373 14847 433 14861
rect 373 14789 386 14847
rect 420 14789 433 14847
rect 373 14779 433 14789
rect 373 14717 386 14779
rect 420 14717 433 14779
rect 373 14711 433 14717
rect 373 14645 386 14711
rect 420 14645 433 14711
rect 373 14643 433 14645
rect 373 14609 386 14643
rect 420 14609 433 14643
rect 373 14607 433 14609
rect 373 14541 386 14607
rect 420 14541 433 14607
rect 373 14535 433 14541
rect 373 14473 386 14535
rect 420 14473 433 14535
rect 373 14463 433 14473
rect 373 14405 386 14463
rect 420 14405 433 14463
rect 373 14391 433 14405
rect 373 14337 386 14391
rect 420 14337 433 14391
rect 373 14319 433 14337
rect 373 14269 386 14319
rect 420 14269 433 14319
rect 373 14247 433 14269
rect 373 14201 386 14247
rect 420 14201 433 14247
rect 373 14175 433 14201
rect 373 14133 386 14175
rect 420 14133 433 14175
rect 373 14103 433 14133
rect 373 14065 386 14103
rect 420 14065 433 14103
rect 373 14031 433 14065
rect 373 13997 386 14031
rect 420 13997 433 14031
rect 373 13963 433 13997
rect 373 13925 386 13963
rect 420 13925 433 13963
rect 373 13895 433 13925
rect 373 13853 386 13895
rect 420 13853 433 13895
rect 373 13827 433 13853
rect 373 13781 386 13827
rect 420 13781 433 13827
rect 373 13759 433 13781
rect 373 13709 386 13759
rect 420 13709 433 13759
rect 373 13691 433 13709
rect 373 13637 386 13691
rect 420 13637 433 13691
rect 373 13623 433 13637
rect 373 13565 386 13623
rect 420 13565 433 13623
rect 373 13555 433 13565
rect 531 15435 565 15474
rect 531 15362 565 15401
rect 531 15289 565 15328
rect 531 15216 565 15255
rect 531 15143 565 15182
rect 531 15070 565 15109
rect 531 14997 565 15036
rect 531 14924 565 14963
rect 531 14851 565 14890
rect 531 14778 565 14817
rect 531 14705 565 14744
rect 531 14632 565 14671
rect 531 14558 565 14598
rect 531 14484 565 14524
rect 531 14410 565 14450
rect 531 14336 565 14376
rect 531 14262 565 14302
rect 531 14188 565 14228
rect 531 14114 565 14154
rect 531 14040 565 14080
rect 531 13966 565 14006
rect 531 13892 565 13932
rect 531 13818 565 13858
rect 531 13744 565 13784
rect 531 13670 565 13710
rect 531 13596 565 13636
rect 767 15435 801 15474
rect 767 15362 801 15401
rect 767 15289 801 15328
rect 767 15216 801 15255
rect 767 15143 801 15182
rect 767 15070 801 15109
rect 767 14997 801 15036
rect 767 14924 801 14963
rect 767 14851 801 14890
rect 767 14778 801 14817
rect 767 14705 801 14744
rect 767 14632 801 14671
rect 767 14558 801 14598
rect 767 14484 801 14524
rect 767 14410 801 14450
rect 767 14336 801 14376
rect 767 14262 801 14302
rect 767 14188 801 14228
rect 767 14114 801 14154
rect 767 14040 801 14080
rect 767 13966 801 14006
rect 767 13892 801 13932
rect 767 13818 801 13858
rect 767 13744 801 13784
rect 767 13670 801 13710
rect 767 13596 801 13636
rect 1003 15435 1037 15474
rect 1003 15362 1037 15401
rect 1003 15289 1037 15328
rect 1003 15216 1037 15255
rect 1003 15143 1037 15182
rect 1003 15070 1037 15109
rect 1003 14997 1037 15036
rect 1003 14924 1037 14963
rect 1003 14851 1037 14890
rect 1003 14778 1037 14817
rect 1003 14705 1037 14744
rect 1003 14632 1037 14671
rect 1003 14558 1037 14598
rect 1003 14484 1037 14524
rect 1003 14410 1037 14450
rect 1003 14336 1037 14376
rect 1003 14262 1037 14302
rect 1003 14188 1037 14228
rect 1003 14114 1037 14154
rect 1003 14040 1037 14080
rect 1003 13966 1037 14006
rect 1003 13892 1037 13932
rect 1003 13818 1037 13858
rect 1003 13744 1037 13784
rect 1003 13670 1037 13710
rect 1003 13596 1037 13636
rect 1239 15435 1273 15474
rect 1239 15362 1273 15401
rect 1239 15289 1273 15328
rect 1239 15216 1273 15255
rect 1239 15143 1273 15182
rect 1239 15070 1273 15109
rect 1239 14997 1273 15036
rect 1239 14924 1273 14963
rect 1239 14851 1273 14890
rect 1239 14778 1273 14817
rect 1239 14705 1273 14744
rect 1239 14632 1273 14671
rect 1239 14558 1273 14598
rect 1239 14484 1273 14524
rect 1239 14410 1273 14450
rect 1239 14336 1273 14376
rect 1239 14262 1273 14302
rect 1239 14188 1273 14228
rect 1239 14114 1273 14154
rect 1239 14040 1273 14080
rect 1239 13966 1273 14006
rect 1239 13892 1273 13932
rect 1239 13818 1273 13858
rect 1239 13744 1273 13784
rect 1239 13670 1273 13710
rect 1239 13596 1273 13636
rect 1475 15435 1509 15474
rect 1475 15362 1509 15401
rect 1475 15289 1509 15328
rect 1475 15216 1509 15255
rect 1475 15143 1509 15182
rect 1475 15070 1509 15109
rect 1475 14997 1509 15036
rect 1475 14924 1509 14963
rect 1475 14851 1509 14890
rect 1475 14778 1509 14817
rect 1475 14705 1509 14744
rect 1475 14632 1509 14671
rect 1475 14558 1509 14598
rect 1475 14484 1509 14524
rect 1475 14410 1509 14450
rect 1475 14336 1509 14376
rect 1475 14262 1509 14302
rect 1475 14188 1509 14228
rect 1475 14114 1509 14154
rect 1475 14040 1509 14080
rect 1475 13966 1509 14006
rect 1475 13892 1509 13932
rect 1475 13818 1509 13858
rect 1475 13744 1509 13784
rect 1475 13670 1509 13710
rect 1475 13596 1509 13636
rect 1711 15435 1745 15474
rect 1711 15362 1745 15401
rect 1711 15289 1745 15328
rect 1711 15216 1745 15255
rect 1711 15143 1745 15182
rect 1711 15070 1745 15109
rect 1711 14997 1745 15036
rect 1711 14924 1745 14963
rect 1711 14851 1745 14890
rect 1711 14778 1745 14817
rect 1711 14705 1745 14744
rect 1711 14632 1745 14671
rect 1711 14558 1745 14598
rect 1711 14484 1745 14524
rect 1711 14410 1745 14450
rect 1711 14336 1745 14376
rect 1711 14262 1745 14302
rect 1711 14188 1745 14228
rect 1711 14114 1745 14154
rect 1711 14040 1745 14080
rect 1711 13966 1745 14006
rect 1711 13892 1745 13932
rect 1711 13818 1745 13858
rect 1711 13744 1745 13784
rect 1711 13670 1745 13710
rect 1711 13596 1745 13636
rect 1947 15435 1981 15474
rect 1947 15362 1981 15401
rect 1947 15289 1981 15328
rect 1947 15216 1981 15255
rect 1947 15143 1981 15182
rect 1947 15070 1981 15109
rect 1947 14997 1981 15036
rect 1947 14924 1981 14963
rect 1947 14851 1981 14890
rect 1947 14778 1981 14817
rect 1947 14705 1981 14744
rect 1947 14632 1981 14671
rect 1947 14558 1981 14598
rect 1947 14484 1981 14524
rect 1947 14410 1981 14450
rect 1947 14336 1981 14376
rect 1947 14262 1981 14302
rect 1947 14188 1981 14228
rect 1947 14114 1981 14154
rect 1947 14040 1981 14080
rect 1947 13966 1981 14006
rect 1947 13892 1981 13932
rect 1947 13818 1981 13858
rect 1947 13744 1981 13784
rect 1947 13670 1981 13710
rect 1947 13596 1981 13636
rect 2183 15435 2217 15474
rect 2183 15362 2217 15401
rect 2183 15289 2217 15328
rect 2183 15216 2217 15255
rect 2183 15143 2217 15182
rect 2183 15070 2217 15109
rect 2183 14997 2217 15036
rect 2183 14924 2217 14963
rect 2183 14851 2217 14890
rect 2183 14778 2217 14817
rect 2183 14705 2217 14744
rect 2183 14632 2217 14671
rect 2183 14558 2217 14598
rect 2183 14484 2217 14524
rect 2183 14410 2217 14450
rect 2183 14336 2217 14376
rect 2183 14262 2217 14302
rect 2183 14188 2217 14228
rect 2183 14114 2217 14154
rect 2183 14040 2217 14080
rect 2183 13966 2217 14006
rect 2183 13892 2217 13932
rect 2183 13818 2217 13858
rect 2183 13744 2217 13784
rect 2183 13670 2217 13710
rect 2183 13596 2217 13636
rect 2419 15435 2453 15474
rect 2419 15362 2453 15401
rect 2419 15289 2453 15328
rect 2419 15216 2453 15255
rect 2419 15143 2453 15182
rect 2419 15070 2453 15109
rect 2419 14997 2453 15036
rect 2419 14924 2453 14963
rect 2419 14851 2453 14890
rect 2419 14778 2453 14817
rect 2419 14705 2453 14744
rect 2419 14632 2453 14671
rect 2419 14558 2453 14598
rect 2419 14484 2453 14524
rect 2419 14410 2453 14450
rect 2419 14336 2453 14376
rect 2419 14262 2453 14302
rect 2419 14188 2453 14228
rect 2419 14114 2453 14154
rect 2419 14040 2453 14080
rect 2419 13966 2453 14006
rect 2419 13892 2453 13932
rect 2419 13818 2453 13858
rect 2419 13744 2453 13784
rect 2419 13670 2453 13710
rect 2419 13596 2453 13636
rect 2655 15435 2689 15474
rect 2655 15362 2689 15401
rect 2655 15289 2689 15328
rect 2655 15216 2689 15255
rect 2655 15143 2689 15182
rect 2655 15070 2689 15109
rect 2655 14997 2689 15036
rect 2655 14924 2689 14963
rect 2655 14851 2689 14890
rect 2655 14778 2689 14817
rect 2655 14705 2689 14744
rect 2655 14632 2689 14671
rect 2655 14558 2689 14598
rect 2655 14484 2689 14524
rect 2655 14410 2689 14450
rect 2655 14336 2689 14376
rect 2655 14262 2689 14302
rect 2655 14188 2689 14228
rect 2655 14114 2689 14154
rect 2655 14040 2689 14080
rect 2655 13966 2689 14006
rect 2655 13892 2689 13932
rect 2655 13818 2689 13858
rect 2655 13744 2689 13784
rect 2655 13670 2689 13710
rect 2655 13596 2689 13636
rect 2891 15435 2925 15474
rect 2891 15362 2925 15401
rect 2891 15289 2925 15328
rect 2891 15216 2925 15255
rect 2891 15143 2925 15182
rect 2891 15070 2925 15109
rect 2891 14997 2925 15036
rect 2891 14924 2925 14963
rect 2891 14851 2925 14890
rect 2891 14778 2925 14817
rect 2891 14705 2925 14744
rect 2891 14632 2925 14671
rect 2891 14558 2925 14598
rect 2891 14484 2925 14524
rect 2891 14410 2925 14450
rect 2891 14336 2925 14376
rect 2891 14262 2925 14302
rect 2891 14188 2925 14228
rect 2891 14114 2925 14154
rect 2891 14040 2925 14080
rect 2891 13966 2925 14006
rect 2891 13892 2925 13932
rect 2891 13818 2925 13858
rect 2891 13744 2925 13784
rect 2891 13670 2925 13710
rect 2891 13596 2925 13636
rect 3023 15456 3036 15514
rect 3070 15456 3083 15514
rect 3023 15446 3083 15456
rect 3023 15384 3036 15446
rect 3070 15384 3083 15446
rect 3023 15378 3083 15384
rect 3023 15312 3036 15378
rect 3070 15312 3083 15378
rect 3023 15310 3083 15312
rect 3023 15276 3036 15310
rect 3070 15276 3083 15310
rect 3023 15274 3083 15276
rect 3023 15208 3036 15274
rect 3070 15208 3083 15274
rect 3023 15202 3083 15208
rect 3023 15140 3036 15202
rect 3070 15140 3083 15202
rect 3023 15130 3083 15140
rect 3023 15072 3036 15130
rect 3070 15072 3083 15130
rect 3023 15058 3083 15072
rect 3023 15004 3036 15058
rect 3070 15004 3083 15058
rect 3023 14986 3083 15004
rect 3023 14936 3036 14986
rect 3070 14936 3083 14986
rect 3023 14914 3083 14936
rect 3023 14868 3036 14914
rect 3070 14868 3083 14914
rect 3023 14842 3083 14868
rect 3023 14800 3036 14842
rect 3070 14800 3083 14842
rect 3023 14770 3083 14800
rect 3023 14732 3036 14770
rect 3070 14732 3083 14770
rect 3023 14698 3083 14732
rect 3023 14664 3036 14698
rect 3070 14664 3083 14698
rect 3023 14630 3083 14664
rect 3023 14592 3036 14630
rect 3070 14592 3083 14630
rect 3023 14562 3083 14592
rect 3023 14520 3036 14562
rect 3070 14520 3083 14562
rect 3023 14494 3083 14520
rect 3023 14448 3036 14494
rect 3070 14448 3083 14494
rect 3023 14426 3083 14448
rect 3023 14376 3036 14426
rect 3070 14376 3083 14426
rect 3023 14358 3083 14376
rect 3023 14304 3036 14358
rect 3070 14304 3083 14358
rect 3023 14290 3083 14304
rect 3023 14232 3036 14290
rect 3070 14232 3083 14290
rect 3023 14222 3083 14232
rect 3023 14160 3036 14222
rect 3070 14160 3083 14222
rect 3023 14154 3083 14160
rect 3023 14088 3036 14154
rect 3070 14088 3083 14154
rect 3023 14086 3083 14088
rect 3023 14052 3036 14086
rect 3070 14052 3083 14086
rect 3023 14050 3083 14052
rect 3023 13984 3036 14050
rect 3070 13984 3083 14050
rect 3023 13978 3083 13984
rect 3023 13916 3036 13978
rect 3070 13916 3083 13978
rect 3023 13906 3083 13916
rect 3023 13848 3036 13906
rect 3070 13848 3083 13906
rect 3023 13834 3083 13848
rect 3023 13780 3036 13834
rect 3070 13780 3083 13834
rect 3023 13762 3083 13780
rect 3023 13712 3036 13762
rect 3070 13712 3083 13762
rect 3023 13690 3083 13712
rect 3023 13644 3036 13690
rect 3070 13644 3083 13690
rect 3023 13618 3083 13644
rect 3023 13576 3036 13618
rect 3070 13576 3083 13618
rect 373 13493 386 13555
rect 420 13493 433 13555
rect 3023 13546 3083 13576
rect 3023 13508 3036 13546
rect 3070 13508 3083 13546
rect 373 13487 433 13493
rect 373 13421 386 13487
rect 420 13421 433 13487
rect 576 13460 592 13494
rect 659 13460 662 13494
rect 696 13460 700 13494
rect 766 13460 775 13494
rect 836 13460 850 13494
rect 906 13460 925 13494
rect 976 13460 1000 13494
rect 1046 13460 1075 13494
rect 1116 13460 1150 13494
rect 1186 13460 1222 13494
rect 1259 13460 1292 13494
rect 1334 13460 1362 13494
rect 1409 13460 1432 13494
rect 1484 13460 1502 13494
rect 1559 13460 1572 13494
rect 1634 13460 1642 13494
rect 1708 13460 1712 13494
rect 1746 13460 1748 13494
rect 1816 13460 1822 13494
rect 1886 13460 1896 13494
rect 1956 13460 1970 13494
rect 2026 13460 2044 13494
rect 2096 13460 2118 13494
rect 2166 13460 2192 13494
rect 2236 13460 2266 13494
rect 2306 13460 2340 13494
rect 2376 13460 2412 13494
rect 2448 13460 2482 13494
rect 2522 13460 2552 13494
rect 2596 13460 2622 13494
rect 2670 13460 2692 13494
rect 2744 13460 2761 13494
rect 2818 13460 2830 13494
rect 2864 13460 2880 13494
rect 3023 13474 3083 13508
rect 373 13419 433 13421
rect 373 13385 386 13419
rect 420 13385 433 13419
rect 3023 13440 3036 13474
rect 3070 13440 3083 13474
rect 3023 13406 3083 13440
rect 373 13383 433 13385
rect 373 13317 386 13383
rect 420 13317 433 13383
rect 373 13311 433 13317
rect 373 13249 386 13311
rect 420 13249 433 13311
rect 373 13239 433 13249
rect 373 13181 386 13239
rect 420 13181 433 13239
rect 373 13167 433 13181
rect 373 13113 386 13167
rect 420 13113 433 13167
rect 373 13095 433 13113
rect 373 13045 386 13095
rect 420 13045 433 13095
rect 373 13023 433 13045
rect 373 12977 386 13023
rect 420 12977 433 13023
rect 373 12951 433 12977
rect 373 12909 386 12951
rect 420 12909 433 12951
rect 373 12879 433 12909
rect 373 12841 386 12879
rect 420 12841 433 12879
rect 373 12807 433 12841
rect 373 12773 386 12807
rect 420 12773 433 12807
rect 373 12739 433 12773
rect 373 12701 386 12739
rect 420 12701 433 12739
rect 373 12671 433 12701
rect 373 12629 386 12671
rect 420 12629 433 12671
rect 373 12603 433 12629
rect 373 12557 386 12603
rect 420 12557 433 12603
rect 373 12535 433 12557
rect 373 12485 386 12535
rect 420 12485 433 12535
rect 373 12467 433 12485
rect 373 12413 386 12467
rect 420 12413 433 12467
rect 373 12399 433 12413
rect 373 12341 386 12399
rect 420 12341 433 12399
rect 373 12331 433 12341
rect 373 12269 386 12331
rect 420 12269 433 12331
rect 373 12263 433 12269
rect 373 12197 386 12263
rect 420 12197 433 12263
rect 373 12195 433 12197
rect 373 12161 386 12195
rect 420 12161 433 12195
rect 373 12159 433 12161
rect 373 12093 386 12159
rect 420 12093 433 12159
rect 373 12087 433 12093
rect 373 12025 386 12087
rect 420 12025 433 12087
rect 373 12015 433 12025
rect 373 11957 386 12015
rect 420 11957 433 12015
rect 373 11943 433 11957
rect 373 11889 386 11943
rect 420 11889 433 11943
rect 373 11871 433 11889
rect 373 11821 386 11871
rect 420 11821 433 11871
rect 373 11799 433 11821
rect 373 11753 386 11799
rect 420 11753 433 11799
rect 373 11727 433 11753
rect 373 11685 386 11727
rect 420 11685 433 11727
rect 373 11655 433 11685
rect 373 11617 386 11655
rect 420 11617 433 11655
rect 373 11583 433 11617
rect 373 11549 386 11583
rect 420 11549 433 11583
rect 373 11515 433 11549
rect 373 11477 386 11515
rect 420 11477 433 11515
rect 373 11447 433 11477
rect 373 11405 386 11447
rect 420 11405 433 11447
rect 531 13319 565 13358
rect 531 13246 565 13285
rect 531 13173 565 13212
rect 531 13100 565 13139
rect 531 13027 565 13066
rect 531 12954 565 12993
rect 531 12881 565 12920
rect 531 12808 565 12847
rect 531 12735 565 12774
rect 531 12662 565 12701
rect 531 12589 565 12628
rect 531 12516 565 12555
rect 531 12442 565 12482
rect 531 12368 565 12408
rect 531 12294 565 12334
rect 531 12220 565 12260
rect 531 12146 565 12186
rect 531 12072 565 12112
rect 531 11998 565 12038
rect 531 11924 565 11964
rect 531 11850 565 11890
rect 531 11776 565 11816
rect 531 11702 565 11742
rect 531 11628 565 11668
rect 531 11554 565 11594
rect 531 11480 565 11520
rect 767 13319 801 13358
rect 767 13246 801 13285
rect 767 13173 801 13212
rect 767 13100 801 13139
rect 767 13027 801 13066
rect 767 12954 801 12993
rect 767 12881 801 12920
rect 767 12808 801 12847
rect 767 12735 801 12774
rect 767 12662 801 12701
rect 767 12589 801 12628
rect 767 12516 801 12555
rect 767 12442 801 12482
rect 767 12368 801 12408
rect 767 12294 801 12334
rect 767 12220 801 12260
rect 767 12146 801 12186
rect 767 12072 801 12112
rect 767 11998 801 12038
rect 767 11924 801 11964
rect 767 11850 801 11890
rect 767 11776 801 11816
rect 767 11702 801 11742
rect 767 11628 801 11668
rect 767 11554 801 11594
rect 767 11480 801 11520
rect 1003 13319 1037 13358
rect 1003 13246 1037 13285
rect 1003 13173 1037 13212
rect 1003 13100 1037 13139
rect 1003 13027 1037 13066
rect 1003 12954 1037 12993
rect 1003 12881 1037 12920
rect 1003 12808 1037 12847
rect 1003 12735 1037 12774
rect 1003 12662 1037 12701
rect 1003 12589 1037 12628
rect 1003 12516 1037 12555
rect 1003 12442 1037 12482
rect 1003 12368 1037 12408
rect 1003 12294 1037 12334
rect 1003 12220 1037 12260
rect 1003 12146 1037 12186
rect 1003 12072 1037 12112
rect 1003 11998 1037 12038
rect 1003 11924 1037 11964
rect 1003 11850 1037 11890
rect 1003 11776 1037 11816
rect 1003 11702 1037 11742
rect 1003 11628 1037 11668
rect 1003 11554 1037 11594
rect 1003 11480 1037 11520
rect 1239 13319 1273 13358
rect 1239 13246 1273 13285
rect 1239 13173 1273 13212
rect 1239 13100 1273 13139
rect 1239 13027 1273 13066
rect 1239 12954 1273 12993
rect 1239 12881 1273 12920
rect 1239 12808 1273 12847
rect 1239 12735 1273 12774
rect 1239 12662 1273 12701
rect 1239 12589 1273 12628
rect 1239 12516 1273 12555
rect 1239 12442 1273 12482
rect 1239 12368 1273 12408
rect 1239 12294 1273 12334
rect 1239 12220 1273 12260
rect 1239 12146 1273 12186
rect 1239 12072 1273 12112
rect 1239 11998 1273 12038
rect 1239 11924 1273 11964
rect 1239 11850 1273 11890
rect 1239 11776 1273 11816
rect 1239 11702 1273 11742
rect 1239 11628 1273 11668
rect 1239 11554 1273 11594
rect 1239 11480 1273 11520
rect 1475 13319 1509 13358
rect 1475 13246 1509 13285
rect 1475 13173 1509 13212
rect 1475 13100 1509 13139
rect 1475 13027 1509 13066
rect 1475 12954 1509 12993
rect 1475 12881 1509 12920
rect 1475 12808 1509 12847
rect 1475 12735 1509 12774
rect 1475 12662 1509 12701
rect 1475 12589 1509 12628
rect 1475 12516 1509 12555
rect 1475 12442 1509 12482
rect 1475 12368 1509 12408
rect 1475 12294 1509 12334
rect 1475 12220 1509 12260
rect 1475 12146 1509 12186
rect 1475 12072 1509 12112
rect 1475 11998 1509 12038
rect 1475 11924 1509 11964
rect 1475 11850 1509 11890
rect 1475 11776 1509 11816
rect 1475 11702 1509 11742
rect 1475 11628 1509 11668
rect 1475 11554 1509 11594
rect 1475 11480 1509 11520
rect 1711 13319 1745 13358
rect 1711 13246 1745 13285
rect 1711 13173 1745 13212
rect 1711 13100 1745 13139
rect 1711 13027 1745 13066
rect 1711 12954 1745 12993
rect 1711 12881 1745 12920
rect 1711 12808 1745 12847
rect 1711 12735 1745 12774
rect 1711 12662 1745 12701
rect 1711 12589 1745 12628
rect 1711 12516 1745 12555
rect 1711 12442 1745 12482
rect 1711 12368 1745 12408
rect 1711 12294 1745 12334
rect 1711 12220 1745 12260
rect 1711 12146 1745 12186
rect 1711 12072 1745 12112
rect 1711 11998 1745 12038
rect 1711 11924 1745 11964
rect 1711 11850 1745 11890
rect 1711 11776 1745 11816
rect 1711 11702 1745 11742
rect 1711 11628 1745 11668
rect 1711 11554 1745 11594
rect 1711 11480 1745 11520
rect 1947 13319 1981 13358
rect 1947 13246 1981 13285
rect 1947 13173 1981 13212
rect 1947 13100 1981 13139
rect 1947 13027 1981 13066
rect 1947 12954 1981 12993
rect 1947 12881 1981 12920
rect 1947 12808 1981 12847
rect 1947 12735 1981 12774
rect 1947 12662 1981 12701
rect 1947 12589 1981 12628
rect 1947 12516 1981 12555
rect 1947 12442 1981 12482
rect 1947 12368 1981 12408
rect 1947 12294 1981 12334
rect 1947 12220 1981 12260
rect 1947 12146 1981 12186
rect 1947 12072 1981 12112
rect 1947 11998 1981 12038
rect 1947 11924 1981 11964
rect 1947 11850 1981 11890
rect 1947 11776 1981 11816
rect 1947 11702 1981 11742
rect 1947 11628 1981 11668
rect 1947 11554 1981 11594
rect 1947 11480 1981 11520
rect 2183 13319 2217 13358
rect 2183 13246 2217 13285
rect 2183 13173 2217 13212
rect 2183 13100 2217 13139
rect 2183 13027 2217 13066
rect 2183 12954 2217 12993
rect 2183 12881 2217 12920
rect 2183 12808 2217 12847
rect 2183 12735 2217 12774
rect 2183 12662 2217 12701
rect 2183 12589 2217 12628
rect 2183 12516 2217 12555
rect 2183 12442 2217 12482
rect 2183 12368 2217 12408
rect 2183 12294 2217 12334
rect 2183 12220 2217 12260
rect 2183 12146 2217 12186
rect 2183 12072 2217 12112
rect 2183 11998 2217 12038
rect 2183 11924 2217 11964
rect 2183 11850 2217 11890
rect 2183 11776 2217 11816
rect 2183 11702 2217 11742
rect 2183 11628 2217 11668
rect 2183 11554 2217 11594
rect 2183 11480 2217 11520
rect 2419 13319 2453 13358
rect 2419 13246 2453 13285
rect 2419 13173 2453 13212
rect 2419 13100 2453 13139
rect 2419 13027 2453 13066
rect 2419 12954 2453 12993
rect 2419 12881 2453 12920
rect 2419 12808 2453 12847
rect 2419 12735 2453 12774
rect 2419 12662 2453 12701
rect 2419 12589 2453 12628
rect 2419 12516 2453 12555
rect 2419 12442 2453 12482
rect 2419 12368 2453 12408
rect 2419 12294 2453 12334
rect 2419 12220 2453 12260
rect 2419 12146 2453 12186
rect 2419 12072 2453 12112
rect 2419 11998 2453 12038
rect 2419 11924 2453 11964
rect 2419 11850 2453 11890
rect 2419 11776 2453 11816
rect 2419 11702 2453 11742
rect 2419 11628 2453 11668
rect 2419 11554 2453 11594
rect 2419 11480 2453 11520
rect 2655 13319 2689 13358
rect 2655 13246 2689 13285
rect 2655 13173 2689 13212
rect 2655 13100 2689 13139
rect 2655 13027 2689 13066
rect 2655 12954 2689 12993
rect 2655 12881 2689 12920
rect 2655 12808 2689 12847
rect 2655 12735 2689 12774
rect 2655 12662 2689 12701
rect 2655 12589 2689 12628
rect 2655 12516 2689 12555
rect 2655 12442 2689 12482
rect 2655 12368 2689 12408
rect 2655 12294 2689 12334
rect 2655 12220 2689 12260
rect 2655 12146 2689 12186
rect 2655 12072 2689 12112
rect 2655 11998 2689 12038
rect 2655 11924 2689 11964
rect 2655 11850 2689 11890
rect 2655 11776 2689 11816
rect 2655 11702 2689 11742
rect 2655 11628 2689 11668
rect 2655 11554 2689 11594
rect 2655 11480 2689 11520
rect 2891 13319 2925 13358
rect 2891 13246 2925 13285
rect 2891 13173 2925 13212
rect 2891 13100 2925 13139
rect 2891 13027 2925 13066
rect 2891 12954 2925 12993
rect 2891 12881 2925 12920
rect 2891 12808 2925 12847
rect 2891 12735 2925 12774
rect 2891 12662 2925 12701
rect 2891 12589 2925 12628
rect 2891 12516 2925 12555
rect 2891 12442 2925 12482
rect 2891 12368 2925 12408
rect 2891 12294 2925 12334
rect 2891 12220 2925 12260
rect 2891 12146 2925 12186
rect 2891 12072 2925 12112
rect 2891 11998 2925 12038
rect 2891 11924 2925 11964
rect 2891 11850 2925 11890
rect 2891 11776 2925 11816
rect 2891 11702 2925 11742
rect 2891 11628 2925 11668
rect 2891 11554 2925 11594
rect 2891 11480 2925 11520
rect 3023 13368 3036 13406
rect 3070 13368 3083 13406
rect 3023 13338 3083 13368
rect 3023 13296 3036 13338
rect 3070 13296 3083 13338
rect 3023 13270 3083 13296
rect 3023 13224 3036 13270
rect 3070 13224 3083 13270
rect 3023 13202 3083 13224
rect 3023 13152 3036 13202
rect 3070 13152 3083 13202
rect 3023 13134 3083 13152
rect 3023 13080 3036 13134
rect 3070 13080 3083 13134
rect 3023 13066 3083 13080
rect 3023 13008 3036 13066
rect 3070 13008 3083 13066
rect 3023 12998 3083 13008
rect 3023 12936 3036 12998
rect 3070 12936 3083 12998
rect 3023 12930 3083 12936
rect 3023 12864 3036 12930
rect 3070 12864 3083 12930
rect 3023 12862 3083 12864
rect 3023 12828 3036 12862
rect 3070 12828 3083 12862
rect 3023 12826 3083 12828
rect 3023 12760 3036 12826
rect 3070 12760 3083 12826
rect 3023 12754 3083 12760
rect 3023 12692 3036 12754
rect 3070 12692 3083 12754
rect 3023 12682 3083 12692
rect 3023 12624 3036 12682
rect 3070 12624 3083 12682
rect 3023 12610 3083 12624
rect 3023 12556 3036 12610
rect 3070 12556 3083 12610
rect 3023 12538 3083 12556
rect 3023 12488 3036 12538
rect 3070 12488 3083 12538
rect 3023 12466 3083 12488
rect 3023 12420 3036 12466
rect 3070 12420 3083 12466
rect 3023 12394 3083 12420
rect 3023 12352 3036 12394
rect 3070 12352 3083 12394
rect 3023 12322 3083 12352
rect 3023 12284 3036 12322
rect 3070 12284 3083 12322
rect 3023 12250 3083 12284
rect 3023 12216 3036 12250
rect 3070 12216 3083 12250
rect 3023 12182 3083 12216
rect 3023 12144 3036 12182
rect 3070 12144 3083 12182
rect 3023 12114 3083 12144
rect 3023 12072 3036 12114
rect 3070 12072 3083 12114
rect 3023 12046 3083 12072
rect 3023 12000 3036 12046
rect 3070 12000 3083 12046
rect 3023 11978 3083 12000
rect 3023 11928 3036 11978
rect 3070 11928 3083 11978
rect 3023 11910 3083 11928
rect 3023 11856 3036 11910
rect 3070 11856 3083 11910
rect 3023 11842 3083 11856
rect 3023 11784 3036 11842
rect 3070 11784 3083 11842
rect 3023 11774 3083 11784
rect 3023 11712 3036 11774
rect 3070 11712 3083 11774
rect 3023 11706 3083 11712
rect 3023 11640 3036 11706
rect 3070 11640 3083 11706
rect 3023 11638 3083 11640
rect 3023 11604 3036 11638
rect 3070 11604 3083 11638
rect 3023 11602 3083 11604
rect 3023 11536 3036 11602
rect 3070 11536 3083 11602
rect 3023 11530 3083 11536
rect 3023 11468 3036 11530
rect 3070 11468 3083 11530
rect 3023 11458 3083 11468
rect 373 11379 433 11405
rect 373 11333 386 11379
rect 420 11333 433 11379
rect 3023 11400 3036 11458
rect 3070 11400 3083 11458
rect 3023 11386 3083 11400
rect 373 11311 433 11333
rect 576 11330 592 11364
rect 659 11330 662 11364
rect 696 11330 700 11364
rect 766 11330 775 11364
rect 836 11330 850 11364
rect 906 11330 925 11364
rect 976 11330 1000 11364
rect 1046 11330 1075 11364
rect 1116 11330 1150 11364
rect 1186 11330 1222 11364
rect 1259 11330 1292 11364
rect 1334 11330 1362 11364
rect 1409 11330 1432 11364
rect 1484 11330 1502 11364
rect 1559 11330 1572 11364
rect 1634 11330 1642 11364
rect 1708 11330 1712 11364
rect 1746 11330 1748 11364
rect 1816 11330 1822 11364
rect 1886 11330 1896 11364
rect 1956 11330 1970 11364
rect 2026 11330 2044 11364
rect 2096 11330 2118 11364
rect 2166 11330 2192 11364
rect 2236 11330 2266 11364
rect 2306 11330 2340 11364
rect 2376 11330 2412 11364
rect 2448 11330 2482 11364
rect 2522 11330 2552 11364
rect 2596 11330 2622 11364
rect 2670 11330 2692 11364
rect 2744 11330 2761 11364
rect 2818 11330 2830 11364
rect 2864 11330 2880 11364
rect 3023 11332 3036 11386
rect 3070 11332 3083 11386
rect 373 11261 386 11311
rect 420 11261 433 11311
rect 373 11243 433 11261
rect 3023 11314 3083 11332
rect 3023 11264 3036 11314
rect 3070 11264 3083 11314
rect 373 11189 386 11243
rect 420 11189 433 11243
rect 373 11175 433 11189
rect 373 11117 386 11175
rect 420 11117 433 11175
rect 373 11107 433 11117
rect 373 11045 386 11107
rect 420 11045 433 11107
rect 373 11039 433 11045
rect 373 10973 386 11039
rect 420 10973 433 11039
rect 373 10971 433 10973
rect 373 10937 386 10971
rect 420 10937 433 10971
rect 373 10935 433 10937
rect 373 10869 386 10935
rect 420 10869 433 10935
rect 373 10863 433 10869
rect 373 10801 386 10863
rect 420 10801 433 10863
rect 373 10791 433 10801
rect 373 10733 386 10791
rect 420 10733 433 10791
rect 373 10719 433 10733
rect 373 10665 386 10719
rect 420 10665 433 10719
rect 373 10647 433 10665
rect 373 10597 386 10647
rect 420 10597 433 10647
rect 373 10575 433 10597
rect 373 10529 386 10575
rect 420 10529 433 10575
rect 373 10503 433 10529
rect 373 10461 386 10503
rect 420 10461 433 10503
rect 373 10431 433 10461
rect 373 10393 386 10431
rect 420 10393 433 10431
rect 373 10359 433 10393
rect 373 10325 386 10359
rect 420 10325 433 10359
rect 373 10291 433 10325
rect 373 10253 386 10291
rect 420 10253 433 10291
rect 373 10223 433 10253
rect 373 10181 386 10223
rect 420 10181 433 10223
rect 373 10155 433 10181
rect 373 10109 386 10155
rect 420 10109 433 10155
rect 373 10087 433 10109
rect 373 10037 386 10087
rect 420 10037 433 10087
rect 373 10019 433 10037
rect 373 9965 386 10019
rect 420 9965 433 10019
rect 373 9951 433 9965
rect 373 9893 386 9951
rect 420 9893 433 9951
rect 373 9883 433 9893
rect 373 9821 386 9883
rect 420 9821 433 9883
rect 373 9815 433 9821
rect 373 9749 386 9815
rect 420 9749 433 9815
rect 373 9747 433 9749
rect 373 9713 386 9747
rect 420 9713 433 9747
rect 373 9711 433 9713
rect 373 9645 386 9711
rect 420 9645 433 9711
rect 373 9639 433 9645
rect 373 9577 386 9639
rect 420 9577 433 9639
rect 373 9567 433 9577
rect 373 9509 386 9567
rect 420 9509 433 9567
rect 373 9495 433 9509
rect 373 9441 386 9495
rect 420 9441 433 9495
rect 373 9423 433 9441
rect 373 9373 386 9423
rect 420 9373 433 9423
rect 373 9351 433 9373
rect 373 9305 386 9351
rect 420 9305 433 9351
rect 373 9279 433 9305
rect 531 11175 565 11214
rect 531 11102 565 11141
rect 531 11029 565 11068
rect 531 10956 565 10995
rect 531 10883 565 10922
rect 531 10810 565 10849
rect 531 10737 565 10776
rect 531 10664 565 10703
rect 531 10591 565 10630
rect 531 10518 565 10557
rect 531 10445 565 10484
rect 531 10372 565 10411
rect 531 10298 565 10338
rect 531 10224 565 10264
rect 531 10150 565 10190
rect 531 10076 565 10116
rect 531 10002 565 10042
rect 531 9928 565 9968
rect 531 9854 565 9894
rect 531 9780 565 9820
rect 531 9706 565 9746
rect 531 9632 565 9672
rect 531 9558 565 9598
rect 531 9484 565 9524
rect 531 9410 565 9450
rect 531 9336 565 9376
rect 767 11175 801 11214
rect 767 11102 801 11141
rect 767 11029 801 11068
rect 767 10956 801 10995
rect 767 10883 801 10922
rect 767 10810 801 10849
rect 767 10737 801 10776
rect 767 10664 801 10703
rect 767 10591 801 10630
rect 767 10518 801 10557
rect 767 10445 801 10484
rect 767 10372 801 10411
rect 767 10298 801 10338
rect 767 10224 801 10264
rect 767 10150 801 10190
rect 767 10076 801 10116
rect 767 10002 801 10042
rect 767 9928 801 9968
rect 767 9854 801 9894
rect 767 9780 801 9820
rect 767 9706 801 9746
rect 767 9632 801 9672
rect 767 9558 801 9598
rect 767 9484 801 9524
rect 767 9410 801 9450
rect 767 9336 801 9376
rect 1003 11175 1037 11214
rect 1003 11102 1037 11141
rect 1003 11029 1037 11068
rect 1003 10956 1037 10995
rect 1003 10883 1037 10922
rect 1003 10810 1037 10849
rect 1003 10737 1037 10776
rect 1003 10664 1037 10703
rect 1003 10591 1037 10630
rect 1003 10518 1037 10557
rect 1003 10445 1037 10484
rect 1003 10372 1037 10411
rect 1003 10298 1037 10338
rect 1003 10224 1037 10264
rect 1003 10150 1037 10190
rect 1003 10076 1037 10116
rect 1003 10002 1037 10042
rect 1003 9928 1037 9968
rect 1003 9854 1037 9894
rect 1003 9780 1037 9820
rect 1003 9706 1037 9746
rect 1003 9632 1037 9672
rect 1003 9558 1037 9598
rect 1003 9484 1037 9524
rect 1003 9410 1037 9450
rect 1003 9336 1037 9376
rect 1239 11175 1273 11214
rect 1239 11102 1273 11141
rect 1239 11029 1273 11068
rect 1239 10956 1273 10995
rect 1239 10883 1273 10922
rect 1239 10810 1273 10849
rect 1239 10737 1273 10776
rect 1239 10664 1273 10703
rect 1239 10591 1273 10630
rect 1239 10518 1273 10557
rect 1239 10445 1273 10484
rect 1239 10372 1273 10411
rect 1239 10298 1273 10338
rect 1239 10224 1273 10264
rect 1239 10150 1273 10190
rect 1239 10076 1273 10116
rect 1239 10002 1273 10042
rect 1239 9928 1273 9968
rect 1239 9854 1273 9894
rect 1239 9780 1273 9820
rect 1239 9706 1273 9746
rect 1239 9632 1273 9672
rect 1239 9558 1273 9598
rect 1239 9484 1273 9524
rect 1239 9410 1273 9450
rect 1239 9336 1273 9376
rect 1475 11175 1509 11214
rect 1475 11102 1509 11141
rect 1475 11029 1509 11068
rect 1475 10956 1509 10995
rect 1475 10883 1509 10922
rect 1475 10810 1509 10849
rect 1475 10737 1509 10776
rect 1475 10664 1509 10703
rect 1475 10591 1509 10630
rect 1475 10518 1509 10557
rect 1475 10445 1509 10484
rect 1475 10372 1509 10411
rect 1475 10298 1509 10338
rect 1475 10224 1509 10264
rect 1475 10150 1509 10190
rect 1475 10076 1509 10116
rect 1475 10002 1509 10042
rect 1475 9928 1509 9968
rect 1475 9854 1509 9894
rect 1475 9780 1509 9820
rect 1475 9706 1509 9746
rect 1475 9632 1509 9672
rect 1475 9558 1509 9598
rect 1475 9484 1509 9524
rect 1475 9410 1509 9450
rect 1475 9336 1509 9376
rect 1711 11175 1745 11214
rect 1711 11102 1745 11141
rect 1711 11029 1745 11068
rect 1711 10956 1745 10995
rect 1711 10883 1745 10922
rect 1711 10810 1745 10849
rect 1711 10737 1745 10776
rect 1711 10664 1745 10703
rect 1711 10591 1745 10630
rect 1711 10518 1745 10557
rect 1711 10445 1745 10484
rect 1711 10372 1745 10411
rect 1711 10298 1745 10338
rect 1711 10224 1745 10264
rect 1711 10150 1745 10190
rect 1711 10076 1745 10116
rect 1711 10002 1745 10042
rect 1711 9928 1745 9968
rect 1711 9854 1745 9894
rect 1711 9780 1745 9820
rect 1711 9706 1745 9746
rect 1711 9632 1745 9672
rect 1711 9558 1745 9598
rect 1711 9484 1745 9524
rect 1711 9410 1745 9450
rect 1711 9336 1745 9376
rect 1947 11175 1981 11214
rect 1947 11102 1981 11141
rect 1947 11029 1981 11068
rect 1947 10956 1981 10995
rect 1947 10883 1981 10922
rect 1947 10810 1981 10849
rect 1947 10737 1981 10776
rect 1947 10664 1981 10703
rect 1947 10591 1981 10630
rect 1947 10518 1981 10557
rect 1947 10445 1981 10484
rect 1947 10372 1981 10411
rect 1947 10298 1981 10338
rect 1947 10224 1981 10264
rect 1947 10150 1981 10190
rect 1947 10076 1981 10116
rect 1947 10002 1981 10042
rect 1947 9928 1981 9968
rect 1947 9854 1981 9894
rect 1947 9780 1981 9820
rect 1947 9706 1981 9746
rect 1947 9632 1981 9672
rect 1947 9558 1981 9598
rect 1947 9484 1981 9524
rect 1947 9410 1981 9450
rect 1947 9336 1981 9376
rect 2183 11175 2217 11214
rect 2183 11102 2217 11141
rect 2183 11029 2217 11068
rect 2183 10956 2217 10995
rect 2183 10883 2217 10922
rect 2183 10810 2217 10849
rect 2183 10737 2217 10776
rect 2183 10664 2217 10703
rect 2183 10591 2217 10630
rect 2183 10518 2217 10557
rect 2183 10445 2217 10484
rect 2183 10372 2217 10411
rect 2183 10298 2217 10338
rect 2183 10224 2217 10264
rect 2183 10150 2217 10190
rect 2183 10076 2217 10116
rect 2183 10002 2217 10042
rect 2183 9928 2217 9968
rect 2183 9854 2217 9894
rect 2183 9780 2217 9820
rect 2183 9706 2217 9746
rect 2183 9632 2217 9672
rect 2183 9558 2217 9598
rect 2183 9484 2217 9524
rect 2183 9410 2217 9450
rect 2183 9336 2217 9376
rect 2419 11175 2453 11214
rect 2419 11102 2453 11141
rect 2419 11029 2453 11068
rect 2419 10956 2453 10995
rect 2419 10883 2453 10922
rect 2419 10810 2453 10849
rect 2419 10737 2453 10776
rect 2419 10664 2453 10703
rect 2419 10591 2453 10630
rect 2419 10518 2453 10557
rect 2419 10445 2453 10484
rect 2419 10372 2453 10411
rect 2419 10298 2453 10338
rect 2419 10224 2453 10264
rect 2419 10150 2453 10190
rect 2419 10076 2453 10116
rect 2419 10002 2453 10042
rect 2419 9928 2453 9968
rect 2419 9854 2453 9894
rect 2419 9780 2453 9820
rect 2419 9706 2453 9746
rect 2419 9632 2453 9672
rect 2419 9558 2453 9598
rect 2419 9484 2453 9524
rect 2419 9410 2453 9450
rect 2419 9336 2453 9376
rect 2655 11175 2689 11214
rect 2655 11102 2689 11141
rect 2655 11029 2689 11068
rect 2655 10956 2689 10995
rect 2655 10883 2689 10922
rect 2655 10810 2689 10849
rect 2655 10737 2689 10776
rect 2655 10664 2689 10703
rect 2655 10591 2689 10630
rect 2655 10518 2689 10557
rect 2655 10445 2689 10484
rect 2655 10372 2689 10411
rect 2655 10298 2689 10338
rect 2655 10224 2689 10264
rect 2655 10150 2689 10190
rect 2655 10076 2689 10116
rect 2655 10002 2689 10042
rect 2655 9928 2689 9968
rect 2655 9854 2689 9894
rect 2655 9780 2689 9820
rect 2655 9706 2689 9746
rect 2655 9632 2689 9672
rect 2655 9558 2689 9598
rect 2655 9484 2689 9524
rect 2655 9410 2689 9450
rect 2655 9336 2689 9376
rect 2891 11175 2925 11214
rect 2891 11102 2925 11141
rect 2891 11029 2925 11068
rect 2891 10956 2925 10995
rect 2891 10883 2925 10922
rect 2891 10810 2925 10849
rect 2891 10737 2925 10776
rect 2891 10664 2925 10703
rect 2891 10591 2925 10630
rect 2891 10518 2925 10557
rect 2891 10445 2925 10484
rect 2891 10372 2925 10411
rect 2891 10298 2925 10338
rect 2891 10224 2925 10264
rect 2891 10150 2925 10190
rect 2891 10076 2925 10116
rect 2891 10002 2925 10042
rect 2891 9928 2925 9968
rect 2891 9854 2925 9894
rect 2891 9780 2925 9820
rect 2891 9706 2925 9746
rect 2891 9632 2925 9672
rect 2891 9558 2925 9598
rect 2891 9484 2925 9524
rect 2891 9410 2925 9450
rect 2891 9336 2925 9376
rect 3023 11242 3083 11264
rect 3023 11196 3036 11242
rect 3070 11196 3083 11242
rect 3023 11170 3083 11196
rect 3023 11128 3036 11170
rect 3070 11128 3083 11170
rect 3023 11098 3083 11128
rect 3023 11060 3036 11098
rect 3070 11060 3083 11098
rect 3023 11026 3083 11060
rect 3023 10992 3036 11026
rect 3070 10992 3083 11026
rect 3023 10958 3083 10992
rect 3023 10920 3036 10958
rect 3070 10920 3083 10958
rect 3023 10890 3083 10920
rect 3023 10848 3036 10890
rect 3070 10848 3083 10890
rect 3023 10822 3083 10848
rect 3023 10776 3036 10822
rect 3070 10776 3083 10822
rect 3023 10754 3083 10776
rect 3023 10704 3036 10754
rect 3070 10704 3083 10754
rect 3023 10686 3083 10704
rect 3023 10632 3036 10686
rect 3070 10632 3083 10686
rect 3023 10618 3083 10632
rect 3023 10560 3036 10618
rect 3070 10560 3083 10618
rect 3023 10550 3083 10560
rect 3023 10488 3036 10550
rect 3070 10488 3083 10550
rect 3023 10482 3083 10488
rect 3023 10416 3036 10482
rect 3070 10416 3083 10482
rect 3023 10414 3083 10416
rect 3023 10380 3036 10414
rect 3070 10380 3083 10414
rect 3023 10378 3083 10380
rect 3023 10312 3036 10378
rect 3070 10312 3083 10378
rect 3023 10306 3083 10312
rect 3023 10244 3036 10306
rect 3070 10244 3083 10306
rect 3023 10234 3083 10244
rect 3023 10176 3036 10234
rect 3070 10176 3083 10234
rect 3023 10162 3083 10176
rect 3023 10108 3036 10162
rect 3070 10108 3083 10162
rect 3023 10090 3083 10108
rect 3023 10040 3036 10090
rect 3070 10040 3083 10090
rect 3023 10018 3083 10040
rect 3023 9972 3036 10018
rect 3070 9972 3083 10018
rect 3023 9946 3083 9972
rect 3023 9904 3036 9946
rect 3070 9904 3083 9946
rect 3023 9874 3083 9904
rect 3023 9836 3036 9874
rect 3070 9836 3083 9874
rect 3023 9802 3083 9836
rect 3023 9768 3036 9802
rect 3070 9768 3083 9802
rect 3023 9734 3083 9768
rect 3023 9696 3036 9734
rect 3070 9696 3083 9734
rect 3023 9666 3083 9696
rect 3023 9624 3036 9666
rect 3070 9624 3083 9666
rect 3023 9598 3083 9624
rect 3023 9552 3036 9598
rect 3070 9552 3083 9598
rect 3023 9530 3083 9552
rect 3023 9480 3036 9530
rect 3070 9480 3083 9530
rect 3023 9462 3083 9480
rect 3023 9408 3036 9462
rect 3070 9408 3083 9462
rect 3023 9394 3083 9408
rect 3023 9336 3036 9394
rect 3070 9336 3083 9394
rect 3023 9326 3083 9336
rect 373 9237 386 9279
rect 420 9237 433 9279
rect 373 9207 433 9237
rect 3023 9264 3036 9326
rect 3070 9264 3083 9326
rect 3023 9258 3083 9264
rect 373 9169 386 9207
rect 420 9169 433 9207
rect 576 9200 592 9234
rect 659 9200 662 9234
rect 696 9200 700 9234
rect 766 9200 775 9234
rect 836 9200 850 9234
rect 906 9200 925 9234
rect 976 9200 1000 9234
rect 1046 9200 1075 9234
rect 1116 9200 1150 9234
rect 1186 9200 1222 9234
rect 1259 9200 1292 9234
rect 1334 9200 1362 9234
rect 1409 9200 1432 9234
rect 1484 9200 1502 9234
rect 1559 9200 1572 9234
rect 1634 9200 1642 9234
rect 1708 9200 1712 9234
rect 1746 9200 1748 9234
rect 1816 9200 1822 9234
rect 1886 9200 1896 9234
rect 1956 9200 1970 9234
rect 2026 9200 2044 9234
rect 2096 9200 2118 9234
rect 2166 9200 2192 9234
rect 2236 9200 2266 9234
rect 2306 9200 2340 9234
rect 2376 9200 2412 9234
rect 2448 9200 2482 9234
rect 2522 9200 2552 9234
rect 2596 9200 2622 9234
rect 2670 9200 2692 9234
rect 2744 9200 2761 9234
rect 2818 9200 2830 9234
rect 2864 9200 2880 9234
rect 373 9135 433 9169
rect 373 9101 386 9135
rect 420 9101 433 9135
rect 3023 9192 3036 9258
rect 3070 9192 3083 9258
rect 3023 9190 3083 9192
rect 3023 9156 3036 9190
rect 3070 9156 3083 9190
rect 3023 9154 3083 9156
rect 373 9067 433 9101
rect 373 9029 386 9067
rect 420 9029 433 9067
rect 373 8999 433 9029
rect 373 8957 386 8999
rect 420 8957 433 8999
rect 373 8931 433 8957
rect 373 8885 386 8931
rect 420 8885 433 8931
rect 373 8863 433 8885
rect 373 8813 386 8863
rect 420 8813 433 8863
rect 373 8795 433 8813
rect 373 8741 386 8795
rect 420 8741 433 8795
rect 373 8727 433 8741
rect 373 8669 386 8727
rect 420 8669 433 8727
rect 373 8659 433 8669
rect 373 8597 386 8659
rect 420 8597 433 8659
rect 373 8591 433 8597
rect 373 8525 386 8591
rect 420 8525 433 8591
rect 373 8523 433 8525
rect 373 8489 386 8523
rect 420 8489 433 8523
rect 373 8487 433 8489
rect 373 8421 386 8487
rect 420 8421 433 8487
rect 373 8415 433 8421
rect 373 8353 386 8415
rect 420 8353 433 8415
rect 373 8343 433 8353
rect 373 8285 386 8343
rect 420 8285 433 8343
rect 373 8271 433 8285
rect 373 8217 386 8271
rect 420 8217 433 8271
rect 373 8199 433 8217
rect 373 8149 386 8199
rect 420 8149 433 8199
rect 373 8127 433 8149
rect 373 8081 386 8127
rect 420 8081 433 8127
rect 373 8055 433 8081
rect 373 8013 386 8055
rect 420 8013 433 8055
rect 373 7983 433 8013
rect 373 7945 386 7983
rect 420 7945 433 7983
rect 373 7911 433 7945
rect 373 7877 386 7911
rect 420 7877 433 7911
rect 373 7843 433 7877
rect 373 7805 386 7843
rect 420 7805 433 7843
rect 373 7775 433 7805
rect 373 7733 386 7775
rect 420 7733 433 7775
rect 373 7707 433 7733
rect 373 7661 386 7707
rect 420 7661 433 7707
rect 373 7639 433 7661
rect 373 7589 386 7639
rect 420 7589 433 7639
rect 373 7571 433 7589
rect 373 7517 386 7571
rect 420 7517 433 7571
rect 373 7503 433 7517
rect 373 7445 386 7503
rect 420 7445 433 7503
rect 373 7435 433 7445
rect 373 7373 386 7435
rect 420 7373 433 7435
rect 373 7367 433 7373
rect 373 7301 386 7367
rect 420 7301 433 7367
rect 373 7299 433 7301
rect 373 7265 386 7299
rect 420 7265 433 7299
rect 373 7263 433 7265
rect 373 7197 386 7263
rect 420 7197 433 7263
rect 373 7191 433 7197
rect 373 7129 386 7191
rect 420 7129 433 7191
rect 531 9059 565 9098
rect 531 8986 565 9025
rect 531 8913 565 8952
rect 531 8840 565 8879
rect 531 8767 565 8806
rect 531 8694 565 8733
rect 531 8621 565 8660
rect 531 8548 565 8587
rect 531 8475 565 8514
rect 531 8402 565 8441
rect 531 8329 565 8368
rect 531 8256 565 8295
rect 531 8182 565 8222
rect 531 8108 565 8148
rect 531 8034 565 8074
rect 531 7960 565 8000
rect 531 7886 565 7926
rect 531 7812 565 7852
rect 531 7738 565 7778
rect 531 7664 565 7704
rect 531 7590 565 7630
rect 531 7516 565 7556
rect 531 7442 565 7482
rect 531 7368 565 7408
rect 531 7294 565 7334
rect 531 7220 565 7260
rect 767 9059 801 9098
rect 767 8986 801 9025
rect 767 8913 801 8952
rect 767 8840 801 8879
rect 767 8767 801 8806
rect 767 8694 801 8733
rect 767 8621 801 8660
rect 767 8548 801 8587
rect 767 8475 801 8514
rect 767 8402 801 8441
rect 767 8329 801 8368
rect 767 8256 801 8295
rect 767 8182 801 8222
rect 767 8108 801 8148
rect 767 8034 801 8074
rect 767 7960 801 8000
rect 767 7886 801 7926
rect 767 7812 801 7852
rect 767 7738 801 7778
rect 767 7664 801 7704
rect 767 7590 801 7630
rect 767 7516 801 7556
rect 767 7442 801 7482
rect 767 7368 801 7408
rect 767 7294 801 7334
rect 767 7220 801 7260
rect 1003 9059 1037 9098
rect 1003 8986 1037 9025
rect 1003 8913 1037 8952
rect 1003 8840 1037 8879
rect 1003 8767 1037 8806
rect 1003 8694 1037 8733
rect 1003 8621 1037 8660
rect 1003 8548 1037 8587
rect 1003 8475 1037 8514
rect 1003 8402 1037 8441
rect 1003 8329 1037 8368
rect 1003 8256 1037 8295
rect 1003 8182 1037 8222
rect 1003 8108 1037 8148
rect 1003 8034 1037 8074
rect 1003 7960 1037 8000
rect 1003 7886 1037 7926
rect 1003 7812 1037 7852
rect 1003 7738 1037 7778
rect 1003 7664 1037 7704
rect 1003 7590 1037 7630
rect 1003 7516 1037 7556
rect 1003 7442 1037 7482
rect 1003 7368 1037 7408
rect 1003 7294 1037 7334
rect 1003 7220 1037 7260
rect 1239 9059 1273 9098
rect 1239 8986 1273 9025
rect 1239 8913 1273 8952
rect 1239 8840 1273 8879
rect 1239 8767 1273 8806
rect 1239 8694 1273 8733
rect 1239 8621 1273 8660
rect 1239 8548 1273 8587
rect 1239 8475 1273 8514
rect 1239 8402 1273 8441
rect 1239 8329 1273 8368
rect 1239 8256 1273 8295
rect 1239 8182 1273 8222
rect 1239 8108 1273 8148
rect 1239 8034 1273 8074
rect 1239 7960 1273 8000
rect 1239 7886 1273 7926
rect 1239 7812 1273 7852
rect 1239 7738 1273 7778
rect 1239 7664 1273 7704
rect 1239 7590 1273 7630
rect 1239 7516 1273 7556
rect 1239 7442 1273 7482
rect 1239 7368 1273 7408
rect 1239 7294 1273 7334
rect 1239 7220 1273 7260
rect 1475 9059 1509 9098
rect 1475 8986 1509 9025
rect 1475 8913 1509 8952
rect 1475 8840 1509 8879
rect 1475 8767 1509 8806
rect 1475 8694 1509 8733
rect 1475 8621 1509 8660
rect 1475 8548 1509 8587
rect 1475 8475 1509 8514
rect 1475 8402 1509 8441
rect 1475 8329 1509 8368
rect 1475 8256 1509 8295
rect 1475 8182 1509 8222
rect 1475 8108 1509 8148
rect 1475 8034 1509 8074
rect 1475 7960 1509 8000
rect 1475 7886 1509 7926
rect 1475 7812 1509 7852
rect 1475 7738 1509 7778
rect 1475 7664 1509 7704
rect 1475 7590 1509 7630
rect 1475 7516 1509 7556
rect 1475 7442 1509 7482
rect 1475 7368 1509 7408
rect 1475 7294 1509 7334
rect 1475 7220 1509 7260
rect 1711 9059 1745 9098
rect 1711 8986 1745 9025
rect 1711 8913 1745 8952
rect 1711 8840 1745 8879
rect 1711 8767 1745 8806
rect 1711 8694 1745 8733
rect 1711 8621 1745 8660
rect 1711 8548 1745 8587
rect 1711 8475 1745 8514
rect 1711 8402 1745 8441
rect 1711 8329 1745 8368
rect 1711 8256 1745 8295
rect 1711 8182 1745 8222
rect 1711 8108 1745 8148
rect 1711 8034 1745 8074
rect 1711 7960 1745 8000
rect 1711 7886 1745 7926
rect 1711 7812 1745 7852
rect 1711 7738 1745 7778
rect 1711 7664 1745 7704
rect 1711 7590 1745 7630
rect 1711 7516 1745 7556
rect 1711 7442 1745 7482
rect 1711 7368 1745 7408
rect 1711 7294 1745 7334
rect 1711 7220 1745 7260
rect 1947 9059 1981 9098
rect 1947 8986 1981 9025
rect 1947 8913 1981 8952
rect 1947 8840 1981 8879
rect 1947 8767 1981 8806
rect 1947 8694 1981 8733
rect 1947 8621 1981 8660
rect 1947 8548 1981 8587
rect 1947 8475 1981 8514
rect 1947 8402 1981 8441
rect 1947 8329 1981 8368
rect 1947 8256 1981 8295
rect 1947 8182 1981 8222
rect 1947 8108 1981 8148
rect 1947 8034 1981 8074
rect 1947 7960 1981 8000
rect 1947 7886 1981 7926
rect 1947 7812 1981 7852
rect 1947 7738 1981 7778
rect 1947 7664 1981 7704
rect 1947 7590 1981 7630
rect 1947 7516 1981 7556
rect 1947 7442 1981 7482
rect 1947 7368 1981 7408
rect 1947 7294 1981 7334
rect 1947 7220 1981 7260
rect 2183 9059 2217 9098
rect 2183 8986 2217 9025
rect 2183 8913 2217 8952
rect 2183 8840 2217 8879
rect 2183 8767 2217 8806
rect 2183 8694 2217 8733
rect 2183 8621 2217 8660
rect 2183 8548 2217 8587
rect 2183 8475 2217 8514
rect 2183 8402 2217 8441
rect 2183 8329 2217 8368
rect 2183 8256 2217 8295
rect 2183 8182 2217 8222
rect 2183 8108 2217 8148
rect 2183 8034 2217 8074
rect 2183 7960 2217 8000
rect 2183 7886 2217 7926
rect 2183 7812 2217 7852
rect 2183 7738 2217 7778
rect 2183 7664 2217 7704
rect 2183 7590 2217 7630
rect 2183 7516 2217 7556
rect 2183 7442 2217 7482
rect 2183 7368 2217 7408
rect 2183 7294 2217 7334
rect 2183 7220 2217 7260
rect 2419 9059 2453 9098
rect 2419 8986 2453 9025
rect 2419 8913 2453 8952
rect 2419 8840 2453 8879
rect 2419 8767 2453 8806
rect 2419 8694 2453 8733
rect 2419 8621 2453 8660
rect 2419 8548 2453 8587
rect 2419 8475 2453 8514
rect 2419 8402 2453 8441
rect 2419 8329 2453 8368
rect 2419 8256 2453 8295
rect 2419 8182 2453 8222
rect 2419 8108 2453 8148
rect 2419 8034 2453 8074
rect 2419 7960 2453 8000
rect 2419 7886 2453 7926
rect 2419 7812 2453 7852
rect 2419 7738 2453 7778
rect 2419 7664 2453 7704
rect 2419 7590 2453 7630
rect 2419 7516 2453 7556
rect 2419 7442 2453 7482
rect 2419 7368 2453 7408
rect 2419 7294 2453 7334
rect 2419 7220 2453 7260
rect 2655 9059 2689 9098
rect 2655 8986 2689 9025
rect 2655 8913 2689 8952
rect 2655 8840 2689 8879
rect 2655 8767 2689 8806
rect 2655 8694 2689 8733
rect 2655 8621 2689 8660
rect 2655 8548 2689 8587
rect 2655 8475 2689 8514
rect 2655 8402 2689 8441
rect 2655 8329 2689 8368
rect 2655 8256 2689 8295
rect 2655 8182 2689 8222
rect 2655 8108 2689 8148
rect 2655 8034 2689 8074
rect 2655 7960 2689 8000
rect 2655 7886 2689 7926
rect 2655 7812 2689 7852
rect 2655 7738 2689 7778
rect 2655 7664 2689 7704
rect 2655 7590 2689 7630
rect 2655 7516 2689 7556
rect 2655 7442 2689 7482
rect 2655 7368 2689 7408
rect 2655 7294 2689 7334
rect 2655 7220 2689 7260
rect 2891 9059 2925 9098
rect 2891 8986 2925 9025
rect 2891 8913 2925 8952
rect 2891 8840 2925 8879
rect 2891 8767 2925 8806
rect 2891 8694 2925 8733
rect 2891 8621 2925 8660
rect 2891 8548 2925 8587
rect 2891 8475 2925 8514
rect 2891 8402 2925 8441
rect 2891 8329 2925 8368
rect 2891 8256 2925 8295
rect 2891 8182 2925 8222
rect 2891 8108 2925 8148
rect 2891 8034 2925 8074
rect 2891 7960 2925 8000
rect 2891 7886 2925 7926
rect 2891 7812 2925 7852
rect 2891 7738 2925 7778
rect 2891 7664 2925 7704
rect 2891 7590 2925 7630
rect 2891 7516 2925 7556
rect 2891 7442 2925 7482
rect 2891 7368 2925 7408
rect 2891 7294 2925 7334
rect 2891 7220 2925 7260
rect 3023 9088 3036 9154
rect 3070 9088 3083 9154
rect 3023 9082 3083 9088
rect 3023 9020 3036 9082
rect 3070 9020 3083 9082
rect 3023 9010 3083 9020
rect 3023 8952 3036 9010
rect 3070 8952 3083 9010
rect 3023 8938 3083 8952
rect 3023 8884 3036 8938
rect 3070 8884 3083 8938
rect 3023 8866 3083 8884
rect 3023 8816 3036 8866
rect 3070 8816 3083 8866
rect 3023 8794 3083 8816
rect 3023 8748 3036 8794
rect 3070 8748 3083 8794
rect 3023 8722 3083 8748
rect 3023 8680 3036 8722
rect 3070 8680 3083 8722
rect 3023 8650 3083 8680
rect 3023 8612 3036 8650
rect 3070 8612 3083 8650
rect 3023 8578 3083 8612
rect 3023 8544 3036 8578
rect 3070 8544 3083 8578
rect 3023 8510 3083 8544
rect 3023 8472 3036 8510
rect 3070 8472 3083 8510
rect 3023 8442 3083 8472
rect 3023 8400 3036 8442
rect 3070 8400 3083 8442
rect 3023 8374 3083 8400
rect 3023 8328 3036 8374
rect 3070 8328 3083 8374
rect 3023 8306 3083 8328
rect 3023 8256 3036 8306
rect 3070 8256 3083 8306
rect 3023 8238 3083 8256
rect 3023 8184 3036 8238
rect 3070 8184 3083 8238
rect 3023 8170 3083 8184
rect 3023 8112 3036 8170
rect 3070 8112 3083 8170
rect 3023 8102 3083 8112
rect 3023 8040 3036 8102
rect 3070 8040 3083 8102
rect 3023 8034 3083 8040
rect 3023 7968 3036 8034
rect 3070 7968 3083 8034
rect 3023 7966 3083 7968
rect 3023 7932 3036 7966
rect 3070 7932 3083 7966
rect 3023 7930 3083 7932
rect 3023 7864 3036 7930
rect 3070 7864 3083 7930
rect 3023 7858 3083 7864
rect 3023 7796 3036 7858
rect 3070 7796 3083 7858
rect 3023 7786 3083 7796
rect 3023 7728 3036 7786
rect 3070 7728 3083 7786
rect 3023 7714 3083 7728
rect 3023 7660 3036 7714
rect 3070 7660 3083 7714
rect 3023 7642 3083 7660
rect 3023 7592 3036 7642
rect 3070 7592 3083 7642
rect 3023 7570 3083 7592
rect 3023 7524 3036 7570
rect 3070 7524 3083 7570
rect 3023 7498 3083 7524
rect 3023 7456 3036 7498
rect 3070 7456 3083 7498
rect 3023 7426 3083 7456
rect 3023 7388 3036 7426
rect 3070 7388 3083 7426
rect 3023 7354 3083 7388
rect 3023 7320 3036 7354
rect 3070 7320 3083 7354
rect 3023 7286 3083 7320
rect 3023 7248 3036 7286
rect 3070 7248 3083 7286
rect 3023 7218 3083 7248
rect 373 7119 433 7129
rect 373 7061 386 7119
rect 420 7061 433 7119
rect 3023 7176 3036 7218
rect 3070 7176 3083 7218
rect 3023 7150 3083 7176
rect 3023 7104 3036 7150
rect 3070 7104 3083 7150
rect 576 7070 592 7104
rect 659 7070 662 7104
rect 696 7070 700 7104
rect 766 7070 775 7104
rect 836 7070 850 7104
rect 906 7070 925 7104
rect 976 7070 1000 7104
rect 1046 7070 1075 7104
rect 1116 7070 1150 7104
rect 1186 7070 1222 7104
rect 1259 7070 1292 7104
rect 1334 7070 1362 7104
rect 1409 7070 1432 7104
rect 1484 7070 1502 7104
rect 1559 7070 1572 7104
rect 1634 7070 1642 7104
rect 1708 7070 1712 7104
rect 1746 7070 1748 7104
rect 1816 7070 1822 7104
rect 1886 7070 1896 7104
rect 1956 7070 1970 7104
rect 2026 7070 2044 7104
rect 2096 7070 2118 7104
rect 2166 7070 2192 7104
rect 2236 7070 2266 7104
rect 2306 7070 2340 7104
rect 2376 7070 2412 7104
rect 2448 7070 2482 7104
rect 2522 7070 2552 7104
rect 2596 7070 2622 7104
rect 2670 7070 2692 7104
rect 2744 7070 2761 7104
rect 2818 7070 2830 7104
rect 2864 7070 2880 7104
rect 3023 7082 3083 7104
rect 373 7047 433 7061
rect 373 6993 386 7047
rect 420 6993 433 7047
rect 373 6975 433 6993
rect 3023 7032 3036 7082
rect 3070 7032 3083 7082
rect 3023 7014 3083 7032
rect 373 6925 386 6975
rect 420 6925 433 6975
rect 373 6903 433 6925
rect 373 6857 386 6903
rect 420 6857 433 6903
rect 373 6831 433 6857
rect 373 6789 386 6831
rect 420 6789 433 6831
rect 373 6759 433 6789
rect 373 6721 386 6759
rect 420 6721 433 6759
rect 373 6687 433 6721
rect 373 6653 386 6687
rect 420 6653 433 6687
rect 373 6619 433 6653
rect 373 6581 386 6619
rect 420 6581 433 6619
rect 373 6551 433 6581
rect 373 6509 386 6551
rect 420 6509 433 6551
rect 373 6483 433 6509
rect 373 6437 386 6483
rect 420 6437 433 6483
rect 373 6415 433 6437
rect 373 6365 386 6415
rect 420 6365 433 6415
rect 373 6347 433 6365
rect 373 6293 386 6347
rect 420 6293 433 6347
rect 373 6279 433 6293
rect 373 6221 386 6279
rect 420 6221 433 6279
rect 373 6211 433 6221
rect 373 6149 386 6211
rect 420 6149 433 6211
rect 373 6143 433 6149
rect 373 6077 386 6143
rect 420 6077 433 6143
rect 373 6075 433 6077
rect 373 6041 386 6075
rect 420 6041 433 6075
rect 373 6039 433 6041
rect 373 5973 386 6039
rect 420 5973 433 6039
rect 373 5967 433 5973
rect 373 5905 386 5967
rect 420 5905 433 5967
rect 373 5895 433 5905
rect 373 5837 386 5895
rect 420 5837 433 5895
rect 373 5823 433 5837
rect 373 5769 386 5823
rect 420 5769 433 5823
rect 373 5751 433 5769
rect 373 5701 386 5751
rect 420 5701 433 5751
rect 373 5679 433 5701
rect 373 5633 386 5679
rect 420 5633 433 5679
rect 373 5607 433 5633
rect 373 5565 386 5607
rect 420 5565 433 5607
rect 373 5535 433 5565
rect 373 5497 386 5535
rect 420 5497 433 5535
rect 373 5463 433 5497
rect 373 5429 386 5463
rect 420 5429 433 5463
rect 373 5395 433 5429
rect 373 5357 386 5395
rect 420 5357 433 5395
rect 373 5327 433 5357
rect 373 5285 386 5327
rect 420 5285 433 5327
rect 373 5259 433 5285
rect 373 5213 386 5259
rect 420 5213 433 5259
rect 373 5191 433 5213
rect 373 5141 386 5191
rect 420 5141 433 5191
rect 373 5123 433 5141
rect 373 5069 386 5123
rect 420 5069 433 5123
rect 373 5055 433 5069
rect 373 4997 386 5055
rect 420 4997 433 5055
rect 531 6915 565 6954
rect 531 6842 565 6881
rect 531 6769 565 6808
rect 531 6696 565 6735
rect 531 6623 565 6662
rect 531 6550 565 6589
rect 531 6477 565 6516
rect 531 6404 565 6443
rect 531 6331 565 6370
rect 531 6258 565 6297
rect 531 6185 565 6224
rect 531 6112 565 6151
rect 531 6038 565 6078
rect 531 5964 565 6004
rect 531 5890 565 5930
rect 531 5816 565 5856
rect 531 5742 565 5782
rect 531 5668 565 5708
rect 531 5594 565 5634
rect 531 5520 565 5560
rect 531 5446 565 5486
rect 531 5372 565 5412
rect 531 5298 565 5338
rect 531 5224 565 5264
rect 531 5150 565 5190
rect 531 5076 565 5116
rect 767 6915 801 6954
rect 767 6842 801 6881
rect 767 6769 801 6808
rect 767 6696 801 6735
rect 767 6623 801 6662
rect 767 6550 801 6589
rect 767 6477 801 6516
rect 767 6404 801 6443
rect 767 6331 801 6370
rect 767 6258 801 6297
rect 767 6185 801 6224
rect 767 6112 801 6151
rect 767 6038 801 6078
rect 767 5964 801 6004
rect 767 5890 801 5930
rect 767 5816 801 5856
rect 767 5742 801 5782
rect 767 5668 801 5708
rect 767 5594 801 5634
rect 767 5520 801 5560
rect 767 5446 801 5486
rect 767 5372 801 5412
rect 767 5298 801 5338
rect 767 5224 801 5264
rect 767 5150 801 5190
rect 767 5076 801 5116
rect 1003 6915 1037 6954
rect 1003 6842 1037 6881
rect 1003 6769 1037 6808
rect 1003 6696 1037 6735
rect 1003 6623 1037 6662
rect 1003 6550 1037 6589
rect 1003 6477 1037 6516
rect 1003 6404 1037 6443
rect 1003 6331 1037 6370
rect 1003 6258 1037 6297
rect 1003 6185 1037 6224
rect 1003 6112 1037 6151
rect 1003 6038 1037 6078
rect 1003 5964 1037 6004
rect 1003 5890 1037 5930
rect 1003 5816 1037 5856
rect 1003 5742 1037 5782
rect 1003 5668 1037 5708
rect 1003 5594 1037 5634
rect 1003 5520 1037 5560
rect 1003 5446 1037 5486
rect 1003 5372 1037 5412
rect 1003 5298 1037 5338
rect 1003 5224 1037 5264
rect 1003 5150 1037 5190
rect 1003 5076 1037 5116
rect 1239 6915 1273 6954
rect 1239 6842 1273 6881
rect 1239 6769 1273 6808
rect 1239 6696 1273 6735
rect 1239 6623 1273 6662
rect 1239 6550 1273 6589
rect 1239 6477 1273 6516
rect 1239 6404 1273 6443
rect 1239 6331 1273 6370
rect 1239 6258 1273 6297
rect 1239 6185 1273 6224
rect 1239 6112 1273 6151
rect 1239 6038 1273 6078
rect 1239 5964 1273 6004
rect 1239 5890 1273 5930
rect 1239 5816 1273 5856
rect 1239 5742 1273 5782
rect 1239 5668 1273 5708
rect 1239 5594 1273 5634
rect 1239 5520 1273 5560
rect 1239 5446 1273 5486
rect 1239 5372 1273 5412
rect 1239 5298 1273 5338
rect 1239 5224 1273 5264
rect 1239 5150 1273 5190
rect 1239 5076 1273 5116
rect 1475 6915 1509 6954
rect 1475 6842 1509 6881
rect 1475 6769 1509 6808
rect 1475 6696 1509 6735
rect 1475 6623 1509 6662
rect 1475 6550 1509 6589
rect 1475 6477 1509 6516
rect 1475 6404 1509 6443
rect 1475 6331 1509 6370
rect 1475 6258 1509 6297
rect 1475 6185 1509 6224
rect 1475 6112 1509 6151
rect 1475 6038 1509 6078
rect 1475 5964 1509 6004
rect 1475 5890 1509 5930
rect 1475 5816 1509 5856
rect 1475 5742 1509 5782
rect 1475 5668 1509 5708
rect 1475 5594 1509 5634
rect 1475 5520 1509 5560
rect 1475 5446 1509 5486
rect 1475 5372 1509 5412
rect 1475 5298 1509 5338
rect 1475 5224 1509 5264
rect 1475 5150 1509 5190
rect 1475 5076 1509 5116
rect 1711 6915 1745 6954
rect 1711 6842 1745 6881
rect 1711 6769 1745 6808
rect 1711 6696 1745 6735
rect 1711 6623 1745 6662
rect 1711 6550 1745 6589
rect 1711 6477 1745 6516
rect 1711 6404 1745 6443
rect 1711 6331 1745 6370
rect 1711 6258 1745 6297
rect 1711 6185 1745 6224
rect 1711 6112 1745 6151
rect 1711 6038 1745 6078
rect 1711 5964 1745 6004
rect 1711 5890 1745 5930
rect 1711 5816 1745 5856
rect 1711 5742 1745 5782
rect 1711 5668 1745 5708
rect 1711 5594 1745 5634
rect 1711 5520 1745 5560
rect 1711 5446 1745 5486
rect 1711 5372 1745 5412
rect 1711 5298 1745 5338
rect 1711 5224 1745 5264
rect 1711 5150 1745 5190
rect 1711 5076 1745 5116
rect 1947 6915 1981 6954
rect 1947 6842 1981 6881
rect 1947 6769 1981 6808
rect 1947 6696 1981 6735
rect 1947 6623 1981 6662
rect 1947 6550 1981 6589
rect 1947 6477 1981 6516
rect 1947 6404 1981 6443
rect 1947 6331 1981 6370
rect 1947 6258 1981 6297
rect 1947 6185 1981 6224
rect 1947 6112 1981 6151
rect 1947 6038 1981 6078
rect 1947 5964 1981 6004
rect 1947 5890 1981 5930
rect 1947 5816 1981 5856
rect 1947 5742 1981 5782
rect 1947 5668 1981 5708
rect 1947 5594 1981 5634
rect 1947 5520 1981 5560
rect 1947 5446 1981 5486
rect 1947 5372 1981 5412
rect 1947 5298 1981 5338
rect 1947 5224 1981 5264
rect 1947 5150 1981 5190
rect 1947 5076 1981 5116
rect 2183 6915 2217 6954
rect 2183 6842 2217 6881
rect 2183 6769 2217 6808
rect 2183 6696 2217 6735
rect 2183 6623 2217 6662
rect 2183 6550 2217 6589
rect 2183 6477 2217 6516
rect 2183 6404 2217 6443
rect 2183 6331 2217 6370
rect 2183 6258 2217 6297
rect 2183 6185 2217 6224
rect 2183 6112 2217 6151
rect 2183 6038 2217 6078
rect 2183 5964 2217 6004
rect 2183 5890 2217 5930
rect 2183 5816 2217 5856
rect 2183 5742 2217 5782
rect 2183 5668 2217 5708
rect 2183 5594 2217 5634
rect 2183 5520 2217 5560
rect 2183 5446 2217 5486
rect 2183 5372 2217 5412
rect 2183 5298 2217 5338
rect 2183 5224 2217 5264
rect 2183 5150 2217 5190
rect 2183 5076 2217 5116
rect 2419 6915 2453 6954
rect 2419 6842 2453 6881
rect 2419 6769 2453 6808
rect 2419 6696 2453 6735
rect 2419 6623 2453 6662
rect 2419 6550 2453 6589
rect 2419 6477 2453 6516
rect 2419 6404 2453 6443
rect 2419 6331 2453 6370
rect 2419 6258 2453 6297
rect 2419 6185 2453 6224
rect 2419 6112 2453 6151
rect 2419 6038 2453 6078
rect 2419 5964 2453 6004
rect 2419 5890 2453 5930
rect 2419 5816 2453 5856
rect 2419 5742 2453 5782
rect 2419 5668 2453 5708
rect 2419 5594 2453 5634
rect 2419 5520 2453 5560
rect 2419 5446 2453 5486
rect 2419 5372 2453 5412
rect 2419 5298 2453 5338
rect 2419 5224 2453 5264
rect 2419 5150 2453 5190
rect 2419 5076 2453 5116
rect 2655 6915 2689 6954
rect 2655 6842 2689 6881
rect 2655 6769 2689 6808
rect 2655 6696 2689 6735
rect 2655 6623 2689 6662
rect 2655 6550 2689 6589
rect 2655 6477 2689 6516
rect 2655 6404 2689 6443
rect 2655 6331 2689 6370
rect 2655 6258 2689 6297
rect 2655 6185 2689 6224
rect 2655 6112 2689 6151
rect 2655 6038 2689 6078
rect 2655 5964 2689 6004
rect 2655 5890 2689 5930
rect 2655 5816 2689 5856
rect 2655 5742 2689 5782
rect 2655 5668 2689 5708
rect 2655 5594 2689 5634
rect 2655 5520 2689 5560
rect 2655 5446 2689 5486
rect 2655 5372 2689 5412
rect 2655 5298 2689 5338
rect 2655 5224 2689 5264
rect 2655 5150 2689 5190
rect 2655 5076 2689 5116
rect 2891 6915 2925 6954
rect 2891 6842 2925 6881
rect 2891 6769 2925 6808
rect 2891 6696 2925 6735
rect 2891 6623 2925 6662
rect 2891 6550 2925 6589
rect 2891 6477 2925 6516
rect 2891 6404 2925 6443
rect 2891 6331 2925 6370
rect 2891 6258 2925 6297
rect 2891 6185 2925 6224
rect 2891 6112 2925 6151
rect 2891 6038 2925 6078
rect 2891 5964 2925 6004
rect 2891 5890 2925 5930
rect 2891 5816 2925 5856
rect 2891 5742 2925 5782
rect 2891 5668 2925 5708
rect 2891 5594 2925 5634
rect 2891 5520 2925 5560
rect 2891 5446 2925 5486
rect 2891 5372 2925 5412
rect 2891 5298 2925 5338
rect 2891 5224 2925 5264
rect 2891 5150 2925 5190
rect 2891 5076 2925 5116
rect 3023 6960 3036 7014
rect 3070 6960 3083 7014
rect 3023 6946 3083 6960
rect 3023 6888 3036 6946
rect 3070 6888 3083 6946
rect 3023 6878 3083 6888
rect 3023 6816 3036 6878
rect 3070 6816 3083 6878
rect 3023 6810 3083 6816
rect 3023 6744 3036 6810
rect 3070 6744 3083 6810
rect 3023 6742 3083 6744
rect 3023 6708 3036 6742
rect 3070 6708 3083 6742
rect 3023 6706 3083 6708
rect 3023 6640 3036 6706
rect 3070 6640 3083 6706
rect 3023 6634 3083 6640
rect 3023 6572 3036 6634
rect 3070 6572 3083 6634
rect 3023 6562 3083 6572
rect 3023 6504 3036 6562
rect 3070 6504 3083 6562
rect 3023 6490 3083 6504
rect 3023 6436 3036 6490
rect 3070 6436 3083 6490
rect 3023 6418 3083 6436
rect 3023 6368 3036 6418
rect 3070 6368 3083 6418
rect 3023 6346 3083 6368
rect 3023 6300 3036 6346
rect 3070 6300 3083 6346
rect 3023 6274 3083 6300
rect 3023 6232 3036 6274
rect 3070 6232 3083 6274
rect 3023 6202 3083 6232
rect 3023 6164 3036 6202
rect 3070 6164 3083 6202
rect 3023 6130 3083 6164
rect 3023 6096 3036 6130
rect 3070 6096 3083 6130
rect 3023 6062 3083 6096
rect 3023 6024 3036 6062
rect 3070 6024 3083 6062
rect 3023 5994 3083 6024
rect 3023 5952 3036 5994
rect 3070 5952 3083 5994
rect 3023 5926 3083 5952
rect 3023 5880 3036 5926
rect 3070 5880 3083 5926
rect 3023 5858 3083 5880
rect 3023 5808 3036 5858
rect 3070 5808 3083 5858
rect 3023 5790 3083 5808
rect 3023 5736 3036 5790
rect 3070 5736 3083 5790
rect 3023 5722 3083 5736
rect 3023 5664 3036 5722
rect 3070 5664 3083 5722
rect 3023 5654 3083 5664
rect 3023 5592 3036 5654
rect 3070 5592 3083 5654
rect 3023 5586 3083 5592
rect 3023 5520 3036 5586
rect 3070 5520 3083 5586
rect 3023 5518 3083 5520
rect 3023 5484 3036 5518
rect 3070 5484 3083 5518
rect 3023 5482 3083 5484
rect 3023 5416 3036 5482
rect 3070 5416 3083 5482
rect 3023 5410 3083 5416
rect 3023 5348 3036 5410
rect 3070 5348 3083 5410
rect 3023 5338 3083 5348
rect 3023 5280 3036 5338
rect 3070 5280 3083 5338
rect 3023 5266 3083 5280
rect 3023 5212 3036 5266
rect 3070 5212 3083 5266
rect 3023 5194 3083 5212
rect 3023 5144 3036 5194
rect 3070 5144 3083 5194
rect 3023 5122 3083 5144
rect 3023 5076 3036 5122
rect 3070 5076 3083 5122
rect 3023 5050 3083 5076
rect 373 4987 433 4997
rect 373 4925 386 4987
rect 420 4925 433 4987
rect 3023 5008 3036 5050
rect 3070 5008 3083 5050
rect 3023 4978 3083 5008
rect 576 4940 592 4974
rect 659 4940 662 4974
rect 696 4940 700 4974
rect 766 4940 775 4974
rect 836 4940 850 4974
rect 906 4940 925 4974
rect 976 4940 1000 4974
rect 1046 4940 1075 4974
rect 1116 4940 1150 4974
rect 1186 4940 1222 4974
rect 1259 4940 1292 4974
rect 1334 4940 1362 4974
rect 1409 4940 1432 4974
rect 1484 4940 1502 4974
rect 1559 4940 1572 4974
rect 1634 4940 1642 4974
rect 1708 4940 1712 4974
rect 1746 4940 1748 4974
rect 1816 4940 1822 4974
rect 1886 4940 1896 4974
rect 1956 4940 1970 4974
rect 2026 4940 2044 4974
rect 2096 4940 2118 4974
rect 2166 4940 2192 4974
rect 2236 4940 2266 4974
rect 2306 4940 2340 4974
rect 2376 4940 2412 4974
rect 2448 4940 2482 4974
rect 2522 4940 2552 4974
rect 2596 4940 2622 4974
rect 2670 4940 2692 4974
rect 2744 4940 2761 4974
rect 2818 4940 2830 4974
rect 2864 4940 2880 4974
rect 3023 4940 3036 4978
rect 3070 4940 3083 4978
rect 373 4919 433 4925
rect 373 4853 386 4919
rect 420 4853 433 4919
rect 3023 4906 3083 4940
rect 3023 4872 3036 4906
rect 3070 4872 3083 4906
rect 373 4851 433 4853
rect 373 4817 386 4851
rect 420 4817 433 4851
rect 373 4815 433 4817
rect 373 4749 386 4815
rect 420 4749 433 4815
rect 373 4743 433 4749
rect 373 4681 386 4743
rect 420 4681 433 4743
rect 373 4671 433 4681
rect 373 4613 386 4671
rect 420 4613 433 4671
rect 373 4599 433 4613
rect 373 4545 386 4599
rect 420 4545 433 4599
rect 373 4527 433 4545
rect 373 4477 386 4527
rect 420 4477 433 4527
rect 373 4455 433 4477
rect 373 4409 386 4455
rect 420 4409 433 4455
rect 373 4383 433 4409
rect 373 4341 386 4383
rect 420 4341 433 4383
rect 373 4311 433 4341
rect 373 4273 386 4311
rect 420 4273 433 4311
rect 373 4239 433 4273
rect 373 4205 386 4239
rect 420 4205 433 4239
rect 373 4171 433 4205
rect 373 4133 386 4171
rect 420 4133 433 4171
rect 373 4103 433 4133
rect 373 4061 386 4103
rect 420 4061 433 4103
rect 373 4035 433 4061
rect 373 3989 386 4035
rect 420 3989 433 4035
rect 373 3967 433 3989
rect 373 3917 386 3967
rect 420 3917 433 3967
rect 373 3899 433 3917
rect 373 3845 386 3899
rect 420 3845 433 3899
rect 373 3831 433 3845
rect 373 3773 386 3831
rect 420 3773 433 3831
rect 373 3763 433 3773
rect 373 3701 386 3763
rect 420 3701 433 3763
rect 373 3695 433 3701
rect 373 3629 386 3695
rect 420 3629 433 3695
rect 373 3627 433 3629
rect 373 3593 386 3627
rect 420 3593 433 3627
rect 373 3591 433 3593
rect 373 3525 386 3591
rect 420 3525 433 3591
rect 373 3519 433 3525
rect 373 3457 386 3519
rect 420 3457 433 3519
rect 373 3447 433 3457
rect 373 3389 386 3447
rect 420 3389 433 3447
rect 373 3375 433 3389
rect 373 3321 386 3375
rect 420 3321 433 3375
rect 373 3303 433 3321
rect 373 3253 386 3303
rect 420 3253 433 3303
rect 373 3231 433 3253
rect 373 3185 386 3231
rect 420 3185 433 3231
rect 373 3159 433 3185
rect 373 3117 386 3159
rect 420 3117 433 3159
rect 373 3087 433 3117
rect 373 3049 386 3087
rect 420 3049 433 3087
rect 373 3015 433 3049
rect 373 2981 386 3015
rect 420 2981 433 3015
rect 373 2947 433 2981
rect 373 2909 386 2947
rect 420 2909 433 2947
rect 531 4799 565 4838
rect 531 4726 565 4765
rect 531 4653 565 4692
rect 531 4580 565 4619
rect 531 4507 565 4546
rect 531 4434 565 4473
rect 531 4361 565 4400
rect 531 4288 565 4327
rect 531 4215 565 4254
rect 531 4142 565 4181
rect 531 4069 565 4108
rect 531 3996 565 4035
rect 531 3922 565 3962
rect 531 3848 565 3888
rect 531 3774 565 3814
rect 531 3700 565 3740
rect 531 3626 565 3666
rect 531 3552 565 3592
rect 531 3478 565 3518
rect 531 3404 565 3444
rect 531 3330 565 3370
rect 531 3256 565 3296
rect 531 3182 565 3222
rect 531 3108 565 3148
rect 531 3034 565 3074
rect 531 2960 565 3000
rect 767 4799 801 4838
rect 767 4726 801 4765
rect 767 4653 801 4692
rect 767 4580 801 4619
rect 767 4507 801 4546
rect 767 4434 801 4473
rect 767 4361 801 4400
rect 767 4288 801 4327
rect 767 4215 801 4254
rect 767 4142 801 4181
rect 767 4069 801 4108
rect 767 3996 801 4035
rect 767 3922 801 3962
rect 767 3848 801 3888
rect 767 3774 801 3814
rect 767 3700 801 3740
rect 767 3626 801 3666
rect 767 3552 801 3592
rect 767 3478 801 3518
rect 767 3404 801 3444
rect 767 3330 801 3370
rect 767 3256 801 3296
rect 767 3182 801 3222
rect 767 3108 801 3148
rect 767 3034 801 3074
rect 767 2960 801 3000
rect 1003 4799 1037 4838
rect 1003 4726 1037 4765
rect 1003 4653 1037 4692
rect 1003 4580 1037 4619
rect 1003 4507 1037 4546
rect 1003 4434 1037 4473
rect 1003 4361 1037 4400
rect 1003 4288 1037 4327
rect 1003 4215 1037 4254
rect 1003 4142 1037 4181
rect 1003 4069 1037 4108
rect 1003 3996 1037 4035
rect 1003 3922 1037 3962
rect 1003 3848 1037 3888
rect 1003 3774 1037 3814
rect 1003 3700 1037 3740
rect 1003 3626 1037 3666
rect 1003 3552 1037 3592
rect 1003 3478 1037 3518
rect 1003 3404 1037 3444
rect 1003 3330 1037 3370
rect 1003 3256 1037 3296
rect 1003 3182 1037 3222
rect 1003 3108 1037 3148
rect 1003 3034 1037 3074
rect 1003 2960 1037 3000
rect 1239 4799 1273 4838
rect 1239 4726 1273 4765
rect 1239 4653 1273 4692
rect 1239 4580 1273 4619
rect 1239 4507 1273 4546
rect 1239 4434 1273 4473
rect 1239 4361 1273 4400
rect 1239 4288 1273 4327
rect 1239 4215 1273 4254
rect 1239 4142 1273 4181
rect 1239 4069 1273 4108
rect 1239 3996 1273 4035
rect 1239 3922 1273 3962
rect 1239 3848 1273 3888
rect 1239 3774 1273 3814
rect 1239 3700 1273 3740
rect 1239 3626 1273 3666
rect 1239 3552 1273 3592
rect 1239 3478 1273 3518
rect 1239 3404 1273 3444
rect 1239 3330 1273 3370
rect 1239 3256 1273 3296
rect 1239 3182 1273 3222
rect 1239 3108 1273 3148
rect 1239 3034 1273 3074
rect 1239 2960 1273 3000
rect 1475 4799 1509 4838
rect 1475 4726 1509 4765
rect 1475 4653 1509 4692
rect 1475 4580 1509 4619
rect 1475 4507 1509 4546
rect 1475 4434 1509 4473
rect 1475 4361 1509 4400
rect 1475 4288 1509 4327
rect 1475 4215 1509 4254
rect 1475 4142 1509 4181
rect 1475 4069 1509 4108
rect 1475 3996 1509 4035
rect 1475 3922 1509 3962
rect 1475 3848 1509 3888
rect 1475 3774 1509 3814
rect 1475 3700 1509 3740
rect 1475 3626 1509 3666
rect 1475 3552 1509 3592
rect 1475 3478 1509 3518
rect 1475 3404 1509 3444
rect 1475 3330 1509 3370
rect 1475 3256 1509 3296
rect 1475 3182 1509 3222
rect 1475 3108 1509 3148
rect 1475 3034 1509 3074
rect 1475 2960 1509 3000
rect 1711 4799 1745 4838
rect 1711 4726 1745 4765
rect 1711 4653 1745 4692
rect 1711 4580 1745 4619
rect 1711 4507 1745 4546
rect 1711 4434 1745 4473
rect 1711 4361 1745 4400
rect 1711 4288 1745 4327
rect 1711 4215 1745 4254
rect 1711 4142 1745 4181
rect 1711 4069 1745 4108
rect 1711 3996 1745 4035
rect 1711 3922 1745 3962
rect 1711 3848 1745 3888
rect 1711 3774 1745 3814
rect 1711 3700 1745 3740
rect 1711 3626 1745 3666
rect 1711 3552 1745 3592
rect 1711 3478 1745 3518
rect 1711 3404 1745 3444
rect 1711 3330 1745 3370
rect 1711 3256 1745 3296
rect 1711 3182 1745 3222
rect 1711 3108 1745 3148
rect 1711 3034 1745 3074
rect 1711 2960 1745 3000
rect 1947 4799 1981 4838
rect 1947 4726 1981 4765
rect 1947 4653 1981 4692
rect 1947 4580 1981 4619
rect 1947 4507 1981 4546
rect 1947 4434 1981 4473
rect 1947 4361 1981 4400
rect 1947 4288 1981 4327
rect 1947 4215 1981 4254
rect 1947 4142 1981 4181
rect 1947 4069 1981 4108
rect 1947 3996 1981 4035
rect 1947 3922 1981 3962
rect 1947 3848 1981 3888
rect 1947 3774 1981 3814
rect 1947 3700 1981 3740
rect 1947 3626 1981 3666
rect 1947 3552 1981 3592
rect 1947 3478 1981 3518
rect 1947 3404 1981 3444
rect 1947 3330 1981 3370
rect 1947 3256 1981 3296
rect 1947 3182 1981 3222
rect 1947 3108 1981 3148
rect 1947 3034 1981 3074
rect 1947 2960 1981 3000
rect 2183 4799 2217 4838
rect 2183 4726 2217 4765
rect 2183 4653 2217 4692
rect 2183 4580 2217 4619
rect 2183 4507 2217 4546
rect 2183 4434 2217 4473
rect 2183 4361 2217 4400
rect 2183 4288 2217 4327
rect 2183 4215 2217 4254
rect 2183 4142 2217 4181
rect 2183 4069 2217 4108
rect 2183 3996 2217 4035
rect 2183 3922 2217 3962
rect 2183 3848 2217 3888
rect 2183 3774 2217 3814
rect 2183 3700 2217 3740
rect 2183 3626 2217 3666
rect 2183 3552 2217 3592
rect 2183 3478 2217 3518
rect 2183 3404 2217 3444
rect 2183 3330 2217 3370
rect 2183 3256 2217 3296
rect 2183 3182 2217 3222
rect 2183 3108 2217 3148
rect 2183 3034 2217 3074
rect 2183 2960 2217 3000
rect 2419 4799 2453 4838
rect 2419 4726 2453 4765
rect 2419 4653 2453 4692
rect 2419 4580 2453 4619
rect 2419 4507 2453 4546
rect 2419 4434 2453 4473
rect 2419 4361 2453 4400
rect 2419 4288 2453 4327
rect 2419 4215 2453 4254
rect 2419 4142 2453 4181
rect 2419 4069 2453 4108
rect 2419 3996 2453 4035
rect 2419 3922 2453 3962
rect 2419 3848 2453 3888
rect 2419 3774 2453 3814
rect 2419 3700 2453 3740
rect 2419 3626 2453 3666
rect 2419 3552 2453 3592
rect 2419 3478 2453 3518
rect 2419 3404 2453 3444
rect 2419 3330 2453 3370
rect 2419 3256 2453 3296
rect 2419 3182 2453 3222
rect 2419 3108 2453 3148
rect 2419 3034 2453 3074
rect 2419 2960 2453 3000
rect 2655 4799 2689 4838
rect 2655 4726 2689 4765
rect 2655 4653 2689 4692
rect 2655 4580 2689 4619
rect 2655 4507 2689 4546
rect 2655 4434 2689 4473
rect 2655 4361 2689 4400
rect 2655 4288 2689 4327
rect 2655 4215 2689 4254
rect 2655 4142 2689 4181
rect 2655 4069 2689 4108
rect 2655 3996 2689 4035
rect 2655 3922 2689 3962
rect 2655 3848 2689 3888
rect 2655 3774 2689 3814
rect 2655 3700 2689 3740
rect 2655 3626 2689 3666
rect 2655 3552 2689 3592
rect 2655 3478 2689 3518
rect 2655 3404 2689 3444
rect 2655 3330 2689 3370
rect 2655 3256 2689 3296
rect 2655 3182 2689 3222
rect 2655 3108 2689 3148
rect 2655 3034 2689 3074
rect 2655 2960 2689 3000
rect 2891 4799 2925 4838
rect 2891 4726 2925 4765
rect 2891 4653 2925 4692
rect 2891 4580 2925 4619
rect 2891 4507 2925 4546
rect 2891 4434 2925 4473
rect 2891 4361 2925 4400
rect 2891 4288 2925 4327
rect 2891 4215 2925 4254
rect 2891 4142 2925 4181
rect 2891 4069 2925 4108
rect 2891 3996 2925 4035
rect 2891 3922 2925 3962
rect 2891 3848 2925 3888
rect 2891 3774 2925 3814
rect 2891 3700 2925 3740
rect 2891 3626 2925 3666
rect 2891 3552 2925 3592
rect 2891 3478 2925 3518
rect 2891 3404 2925 3444
rect 2891 3330 2925 3370
rect 2891 3256 2925 3296
rect 2891 3182 2925 3222
rect 2891 3108 2925 3148
rect 2891 3034 2925 3074
rect 2891 2960 2925 3000
rect 3023 4838 3083 4872
rect 3023 4800 3036 4838
rect 3070 4800 3083 4838
rect 3023 4770 3083 4800
rect 3023 4728 3036 4770
rect 3070 4728 3083 4770
rect 3023 4702 3083 4728
rect 3023 4656 3036 4702
rect 3070 4656 3083 4702
rect 3023 4634 3083 4656
rect 3023 4584 3036 4634
rect 3070 4584 3083 4634
rect 3023 4566 3083 4584
rect 3023 4512 3036 4566
rect 3070 4512 3083 4566
rect 3023 4498 3083 4512
rect 3023 4440 3036 4498
rect 3070 4440 3083 4498
rect 3023 4430 3083 4440
rect 3023 4368 3036 4430
rect 3070 4368 3083 4430
rect 3023 4362 3083 4368
rect 3023 4296 3036 4362
rect 3070 4296 3083 4362
rect 3023 4294 3083 4296
rect 3023 4260 3036 4294
rect 3070 4260 3083 4294
rect 3023 4258 3083 4260
rect 3023 4192 3036 4258
rect 3070 4192 3083 4258
rect 3023 4186 3083 4192
rect 3023 4124 3036 4186
rect 3070 4124 3083 4186
rect 3023 4114 3083 4124
rect 3023 4056 3036 4114
rect 3070 4056 3083 4114
rect 3023 4042 3083 4056
rect 3023 3988 3036 4042
rect 3070 3988 3083 4042
rect 3023 3970 3083 3988
rect 3023 3920 3036 3970
rect 3070 3920 3083 3970
rect 3023 3898 3083 3920
rect 3023 3852 3036 3898
rect 3070 3852 3083 3898
rect 3023 3826 3083 3852
rect 3023 3784 3036 3826
rect 3070 3784 3083 3826
rect 3023 3754 3083 3784
rect 3023 3716 3036 3754
rect 3070 3716 3083 3754
rect 3023 3682 3083 3716
rect 3023 3648 3036 3682
rect 3070 3648 3083 3682
rect 3023 3614 3083 3648
rect 3023 3576 3036 3614
rect 3070 3576 3083 3614
rect 3023 3546 3083 3576
rect 3023 3504 3036 3546
rect 3070 3504 3083 3546
rect 3023 3478 3083 3504
rect 3023 3432 3036 3478
rect 3070 3432 3083 3478
rect 3023 3410 3083 3432
rect 3023 3360 3036 3410
rect 3070 3360 3083 3410
rect 3023 3342 3083 3360
rect 3023 3288 3036 3342
rect 3070 3288 3083 3342
rect 3023 3274 3083 3288
rect 3023 3216 3036 3274
rect 3070 3216 3083 3274
rect 3023 3206 3083 3216
rect 3023 3144 3036 3206
rect 3070 3144 3083 3206
rect 3023 3138 3083 3144
rect 3023 3072 3036 3138
rect 3070 3072 3083 3138
rect 3023 3070 3083 3072
rect 3023 3036 3036 3070
rect 3070 3036 3083 3070
rect 3023 3034 3083 3036
rect 3023 2968 3036 3034
rect 3070 2968 3083 3034
rect 3023 2962 3083 2968
rect 373 2879 433 2909
rect 373 2837 386 2879
rect 420 2837 433 2879
rect 3023 2900 3036 2962
rect 3070 2900 3083 2962
rect 3023 2890 3083 2900
rect 373 2811 433 2837
rect 373 2765 386 2811
rect 420 2765 433 2811
rect 576 2810 592 2844
rect 659 2810 662 2844
rect 696 2810 700 2844
rect 766 2810 775 2844
rect 836 2810 850 2844
rect 906 2810 925 2844
rect 976 2810 1000 2844
rect 1046 2810 1075 2844
rect 1116 2810 1150 2844
rect 1186 2810 1222 2844
rect 1259 2810 1292 2844
rect 1334 2810 1362 2844
rect 1409 2810 1432 2844
rect 1484 2810 1502 2844
rect 1559 2810 1572 2844
rect 1634 2810 1642 2844
rect 1708 2810 1712 2844
rect 1746 2810 1748 2844
rect 1816 2810 1822 2844
rect 1886 2810 1896 2844
rect 1956 2810 1970 2844
rect 2026 2810 2044 2844
rect 2096 2810 2118 2844
rect 2166 2810 2192 2844
rect 2236 2810 2266 2844
rect 2306 2810 2340 2844
rect 2376 2810 2412 2844
rect 2448 2810 2482 2844
rect 2522 2810 2552 2844
rect 2596 2810 2622 2844
rect 2670 2810 2692 2844
rect 2744 2810 2761 2844
rect 2818 2810 2830 2844
rect 2864 2810 2880 2844
rect 3023 2832 3036 2890
rect 3070 2832 3083 2890
rect 3023 2818 3083 2832
rect 373 2743 433 2765
rect 373 2693 386 2743
rect 420 2693 433 2743
rect 3023 2764 3036 2818
rect 3070 2764 3083 2818
rect 3023 2746 3083 2764
rect 373 2675 433 2693
rect 373 2621 386 2675
rect 420 2621 433 2675
rect 373 2607 433 2621
rect 373 2549 386 2607
rect 420 2549 433 2607
rect 373 2539 433 2549
rect 373 2477 386 2539
rect 420 2477 433 2539
rect 373 2471 433 2477
rect 373 2405 386 2471
rect 420 2405 433 2471
rect 373 2403 433 2405
rect 373 2369 386 2403
rect 420 2369 433 2403
rect 373 2367 433 2369
rect 373 2301 386 2367
rect 420 2301 433 2367
rect 373 2295 433 2301
rect 373 2233 386 2295
rect 420 2233 433 2295
rect 373 2223 433 2233
rect 373 2165 386 2223
rect 420 2165 433 2223
rect 373 2151 433 2165
rect 373 2097 386 2151
rect 420 2097 433 2151
rect 373 2079 433 2097
rect 373 2029 386 2079
rect 420 2029 433 2079
rect 373 2007 433 2029
rect 373 1961 386 2007
rect 420 1961 433 2007
rect 373 1935 433 1961
rect 373 1893 386 1935
rect 420 1893 433 1935
rect 373 1863 433 1893
rect 373 1825 386 1863
rect 420 1825 433 1863
rect 373 1791 433 1825
rect 373 1757 386 1791
rect 420 1757 433 1791
rect 373 1723 433 1757
rect 373 1685 386 1723
rect 420 1685 433 1723
rect 373 1655 433 1685
rect 373 1613 386 1655
rect 420 1613 433 1655
rect 373 1587 433 1613
rect 373 1541 386 1587
rect 420 1541 433 1587
rect 373 1519 433 1541
rect 373 1469 386 1519
rect 420 1469 433 1519
rect 373 1451 433 1469
rect 373 1397 386 1451
rect 420 1397 433 1451
rect 373 1383 433 1397
rect 373 1325 386 1383
rect 420 1325 433 1383
rect 373 1315 433 1325
rect 373 1253 386 1315
rect 420 1253 433 1315
rect 373 1247 433 1253
rect 373 1181 386 1247
rect 420 1181 433 1247
rect 373 1179 433 1181
rect 373 1145 386 1179
rect 420 1145 433 1179
rect 373 1143 433 1145
rect 373 1077 386 1143
rect 420 1077 433 1143
rect 373 1071 433 1077
rect 373 1009 386 1071
rect 420 1009 433 1071
rect 373 999 433 1009
rect 373 941 386 999
rect 420 941 433 999
rect 373 927 433 941
rect 373 873 386 927
rect 420 873 433 927
rect 373 855 433 873
rect 373 805 386 855
rect 420 805 433 855
rect 373 783 433 805
rect 373 737 386 783
rect 420 737 433 783
rect 531 2647 565 2686
rect 531 2574 565 2613
rect 531 2501 565 2540
rect 531 2428 565 2467
rect 531 2355 565 2394
rect 531 2282 565 2321
rect 531 2209 565 2248
rect 531 2136 565 2175
rect 531 2063 565 2102
rect 531 1990 565 2029
rect 531 1917 565 1956
rect 531 1844 565 1883
rect 531 1770 565 1810
rect 531 1696 565 1736
rect 531 1622 565 1662
rect 531 1548 565 1588
rect 531 1474 565 1514
rect 531 1400 565 1440
rect 531 1326 565 1366
rect 531 1252 565 1292
rect 531 1178 565 1218
rect 531 1104 565 1144
rect 531 1030 565 1070
rect 531 956 565 996
rect 531 882 565 922
rect 531 808 565 848
rect 767 2647 801 2686
rect 767 2574 801 2613
rect 767 2501 801 2540
rect 767 2428 801 2467
rect 767 2355 801 2394
rect 767 2282 801 2321
rect 767 2209 801 2248
rect 767 2136 801 2175
rect 767 2063 801 2102
rect 767 1990 801 2029
rect 767 1917 801 1956
rect 767 1844 801 1883
rect 767 1770 801 1810
rect 767 1696 801 1736
rect 767 1622 801 1662
rect 767 1548 801 1588
rect 767 1474 801 1514
rect 767 1400 801 1440
rect 767 1326 801 1366
rect 767 1252 801 1292
rect 767 1178 801 1218
rect 767 1104 801 1144
rect 767 1030 801 1070
rect 767 956 801 996
rect 767 882 801 922
rect 767 808 801 848
rect 1003 2647 1037 2686
rect 1003 2574 1037 2613
rect 1003 2501 1037 2540
rect 1003 2428 1037 2467
rect 1003 2355 1037 2394
rect 1003 2282 1037 2321
rect 1003 2209 1037 2248
rect 1003 2136 1037 2175
rect 1003 2063 1037 2102
rect 1003 1990 1037 2029
rect 1003 1917 1037 1956
rect 1003 1844 1037 1883
rect 1003 1770 1037 1810
rect 1003 1696 1037 1736
rect 1003 1622 1037 1662
rect 1003 1548 1037 1588
rect 1003 1474 1037 1514
rect 1003 1400 1037 1440
rect 1003 1326 1037 1366
rect 1003 1252 1037 1292
rect 1003 1178 1037 1218
rect 1003 1104 1037 1144
rect 1003 1030 1037 1070
rect 1003 956 1037 996
rect 1003 882 1037 922
rect 1003 808 1037 848
rect 1239 2647 1273 2686
rect 1239 2574 1273 2613
rect 1239 2501 1273 2540
rect 1239 2428 1273 2467
rect 1239 2355 1273 2394
rect 1239 2282 1273 2321
rect 1239 2209 1273 2248
rect 1239 2136 1273 2175
rect 1239 2063 1273 2102
rect 1239 1990 1273 2029
rect 1239 1917 1273 1956
rect 1239 1844 1273 1883
rect 1239 1770 1273 1810
rect 1239 1696 1273 1736
rect 1239 1622 1273 1662
rect 1239 1548 1273 1588
rect 1239 1474 1273 1514
rect 1239 1400 1273 1440
rect 1239 1326 1273 1366
rect 1239 1252 1273 1292
rect 1239 1178 1273 1218
rect 1239 1104 1273 1144
rect 1239 1030 1273 1070
rect 1239 956 1273 996
rect 1239 882 1273 922
rect 1239 808 1273 848
rect 1475 2647 1509 2686
rect 1475 2574 1509 2613
rect 1475 2501 1509 2540
rect 1475 2428 1509 2467
rect 1475 2355 1509 2394
rect 1475 2282 1509 2321
rect 1475 2209 1509 2248
rect 1475 2136 1509 2175
rect 1475 2063 1509 2102
rect 1475 1990 1509 2029
rect 1475 1917 1509 1956
rect 1475 1844 1509 1883
rect 1475 1770 1509 1810
rect 1475 1696 1509 1736
rect 1475 1622 1509 1662
rect 1475 1548 1509 1588
rect 1475 1474 1509 1514
rect 1475 1400 1509 1440
rect 1475 1326 1509 1366
rect 1475 1252 1509 1292
rect 1475 1178 1509 1218
rect 1475 1104 1509 1144
rect 1475 1030 1509 1070
rect 1475 956 1509 996
rect 1475 882 1509 922
rect 1475 808 1509 848
rect 1711 2647 1745 2686
rect 1711 2574 1745 2613
rect 1711 2501 1745 2540
rect 1711 2428 1745 2467
rect 1711 2355 1745 2394
rect 1711 2282 1745 2321
rect 1711 2209 1745 2248
rect 1711 2136 1745 2175
rect 1711 2063 1745 2102
rect 1711 1990 1745 2029
rect 1711 1917 1745 1956
rect 1711 1844 1745 1883
rect 1711 1770 1745 1810
rect 1711 1696 1745 1736
rect 1711 1622 1745 1662
rect 1711 1548 1745 1588
rect 1711 1474 1745 1514
rect 1711 1400 1745 1440
rect 1711 1326 1745 1366
rect 1711 1252 1745 1292
rect 1711 1178 1745 1218
rect 1711 1104 1745 1144
rect 1711 1030 1745 1070
rect 1711 956 1745 996
rect 1711 882 1745 922
rect 1711 808 1745 848
rect 1947 2647 1981 2686
rect 1947 2574 1981 2613
rect 1947 2501 1981 2540
rect 1947 2428 1981 2467
rect 1947 2355 1981 2394
rect 1947 2282 1981 2321
rect 1947 2209 1981 2248
rect 1947 2136 1981 2175
rect 1947 2063 1981 2102
rect 1947 1990 1981 2029
rect 1947 1917 1981 1956
rect 1947 1844 1981 1883
rect 1947 1770 1981 1810
rect 1947 1696 1981 1736
rect 1947 1622 1981 1662
rect 1947 1548 1981 1588
rect 1947 1474 1981 1514
rect 1947 1400 1981 1440
rect 1947 1326 1981 1366
rect 1947 1252 1981 1292
rect 1947 1178 1981 1218
rect 1947 1104 1981 1144
rect 1947 1030 1981 1070
rect 1947 956 1981 996
rect 1947 882 1981 922
rect 1947 808 1981 848
rect 2183 2647 2217 2686
rect 2183 2574 2217 2613
rect 2183 2501 2217 2540
rect 2183 2428 2217 2467
rect 2183 2355 2217 2394
rect 2183 2282 2217 2321
rect 2183 2209 2217 2248
rect 2183 2136 2217 2175
rect 2183 2063 2217 2102
rect 2183 1990 2217 2029
rect 2183 1917 2217 1956
rect 2183 1844 2217 1883
rect 2183 1770 2217 1810
rect 2183 1696 2217 1736
rect 2183 1622 2217 1662
rect 2183 1548 2217 1588
rect 2183 1474 2217 1514
rect 2183 1400 2217 1440
rect 2183 1326 2217 1366
rect 2183 1252 2217 1292
rect 2183 1178 2217 1218
rect 2183 1104 2217 1144
rect 2183 1030 2217 1070
rect 2183 956 2217 996
rect 2183 882 2217 922
rect 2183 808 2217 848
rect 2419 2647 2453 2686
rect 2419 2574 2453 2613
rect 2419 2501 2453 2540
rect 2419 2428 2453 2467
rect 2419 2355 2453 2394
rect 2419 2282 2453 2321
rect 2419 2209 2453 2248
rect 2419 2136 2453 2175
rect 2419 2063 2453 2102
rect 2419 1990 2453 2029
rect 2419 1917 2453 1956
rect 2419 1844 2453 1883
rect 2419 1770 2453 1810
rect 2419 1696 2453 1736
rect 2419 1622 2453 1662
rect 2419 1548 2453 1588
rect 2419 1474 2453 1514
rect 2419 1400 2453 1440
rect 2419 1326 2453 1366
rect 2419 1252 2453 1292
rect 2419 1178 2453 1218
rect 2419 1104 2453 1144
rect 2419 1030 2453 1070
rect 2419 956 2453 996
rect 2419 882 2453 922
rect 2419 808 2453 848
rect 2655 2647 2689 2686
rect 2655 2574 2689 2613
rect 2655 2501 2689 2540
rect 2655 2428 2689 2467
rect 2655 2355 2689 2394
rect 2655 2282 2689 2321
rect 2655 2209 2689 2248
rect 2655 2136 2689 2175
rect 2655 2063 2689 2102
rect 2655 1990 2689 2029
rect 2655 1917 2689 1956
rect 2655 1844 2689 1883
rect 2655 1770 2689 1810
rect 2655 1696 2689 1736
rect 2655 1622 2689 1662
rect 2655 1548 2689 1588
rect 2655 1474 2689 1514
rect 2655 1400 2689 1440
rect 2655 1326 2689 1366
rect 2655 1252 2689 1292
rect 2655 1178 2689 1218
rect 2655 1104 2689 1144
rect 2655 1030 2689 1070
rect 2655 956 2689 996
rect 2655 882 2689 922
rect 2655 808 2689 848
rect 2891 2639 2925 2678
rect 2891 2566 2925 2605
rect 2891 2493 2925 2532
rect 2891 2420 2925 2459
rect 2891 2347 2925 2386
rect 2891 2274 2925 2313
rect 2891 2201 2925 2240
rect 2891 2128 2925 2167
rect 2891 2055 2925 2094
rect 2891 1982 2925 2021
rect 2891 1909 2925 1948
rect 2891 1836 2925 1875
rect 2891 1762 2925 1802
rect 2891 1688 2925 1728
rect 2891 1614 2925 1654
rect 2891 1540 2925 1580
rect 2891 1466 2925 1506
rect 2891 1392 2925 1432
rect 2891 1318 2925 1358
rect 2891 1244 2925 1284
rect 2891 1170 2925 1210
rect 2891 1096 2925 1136
rect 2891 1022 2925 1062
rect 2891 948 2925 988
rect 2891 874 2925 914
rect 2891 800 2925 840
rect 3023 2696 3036 2746
rect 3070 2696 3083 2746
rect 3023 2674 3083 2696
rect 3023 2628 3036 2674
rect 3070 2628 3083 2674
rect 3023 2602 3083 2628
rect 3023 2560 3036 2602
rect 3070 2560 3083 2602
rect 3023 2530 3083 2560
rect 3023 2492 3036 2530
rect 3070 2492 3083 2530
rect 3023 2458 3083 2492
rect 3023 2424 3036 2458
rect 3070 2424 3083 2458
rect 3023 2390 3083 2424
rect 3023 2352 3036 2390
rect 3070 2352 3083 2390
rect 3023 2322 3083 2352
rect 3023 2280 3036 2322
rect 3070 2280 3083 2322
rect 3023 2254 3083 2280
rect 3023 2208 3036 2254
rect 3070 2208 3083 2254
rect 3023 2186 3083 2208
rect 3023 2136 3036 2186
rect 3070 2136 3083 2186
rect 3023 2118 3083 2136
rect 3023 2064 3036 2118
rect 3070 2064 3083 2118
rect 3023 2050 3083 2064
rect 3023 1992 3036 2050
rect 3070 1992 3083 2050
rect 3023 1982 3083 1992
rect 3023 1919 3036 1982
rect 3070 1919 3083 1982
rect 3023 1914 3083 1919
rect 3023 1812 3036 1914
rect 3070 1812 3083 1914
rect 3023 1807 3083 1812
rect 3023 1744 3036 1807
rect 3070 1744 3083 1807
rect 3023 1734 3083 1744
rect 3023 1676 3036 1734
rect 3070 1676 3083 1734
rect 3023 1661 3083 1676
rect 3023 1608 3036 1661
rect 3070 1608 3083 1661
rect 3023 1588 3083 1608
rect 3023 1540 3036 1588
rect 3070 1540 3083 1588
rect 3023 1515 3083 1540
rect 3023 1472 3036 1515
rect 3070 1472 3083 1515
rect 3023 1442 3083 1472
rect 3023 1404 3036 1442
rect 3070 1404 3083 1442
rect 3023 1370 3083 1404
rect 3023 1335 3036 1370
rect 3070 1335 3083 1370
rect 3023 1302 3083 1335
rect 3023 1262 3036 1302
rect 3070 1262 3083 1302
rect 3023 1234 3083 1262
rect 3023 1189 3036 1234
rect 3070 1189 3083 1234
rect 3023 1166 3083 1189
rect 3023 1116 3036 1166
rect 3070 1116 3083 1166
rect 3023 1098 3083 1116
rect 3023 1043 3036 1098
rect 3070 1043 3083 1098
rect 3023 1030 3083 1043
rect 3023 970 3036 1030
rect 3070 970 3083 1030
rect 3023 962 3083 970
rect 3023 897 3036 962
rect 3070 897 3083 962
rect 3023 894 3083 897
rect 3023 860 3036 894
rect 3070 860 3083 894
rect 3023 858 3083 860
rect 3023 792 3036 858
rect 3070 792 3083 858
rect 3023 785 3083 792
rect 373 711 433 737
rect 3023 724 3036 785
rect 3070 724 3083 785
rect 373 669 386 711
rect 420 669 433 711
rect 576 680 592 714
rect 659 680 662 714
rect 696 680 700 714
rect 766 680 775 714
rect 836 680 850 714
rect 906 680 925 714
rect 976 680 1000 714
rect 1046 680 1075 714
rect 1116 680 1150 714
rect 1186 680 1222 714
rect 1259 680 1292 714
rect 1334 680 1362 714
rect 1409 680 1432 714
rect 1484 680 1502 714
rect 1559 680 1572 714
rect 1634 680 1642 714
rect 1708 680 1712 714
rect 1746 680 1748 714
rect 1816 680 1822 714
rect 1886 680 1896 714
rect 1956 680 1970 714
rect 2026 680 2044 714
rect 2096 680 2118 714
rect 2166 680 2192 714
rect 2236 680 2266 714
rect 2306 680 2340 714
rect 2376 680 2412 714
rect 2448 680 2482 714
rect 2522 680 2552 714
rect 2596 680 2622 714
rect 2670 680 2692 714
rect 2744 680 2761 714
rect 2818 680 2830 714
rect 2864 680 2880 714
rect 3023 712 3083 724
rect 373 639 433 669
rect 373 605 386 639
rect 420 605 433 639
rect 373 580 433 605
rect 3023 656 3036 712
rect 3070 656 3083 712
rect 3023 639 3083 656
rect 3023 588 3036 639
rect 3070 588 3083 639
rect 3023 580 3083 588
rect 373 567 3083 580
rect 373 533 441 567
rect 492 533 509 567
rect 566 533 577 567
rect 640 533 645 567
rect 679 533 680 567
rect 747 533 754 567
rect 815 533 828 567
rect 883 533 902 567
rect 951 533 976 567
rect 1019 533 1050 567
rect 1087 533 1121 567
rect 1158 533 1189 567
rect 1232 533 1257 567
rect 1306 533 1325 567
rect 1380 533 1393 567
rect 1454 533 1461 567
rect 1528 533 1529 567
rect 1563 533 1568 567
rect 1631 533 1642 567
rect 1699 533 1716 567
rect 1767 533 1790 567
rect 1835 533 1864 567
rect 1903 533 1937 567
rect 1972 533 2005 567
rect 2046 533 2073 567
rect 2120 533 2141 567
rect 2194 533 2209 567
rect 2267 533 2277 567
rect 2340 533 2345 567
rect 2447 533 2452 567
rect 2515 533 2525 567
rect 2583 533 2598 567
rect 2651 533 2671 567
rect 2719 533 2744 567
rect 2787 533 2817 567
rect 2855 533 2889 567
rect 2924 533 2957 567
rect 2997 533 3083 567
rect 373 520 3083 533
rect 3290 39158 3296 39260
rect 3330 39158 3336 39260
rect 3290 39154 3336 39158
rect 3290 39090 3296 39154
rect 3330 39090 3336 39154
rect 3290 39082 3336 39090
rect 3290 39022 3296 39082
rect 3330 39022 3336 39082
rect 3290 39010 3336 39022
rect 3290 38954 3296 39010
rect 3330 38954 3336 39010
rect 3290 38938 3336 38954
rect 3290 38886 3296 38938
rect 3330 38886 3336 38938
rect 3290 38866 3336 38886
rect 3290 38818 3296 38866
rect 3330 38818 3336 38866
rect 3290 38794 3336 38818
rect 3290 38750 3296 38794
rect 3330 38750 3336 38794
rect 3290 38722 3336 38750
rect 3290 38682 3296 38722
rect 3330 38682 3336 38722
rect 3290 38650 3336 38682
rect 3290 38614 3296 38650
rect 3330 38614 3336 38650
rect 3290 38580 3336 38614
rect 3290 38544 3296 38580
rect 3330 38544 3336 38580
rect 3290 38512 3336 38544
rect 3290 38472 3296 38512
rect 3330 38472 3336 38512
rect 3290 38444 3336 38472
rect 3290 38400 3296 38444
rect 3330 38400 3336 38444
rect 3290 38376 3336 38400
rect 3290 38328 3296 38376
rect 3330 38328 3336 38376
rect 3290 38308 3336 38328
rect 3290 38256 3296 38308
rect 3330 38256 3336 38308
rect 3290 38240 3336 38256
rect 3290 38184 3296 38240
rect 3330 38184 3336 38240
rect 3290 38172 3336 38184
rect 3290 38112 3296 38172
rect 3330 38112 3336 38172
rect 3290 38104 3336 38112
rect 3290 38040 3296 38104
rect 3330 38040 3336 38104
rect 3290 38036 3336 38040
rect 3290 37934 3296 38036
rect 3330 37934 3336 38036
rect 3290 37930 3336 37934
rect 3290 37866 3296 37930
rect 3330 37866 3336 37930
rect 3290 37858 3336 37866
rect 3290 37798 3296 37858
rect 3330 37798 3336 37858
rect 3290 37786 3336 37798
rect 3290 37730 3296 37786
rect 3330 37730 3336 37786
rect 3290 37714 3336 37730
rect 3290 37662 3296 37714
rect 3330 37662 3336 37714
rect 3290 37642 3336 37662
rect 3290 37594 3296 37642
rect 3330 37594 3336 37642
rect 3290 37570 3336 37594
rect 3290 37526 3296 37570
rect 3330 37526 3336 37570
rect 3290 37498 3336 37526
rect 3290 37458 3296 37498
rect 3330 37458 3336 37498
rect 3290 37426 3336 37458
rect 3290 37390 3296 37426
rect 3330 37390 3336 37426
rect 3290 37356 3336 37390
rect 3290 37320 3296 37356
rect 3330 37320 3336 37356
rect 3290 37288 3336 37320
rect 3290 37248 3296 37288
rect 3330 37248 3336 37288
rect 3290 37220 3336 37248
rect 3290 37176 3296 37220
rect 3330 37176 3336 37220
rect 3290 37152 3336 37176
rect 3290 37104 3296 37152
rect 3330 37104 3336 37152
rect 3290 37084 3336 37104
rect 3290 37032 3296 37084
rect 3330 37032 3336 37084
rect 3290 37016 3336 37032
rect 3290 36960 3296 37016
rect 3330 36960 3336 37016
rect 3290 36948 3336 36960
rect 3290 36888 3296 36948
rect 3330 36888 3336 36948
rect 3290 36880 3336 36888
rect 3290 36816 3296 36880
rect 3330 36816 3336 36880
rect 3290 36812 3336 36816
rect 3290 36710 3296 36812
rect 3330 36710 3336 36812
rect 3290 36706 3336 36710
rect 3290 36642 3296 36706
rect 3330 36642 3336 36706
rect 3290 36634 3336 36642
rect 3290 36574 3296 36634
rect 3330 36574 3336 36634
rect 3290 36562 3336 36574
rect 3290 36506 3296 36562
rect 3330 36506 3336 36562
rect 3290 36490 3336 36506
rect 3290 36438 3296 36490
rect 3330 36438 3336 36490
rect 3290 36418 3336 36438
rect 3290 36370 3296 36418
rect 3330 36370 3336 36418
rect 3290 36346 3336 36370
rect 3290 36302 3296 36346
rect 3330 36302 3336 36346
rect 3290 36274 3336 36302
rect 3290 36234 3296 36274
rect 3330 36234 3336 36274
rect 3290 36202 3336 36234
rect 3290 36166 3296 36202
rect 3330 36166 3336 36202
rect 3290 36132 3336 36166
rect 3290 36096 3296 36132
rect 3330 36096 3336 36132
rect 3290 36064 3336 36096
rect 3290 36024 3296 36064
rect 3330 36024 3336 36064
rect 3290 35996 3336 36024
rect 3290 35952 3296 35996
rect 3330 35952 3336 35996
rect 3290 35928 3336 35952
rect 3290 35880 3296 35928
rect 3330 35880 3336 35928
rect 3290 35860 3336 35880
rect 3290 35808 3296 35860
rect 3330 35808 3336 35860
rect 3290 35792 3336 35808
rect 3290 35736 3296 35792
rect 3330 35736 3336 35792
rect 3290 35724 3336 35736
rect 3290 35664 3296 35724
rect 3330 35664 3336 35724
rect 3290 35656 3336 35664
rect 3290 35592 3296 35656
rect 3330 35592 3336 35656
rect 3290 35588 3336 35592
rect 3290 35486 3296 35588
rect 3330 35486 3336 35588
rect 3290 35482 3336 35486
rect 3290 35418 3296 35482
rect 3330 35418 3336 35482
rect 3290 35410 3336 35418
rect 3290 35350 3296 35410
rect 3330 35350 3336 35410
rect 3290 35338 3336 35350
rect 3290 35282 3296 35338
rect 3330 35282 3336 35338
rect 3290 35266 3336 35282
rect 3290 35214 3296 35266
rect 3330 35214 3336 35266
rect 3290 35194 3336 35214
rect 3290 35146 3296 35194
rect 3330 35146 3336 35194
rect 3290 35122 3336 35146
rect 3290 35078 3296 35122
rect 3330 35078 3336 35122
rect 3290 35050 3336 35078
rect 3290 35010 3296 35050
rect 3330 35010 3336 35050
rect 3290 34978 3336 35010
rect 3290 34942 3296 34978
rect 3330 34942 3336 34978
rect 3290 34908 3336 34942
rect 3290 34872 3296 34908
rect 3330 34872 3336 34908
rect 3290 34840 3336 34872
rect 3290 34800 3296 34840
rect 3330 34800 3336 34840
rect 3290 34772 3336 34800
rect 3290 34728 3296 34772
rect 3330 34728 3336 34772
rect 3290 34704 3336 34728
rect 3290 34656 3296 34704
rect 3330 34656 3336 34704
rect 3290 34636 3336 34656
rect 3290 34584 3296 34636
rect 3330 34584 3336 34636
rect 3290 34568 3336 34584
rect 3290 34512 3296 34568
rect 3330 34512 3336 34568
rect 3290 34500 3336 34512
rect 3290 34440 3296 34500
rect 3330 34440 3336 34500
rect 3290 34432 3336 34440
rect 3290 34368 3296 34432
rect 3330 34368 3336 34432
rect 3290 34364 3336 34368
rect 3290 34262 3296 34364
rect 3330 34262 3336 34364
rect 3290 34258 3336 34262
rect 3290 34194 3296 34258
rect 3330 34194 3336 34258
rect 3290 34186 3336 34194
rect 3290 34126 3296 34186
rect 3330 34126 3336 34186
rect 3290 34114 3336 34126
rect 3290 34058 3296 34114
rect 3330 34058 3336 34114
rect 3290 34042 3336 34058
rect 3290 33990 3296 34042
rect 3330 33990 3336 34042
rect 3290 33970 3336 33990
rect 3290 33922 3296 33970
rect 3330 33922 3336 33970
rect 3290 33898 3336 33922
rect 3290 33854 3296 33898
rect 3330 33854 3336 33898
rect 3290 33826 3336 33854
rect 3290 33786 3296 33826
rect 3330 33786 3336 33826
rect 3290 33754 3336 33786
rect 3290 33718 3296 33754
rect 3330 33718 3336 33754
rect 3290 33684 3336 33718
rect 3290 33648 3296 33684
rect 3330 33648 3336 33684
rect 3290 33616 3336 33648
rect 3290 33576 3296 33616
rect 3330 33576 3336 33616
rect 3290 33548 3336 33576
rect 3290 33504 3296 33548
rect 3330 33504 3336 33548
rect 3290 33480 3336 33504
rect 3290 33432 3296 33480
rect 3330 33432 3336 33480
rect 3290 33412 3336 33432
rect 3290 33360 3296 33412
rect 3330 33360 3336 33412
rect 3290 33344 3336 33360
rect 3290 33288 3296 33344
rect 3330 33288 3336 33344
rect 3290 33276 3336 33288
rect 3290 33216 3296 33276
rect 3330 33216 3336 33276
rect 3290 33208 3336 33216
rect 3290 33144 3296 33208
rect 3330 33144 3336 33208
rect 3290 33140 3336 33144
rect 3290 33038 3296 33140
rect 3330 33038 3336 33140
rect 3290 33034 3336 33038
rect 3290 32970 3296 33034
rect 3330 32970 3336 33034
rect 3290 32962 3336 32970
rect 3290 32902 3296 32962
rect 3330 32902 3336 32962
rect 3290 32890 3336 32902
rect 3290 32834 3296 32890
rect 3330 32834 3336 32890
rect 3290 32818 3336 32834
rect 3290 32766 3296 32818
rect 3330 32766 3336 32818
rect 3290 32746 3336 32766
rect 3290 32698 3296 32746
rect 3330 32698 3336 32746
rect 3290 32674 3336 32698
rect 3290 32630 3296 32674
rect 3330 32630 3336 32674
rect 3290 32602 3336 32630
rect 3290 32562 3296 32602
rect 3330 32562 3336 32602
rect 3290 32530 3336 32562
rect 3290 32494 3296 32530
rect 3330 32494 3336 32530
rect 3290 32460 3336 32494
rect 3290 32424 3296 32460
rect 3330 32424 3336 32460
rect 3290 32392 3336 32424
rect 3290 32352 3296 32392
rect 3330 32352 3336 32392
rect 3290 32324 3336 32352
rect 3290 32280 3296 32324
rect 3330 32280 3336 32324
rect 3290 32256 3336 32280
rect 3290 32208 3296 32256
rect 3330 32208 3336 32256
rect 3290 32188 3336 32208
rect 3290 32136 3296 32188
rect 3330 32136 3336 32188
rect 3290 32120 3336 32136
rect 3290 32064 3296 32120
rect 3330 32064 3336 32120
rect 3290 32052 3336 32064
rect 3290 31992 3296 32052
rect 3330 31992 3336 32052
rect 3290 31984 3336 31992
rect 3290 31920 3296 31984
rect 3330 31920 3336 31984
rect 3290 31916 3336 31920
rect 3290 31814 3296 31916
rect 3330 31814 3336 31916
rect 3290 31810 3336 31814
rect 3290 31746 3296 31810
rect 3330 31746 3336 31810
rect 3290 31738 3336 31746
rect 3290 31678 3296 31738
rect 3330 31678 3336 31738
rect 3290 31666 3336 31678
rect 3290 31610 3296 31666
rect 3330 31610 3336 31666
rect 3290 31594 3336 31610
rect 3290 31542 3296 31594
rect 3330 31542 3336 31594
rect 3290 31522 3336 31542
rect 3290 31474 3296 31522
rect 3330 31474 3336 31522
rect 3290 31450 3336 31474
rect 3290 31406 3296 31450
rect 3330 31406 3336 31450
rect 3290 31378 3336 31406
rect 3290 31338 3296 31378
rect 3330 31338 3336 31378
rect 3290 31306 3336 31338
rect 3290 31270 3296 31306
rect 3330 31270 3336 31306
rect 3290 31236 3336 31270
rect 3290 31200 3296 31236
rect 3330 31200 3336 31236
rect 3290 31168 3336 31200
rect 3290 31128 3296 31168
rect 3330 31128 3336 31168
rect 3290 31100 3336 31128
rect 3290 31056 3296 31100
rect 3330 31056 3336 31100
rect 3290 31032 3336 31056
rect 3290 30984 3296 31032
rect 3330 30984 3336 31032
rect 3290 30964 3336 30984
rect 3290 30912 3296 30964
rect 3330 30912 3336 30964
rect 3290 30896 3336 30912
rect 3290 30840 3296 30896
rect 3330 30840 3336 30896
rect 3290 30828 3336 30840
rect 3290 30768 3296 30828
rect 3330 30768 3336 30828
rect 3290 30760 3336 30768
rect 3290 30696 3296 30760
rect 3330 30696 3336 30760
rect 3290 30692 3336 30696
rect 3290 30590 3296 30692
rect 3330 30590 3336 30692
rect 3290 30586 3336 30590
rect 3290 30522 3296 30586
rect 3330 30522 3336 30586
rect 3290 30514 3336 30522
rect 3290 30454 3296 30514
rect 3330 30454 3336 30514
rect 3290 30442 3336 30454
rect 3290 30386 3296 30442
rect 3330 30386 3336 30442
rect 3290 30370 3336 30386
rect 3290 30318 3296 30370
rect 3330 30318 3336 30370
rect 3290 30298 3336 30318
rect 3290 30250 3296 30298
rect 3330 30250 3336 30298
rect 3290 30226 3336 30250
rect 3290 30182 3296 30226
rect 3330 30182 3336 30226
rect 3290 30154 3336 30182
rect 3290 30114 3296 30154
rect 3330 30114 3336 30154
rect 3290 30082 3336 30114
rect 3290 30046 3296 30082
rect 3330 30046 3336 30082
rect 3290 30012 3336 30046
rect 3290 29976 3296 30012
rect 3330 29976 3336 30012
rect 3290 29944 3336 29976
rect 3290 29904 3296 29944
rect 3330 29904 3336 29944
rect 3290 29876 3336 29904
rect 3290 29832 3296 29876
rect 3330 29832 3336 29876
rect 3290 29808 3336 29832
rect 3290 29760 3296 29808
rect 3330 29760 3336 29808
rect 3290 29740 3336 29760
rect 3290 29688 3296 29740
rect 3330 29688 3336 29740
rect 3290 29672 3336 29688
rect 3290 29616 3296 29672
rect 3330 29616 3336 29672
rect 3290 29604 3336 29616
rect 3290 29544 3296 29604
rect 3330 29544 3336 29604
rect 3290 29536 3336 29544
rect 3290 29472 3296 29536
rect 3330 29472 3336 29536
rect 3290 29468 3336 29472
rect 3290 29366 3296 29468
rect 3330 29366 3336 29468
rect 3290 29362 3336 29366
rect 3290 29298 3296 29362
rect 3330 29298 3336 29362
rect 3290 29290 3336 29298
rect 3290 29230 3296 29290
rect 3330 29230 3336 29290
rect 3290 29218 3336 29230
rect 3290 29162 3296 29218
rect 3330 29162 3336 29218
rect 3290 29146 3336 29162
rect 3290 29094 3296 29146
rect 3330 29094 3336 29146
rect 3290 29074 3336 29094
rect 3290 29026 3296 29074
rect 3330 29026 3336 29074
rect 3290 29002 3336 29026
rect 3290 28958 3296 29002
rect 3330 28958 3336 29002
rect 3290 28930 3336 28958
rect 3290 28890 3296 28930
rect 3330 28890 3336 28930
rect 3290 28858 3336 28890
rect 3290 28822 3296 28858
rect 3330 28822 3336 28858
rect 3290 28788 3336 28822
rect 3290 28752 3296 28788
rect 3330 28752 3336 28788
rect 3290 28720 3336 28752
rect 3290 28680 3296 28720
rect 3330 28680 3336 28720
rect 3290 28652 3336 28680
rect 3290 28608 3296 28652
rect 3330 28608 3336 28652
rect 3290 28584 3336 28608
rect 3290 28536 3296 28584
rect 3330 28536 3336 28584
rect 3290 28516 3336 28536
rect 3290 28464 3296 28516
rect 3330 28464 3336 28516
rect 3290 28448 3336 28464
rect 3290 28392 3296 28448
rect 3330 28392 3336 28448
rect 3290 28380 3336 28392
rect 3290 28320 3296 28380
rect 3330 28320 3336 28380
rect 3290 28312 3336 28320
rect 3290 28248 3296 28312
rect 3330 28248 3336 28312
rect 3290 28244 3336 28248
rect 3290 28142 3296 28244
rect 3330 28142 3336 28244
rect 3290 28138 3336 28142
rect 3290 28074 3296 28138
rect 3330 28074 3336 28138
rect 3290 28066 3336 28074
rect 3290 28006 3296 28066
rect 3330 28006 3336 28066
rect 3290 27994 3336 28006
rect 3290 27938 3296 27994
rect 3330 27938 3336 27994
rect 3290 27922 3336 27938
rect 3290 27870 3296 27922
rect 3330 27870 3336 27922
rect 3290 27850 3336 27870
rect 3290 27802 3296 27850
rect 3330 27802 3336 27850
rect 3290 27778 3336 27802
rect 3290 27734 3296 27778
rect 3330 27734 3336 27778
rect 3290 27706 3336 27734
rect 3290 27666 3296 27706
rect 3330 27666 3336 27706
rect 3290 27634 3336 27666
rect 3290 27598 3296 27634
rect 3330 27598 3336 27634
rect 3290 27564 3336 27598
rect 3290 27528 3296 27564
rect 3330 27528 3336 27564
rect 3290 27496 3336 27528
rect 3290 27456 3296 27496
rect 3330 27456 3336 27496
rect 3290 27428 3336 27456
rect 3290 27384 3296 27428
rect 3330 27384 3336 27428
rect 3290 27360 3336 27384
rect 3290 27312 3296 27360
rect 3330 27312 3336 27360
rect 3290 27292 3336 27312
rect 3290 27240 3296 27292
rect 3330 27240 3336 27292
rect 3290 27224 3336 27240
rect 3290 27168 3296 27224
rect 3330 27168 3336 27224
rect 3290 27156 3336 27168
rect 3290 27096 3296 27156
rect 3330 27096 3336 27156
rect 3290 27088 3336 27096
rect 3290 27024 3296 27088
rect 3330 27024 3336 27088
rect 3290 27020 3336 27024
rect 3290 26918 3296 27020
rect 3330 26918 3336 27020
rect 3290 26914 3336 26918
rect 3290 26850 3296 26914
rect 3330 26850 3336 26914
rect 3290 26842 3336 26850
rect 3290 26782 3296 26842
rect 3330 26782 3336 26842
rect 3290 26770 3336 26782
rect 3290 26714 3296 26770
rect 3330 26714 3336 26770
rect 3290 26698 3336 26714
rect 3290 26646 3296 26698
rect 3330 26646 3336 26698
rect 3290 26626 3336 26646
rect 3290 26578 3296 26626
rect 3330 26578 3336 26626
rect 3290 26554 3336 26578
rect 3290 26510 3296 26554
rect 3330 26510 3336 26554
rect 3290 26482 3336 26510
rect 3290 26442 3296 26482
rect 3330 26442 3336 26482
rect 3290 26410 3336 26442
rect 3290 26374 3296 26410
rect 3330 26374 3336 26410
rect 3290 26340 3336 26374
rect 3290 26304 3296 26340
rect 3330 26304 3336 26340
rect 3290 26272 3336 26304
rect 3290 26232 3296 26272
rect 3330 26232 3336 26272
rect 3290 26204 3336 26232
rect 3290 26160 3296 26204
rect 3330 26160 3336 26204
rect 3290 26136 3336 26160
rect 3290 26088 3296 26136
rect 3330 26088 3336 26136
rect 3290 26068 3336 26088
rect 3290 26016 3296 26068
rect 3330 26016 3336 26068
rect 3290 26000 3336 26016
rect 3290 25944 3296 26000
rect 3330 25944 3336 26000
rect 3290 25932 3336 25944
rect 3290 25872 3296 25932
rect 3330 25872 3336 25932
rect 3290 25864 3336 25872
rect 3290 25800 3296 25864
rect 3330 25800 3336 25864
rect 3290 25796 3336 25800
rect 3290 25694 3296 25796
rect 3330 25694 3336 25796
rect 3290 25690 3336 25694
rect 3290 25626 3296 25690
rect 3330 25626 3336 25690
rect 3290 25618 3336 25626
rect 3290 25558 3296 25618
rect 3330 25558 3336 25618
rect 3290 25546 3336 25558
rect 3290 25490 3296 25546
rect 3330 25490 3336 25546
rect 3290 25474 3336 25490
rect 3290 25422 3296 25474
rect 3330 25422 3336 25474
rect 3290 25402 3336 25422
rect 3290 25354 3296 25402
rect 3330 25354 3336 25402
rect 3290 25330 3336 25354
rect 3290 25286 3296 25330
rect 3330 25286 3336 25330
rect 3290 25258 3336 25286
rect 3290 25218 3296 25258
rect 3330 25218 3336 25258
rect 3290 25186 3336 25218
rect 3290 25150 3296 25186
rect 3330 25150 3336 25186
rect 3290 25116 3336 25150
rect 3290 25080 3296 25116
rect 3330 25080 3336 25116
rect 3290 25048 3336 25080
rect 3290 25008 3296 25048
rect 3330 25008 3336 25048
rect 3290 24980 3336 25008
rect 3290 24936 3296 24980
rect 3330 24936 3336 24980
rect 3290 24912 3336 24936
rect 3290 24864 3296 24912
rect 3330 24864 3336 24912
rect 3290 24844 3336 24864
rect 3290 24792 3296 24844
rect 3330 24792 3336 24844
rect 3290 24776 3336 24792
rect 3290 24720 3296 24776
rect 3330 24720 3336 24776
rect 3290 24708 3336 24720
rect 3290 24648 3296 24708
rect 3330 24648 3336 24708
rect 3290 24640 3336 24648
rect 3290 24576 3296 24640
rect 3330 24576 3336 24640
rect 3290 24572 3336 24576
rect 3290 24470 3296 24572
rect 3330 24470 3336 24572
rect 3290 24466 3336 24470
rect 3290 24402 3296 24466
rect 3330 24402 3336 24466
rect 3290 24394 3336 24402
rect 3290 24334 3296 24394
rect 3330 24334 3336 24394
rect 3290 24322 3336 24334
rect 3290 24266 3296 24322
rect 3330 24266 3336 24322
rect 3290 24250 3336 24266
rect 3290 24198 3296 24250
rect 3330 24198 3336 24250
rect 3290 24178 3336 24198
rect 3290 24130 3296 24178
rect 3330 24130 3336 24178
rect 3290 24106 3336 24130
rect 3290 24062 3296 24106
rect 3330 24062 3336 24106
rect 3290 24034 3336 24062
rect 3290 23994 3296 24034
rect 3330 23994 3336 24034
rect 3290 23962 3336 23994
rect 3290 23926 3296 23962
rect 3330 23926 3336 23962
rect 3290 23892 3336 23926
rect 3290 23856 3296 23892
rect 3330 23856 3336 23892
rect 3290 23824 3336 23856
rect 3290 23784 3296 23824
rect 3330 23784 3336 23824
rect 3290 23756 3336 23784
rect 3290 23712 3296 23756
rect 3330 23712 3336 23756
rect 3290 23688 3336 23712
rect 3290 23640 3296 23688
rect 3330 23640 3336 23688
rect 3290 23620 3336 23640
rect 3290 23568 3296 23620
rect 3330 23568 3336 23620
rect 3290 23552 3336 23568
rect 3290 23496 3296 23552
rect 3330 23496 3336 23552
rect 3290 23484 3336 23496
rect 3290 23424 3296 23484
rect 3330 23424 3336 23484
rect 3290 23416 3336 23424
rect 3290 23352 3296 23416
rect 3330 23352 3336 23416
rect 3290 23348 3336 23352
rect 3290 23246 3296 23348
rect 3330 23246 3336 23348
rect 3290 23242 3336 23246
rect 3290 23178 3296 23242
rect 3330 23178 3336 23242
rect 3290 23170 3336 23178
rect 3290 23110 3296 23170
rect 3330 23110 3336 23170
rect 3290 23098 3336 23110
rect 3290 23042 3296 23098
rect 3330 23042 3336 23098
rect 3290 23026 3336 23042
rect 3290 22974 3296 23026
rect 3330 22974 3336 23026
rect 3290 22954 3336 22974
rect 3290 22906 3296 22954
rect 3330 22906 3336 22954
rect 3290 22882 3336 22906
rect 3290 22838 3296 22882
rect 3330 22838 3336 22882
rect 3290 22810 3336 22838
rect 3290 22770 3296 22810
rect 3330 22770 3336 22810
rect 3290 22738 3336 22770
rect 3290 22702 3296 22738
rect 3330 22702 3336 22738
rect 3290 22668 3336 22702
rect 3290 22632 3296 22668
rect 3330 22632 3336 22668
rect 3290 22600 3336 22632
rect 3290 22560 3296 22600
rect 3330 22560 3336 22600
rect 3290 22532 3336 22560
rect 3290 22488 3296 22532
rect 3330 22488 3336 22532
rect 3290 22464 3336 22488
rect 3290 22416 3296 22464
rect 3330 22416 3336 22464
rect 3290 22396 3336 22416
rect 3290 22344 3296 22396
rect 3330 22344 3336 22396
rect 3290 22328 3336 22344
rect 3290 22272 3296 22328
rect 3330 22272 3336 22328
rect 3290 22260 3336 22272
rect 3290 22200 3296 22260
rect 3330 22200 3336 22260
rect 3290 22192 3336 22200
rect 3290 22128 3296 22192
rect 3330 22128 3336 22192
rect 3290 22124 3336 22128
rect 3290 22022 3296 22124
rect 3330 22022 3336 22124
rect 3290 22018 3336 22022
rect 3290 21954 3296 22018
rect 3330 21954 3336 22018
rect 3290 21946 3336 21954
rect 3290 21886 3296 21946
rect 3330 21886 3336 21946
rect 3290 21874 3336 21886
rect 3290 21818 3296 21874
rect 3330 21818 3336 21874
rect 3290 21802 3336 21818
rect 3290 21750 3296 21802
rect 3330 21750 3336 21802
rect 3290 21730 3336 21750
rect 3290 21682 3296 21730
rect 3330 21682 3336 21730
rect 3290 21658 3336 21682
rect 3290 21614 3296 21658
rect 3330 21614 3336 21658
rect 3290 21586 3336 21614
rect 3290 21546 3296 21586
rect 3330 21546 3336 21586
rect 3290 21514 3336 21546
rect 3290 21478 3296 21514
rect 3330 21478 3336 21514
rect 3290 21444 3336 21478
rect 3290 21408 3296 21444
rect 3330 21408 3336 21444
rect 3290 21376 3336 21408
rect 3290 21336 3296 21376
rect 3330 21336 3336 21376
rect 3290 21308 3336 21336
rect 3290 21264 3296 21308
rect 3330 21264 3336 21308
rect 3290 21240 3336 21264
rect 3290 21192 3296 21240
rect 3330 21192 3336 21240
rect 3290 21172 3336 21192
rect 3290 21120 3296 21172
rect 3330 21120 3336 21172
rect 3290 21104 3336 21120
rect 3290 21048 3296 21104
rect 3330 21048 3336 21104
rect 3290 21036 3336 21048
rect 3290 20976 3296 21036
rect 3330 20976 3336 21036
rect 3290 20968 3336 20976
rect 3290 20904 3296 20968
rect 3330 20904 3336 20968
rect 3290 20900 3336 20904
rect 3290 20798 3296 20900
rect 3330 20798 3336 20900
rect 3290 20794 3336 20798
rect 3290 20730 3296 20794
rect 3330 20730 3336 20794
rect 3290 20722 3336 20730
rect 3290 20662 3296 20722
rect 3330 20662 3336 20722
rect 3290 20650 3336 20662
rect 3290 20594 3296 20650
rect 3330 20594 3336 20650
rect 3290 20578 3336 20594
rect 3290 20526 3296 20578
rect 3330 20526 3336 20578
rect 3290 20506 3336 20526
rect 3290 20458 3296 20506
rect 3330 20458 3336 20506
rect 3290 20434 3336 20458
rect 3290 20390 3296 20434
rect 3330 20390 3336 20434
rect 3290 20362 3336 20390
rect 3290 20322 3296 20362
rect 3330 20322 3336 20362
rect 3290 20290 3336 20322
rect 3290 20254 3296 20290
rect 3330 20254 3336 20290
rect 3290 20220 3336 20254
rect 3290 20184 3296 20220
rect 3330 20184 3336 20220
rect 3290 20152 3336 20184
rect 3290 20112 3296 20152
rect 3330 20112 3336 20152
rect 3290 20084 3336 20112
rect 3290 20040 3296 20084
rect 3330 20040 3336 20084
rect 3290 20016 3336 20040
rect 3290 19968 3296 20016
rect 3330 19968 3336 20016
rect 3290 19948 3336 19968
rect 3290 19896 3296 19948
rect 3330 19896 3336 19948
rect 3290 19880 3336 19896
rect 3290 19824 3296 19880
rect 3330 19824 3336 19880
rect 3290 19812 3336 19824
rect 3290 19752 3296 19812
rect 3330 19752 3336 19812
rect 3290 19744 3336 19752
rect 3290 19680 3296 19744
rect 3330 19680 3336 19744
rect 3290 19676 3336 19680
rect 3290 19574 3296 19676
rect 3330 19574 3336 19676
rect 3290 19570 3336 19574
rect 3290 19506 3296 19570
rect 3330 19506 3336 19570
rect 3290 19498 3336 19506
rect 3290 19438 3296 19498
rect 3330 19438 3336 19498
rect 3290 19426 3336 19438
rect 3290 19370 3296 19426
rect 3330 19370 3336 19426
rect 3290 19354 3336 19370
rect 3290 19302 3296 19354
rect 3330 19302 3336 19354
rect 3290 19282 3336 19302
rect 3290 19234 3296 19282
rect 3330 19234 3336 19282
rect 3290 19210 3336 19234
rect 3290 19166 3296 19210
rect 3330 19166 3336 19210
rect 3290 19138 3336 19166
rect 3290 19098 3296 19138
rect 3330 19098 3336 19138
rect 3290 19066 3336 19098
rect 3290 19030 3296 19066
rect 3330 19030 3336 19066
rect 3290 18996 3336 19030
rect 3290 18960 3296 18996
rect 3330 18960 3336 18996
rect 3290 18928 3336 18960
rect 3290 18888 3296 18928
rect 3330 18888 3336 18928
rect 3290 18860 3336 18888
rect 3290 18816 3296 18860
rect 3330 18816 3336 18860
rect 3290 18792 3336 18816
rect 3290 18744 3296 18792
rect 3330 18744 3336 18792
rect 3290 18724 3336 18744
rect 3290 18672 3296 18724
rect 3330 18672 3336 18724
rect 3290 18656 3336 18672
rect 3290 18600 3296 18656
rect 3330 18600 3336 18656
rect 3290 18588 3336 18600
rect 3290 18528 3296 18588
rect 3330 18528 3336 18588
rect 3290 18520 3336 18528
rect 3290 18456 3296 18520
rect 3330 18456 3336 18520
rect 3290 18452 3336 18456
rect 3290 18350 3296 18452
rect 3330 18350 3336 18452
rect 3290 18346 3336 18350
rect 3290 18282 3296 18346
rect 3330 18282 3336 18346
rect 3290 18274 3336 18282
rect 3290 18214 3296 18274
rect 3330 18214 3336 18274
rect 3290 18202 3336 18214
rect 3290 18146 3296 18202
rect 3330 18146 3336 18202
rect 3290 18130 3336 18146
rect 3290 18078 3296 18130
rect 3330 18078 3336 18130
rect 3290 18058 3336 18078
rect 3290 18010 3296 18058
rect 3330 18010 3336 18058
rect 3290 17986 3336 18010
rect 3290 17942 3296 17986
rect 3330 17942 3336 17986
rect 3290 17914 3336 17942
rect 3290 17874 3296 17914
rect 3330 17874 3336 17914
rect 3290 17842 3336 17874
rect 3290 17806 3296 17842
rect 3330 17806 3336 17842
rect 3290 17772 3336 17806
rect 3290 17736 3296 17772
rect 3330 17736 3336 17772
rect 3290 17704 3336 17736
rect 3290 17664 3296 17704
rect 3330 17664 3336 17704
rect 3290 17636 3336 17664
rect 3290 17592 3296 17636
rect 3330 17592 3336 17636
rect 3290 17568 3336 17592
rect 3290 17520 3296 17568
rect 3330 17520 3336 17568
rect 3290 17500 3336 17520
rect 3290 17448 3296 17500
rect 3330 17448 3336 17500
rect 3290 17432 3336 17448
rect 3290 17376 3296 17432
rect 3330 17376 3336 17432
rect 3290 17364 3336 17376
rect 3290 17304 3296 17364
rect 3330 17304 3336 17364
rect 3290 17296 3336 17304
rect 3290 17232 3296 17296
rect 3330 17232 3336 17296
rect 3290 17228 3336 17232
rect 3290 17126 3296 17228
rect 3330 17126 3336 17228
rect 3290 17122 3336 17126
rect 3290 17058 3296 17122
rect 3330 17058 3336 17122
rect 3290 17050 3336 17058
rect 3290 16990 3296 17050
rect 3330 16990 3336 17050
rect 3290 16978 3336 16990
rect 3290 16922 3296 16978
rect 3330 16922 3336 16978
rect 3290 16906 3336 16922
rect 3290 16854 3296 16906
rect 3330 16854 3336 16906
rect 3290 16834 3336 16854
rect 3290 16786 3296 16834
rect 3330 16786 3336 16834
rect 3290 16762 3336 16786
rect 3290 16718 3296 16762
rect 3330 16718 3336 16762
rect 3290 16690 3336 16718
rect 3290 16650 3296 16690
rect 3330 16650 3336 16690
rect 3290 16618 3336 16650
rect 3290 16582 3296 16618
rect 3330 16582 3336 16618
rect 3290 16548 3336 16582
rect 3290 16512 3296 16548
rect 3330 16512 3336 16548
rect 3290 16480 3336 16512
rect 3290 16440 3296 16480
rect 3330 16440 3336 16480
rect 3290 16412 3336 16440
rect 3290 16368 3296 16412
rect 3330 16368 3336 16412
rect 3290 16344 3336 16368
rect 3290 16296 3296 16344
rect 3330 16296 3336 16344
rect 3290 16276 3336 16296
rect 3290 16224 3296 16276
rect 3330 16224 3336 16276
rect 3290 16208 3336 16224
rect 3290 16152 3296 16208
rect 3330 16152 3336 16208
rect 3290 16140 3336 16152
rect 3290 16080 3296 16140
rect 3330 16080 3336 16140
rect 3290 16072 3336 16080
rect 3290 16008 3296 16072
rect 3330 16008 3336 16072
rect 3290 16004 3336 16008
rect 3290 15902 3296 16004
rect 3330 15902 3336 16004
rect 3290 15898 3336 15902
rect 3290 15834 3296 15898
rect 3330 15834 3336 15898
rect 3290 15826 3336 15834
rect 3290 15766 3296 15826
rect 3330 15766 3336 15826
rect 3290 15754 3336 15766
rect 3290 15698 3296 15754
rect 3330 15698 3336 15754
rect 3290 15682 3336 15698
rect 3290 15630 3296 15682
rect 3330 15630 3336 15682
rect 3290 15610 3336 15630
rect 3290 15562 3296 15610
rect 3330 15562 3336 15610
rect 3290 15538 3336 15562
rect 3290 15494 3296 15538
rect 3330 15494 3336 15538
rect 3290 15466 3336 15494
rect 3290 15426 3296 15466
rect 3330 15426 3336 15466
rect 3290 15394 3336 15426
rect 3290 15358 3296 15394
rect 3330 15358 3336 15394
rect 3290 15324 3336 15358
rect 3290 15288 3296 15324
rect 3330 15288 3336 15324
rect 3290 15256 3336 15288
rect 3290 15216 3296 15256
rect 3330 15216 3336 15256
rect 3290 15188 3336 15216
rect 3290 15144 3296 15188
rect 3330 15144 3336 15188
rect 3290 15120 3336 15144
rect 3290 15072 3296 15120
rect 3330 15072 3336 15120
rect 3290 15052 3336 15072
rect 3290 15000 3296 15052
rect 3330 15000 3336 15052
rect 3290 14984 3336 15000
rect 3290 14928 3296 14984
rect 3330 14928 3336 14984
rect 3290 14916 3336 14928
rect 3290 14856 3296 14916
rect 3330 14856 3336 14916
rect 3290 14848 3336 14856
rect 3290 14784 3296 14848
rect 3330 14784 3336 14848
rect 3290 14780 3336 14784
rect 3290 14678 3296 14780
rect 3330 14678 3336 14780
rect 3290 14674 3336 14678
rect 3290 14610 3296 14674
rect 3330 14610 3336 14674
rect 3290 14602 3336 14610
rect 3290 14542 3296 14602
rect 3330 14542 3336 14602
rect 3290 14530 3336 14542
rect 3290 14474 3296 14530
rect 3330 14474 3336 14530
rect 3290 14458 3336 14474
rect 3290 14406 3296 14458
rect 3330 14406 3336 14458
rect 3290 14386 3336 14406
rect 3290 14338 3296 14386
rect 3330 14338 3336 14386
rect 3290 14314 3336 14338
rect 3290 14270 3296 14314
rect 3330 14270 3336 14314
rect 3290 14242 3336 14270
rect 3290 14202 3296 14242
rect 3330 14202 3336 14242
rect 3290 14170 3336 14202
rect 3290 14134 3296 14170
rect 3330 14134 3336 14170
rect 3290 14100 3336 14134
rect 3290 14064 3296 14100
rect 3330 14064 3336 14100
rect 3290 14032 3336 14064
rect 3290 13992 3296 14032
rect 3330 13992 3336 14032
rect 3290 13964 3336 13992
rect 3290 13920 3296 13964
rect 3330 13920 3336 13964
rect 3290 13896 3336 13920
rect 3290 13848 3296 13896
rect 3330 13848 3336 13896
rect 3290 13828 3336 13848
rect 3290 13776 3296 13828
rect 3330 13776 3336 13828
rect 3290 13760 3336 13776
rect 3290 13704 3296 13760
rect 3330 13704 3336 13760
rect 3290 13692 3336 13704
rect 3290 13632 3296 13692
rect 3330 13632 3336 13692
rect 3290 13624 3336 13632
rect 3290 13560 3296 13624
rect 3330 13560 3336 13624
rect 3290 13556 3336 13560
rect 3290 13454 3296 13556
rect 3330 13454 3336 13556
rect 3290 13450 3336 13454
rect 3290 13386 3296 13450
rect 3330 13386 3336 13450
rect 3290 13378 3336 13386
rect 3290 13318 3296 13378
rect 3330 13318 3336 13378
rect 3290 13306 3336 13318
rect 3290 13250 3296 13306
rect 3330 13250 3336 13306
rect 3290 13234 3336 13250
rect 3290 13182 3296 13234
rect 3330 13182 3336 13234
rect 3290 13162 3336 13182
rect 3290 13114 3296 13162
rect 3330 13114 3336 13162
rect 3290 13090 3336 13114
rect 3290 13046 3296 13090
rect 3330 13046 3336 13090
rect 3290 13018 3336 13046
rect 3290 12978 3296 13018
rect 3330 12978 3336 13018
rect 3290 12946 3336 12978
rect 3290 12910 3296 12946
rect 3330 12910 3336 12946
rect 3290 12876 3336 12910
rect 3290 12840 3296 12876
rect 3330 12840 3336 12876
rect 3290 12808 3336 12840
rect 3290 12768 3296 12808
rect 3330 12768 3336 12808
rect 3290 12740 3336 12768
rect 3290 12696 3296 12740
rect 3330 12696 3336 12740
rect 3290 12672 3336 12696
rect 3290 12624 3296 12672
rect 3330 12624 3336 12672
rect 3290 12604 3336 12624
rect 3290 12552 3296 12604
rect 3330 12552 3336 12604
rect 3290 12536 3336 12552
rect 3290 12480 3296 12536
rect 3330 12480 3336 12536
rect 3290 12468 3336 12480
rect 3290 12408 3296 12468
rect 3330 12408 3336 12468
rect 3290 12400 3336 12408
rect 3290 12336 3296 12400
rect 3330 12336 3336 12400
rect 3290 12332 3336 12336
rect 3290 12230 3296 12332
rect 3330 12230 3336 12332
rect 3290 12226 3336 12230
rect 3290 12162 3296 12226
rect 3330 12162 3336 12226
rect 3290 12154 3336 12162
rect 3290 12094 3296 12154
rect 3330 12094 3336 12154
rect 3290 12082 3336 12094
rect 3290 12026 3296 12082
rect 3330 12026 3336 12082
rect 3290 12010 3336 12026
rect 3290 11958 3296 12010
rect 3330 11958 3336 12010
rect 3290 11938 3336 11958
rect 3290 11890 3296 11938
rect 3330 11890 3336 11938
rect 3290 11866 3336 11890
rect 3290 11822 3296 11866
rect 3330 11822 3336 11866
rect 3290 11794 3336 11822
rect 3290 11754 3296 11794
rect 3330 11754 3336 11794
rect 3290 11722 3336 11754
rect 3290 11686 3296 11722
rect 3330 11686 3336 11722
rect 3290 11652 3336 11686
rect 3290 11616 3296 11652
rect 3330 11616 3336 11652
rect 3290 11584 3336 11616
rect 3290 11544 3296 11584
rect 3330 11544 3336 11584
rect 3290 11516 3336 11544
rect 3290 11472 3296 11516
rect 3330 11472 3336 11516
rect 3290 11448 3336 11472
rect 3290 11400 3296 11448
rect 3330 11400 3336 11448
rect 3290 11380 3336 11400
rect 3290 11328 3296 11380
rect 3330 11328 3336 11380
rect 3290 11312 3336 11328
rect 3290 11256 3296 11312
rect 3330 11256 3336 11312
rect 3290 11244 3336 11256
rect 3290 11184 3296 11244
rect 3330 11184 3336 11244
rect 3290 11176 3336 11184
rect 3290 11112 3296 11176
rect 3330 11112 3336 11176
rect 3290 11108 3336 11112
rect 3290 11006 3296 11108
rect 3330 11006 3336 11108
rect 3290 11002 3336 11006
rect 3290 10938 3296 11002
rect 3330 10938 3336 11002
rect 3290 10930 3336 10938
rect 3290 10870 3296 10930
rect 3330 10870 3336 10930
rect 3290 10858 3336 10870
rect 3290 10802 3296 10858
rect 3330 10802 3336 10858
rect 3290 10786 3336 10802
rect 3290 10734 3296 10786
rect 3330 10734 3336 10786
rect 3290 10714 3336 10734
rect 3290 10666 3296 10714
rect 3330 10666 3336 10714
rect 3290 10642 3336 10666
rect 3290 10598 3296 10642
rect 3330 10598 3336 10642
rect 3290 10570 3336 10598
rect 3290 10530 3296 10570
rect 3330 10530 3336 10570
rect 3290 10498 3336 10530
rect 3290 10462 3296 10498
rect 3330 10462 3336 10498
rect 3290 10428 3336 10462
rect 3290 10392 3296 10428
rect 3330 10392 3336 10428
rect 3290 10360 3336 10392
rect 3290 10320 3296 10360
rect 3330 10320 3336 10360
rect 3290 10292 3336 10320
rect 3290 10248 3296 10292
rect 3330 10248 3336 10292
rect 3290 10224 3336 10248
rect 3290 10176 3296 10224
rect 3330 10176 3336 10224
rect 3290 10156 3336 10176
rect 3290 10104 3296 10156
rect 3330 10104 3336 10156
rect 3290 10088 3336 10104
rect 3290 10032 3296 10088
rect 3330 10032 3336 10088
rect 3290 10020 3336 10032
rect 3290 9960 3296 10020
rect 3330 9960 3336 10020
rect 3290 9952 3336 9960
rect 3290 9888 3296 9952
rect 3330 9888 3336 9952
rect 3290 9884 3336 9888
rect 3290 9782 3296 9884
rect 3330 9782 3336 9884
rect 3290 9778 3336 9782
rect 3290 9714 3296 9778
rect 3330 9714 3336 9778
rect 3290 9706 3336 9714
rect 3290 9646 3296 9706
rect 3330 9646 3336 9706
rect 3290 9634 3336 9646
rect 3290 9578 3296 9634
rect 3330 9578 3336 9634
rect 3290 9562 3336 9578
rect 3290 9510 3296 9562
rect 3330 9510 3336 9562
rect 3290 9490 3336 9510
rect 3290 9442 3296 9490
rect 3330 9442 3336 9490
rect 3290 9418 3336 9442
rect 3290 9374 3296 9418
rect 3330 9374 3336 9418
rect 3290 9346 3336 9374
rect 3290 9306 3296 9346
rect 3330 9306 3336 9346
rect 3290 9274 3336 9306
rect 3290 9238 3296 9274
rect 3330 9238 3336 9274
rect 3290 9204 3336 9238
rect 3290 9168 3296 9204
rect 3330 9168 3336 9204
rect 3290 9136 3336 9168
rect 3290 9096 3296 9136
rect 3330 9096 3336 9136
rect 3290 9068 3336 9096
rect 3290 9024 3296 9068
rect 3330 9024 3336 9068
rect 3290 9000 3336 9024
rect 3290 8952 3296 9000
rect 3330 8952 3336 9000
rect 3290 8932 3336 8952
rect 3290 8880 3296 8932
rect 3330 8880 3336 8932
rect 3290 8864 3336 8880
rect 3290 8808 3296 8864
rect 3330 8808 3336 8864
rect 3290 8796 3336 8808
rect 3290 8736 3296 8796
rect 3330 8736 3336 8796
rect 3290 8728 3336 8736
rect 3290 8664 3296 8728
rect 3330 8664 3336 8728
rect 3290 8660 3336 8664
rect 3290 8558 3296 8660
rect 3330 8558 3336 8660
rect 3290 8554 3336 8558
rect 3290 8490 3296 8554
rect 3330 8490 3336 8554
rect 3290 8482 3336 8490
rect 3290 8422 3296 8482
rect 3330 8422 3336 8482
rect 3290 8410 3336 8422
rect 3290 8354 3296 8410
rect 3330 8354 3336 8410
rect 3290 8338 3336 8354
rect 3290 8286 3296 8338
rect 3330 8286 3336 8338
rect 3290 8266 3336 8286
rect 3290 8218 3296 8266
rect 3330 8218 3336 8266
rect 3290 8194 3336 8218
rect 3290 8150 3296 8194
rect 3330 8150 3336 8194
rect 3290 8122 3336 8150
rect 3290 8082 3296 8122
rect 3330 8082 3336 8122
rect 3290 8050 3336 8082
rect 3290 8014 3296 8050
rect 3330 8014 3336 8050
rect 3290 7980 3336 8014
rect 3290 7944 3296 7980
rect 3330 7944 3336 7980
rect 3290 7912 3336 7944
rect 3290 7872 3296 7912
rect 3330 7872 3336 7912
rect 3290 7844 3336 7872
rect 3290 7800 3296 7844
rect 3330 7800 3336 7844
rect 3290 7776 3336 7800
rect 3290 7728 3296 7776
rect 3330 7728 3336 7776
rect 3290 7708 3336 7728
rect 3290 7656 3296 7708
rect 3330 7656 3336 7708
rect 3290 7640 3336 7656
rect 3290 7584 3296 7640
rect 3330 7584 3336 7640
rect 3290 7572 3336 7584
rect 3290 7512 3296 7572
rect 3330 7512 3336 7572
rect 3290 7504 3336 7512
rect 3290 7440 3296 7504
rect 3330 7440 3336 7504
rect 3290 7436 3336 7440
rect 3290 7334 3296 7436
rect 3330 7334 3336 7436
rect 3290 7330 3336 7334
rect 3290 7266 3296 7330
rect 3330 7266 3336 7330
rect 3290 7258 3336 7266
rect 3290 7198 3296 7258
rect 3330 7198 3336 7258
rect 3290 7186 3336 7198
rect 3290 7130 3296 7186
rect 3330 7130 3336 7186
rect 3290 7114 3336 7130
rect 3290 7062 3296 7114
rect 3330 7062 3336 7114
rect 3290 7042 3336 7062
rect 3290 6994 3296 7042
rect 3330 6994 3336 7042
rect 3290 6970 3336 6994
rect 3290 6926 3296 6970
rect 3330 6926 3336 6970
rect 3290 6898 3336 6926
rect 3290 6858 3296 6898
rect 3330 6858 3336 6898
rect 3290 6826 3336 6858
rect 3290 6790 3296 6826
rect 3330 6790 3336 6826
rect 3290 6756 3336 6790
rect 3290 6720 3296 6756
rect 3330 6720 3336 6756
rect 3290 6688 3336 6720
rect 3290 6648 3296 6688
rect 3330 6648 3336 6688
rect 3290 6620 3336 6648
rect 3290 6576 3296 6620
rect 3330 6576 3336 6620
rect 3290 6552 3336 6576
rect 3290 6504 3296 6552
rect 3330 6504 3336 6552
rect 3290 6484 3336 6504
rect 3290 6432 3296 6484
rect 3330 6432 3336 6484
rect 3290 6416 3336 6432
rect 3290 6360 3296 6416
rect 3330 6360 3336 6416
rect 3290 6348 3336 6360
rect 3290 6288 3296 6348
rect 3330 6288 3336 6348
rect 3290 6280 3336 6288
rect 3290 6216 3296 6280
rect 3330 6216 3336 6280
rect 3290 6212 3336 6216
rect 3290 6110 3296 6212
rect 3330 6110 3336 6212
rect 3290 6106 3336 6110
rect 3290 6042 3296 6106
rect 3330 6042 3336 6106
rect 3290 6034 3336 6042
rect 3290 5974 3296 6034
rect 3330 5974 3336 6034
rect 3290 5962 3336 5974
rect 3290 5906 3296 5962
rect 3330 5906 3336 5962
rect 3290 5890 3336 5906
rect 3290 5838 3296 5890
rect 3330 5838 3336 5890
rect 3290 5818 3336 5838
rect 3290 5770 3296 5818
rect 3330 5770 3336 5818
rect 3290 5746 3336 5770
rect 3290 5702 3296 5746
rect 3330 5702 3336 5746
rect 3290 5674 3336 5702
rect 3290 5634 3296 5674
rect 3330 5634 3336 5674
rect 3290 5602 3336 5634
rect 3290 5566 3296 5602
rect 3330 5566 3336 5602
rect 3290 5532 3336 5566
rect 3290 5496 3296 5532
rect 3330 5496 3336 5532
rect 3290 5464 3336 5496
rect 3290 5424 3296 5464
rect 3330 5424 3336 5464
rect 3290 5396 3336 5424
rect 3290 5352 3296 5396
rect 3330 5352 3336 5396
rect 3290 5328 3336 5352
rect 3290 5280 3296 5328
rect 3330 5280 3336 5328
rect 3290 5260 3336 5280
rect 3290 5208 3296 5260
rect 3330 5208 3336 5260
rect 3290 5192 3336 5208
rect 3290 5136 3296 5192
rect 3330 5136 3336 5192
rect 3290 5124 3336 5136
rect 3290 5064 3296 5124
rect 3330 5064 3336 5124
rect 3290 5056 3336 5064
rect 3290 4992 3296 5056
rect 3330 4992 3336 5056
rect 3290 4988 3336 4992
rect 3290 4886 3296 4988
rect 3330 4886 3336 4988
rect 3290 4882 3336 4886
rect 3290 4818 3296 4882
rect 3330 4818 3336 4882
rect 3290 4810 3336 4818
rect 3290 4750 3296 4810
rect 3330 4750 3336 4810
rect 3290 4738 3336 4750
rect 3290 4682 3296 4738
rect 3330 4682 3336 4738
rect 3290 4666 3336 4682
rect 3290 4614 3296 4666
rect 3330 4614 3336 4666
rect 3290 4594 3336 4614
rect 3290 4546 3296 4594
rect 3330 4546 3336 4594
rect 3290 4522 3336 4546
rect 3290 4478 3296 4522
rect 3330 4478 3336 4522
rect 3290 4450 3336 4478
rect 3290 4410 3296 4450
rect 3330 4410 3336 4450
rect 3290 4378 3336 4410
rect 3290 4342 3296 4378
rect 3330 4342 3336 4378
rect 3290 4308 3336 4342
rect 3290 4272 3296 4308
rect 3330 4272 3336 4308
rect 3290 4240 3336 4272
rect 3290 4200 3296 4240
rect 3330 4200 3336 4240
rect 3290 4172 3336 4200
rect 3290 4128 3296 4172
rect 3330 4128 3336 4172
rect 3290 4104 3336 4128
rect 3290 4056 3296 4104
rect 3330 4056 3336 4104
rect 3290 4036 3336 4056
rect 3290 3984 3296 4036
rect 3330 3984 3336 4036
rect 3290 3968 3336 3984
rect 3290 3912 3296 3968
rect 3330 3912 3336 3968
rect 3290 3900 3336 3912
rect 3290 3840 3296 3900
rect 3330 3840 3336 3900
rect 3290 3832 3336 3840
rect 3290 3768 3296 3832
rect 3330 3768 3336 3832
rect 3290 3764 3336 3768
rect 3290 3662 3296 3764
rect 3330 3662 3336 3764
rect 3290 3658 3336 3662
rect 3290 3594 3296 3658
rect 3330 3594 3336 3658
rect 3290 3586 3336 3594
rect 3290 3526 3296 3586
rect 3330 3526 3336 3586
rect 3290 3514 3336 3526
rect 3290 3458 3296 3514
rect 3330 3458 3336 3514
rect 3290 3442 3336 3458
rect 3290 3390 3296 3442
rect 3330 3390 3336 3442
rect 3290 3370 3336 3390
rect 3290 3322 3296 3370
rect 3330 3322 3336 3370
rect 3290 3298 3336 3322
rect 3290 3254 3296 3298
rect 3330 3254 3336 3298
rect 3290 3225 3336 3254
rect 3290 3186 3296 3225
rect 3330 3186 3336 3225
rect 3290 3152 3336 3186
rect 3290 3118 3296 3152
rect 3330 3118 3336 3152
rect 3290 3084 3336 3118
rect 3290 3045 3296 3084
rect 3330 3045 3336 3084
rect 3290 3016 3336 3045
rect 3290 2972 3296 3016
rect 3330 2972 3336 3016
rect 3290 2948 3336 2972
rect 3290 2899 3296 2948
rect 3330 2899 3336 2948
rect 3290 2880 3336 2899
rect 3290 2826 3296 2880
rect 3330 2826 3336 2880
rect 3290 2812 3336 2826
rect 3290 2753 3296 2812
rect 3330 2753 3336 2812
rect 3290 2744 3336 2753
rect 3290 2680 3296 2744
rect 3330 2680 3336 2744
rect 3290 2676 3336 2680
rect 3290 2642 3296 2676
rect 3330 2642 3336 2676
rect 3290 2641 3336 2642
rect 3290 2574 3296 2641
rect 3330 2574 3336 2641
rect 3290 2568 3336 2574
rect 3290 2506 3296 2568
rect 3330 2506 3336 2568
rect 3290 2495 3336 2506
rect 3290 2438 3296 2495
rect 3330 2438 3336 2495
rect 3290 2422 3336 2438
rect 3290 2370 3296 2422
rect 3330 2370 3336 2422
rect 3290 2349 3336 2370
rect 3290 2302 3296 2349
rect 3330 2302 3336 2349
rect 3290 2276 3336 2302
rect 3290 2234 3296 2276
rect 3330 2234 3336 2276
rect 3290 2203 3336 2234
rect 3290 2166 3296 2203
rect 3330 2166 3336 2203
rect 3290 2132 3336 2166
rect 3290 2096 3296 2132
rect 3330 2096 3336 2132
rect 3290 2064 3336 2096
rect 3290 2023 3296 2064
rect 3330 2023 3336 2064
rect 3290 1996 3336 2023
rect 3290 1950 3296 1996
rect 3330 1950 3336 1996
rect 3290 1928 3336 1950
rect 3290 1877 3296 1928
rect 3330 1877 3336 1928
rect 3290 1860 3336 1877
rect 3290 1804 3296 1860
rect 3330 1804 3336 1860
rect 3290 1792 3336 1804
rect 3290 1731 3296 1792
rect 3330 1731 3336 1792
rect 3290 1724 3336 1731
rect 3290 1658 3296 1724
rect 3330 1658 3336 1724
rect 3290 1656 3336 1658
rect 3290 1622 3296 1656
rect 3330 1622 3336 1656
rect 3290 1619 3336 1622
rect 3290 1554 3296 1619
rect 3330 1554 3336 1619
rect 3290 1546 3336 1554
rect 3290 1486 3296 1546
rect 3330 1486 3336 1546
rect 3290 1473 3336 1486
rect 3290 1418 3296 1473
rect 3330 1418 3336 1473
rect 3290 1400 3336 1418
rect 3290 1350 3296 1400
rect 3330 1350 3336 1400
rect 3290 1327 3336 1350
rect 3290 1282 3296 1327
rect 3330 1282 3336 1327
rect 3290 1254 3336 1282
rect 3290 1214 3296 1254
rect 3330 1214 3336 1254
rect 3290 1181 3336 1214
rect 3290 1146 3296 1181
rect 3330 1146 3336 1181
rect 3290 1112 3336 1146
rect 3290 1074 3296 1112
rect 3330 1074 3336 1112
rect 3290 1044 3336 1074
rect 3290 1001 3296 1044
rect 3330 1001 3336 1044
rect 3290 976 3336 1001
rect 3290 928 3296 976
rect 3330 928 3336 976
rect 3290 908 3336 928
rect 3290 855 3296 908
rect 3330 855 3336 908
rect 3290 840 3336 855
rect 3290 782 3296 840
rect 3330 782 3336 840
rect 3290 772 3336 782
rect 3290 709 3296 772
rect 3330 709 3336 772
rect 3290 704 3336 709
rect 3290 602 3296 704
rect 3330 602 3336 704
rect 3290 597 3336 602
rect 3290 534 3296 597
rect 3330 534 3336 597
rect 3290 524 3336 534
rect 120 468 126 520
rect 160 468 166 520
rect 120 448 166 468
rect 120 400 126 448
rect 160 400 166 448
rect 120 376 166 400
rect 120 332 126 376
rect 160 332 166 376
rect 120 304 166 332
rect 120 270 126 304
rect 160 270 166 304
rect 120 252 166 270
rect 120 198 126 252
rect 160 198 166 252
rect 120 166 166 198
rect 3290 466 3296 524
rect 3330 466 3336 524
rect 3290 451 3336 466
rect 3290 398 3296 451
rect 3330 398 3336 451
rect 3290 378 3336 398
rect 3290 330 3296 378
rect 3330 330 3336 378
rect 3290 305 3336 330
rect 3290 262 3296 305
rect 3330 262 3336 305
rect 3290 232 3336 262
rect 3290 194 3296 232
rect 3330 194 3336 232
rect 3290 166 3336 194
rect 120 160 3336 166
rect 120 126 194 160
rect 232 126 262 160
rect 305 126 330 160
rect 378 126 398 160
rect 450 126 466 160
rect 522 126 534 160
rect 594 126 602 160
rect 666 126 670 160
rect 772 126 776 160
rect 840 126 848 160
rect 908 126 920 160
rect 976 126 992 160
rect 1044 126 1064 160
rect 1112 126 1136 160
rect 1180 126 1208 160
rect 1248 126 1280 160
rect 1316 126 1350 160
rect 1386 126 1418 160
rect 1458 126 1486 160
rect 1530 126 1554 160
rect 1602 126 1622 160
rect 1674 126 1690 160
rect 1746 126 1758 160
rect 1818 126 1826 160
rect 1890 126 1894 160
rect 1996 126 2000 160
rect 2064 126 2072 160
rect 2132 126 2144 160
rect 2200 126 2216 160
rect 2268 126 2288 160
rect 2336 126 2360 160
rect 2404 126 2432 160
rect 2472 126 2504 160
rect 2540 126 2574 160
rect 2610 126 2642 160
rect 2682 126 2710 160
rect 2754 126 2778 160
rect 2826 126 2846 160
rect 2898 126 2914 160
rect 2970 126 2982 160
rect 3042 126 3050 160
rect 3114 126 3118 160
rect 3220 126 3224 160
rect 3258 126 3336 160
rect 120 120 3336 126
<< viali >>
rect 206 39840 236 39874
rect 236 39840 240 39874
rect 286 39840 304 39874
rect 304 39840 320 39874
rect 366 39840 372 39874
rect 372 39840 400 39874
rect 447 39840 474 39874
rect 474 39840 481 39874
rect 528 39840 542 39874
rect 542 39840 562 39874
rect 609 39840 610 39874
rect 610 39840 643 39874
rect 690 39840 712 39874
rect 712 39840 724 39874
rect 800 39840 814 39874
rect 814 39840 834 39874
rect 873 39840 882 39874
rect 882 39840 907 39874
rect 946 39840 950 39874
rect 950 39840 980 39874
rect 1019 39840 1052 39874
rect 1052 39840 1053 39874
rect 1092 39840 1120 39874
rect 1120 39840 1126 39874
rect 1165 39840 1188 39874
rect 1188 39840 1199 39874
rect 1238 39840 1256 39874
rect 1256 39840 1272 39874
rect 1311 39840 1324 39874
rect 1324 39840 1345 39874
rect 1384 39840 1392 39874
rect 1392 39840 1418 39874
rect 1457 39840 1460 39874
rect 1460 39840 1491 39874
rect 1530 39840 1562 39874
rect 1562 39840 1564 39874
rect 1603 39840 1630 39874
rect 1630 39840 1637 39874
rect 1676 39840 1698 39874
rect 1698 39840 1710 39874
rect 1749 39840 1766 39874
rect 1766 39840 1783 39874
rect 1822 39840 1834 39874
rect 1834 39840 1856 39874
rect 1895 39840 1902 39874
rect 1902 39840 1929 39874
rect 1968 39840 1970 39874
rect 1970 39840 2002 39874
rect 2041 39840 2072 39874
rect 2072 39840 2075 39874
rect 2114 39840 2140 39874
rect 2140 39840 2148 39874
rect 2188 39840 2208 39874
rect 2208 39840 2222 39874
rect 2262 39840 2276 39874
rect 2276 39840 2296 39874
rect 2336 39840 2344 39874
rect 2344 39840 2370 39874
rect 2410 39840 2412 39874
rect 2412 39840 2444 39874
rect 2484 39840 2514 39874
rect 2514 39840 2518 39874
rect 2558 39840 2582 39874
rect 2582 39840 2592 39874
rect 2632 39840 2650 39874
rect 2650 39840 2666 39874
rect 2706 39840 2718 39874
rect 2718 39840 2740 39874
rect 2780 39840 2786 39874
rect 2786 39840 2814 39874
rect 2854 39840 2888 39874
rect 2928 39840 2956 39874
rect 2956 39840 2962 39874
rect 3002 39840 3024 39874
rect 3024 39840 3036 39874
rect 3076 39840 3092 39874
rect 3092 39840 3110 39874
rect 3150 39840 3160 39874
rect 3160 39840 3184 39874
rect 3224 39840 3228 39874
rect 3228 39840 3258 39874
rect 126 39772 160 39802
rect 126 39768 160 39772
rect 126 39704 160 39729
rect 126 39695 160 39704
rect 126 39636 160 39656
rect 126 39622 160 39636
rect 126 39568 160 39583
rect 126 39549 160 39568
rect 126 39500 160 39510
rect 126 39476 160 39500
rect 126 39432 160 39437
rect 126 39403 160 39432
rect 126 39330 160 39364
rect 126 39262 160 39291
rect 126 39257 160 39262
rect 126 39194 160 39218
rect 126 39184 160 39194
rect 3296 39770 3330 39802
rect 3296 39768 3330 39770
rect 3296 39702 3330 39730
rect 3296 39696 3330 39702
rect 3296 39634 3330 39658
rect 3296 39624 3330 39634
rect 3296 39566 3330 39586
rect 3296 39552 3330 39566
rect 3296 39498 3330 39514
rect 3296 39480 3330 39498
rect 3296 39430 3330 39442
rect 3296 39408 3330 39430
rect 3296 39362 3330 39370
rect 3296 39336 3330 39362
rect 3296 39294 3330 39298
rect 3296 39264 3330 39294
rect 126 39126 160 39145
rect 126 39111 160 39126
rect 126 39058 160 39072
rect 126 39038 160 39058
rect 126 38990 160 38999
rect 126 38965 160 38990
rect 126 38922 160 38926
rect 126 38892 160 38922
rect 126 38820 160 38853
rect 126 38819 160 38820
rect 126 38752 160 38780
rect 126 38746 160 38752
rect 126 38684 160 38707
rect 126 38673 160 38684
rect 126 38616 160 38634
rect 126 38600 160 38616
rect 126 38548 160 38561
rect 126 38527 160 38548
rect 126 38480 160 38488
rect 126 38454 160 38480
rect 126 38412 160 38415
rect 126 38381 160 38412
rect 126 38310 160 38342
rect 126 38308 160 38310
rect 126 38242 160 38269
rect 126 38235 160 38242
rect 126 38174 160 38196
rect 126 38162 160 38174
rect 126 38106 160 38123
rect 126 38089 160 38106
rect 126 38038 160 38050
rect 126 38016 160 38038
rect 126 37970 160 37977
rect 126 37943 160 37970
rect 126 37902 160 37904
rect 126 37870 160 37902
rect 126 37800 160 37831
rect 126 37797 160 37800
rect 126 37732 160 37758
rect 126 37724 160 37732
rect 126 37664 160 37685
rect 126 37651 160 37664
rect 126 37596 160 37612
rect 126 37578 160 37596
rect 126 37528 160 37539
rect 126 37505 160 37528
rect 126 37460 160 37466
rect 126 37432 160 37460
rect 126 37392 160 37393
rect 126 37359 160 37392
rect 126 37290 160 37320
rect 126 37286 160 37290
rect 126 37222 160 37247
rect 126 37213 160 37222
rect 126 37154 160 37174
rect 126 37140 160 37154
rect 126 37086 160 37101
rect 126 37067 160 37086
rect 126 37018 160 37028
rect 126 36994 160 37018
rect 126 36950 160 36955
rect 126 36921 160 36950
rect 126 36848 160 36882
rect 126 36780 160 36809
rect 126 36775 160 36780
rect 126 36712 160 36736
rect 126 36702 160 36712
rect 126 36644 160 36664
rect 126 36630 160 36644
rect 126 36576 160 36592
rect 126 36558 160 36576
rect 126 36508 160 36520
rect 126 36486 160 36508
rect 126 36440 160 36448
rect 126 36414 160 36440
rect 126 36372 160 36376
rect 126 36342 160 36372
rect 126 36270 160 36304
rect 126 36202 160 36232
rect 126 36198 160 36202
rect 126 36134 160 36160
rect 126 36126 160 36134
rect 126 36066 160 36088
rect 126 36054 160 36066
rect 126 35998 160 36016
rect 126 35982 160 35998
rect 126 35930 160 35944
rect 126 35910 160 35930
rect 126 35862 160 35872
rect 126 35838 160 35862
rect 126 35794 160 35800
rect 126 35766 160 35794
rect 126 35726 160 35728
rect 126 35694 160 35726
rect 126 35624 160 35656
rect 126 35622 160 35624
rect 126 35556 160 35584
rect 126 35550 160 35556
rect 126 35488 160 35512
rect 126 35478 160 35488
rect 126 35420 160 35440
rect 126 35406 160 35420
rect 126 35352 160 35368
rect 126 35334 160 35352
rect 126 35284 160 35296
rect 126 35262 160 35284
rect 126 35216 160 35224
rect 126 35190 160 35216
rect 126 35148 160 35152
rect 126 35118 160 35148
rect 126 35046 160 35080
rect 126 34978 160 35008
rect 126 34974 160 34978
rect 126 34910 160 34936
rect 126 34902 160 34910
rect 126 34842 160 34864
rect 126 34830 160 34842
rect 126 34774 160 34792
rect 126 34758 160 34774
rect 126 34706 160 34720
rect 126 34686 160 34706
rect 126 34638 160 34648
rect 126 34614 160 34638
rect 126 34570 160 34576
rect 126 34542 160 34570
rect 126 34502 160 34504
rect 126 34470 160 34502
rect 126 34400 160 34432
rect 126 34398 160 34400
rect 126 34332 160 34360
rect 126 34326 160 34332
rect 126 34264 160 34288
rect 126 34254 160 34264
rect 126 34196 160 34216
rect 126 34182 160 34196
rect 126 34128 160 34144
rect 126 34110 160 34128
rect 126 34060 160 34072
rect 126 34038 160 34060
rect 126 33992 160 34000
rect 126 33966 160 33992
rect 126 33924 160 33928
rect 126 33894 160 33924
rect 126 33822 160 33856
rect 126 33754 160 33784
rect 126 33750 160 33754
rect 126 33686 160 33712
rect 126 33678 160 33686
rect 126 33618 160 33640
rect 126 33606 160 33618
rect 126 33550 160 33568
rect 126 33534 160 33550
rect 126 33482 160 33496
rect 126 33462 160 33482
rect 126 33414 160 33424
rect 126 33390 160 33414
rect 126 33346 160 33352
rect 126 33318 160 33346
rect 126 33278 160 33280
rect 126 33246 160 33278
rect 126 33176 160 33208
rect 126 33174 160 33176
rect 126 33108 160 33136
rect 126 33102 160 33108
rect 126 33040 160 33064
rect 126 33030 160 33040
rect 126 32972 160 32992
rect 126 32958 160 32972
rect 126 32904 160 32920
rect 126 32886 160 32904
rect 126 32836 160 32848
rect 126 32814 160 32836
rect 126 32768 160 32776
rect 126 32742 160 32768
rect 126 32700 160 32704
rect 126 32670 160 32700
rect 126 32598 160 32632
rect 126 32530 160 32560
rect 126 32526 160 32530
rect 126 32462 160 32488
rect 126 32454 160 32462
rect 126 32394 160 32416
rect 126 32382 160 32394
rect 126 32326 160 32344
rect 126 32310 160 32326
rect 126 32258 160 32272
rect 126 32238 160 32258
rect 126 32190 160 32200
rect 126 32166 160 32190
rect 126 32122 160 32128
rect 126 32094 160 32122
rect 126 32054 160 32056
rect 126 32022 160 32054
rect 126 31952 160 31984
rect 126 31950 160 31952
rect 126 31884 160 31912
rect 126 31878 160 31884
rect 126 31816 160 31840
rect 126 31806 160 31816
rect 126 31748 160 31768
rect 126 31734 160 31748
rect 126 31680 160 31696
rect 126 31662 160 31680
rect 126 31612 160 31624
rect 126 31590 160 31612
rect 126 31544 160 31552
rect 126 31518 160 31544
rect 126 31476 160 31480
rect 126 31446 160 31476
rect 126 31374 160 31408
rect 126 31306 160 31336
rect 126 31302 160 31306
rect 126 31238 160 31264
rect 126 31230 160 31238
rect 126 31170 160 31192
rect 126 31158 160 31170
rect 126 31102 160 31120
rect 126 31086 160 31102
rect 126 31034 160 31048
rect 126 31014 160 31034
rect 126 30966 160 30976
rect 126 30942 160 30966
rect 126 30898 160 30904
rect 126 30870 160 30898
rect 126 30830 160 30832
rect 126 30798 160 30830
rect 126 30728 160 30760
rect 126 30726 160 30728
rect 126 30660 160 30688
rect 126 30654 160 30660
rect 126 30592 160 30616
rect 126 30582 160 30592
rect 126 30524 160 30544
rect 126 30510 160 30524
rect 126 30456 160 30472
rect 126 30438 160 30456
rect 126 30388 160 30400
rect 126 30366 160 30388
rect 126 30320 160 30328
rect 126 30294 160 30320
rect 126 30252 160 30256
rect 126 30222 160 30252
rect 126 30150 160 30184
rect 126 30082 160 30112
rect 126 30078 160 30082
rect 126 30014 160 30040
rect 126 30006 160 30014
rect 126 29946 160 29968
rect 126 29934 160 29946
rect 126 29878 160 29896
rect 126 29862 160 29878
rect 126 29810 160 29824
rect 126 29790 160 29810
rect 126 29742 160 29752
rect 126 29718 160 29742
rect 126 29674 160 29680
rect 126 29646 160 29674
rect 126 29606 160 29608
rect 126 29574 160 29606
rect 126 29504 160 29536
rect 126 29502 160 29504
rect 126 29436 160 29464
rect 126 29430 160 29436
rect 126 29368 160 29392
rect 126 29358 160 29368
rect 126 29300 160 29320
rect 126 29286 160 29300
rect 126 29232 160 29248
rect 126 29214 160 29232
rect 126 29164 160 29176
rect 126 29142 160 29164
rect 126 29096 160 29104
rect 126 29070 160 29096
rect 126 29028 160 29032
rect 126 28998 160 29028
rect 126 28926 160 28960
rect 126 28858 160 28888
rect 126 28854 160 28858
rect 126 28790 160 28816
rect 126 28782 160 28790
rect 126 28722 160 28744
rect 126 28710 160 28722
rect 126 28654 160 28672
rect 126 28638 160 28654
rect 126 28586 160 28600
rect 126 28566 160 28586
rect 126 28518 160 28528
rect 126 28494 160 28518
rect 126 28450 160 28456
rect 126 28422 160 28450
rect 126 28382 160 28384
rect 126 28350 160 28382
rect 126 28280 160 28312
rect 126 28278 160 28280
rect 126 28212 160 28240
rect 126 28206 160 28212
rect 126 28144 160 28168
rect 126 28134 160 28144
rect 126 28076 160 28096
rect 126 28062 160 28076
rect 126 28008 160 28024
rect 126 27990 160 28008
rect 126 27940 160 27952
rect 126 27918 160 27940
rect 126 27872 160 27880
rect 126 27846 160 27872
rect 126 27804 160 27808
rect 126 27774 160 27804
rect 126 27702 160 27736
rect 126 27634 160 27664
rect 126 27630 160 27634
rect 126 27566 160 27592
rect 126 27558 160 27566
rect 126 27498 160 27520
rect 126 27486 160 27498
rect 126 27430 160 27448
rect 126 27414 160 27430
rect 126 27362 160 27376
rect 126 27342 160 27362
rect 126 27294 160 27304
rect 126 27270 160 27294
rect 126 27226 160 27232
rect 126 27198 160 27226
rect 126 27158 160 27160
rect 126 27126 160 27158
rect 126 27056 160 27088
rect 126 27054 160 27056
rect 126 26988 160 27016
rect 126 26982 160 26988
rect 126 26920 160 26944
rect 126 26910 160 26920
rect 126 26852 160 26872
rect 126 26838 160 26852
rect 126 26784 160 26800
rect 126 26766 160 26784
rect 126 26716 160 26728
rect 126 26694 160 26716
rect 126 26648 160 26656
rect 126 26622 160 26648
rect 126 26580 160 26584
rect 126 26550 160 26580
rect 126 26478 160 26512
rect 126 26410 160 26440
rect 126 26406 160 26410
rect 126 26342 160 26368
rect 126 26334 160 26342
rect 126 26274 160 26296
rect 126 26262 160 26274
rect 126 26206 160 26224
rect 126 26190 160 26206
rect 126 26138 160 26152
rect 126 26118 160 26138
rect 126 26070 160 26080
rect 126 26046 160 26070
rect 126 26002 160 26008
rect 126 25974 160 26002
rect 126 25934 160 25936
rect 126 25902 160 25934
rect 126 25832 160 25864
rect 126 25830 160 25832
rect 126 25764 160 25792
rect 126 25758 160 25764
rect 126 25696 160 25720
rect 126 25686 160 25696
rect 126 25628 160 25648
rect 126 25614 160 25628
rect 126 25560 160 25576
rect 126 25542 160 25560
rect 126 25492 160 25504
rect 126 25470 160 25492
rect 126 25424 160 25432
rect 126 25398 160 25424
rect 126 25356 160 25360
rect 126 25326 160 25356
rect 126 25254 160 25288
rect 126 25186 160 25216
rect 126 25182 160 25186
rect 126 25118 160 25144
rect 126 25110 160 25118
rect 126 25050 160 25072
rect 126 25038 160 25050
rect 126 24982 160 25000
rect 126 24966 160 24982
rect 126 24914 160 24928
rect 126 24894 160 24914
rect 126 24846 160 24856
rect 126 24822 160 24846
rect 126 24778 160 24784
rect 126 24750 160 24778
rect 126 24710 160 24712
rect 126 24678 160 24710
rect 126 24608 160 24640
rect 126 24606 160 24608
rect 126 24540 160 24568
rect 126 24534 160 24540
rect 126 24472 160 24496
rect 126 24462 160 24472
rect 126 24404 160 24424
rect 126 24390 160 24404
rect 126 24336 160 24352
rect 126 24318 160 24336
rect 126 24268 160 24280
rect 126 24246 160 24268
rect 126 24200 160 24208
rect 126 24174 160 24200
rect 126 24132 160 24136
rect 126 24102 160 24132
rect 126 24030 160 24064
rect 126 23962 160 23992
rect 126 23958 160 23962
rect 126 23894 160 23920
rect 126 23886 160 23894
rect 126 23826 160 23848
rect 126 23814 160 23826
rect 126 23758 160 23776
rect 126 23742 160 23758
rect 126 23690 160 23704
rect 126 23670 160 23690
rect 126 23622 160 23632
rect 126 23598 160 23622
rect 126 23554 160 23560
rect 126 23526 160 23554
rect 126 23486 160 23488
rect 126 23454 160 23486
rect 126 23384 160 23416
rect 126 23382 160 23384
rect 126 23316 160 23344
rect 126 23310 160 23316
rect 126 23248 160 23272
rect 126 23238 160 23248
rect 126 23180 160 23200
rect 126 23166 160 23180
rect 126 23112 160 23128
rect 126 23094 160 23112
rect 126 23044 160 23056
rect 126 23022 160 23044
rect 126 22976 160 22984
rect 126 22950 160 22976
rect 126 22908 160 22912
rect 126 22878 160 22908
rect 126 22806 160 22840
rect 126 22738 160 22768
rect 126 22734 160 22738
rect 126 22670 160 22696
rect 126 22662 160 22670
rect 126 22602 160 22624
rect 126 22590 160 22602
rect 126 22534 160 22552
rect 126 22518 160 22534
rect 126 22466 160 22480
rect 126 22446 160 22466
rect 126 22398 160 22408
rect 126 22374 160 22398
rect 126 22330 160 22336
rect 126 22302 160 22330
rect 126 22262 160 22264
rect 126 22230 160 22262
rect 126 22160 160 22192
rect 126 22158 160 22160
rect 126 22092 160 22120
rect 126 22086 160 22092
rect 126 22024 160 22048
rect 126 22014 160 22024
rect 126 21956 160 21976
rect 126 21942 160 21956
rect 126 21888 160 21904
rect 126 21870 160 21888
rect 126 21820 160 21832
rect 126 21798 160 21820
rect 126 21752 160 21760
rect 126 21726 160 21752
rect 126 21684 160 21688
rect 126 21654 160 21684
rect 126 21582 160 21616
rect 126 21514 160 21544
rect 126 21510 160 21514
rect 126 21446 160 21472
rect 126 21438 160 21446
rect 126 21378 160 21400
rect 126 21366 160 21378
rect 126 21310 160 21328
rect 126 21294 160 21310
rect 126 21242 160 21256
rect 126 21222 160 21242
rect 126 21174 160 21184
rect 126 21150 160 21174
rect 126 21106 160 21112
rect 126 21078 160 21106
rect 126 21038 160 21040
rect 126 21006 160 21038
rect 126 20936 160 20968
rect 126 20934 160 20936
rect 126 20868 160 20896
rect 126 20862 160 20868
rect 126 20800 160 20824
rect 126 20790 160 20800
rect 126 20732 160 20752
rect 126 20718 160 20732
rect 126 20664 160 20680
rect 126 20646 160 20664
rect 126 20596 160 20608
rect 126 20574 160 20596
rect 126 20528 160 20536
rect 126 20502 160 20528
rect 126 20460 160 20464
rect 126 20430 160 20460
rect 126 20358 160 20392
rect 126 20290 160 20320
rect 126 20286 160 20290
rect 126 20222 160 20248
rect 126 20214 160 20222
rect 126 20154 160 20176
rect 126 20142 160 20154
rect 126 20086 160 20104
rect 126 20070 160 20086
rect 126 20018 160 20032
rect 126 19998 160 20018
rect 126 19950 160 19960
rect 126 19926 160 19950
rect 126 19882 160 19888
rect 126 19854 160 19882
rect 126 19814 160 19816
rect 126 19782 160 19814
rect 126 19712 160 19744
rect 126 19710 160 19712
rect 126 19644 160 19672
rect 126 19638 160 19644
rect 126 19576 160 19600
rect 126 19566 160 19576
rect 126 19508 160 19528
rect 126 19494 160 19508
rect 126 19440 160 19456
rect 126 19422 160 19440
rect 126 19372 160 19384
rect 126 19350 160 19372
rect 126 19304 160 19312
rect 126 19278 160 19304
rect 126 19236 160 19240
rect 126 19206 160 19236
rect 126 19134 160 19168
rect 126 19066 160 19096
rect 126 19062 160 19066
rect 126 18998 160 19024
rect 126 18990 160 18998
rect 126 18930 160 18952
rect 126 18918 160 18930
rect 126 18862 160 18880
rect 126 18846 160 18862
rect 126 18794 160 18808
rect 126 18774 160 18794
rect 126 18726 160 18736
rect 126 18702 160 18726
rect 126 18658 160 18664
rect 126 18630 160 18658
rect 126 18590 160 18592
rect 126 18558 160 18590
rect 126 18488 160 18520
rect 126 18486 160 18488
rect 126 18420 160 18448
rect 126 18414 160 18420
rect 126 18352 160 18376
rect 126 18342 160 18352
rect 126 18284 160 18304
rect 126 18270 160 18284
rect 126 18216 160 18232
rect 126 18198 160 18216
rect 126 18148 160 18160
rect 126 18126 160 18148
rect 126 18080 160 18088
rect 126 18054 160 18080
rect 126 18012 160 18016
rect 126 17982 160 18012
rect 126 17910 160 17944
rect 126 17842 160 17872
rect 126 17838 160 17842
rect 126 17774 160 17800
rect 126 17766 160 17774
rect 126 17706 160 17728
rect 126 17694 160 17706
rect 126 17638 160 17656
rect 126 17622 160 17638
rect 126 17570 160 17584
rect 126 17550 160 17570
rect 126 17502 160 17512
rect 126 17478 160 17502
rect 126 17434 160 17440
rect 126 17406 160 17434
rect 126 17366 160 17368
rect 126 17334 160 17366
rect 126 17264 160 17296
rect 126 17262 160 17264
rect 126 17196 160 17224
rect 126 17190 160 17196
rect 126 17128 160 17152
rect 126 17118 160 17128
rect 126 17060 160 17080
rect 126 17046 160 17060
rect 126 16992 160 17008
rect 126 16974 160 16992
rect 126 16924 160 16936
rect 126 16902 160 16924
rect 126 16856 160 16864
rect 126 16830 160 16856
rect 126 16788 160 16792
rect 126 16758 160 16788
rect 126 16686 160 16720
rect 126 16618 160 16648
rect 126 16614 160 16618
rect 126 16550 160 16576
rect 126 16542 160 16550
rect 126 16482 160 16504
rect 126 16470 160 16482
rect 126 16414 160 16432
rect 126 16398 160 16414
rect 126 16346 160 16360
rect 126 16326 160 16346
rect 126 16278 160 16288
rect 126 16254 160 16278
rect 126 16210 160 16216
rect 126 16182 160 16210
rect 126 16142 160 16144
rect 126 16110 160 16142
rect 126 16040 160 16072
rect 126 16038 160 16040
rect 126 15972 160 16000
rect 126 15966 160 15972
rect 126 15904 160 15928
rect 126 15894 160 15904
rect 126 15836 160 15856
rect 126 15822 160 15836
rect 126 15768 160 15784
rect 126 15750 160 15768
rect 126 15700 160 15712
rect 126 15678 160 15700
rect 126 15632 160 15640
rect 126 15606 160 15632
rect 126 15564 160 15568
rect 126 15534 160 15564
rect 126 15462 160 15496
rect 126 15394 160 15424
rect 126 15390 160 15394
rect 126 15326 160 15352
rect 126 15318 160 15326
rect 126 15258 160 15280
rect 126 15246 160 15258
rect 126 15190 160 15208
rect 126 15174 160 15190
rect 126 15122 160 15136
rect 126 15102 160 15122
rect 126 15054 160 15064
rect 126 15030 160 15054
rect 126 14986 160 14992
rect 126 14958 160 14986
rect 126 14918 160 14920
rect 126 14886 160 14918
rect 126 14816 160 14848
rect 126 14814 160 14816
rect 126 14748 160 14776
rect 126 14742 160 14748
rect 126 14680 160 14704
rect 126 14670 160 14680
rect 126 14612 160 14632
rect 126 14598 160 14612
rect 126 14544 160 14560
rect 126 14526 160 14544
rect 126 14476 160 14488
rect 126 14454 160 14476
rect 126 14408 160 14416
rect 126 14382 160 14408
rect 126 14340 160 14344
rect 126 14310 160 14340
rect 126 14238 160 14272
rect 126 14170 160 14200
rect 126 14166 160 14170
rect 126 14102 160 14128
rect 126 14094 160 14102
rect 126 14034 160 14056
rect 126 14022 160 14034
rect 126 13966 160 13984
rect 126 13950 160 13966
rect 126 13898 160 13912
rect 126 13878 160 13898
rect 126 13830 160 13840
rect 126 13806 160 13830
rect 126 13762 160 13768
rect 126 13734 160 13762
rect 126 13694 160 13696
rect 126 13662 160 13694
rect 126 13592 160 13624
rect 126 13590 160 13592
rect 126 13524 160 13552
rect 126 13518 160 13524
rect 126 13456 160 13480
rect 126 13446 160 13456
rect 126 13388 160 13408
rect 126 13374 160 13388
rect 126 13320 160 13336
rect 126 13302 160 13320
rect 126 13252 160 13264
rect 126 13230 160 13252
rect 126 13184 160 13192
rect 126 13158 160 13184
rect 126 13116 160 13120
rect 126 13086 160 13116
rect 126 13014 160 13048
rect 126 12946 160 12976
rect 126 12942 160 12946
rect 126 12878 160 12904
rect 126 12870 160 12878
rect 126 12810 160 12832
rect 126 12798 160 12810
rect 126 12742 160 12760
rect 126 12726 160 12742
rect 126 12674 160 12688
rect 126 12654 160 12674
rect 126 12606 160 12616
rect 126 12582 160 12606
rect 126 12538 160 12544
rect 126 12510 160 12538
rect 126 12470 160 12472
rect 126 12438 160 12470
rect 126 12368 160 12400
rect 126 12366 160 12368
rect 126 12300 160 12328
rect 126 12294 160 12300
rect 126 12232 160 12256
rect 126 12222 160 12232
rect 126 12164 160 12184
rect 126 12150 160 12164
rect 126 12096 160 12112
rect 126 12078 160 12096
rect 126 12028 160 12040
rect 126 12006 160 12028
rect 126 11960 160 11968
rect 126 11934 160 11960
rect 126 11892 160 11896
rect 126 11862 160 11892
rect 126 11790 160 11824
rect 126 11722 160 11752
rect 126 11718 160 11722
rect 126 11654 160 11680
rect 126 11646 160 11654
rect 126 11586 160 11608
rect 126 11574 160 11586
rect 126 11518 160 11536
rect 126 11502 160 11518
rect 126 11450 160 11464
rect 126 11430 160 11450
rect 126 11382 160 11392
rect 126 11358 160 11382
rect 126 11314 160 11320
rect 126 11286 160 11314
rect 126 11246 160 11248
rect 126 11214 160 11246
rect 126 11144 160 11176
rect 126 11142 160 11144
rect 126 11076 160 11104
rect 126 11070 160 11076
rect 126 11008 160 11032
rect 126 10998 160 11008
rect 126 10940 160 10960
rect 126 10926 160 10940
rect 126 10872 160 10888
rect 126 10854 160 10872
rect 126 10804 160 10816
rect 126 10782 160 10804
rect 126 10736 160 10744
rect 126 10710 160 10736
rect 126 10668 160 10672
rect 126 10638 160 10668
rect 126 10566 160 10600
rect 126 10498 160 10528
rect 126 10494 160 10498
rect 126 10430 160 10456
rect 126 10422 160 10430
rect 126 10362 160 10384
rect 126 10350 160 10362
rect 126 10294 160 10312
rect 126 10278 160 10294
rect 126 10226 160 10240
rect 126 10206 160 10226
rect 126 10158 160 10168
rect 126 10134 160 10158
rect 126 10090 160 10096
rect 126 10062 160 10090
rect 126 10022 160 10024
rect 126 9990 160 10022
rect 126 9920 160 9952
rect 126 9918 160 9920
rect 126 9852 160 9880
rect 126 9846 160 9852
rect 126 9784 160 9808
rect 126 9774 160 9784
rect 126 9716 160 9736
rect 126 9702 160 9716
rect 126 9648 160 9664
rect 126 9630 160 9648
rect 126 9580 160 9592
rect 126 9558 160 9580
rect 126 9512 160 9520
rect 126 9486 160 9512
rect 126 9444 160 9448
rect 126 9414 160 9444
rect 126 9342 160 9376
rect 126 9274 160 9304
rect 126 9270 160 9274
rect 126 9206 160 9232
rect 126 9198 160 9206
rect 126 9138 160 9160
rect 126 9126 160 9138
rect 126 9070 160 9088
rect 126 9054 160 9070
rect 126 9002 160 9016
rect 126 8982 160 9002
rect 126 8934 160 8944
rect 126 8910 160 8934
rect 126 8866 160 8872
rect 126 8838 160 8866
rect 126 8798 160 8800
rect 126 8766 160 8798
rect 126 8696 160 8728
rect 126 8694 160 8696
rect 126 8628 160 8656
rect 126 8622 160 8628
rect 126 8560 160 8584
rect 126 8550 160 8560
rect 126 8492 160 8512
rect 126 8478 160 8492
rect 126 8424 160 8440
rect 126 8406 160 8424
rect 126 8356 160 8368
rect 126 8334 160 8356
rect 126 8288 160 8296
rect 126 8262 160 8288
rect 126 8220 160 8224
rect 126 8190 160 8220
rect 126 8118 160 8152
rect 126 8050 160 8080
rect 126 8046 160 8050
rect 126 7982 160 8008
rect 126 7974 160 7982
rect 126 7914 160 7936
rect 126 7902 160 7914
rect 126 7846 160 7864
rect 126 7830 160 7846
rect 126 7778 160 7792
rect 126 7758 160 7778
rect 126 7710 160 7720
rect 126 7686 160 7710
rect 126 7642 160 7648
rect 126 7614 160 7642
rect 126 7574 160 7576
rect 126 7542 160 7574
rect 126 7472 160 7504
rect 126 7470 160 7472
rect 126 7404 160 7432
rect 126 7398 160 7404
rect 126 7336 160 7360
rect 126 7326 160 7336
rect 126 7268 160 7288
rect 126 7254 160 7268
rect 126 7200 160 7216
rect 126 7182 160 7200
rect 126 7132 160 7144
rect 126 7110 160 7132
rect 126 7064 160 7072
rect 126 7038 160 7064
rect 126 6996 160 7000
rect 126 6966 160 6996
rect 126 6894 160 6928
rect 126 6826 160 6856
rect 126 6822 160 6826
rect 126 6758 160 6784
rect 126 6750 160 6758
rect 126 6690 160 6712
rect 126 6678 160 6690
rect 126 6622 160 6640
rect 126 6606 160 6622
rect 126 6554 160 6568
rect 126 6534 160 6554
rect 126 6486 160 6496
rect 126 6462 160 6486
rect 126 6418 160 6424
rect 126 6390 160 6418
rect 126 6350 160 6352
rect 126 6318 160 6350
rect 126 6248 160 6280
rect 126 6246 160 6248
rect 126 6180 160 6208
rect 126 6174 160 6180
rect 126 6112 160 6136
rect 126 6102 160 6112
rect 126 6044 160 6064
rect 126 6030 160 6044
rect 126 5976 160 5992
rect 126 5958 160 5976
rect 126 5908 160 5920
rect 126 5886 160 5908
rect 126 5840 160 5848
rect 126 5814 160 5840
rect 126 5772 160 5776
rect 126 5742 160 5772
rect 126 5670 160 5704
rect 126 5602 160 5632
rect 126 5598 160 5602
rect 126 5534 160 5560
rect 126 5526 160 5534
rect 126 5466 160 5488
rect 126 5454 160 5466
rect 126 5398 160 5416
rect 126 5382 160 5398
rect 126 5330 160 5344
rect 126 5310 160 5330
rect 126 5262 160 5272
rect 126 5238 160 5262
rect 126 5194 160 5200
rect 126 5166 160 5194
rect 126 5126 160 5128
rect 126 5094 160 5126
rect 126 5024 160 5056
rect 126 5022 160 5024
rect 126 4956 160 4984
rect 126 4950 160 4956
rect 126 4888 160 4912
rect 126 4878 160 4888
rect 126 4820 160 4840
rect 126 4806 160 4820
rect 126 4752 160 4768
rect 126 4734 160 4752
rect 126 4684 160 4696
rect 126 4662 160 4684
rect 126 4616 160 4624
rect 126 4590 160 4616
rect 126 4548 160 4552
rect 126 4518 160 4548
rect 126 4446 160 4480
rect 126 4378 160 4408
rect 126 4374 160 4378
rect 126 4310 160 4336
rect 126 4302 160 4310
rect 126 4242 160 4264
rect 126 4230 160 4242
rect 126 4174 160 4192
rect 126 4158 160 4174
rect 126 4106 160 4120
rect 126 4086 160 4106
rect 126 4038 160 4048
rect 126 4014 160 4038
rect 126 3970 160 3976
rect 126 3942 160 3970
rect 126 3902 160 3904
rect 126 3870 160 3902
rect 126 3800 160 3832
rect 126 3798 160 3800
rect 126 3732 160 3760
rect 126 3726 160 3732
rect 126 3664 160 3688
rect 126 3654 160 3664
rect 126 3596 160 3616
rect 126 3582 160 3596
rect 126 3528 160 3544
rect 126 3510 160 3528
rect 126 3460 160 3472
rect 126 3438 160 3460
rect 126 3392 160 3400
rect 126 3366 160 3392
rect 126 3324 160 3328
rect 126 3294 160 3324
rect 126 3222 160 3256
rect 126 3154 160 3184
rect 126 3150 160 3154
rect 126 3086 160 3112
rect 126 3078 160 3086
rect 126 3018 160 3040
rect 126 3006 160 3018
rect 126 2950 160 2968
rect 126 2934 160 2950
rect 126 2882 160 2896
rect 126 2862 160 2882
rect 126 2814 160 2824
rect 126 2790 160 2814
rect 126 2746 160 2752
rect 126 2718 160 2746
rect 126 2678 160 2680
rect 126 2646 160 2678
rect 126 2576 160 2608
rect 126 2574 160 2576
rect 126 2508 160 2536
rect 126 2502 160 2508
rect 126 2440 160 2464
rect 126 2430 160 2440
rect 126 2372 160 2392
rect 126 2358 160 2372
rect 126 2304 160 2320
rect 126 2286 160 2304
rect 126 2236 160 2248
rect 126 2214 160 2236
rect 126 2168 160 2176
rect 126 2142 160 2168
rect 126 2100 160 2104
rect 126 2070 160 2100
rect 126 1998 160 2032
rect 126 1930 160 1960
rect 126 1926 160 1930
rect 126 1862 160 1888
rect 126 1854 160 1862
rect 126 1794 160 1816
rect 126 1782 160 1794
rect 126 1726 160 1744
rect 126 1710 160 1726
rect 126 1658 160 1672
rect 126 1638 160 1658
rect 126 1590 160 1600
rect 126 1566 160 1590
rect 126 1522 160 1528
rect 126 1494 160 1522
rect 126 1454 160 1456
rect 126 1422 160 1454
rect 126 1352 160 1384
rect 126 1350 160 1352
rect 126 1284 160 1312
rect 126 1278 160 1284
rect 126 1216 160 1240
rect 126 1206 160 1216
rect 126 1148 160 1168
rect 126 1134 160 1148
rect 126 1080 160 1096
rect 126 1062 160 1080
rect 126 1012 160 1024
rect 126 990 160 1012
rect 126 944 160 952
rect 126 918 160 944
rect 126 876 160 880
rect 126 846 160 876
rect 126 774 160 808
rect 126 706 160 736
rect 126 702 160 706
rect 126 638 160 664
rect 126 630 160 638
rect 126 570 160 592
rect 126 558 160 570
rect 462 39144 465 39178
rect 465 39144 496 39178
rect 538 39144 567 39178
rect 567 39144 572 39178
rect 648 39144 669 39178
rect 669 39144 682 39178
rect 720 39144 737 39178
rect 737 39144 754 39178
rect 792 39144 805 39178
rect 805 39144 826 39178
rect 864 39144 873 39178
rect 873 39144 898 39178
rect 936 39144 941 39178
rect 941 39144 970 39178
rect 1008 39144 1009 39178
rect 1009 39144 1042 39178
rect 1080 39144 1111 39178
rect 1111 39144 1114 39178
rect 1152 39144 1179 39178
rect 1179 39144 1186 39178
rect 1224 39144 1247 39178
rect 1247 39144 1258 39178
rect 1296 39144 1315 39178
rect 1315 39144 1330 39178
rect 1368 39144 1383 39178
rect 1383 39144 1402 39178
rect 1440 39144 1451 39178
rect 1451 39144 1474 39178
rect 1512 39144 1519 39178
rect 1519 39144 1546 39178
rect 1584 39144 1587 39178
rect 1587 39144 1618 39178
rect 1656 39144 1689 39178
rect 1689 39144 1690 39178
rect 1728 39144 1757 39178
rect 1757 39144 1762 39178
rect 1800 39144 1825 39178
rect 1825 39144 1834 39178
rect 1872 39144 1893 39178
rect 1893 39144 1906 39178
rect 1944 39144 1961 39178
rect 1961 39144 1978 39178
rect 2016 39144 2029 39178
rect 2029 39144 2050 39178
rect 2088 39144 2097 39178
rect 2097 39144 2122 39178
rect 2161 39144 2165 39178
rect 2165 39144 2195 39178
rect 2234 39144 2267 39178
rect 2267 39144 2268 39178
rect 2307 39144 2335 39178
rect 2335 39144 2341 39178
rect 2380 39144 2403 39178
rect 2403 39144 2414 39178
rect 2453 39144 2471 39178
rect 2471 39144 2487 39178
rect 2526 39144 2539 39178
rect 2539 39144 2560 39178
rect 2599 39144 2607 39178
rect 2607 39144 2633 39178
rect 2672 39144 2675 39178
rect 2675 39144 2706 39178
rect 2745 39144 2777 39178
rect 2777 39144 2779 39178
rect 2818 39144 2845 39178
rect 2845 39144 2852 39178
rect 2891 39144 2913 39178
rect 2913 39144 2925 39178
rect 2964 39144 2981 39178
rect 2981 39144 2998 39178
rect 386 39089 420 39106
rect 386 39072 420 39089
rect 386 39021 420 39033
rect 386 38999 420 39021
rect 3036 39076 3070 39106
rect 3036 39072 3070 39076
rect 386 38953 420 38960
rect 386 38926 420 38953
rect 3036 39008 3070 39034
rect 3036 39000 3070 39008
rect 386 38885 420 38887
rect 386 38853 420 38885
rect 386 38783 420 38814
rect 386 38780 420 38783
rect 386 38715 420 38741
rect 386 38707 420 38715
rect 386 38647 420 38668
rect 386 38634 420 38647
rect 386 38579 420 38595
rect 386 38561 420 38579
rect 386 38511 420 38522
rect 386 38488 420 38511
rect 386 38443 420 38449
rect 386 38415 420 38443
rect 386 38375 420 38376
rect 386 38342 420 38375
rect 386 38273 420 38303
rect 386 38269 420 38273
rect 386 38205 420 38230
rect 386 38196 420 38205
rect 386 38137 420 38157
rect 386 38123 420 38137
rect 386 38069 420 38084
rect 386 38050 420 38069
rect 386 38001 420 38011
rect 386 37977 420 38001
rect 386 37933 420 37938
rect 386 37904 420 37933
rect 386 37831 420 37865
rect 386 37763 420 37792
rect 386 37758 420 37763
rect 386 37695 420 37719
rect 386 37685 420 37695
rect 386 37627 420 37647
rect 386 37613 420 37627
rect 386 37559 420 37575
rect 386 37541 420 37559
rect 386 37491 420 37503
rect 386 37469 420 37491
rect 386 37423 420 37431
rect 386 37397 420 37423
rect 386 37355 420 37359
rect 386 37325 420 37355
rect 386 37253 420 37287
rect 386 37185 420 37215
rect 386 37181 420 37185
rect 386 37117 420 37143
rect 386 37109 420 37117
rect 386 37049 420 37071
rect 386 37037 420 37049
rect 531 38930 565 38964
rect 531 38857 565 38891
rect 531 38784 565 38818
rect 531 38711 565 38745
rect 531 38638 565 38672
rect 531 38565 565 38599
rect 531 38492 565 38526
rect 531 38419 565 38453
rect 531 38346 565 38380
rect 531 38273 565 38307
rect 531 38200 565 38234
rect 531 38127 565 38161
rect 531 38054 565 38088
rect 531 37980 565 38014
rect 531 37906 565 37940
rect 531 37832 565 37866
rect 531 37758 565 37792
rect 531 37684 565 37718
rect 531 37610 565 37644
rect 531 37536 565 37570
rect 531 37462 565 37496
rect 531 37388 565 37422
rect 531 37314 565 37348
rect 531 37240 565 37274
rect 531 37166 565 37200
rect 531 37092 565 37126
rect 531 37018 565 37052
rect 767 38930 801 38964
rect 767 38857 801 38891
rect 767 38784 801 38818
rect 767 38711 801 38745
rect 767 38638 801 38672
rect 767 38565 801 38599
rect 767 38492 801 38526
rect 767 38419 801 38453
rect 767 38346 801 38380
rect 767 38273 801 38307
rect 767 38200 801 38234
rect 767 38127 801 38161
rect 767 38054 801 38088
rect 767 37980 801 38014
rect 767 37906 801 37940
rect 767 37832 801 37866
rect 767 37758 801 37792
rect 767 37684 801 37718
rect 767 37610 801 37644
rect 767 37536 801 37570
rect 767 37462 801 37496
rect 767 37388 801 37422
rect 767 37314 801 37348
rect 767 37240 801 37274
rect 767 37166 801 37200
rect 767 37092 801 37126
rect 767 37018 801 37052
rect 1003 38930 1037 38964
rect 1003 38857 1037 38891
rect 1003 38784 1037 38818
rect 1003 38711 1037 38745
rect 1003 38638 1037 38672
rect 1003 38565 1037 38599
rect 1003 38492 1037 38526
rect 1003 38419 1037 38453
rect 1003 38346 1037 38380
rect 1003 38273 1037 38307
rect 1003 38200 1037 38234
rect 1003 38127 1037 38161
rect 1003 38054 1037 38088
rect 1003 37980 1037 38014
rect 1003 37906 1037 37940
rect 1003 37832 1037 37866
rect 1003 37758 1037 37792
rect 1003 37684 1037 37718
rect 1003 37610 1037 37644
rect 1003 37536 1037 37570
rect 1003 37462 1037 37496
rect 1003 37388 1037 37422
rect 1003 37314 1037 37348
rect 1003 37240 1037 37274
rect 1003 37166 1037 37200
rect 1003 37092 1037 37126
rect 1003 37018 1037 37052
rect 1239 38930 1273 38964
rect 1239 38857 1273 38891
rect 1239 38784 1273 38818
rect 1239 38711 1273 38745
rect 1239 38638 1273 38672
rect 1239 38565 1273 38599
rect 1239 38492 1273 38526
rect 1239 38419 1273 38453
rect 1239 38346 1273 38380
rect 1239 38273 1273 38307
rect 1239 38200 1273 38234
rect 1239 38127 1273 38161
rect 1239 38054 1273 38088
rect 1239 37980 1273 38014
rect 1239 37906 1273 37940
rect 1239 37832 1273 37866
rect 1239 37758 1273 37792
rect 1239 37684 1273 37718
rect 1239 37610 1273 37644
rect 1239 37536 1273 37570
rect 1239 37462 1273 37496
rect 1239 37388 1273 37422
rect 1239 37314 1273 37348
rect 1239 37240 1273 37274
rect 1239 37166 1273 37200
rect 1239 37092 1273 37126
rect 1239 37018 1273 37052
rect 1475 38930 1509 38964
rect 1475 38857 1509 38891
rect 1475 38784 1509 38818
rect 1475 38711 1509 38745
rect 1475 38638 1509 38672
rect 1475 38565 1509 38599
rect 1475 38492 1509 38526
rect 1475 38419 1509 38453
rect 1475 38346 1509 38380
rect 1475 38273 1509 38307
rect 1475 38200 1509 38234
rect 1475 38127 1509 38161
rect 1475 38054 1509 38088
rect 1475 37980 1509 38014
rect 1475 37906 1509 37940
rect 1475 37832 1509 37866
rect 1475 37758 1509 37792
rect 1475 37684 1509 37718
rect 1475 37610 1509 37644
rect 1475 37536 1509 37570
rect 1475 37462 1509 37496
rect 1475 37388 1509 37422
rect 1475 37314 1509 37348
rect 1475 37240 1509 37274
rect 1475 37166 1509 37200
rect 1475 37092 1509 37126
rect 1475 37018 1509 37052
rect 1711 38930 1745 38964
rect 1711 38857 1745 38891
rect 1711 38784 1745 38818
rect 1711 38711 1745 38745
rect 1711 38638 1745 38672
rect 1711 38565 1745 38599
rect 1711 38492 1745 38526
rect 1711 38419 1745 38453
rect 1711 38346 1745 38380
rect 1711 38273 1745 38307
rect 1711 38200 1745 38234
rect 1711 38127 1745 38161
rect 1711 38054 1745 38088
rect 1711 37980 1745 38014
rect 1711 37906 1745 37940
rect 1711 37832 1745 37866
rect 1711 37758 1745 37792
rect 1711 37684 1745 37718
rect 1711 37610 1745 37644
rect 1711 37536 1745 37570
rect 1711 37462 1745 37496
rect 1711 37388 1745 37422
rect 1711 37314 1745 37348
rect 1711 37240 1745 37274
rect 1711 37166 1745 37200
rect 1711 37092 1745 37126
rect 1711 37018 1745 37052
rect 1947 38930 1981 38964
rect 1947 38857 1981 38891
rect 1947 38784 1981 38818
rect 1947 38711 1981 38745
rect 1947 38638 1981 38672
rect 1947 38565 1981 38599
rect 1947 38492 1981 38526
rect 1947 38419 1981 38453
rect 1947 38346 1981 38380
rect 1947 38273 1981 38307
rect 1947 38200 1981 38234
rect 1947 38127 1981 38161
rect 1947 38054 1981 38088
rect 1947 37980 1981 38014
rect 1947 37906 1981 37940
rect 1947 37832 1981 37866
rect 1947 37758 1981 37792
rect 1947 37684 1981 37718
rect 1947 37610 1981 37644
rect 1947 37536 1981 37570
rect 1947 37462 1981 37496
rect 1947 37388 1981 37422
rect 1947 37314 1981 37348
rect 1947 37240 1981 37274
rect 1947 37166 1981 37200
rect 1947 37092 1981 37126
rect 1947 37018 1981 37052
rect 2183 38930 2217 38964
rect 2183 38857 2217 38891
rect 2183 38784 2217 38818
rect 2183 38711 2217 38745
rect 2183 38638 2217 38672
rect 2183 38565 2217 38599
rect 2183 38492 2217 38526
rect 2183 38419 2217 38453
rect 2183 38346 2217 38380
rect 2183 38273 2217 38307
rect 2183 38200 2217 38234
rect 2183 38127 2217 38161
rect 2183 38054 2217 38088
rect 2183 37980 2217 38014
rect 2183 37906 2217 37940
rect 2183 37832 2217 37866
rect 2183 37758 2217 37792
rect 2183 37684 2217 37718
rect 2183 37610 2217 37644
rect 2183 37536 2217 37570
rect 2183 37462 2217 37496
rect 2183 37388 2217 37422
rect 2183 37314 2217 37348
rect 2183 37240 2217 37274
rect 2183 37166 2217 37200
rect 2183 37092 2217 37126
rect 2183 37018 2217 37052
rect 2419 38930 2453 38964
rect 2419 38857 2453 38891
rect 2419 38784 2453 38818
rect 2419 38711 2453 38745
rect 2419 38638 2453 38672
rect 2419 38565 2453 38599
rect 2419 38492 2453 38526
rect 2419 38419 2453 38453
rect 2419 38346 2453 38380
rect 2419 38273 2453 38307
rect 2419 38200 2453 38234
rect 2419 38127 2453 38161
rect 2419 38054 2453 38088
rect 2419 37980 2453 38014
rect 2419 37906 2453 37940
rect 2419 37832 2453 37866
rect 2419 37758 2453 37792
rect 2419 37684 2453 37718
rect 2419 37610 2453 37644
rect 2419 37536 2453 37570
rect 2419 37462 2453 37496
rect 2419 37388 2453 37422
rect 2419 37314 2453 37348
rect 2419 37240 2453 37274
rect 2419 37166 2453 37200
rect 2419 37092 2453 37126
rect 2419 37018 2453 37052
rect 2655 38930 2689 38964
rect 2655 38857 2689 38891
rect 2655 38784 2689 38818
rect 2655 38711 2689 38745
rect 2655 38638 2689 38672
rect 2655 38565 2689 38599
rect 2655 38492 2689 38526
rect 2655 38419 2689 38453
rect 2655 38346 2689 38380
rect 2655 38273 2689 38307
rect 2655 38200 2689 38234
rect 2655 38127 2689 38161
rect 2655 38054 2689 38088
rect 2655 37980 2689 38014
rect 2655 37906 2689 37940
rect 2655 37832 2689 37866
rect 2655 37758 2689 37792
rect 2655 37684 2689 37718
rect 2655 37610 2689 37644
rect 2655 37536 2689 37570
rect 2655 37462 2689 37496
rect 2655 37388 2689 37422
rect 2655 37314 2689 37348
rect 2655 37240 2689 37274
rect 2655 37166 2689 37200
rect 2655 37092 2689 37126
rect 2655 37018 2689 37052
rect 2891 38930 2925 38964
rect 2891 38857 2925 38891
rect 2891 38784 2925 38818
rect 2891 38711 2925 38745
rect 2891 38638 2925 38672
rect 2891 38565 2925 38599
rect 2891 38492 2925 38526
rect 2891 38419 2925 38453
rect 2891 38346 2925 38380
rect 2891 38273 2925 38307
rect 2891 38200 2925 38234
rect 2891 38127 2925 38161
rect 2891 38054 2925 38088
rect 2891 37980 2925 38014
rect 2891 37906 2925 37940
rect 2891 37832 2925 37866
rect 2891 37758 2925 37792
rect 2891 37684 2925 37718
rect 2891 37610 2925 37644
rect 2891 37536 2925 37570
rect 2891 37462 2925 37496
rect 2891 37388 2925 37422
rect 2891 37314 2925 37348
rect 2891 37240 2925 37274
rect 2891 37166 2925 37200
rect 2891 37092 2925 37126
rect 2891 37018 2925 37052
rect 3036 38940 3070 38962
rect 3036 38928 3070 38940
rect 3036 38872 3070 38890
rect 3036 38856 3070 38872
rect 3036 38804 3070 38818
rect 3036 38784 3070 38804
rect 3036 38736 3070 38746
rect 3036 38712 3070 38736
rect 3036 38668 3070 38674
rect 3036 38640 3070 38668
rect 3036 38600 3070 38602
rect 3036 38568 3070 38600
rect 3036 38498 3070 38530
rect 3036 38496 3070 38498
rect 3036 38430 3070 38458
rect 3036 38424 3070 38430
rect 3036 38362 3070 38386
rect 3036 38352 3070 38362
rect 3036 38294 3070 38314
rect 3036 38280 3070 38294
rect 3036 38226 3070 38242
rect 3036 38208 3070 38226
rect 3036 38158 3070 38170
rect 3036 38136 3070 38158
rect 3036 38090 3070 38098
rect 3036 38064 3070 38090
rect 3036 38022 3070 38026
rect 3036 37992 3070 38022
rect 3036 37920 3070 37954
rect 3036 37852 3070 37882
rect 3036 37848 3070 37852
rect 3036 37784 3070 37810
rect 3036 37776 3070 37784
rect 3036 37716 3070 37738
rect 3036 37704 3070 37716
rect 3036 37648 3070 37666
rect 3036 37632 3070 37648
rect 3036 37580 3070 37594
rect 3036 37560 3070 37580
rect 3036 37512 3070 37522
rect 3036 37488 3070 37512
rect 3036 37444 3070 37450
rect 3036 37416 3070 37444
rect 3036 37376 3070 37378
rect 3036 37344 3070 37376
rect 3036 37274 3070 37306
rect 3036 37272 3070 37274
rect 3036 37206 3070 37234
rect 3036 37200 3070 37206
rect 3036 37138 3070 37162
rect 3036 37128 3070 37138
rect 3036 37070 3070 37090
rect 3036 37056 3070 37070
rect 386 36981 420 36999
rect 386 36965 420 36981
rect 386 36913 420 36927
rect 386 36893 420 36913
rect 3036 37002 3070 37018
rect 3036 36984 3070 37002
rect 625 36890 626 36924
rect 626 36890 659 36924
rect 700 36890 732 36924
rect 732 36890 734 36924
rect 775 36890 802 36924
rect 802 36890 809 36924
rect 850 36890 872 36924
rect 872 36890 884 36924
rect 925 36890 942 36924
rect 942 36890 959 36924
rect 1000 36890 1012 36924
rect 1012 36890 1034 36924
rect 1075 36890 1082 36924
rect 1082 36890 1109 36924
rect 1150 36890 1152 36924
rect 1152 36890 1184 36924
rect 1225 36890 1256 36924
rect 1256 36890 1259 36924
rect 1300 36890 1326 36924
rect 1326 36890 1334 36924
rect 1375 36890 1396 36924
rect 1396 36890 1409 36924
rect 1450 36890 1466 36924
rect 1466 36890 1484 36924
rect 1525 36890 1536 36924
rect 1536 36890 1559 36924
rect 1600 36890 1606 36924
rect 1606 36890 1634 36924
rect 1674 36890 1676 36924
rect 1676 36890 1708 36924
rect 1748 36890 1782 36924
rect 1822 36890 1852 36924
rect 1852 36890 1856 36924
rect 1896 36890 1922 36924
rect 1922 36890 1930 36924
rect 1970 36890 1992 36924
rect 1992 36890 2004 36924
rect 2044 36890 2062 36924
rect 2062 36890 2078 36924
rect 2118 36890 2132 36924
rect 2132 36890 2152 36924
rect 2192 36890 2202 36924
rect 2202 36890 2226 36924
rect 2266 36890 2272 36924
rect 2272 36890 2300 36924
rect 2340 36890 2342 36924
rect 2342 36890 2374 36924
rect 2414 36890 2446 36924
rect 2446 36890 2448 36924
rect 2488 36890 2516 36924
rect 2516 36890 2522 36924
rect 2562 36890 2586 36924
rect 2586 36890 2596 36924
rect 2636 36890 2656 36924
rect 2656 36890 2670 36924
rect 2710 36890 2726 36924
rect 2726 36890 2744 36924
rect 2784 36890 2795 36924
rect 2795 36890 2818 36924
rect 3036 36934 3070 36946
rect 3036 36912 3070 36934
rect 386 36845 420 36855
rect 386 36821 420 36845
rect 3036 36866 3070 36874
rect 3036 36840 3070 36866
rect 386 36777 420 36783
rect 386 36749 420 36777
rect 386 36709 420 36711
rect 386 36677 420 36709
rect 386 36607 420 36639
rect 386 36605 420 36607
rect 386 36539 420 36567
rect 386 36533 420 36539
rect 386 36471 420 36495
rect 386 36461 420 36471
rect 386 36403 420 36423
rect 386 36389 420 36403
rect 386 36335 420 36351
rect 386 36317 420 36335
rect 386 36267 420 36279
rect 386 36245 420 36267
rect 386 36199 420 36207
rect 386 36173 420 36199
rect 386 36131 420 36135
rect 386 36101 420 36131
rect 386 36029 420 36063
rect 386 35961 420 35991
rect 386 35957 420 35961
rect 386 35893 420 35919
rect 386 35885 420 35893
rect 386 35825 420 35847
rect 386 35813 420 35825
rect 386 35757 420 35775
rect 386 35741 420 35757
rect 386 35689 420 35703
rect 386 35669 420 35689
rect 386 35621 420 35631
rect 386 35597 420 35621
rect 386 35553 420 35559
rect 386 35525 420 35553
rect 386 35485 420 35487
rect 386 35453 420 35485
rect 386 35383 420 35415
rect 386 35381 420 35383
rect 386 35315 420 35343
rect 386 35309 420 35315
rect 386 35247 420 35271
rect 386 35237 420 35247
rect 386 35179 420 35199
rect 386 35165 420 35179
rect 386 35111 420 35127
rect 386 35093 420 35111
rect 386 35043 420 35055
rect 386 35021 420 35043
rect 386 34975 420 34983
rect 386 34949 420 34975
rect 386 34907 420 34911
rect 386 34877 420 34907
rect 531 36788 565 36822
rect 531 36715 565 36749
rect 531 36642 565 36676
rect 531 36569 565 36603
rect 531 36496 565 36530
rect 531 36423 565 36457
rect 531 36350 565 36384
rect 531 36277 565 36311
rect 531 36204 565 36238
rect 531 36131 565 36165
rect 531 36058 565 36092
rect 531 35985 565 36019
rect 531 35912 565 35946
rect 531 35838 565 35872
rect 531 35764 565 35798
rect 531 35690 565 35724
rect 531 35616 565 35650
rect 531 35542 565 35576
rect 531 35468 565 35502
rect 531 35394 565 35428
rect 531 35320 565 35354
rect 531 35246 565 35280
rect 531 35172 565 35206
rect 531 35098 565 35132
rect 531 35024 565 35058
rect 531 34950 565 34984
rect 531 34876 565 34910
rect 767 36788 801 36822
rect 767 36715 801 36749
rect 767 36642 801 36676
rect 767 36569 801 36603
rect 767 36496 801 36530
rect 767 36423 801 36457
rect 767 36350 801 36384
rect 767 36277 801 36311
rect 767 36204 801 36238
rect 767 36131 801 36165
rect 767 36058 801 36092
rect 767 35985 801 36019
rect 767 35912 801 35946
rect 767 35838 801 35872
rect 767 35764 801 35798
rect 767 35690 801 35724
rect 767 35616 801 35650
rect 767 35542 801 35576
rect 767 35468 801 35502
rect 767 35394 801 35428
rect 767 35320 801 35354
rect 767 35246 801 35280
rect 767 35172 801 35206
rect 767 35098 801 35132
rect 767 35024 801 35058
rect 767 34950 801 34984
rect 767 34876 801 34910
rect 1003 36788 1037 36822
rect 1003 36715 1037 36749
rect 1003 36642 1037 36676
rect 1003 36569 1037 36603
rect 1003 36496 1037 36530
rect 1003 36423 1037 36457
rect 1003 36350 1037 36384
rect 1003 36277 1037 36311
rect 1003 36204 1037 36238
rect 1003 36131 1037 36165
rect 1003 36058 1037 36092
rect 1003 35985 1037 36019
rect 1003 35912 1037 35946
rect 1003 35838 1037 35872
rect 1003 35764 1037 35798
rect 1003 35690 1037 35724
rect 1003 35616 1037 35650
rect 1003 35542 1037 35576
rect 1003 35468 1037 35502
rect 1003 35394 1037 35428
rect 1003 35320 1037 35354
rect 1003 35246 1037 35280
rect 1003 35172 1037 35206
rect 1003 35098 1037 35132
rect 1003 35024 1037 35058
rect 1003 34950 1037 34984
rect 1003 34876 1037 34910
rect 1239 36788 1273 36822
rect 1239 36715 1273 36749
rect 1239 36642 1273 36676
rect 1239 36569 1273 36603
rect 1239 36496 1273 36530
rect 1239 36423 1273 36457
rect 1239 36350 1273 36384
rect 1239 36277 1273 36311
rect 1239 36204 1273 36238
rect 1239 36131 1273 36165
rect 1239 36058 1273 36092
rect 1239 35985 1273 36019
rect 1239 35912 1273 35946
rect 1239 35838 1273 35872
rect 1239 35764 1273 35798
rect 1239 35690 1273 35724
rect 1239 35616 1273 35650
rect 1239 35542 1273 35576
rect 1239 35468 1273 35502
rect 1239 35394 1273 35428
rect 1239 35320 1273 35354
rect 1239 35246 1273 35280
rect 1239 35172 1273 35206
rect 1239 35098 1273 35132
rect 1239 35024 1273 35058
rect 1239 34950 1273 34984
rect 1239 34876 1273 34910
rect 1475 36788 1509 36822
rect 1475 36715 1509 36749
rect 1475 36642 1509 36676
rect 1475 36569 1509 36603
rect 1475 36496 1509 36530
rect 1475 36423 1509 36457
rect 1475 36350 1509 36384
rect 1475 36277 1509 36311
rect 1475 36204 1509 36238
rect 1475 36131 1509 36165
rect 1475 36058 1509 36092
rect 1475 35985 1509 36019
rect 1475 35912 1509 35946
rect 1475 35838 1509 35872
rect 1475 35764 1509 35798
rect 1475 35690 1509 35724
rect 1475 35616 1509 35650
rect 1475 35542 1509 35576
rect 1475 35468 1509 35502
rect 1475 35394 1509 35428
rect 1475 35320 1509 35354
rect 1475 35246 1509 35280
rect 1475 35172 1509 35206
rect 1475 35098 1509 35132
rect 1475 35024 1509 35058
rect 1475 34950 1509 34984
rect 1475 34876 1509 34910
rect 1711 36788 1745 36822
rect 1711 36715 1745 36749
rect 1711 36642 1745 36676
rect 1711 36569 1745 36603
rect 1711 36496 1745 36530
rect 1711 36423 1745 36457
rect 1711 36350 1745 36384
rect 1711 36277 1745 36311
rect 1711 36204 1745 36238
rect 1711 36131 1745 36165
rect 1711 36058 1745 36092
rect 1711 35985 1745 36019
rect 1711 35912 1745 35946
rect 1711 35838 1745 35872
rect 1711 35764 1745 35798
rect 1711 35690 1745 35724
rect 1711 35616 1745 35650
rect 1711 35542 1745 35576
rect 1711 35468 1745 35502
rect 1711 35394 1745 35428
rect 1711 35320 1745 35354
rect 1711 35246 1745 35280
rect 1711 35172 1745 35206
rect 1711 35098 1745 35132
rect 1711 35024 1745 35058
rect 1711 34950 1745 34984
rect 1711 34876 1745 34910
rect 1947 36788 1981 36822
rect 1947 36715 1981 36749
rect 1947 36642 1981 36676
rect 1947 36569 1981 36603
rect 1947 36496 1981 36530
rect 1947 36423 1981 36457
rect 1947 36350 1981 36384
rect 1947 36277 1981 36311
rect 1947 36204 1981 36238
rect 1947 36131 1981 36165
rect 1947 36058 1981 36092
rect 1947 35985 1981 36019
rect 1947 35912 1981 35946
rect 1947 35838 1981 35872
rect 1947 35764 1981 35798
rect 1947 35690 1981 35724
rect 1947 35616 1981 35650
rect 1947 35542 1981 35576
rect 1947 35468 1981 35502
rect 1947 35394 1981 35428
rect 1947 35320 1981 35354
rect 1947 35246 1981 35280
rect 1947 35172 1981 35206
rect 1947 35098 1981 35132
rect 1947 35024 1981 35058
rect 1947 34950 1981 34984
rect 1947 34876 1981 34910
rect 2183 36788 2217 36822
rect 2183 36715 2217 36749
rect 2183 36642 2217 36676
rect 2183 36569 2217 36603
rect 2183 36496 2217 36530
rect 2183 36423 2217 36457
rect 2183 36350 2217 36384
rect 2183 36277 2217 36311
rect 2183 36204 2217 36238
rect 2183 36131 2217 36165
rect 2183 36058 2217 36092
rect 2183 35985 2217 36019
rect 2183 35912 2217 35946
rect 2183 35838 2217 35872
rect 2183 35764 2217 35798
rect 2183 35690 2217 35724
rect 2183 35616 2217 35650
rect 2183 35542 2217 35576
rect 2183 35468 2217 35502
rect 2183 35394 2217 35428
rect 2183 35320 2217 35354
rect 2183 35246 2217 35280
rect 2183 35172 2217 35206
rect 2183 35098 2217 35132
rect 2183 35024 2217 35058
rect 2183 34950 2217 34984
rect 2183 34876 2217 34910
rect 2419 36788 2453 36822
rect 2419 36715 2453 36749
rect 2419 36642 2453 36676
rect 2419 36569 2453 36603
rect 2419 36496 2453 36530
rect 2419 36423 2453 36457
rect 2419 36350 2453 36384
rect 2419 36277 2453 36311
rect 2419 36204 2453 36238
rect 2419 36131 2453 36165
rect 2419 36058 2453 36092
rect 2419 35985 2453 36019
rect 2419 35912 2453 35946
rect 2419 35838 2453 35872
rect 2419 35764 2453 35798
rect 2419 35690 2453 35724
rect 2419 35616 2453 35650
rect 2419 35542 2453 35576
rect 2419 35468 2453 35502
rect 2419 35394 2453 35428
rect 2419 35320 2453 35354
rect 2419 35246 2453 35280
rect 2419 35172 2453 35206
rect 2419 35098 2453 35132
rect 2419 35024 2453 35058
rect 2419 34950 2453 34984
rect 2419 34876 2453 34910
rect 2655 36788 2689 36822
rect 2655 36715 2689 36749
rect 2655 36642 2689 36676
rect 2655 36569 2689 36603
rect 2655 36496 2689 36530
rect 2655 36423 2689 36457
rect 2655 36350 2689 36384
rect 2655 36277 2689 36311
rect 2655 36204 2689 36238
rect 2655 36131 2689 36165
rect 2655 36058 2689 36092
rect 2655 35985 2689 36019
rect 2655 35912 2689 35946
rect 2655 35838 2689 35872
rect 2655 35764 2689 35798
rect 2655 35690 2689 35724
rect 2655 35616 2689 35650
rect 2655 35542 2689 35576
rect 2655 35468 2689 35502
rect 2655 35394 2689 35428
rect 2655 35320 2689 35354
rect 2655 35246 2689 35280
rect 2655 35172 2689 35206
rect 2655 35098 2689 35132
rect 2655 35024 2689 35058
rect 2655 34950 2689 34984
rect 2655 34876 2689 34910
rect 2891 36788 2925 36822
rect 2891 36715 2925 36749
rect 2891 36642 2925 36676
rect 2891 36569 2925 36603
rect 2891 36496 2925 36530
rect 2891 36423 2925 36457
rect 2891 36350 2925 36384
rect 2891 36277 2925 36311
rect 2891 36204 2925 36238
rect 2891 36131 2925 36165
rect 2891 36058 2925 36092
rect 2891 35985 2925 36019
rect 2891 35912 2925 35946
rect 2891 35838 2925 35872
rect 2891 35764 2925 35798
rect 2891 35690 2925 35724
rect 2891 35616 2925 35650
rect 2891 35542 2925 35576
rect 2891 35468 2925 35502
rect 2891 35394 2925 35428
rect 2891 35320 2925 35354
rect 2891 35246 2925 35280
rect 2891 35172 2925 35206
rect 2891 35098 2925 35132
rect 2891 35024 2925 35058
rect 2891 34950 2925 34984
rect 2891 34876 2925 34910
rect 3036 36798 3070 36802
rect 3036 36768 3070 36798
rect 3036 36696 3070 36730
rect 3036 36628 3070 36658
rect 3036 36624 3070 36628
rect 3036 36560 3070 36586
rect 3036 36552 3070 36560
rect 3036 36492 3070 36514
rect 3036 36480 3070 36492
rect 3036 36424 3070 36442
rect 3036 36408 3070 36424
rect 3036 36356 3070 36370
rect 3036 36336 3070 36356
rect 3036 36288 3070 36298
rect 3036 36264 3070 36288
rect 3036 36220 3070 36226
rect 3036 36192 3070 36220
rect 3036 36152 3070 36154
rect 3036 36120 3070 36152
rect 3036 36050 3070 36082
rect 3036 36048 3070 36050
rect 3036 35982 3070 36010
rect 3036 35976 3070 35982
rect 3036 35914 3070 35938
rect 3036 35904 3070 35914
rect 3036 35846 3070 35866
rect 3036 35832 3070 35846
rect 3036 35778 3070 35794
rect 3036 35760 3070 35778
rect 3036 35710 3070 35722
rect 3036 35688 3070 35710
rect 3036 35642 3070 35650
rect 3036 35616 3070 35642
rect 3036 35574 3070 35578
rect 3036 35544 3070 35574
rect 3036 35472 3070 35506
rect 3036 35404 3070 35434
rect 3036 35400 3070 35404
rect 3036 35336 3070 35362
rect 3036 35328 3070 35336
rect 3036 35268 3070 35290
rect 3036 35256 3070 35268
rect 3036 35200 3070 35218
rect 3036 35184 3070 35200
rect 3036 35132 3070 35146
rect 3036 35112 3070 35132
rect 3036 35064 3070 35074
rect 3036 35040 3070 35064
rect 3036 34996 3070 35002
rect 3036 34968 3070 34996
rect 3036 34928 3070 34930
rect 3036 34896 3070 34928
rect 386 34805 420 34839
rect 386 34737 420 34767
rect 386 34733 420 34737
rect 625 34760 626 34794
rect 626 34760 659 34794
rect 700 34760 732 34794
rect 732 34760 734 34794
rect 775 34760 802 34794
rect 802 34760 809 34794
rect 850 34760 872 34794
rect 872 34760 884 34794
rect 925 34760 942 34794
rect 942 34760 959 34794
rect 1000 34760 1012 34794
rect 1012 34760 1034 34794
rect 1075 34760 1082 34794
rect 1082 34760 1109 34794
rect 1150 34760 1152 34794
rect 1152 34760 1184 34794
rect 1225 34760 1256 34794
rect 1256 34760 1259 34794
rect 1300 34760 1326 34794
rect 1326 34760 1334 34794
rect 1375 34760 1396 34794
rect 1396 34760 1409 34794
rect 1450 34760 1466 34794
rect 1466 34760 1484 34794
rect 1525 34760 1536 34794
rect 1536 34760 1559 34794
rect 1600 34760 1606 34794
rect 1606 34760 1634 34794
rect 1674 34760 1676 34794
rect 1676 34760 1708 34794
rect 1748 34760 1782 34794
rect 1822 34760 1852 34794
rect 1852 34760 1856 34794
rect 1896 34760 1922 34794
rect 1922 34760 1930 34794
rect 1970 34760 1992 34794
rect 1992 34760 2004 34794
rect 2044 34760 2062 34794
rect 2062 34760 2078 34794
rect 2118 34760 2132 34794
rect 2132 34760 2152 34794
rect 2192 34760 2202 34794
rect 2202 34760 2226 34794
rect 2266 34760 2272 34794
rect 2272 34760 2300 34794
rect 2340 34760 2342 34794
rect 2342 34760 2374 34794
rect 2414 34760 2446 34794
rect 2446 34760 2448 34794
rect 2488 34760 2516 34794
rect 2516 34760 2522 34794
rect 2562 34760 2586 34794
rect 2586 34760 2596 34794
rect 2636 34760 2656 34794
rect 2656 34760 2670 34794
rect 2710 34760 2726 34794
rect 2726 34760 2744 34794
rect 2784 34760 2795 34794
rect 2795 34760 2818 34794
rect 3036 34826 3070 34858
rect 3036 34824 3070 34826
rect 386 34669 420 34695
rect 386 34661 420 34669
rect 3036 34758 3070 34786
rect 3036 34752 3070 34758
rect 386 34601 420 34623
rect 386 34589 420 34601
rect 386 34533 420 34551
rect 386 34517 420 34533
rect 386 34465 420 34479
rect 386 34445 420 34465
rect 386 34397 420 34407
rect 386 34373 420 34397
rect 386 34329 420 34335
rect 386 34301 420 34329
rect 386 34261 420 34263
rect 386 34229 420 34261
rect 386 34159 420 34191
rect 386 34157 420 34159
rect 386 34091 420 34119
rect 386 34085 420 34091
rect 386 34023 420 34047
rect 386 34013 420 34023
rect 386 33955 420 33975
rect 386 33941 420 33955
rect 386 33887 420 33903
rect 386 33869 420 33887
rect 386 33819 420 33831
rect 386 33797 420 33819
rect 386 33751 420 33759
rect 386 33725 420 33751
rect 386 33683 420 33687
rect 386 33653 420 33683
rect 386 33581 420 33615
rect 386 33513 420 33543
rect 386 33509 420 33513
rect 386 33445 420 33471
rect 386 33437 420 33445
rect 386 33377 420 33399
rect 386 33365 420 33377
rect 386 33309 420 33327
rect 386 33293 420 33309
rect 386 33241 420 33255
rect 386 33221 420 33241
rect 386 33173 420 33183
rect 386 33149 420 33173
rect 386 33105 420 33111
rect 386 33077 420 33105
rect 386 33037 420 33039
rect 386 33005 420 33037
rect 386 32935 420 32967
rect 386 32933 420 32935
rect 386 32867 420 32895
rect 386 32861 420 32867
rect 386 32799 420 32823
rect 386 32789 420 32799
rect 386 32731 420 32751
rect 386 32717 420 32731
rect 531 34658 565 34692
rect 531 34585 565 34619
rect 531 34512 565 34546
rect 531 34439 565 34473
rect 531 34366 565 34400
rect 531 34293 565 34327
rect 531 34220 565 34254
rect 531 34147 565 34181
rect 531 34074 565 34108
rect 531 34001 565 34035
rect 531 33928 565 33962
rect 531 33855 565 33889
rect 531 33782 565 33816
rect 531 33708 565 33742
rect 531 33634 565 33668
rect 531 33560 565 33594
rect 531 33486 565 33520
rect 531 33412 565 33446
rect 531 33338 565 33372
rect 531 33264 565 33298
rect 531 33190 565 33224
rect 531 33116 565 33150
rect 531 33042 565 33076
rect 531 32968 565 33002
rect 531 32894 565 32928
rect 531 32820 565 32854
rect 531 32746 565 32780
rect 767 34658 801 34692
rect 767 34585 801 34619
rect 767 34512 801 34546
rect 767 34439 801 34473
rect 767 34366 801 34400
rect 767 34293 801 34327
rect 767 34220 801 34254
rect 767 34147 801 34181
rect 767 34074 801 34108
rect 767 34001 801 34035
rect 767 33928 801 33962
rect 767 33855 801 33889
rect 767 33782 801 33816
rect 767 33708 801 33742
rect 767 33634 801 33668
rect 767 33560 801 33594
rect 767 33486 801 33520
rect 767 33412 801 33446
rect 767 33338 801 33372
rect 767 33264 801 33298
rect 767 33190 801 33224
rect 767 33116 801 33150
rect 767 33042 801 33076
rect 767 32968 801 33002
rect 767 32894 801 32928
rect 767 32820 801 32854
rect 767 32746 801 32780
rect 1003 34658 1037 34692
rect 1003 34585 1037 34619
rect 1003 34512 1037 34546
rect 1003 34439 1037 34473
rect 1003 34366 1037 34400
rect 1003 34293 1037 34327
rect 1003 34220 1037 34254
rect 1003 34147 1037 34181
rect 1003 34074 1037 34108
rect 1003 34001 1037 34035
rect 1003 33928 1037 33962
rect 1003 33855 1037 33889
rect 1003 33782 1037 33816
rect 1003 33708 1037 33742
rect 1003 33634 1037 33668
rect 1003 33560 1037 33594
rect 1003 33486 1037 33520
rect 1003 33412 1037 33446
rect 1003 33338 1037 33372
rect 1003 33264 1037 33298
rect 1003 33190 1037 33224
rect 1003 33116 1037 33150
rect 1003 33042 1037 33076
rect 1003 32968 1037 33002
rect 1003 32894 1037 32928
rect 1003 32820 1037 32854
rect 1003 32746 1037 32780
rect 1239 34658 1273 34692
rect 1239 34585 1273 34619
rect 1239 34512 1273 34546
rect 1239 34439 1273 34473
rect 1239 34366 1273 34400
rect 1239 34293 1273 34327
rect 1239 34220 1273 34254
rect 1239 34147 1273 34181
rect 1239 34074 1273 34108
rect 1239 34001 1273 34035
rect 1239 33928 1273 33962
rect 1239 33855 1273 33889
rect 1239 33782 1273 33816
rect 1239 33708 1273 33742
rect 1239 33634 1273 33668
rect 1239 33560 1273 33594
rect 1239 33486 1273 33520
rect 1239 33412 1273 33446
rect 1239 33338 1273 33372
rect 1239 33264 1273 33298
rect 1239 33190 1273 33224
rect 1239 33116 1273 33150
rect 1239 33042 1273 33076
rect 1239 32968 1273 33002
rect 1239 32894 1273 32928
rect 1239 32820 1273 32854
rect 1239 32746 1273 32780
rect 1475 34658 1509 34692
rect 1475 34585 1509 34619
rect 1475 34512 1509 34546
rect 1475 34439 1509 34473
rect 1475 34366 1509 34400
rect 1475 34293 1509 34327
rect 1475 34220 1509 34254
rect 1475 34147 1509 34181
rect 1475 34074 1509 34108
rect 1475 34001 1509 34035
rect 1475 33928 1509 33962
rect 1475 33855 1509 33889
rect 1475 33782 1509 33816
rect 1475 33708 1509 33742
rect 1475 33634 1509 33668
rect 1475 33560 1509 33594
rect 1475 33486 1509 33520
rect 1475 33412 1509 33446
rect 1475 33338 1509 33372
rect 1475 33264 1509 33298
rect 1475 33190 1509 33224
rect 1475 33116 1509 33150
rect 1475 33042 1509 33076
rect 1475 32968 1509 33002
rect 1475 32894 1509 32928
rect 1475 32820 1509 32854
rect 1475 32746 1509 32780
rect 1711 34658 1745 34692
rect 1711 34585 1745 34619
rect 1711 34512 1745 34546
rect 1711 34439 1745 34473
rect 1711 34366 1745 34400
rect 1711 34293 1745 34327
rect 1711 34220 1745 34254
rect 1711 34147 1745 34181
rect 1711 34074 1745 34108
rect 1711 34001 1745 34035
rect 1711 33928 1745 33962
rect 1711 33855 1745 33889
rect 1711 33782 1745 33816
rect 1711 33708 1745 33742
rect 1711 33634 1745 33668
rect 1711 33560 1745 33594
rect 1711 33486 1745 33520
rect 1711 33412 1745 33446
rect 1711 33338 1745 33372
rect 1711 33264 1745 33298
rect 1711 33190 1745 33224
rect 1711 33116 1745 33150
rect 1711 33042 1745 33076
rect 1711 32968 1745 33002
rect 1711 32894 1745 32928
rect 1711 32820 1745 32854
rect 1711 32746 1745 32780
rect 1947 34658 1981 34692
rect 1947 34585 1981 34619
rect 1947 34512 1981 34546
rect 1947 34439 1981 34473
rect 1947 34366 1981 34400
rect 1947 34293 1981 34327
rect 1947 34220 1981 34254
rect 1947 34147 1981 34181
rect 1947 34074 1981 34108
rect 1947 34001 1981 34035
rect 1947 33928 1981 33962
rect 1947 33855 1981 33889
rect 1947 33782 1981 33816
rect 1947 33708 1981 33742
rect 1947 33634 1981 33668
rect 1947 33560 1981 33594
rect 1947 33486 1981 33520
rect 1947 33412 1981 33446
rect 1947 33338 1981 33372
rect 1947 33264 1981 33298
rect 1947 33190 1981 33224
rect 1947 33116 1981 33150
rect 1947 33042 1981 33076
rect 1947 32968 1981 33002
rect 1947 32894 1981 32928
rect 1947 32820 1981 32854
rect 1947 32746 1981 32780
rect 2183 34658 2217 34692
rect 2183 34585 2217 34619
rect 2183 34512 2217 34546
rect 2183 34439 2217 34473
rect 2183 34366 2217 34400
rect 2183 34293 2217 34327
rect 2183 34220 2217 34254
rect 2183 34147 2217 34181
rect 2183 34074 2217 34108
rect 2183 34001 2217 34035
rect 2183 33928 2217 33962
rect 2183 33855 2217 33889
rect 2183 33782 2217 33816
rect 2183 33708 2217 33742
rect 2183 33634 2217 33668
rect 2183 33560 2217 33594
rect 2183 33486 2217 33520
rect 2183 33412 2217 33446
rect 2183 33338 2217 33372
rect 2183 33264 2217 33298
rect 2183 33190 2217 33224
rect 2183 33116 2217 33150
rect 2183 33042 2217 33076
rect 2183 32968 2217 33002
rect 2183 32894 2217 32928
rect 2183 32820 2217 32854
rect 2183 32746 2217 32780
rect 2419 34658 2453 34692
rect 2419 34585 2453 34619
rect 2419 34512 2453 34546
rect 2419 34439 2453 34473
rect 2419 34366 2453 34400
rect 2419 34293 2453 34327
rect 2419 34220 2453 34254
rect 2419 34147 2453 34181
rect 2419 34074 2453 34108
rect 2419 34001 2453 34035
rect 2419 33928 2453 33962
rect 2419 33855 2453 33889
rect 2419 33782 2453 33816
rect 2419 33708 2453 33742
rect 2419 33634 2453 33668
rect 2419 33560 2453 33594
rect 2419 33486 2453 33520
rect 2419 33412 2453 33446
rect 2419 33338 2453 33372
rect 2419 33264 2453 33298
rect 2419 33190 2453 33224
rect 2419 33116 2453 33150
rect 2419 33042 2453 33076
rect 2419 32968 2453 33002
rect 2419 32894 2453 32928
rect 2419 32820 2453 32854
rect 2419 32746 2453 32780
rect 2655 34658 2689 34692
rect 2655 34585 2689 34619
rect 2655 34512 2689 34546
rect 2655 34439 2689 34473
rect 2655 34366 2689 34400
rect 2655 34293 2689 34327
rect 2655 34220 2689 34254
rect 2655 34147 2689 34181
rect 2655 34074 2689 34108
rect 2655 34001 2689 34035
rect 2655 33928 2689 33962
rect 2655 33855 2689 33889
rect 2655 33782 2689 33816
rect 2655 33708 2689 33742
rect 2655 33634 2689 33668
rect 2655 33560 2689 33594
rect 2655 33486 2689 33520
rect 2655 33412 2689 33446
rect 2655 33338 2689 33372
rect 2655 33264 2689 33298
rect 2655 33190 2689 33224
rect 2655 33116 2689 33150
rect 2655 33042 2689 33076
rect 2655 32968 2689 33002
rect 2655 32894 2689 32928
rect 2655 32820 2689 32854
rect 2655 32746 2689 32780
rect 2891 34658 2925 34692
rect 2891 34585 2925 34619
rect 2891 34512 2925 34546
rect 2891 34439 2925 34473
rect 2891 34366 2925 34400
rect 2891 34293 2925 34327
rect 2891 34220 2925 34254
rect 2891 34147 2925 34181
rect 2891 34074 2925 34108
rect 2891 34001 2925 34035
rect 2891 33928 2925 33962
rect 2891 33855 2925 33889
rect 2891 33782 2925 33816
rect 2891 33708 2925 33742
rect 2891 33634 2925 33668
rect 2891 33560 2925 33594
rect 2891 33486 2925 33520
rect 2891 33412 2925 33446
rect 2891 33338 2925 33372
rect 2891 33264 2925 33298
rect 2891 33190 2925 33224
rect 2891 33116 2925 33150
rect 2891 33042 2925 33076
rect 2891 32968 2925 33002
rect 2891 32894 2925 32928
rect 2891 32820 2925 32854
rect 2891 32746 2925 32780
rect 3036 34690 3070 34714
rect 3036 34680 3070 34690
rect 3036 34622 3070 34642
rect 3036 34608 3070 34622
rect 3036 34554 3070 34570
rect 3036 34536 3070 34554
rect 3036 34486 3070 34498
rect 3036 34464 3070 34486
rect 3036 34418 3070 34426
rect 3036 34392 3070 34418
rect 3036 34350 3070 34354
rect 3036 34320 3070 34350
rect 3036 34248 3070 34282
rect 3036 34180 3070 34210
rect 3036 34176 3070 34180
rect 3036 34112 3070 34138
rect 3036 34104 3070 34112
rect 3036 34044 3070 34066
rect 3036 34032 3070 34044
rect 3036 33976 3070 33994
rect 3036 33960 3070 33976
rect 3036 33908 3070 33922
rect 3036 33888 3070 33908
rect 3036 33840 3070 33850
rect 3036 33816 3070 33840
rect 3036 33772 3070 33778
rect 3036 33744 3070 33772
rect 3036 33704 3070 33706
rect 3036 33672 3070 33704
rect 3036 33602 3070 33634
rect 3036 33600 3070 33602
rect 3036 33534 3070 33562
rect 3036 33528 3070 33534
rect 3036 33466 3070 33490
rect 3036 33456 3070 33466
rect 3036 33398 3070 33418
rect 3036 33384 3070 33398
rect 3036 33330 3070 33346
rect 3036 33312 3070 33330
rect 3036 33262 3070 33274
rect 3036 33240 3070 33262
rect 3036 33194 3070 33202
rect 3036 33168 3070 33194
rect 3036 33126 3070 33130
rect 3036 33096 3070 33126
rect 3036 33024 3070 33058
rect 3036 32956 3070 32986
rect 3036 32952 3070 32956
rect 3036 32888 3070 32914
rect 3036 32880 3070 32888
rect 3036 32820 3070 32842
rect 3036 32808 3070 32820
rect 386 32663 420 32679
rect 386 32645 420 32663
rect 3036 32752 3070 32770
rect 3036 32736 3070 32752
rect 3036 32684 3070 32698
rect 3036 32664 3070 32684
rect 625 32630 626 32664
rect 626 32630 659 32664
rect 700 32630 732 32664
rect 732 32630 734 32664
rect 775 32630 802 32664
rect 802 32630 809 32664
rect 850 32630 872 32664
rect 872 32630 884 32664
rect 925 32630 942 32664
rect 942 32630 959 32664
rect 1000 32630 1012 32664
rect 1012 32630 1034 32664
rect 1075 32630 1082 32664
rect 1082 32630 1109 32664
rect 1150 32630 1152 32664
rect 1152 32630 1184 32664
rect 1225 32630 1256 32664
rect 1256 32630 1259 32664
rect 1300 32630 1326 32664
rect 1326 32630 1334 32664
rect 1375 32630 1396 32664
rect 1396 32630 1409 32664
rect 1450 32630 1466 32664
rect 1466 32630 1484 32664
rect 1525 32630 1536 32664
rect 1536 32630 1559 32664
rect 1600 32630 1606 32664
rect 1606 32630 1634 32664
rect 1674 32630 1676 32664
rect 1676 32630 1708 32664
rect 1748 32630 1782 32664
rect 1822 32630 1852 32664
rect 1852 32630 1856 32664
rect 1896 32630 1922 32664
rect 1922 32630 1930 32664
rect 1970 32630 1992 32664
rect 1992 32630 2004 32664
rect 2044 32630 2062 32664
rect 2062 32630 2078 32664
rect 2118 32630 2132 32664
rect 2132 32630 2152 32664
rect 2192 32630 2202 32664
rect 2202 32630 2226 32664
rect 2266 32630 2272 32664
rect 2272 32630 2300 32664
rect 2340 32630 2342 32664
rect 2342 32630 2374 32664
rect 2414 32630 2446 32664
rect 2446 32630 2448 32664
rect 2488 32630 2516 32664
rect 2516 32630 2522 32664
rect 2562 32630 2586 32664
rect 2586 32630 2596 32664
rect 2636 32630 2656 32664
rect 2656 32630 2670 32664
rect 2710 32630 2726 32664
rect 2726 32630 2744 32664
rect 2784 32630 2795 32664
rect 2795 32630 2818 32664
rect 386 32595 420 32607
rect 386 32573 420 32595
rect 3036 32616 3070 32626
rect 3036 32592 3070 32616
rect 386 32527 420 32535
rect 386 32501 420 32527
rect 386 32459 420 32463
rect 386 32429 420 32459
rect 386 32357 420 32391
rect 386 32289 420 32319
rect 386 32285 420 32289
rect 386 32221 420 32247
rect 386 32213 420 32221
rect 386 32153 420 32175
rect 386 32141 420 32153
rect 386 32085 420 32103
rect 386 32069 420 32085
rect 386 32017 420 32031
rect 386 31997 420 32017
rect 386 31949 420 31959
rect 386 31925 420 31949
rect 386 31881 420 31887
rect 386 31853 420 31881
rect 386 31813 420 31815
rect 386 31781 420 31813
rect 386 31711 420 31743
rect 386 31709 420 31711
rect 386 31643 420 31671
rect 386 31637 420 31643
rect 386 31575 420 31599
rect 386 31565 420 31575
rect 386 31507 420 31527
rect 386 31493 420 31507
rect 386 31439 420 31455
rect 386 31421 420 31439
rect 386 31371 420 31383
rect 386 31349 420 31371
rect 386 31303 420 31311
rect 386 31277 420 31303
rect 386 31235 420 31239
rect 386 31205 420 31235
rect 386 31133 420 31167
rect 386 31065 420 31095
rect 386 31061 420 31065
rect 386 30997 420 31023
rect 386 30989 420 30997
rect 386 30929 420 30951
rect 386 30917 420 30929
rect 386 30861 420 30879
rect 386 30845 420 30861
rect 386 30793 420 30807
rect 386 30773 420 30793
rect 386 30725 420 30735
rect 386 30701 420 30725
rect 386 30657 420 30663
rect 386 30629 420 30657
rect 386 30589 420 30591
rect 386 30557 420 30589
rect 531 32514 565 32548
rect 531 32441 565 32475
rect 531 32368 565 32402
rect 531 32295 565 32329
rect 531 32222 565 32256
rect 531 32149 565 32183
rect 531 32076 565 32110
rect 531 32003 565 32037
rect 531 31930 565 31964
rect 531 31857 565 31891
rect 531 31784 565 31818
rect 531 31711 565 31745
rect 531 31638 565 31672
rect 531 31564 565 31598
rect 531 31490 565 31524
rect 531 31416 565 31450
rect 531 31342 565 31376
rect 531 31268 565 31302
rect 531 31194 565 31228
rect 531 31120 565 31154
rect 531 31046 565 31080
rect 531 30972 565 31006
rect 531 30898 565 30932
rect 531 30824 565 30858
rect 531 30750 565 30784
rect 531 30676 565 30710
rect 531 30602 565 30636
rect 767 32514 801 32548
rect 767 32441 801 32475
rect 767 32368 801 32402
rect 767 32295 801 32329
rect 767 32222 801 32256
rect 767 32149 801 32183
rect 767 32076 801 32110
rect 767 32003 801 32037
rect 767 31930 801 31964
rect 767 31857 801 31891
rect 767 31784 801 31818
rect 767 31711 801 31745
rect 767 31638 801 31672
rect 767 31564 801 31598
rect 767 31490 801 31524
rect 767 31416 801 31450
rect 767 31342 801 31376
rect 767 31268 801 31302
rect 767 31194 801 31228
rect 767 31120 801 31154
rect 767 31046 801 31080
rect 767 30972 801 31006
rect 767 30898 801 30932
rect 767 30824 801 30858
rect 767 30750 801 30784
rect 767 30676 801 30710
rect 767 30602 801 30636
rect 1003 32514 1037 32548
rect 1003 32441 1037 32475
rect 1003 32368 1037 32402
rect 1003 32295 1037 32329
rect 1003 32222 1037 32256
rect 1003 32149 1037 32183
rect 1003 32076 1037 32110
rect 1003 32003 1037 32037
rect 1003 31930 1037 31964
rect 1003 31857 1037 31891
rect 1003 31784 1037 31818
rect 1003 31711 1037 31745
rect 1003 31638 1037 31672
rect 1003 31564 1037 31598
rect 1003 31490 1037 31524
rect 1003 31416 1037 31450
rect 1003 31342 1037 31376
rect 1003 31268 1037 31302
rect 1003 31194 1037 31228
rect 1003 31120 1037 31154
rect 1003 31046 1037 31080
rect 1003 30972 1037 31006
rect 1003 30898 1037 30932
rect 1003 30824 1037 30858
rect 1003 30750 1037 30784
rect 1003 30676 1037 30710
rect 1003 30602 1037 30636
rect 1239 32514 1273 32548
rect 1239 32441 1273 32475
rect 1239 32368 1273 32402
rect 1239 32295 1273 32329
rect 1239 32222 1273 32256
rect 1239 32149 1273 32183
rect 1239 32076 1273 32110
rect 1239 32003 1273 32037
rect 1239 31930 1273 31964
rect 1239 31857 1273 31891
rect 1239 31784 1273 31818
rect 1239 31711 1273 31745
rect 1239 31638 1273 31672
rect 1239 31564 1273 31598
rect 1239 31490 1273 31524
rect 1239 31416 1273 31450
rect 1239 31342 1273 31376
rect 1239 31268 1273 31302
rect 1239 31194 1273 31228
rect 1239 31120 1273 31154
rect 1239 31046 1273 31080
rect 1239 30972 1273 31006
rect 1239 30898 1273 30932
rect 1239 30824 1273 30858
rect 1239 30750 1273 30784
rect 1239 30676 1273 30710
rect 1239 30602 1273 30636
rect 1475 32514 1509 32548
rect 1475 32441 1509 32475
rect 1475 32368 1509 32402
rect 1475 32295 1509 32329
rect 1475 32222 1509 32256
rect 1475 32149 1509 32183
rect 1475 32076 1509 32110
rect 1475 32003 1509 32037
rect 1475 31930 1509 31964
rect 1475 31857 1509 31891
rect 1475 31784 1509 31818
rect 1475 31711 1509 31745
rect 1475 31638 1509 31672
rect 1475 31564 1509 31598
rect 1475 31490 1509 31524
rect 1475 31416 1509 31450
rect 1475 31342 1509 31376
rect 1475 31268 1509 31302
rect 1475 31194 1509 31228
rect 1475 31120 1509 31154
rect 1475 31046 1509 31080
rect 1475 30972 1509 31006
rect 1475 30898 1509 30932
rect 1475 30824 1509 30858
rect 1475 30750 1509 30784
rect 1475 30676 1509 30710
rect 1475 30602 1509 30636
rect 1711 32514 1745 32548
rect 1711 32441 1745 32475
rect 1711 32368 1745 32402
rect 1711 32295 1745 32329
rect 1711 32222 1745 32256
rect 1711 32149 1745 32183
rect 1711 32076 1745 32110
rect 1711 32003 1745 32037
rect 1711 31930 1745 31964
rect 1711 31857 1745 31891
rect 1711 31784 1745 31818
rect 1711 31711 1745 31745
rect 1711 31638 1745 31672
rect 1711 31564 1745 31598
rect 1711 31490 1745 31524
rect 1711 31416 1745 31450
rect 1711 31342 1745 31376
rect 1711 31268 1745 31302
rect 1711 31194 1745 31228
rect 1711 31120 1745 31154
rect 1711 31046 1745 31080
rect 1711 30972 1745 31006
rect 1711 30898 1745 30932
rect 1711 30824 1745 30858
rect 1711 30750 1745 30784
rect 1711 30676 1745 30710
rect 1711 30602 1745 30636
rect 1947 32514 1981 32548
rect 1947 32441 1981 32475
rect 1947 32368 1981 32402
rect 1947 32295 1981 32329
rect 1947 32222 1981 32256
rect 1947 32149 1981 32183
rect 1947 32076 1981 32110
rect 1947 32003 1981 32037
rect 1947 31930 1981 31964
rect 1947 31857 1981 31891
rect 1947 31784 1981 31818
rect 1947 31711 1981 31745
rect 1947 31638 1981 31672
rect 1947 31564 1981 31598
rect 1947 31490 1981 31524
rect 1947 31416 1981 31450
rect 1947 31342 1981 31376
rect 1947 31268 1981 31302
rect 1947 31194 1981 31228
rect 1947 31120 1981 31154
rect 1947 31046 1981 31080
rect 1947 30972 1981 31006
rect 1947 30898 1981 30932
rect 1947 30824 1981 30858
rect 1947 30750 1981 30784
rect 1947 30676 1981 30710
rect 1947 30602 1981 30636
rect 2183 32514 2217 32548
rect 2183 32441 2217 32475
rect 2183 32368 2217 32402
rect 2183 32295 2217 32329
rect 2183 32222 2217 32256
rect 2183 32149 2217 32183
rect 2183 32076 2217 32110
rect 2183 32003 2217 32037
rect 2183 31930 2217 31964
rect 2183 31857 2217 31891
rect 2183 31784 2217 31818
rect 2183 31711 2217 31745
rect 2183 31638 2217 31672
rect 2183 31564 2217 31598
rect 2183 31490 2217 31524
rect 2183 31416 2217 31450
rect 2183 31342 2217 31376
rect 2183 31268 2217 31302
rect 2183 31194 2217 31228
rect 2183 31120 2217 31154
rect 2183 31046 2217 31080
rect 2183 30972 2217 31006
rect 2183 30898 2217 30932
rect 2183 30824 2217 30858
rect 2183 30750 2217 30784
rect 2183 30676 2217 30710
rect 2183 30602 2217 30636
rect 2419 32514 2453 32548
rect 2419 32441 2453 32475
rect 2419 32368 2453 32402
rect 2419 32295 2453 32329
rect 2419 32222 2453 32256
rect 2419 32149 2453 32183
rect 2419 32076 2453 32110
rect 2419 32003 2453 32037
rect 2419 31930 2453 31964
rect 2419 31857 2453 31891
rect 2419 31784 2453 31818
rect 2419 31711 2453 31745
rect 2419 31638 2453 31672
rect 2419 31564 2453 31598
rect 2419 31490 2453 31524
rect 2419 31416 2453 31450
rect 2419 31342 2453 31376
rect 2419 31268 2453 31302
rect 2419 31194 2453 31228
rect 2419 31120 2453 31154
rect 2419 31046 2453 31080
rect 2419 30972 2453 31006
rect 2419 30898 2453 30932
rect 2419 30824 2453 30858
rect 2419 30750 2453 30784
rect 2419 30676 2453 30710
rect 2419 30602 2453 30636
rect 2655 32514 2689 32548
rect 2655 32441 2689 32475
rect 2655 32368 2689 32402
rect 2655 32295 2689 32329
rect 2655 32222 2689 32256
rect 2655 32149 2689 32183
rect 2655 32076 2689 32110
rect 2655 32003 2689 32037
rect 2655 31930 2689 31964
rect 2655 31857 2689 31891
rect 2655 31784 2689 31818
rect 2655 31711 2689 31745
rect 2655 31638 2689 31672
rect 2655 31564 2689 31598
rect 2655 31490 2689 31524
rect 2655 31416 2689 31450
rect 2655 31342 2689 31376
rect 2655 31268 2689 31302
rect 2655 31194 2689 31228
rect 2655 31120 2689 31154
rect 2655 31046 2689 31080
rect 2655 30972 2689 31006
rect 2655 30898 2689 30932
rect 2655 30824 2689 30858
rect 2655 30750 2689 30784
rect 2655 30676 2689 30710
rect 2655 30602 2689 30636
rect 2891 32514 2925 32548
rect 2891 32441 2925 32475
rect 2891 32368 2925 32402
rect 2891 32295 2925 32329
rect 2891 32222 2925 32256
rect 2891 32149 2925 32183
rect 2891 32076 2925 32110
rect 2891 32003 2925 32037
rect 2891 31930 2925 31964
rect 2891 31857 2925 31891
rect 2891 31784 2925 31818
rect 2891 31711 2925 31745
rect 2891 31638 2925 31672
rect 2891 31564 2925 31598
rect 2891 31490 2925 31524
rect 2891 31416 2925 31450
rect 2891 31342 2925 31376
rect 2891 31268 2925 31302
rect 2891 31194 2925 31228
rect 2891 31120 2925 31154
rect 2891 31046 2925 31080
rect 2891 30972 2925 31006
rect 2891 30898 2925 30932
rect 2891 30824 2925 30858
rect 2891 30750 2925 30784
rect 2891 30676 2925 30710
rect 2891 30602 2925 30636
rect 3036 32548 3070 32554
rect 3036 32520 3070 32548
rect 3036 32480 3070 32482
rect 3036 32448 3070 32480
rect 3036 32378 3070 32410
rect 3036 32376 3070 32378
rect 3036 32310 3070 32338
rect 3036 32304 3070 32310
rect 3036 32242 3070 32266
rect 3036 32232 3070 32242
rect 3036 32174 3070 32194
rect 3036 32160 3070 32174
rect 3036 32106 3070 32122
rect 3036 32088 3070 32106
rect 3036 32038 3070 32050
rect 3036 32016 3070 32038
rect 3036 31970 3070 31978
rect 3036 31944 3070 31970
rect 3036 31902 3070 31906
rect 3036 31872 3070 31902
rect 3036 31800 3070 31834
rect 3036 31732 3070 31762
rect 3036 31728 3070 31732
rect 3036 31664 3070 31690
rect 3036 31656 3070 31664
rect 3036 31596 3070 31618
rect 3036 31584 3070 31596
rect 3036 31528 3070 31546
rect 3036 31512 3070 31528
rect 3036 31460 3070 31474
rect 3036 31440 3070 31460
rect 3036 31392 3070 31402
rect 3036 31368 3070 31392
rect 3036 31324 3070 31330
rect 3036 31296 3070 31324
rect 3036 31256 3070 31258
rect 3036 31224 3070 31256
rect 3036 31154 3070 31186
rect 3036 31152 3070 31154
rect 3036 31086 3070 31114
rect 3036 31080 3070 31086
rect 3036 31018 3070 31042
rect 3036 31008 3070 31018
rect 3036 30950 3070 30970
rect 3036 30936 3070 30950
rect 3036 30882 3070 30898
rect 3036 30864 3070 30882
rect 3036 30814 3070 30826
rect 3036 30792 3070 30814
rect 3036 30746 3070 30754
rect 3036 30720 3070 30746
rect 3036 30678 3070 30682
rect 3036 30648 3070 30678
rect 3036 30576 3070 30610
rect 386 30487 420 30519
rect 386 30485 420 30487
rect 625 30500 626 30534
rect 626 30500 659 30534
rect 700 30500 732 30534
rect 732 30500 734 30534
rect 775 30500 802 30534
rect 802 30500 809 30534
rect 850 30500 872 30534
rect 872 30500 884 30534
rect 925 30500 942 30534
rect 942 30500 959 30534
rect 1000 30500 1012 30534
rect 1012 30500 1034 30534
rect 1075 30500 1082 30534
rect 1082 30500 1109 30534
rect 1150 30500 1152 30534
rect 1152 30500 1184 30534
rect 1225 30500 1256 30534
rect 1256 30500 1259 30534
rect 1300 30500 1326 30534
rect 1326 30500 1334 30534
rect 1375 30500 1396 30534
rect 1396 30500 1409 30534
rect 1450 30500 1466 30534
rect 1466 30500 1484 30534
rect 1525 30500 1536 30534
rect 1536 30500 1559 30534
rect 1600 30500 1606 30534
rect 1606 30500 1634 30534
rect 1674 30500 1676 30534
rect 1676 30500 1708 30534
rect 1748 30500 1782 30534
rect 1822 30500 1852 30534
rect 1852 30500 1856 30534
rect 1896 30500 1922 30534
rect 1922 30500 1930 30534
rect 1970 30500 1992 30534
rect 1992 30500 2004 30534
rect 2044 30500 2062 30534
rect 2062 30500 2078 30534
rect 2118 30500 2132 30534
rect 2132 30500 2152 30534
rect 2192 30500 2202 30534
rect 2202 30500 2226 30534
rect 2266 30500 2272 30534
rect 2272 30500 2300 30534
rect 2340 30500 2342 30534
rect 2342 30500 2374 30534
rect 2414 30500 2446 30534
rect 2446 30500 2448 30534
rect 2488 30500 2516 30534
rect 2516 30500 2522 30534
rect 2562 30500 2586 30534
rect 2586 30500 2596 30534
rect 2636 30500 2656 30534
rect 2656 30500 2670 30534
rect 2710 30500 2726 30534
rect 2726 30500 2744 30534
rect 2784 30500 2795 30534
rect 2795 30500 2818 30534
rect 3036 30508 3070 30538
rect 3036 30504 3070 30508
rect 386 30419 420 30447
rect 386 30413 420 30419
rect 3036 30440 3070 30466
rect 3036 30432 3070 30440
rect 386 30351 420 30375
rect 386 30341 420 30351
rect 386 30283 420 30303
rect 386 30269 420 30283
rect 386 30215 420 30231
rect 386 30197 420 30215
rect 386 30147 420 30159
rect 386 30125 420 30147
rect 386 30079 420 30087
rect 386 30053 420 30079
rect 386 30011 420 30015
rect 386 29981 420 30011
rect 386 29909 420 29943
rect 386 29841 420 29871
rect 386 29837 420 29841
rect 386 29773 420 29799
rect 386 29765 420 29773
rect 386 29705 420 29727
rect 386 29693 420 29705
rect 386 29637 420 29655
rect 386 29621 420 29637
rect 386 29569 420 29583
rect 386 29549 420 29569
rect 386 29501 420 29511
rect 386 29477 420 29501
rect 386 29433 420 29439
rect 386 29405 420 29433
rect 386 29365 420 29367
rect 386 29333 420 29365
rect 386 29263 420 29295
rect 386 29261 420 29263
rect 386 29195 420 29223
rect 386 29189 420 29195
rect 386 29127 420 29151
rect 386 29117 420 29127
rect 386 29059 420 29079
rect 386 29045 420 29059
rect 386 28991 420 29007
rect 386 28973 420 28991
rect 386 28923 420 28935
rect 386 28901 420 28923
rect 386 28855 420 28863
rect 386 28829 420 28855
rect 386 28787 420 28791
rect 386 28757 420 28787
rect 386 28685 420 28719
rect 386 28617 420 28647
rect 386 28613 420 28617
rect 386 28549 420 28575
rect 386 28541 420 28549
rect 386 28481 420 28503
rect 386 28469 420 28481
rect 531 30398 565 30432
rect 531 30325 565 30359
rect 531 30252 565 30286
rect 531 30179 565 30213
rect 531 30106 565 30140
rect 531 30033 565 30067
rect 531 29960 565 29994
rect 531 29887 565 29921
rect 531 29814 565 29848
rect 531 29741 565 29775
rect 531 29668 565 29702
rect 531 29595 565 29629
rect 531 29522 565 29556
rect 531 29448 565 29482
rect 531 29374 565 29408
rect 531 29300 565 29334
rect 531 29226 565 29260
rect 531 29152 565 29186
rect 531 29078 565 29112
rect 531 29004 565 29038
rect 531 28930 565 28964
rect 531 28856 565 28890
rect 531 28782 565 28816
rect 531 28708 565 28742
rect 531 28634 565 28668
rect 531 28560 565 28594
rect 531 28486 565 28520
rect 767 30398 801 30432
rect 767 30325 801 30359
rect 767 30252 801 30286
rect 767 30179 801 30213
rect 767 30106 801 30140
rect 767 30033 801 30067
rect 767 29960 801 29994
rect 767 29887 801 29921
rect 767 29814 801 29848
rect 767 29741 801 29775
rect 767 29668 801 29702
rect 767 29595 801 29629
rect 767 29522 801 29556
rect 767 29448 801 29482
rect 767 29374 801 29408
rect 767 29300 801 29334
rect 767 29226 801 29260
rect 767 29152 801 29186
rect 767 29078 801 29112
rect 767 29004 801 29038
rect 767 28930 801 28964
rect 767 28856 801 28890
rect 767 28782 801 28816
rect 767 28708 801 28742
rect 767 28634 801 28668
rect 767 28560 801 28594
rect 767 28486 801 28520
rect 1003 30398 1037 30432
rect 1003 30325 1037 30359
rect 1003 30252 1037 30286
rect 1003 30179 1037 30213
rect 1003 30106 1037 30140
rect 1003 30033 1037 30067
rect 1003 29960 1037 29994
rect 1003 29887 1037 29921
rect 1003 29814 1037 29848
rect 1003 29741 1037 29775
rect 1003 29668 1037 29702
rect 1003 29595 1037 29629
rect 1003 29522 1037 29556
rect 1003 29448 1037 29482
rect 1003 29374 1037 29408
rect 1003 29300 1037 29334
rect 1003 29226 1037 29260
rect 1003 29152 1037 29186
rect 1003 29078 1037 29112
rect 1003 29004 1037 29038
rect 1003 28930 1037 28964
rect 1003 28856 1037 28890
rect 1003 28782 1037 28816
rect 1003 28708 1037 28742
rect 1003 28634 1037 28668
rect 1003 28560 1037 28594
rect 1003 28486 1037 28520
rect 1239 30398 1273 30432
rect 1239 30325 1273 30359
rect 1239 30252 1273 30286
rect 1239 30179 1273 30213
rect 1239 30106 1273 30140
rect 1239 30033 1273 30067
rect 1239 29960 1273 29994
rect 1239 29887 1273 29921
rect 1239 29814 1273 29848
rect 1239 29741 1273 29775
rect 1239 29668 1273 29702
rect 1239 29595 1273 29629
rect 1239 29522 1273 29556
rect 1239 29448 1273 29482
rect 1239 29374 1273 29408
rect 1239 29300 1273 29334
rect 1239 29226 1273 29260
rect 1239 29152 1273 29186
rect 1239 29078 1273 29112
rect 1239 29004 1273 29038
rect 1239 28930 1273 28964
rect 1239 28856 1273 28890
rect 1239 28782 1273 28816
rect 1239 28708 1273 28742
rect 1239 28634 1273 28668
rect 1239 28560 1273 28594
rect 1239 28486 1273 28520
rect 1475 30398 1509 30432
rect 1475 30325 1509 30359
rect 1475 30252 1509 30286
rect 1475 30179 1509 30213
rect 1475 30106 1509 30140
rect 1475 30033 1509 30067
rect 1475 29960 1509 29994
rect 1475 29887 1509 29921
rect 1475 29814 1509 29848
rect 1475 29741 1509 29775
rect 1475 29668 1509 29702
rect 1475 29595 1509 29629
rect 1475 29522 1509 29556
rect 1475 29448 1509 29482
rect 1475 29374 1509 29408
rect 1475 29300 1509 29334
rect 1475 29226 1509 29260
rect 1475 29152 1509 29186
rect 1475 29078 1509 29112
rect 1475 29004 1509 29038
rect 1475 28930 1509 28964
rect 1475 28856 1509 28890
rect 1475 28782 1509 28816
rect 1475 28708 1509 28742
rect 1475 28634 1509 28668
rect 1475 28560 1509 28594
rect 1475 28486 1509 28520
rect 1711 30398 1745 30432
rect 1711 30325 1745 30359
rect 1711 30252 1745 30286
rect 1711 30179 1745 30213
rect 1711 30106 1745 30140
rect 1711 30033 1745 30067
rect 1711 29960 1745 29994
rect 1711 29887 1745 29921
rect 1711 29814 1745 29848
rect 1711 29741 1745 29775
rect 1711 29668 1745 29702
rect 1711 29595 1745 29629
rect 1711 29522 1745 29556
rect 1711 29448 1745 29482
rect 1711 29374 1745 29408
rect 1711 29300 1745 29334
rect 1711 29226 1745 29260
rect 1711 29152 1745 29186
rect 1711 29078 1745 29112
rect 1711 29004 1745 29038
rect 1711 28930 1745 28964
rect 1711 28856 1745 28890
rect 1711 28782 1745 28816
rect 1711 28708 1745 28742
rect 1711 28634 1745 28668
rect 1711 28560 1745 28594
rect 1711 28486 1745 28520
rect 1947 30398 1981 30432
rect 1947 30325 1981 30359
rect 1947 30252 1981 30286
rect 1947 30179 1981 30213
rect 1947 30106 1981 30140
rect 1947 30033 1981 30067
rect 1947 29960 1981 29994
rect 1947 29887 1981 29921
rect 1947 29814 1981 29848
rect 1947 29741 1981 29775
rect 1947 29668 1981 29702
rect 1947 29595 1981 29629
rect 1947 29522 1981 29556
rect 1947 29448 1981 29482
rect 1947 29374 1981 29408
rect 1947 29300 1981 29334
rect 1947 29226 1981 29260
rect 1947 29152 1981 29186
rect 1947 29078 1981 29112
rect 1947 29004 1981 29038
rect 1947 28930 1981 28964
rect 1947 28856 1981 28890
rect 1947 28782 1981 28816
rect 1947 28708 1981 28742
rect 1947 28634 1981 28668
rect 1947 28560 1981 28594
rect 1947 28486 1981 28520
rect 2183 30398 2217 30432
rect 2183 30325 2217 30359
rect 2183 30252 2217 30286
rect 2183 30179 2217 30213
rect 2183 30106 2217 30140
rect 2183 30033 2217 30067
rect 2183 29960 2217 29994
rect 2183 29887 2217 29921
rect 2183 29814 2217 29848
rect 2183 29741 2217 29775
rect 2183 29668 2217 29702
rect 2183 29595 2217 29629
rect 2183 29522 2217 29556
rect 2183 29448 2217 29482
rect 2183 29374 2217 29408
rect 2183 29300 2217 29334
rect 2183 29226 2217 29260
rect 2183 29152 2217 29186
rect 2183 29078 2217 29112
rect 2183 29004 2217 29038
rect 2183 28930 2217 28964
rect 2183 28856 2217 28890
rect 2183 28782 2217 28816
rect 2183 28708 2217 28742
rect 2183 28634 2217 28668
rect 2183 28560 2217 28594
rect 2183 28486 2217 28520
rect 2419 30398 2453 30432
rect 2419 30325 2453 30359
rect 2419 30252 2453 30286
rect 2419 30179 2453 30213
rect 2419 30106 2453 30140
rect 2419 30033 2453 30067
rect 2419 29960 2453 29994
rect 2419 29887 2453 29921
rect 2419 29814 2453 29848
rect 2419 29741 2453 29775
rect 2419 29668 2453 29702
rect 2419 29595 2453 29629
rect 2419 29522 2453 29556
rect 2419 29448 2453 29482
rect 2419 29374 2453 29408
rect 2419 29300 2453 29334
rect 2419 29226 2453 29260
rect 2419 29152 2453 29186
rect 2419 29078 2453 29112
rect 2419 29004 2453 29038
rect 2419 28930 2453 28964
rect 2419 28856 2453 28890
rect 2419 28782 2453 28816
rect 2419 28708 2453 28742
rect 2419 28634 2453 28668
rect 2419 28560 2453 28594
rect 2419 28486 2453 28520
rect 2655 30398 2689 30432
rect 2655 30325 2689 30359
rect 2655 30252 2689 30286
rect 2655 30179 2689 30213
rect 2655 30106 2689 30140
rect 2655 30033 2689 30067
rect 2655 29960 2689 29994
rect 2655 29887 2689 29921
rect 2655 29814 2689 29848
rect 2655 29741 2689 29775
rect 2655 29668 2689 29702
rect 2655 29595 2689 29629
rect 2655 29522 2689 29556
rect 2655 29448 2689 29482
rect 2655 29374 2689 29408
rect 2655 29300 2689 29334
rect 2655 29226 2689 29260
rect 2655 29152 2689 29186
rect 2655 29078 2689 29112
rect 2655 29004 2689 29038
rect 2655 28930 2689 28964
rect 2655 28856 2689 28890
rect 2655 28782 2689 28816
rect 2655 28708 2689 28742
rect 2655 28634 2689 28668
rect 2655 28560 2689 28594
rect 2655 28486 2689 28520
rect 2891 30398 2925 30432
rect 2891 30325 2925 30359
rect 2891 30252 2925 30286
rect 2891 30179 2925 30213
rect 2891 30106 2925 30140
rect 2891 30033 2925 30067
rect 2891 29960 2925 29994
rect 2891 29887 2925 29921
rect 2891 29814 2925 29848
rect 2891 29741 2925 29775
rect 2891 29668 2925 29702
rect 2891 29595 2925 29629
rect 2891 29522 2925 29556
rect 2891 29448 2925 29482
rect 2891 29374 2925 29408
rect 2891 29300 2925 29334
rect 2891 29226 2925 29260
rect 2891 29152 2925 29186
rect 2891 29078 2925 29112
rect 2891 29004 2925 29038
rect 2891 28930 2925 28964
rect 2891 28856 2925 28890
rect 2891 28782 2925 28816
rect 2891 28708 2925 28742
rect 2891 28634 2925 28668
rect 2891 28560 2925 28594
rect 2891 28486 2925 28520
rect 3036 30372 3070 30394
rect 3036 30360 3070 30372
rect 3036 30304 3070 30322
rect 3036 30288 3070 30304
rect 3036 30236 3070 30250
rect 3036 30216 3070 30236
rect 3036 30168 3070 30178
rect 3036 30144 3070 30168
rect 3036 30100 3070 30106
rect 3036 30072 3070 30100
rect 3036 30032 3070 30034
rect 3036 30000 3070 30032
rect 3036 29930 3070 29962
rect 3036 29928 3070 29930
rect 3036 29862 3070 29890
rect 3036 29856 3070 29862
rect 3036 29794 3070 29818
rect 3036 29784 3070 29794
rect 3036 29726 3070 29746
rect 3036 29712 3070 29726
rect 3036 29658 3070 29674
rect 3036 29640 3070 29658
rect 3036 29590 3070 29602
rect 3036 29568 3070 29590
rect 3036 29522 3070 29530
rect 3036 29496 3070 29522
rect 3036 29454 3070 29458
rect 3036 29424 3070 29454
rect 3036 29352 3070 29386
rect 3036 29284 3070 29314
rect 3036 29280 3070 29284
rect 3036 29216 3070 29242
rect 3036 29208 3070 29216
rect 3036 29148 3070 29170
rect 3036 29136 3070 29148
rect 3036 29080 3070 29098
rect 3036 29064 3070 29080
rect 3036 29012 3070 29026
rect 3036 28992 3070 29012
rect 3036 28944 3070 28954
rect 3036 28920 3070 28944
rect 3036 28876 3070 28882
rect 3036 28848 3070 28876
rect 3036 28808 3070 28810
rect 3036 28776 3070 28808
rect 3036 28706 3070 28738
rect 3036 28704 3070 28706
rect 3036 28638 3070 28666
rect 3036 28632 3070 28638
rect 3036 28570 3070 28594
rect 3036 28560 3070 28570
rect 386 28413 420 28431
rect 386 28397 420 28413
rect 3036 28502 3070 28522
rect 3036 28488 3070 28502
rect 386 28345 420 28359
rect 386 28325 420 28345
rect 625 28370 626 28404
rect 626 28370 659 28404
rect 700 28370 732 28404
rect 732 28370 734 28404
rect 775 28370 802 28404
rect 802 28370 809 28404
rect 850 28370 872 28404
rect 872 28370 884 28404
rect 925 28370 942 28404
rect 942 28370 959 28404
rect 1000 28370 1012 28404
rect 1012 28370 1034 28404
rect 1075 28370 1082 28404
rect 1082 28370 1109 28404
rect 1150 28370 1152 28404
rect 1152 28370 1184 28404
rect 1225 28370 1256 28404
rect 1256 28370 1259 28404
rect 1300 28370 1326 28404
rect 1326 28370 1334 28404
rect 1375 28370 1396 28404
rect 1396 28370 1409 28404
rect 1450 28370 1466 28404
rect 1466 28370 1484 28404
rect 1525 28370 1536 28404
rect 1536 28370 1559 28404
rect 1600 28370 1606 28404
rect 1606 28370 1634 28404
rect 1674 28370 1676 28404
rect 1676 28370 1708 28404
rect 1748 28370 1782 28404
rect 1822 28370 1852 28404
rect 1852 28370 1856 28404
rect 1896 28370 1922 28404
rect 1922 28370 1930 28404
rect 1970 28370 1992 28404
rect 1992 28370 2004 28404
rect 2044 28370 2062 28404
rect 2062 28370 2078 28404
rect 2118 28370 2132 28404
rect 2132 28370 2152 28404
rect 2192 28370 2202 28404
rect 2202 28370 2226 28404
rect 2266 28370 2272 28404
rect 2272 28370 2300 28404
rect 2340 28370 2342 28404
rect 2342 28370 2374 28404
rect 2414 28370 2446 28404
rect 2446 28370 2448 28404
rect 2488 28370 2516 28404
rect 2516 28370 2522 28404
rect 2562 28370 2586 28404
rect 2586 28370 2596 28404
rect 2636 28370 2656 28404
rect 2656 28370 2670 28404
rect 2710 28370 2726 28404
rect 2726 28370 2744 28404
rect 2784 28370 2795 28404
rect 2795 28370 2818 28404
rect 3036 28434 3070 28450
rect 3036 28416 3070 28434
rect 386 28277 420 28287
rect 386 28253 420 28277
rect 3036 28366 3070 28378
rect 3036 28344 3070 28366
rect 386 28209 420 28215
rect 386 28181 420 28209
rect 386 28141 420 28143
rect 386 28109 420 28141
rect 386 28039 420 28071
rect 386 28037 420 28039
rect 386 27971 420 27999
rect 386 27965 420 27971
rect 386 27903 420 27927
rect 386 27893 420 27903
rect 386 27835 420 27855
rect 386 27821 420 27835
rect 386 27767 420 27783
rect 386 27749 420 27767
rect 386 27699 420 27711
rect 386 27677 420 27699
rect 386 27631 420 27639
rect 386 27605 420 27631
rect 386 27563 420 27567
rect 386 27533 420 27563
rect 386 27461 420 27495
rect 386 27393 420 27423
rect 386 27389 420 27393
rect 386 27325 420 27351
rect 386 27317 420 27325
rect 386 27257 420 27279
rect 386 27245 420 27257
rect 386 27189 420 27207
rect 386 27173 420 27189
rect 386 27121 420 27135
rect 386 27101 420 27121
rect 386 27053 420 27063
rect 386 27029 420 27053
rect 386 26985 420 26991
rect 386 26957 420 26985
rect 386 26917 420 26919
rect 386 26885 420 26917
rect 386 26815 420 26847
rect 386 26813 420 26815
rect 386 26747 420 26775
rect 386 26741 420 26747
rect 386 26679 420 26703
rect 386 26669 420 26679
rect 386 26611 420 26631
rect 386 26597 420 26611
rect 386 26543 420 26559
rect 386 26525 420 26543
rect 386 26475 420 26487
rect 386 26453 420 26475
rect 386 26407 420 26415
rect 386 26381 420 26407
rect 386 26339 420 26343
rect 386 26309 420 26339
rect 531 28254 565 28288
rect 531 28181 565 28215
rect 531 28108 565 28142
rect 531 28035 565 28069
rect 531 27962 565 27996
rect 531 27889 565 27923
rect 531 27816 565 27850
rect 531 27743 565 27777
rect 531 27670 565 27704
rect 531 27597 565 27631
rect 531 27524 565 27558
rect 531 27451 565 27485
rect 531 27378 565 27412
rect 531 27304 565 27338
rect 531 27230 565 27264
rect 531 27156 565 27190
rect 531 27082 565 27116
rect 531 27008 565 27042
rect 531 26934 565 26968
rect 531 26860 565 26894
rect 531 26786 565 26820
rect 531 26712 565 26746
rect 531 26638 565 26672
rect 531 26564 565 26598
rect 531 26490 565 26524
rect 531 26416 565 26450
rect 531 26342 565 26376
rect 767 28254 801 28288
rect 767 28181 801 28215
rect 767 28108 801 28142
rect 767 28035 801 28069
rect 767 27962 801 27996
rect 767 27889 801 27923
rect 767 27816 801 27850
rect 767 27743 801 27777
rect 767 27670 801 27704
rect 767 27597 801 27631
rect 767 27524 801 27558
rect 767 27451 801 27485
rect 767 27378 801 27412
rect 767 27304 801 27338
rect 767 27230 801 27264
rect 767 27156 801 27190
rect 767 27082 801 27116
rect 767 27008 801 27042
rect 767 26934 801 26968
rect 767 26860 801 26894
rect 767 26786 801 26820
rect 767 26712 801 26746
rect 767 26638 801 26672
rect 767 26564 801 26598
rect 767 26490 801 26524
rect 767 26416 801 26450
rect 767 26342 801 26376
rect 1003 28254 1037 28288
rect 1003 28181 1037 28215
rect 1003 28108 1037 28142
rect 1003 28035 1037 28069
rect 1003 27962 1037 27996
rect 1003 27889 1037 27923
rect 1003 27816 1037 27850
rect 1003 27743 1037 27777
rect 1003 27670 1037 27704
rect 1003 27597 1037 27631
rect 1003 27524 1037 27558
rect 1003 27451 1037 27485
rect 1003 27378 1037 27412
rect 1003 27304 1037 27338
rect 1003 27230 1037 27264
rect 1003 27156 1037 27190
rect 1003 27082 1037 27116
rect 1003 27008 1037 27042
rect 1003 26934 1037 26968
rect 1003 26860 1037 26894
rect 1003 26786 1037 26820
rect 1003 26712 1037 26746
rect 1003 26638 1037 26672
rect 1003 26564 1037 26598
rect 1003 26490 1037 26524
rect 1003 26416 1037 26450
rect 1003 26342 1037 26376
rect 1239 28254 1273 28288
rect 1239 28181 1273 28215
rect 1239 28108 1273 28142
rect 1239 28035 1273 28069
rect 1239 27962 1273 27996
rect 1239 27889 1273 27923
rect 1239 27816 1273 27850
rect 1239 27743 1273 27777
rect 1239 27670 1273 27704
rect 1239 27597 1273 27631
rect 1239 27524 1273 27558
rect 1239 27451 1273 27485
rect 1239 27378 1273 27412
rect 1239 27304 1273 27338
rect 1239 27230 1273 27264
rect 1239 27156 1273 27190
rect 1239 27082 1273 27116
rect 1239 27008 1273 27042
rect 1239 26934 1273 26968
rect 1239 26860 1273 26894
rect 1239 26786 1273 26820
rect 1239 26712 1273 26746
rect 1239 26638 1273 26672
rect 1239 26564 1273 26598
rect 1239 26490 1273 26524
rect 1239 26416 1273 26450
rect 1239 26342 1273 26376
rect 1475 28254 1509 28288
rect 1475 28181 1509 28215
rect 1475 28108 1509 28142
rect 1475 28035 1509 28069
rect 1475 27962 1509 27996
rect 1475 27889 1509 27923
rect 1475 27816 1509 27850
rect 1475 27743 1509 27777
rect 1475 27670 1509 27704
rect 1475 27597 1509 27631
rect 1475 27524 1509 27558
rect 1475 27451 1509 27485
rect 1475 27378 1509 27412
rect 1475 27304 1509 27338
rect 1475 27230 1509 27264
rect 1475 27156 1509 27190
rect 1475 27082 1509 27116
rect 1475 27008 1509 27042
rect 1475 26934 1509 26968
rect 1475 26860 1509 26894
rect 1475 26786 1509 26820
rect 1475 26712 1509 26746
rect 1475 26638 1509 26672
rect 1475 26564 1509 26598
rect 1475 26490 1509 26524
rect 1475 26416 1509 26450
rect 1475 26342 1509 26376
rect 1711 28254 1745 28288
rect 1711 28181 1745 28215
rect 1711 28108 1745 28142
rect 1711 28035 1745 28069
rect 1711 27962 1745 27996
rect 1711 27889 1745 27923
rect 1711 27816 1745 27850
rect 1711 27743 1745 27777
rect 1711 27670 1745 27704
rect 1711 27597 1745 27631
rect 1711 27524 1745 27558
rect 1711 27451 1745 27485
rect 1711 27378 1745 27412
rect 1711 27304 1745 27338
rect 1711 27230 1745 27264
rect 1711 27156 1745 27190
rect 1711 27082 1745 27116
rect 1711 27008 1745 27042
rect 1711 26934 1745 26968
rect 1711 26860 1745 26894
rect 1711 26786 1745 26820
rect 1711 26712 1745 26746
rect 1711 26638 1745 26672
rect 1711 26564 1745 26598
rect 1711 26490 1745 26524
rect 1711 26416 1745 26450
rect 1711 26342 1745 26376
rect 1947 28254 1981 28288
rect 1947 28181 1981 28215
rect 1947 28108 1981 28142
rect 1947 28035 1981 28069
rect 1947 27962 1981 27996
rect 1947 27889 1981 27923
rect 1947 27816 1981 27850
rect 1947 27743 1981 27777
rect 1947 27670 1981 27704
rect 1947 27597 1981 27631
rect 1947 27524 1981 27558
rect 1947 27451 1981 27485
rect 1947 27378 1981 27412
rect 1947 27304 1981 27338
rect 1947 27230 1981 27264
rect 1947 27156 1981 27190
rect 1947 27082 1981 27116
rect 1947 27008 1981 27042
rect 1947 26934 1981 26968
rect 1947 26860 1981 26894
rect 1947 26786 1981 26820
rect 1947 26712 1981 26746
rect 1947 26638 1981 26672
rect 1947 26564 1981 26598
rect 1947 26490 1981 26524
rect 1947 26416 1981 26450
rect 1947 26342 1981 26376
rect 2183 28254 2217 28288
rect 2183 28181 2217 28215
rect 2183 28108 2217 28142
rect 2183 28035 2217 28069
rect 2183 27962 2217 27996
rect 2183 27889 2217 27923
rect 2183 27816 2217 27850
rect 2183 27743 2217 27777
rect 2183 27670 2217 27704
rect 2183 27597 2217 27631
rect 2183 27524 2217 27558
rect 2183 27451 2217 27485
rect 2183 27378 2217 27412
rect 2183 27304 2217 27338
rect 2183 27230 2217 27264
rect 2183 27156 2217 27190
rect 2183 27082 2217 27116
rect 2183 27008 2217 27042
rect 2183 26934 2217 26968
rect 2183 26860 2217 26894
rect 2183 26786 2217 26820
rect 2183 26712 2217 26746
rect 2183 26638 2217 26672
rect 2183 26564 2217 26598
rect 2183 26490 2217 26524
rect 2183 26416 2217 26450
rect 2183 26342 2217 26376
rect 2419 28254 2453 28288
rect 2419 28181 2453 28215
rect 2419 28108 2453 28142
rect 2419 28035 2453 28069
rect 2419 27962 2453 27996
rect 2419 27889 2453 27923
rect 2419 27816 2453 27850
rect 2419 27743 2453 27777
rect 2419 27670 2453 27704
rect 2419 27597 2453 27631
rect 2419 27524 2453 27558
rect 2419 27451 2453 27485
rect 2419 27378 2453 27412
rect 2419 27304 2453 27338
rect 2419 27230 2453 27264
rect 2419 27156 2453 27190
rect 2419 27082 2453 27116
rect 2419 27008 2453 27042
rect 2419 26934 2453 26968
rect 2419 26860 2453 26894
rect 2419 26786 2453 26820
rect 2419 26712 2453 26746
rect 2419 26638 2453 26672
rect 2419 26564 2453 26598
rect 2419 26490 2453 26524
rect 2419 26416 2453 26450
rect 2419 26342 2453 26376
rect 2655 28254 2689 28288
rect 2655 28181 2689 28215
rect 2655 28108 2689 28142
rect 2655 28035 2689 28069
rect 2655 27962 2689 27996
rect 2655 27889 2689 27923
rect 2655 27816 2689 27850
rect 2655 27743 2689 27777
rect 2655 27670 2689 27704
rect 2655 27597 2689 27631
rect 2655 27524 2689 27558
rect 2655 27451 2689 27485
rect 2655 27378 2689 27412
rect 2655 27304 2689 27338
rect 2655 27230 2689 27264
rect 2655 27156 2689 27190
rect 2655 27082 2689 27116
rect 2655 27008 2689 27042
rect 2655 26934 2689 26968
rect 2655 26860 2689 26894
rect 2655 26786 2689 26820
rect 2655 26712 2689 26746
rect 2655 26638 2689 26672
rect 2655 26564 2689 26598
rect 2655 26490 2689 26524
rect 2655 26416 2689 26450
rect 2655 26342 2689 26376
rect 2891 28254 2925 28288
rect 2891 28181 2925 28215
rect 2891 28108 2925 28142
rect 2891 28035 2925 28069
rect 2891 27962 2925 27996
rect 2891 27889 2925 27923
rect 2891 27816 2925 27850
rect 2891 27743 2925 27777
rect 2891 27670 2925 27704
rect 2891 27597 2925 27631
rect 2891 27524 2925 27558
rect 2891 27451 2925 27485
rect 2891 27378 2925 27412
rect 2891 27304 2925 27338
rect 2891 27230 2925 27264
rect 2891 27156 2925 27190
rect 2891 27082 2925 27116
rect 2891 27008 2925 27042
rect 2891 26934 2925 26968
rect 2891 26860 2925 26894
rect 2891 26786 2925 26820
rect 2891 26712 2925 26746
rect 2891 26638 2925 26672
rect 2891 26564 2925 26598
rect 2891 26490 2925 26524
rect 2891 26416 2925 26450
rect 2891 26342 2925 26376
rect 3036 28298 3070 28306
rect 3036 28272 3070 28298
rect 3036 28230 3070 28234
rect 3036 28200 3070 28230
rect 3036 28128 3070 28162
rect 3036 28060 3070 28090
rect 3036 28056 3070 28060
rect 3036 27992 3070 28018
rect 3036 27984 3070 27992
rect 3036 27924 3070 27946
rect 3036 27912 3070 27924
rect 3036 27856 3070 27874
rect 3036 27840 3070 27856
rect 3036 27788 3070 27802
rect 3036 27768 3070 27788
rect 3036 27720 3070 27730
rect 3036 27696 3070 27720
rect 3036 27652 3070 27658
rect 3036 27624 3070 27652
rect 3036 27584 3070 27586
rect 3036 27552 3070 27584
rect 3036 27482 3070 27514
rect 3036 27480 3070 27482
rect 3036 27414 3070 27442
rect 3036 27408 3070 27414
rect 3036 27346 3070 27370
rect 3036 27336 3070 27346
rect 3036 27278 3070 27298
rect 3036 27264 3070 27278
rect 3036 27210 3070 27226
rect 3036 27192 3070 27210
rect 3036 27142 3070 27154
rect 3036 27120 3070 27142
rect 3036 27074 3070 27082
rect 3036 27048 3070 27074
rect 3036 27006 3070 27010
rect 3036 26976 3070 27006
rect 3036 26904 3070 26938
rect 3036 26836 3070 26866
rect 3036 26832 3070 26836
rect 3036 26768 3070 26794
rect 3036 26760 3070 26768
rect 3036 26700 3070 26722
rect 3036 26688 3070 26700
rect 3036 26632 3070 26650
rect 3036 26616 3070 26632
rect 3036 26564 3070 26578
rect 3036 26544 3070 26564
rect 3036 26496 3070 26506
rect 3036 26472 3070 26496
rect 3036 26428 3070 26434
rect 3036 26400 3070 26428
rect 3036 26360 3070 26362
rect 3036 26328 3070 26360
rect 386 26237 420 26271
rect 625 26240 626 26274
rect 626 26240 659 26274
rect 700 26240 732 26274
rect 732 26240 734 26274
rect 775 26240 802 26274
rect 802 26240 809 26274
rect 850 26240 872 26274
rect 872 26240 884 26274
rect 925 26240 942 26274
rect 942 26240 959 26274
rect 1000 26240 1012 26274
rect 1012 26240 1034 26274
rect 1075 26240 1082 26274
rect 1082 26240 1109 26274
rect 1150 26240 1152 26274
rect 1152 26240 1184 26274
rect 1225 26240 1256 26274
rect 1256 26240 1259 26274
rect 1300 26240 1326 26274
rect 1326 26240 1334 26274
rect 1375 26240 1396 26274
rect 1396 26240 1409 26274
rect 1450 26240 1466 26274
rect 1466 26240 1484 26274
rect 1525 26240 1536 26274
rect 1536 26240 1559 26274
rect 1600 26240 1606 26274
rect 1606 26240 1634 26274
rect 1674 26240 1676 26274
rect 1676 26240 1708 26274
rect 1748 26240 1782 26274
rect 1822 26240 1852 26274
rect 1852 26240 1856 26274
rect 1896 26240 1922 26274
rect 1922 26240 1930 26274
rect 1970 26240 1992 26274
rect 1992 26240 2004 26274
rect 2044 26240 2062 26274
rect 2062 26240 2078 26274
rect 2118 26240 2132 26274
rect 2132 26240 2152 26274
rect 2192 26240 2202 26274
rect 2202 26240 2226 26274
rect 2266 26240 2272 26274
rect 2272 26240 2300 26274
rect 2340 26240 2342 26274
rect 2342 26240 2374 26274
rect 2414 26240 2446 26274
rect 2446 26240 2448 26274
rect 2488 26240 2516 26274
rect 2516 26240 2522 26274
rect 2562 26240 2586 26274
rect 2586 26240 2596 26274
rect 2636 26240 2656 26274
rect 2656 26240 2670 26274
rect 2710 26240 2726 26274
rect 2726 26240 2744 26274
rect 2784 26240 2795 26274
rect 2795 26240 2818 26274
rect 386 26169 420 26199
rect 386 26165 420 26169
rect 3036 26258 3070 26290
rect 3036 26256 3070 26258
rect 386 26101 420 26127
rect 386 26093 420 26101
rect 386 26033 420 26055
rect 386 26021 420 26033
rect 386 25965 420 25983
rect 386 25949 420 25965
rect 386 25897 420 25911
rect 386 25877 420 25897
rect 386 25829 420 25839
rect 386 25805 420 25829
rect 386 25761 420 25767
rect 386 25733 420 25761
rect 386 25693 420 25695
rect 386 25661 420 25693
rect 386 25591 420 25623
rect 386 25589 420 25591
rect 386 25523 420 25551
rect 386 25517 420 25523
rect 386 25455 420 25479
rect 386 25445 420 25455
rect 386 25387 420 25407
rect 386 25373 420 25387
rect 386 25319 420 25335
rect 386 25301 420 25319
rect 386 25251 420 25263
rect 386 25229 420 25251
rect 386 25183 420 25191
rect 386 25157 420 25183
rect 386 25115 420 25119
rect 386 25085 420 25115
rect 386 25013 420 25047
rect 386 24945 420 24975
rect 386 24941 420 24945
rect 386 24877 420 24903
rect 386 24869 420 24877
rect 386 24809 420 24831
rect 386 24797 420 24809
rect 386 24741 420 24759
rect 386 24725 420 24741
rect 386 24673 420 24687
rect 386 24653 420 24673
rect 386 24605 420 24615
rect 386 24581 420 24605
rect 386 24537 420 24543
rect 386 24509 420 24537
rect 386 24469 420 24471
rect 386 24437 420 24469
rect 386 24367 420 24399
rect 386 24365 420 24367
rect 386 24299 420 24327
rect 386 24293 420 24299
rect 386 24231 420 24255
rect 386 24221 420 24231
rect 531 26138 565 26172
rect 531 26065 565 26099
rect 531 25992 565 26026
rect 531 25919 565 25953
rect 531 25846 565 25880
rect 531 25773 565 25807
rect 531 25700 565 25734
rect 531 25627 565 25661
rect 531 25554 565 25588
rect 531 25481 565 25515
rect 531 25408 565 25442
rect 531 25335 565 25369
rect 531 25262 565 25296
rect 531 25188 565 25222
rect 531 25114 565 25148
rect 531 25040 565 25074
rect 531 24966 565 25000
rect 531 24892 565 24926
rect 531 24818 565 24852
rect 531 24744 565 24778
rect 531 24670 565 24704
rect 531 24596 565 24630
rect 531 24522 565 24556
rect 531 24448 565 24482
rect 531 24374 565 24408
rect 531 24300 565 24334
rect 531 24226 565 24260
rect 767 26138 801 26172
rect 767 26065 801 26099
rect 767 25992 801 26026
rect 767 25919 801 25953
rect 767 25846 801 25880
rect 767 25773 801 25807
rect 767 25700 801 25734
rect 767 25627 801 25661
rect 767 25554 801 25588
rect 767 25481 801 25515
rect 767 25408 801 25442
rect 767 25335 801 25369
rect 767 25262 801 25296
rect 767 25188 801 25222
rect 767 25114 801 25148
rect 767 25040 801 25074
rect 767 24966 801 25000
rect 767 24892 801 24926
rect 767 24818 801 24852
rect 767 24744 801 24778
rect 767 24670 801 24704
rect 767 24596 801 24630
rect 767 24522 801 24556
rect 767 24448 801 24482
rect 767 24374 801 24408
rect 767 24300 801 24334
rect 767 24226 801 24260
rect 1003 26138 1037 26172
rect 1003 26065 1037 26099
rect 1003 25992 1037 26026
rect 1003 25919 1037 25953
rect 1003 25846 1037 25880
rect 1003 25773 1037 25807
rect 1003 25700 1037 25734
rect 1003 25627 1037 25661
rect 1003 25554 1037 25588
rect 1003 25481 1037 25515
rect 1003 25408 1037 25442
rect 1003 25335 1037 25369
rect 1003 25262 1037 25296
rect 1003 25188 1037 25222
rect 1003 25114 1037 25148
rect 1003 25040 1037 25074
rect 1003 24966 1037 25000
rect 1003 24892 1037 24926
rect 1003 24818 1037 24852
rect 1003 24744 1037 24778
rect 1003 24670 1037 24704
rect 1003 24596 1037 24630
rect 1003 24522 1037 24556
rect 1003 24448 1037 24482
rect 1003 24374 1037 24408
rect 1003 24300 1037 24334
rect 1003 24226 1037 24260
rect 1239 26138 1273 26172
rect 1239 26065 1273 26099
rect 1239 25992 1273 26026
rect 1239 25919 1273 25953
rect 1239 25846 1273 25880
rect 1239 25773 1273 25807
rect 1239 25700 1273 25734
rect 1239 25627 1273 25661
rect 1239 25554 1273 25588
rect 1239 25481 1273 25515
rect 1239 25408 1273 25442
rect 1239 25335 1273 25369
rect 1239 25262 1273 25296
rect 1239 25188 1273 25222
rect 1239 25114 1273 25148
rect 1239 25040 1273 25074
rect 1239 24966 1273 25000
rect 1239 24892 1273 24926
rect 1239 24818 1273 24852
rect 1239 24744 1273 24778
rect 1239 24670 1273 24704
rect 1239 24596 1273 24630
rect 1239 24522 1273 24556
rect 1239 24448 1273 24482
rect 1239 24374 1273 24408
rect 1239 24300 1273 24334
rect 1239 24226 1273 24260
rect 1475 26138 1509 26172
rect 1475 26065 1509 26099
rect 1475 25992 1509 26026
rect 1475 25919 1509 25953
rect 1475 25846 1509 25880
rect 1475 25773 1509 25807
rect 1475 25700 1509 25734
rect 1475 25627 1509 25661
rect 1475 25554 1509 25588
rect 1475 25481 1509 25515
rect 1475 25408 1509 25442
rect 1475 25335 1509 25369
rect 1475 25262 1509 25296
rect 1475 25188 1509 25222
rect 1475 25114 1509 25148
rect 1475 25040 1509 25074
rect 1475 24966 1509 25000
rect 1475 24892 1509 24926
rect 1475 24818 1509 24852
rect 1475 24744 1509 24778
rect 1475 24670 1509 24704
rect 1475 24596 1509 24630
rect 1475 24522 1509 24556
rect 1475 24448 1509 24482
rect 1475 24374 1509 24408
rect 1475 24300 1509 24334
rect 1475 24226 1509 24260
rect 1711 26138 1745 26172
rect 1711 26065 1745 26099
rect 1711 25992 1745 26026
rect 1711 25919 1745 25953
rect 1711 25846 1745 25880
rect 1711 25773 1745 25807
rect 1711 25700 1745 25734
rect 1711 25627 1745 25661
rect 1711 25554 1745 25588
rect 1711 25481 1745 25515
rect 1711 25408 1745 25442
rect 1711 25335 1745 25369
rect 1711 25262 1745 25296
rect 1711 25188 1745 25222
rect 1711 25114 1745 25148
rect 1711 25040 1745 25074
rect 1711 24966 1745 25000
rect 1711 24892 1745 24926
rect 1711 24818 1745 24852
rect 1711 24744 1745 24778
rect 1711 24670 1745 24704
rect 1711 24596 1745 24630
rect 1711 24522 1745 24556
rect 1711 24448 1745 24482
rect 1711 24374 1745 24408
rect 1711 24300 1745 24334
rect 1711 24226 1745 24260
rect 1947 26138 1981 26172
rect 1947 26065 1981 26099
rect 1947 25992 1981 26026
rect 1947 25919 1981 25953
rect 1947 25846 1981 25880
rect 1947 25773 1981 25807
rect 1947 25700 1981 25734
rect 1947 25627 1981 25661
rect 1947 25554 1981 25588
rect 1947 25481 1981 25515
rect 1947 25408 1981 25442
rect 1947 25335 1981 25369
rect 1947 25262 1981 25296
rect 1947 25188 1981 25222
rect 1947 25114 1981 25148
rect 1947 25040 1981 25074
rect 1947 24966 1981 25000
rect 1947 24892 1981 24926
rect 1947 24818 1981 24852
rect 1947 24744 1981 24778
rect 1947 24670 1981 24704
rect 1947 24596 1981 24630
rect 1947 24522 1981 24556
rect 1947 24448 1981 24482
rect 1947 24374 1981 24408
rect 1947 24300 1981 24334
rect 1947 24226 1981 24260
rect 2183 26138 2217 26172
rect 2183 26065 2217 26099
rect 2183 25992 2217 26026
rect 2183 25919 2217 25953
rect 2183 25846 2217 25880
rect 2183 25773 2217 25807
rect 2183 25700 2217 25734
rect 2183 25627 2217 25661
rect 2183 25554 2217 25588
rect 2183 25481 2217 25515
rect 2183 25408 2217 25442
rect 2183 25335 2217 25369
rect 2183 25262 2217 25296
rect 2183 25188 2217 25222
rect 2183 25114 2217 25148
rect 2183 25040 2217 25074
rect 2183 24966 2217 25000
rect 2183 24892 2217 24926
rect 2183 24818 2217 24852
rect 2183 24744 2217 24778
rect 2183 24670 2217 24704
rect 2183 24596 2217 24630
rect 2183 24522 2217 24556
rect 2183 24448 2217 24482
rect 2183 24374 2217 24408
rect 2183 24300 2217 24334
rect 2183 24226 2217 24260
rect 2419 26138 2453 26172
rect 2419 26065 2453 26099
rect 2419 25992 2453 26026
rect 2419 25919 2453 25953
rect 2419 25846 2453 25880
rect 2419 25773 2453 25807
rect 2419 25700 2453 25734
rect 2419 25627 2453 25661
rect 2419 25554 2453 25588
rect 2419 25481 2453 25515
rect 2419 25408 2453 25442
rect 2419 25335 2453 25369
rect 2419 25262 2453 25296
rect 2419 25188 2453 25222
rect 2419 25114 2453 25148
rect 2419 25040 2453 25074
rect 2419 24966 2453 25000
rect 2419 24892 2453 24926
rect 2419 24818 2453 24852
rect 2419 24744 2453 24778
rect 2419 24670 2453 24704
rect 2419 24596 2453 24630
rect 2419 24522 2453 24556
rect 2419 24448 2453 24482
rect 2419 24374 2453 24408
rect 2419 24300 2453 24334
rect 2419 24226 2453 24260
rect 2655 26138 2689 26172
rect 2655 26065 2689 26099
rect 2655 25992 2689 26026
rect 2655 25919 2689 25953
rect 2655 25846 2689 25880
rect 2655 25773 2689 25807
rect 2655 25700 2689 25734
rect 2655 25627 2689 25661
rect 2655 25554 2689 25588
rect 2655 25481 2689 25515
rect 2655 25408 2689 25442
rect 2655 25335 2689 25369
rect 2655 25262 2689 25296
rect 2655 25188 2689 25222
rect 2655 25114 2689 25148
rect 2655 25040 2689 25074
rect 2655 24966 2689 25000
rect 2655 24892 2689 24926
rect 2655 24818 2689 24852
rect 2655 24744 2689 24778
rect 2655 24670 2689 24704
rect 2655 24596 2689 24630
rect 2655 24522 2689 24556
rect 2655 24448 2689 24482
rect 2655 24374 2689 24408
rect 2655 24300 2689 24334
rect 2655 24226 2689 24260
rect 2891 26138 2925 26172
rect 2891 26065 2925 26099
rect 2891 25992 2925 26026
rect 2891 25919 2925 25953
rect 2891 25846 2925 25880
rect 2891 25773 2925 25807
rect 2891 25700 2925 25734
rect 2891 25627 2925 25661
rect 2891 25554 2925 25588
rect 2891 25481 2925 25515
rect 2891 25408 2925 25442
rect 2891 25335 2925 25369
rect 2891 25262 2925 25296
rect 2891 25188 2925 25222
rect 2891 25114 2925 25148
rect 2891 25040 2925 25074
rect 2891 24966 2925 25000
rect 2891 24892 2925 24926
rect 2891 24818 2925 24852
rect 2891 24744 2925 24778
rect 2891 24670 2925 24704
rect 2891 24596 2925 24630
rect 2891 24522 2925 24556
rect 2891 24448 2925 24482
rect 2891 24374 2925 24408
rect 2891 24300 2925 24334
rect 2891 24226 2925 24260
rect 3036 26190 3070 26218
rect 3036 26184 3070 26190
rect 3036 26122 3070 26146
rect 3036 26112 3070 26122
rect 3036 26054 3070 26074
rect 3036 26040 3070 26054
rect 3036 25986 3070 26002
rect 3036 25968 3070 25986
rect 3036 25918 3070 25930
rect 3036 25896 3070 25918
rect 3036 25850 3070 25858
rect 3036 25824 3070 25850
rect 3036 25782 3070 25786
rect 3036 25752 3070 25782
rect 3036 25680 3070 25714
rect 3036 25612 3070 25642
rect 3036 25608 3070 25612
rect 3036 25544 3070 25570
rect 3036 25536 3070 25544
rect 3036 25476 3070 25498
rect 3036 25464 3070 25476
rect 3036 25408 3070 25426
rect 3036 25392 3070 25408
rect 3036 25340 3070 25354
rect 3036 25320 3070 25340
rect 3036 25272 3070 25282
rect 3036 25248 3070 25272
rect 3036 25204 3070 25210
rect 3036 25176 3070 25204
rect 3036 25136 3070 25138
rect 3036 25104 3070 25136
rect 3036 25034 3070 25066
rect 3036 25032 3070 25034
rect 3036 24966 3070 24994
rect 3036 24960 3070 24966
rect 3036 24898 3070 24922
rect 3036 24888 3070 24898
rect 3036 24830 3070 24850
rect 3036 24816 3070 24830
rect 3036 24762 3070 24778
rect 3036 24744 3070 24762
rect 3036 24694 3070 24706
rect 3036 24672 3070 24694
rect 3036 24626 3070 24634
rect 3036 24600 3070 24626
rect 3036 24558 3070 24562
rect 3036 24528 3070 24558
rect 3036 24456 3070 24490
rect 3036 24388 3070 24418
rect 3036 24384 3070 24388
rect 3036 24320 3070 24346
rect 3036 24312 3070 24320
rect 3036 24252 3070 24274
rect 3036 24240 3070 24252
rect 386 24163 420 24183
rect 386 24149 420 24163
rect 3036 24184 3070 24202
rect 3036 24168 3070 24184
rect 386 24095 420 24111
rect 386 24077 420 24095
rect 625 24110 626 24144
rect 626 24110 659 24144
rect 700 24110 732 24144
rect 732 24110 734 24144
rect 775 24110 802 24144
rect 802 24110 809 24144
rect 850 24110 872 24144
rect 872 24110 884 24144
rect 925 24110 942 24144
rect 942 24110 959 24144
rect 1000 24110 1012 24144
rect 1012 24110 1034 24144
rect 1075 24110 1082 24144
rect 1082 24110 1109 24144
rect 1150 24110 1152 24144
rect 1152 24110 1184 24144
rect 1225 24110 1256 24144
rect 1256 24110 1259 24144
rect 1300 24110 1326 24144
rect 1326 24110 1334 24144
rect 1375 24110 1396 24144
rect 1396 24110 1409 24144
rect 1450 24110 1466 24144
rect 1466 24110 1484 24144
rect 1525 24110 1536 24144
rect 1536 24110 1559 24144
rect 1600 24110 1606 24144
rect 1606 24110 1634 24144
rect 1674 24110 1676 24144
rect 1676 24110 1708 24144
rect 1748 24110 1782 24144
rect 1822 24110 1852 24144
rect 1852 24110 1856 24144
rect 1896 24110 1922 24144
rect 1922 24110 1930 24144
rect 1970 24110 1992 24144
rect 1992 24110 2004 24144
rect 2044 24110 2062 24144
rect 2062 24110 2078 24144
rect 2118 24110 2132 24144
rect 2132 24110 2152 24144
rect 2192 24110 2202 24144
rect 2202 24110 2226 24144
rect 2266 24110 2272 24144
rect 2272 24110 2300 24144
rect 2340 24110 2342 24144
rect 2342 24110 2374 24144
rect 2414 24110 2446 24144
rect 2446 24110 2448 24144
rect 2488 24110 2516 24144
rect 2516 24110 2522 24144
rect 2562 24110 2586 24144
rect 2586 24110 2596 24144
rect 2636 24110 2656 24144
rect 2656 24110 2670 24144
rect 2710 24110 2726 24144
rect 2726 24110 2744 24144
rect 2784 24110 2795 24144
rect 2795 24110 2818 24144
rect 386 24027 420 24039
rect 386 24005 420 24027
rect 3036 24116 3070 24130
rect 3036 24096 3070 24116
rect 386 23959 420 23967
rect 386 23933 420 23959
rect 386 23891 420 23895
rect 386 23861 420 23891
rect 386 23789 420 23823
rect 386 23721 420 23751
rect 386 23717 420 23721
rect 386 23653 420 23679
rect 386 23645 420 23653
rect 386 23585 420 23607
rect 386 23573 420 23585
rect 386 23517 420 23535
rect 386 23501 420 23517
rect 386 23449 420 23463
rect 386 23429 420 23449
rect 386 23381 420 23391
rect 386 23357 420 23381
rect 386 23313 420 23319
rect 386 23285 420 23313
rect 386 23245 420 23247
rect 386 23213 420 23245
rect 386 23143 420 23175
rect 386 23141 420 23143
rect 386 23075 420 23103
rect 386 23069 420 23075
rect 386 23007 420 23031
rect 386 22997 420 23007
rect 386 22939 420 22959
rect 386 22925 420 22939
rect 386 22871 420 22887
rect 386 22853 420 22871
rect 386 22803 420 22815
rect 386 22781 420 22803
rect 386 22735 420 22743
rect 386 22709 420 22735
rect 386 22667 420 22671
rect 386 22637 420 22667
rect 386 22565 420 22599
rect 386 22497 420 22527
rect 386 22493 420 22497
rect 386 22429 420 22455
rect 386 22421 420 22429
rect 386 22361 420 22383
rect 386 22349 420 22361
rect 386 22293 420 22311
rect 386 22277 420 22293
rect 386 22225 420 22239
rect 386 22205 420 22225
rect 386 22157 420 22167
rect 386 22133 420 22157
rect 386 22089 420 22095
rect 386 22061 420 22089
rect 531 23994 565 24028
rect 531 23921 565 23955
rect 531 23848 565 23882
rect 531 23775 565 23809
rect 531 23702 565 23736
rect 531 23629 565 23663
rect 531 23556 565 23590
rect 531 23483 565 23517
rect 531 23410 565 23444
rect 531 23337 565 23371
rect 531 23264 565 23298
rect 531 23191 565 23225
rect 531 23118 565 23152
rect 531 23044 565 23078
rect 531 22970 565 23004
rect 531 22896 565 22930
rect 531 22822 565 22856
rect 531 22748 565 22782
rect 531 22674 565 22708
rect 531 22600 565 22634
rect 531 22526 565 22560
rect 531 22452 565 22486
rect 531 22378 565 22412
rect 531 22304 565 22338
rect 531 22230 565 22264
rect 531 22156 565 22190
rect 531 22082 565 22116
rect 767 23994 801 24028
rect 767 23921 801 23955
rect 767 23848 801 23882
rect 767 23775 801 23809
rect 767 23702 801 23736
rect 767 23629 801 23663
rect 767 23556 801 23590
rect 767 23483 801 23517
rect 767 23410 801 23444
rect 767 23337 801 23371
rect 767 23264 801 23298
rect 767 23191 801 23225
rect 767 23118 801 23152
rect 767 23044 801 23078
rect 767 22970 801 23004
rect 767 22896 801 22930
rect 767 22822 801 22856
rect 767 22748 801 22782
rect 767 22674 801 22708
rect 767 22600 801 22634
rect 767 22526 801 22560
rect 767 22452 801 22486
rect 767 22378 801 22412
rect 767 22304 801 22338
rect 767 22230 801 22264
rect 767 22156 801 22190
rect 767 22082 801 22116
rect 1003 23994 1037 24028
rect 1003 23921 1037 23955
rect 1003 23848 1037 23882
rect 1003 23775 1037 23809
rect 1003 23702 1037 23736
rect 1003 23629 1037 23663
rect 1003 23556 1037 23590
rect 1003 23483 1037 23517
rect 1003 23410 1037 23444
rect 1003 23337 1037 23371
rect 1003 23264 1037 23298
rect 1003 23191 1037 23225
rect 1003 23118 1037 23152
rect 1003 23044 1037 23078
rect 1003 22970 1037 23004
rect 1003 22896 1037 22930
rect 1003 22822 1037 22856
rect 1003 22748 1037 22782
rect 1003 22674 1037 22708
rect 1003 22600 1037 22634
rect 1003 22526 1037 22560
rect 1003 22452 1037 22486
rect 1003 22378 1037 22412
rect 1003 22304 1037 22338
rect 1003 22230 1037 22264
rect 1003 22156 1037 22190
rect 1003 22082 1037 22116
rect 1239 23994 1273 24028
rect 1239 23921 1273 23955
rect 1239 23848 1273 23882
rect 1239 23775 1273 23809
rect 1239 23702 1273 23736
rect 1239 23629 1273 23663
rect 1239 23556 1273 23590
rect 1239 23483 1273 23517
rect 1239 23410 1273 23444
rect 1239 23337 1273 23371
rect 1239 23264 1273 23298
rect 1239 23191 1273 23225
rect 1239 23118 1273 23152
rect 1239 23044 1273 23078
rect 1239 22970 1273 23004
rect 1239 22896 1273 22930
rect 1239 22822 1273 22856
rect 1239 22748 1273 22782
rect 1239 22674 1273 22708
rect 1239 22600 1273 22634
rect 1239 22526 1273 22560
rect 1239 22452 1273 22486
rect 1239 22378 1273 22412
rect 1239 22304 1273 22338
rect 1239 22230 1273 22264
rect 1239 22156 1273 22190
rect 1239 22082 1273 22116
rect 1475 23994 1509 24028
rect 1475 23921 1509 23955
rect 1475 23848 1509 23882
rect 1475 23775 1509 23809
rect 1475 23702 1509 23736
rect 1475 23629 1509 23663
rect 1475 23556 1509 23590
rect 1475 23483 1509 23517
rect 1475 23410 1509 23444
rect 1475 23337 1509 23371
rect 1475 23264 1509 23298
rect 1475 23191 1509 23225
rect 1475 23118 1509 23152
rect 1475 23044 1509 23078
rect 1475 22970 1509 23004
rect 1475 22896 1509 22930
rect 1475 22822 1509 22856
rect 1475 22748 1509 22782
rect 1475 22674 1509 22708
rect 1475 22600 1509 22634
rect 1475 22526 1509 22560
rect 1475 22452 1509 22486
rect 1475 22378 1509 22412
rect 1475 22304 1509 22338
rect 1475 22230 1509 22264
rect 1475 22156 1509 22190
rect 1475 22082 1509 22116
rect 1711 23994 1745 24028
rect 1711 23921 1745 23955
rect 1711 23848 1745 23882
rect 1711 23775 1745 23809
rect 1711 23702 1745 23736
rect 1711 23629 1745 23663
rect 1711 23556 1745 23590
rect 1711 23483 1745 23517
rect 1711 23410 1745 23444
rect 1711 23337 1745 23371
rect 1711 23264 1745 23298
rect 1711 23191 1745 23225
rect 1711 23118 1745 23152
rect 1711 23044 1745 23078
rect 1711 22970 1745 23004
rect 1711 22896 1745 22930
rect 1711 22822 1745 22856
rect 1711 22748 1745 22782
rect 1711 22674 1745 22708
rect 1711 22600 1745 22634
rect 1711 22526 1745 22560
rect 1711 22452 1745 22486
rect 1711 22378 1745 22412
rect 1711 22304 1745 22338
rect 1711 22230 1745 22264
rect 1711 22156 1745 22190
rect 1711 22082 1745 22116
rect 1947 23994 1981 24028
rect 1947 23921 1981 23955
rect 1947 23848 1981 23882
rect 1947 23775 1981 23809
rect 1947 23702 1981 23736
rect 1947 23629 1981 23663
rect 1947 23556 1981 23590
rect 1947 23483 1981 23517
rect 1947 23410 1981 23444
rect 1947 23337 1981 23371
rect 1947 23264 1981 23298
rect 1947 23191 1981 23225
rect 1947 23118 1981 23152
rect 1947 23044 1981 23078
rect 1947 22970 1981 23004
rect 1947 22896 1981 22930
rect 1947 22822 1981 22856
rect 1947 22748 1981 22782
rect 1947 22674 1981 22708
rect 1947 22600 1981 22634
rect 1947 22526 1981 22560
rect 1947 22452 1981 22486
rect 1947 22378 1981 22412
rect 1947 22304 1981 22338
rect 1947 22230 1981 22264
rect 1947 22156 1981 22190
rect 1947 22082 1981 22116
rect 2183 23994 2217 24028
rect 2183 23921 2217 23955
rect 2183 23848 2217 23882
rect 2183 23775 2217 23809
rect 2183 23702 2217 23736
rect 2183 23629 2217 23663
rect 2183 23556 2217 23590
rect 2183 23483 2217 23517
rect 2183 23410 2217 23444
rect 2183 23337 2217 23371
rect 2183 23264 2217 23298
rect 2183 23191 2217 23225
rect 2183 23118 2217 23152
rect 2183 23044 2217 23078
rect 2183 22970 2217 23004
rect 2183 22896 2217 22930
rect 2183 22822 2217 22856
rect 2183 22748 2217 22782
rect 2183 22674 2217 22708
rect 2183 22600 2217 22634
rect 2183 22526 2217 22560
rect 2183 22452 2217 22486
rect 2183 22378 2217 22412
rect 2183 22304 2217 22338
rect 2183 22230 2217 22264
rect 2183 22156 2217 22190
rect 2183 22082 2217 22116
rect 2419 23994 2453 24028
rect 2419 23921 2453 23955
rect 2419 23848 2453 23882
rect 2419 23775 2453 23809
rect 2419 23702 2453 23736
rect 2419 23629 2453 23663
rect 2419 23556 2453 23590
rect 2419 23483 2453 23517
rect 2419 23410 2453 23444
rect 2419 23337 2453 23371
rect 2419 23264 2453 23298
rect 2419 23191 2453 23225
rect 2419 23118 2453 23152
rect 2419 23044 2453 23078
rect 2419 22970 2453 23004
rect 2419 22896 2453 22930
rect 2419 22822 2453 22856
rect 2419 22748 2453 22782
rect 2419 22674 2453 22708
rect 2419 22600 2453 22634
rect 2419 22526 2453 22560
rect 2419 22452 2453 22486
rect 2419 22378 2453 22412
rect 2419 22304 2453 22338
rect 2419 22230 2453 22264
rect 2419 22156 2453 22190
rect 2419 22082 2453 22116
rect 2655 23994 2689 24028
rect 2655 23921 2689 23955
rect 2655 23848 2689 23882
rect 2655 23775 2689 23809
rect 2655 23702 2689 23736
rect 2655 23629 2689 23663
rect 2655 23556 2689 23590
rect 2655 23483 2689 23517
rect 2655 23410 2689 23444
rect 2655 23337 2689 23371
rect 2655 23264 2689 23298
rect 2655 23191 2689 23225
rect 2655 23118 2689 23152
rect 2655 23044 2689 23078
rect 2655 22970 2689 23004
rect 2655 22896 2689 22930
rect 2655 22822 2689 22856
rect 2655 22748 2689 22782
rect 2655 22674 2689 22708
rect 2655 22600 2689 22634
rect 2655 22526 2689 22560
rect 2655 22452 2689 22486
rect 2655 22378 2689 22412
rect 2655 22304 2689 22338
rect 2655 22230 2689 22264
rect 2655 22156 2689 22190
rect 2655 22082 2689 22116
rect 2891 23994 2925 24028
rect 2891 23921 2925 23955
rect 2891 23848 2925 23882
rect 2891 23775 2925 23809
rect 2891 23702 2925 23736
rect 2891 23629 2925 23663
rect 2891 23556 2925 23590
rect 2891 23483 2925 23517
rect 2891 23410 2925 23444
rect 2891 23337 2925 23371
rect 2891 23264 2925 23298
rect 2891 23191 2925 23225
rect 2891 23118 2925 23152
rect 2891 23044 2925 23078
rect 2891 22970 2925 23004
rect 2891 22896 2925 22930
rect 2891 22822 2925 22856
rect 2891 22748 2925 22782
rect 2891 22674 2925 22708
rect 2891 22600 2925 22634
rect 2891 22526 2925 22560
rect 2891 22452 2925 22486
rect 2891 22378 2925 22412
rect 2891 22304 2925 22338
rect 2891 22230 2925 22264
rect 2891 22156 2925 22190
rect 2891 22082 2925 22116
rect 3036 24048 3070 24058
rect 3036 24024 3070 24048
rect 3036 23980 3070 23986
rect 3036 23952 3070 23980
rect 3036 23912 3070 23914
rect 3036 23880 3070 23912
rect 3036 23810 3070 23842
rect 3036 23808 3070 23810
rect 3036 23742 3070 23770
rect 3036 23736 3070 23742
rect 3036 23674 3070 23698
rect 3036 23664 3070 23674
rect 3036 23606 3070 23626
rect 3036 23592 3070 23606
rect 3036 23538 3070 23554
rect 3036 23520 3070 23538
rect 3036 23470 3070 23482
rect 3036 23448 3070 23470
rect 3036 23402 3070 23410
rect 3036 23376 3070 23402
rect 3036 23334 3070 23338
rect 3036 23304 3070 23334
rect 3036 23232 3070 23266
rect 3036 23164 3070 23194
rect 3036 23160 3070 23164
rect 3036 23096 3070 23122
rect 3036 23088 3070 23096
rect 3036 23028 3070 23050
rect 3036 23016 3070 23028
rect 3036 22960 3070 22978
rect 3036 22944 3070 22960
rect 3036 22892 3070 22906
rect 3036 22872 3070 22892
rect 3036 22824 3070 22834
rect 3036 22800 3070 22824
rect 3036 22756 3070 22762
rect 3036 22728 3070 22756
rect 3036 22688 3070 22690
rect 3036 22656 3070 22688
rect 3036 22586 3070 22618
rect 3036 22584 3070 22586
rect 3036 22518 3070 22546
rect 3036 22512 3070 22518
rect 3036 22450 3070 22474
rect 3036 22440 3070 22450
rect 3036 22382 3070 22402
rect 3036 22368 3070 22382
rect 3036 22314 3070 22330
rect 3036 22296 3070 22314
rect 3036 22246 3070 22258
rect 3036 22224 3070 22246
rect 3036 22178 3070 22186
rect 3036 22152 3070 22178
rect 386 22021 420 22023
rect 386 21989 420 22021
rect 3036 22110 3070 22114
rect 3036 22080 3070 22110
rect 625 21980 626 22014
rect 626 21980 659 22014
rect 700 21980 732 22014
rect 732 21980 734 22014
rect 775 21980 802 22014
rect 802 21980 809 22014
rect 850 21980 872 22014
rect 872 21980 884 22014
rect 925 21980 942 22014
rect 942 21980 959 22014
rect 1000 21980 1012 22014
rect 1012 21980 1034 22014
rect 1075 21980 1082 22014
rect 1082 21980 1109 22014
rect 1150 21980 1152 22014
rect 1152 21980 1184 22014
rect 1225 21980 1256 22014
rect 1256 21980 1259 22014
rect 1300 21980 1326 22014
rect 1326 21980 1334 22014
rect 1375 21980 1396 22014
rect 1396 21980 1409 22014
rect 1450 21980 1466 22014
rect 1466 21980 1484 22014
rect 1525 21980 1536 22014
rect 1536 21980 1559 22014
rect 1600 21980 1606 22014
rect 1606 21980 1634 22014
rect 1674 21980 1676 22014
rect 1676 21980 1708 22014
rect 1748 21980 1782 22014
rect 1822 21980 1852 22014
rect 1852 21980 1856 22014
rect 1896 21980 1922 22014
rect 1922 21980 1930 22014
rect 1970 21980 1992 22014
rect 1992 21980 2004 22014
rect 2044 21980 2062 22014
rect 2062 21980 2078 22014
rect 2118 21980 2132 22014
rect 2132 21980 2152 22014
rect 2192 21980 2202 22014
rect 2202 21980 2226 22014
rect 2266 21980 2272 22014
rect 2272 21980 2300 22014
rect 2340 21980 2342 22014
rect 2342 21980 2374 22014
rect 2414 21980 2446 22014
rect 2446 21980 2448 22014
rect 2488 21980 2516 22014
rect 2516 21980 2522 22014
rect 2562 21980 2586 22014
rect 2586 21980 2596 22014
rect 2636 21980 2656 22014
rect 2656 21980 2670 22014
rect 2710 21980 2726 22014
rect 2726 21980 2744 22014
rect 2784 21980 2795 22014
rect 2795 21980 2818 22014
rect 3036 22008 3070 22042
rect 386 21919 420 21951
rect 386 21917 420 21919
rect 3036 21940 3070 21970
rect 3036 21936 3070 21940
rect 386 21851 420 21879
rect 386 21845 420 21851
rect 386 21783 420 21807
rect 386 21773 420 21783
rect 386 21715 420 21735
rect 386 21701 420 21715
rect 386 21647 420 21663
rect 386 21629 420 21647
rect 386 21579 420 21591
rect 386 21557 420 21579
rect 386 21511 420 21519
rect 386 21485 420 21511
rect 386 21443 420 21447
rect 386 21413 420 21443
rect 386 21341 420 21375
rect 386 21273 420 21303
rect 386 21269 420 21273
rect 386 21205 420 21231
rect 386 21197 420 21205
rect 386 21137 420 21159
rect 386 21125 420 21137
rect 386 21069 420 21087
rect 386 21053 420 21069
rect 386 21001 420 21015
rect 386 20981 420 21001
rect 386 20933 420 20943
rect 386 20909 420 20933
rect 386 20865 420 20871
rect 386 20837 420 20865
rect 386 20797 420 20799
rect 386 20765 420 20797
rect 386 20695 420 20727
rect 386 20693 420 20695
rect 386 20627 420 20655
rect 386 20621 420 20627
rect 386 20559 420 20583
rect 386 20549 420 20559
rect 386 20491 420 20511
rect 386 20477 420 20491
rect 386 20423 420 20439
rect 386 20405 420 20423
rect 386 20355 420 20367
rect 386 20333 420 20355
rect 386 20287 420 20295
rect 386 20261 420 20287
rect 386 20219 420 20223
rect 386 20189 420 20219
rect 386 20117 420 20151
rect 386 20049 420 20079
rect 386 20045 420 20049
rect 386 19981 420 20007
rect 386 19973 420 19981
rect 531 21878 565 21912
rect 531 21805 565 21839
rect 531 21732 565 21766
rect 531 21659 565 21693
rect 531 21586 565 21620
rect 531 21513 565 21547
rect 531 21440 565 21474
rect 531 21367 565 21401
rect 531 21294 565 21328
rect 531 21221 565 21255
rect 531 21148 565 21182
rect 531 21075 565 21109
rect 531 21002 565 21036
rect 531 20928 565 20962
rect 531 20854 565 20888
rect 531 20780 565 20814
rect 531 20706 565 20740
rect 531 20632 565 20666
rect 531 20558 565 20592
rect 531 20484 565 20518
rect 531 20410 565 20444
rect 531 20336 565 20370
rect 531 20262 565 20296
rect 531 20188 565 20222
rect 531 20114 565 20148
rect 531 20040 565 20074
rect 531 19966 565 20000
rect 767 21878 801 21912
rect 767 21805 801 21839
rect 767 21732 801 21766
rect 767 21659 801 21693
rect 767 21586 801 21620
rect 767 21513 801 21547
rect 767 21440 801 21474
rect 767 21367 801 21401
rect 767 21294 801 21328
rect 767 21221 801 21255
rect 767 21148 801 21182
rect 767 21075 801 21109
rect 767 21002 801 21036
rect 767 20928 801 20962
rect 767 20854 801 20888
rect 767 20780 801 20814
rect 767 20706 801 20740
rect 767 20632 801 20666
rect 767 20558 801 20592
rect 767 20484 801 20518
rect 767 20410 801 20444
rect 767 20336 801 20370
rect 767 20262 801 20296
rect 767 20188 801 20222
rect 767 20114 801 20148
rect 767 20040 801 20074
rect 767 19966 801 20000
rect 1003 21878 1037 21912
rect 1003 21805 1037 21839
rect 1003 21732 1037 21766
rect 1003 21659 1037 21693
rect 1003 21586 1037 21620
rect 1003 21513 1037 21547
rect 1003 21440 1037 21474
rect 1003 21367 1037 21401
rect 1003 21294 1037 21328
rect 1003 21221 1037 21255
rect 1003 21148 1037 21182
rect 1003 21075 1037 21109
rect 1003 21002 1037 21036
rect 1003 20928 1037 20962
rect 1003 20854 1037 20888
rect 1003 20780 1037 20814
rect 1003 20706 1037 20740
rect 1003 20632 1037 20666
rect 1003 20558 1037 20592
rect 1003 20484 1037 20518
rect 1003 20410 1037 20444
rect 1003 20336 1037 20370
rect 1003 20262 1037 20296
rect 1003 20188 1037 20222
rect 1003 20114 1037 20148
rect 1003 20040 1037 20074
rect 1003 19966 1037 20000
rect 1239 21878 1273 21912
rect 1239 21805 1273 21839
rect 1239 21732 1273 21766
rect 1239 21659 1273 21693
rect 1239 21586 1273 21620
rect 1239 21513 1273 21547
rect 1239 21440 1273 21474
rect 1239 21367 1273 21401
rect 1239 21294 1273 21328
rect 1239 21221 1273 21255
rect 1239 21148 1273 21182
rect 1239 21075 1273 21109
rect 1239 21002 1273 21036
rect 1239 20928 1273 20962
rect 1239 20854 1273 20888
rect 1239 20780 1273 20814
rect 1239 20706 1273 20740
rect 1239 20632 1273 20666
rect 1239 20558 1273 20592
rect 1239 20484 1273 20518
rect 1239 20410 1273 20444
rect 1239 20336 1273 20370
rect 1239 20262 1273 20296
rect 1239 20188 1273 20222
rect 1239 20114 1273 20148
rect 1239 20040 1273 20074
rect 1239 19966 1273 20000
rect 1475 21878 1509 21912
rect 1475 21805 1509 21839
rect 1475 21732 1509 21766
rect 1475 21659 1509 21693
rect 1475 21586 1509 21620
rect 1475 21513 1509 21547
rect 1475 21440 1509 21474
rect 1475 21367 1509 21401
rect 1475 21294 1509 21328
rect 1475 21221 1509 21255
rect 1475 21148 1509 21182
rect 1475 21075 1509 21109
rect 1475 21002 1509 21036
rect 1475 20928 1509 20962
rect 1475 20854 1509 20888
rect 1475 20780 1509 20814
rect 1475 20706 1509 20740
rect 1475 20632 1509 20666
rect 1475 20558 1509 20592
rect 1475 20484 1509 20518
rect 1475 20410 1509 20444
rect 1475 20336 1509 20370
rect 1475 20262 1509 20296
rect 1475 20188 1509 20222
rect 1475 20114 1509 20148
rect 1475 20040 1509 20074
rect 1475 19966 1509 20000
rect 1711 21878 1745 21912
rect 1711 21805 1745 21839
rect 1711 21732 1745 21766
rect 1711 21659 1745 21693
rect 1711 21586 1745 21620
rect 1711 21513 1745 21547
rect 1711 21440 1745 21474
rect 1711 21367 1745 21401
rect 1711 21294 1745 21328
rect 1711 21221 1745 21255
rect 1711 21148 1745 21182
rect 1711 21075 1745 21109
rect 1711 21002 1745 21036
rect 1711 20928 1745 20962
rect 1711 20854 1745 20888
rect 1711 20780 1745 20814
rect 1711 20706 1745 20740
rect 1711 20632 1745 20666
rect 1711 20558 1745 20592
rect 1711 20484 1745 20518
rect 1711 20410 1745 20444
rect 1711 20336 1745 20370
rect 1711 20262 1745 20296
rect 1711 20188 1745 20222
rect 1711 20114 1745 20148
rect 1711 20040 1745 20074
rect 1711 19966 1745 20000
rect 1947 21878 1981 21912
rect 1947 21805 1981 21839
rect 1947 21732 1981 21766
rect 1947 21659 1981 21693
rect 1947 21586 1981 21620
rect 1947 21513 1981 21547
rect 1947 21440 1981 21474
rect 1947 21367 1981 21401
rect 1947 21294 1981 21328
rect 1947 21221 1981 21255
rect 1947 21148 1981 21182
rect 1947 21075 1981 21109
rect 1947 21002 1981 21036
rect 1947 20928 1981 20962
rect 1947 20854 1981 20888
rect 1947 20780 1981 20814
rect 1947 20706 1981 20740
rect 1947 20632 1981 20666
rect 1947 20558 1981 20592
rect 1947 20484 1981 20518
rect 1947 20410 1981 20444
rect 1947 20336 1981 20370
rect 1947 20262 1981 20296
rect 1947 20188 1981 20222
rect 1947 20114 1981 20148
rect 1947 20040 1981 20074
rect 1947 19966 1981 20000
rect 2183 21878 2217 21912
rect 2183 21805 2217 21839
rect 2183 21732 2217 21766
rect 2183 21659 2217 21693
rect 2183 21586 2217 21620
rect 2183 21513 2217 21547
rect 2183 21440 2217 21474
rect 2183 21367 2217 21401
rect 2183 21294 2217 21328
rect 2183 21221 2217 21255
rect 2183 21148 2217 21182
rect 2183 21075 2217 21109
rect 2183 21002 2217 21036
rect 2183 20928 2217 20962
rect 2183 20854 2217 20888
rect 2183 20780 2217 20814
rect 2183 20706 2217 20740
rect 2183 20632 2217 20666
rect 2183 20558 2217 20592
rect 2183 20484 2217 20518
rect 2183 20410 2217 20444
rect 2183 20336 2217 20370
rect 2183 20262 2217 20296
rect 2183 20188 2217 20222
rect 2183 20114 2217 20148
rect 2183 20040 2217 20074
rect 2183 19966 2217 20000
rect 2419 21878 2453 21912
rect 2419 21805 2453 21839
rect 2419 21732 2453 21766
rect 2419 21659 2453 21693
rect 2419 21586 2453 21620
rect 2419 21513 2453 21547
rect 2419 21440 2453 21474
rect 2419 21367 2453 21401
rect 2419 21294 2453 21328
rect 2419 21221 2453 21255
rect 2419 21148 2453 21182
rect 2419 21075 2453 21109
rect 2419 21002 2453 21036
rect 2419 20928 2453 20962
rect 2419 20854 2453 20888
rect 2419 20780 2453 20814
rect 2419 20706 2453 20740
rect 2419 20632 2453 20666
rect 2419 20558 2453 20592
rect 2419 20484 2453 20518
rect 2419 20410 2453 20444
rect 2419 20336 2453 20370
rect 2419 20262 2453 20296
rect 2419 20188 2453 20222
rect 2419 20114 2453 20148
rect 2419 20040 2453 20074
rect 2419 19966 2453 20000
rect 2655 21878 2689 21912
rect 2655 21805 2689 21839
rect 2655 21732 2689 21766
rect 2655 21659 2689 21693
rect 2655 21586 2689 21620
rect 2655 21513 2689 21547
rect 2655 21440 2689 21474
rect 2655 21367 2689 21401
rect 2655 21294 2689 21328
rect 2655 21221 2689 21255
rect 2655 21148 2689 21182
rect 2655 21075 2689 21109
rect 2655 21002 2689 21036
rect 2655 20928 2689 20962
rect 2655 20854 2689 20888
rect 2655 20780 2689 20814
rect 2655 20706 2689 20740
rect 2655 20632 2689 20666
rect 2655 20558 2689 20592
rect 2655 20484 2689 20518
rect 2655 20410 2689 20444
rect 2655 20336 2689 20370
rect 2655 20262 2689 20296
rect 2655 20188 2689 20222
rect 2655 20114 2689 20148
rect 2655 20040 2689 20074
rect 2655 19966 2689 20000
rect 2891 21878 2925 21912
rect 2891 21805 2925 21839
rect 2891 21732 2925 21766
rect 2891 21659 2925 21693
rect 2891 21586 2925 21620
rect 2891 21513 2925 21547
rect 2891 21440 2925 21474
rect 2891 21367 2925 21401
rect 2891 21294 2925 21328
rect 2891 21221 2925 21255
rect 2891 21148 2925 21182
rect 2891 21075 2925 21109
rect 2891 21002 2925 21036
rect 2891 20928 2925 20962
rect 2891 20854 2925 20888
rect 2891 20780 2925 20814
rect 2891 20706 2925 20740
rect 2891 20632 2925 20666
rect 2891 20558 2925 20592
rect 2891 20484 2925 20518
rect 2891 20410 2925 20444
rect 2891 20336 2925 20370
rect 2891 20262 2925 20296
rect 2891 20188 2925 20222
rect 2891 20114 2925 20148
rect 2891 20040 2925 20074
rect 2891 19966 2925 20000
rect 3036 21872 3070 21898
rect 3036 21864 3070 21872
rect 3036 21804 3070 21826
rect 3036 21792 3070 21804
rect 3036 21736 3070 21754
rect 3036 21720 3070 21736
rect 3036 21668 3070 21682
rect 3036 21648 3070 21668
rect 3036 21600 3070 21610
rect 3036 21576 3070 21600
rect 3036 21532 3070 21538
rect 3036 21504 3070 21532
rect 3036 21464 3070 21466
rect 3036 21432 3070 21464
rect 3036 21362 3070 21394
rect 3036 21360 3070 21362
rect 3036 21294 3070 21322
rect 3036 21288 3070 21294
rect 3036 21226 3070 21250
rect 3036 21216 3070 21226
rect 3036 21158 3070 21178
rect 3036 21144 3070 21158
rect 3036 21090 3070 21106
rect 3036 21072 3070 21090
rect 3036 21022 3070 21034
rect 3036 21000 3070 21022
rect 3036 20954 3070 20962
rect 3036 20928 3070 20954
rect 3036 20886 3070 20890
rect 3036 20856 3070 20886
rect 3036 20784 3070 20818
rect 3036 20716 3070 20746
rect 3036 20712 3070 20716
rect 3036 20648 3070 20674
rect 3036 20640 3070 20648
rect 3036 20580 3070 20602
rect 3036 20568 3070 20580
rect 3036 20512 3070 20530
rect 3036 20496 3070 20512
rect 3036 20444 3070 20458
rect 3036 20424 3070 20444
rect 3036 20376 3070 20386
rect 3036 20352 3070 20376
rect 3036 20308 3070 20314
rect 3036 20280 3070 20308
rect 3036 20240 3070 20242
rect 3036 20208 3070 20240
rect 3036 20138 3070 20170
rect 3036 20136 3070 20138
rect 3036 20070 3070 20098
rect 3036 20064 3070 20070
rect 3036 20002 3070 20026
rect 3036 19992 3070 20002
rect 386 19913 420 19935
rect 386 19901 420 19913
rect 3036 19934 3070 19954
rect 3036 19920 3070 19934
rect 386 19845 420 19863
rect 386 19829 420 19845
rect 625 19850 626 19884
rect 626 19850 659 19884
rect 700 19850 732 19884
rect 732 19850 734 19884
rect 775 19850 802 19884
rect 802 19850 809 19884
rect 850 19850 872 19884
rect 872 19850 884 19884
rect 925 19850 942 19884
rect 942 19850 959 19884
rect 1000 19850 1012 19884
rect 1012 19850 1034 19884
rect 1075 19850 1082 19884
rect 1082 19850 1109 19884
rect 1150 19850 1152 19884
rect 1152 19850 1184 19884
rect 1225 19850 1256 19884
rect 1256 19850 1259 19884
rect 1300 19850 1326 19884
rect 1326 19850 1334 19884
rect 1375 19850 1396 19884
rect 1396 19850 1409 19884
rect 1450 19850 1466 19884
rect 1466 19850 1484 19884
rect 1525 19850 1536 19884
rect 1536 19850 1559 19884
rect 1600 19850 1606 19884
rect 1606 19850 1634 19884
rect 1674 19850 1676 19884
rect 1676 19850 1708 19884
rect 1748 19850 1782 19884
rect 1822 19850 1852 19884
rect 1852 19850 1856 19884
rect 1896 19850 1922 19884
rect 1922 19850 1930 19884
rect 1970 19850 1992 19884
rect 1992 19850 2004 19884
rect 2044 19850 2062 19884
rect 2062 19850 2078 19884
rect 2118 19850 2132 19884
rect 2132 19850 2152 19884
rect 2192 19850 2202 19884
rect 2202 19850 2226 19884
rect 2266 19850 2272 19884
rect 2272 19850 2300 19884
rect 2340 19850 2342 19884
rect 2342 19850 2374 19884
rect 2414 19850 2446 19884
rect 2446 19850 2448 19884
rect 2488 19850 2516 19884
rect 2516 19850 2522 19884
rect 2562 19850 2586 19884
rect 2586 19850 2596 19884
rect 2636 19850 2656 19884
rect 2656 19850 2670 19884
rect 2710 19850 2726 19884
rect 2726 19850 2744 19884
rect 2784 19850 2795 19884
rect 2795 19850 2818 19884
rect 386 19777 420 19791
rect 386 19757 420 19777
rect 3036 19866 3070 19882
rect 3036 19848 3070 19866
rect 386 19709 420 19719
rect 386 19685 420 19709
rect 386 19641 420 19647
rect 386 19613 420 19641
rect 386 19573 420 19575
rect 386 19541 420 19573
rect 386 19471 420 19503
rect 386 19469 420 19471
rect 386 19403 420 19431
rect 386 19397 420 19403
rect 386 19335 420 19359
rect 386 19325 420 19335
rect 386 19267 420 19287
rect 386 19253 420 19267
rect 386 19199 420 19215
rect 386 19181 420 19199
rect 386 19131 420 19143
rect 386 19109 420 19131
rect 386 19063 420 19071
rect 386 19037 420 19063
rect 386 18995 420 18999
rect 386 18965 420 18995
rect 386 18893 420 18927
rect 386 18825 420 18855
rect 386 18821 420 18825
rect 386 18757 420 18783
rect 386 18749 420 18757
rect 386 18689 420 18711
rect 386 18677 420 18689
rect 386 18621 420 18639
rect 386 18605 420 18621
rect 386 18553 420 18567
rect 386 18533 420 18553
rect 386 18485 420 18495
rect 386 18461 420 18485
rect 386 18417 420 18423
rect 386 18389 420 18417
rect 386 18349 420 18351
rect 386 18317 420 18349
rect 386 18247 420 18279
rect 386 18245 420 18247
rect 386 18179 420 18207
rect 386 18173 420 18179
rect 386 18111 420 18135
rect 386 18101 420 18111
rect 386 18043 420 18063
rect 386 18029 420 18043
rect 386 17975 420 17991
rect 386 17957 420 17975
rect 386 17907 420 17919
rect 386 17885 420 17907
rect 386 17839 420 17847
rect 386 17813 420 17839
rect 531 19734 565 19768
rect 531 19661 565 19695
rect 531 19588 565 19622
rect 531 19515 565 19549
rect 531 19442 565 19476
rect 531 19369 565 19403
rect 531 19296 565 19330
rect 531 19223 565 19257
rect 531 19150 565 19184
rect 531 19077 565 19111
rect 531 19004 565 19038
rect 531 18931 565 18965
rect 531 18858 565 18892
rect 531 18784 565 18818
rect 531 18710 565 18744
rect 531 18636 565 18670
rect 531 18562 565 18596
rect 531 18488 565 18522
rect 531 18414 565 18448
rect 531 18340 565 18374
rect 531 18266 565 18300
rect 531 18192 565 18226
rect 531 18118 565 18152
rect 531 18044 565 18078
rect 531 17970 565 18004
rect 531 17896 565 17930
rect 531 17822 565 17856
rect 767 19734 801 19768
rect 767 19661 801 19695
rect 767 19588 801 19622
rect 767 19515 801 19549
rect 767 19442 801 19476
rect 767 19369 801 19403
rect 767 19296 801 19330
rect 767 19223 801 19257
rect 767 19150 801 19184
rect 767 19077 801 19111
rect 767 19004 801 19038
rect 767 18931 801 18965
rect 767 18858 801 18892
rect 767 18784 801 18818
rect 767 18710 801 18744
rect 767 18636 801 18670
rect 767 18562 801 18596
rect 767 18488 801 18522
rect 767 18414 801 18448
rect 767 18340 801 18374
rect 767 18266 801 18300
rect 767 18192 801 18226
rect 767 18118 801 18152
rect 767 18044 801 18078
rect 767 17970 801 18004
rect 767 17896 801 17930
rect 767 17822 801 17856
rect 1003 19734 1037 19768
rect 1003 19661 1037 19695
rect 1003 19588 1037 19622
rect 1003 19515 1037 19549
rect 1003 19442 1037 19476
rect 1003 19369 1037 19403
rect 1003 19296 1037 19330
rect 1003 19223 1037 19257
rect 1003 19150 1037 19184
rect 1003 19077 1037 19111
rect 1003 19004 1037 19038
rect 1003 18931 1037 18965
rect 1003 18858 1037 18892
rect 1003 18784 1037 18818
rect 1003 18710 1037 18744
rect 1003 18636 1037 18670
rect 1003 18562 1037 18596
rect 1003 18488 1037 18522
rect 1003 18414 1037 18448
rect 1003 18340 1037 18374
rect 1003 18266 1037 18300
rect 1003 18192 1037 18226
rect 1003 18118 1037 18152
rect 1003 18044 1037 18078
rect 1003 17970 1037 18004
rect 1003 17896 1037 17930
rect 1003 17822 1037 17856
rect 1239 19734 1273 19768
rect 1239 19661 1273 19695
rect 1239 19588 1273 19622
rect 1239 19515 1273 19549
rect 1239 19442 1273 19476
rect 1239 19369 1273 19403
rect 1239 19296 1273 19330
rect 1239 19223 1273 19257
rect 1239 19150 1273 19184
rect 1239 19077 1273 19111
rect 1239 19004 1273 19038
rect 1239 18931 1273 18965
rect 1239 18858 1273 18892
rect 1239 18784 1273 18818
rect 1239 18710 1273 18744
rect 1239 18636 1273 18670
rect 1239 18562 1273 18596
rect 1239 18488 1273 18522
rect 1239 18414 1273 18448
rect 1239 18340 1273 18374
rect 1239 18266 1273 18300
rect 1239 18192 1273 18226
rect 1239 18118 1273 18152
rect 1239 18044 1273 18078
rect 1239 17970 1273 18004
rect 1239 17896 1273 17930
rect 1239 17822 1273 17856
rect 1475 19734 1509 19768
rect 1475 19661 1509 19695
rect 1475 19588 1509 19622
rect 1475 19515 1509 19549
rect 1475 19442 1509 19476
rect 1475 19369 1509 19403
rect 1475 19296 1509 19330
rect 1475 19223 1509 19257
rect 1475 19150 1509 19184
rect 1475 19077 1509 19111
rect 1475 19004 1509 19038
rect 1475 18931 1509 18965
rect 1475 18858 1509 18892
rect 1475 18784 1509 18818
rect 1475 18710 1509 18744
rect 1475 18636 1509 18670
rect 1475 18562 1509 18596
rect 1475 18488 1509 18522
rect 1475 18414 1509 18448
rect 1475 18340 1509 18374
rect 1475 18266 1509 18300
rect 1475 18192 1509 18226
rect 1475 18118 1509 18152
rect 1475 18044 1509 18078
rect 1475 17970 1509 18004
rect 1475 17896 1509 17930
rect 1475 17822 1509 17856
rect 1711 19734 1745 19768
rect 1711 19661 1745 19695
rect 1711 19588 1745 19622
rect 1711 19515 1745 19549
rect 1711 19442 1745 19476
rect 1711 19369 1745 19403
rect 1711 19296 1745 19330
rect 1711 19223 1745 19257
rect 1711 19150 1745 19184
rect 1711 19077 1745 19111
rect 1711 19004 1745 19038
rect 1711 18931 1745 18965
rect 1711 18858 1745 18892
rect 1711 18784 1745 18818
rect 1711 18710 1745 18744
rect 1711 18636 1745 18670
rect 1711 18562 1745 18596
rect 1711 18488 1745 18522
rect 1711 18414 1745 18448
rect 1711 18340 1745 18374
rect 1711 18266 1745 18300
rect 1711 18192 1745 18226
rect 1711 18118 1745 18152
rect 1711 18044 1745 18078
rect 1711 17970 1745 18004
rect 1711 17896 1745 17930
rect 1711 17822 1745 17856
rect 1947 19734 1981 19768
rect 1947 19661 1981 19695
rect 1947 19588 1981 19622
rect 1947 19515 1981 19549
rect 1947 19442 1981 19476
rect 1947 19369 1981 19403
rect 1947 19296 1981 19330
rect 1947 19223 1981 19257
rect 1947 19150 1981 19184
rect 1947 19077 1981 19111
rect 1947 19004 1981 19038
rect 1947 18931 1981 18965
rect 1947 18858 1981 18892
rect 1947 18784 1981 18818
rect 1947 18710 1981 18744
rect 1947 18636 1981 18670
rect 1947 18562 1981 18596
rect 1947 18488 1981 18522
rect 1947 18414 1981 18448
rect 1947 18340 1981 18374
rect 1947 18266 1981 18300
rect 1947 18192 1981 18226
rect 1947 18118 1981 18152
rect 1947 18044 1981 18078
rect 1947 17970 1981 18004
rect 1947 17896 1981 17930
rect 1947 17822 1981 17856
rect 2183 19734 2217 19768
rect 2183 19661 2217 19695
rect 2183 19588 2217 19622
rect 2183 19515 2217 19549
rect 2183 19442 2217 19476
rect 2183 19369 2217 19403
rect 2183 19296 2217 19330
rect 2183 19223 2217 19257
rect 2183 19150 2217 19184
rect 2183 19077 2217 19111
rect 2183 19004 2217 19038
rect 2183 18931 2217 18965
rect 2183 18858 2217 18892
rect 2183 18784 2217 18818
rect 2183 18710 2217 18744
rect 2183 18636 2217 18670
rect 2183 18562 2217 18596
rect 2183 18488 2217 18522
rect 2183 18414 2217 18448
rect 2183 18340 2217 18374
rect 2183 18266 2217 18300
rect 2183 18192 2217 18226
rect 2183 18118 2217 18152
rect 2183 18044 2217 18078
rect 2183 17970 2217 18004
rect 2183 17896 2217 17930
rect 2183 17822 2217 17856
rect 2419 19734 2453 19768
rect 2419 19661 2453 19695
rect 2419 19588 2453 19622
rect 2419 19515 2453 19549
rect 2419 19442 2453 19476
rect 2419 19369 2453 19403
rect 2419 19296 2453 19330
rect 2419 19223 2453 19257
rect 2419 19150 2453 19184
rect 2419 19077 2453 19111
rect 2419 19004 2453 19038
rect 2419 18931 2453 18965
rect 2419 18858 2453 18892
rect 2419 18784 2453 18818
rect 2419 18710 2453 18744
rect 2419 18636 2453 18670
rect 2419 18562 2453 18596
rect 2419 18488 2453 18522
rect 2419 18414 2453 18448
rect 2419 18340 2453 18374
rect 2419 18266 2453 18300
rect 2419 18192 2453 18226
rect 2419 18118 2453 18152
rect 2419 18044 2453 18078
rect 2419 17970 2453 18004
rect 2419 17896 2453 17930
rect 2419 17822 2453 17856
rect 2655 19734 2689 19768
rect 2655 19661 2689 19695
rect 2655 19588 2689 19622
rect 2655 19515 2689 19549
rect 2655 19442 2689 19476
rect 2655 19369 2689 19403
rect 2655 19296 2689 19330
rect 2655 19223 2689 19257
rect 2655 19150 2689 19184
rect 2655 19077 2689 19111
rect 2655 19004 2689 19038
rect 2655 18931 2689 18965
rect 2655 18858 2689 18892
rect 2655 18784 2689 18818
rect 2655 18710 2689 18744
rect 2655 18636 2689 18670
rect 2655 18562 2689 18596
rect 2655 18488 2689 18522
rect 2655 18414 2689 18448
rect 2655 18340 2689 18374
rect 2655 18266 2689 18300
rect 2655 18192 2689 18226
rect 2655 18118 2689 18152
rect 2655 18044 2689 18078
rect 2655 17970 2689 18004
rect 2655 17896 2689 17930
rect 2655 17822 2689 17856
rect 2891 19734 2925 19768
rect 2891 19661 2925 19695
rect 2891 19588 2925 19622
rect 2891 19515 2925 19549
rect 2891 19442 2925 19476
rect 2891 19369 2925 19403
rect 2891 19296 2925 19330
rect 2891 19223 2925 19257
rect 2891 19150 2925 19184
rect 2891 19077 2925 19111
rect 2891 19004 2925 19038
rect 2891 18931 2925 18965
rect 2891 18858 2925 18892
rect 2891 18784 2925 18818
rect 2891 18710 2925 18744
rect 2891 18636 2925 18670
rect 2891 18562 2925 18596
rect 2891 18488 2925 18522
rect 2891 18414 2925 18448
rect 2891 18340 2925 18374
rect 2891 18266 2925 18300
rect 2891 18192 2925 18226
rect 2891 18118 2925 18152
rect 2891 18044 2925 18078
rect 2891 17970 2925 18004
rect 2891 17896 2925 17930
rect 2891 17822 2925 17856
rect 3036 19798 3070 19810
rect 3036 19776 3070 19798
rect 3036 19730 3070 19738
rect 3036 19704 3070 19730
rect 3036 19662 3070 19666
rect 3036 19632 3070 19662
rect 3036 19560 3070 19594
rect 3036 19492 3070 19522
rect 3036 19488 3070 19492
rect 3036 19424 3070 19450
rect 3036 19416 3070 19424
rect 3036 19356 3070 19378
rect 3036 19344 3070 19356
rect 3036 19288 3070 19306
rect 3036 19272 3070 19288
rect 3036 19220 3070 19234
rect 3036 19200 3070 19220
rect 3036 19152 3070 19162
rect 3036 19128 3070 19152
rect 3036 19084 3070 19090
rect 3036 19056 3070 19084
rect 3036 19016 3070 19018
rect 3036 18984 3070 19016
rect 3036 18914 3070 18946
rect 3036 18912 3070 18914
rect 3036 18846 3070 18874
rect 3036 18840 3070 18846
rect 3036 18778 3070 18802
rect 3036 18768 3070 18778
rect 3036 18710 3070 18730
rect 3036 18696 3070 18710
rect 3036 18642 3070 18658
rect 3036 18624 3070 18642
rect 3036 18574 3070 18586
rect 3036 18552 3070 18574
rect 3036 18506 3070 18514
rect 3036 18480 3070 18506
rect 3036 18438 3070 18442
rect 3036 18408 3070 18438
rect 3036 18336 3070 18370
rect 3036 18268 3070 18298
rect 3036 18264 3070 18268
rect 3036 18200 3070 18226
rect 3036 18192 3070 18200
rect 3036 18132 3070 18154
rect 3036 18120 3070 18132
rect 3036 18064 3070 18082
rect 3036 18048 3070 18064
rect 3036 17996 3070 18010
rect 3036 17976 3070 17996
rect 3036 17928 3070 17938
rect 3036 17904 3070 17928
rect 3036 17860 3070 17866
rect 3036 17832 3070 17860
rect 386 17771 420 17775
rect 386 17741 420 17771
rect 3036 17792 3070 17794
rect 3036 17760 3070 17792
rect 625 17720 626 17754
rect 626 17720 659 17754
rect 700 17720 732 17754
rect 732 17720 734 17754
rect 775 17720 802 17754
rect 802 17720 809 17754
rect 850 17720 872 17754
rect 872 17720 884 17754
rect 925 17720 942 17754
rect 942 17720 959 17754
rect 1000 17720 1012 17754
rect 1012 17720 1034 17754
rect 1075 17720 1082 17754
rect 1082 17720 1109 17754
rect 1150 17720 1152 17754
rect 1152 17720 1184 17754
rect 1225 17720 1256 17754
rect 1256 17720 1259 17754
rect 1300 17720 1326 17754
rect 1326 17720 1334 17754
rect 1375 17720 1396 17754
rect 1396 17720 1409 17754
rect 1450 17720 1466 17754
rect 1466 17720 1484 17754
rect 1525 17720 1536 17754
rect 1536 17720 1559 17754
rect 1600 17720 1606 17754
rect 1606 17720 1634 17754
rect 1674 17720 1676 17754
rect 1676 17720 1708 17754
rect 1748 17720 1782 17754
rect 1822 17720 1852 17754
rect 1852 17720 1856 17754
rect 1896 17720 1922 17754
rect 1922 17720 1930 17754
rect 1970 17720 1992 17754
rect 1992 17720 2004 17754
rect 2044 17720 2062 17754
rect 2062 17720 2078 17754
rect 2118 17720 2132 17754
rect 2132 17720 2152 17754
rect 2192 17720 2202 17754
rect 2202 17720 2226 17754
rect 2266 17720 2272 17754
rect 2272 17720 2300 17754
rect 2340 17720 2342 17754
rect 2342 17720 2374 17754
rect 2414 17720 2446 17754
rect 2446 17720 2448 17754
rect 2488 17720 2516 17754
rect 2516 17720 2522 17754
rect 2562 17720 2586 17754
rect 2586 17720 2596 17754
rect 2636 17720 2656 17754
rect 2656 17720 2670 17754
rect 2710 17720 2726 17754
rect 2726 17720 2744 17754
rect 2784 17720 2795 17754
rect 2795 17720 2818 17754
rect 386 17669 420 17703
rect 3036 17690 3070 17722
rect 3036 17688 3070 17690
rect 386 17601 420 17631
rect 386 17597 420 17601
rect 386 17533 420 17559
rect 386 17525 420 17533
rect 386 17465 420 17487
rect 386 17453 420 17465
rect 386 17397 420 17415
rect 386 17381 420 17397
rect 386 17329 420 17343
rect 386 17309 420 17329
rect 386 17261 420 17271
rect 386 17237 420 17261
rect 386 17193 420 17199
rect 386 17165 420 17193
rect 386 17125 420 17127
rect 386 17093 420 17125
rect 386 17023 420 17055
rect 386 17021 420 17023
rect 386 16955 420 16983
rect 386 16949 420 16955
rect 386 16887 420 16911
rect 386 16877 420 16887
rect 386 16819 420 16839
rect 386 16805 420 16819
rect 386 16751 420 16767
rect 386 16733 420 16751
rect 386 16683 420 16695
rect 386 16661 420 16683
rect 386 16615 420 16623
rect 386 16589 420 16615
rect 386 16547 420 16551
rect 386 16517 420 16547
rect 386 16445 420 16479
rect 386 16377 420 16407
rect 386 16373 420 16377
rect 386 16309 420 16335
rect 386 16301 420 16309
rect 386 16241 420 16263
rect 386 16229 420 16241
rect 386 16173 420 16191
rect 386 16157 420 16173
rect 386 16105 420 16119
rect 386 16085 420 16105
rect 386 16037 420 16047
rect 386 16013 420 16037
rect 386 15969 420 15975
rect 386 15941 420 15969
rect 386 15901 420 15903
rect 386 15869 420 15901
rect 386 15799 420 15831
rect 386 15797 420 15799
rect 386 15731 420 15759
rect 386 15725 420 15731
rect 531 17618 565 17652
rect 531 17545 565 17579
rect 531 17472 565 17506
rect 531 17399 565 17433
rect 531 17326 565 17360
rect 531 17253 565 17287
rect 531 17180 565 17214
rect 531 17107 565 17141
rect 531 17034 565 17068
rect 531 16961 565 16995
rect 531 16888 565 16922
rect 531 16815 565 16849
rect 531 16742 565 16776
rect 531 16668 565 16702
rect 531 16594 565 16628
rect 531 16520 565 16554
rect 531 16446 565 16480
rect 531 16372 565 16406
rect 531 16298 565 16332
rect 531 16224 565 16258
rect 531 16150 565 16184
rect 531 16076 565 16110
rect 531 16002 565 16036
rect 531 15928 565 15962
rect 531 15854 565 15888
rect 531 15780 565 15814
rect 531 15706 565 15740
rect 767 17618 801 17652
rect 767 17545 801 17579
rect 767 17472 801 17506
rect 767 17399 801 17433
rect 767 17326 801 17360
rect 767 17253 801 17287
rect 767 17180 801 17214
rect 767 17107 801 17141
rect 767 17034 801 17068
rect 767 16961 801 16995
rect 767 16888 801 16922
rect 767 16815 801 16849
rect 767 16742 801 16776
rect 767 16668 801 16702
rect 767 16594 801 16628
rect 767 16520 801 16554
rect 767 16446 801 16480
rect 767 16372 801 16406
rect 767 16298 801 16332
rect 767 16224 801 16258
rect 767 16150 801 16184
rect 767 16076 801 16110
rect 767 16002 801 16036
rect 767 15928 801 15962
rect 767 15854 801 15888
rect 767 15780 801 15814
rect 767 15706 801 15740
rect 1003 17618 1037 17652
rect 1003 17545 1037 17579
rect 1003 17472 1037 17506
rect 1003 17399 1037 17433
rect 1003 17326 1037 17360
rect 1003 17253 1037 17287
rect 1003 17180 1037 17214
rect 1003 17107 1037 17141
rect 1003 17034 1037 17068
rect 1003 16961 1037 16995
rect 1003 16888 1037 16922
rect 1003 16815 1037 16849
rect 1003 16742 1037 16776
rect 1003 16668 1037 16702
rect 1003 16594 1037 16628
rect 1003 16520 1037 16554
rect 1003 16446 1037 16480
rect 1003 16372 1037 16406
rect 1003 16298 1037 16332
rect 1003 16224 1037 16258
rect 1003 16150 1037 16184
rect 1003 16076 1037 16110
rect 1003 16002 1037 16036
rect 1003 15928 1037 15962
rect 1003 15854 1037 15888
rect 1003 15780 1037 15814
rect 1003 15706 1037 15740
rect 1239 17618 1273 17652
rect 1239 17545 1273 17579
rect 1239 17472 1273 17506
rect 1239 17399 1273 17433
rect 1239 17326 1273 17360
rect 1239 17253 1273 17287
rect 1239 17180 1273 17214
rect 1239 17107 1273 17141
rect 1239 17034 1273 17068
rect 1239 16961 1273 16995
rect 1239 16888 1273 16922
rect 1239 16815 1273 16849
rect 1239 16742 1273 16776
rect 1239 16668 1273 16702
rect 1239 16594 1273 16628
rect 1239 16520 1273 16554
rect 1239 16446 1273 16480
rect 1239 16372 1273 16406
rect 1239 16298 1273 16332
rect 1239 16224 1273 16258
rect 1239 16150 1273 16184
rect 1239 16076 1273 16110
rect 1239 16002 1273 16036
rect 1239 15928 1273 15962
rect 1239 15854 1273 15888
rect 1239 15780 1273 15814
rect 1239 15706 1273 15740
rect 1475 17618 1509 17652
rect 1475 17545 1509 17579
rect 1475 17472 1509 17506
rect 1475 17399 1509 17433
rect 1475 17326 1509 17360
rect 1475 17253 1509 17287
rect 1475 17180 1509 17214
rect 1475 17107 1509 17141
rect 1475 17034 1509 17068
rect 1475 16961 1509 16995
rect 1475 16888 1509 16922
rect 1475 16815 1509 16849
rect 1475 16742 1509 16776
rect 1475 16668 1509 16702
rect 1475 16594 1509 16628
rect 1475 16520 1509 16554
rect 1475 16446 1509 16480
rect 1475 16372 1509 16406
rect 1475 16298 1509 16332
rect 1475 16224 1509 16258
rect 1475 16150 1509 16184
rect 1475 16076 1509 16110
rect 1475 16002 1509 16036
rect 1475 15928 1509 15962
rect 1475 15854 1509 15888
rect 1475 15780 1509 15814
rect 1475 15706 1509 15740
rect 1711 17618 1745 17652
rect 1711 17545 1745 17579
rect 1711 17472 1745 17506
rect 1711 17399 1745 17433
rect 1711 17326 1745 17360
rect 1711 17253 1745 17287
rect 1711 17180 1745 17214
rect 1711 17107 1745 17141
rect 1711 17034 1745 17068
rect 1711 16961 1745 16995
rect 1711 16888 1745 16922
rect 1711 16815 1745 16849
rect 1711 16742 1745 16776
rect 1711 16668 1745 16702
rect 1711 16594 1745 16628
rect 1711 16520 1745 16554
rect 1711 16446 1745 16480
rect 1711 16372 1745 16406
rect 1711 16298 1745 16332
rect 1711 16224 1745 16258
rect 1711 16150 1745 16184
rect 1711 16076 1745 16110
rect 1711 16002 1745 16036
rect 1711 15928 1745 15962
rect 1711 15854 1745 15888
rect 1711 15780 1745 15814
rect 1711 15706 1745 15740
rect 1947 17618 1981 17652
rect 1947 17545 1981 17579
rect 1947 17472 1981 17506
rect 1947 17399 1981 17433
rect 1947 17326 1981 17360
rect 1947 17253 1981 17287
rect 1947 17180 1981 17214
rect 1947 17107 1981 17141
rect 1947 17034 1981 17068
rect 1947 16961 1981 16995
rect 1947 16888 1981 16922
rect 1947 16815 1981 16849
rect 1947 16742 1981 16776
rect 1947 16668 1981 16702
rect 1947 16594 1981 16628
rect 1947 16520 1981 16554
rect 1947 16446 1981 16480
rect 1947 16372 1981 16406
rect 1947 16298 1981 16332
rect 1947 16224 1981 16258
rect 1947 16150 1981 16184
rect 1947 16076 1981 16110
rect 1947 16002 1981 16036
rect 1947 15928 1981 15962
rect 1947 15854 1981 15888
rect 1947 15780 1981 15814
rect 1947 15706 1981 15740
rect 2183 17618 2217 17652
rect 2183 17545 2217 17579
rect 2183 17472 2217 17506
rect 2183 17399 2217 17433
rect 2183 17326 2217 17360
rect 2183 17253 2217 17287
rect 2183 17180 2217 17214
rect 2183 17107 2217 17141
rect 2183 17034 2217 17068
rect 2183 16961 2217 16995
rect 2183 16888 2217 16922
rect 2183 16815 2217 16849
rect 2183 16742 2217 16776
rect 2183 16668 2217 16702
rect 2183 16594 2217 16628
rect 2183 16520 2217 16554
rect 2183 16446 2217 16480
rect 2183 16372 2217 16406
rect 2183 16298 2217 16332
rect 2183 16224 2217 16258
rect 2183 16150 2217 16184
rect 2183 16076 2217 16110
rect 2183 16002 2217 16036
rect 2183 15928 2217 15962
rect 2183 15854 2217 15888
rect 2183 15780 2217 15814
rect 2183 15706 2217 15740
rect 2419 17618 2453 17652
rect 2419 17545 2453 17579
rect 2419 17472 2453 17506
rect 2419 17399 2453 17433
rect 2419 17326 2453 17360
rect 2419 17253 2453 17287
rect 2419 17180 2453 17214
rect 2419 17107 2453 17141
rect 2419 17034 2453 17068
rect 2419 16961 2453 16995
rect 2419 16888 2453 16922
rect 2419 16815 2453 16849
rect 2419 16742 2453 16776
rect 2419 16668 2453 16702
rect 2419 16594 2453 16628
rect 2419 16520 2453 16554
rect 2419 16446 2453 16480
rect 2419 16372 2453 16406
rect 2419 16298 2453 16332
rect 2419 16224 2453 16258
rect 2419 16150 2453 16184
rect 2419 16076 2453 16110
rect 2419 16002 2453 16036
rect 2419 15928 2453 15962
rect 2419 15854 2453 15888
rect 2419 15780 2453 15814
rect 2419 15706 2453 15740
rect 2655 17618 2689 17652
rect 2655 17545 2689 17579
rect 2655 17472 2689 17506
rect 2655 17399 2689 17433
rect 2655 17326 2689 17360
rect 2655 17253 2689 17287
rect 2655 17180 2689 17214
rect 2655 17107 2689 17141
rect 2655 17034 2689 17068
rect 2655 16961 2689 16995
rect 2655 16888 2689 16922
rect 2655 16815 2689 16849
rect 2655 16742 2689 16776
rect 2655 16668 2689 16702
rect 2655 16594 2689 16628
rect 2655 16520 2689 16554
rect 2655 16446 2689 16480
rect 2655 16372 2689 16406
rect 2655 16298 2689 16332
rect 2655 16224 2689 16258
rect 2655 16150 2689 16184
rect 2655 16076 2689 16110
rect 2655 16002 2689 16036
rect 2655 15928 2689 15962
rect 2655 15854 2689 15888
rect 2655 15780 2689 15814
rect 2655 15706 2689 15740
rect 2891 17618 2925 17652
rect 2891 17545 2925 17579
rect 2891 17472 2925 17506
rect 2891 17399 2925 17433
rect 2891 17326 2925 17360
rect 2891 17253 2925 17287
rect 2891 17180 2925 17214
rect 2891 17107 2925 17141
rect 2891 17034 2925 17068
rect 2891 16961 2925 16995
rect 2891 16888 2925 16922
rect 2891 16815 2925 16849
rect 2891 16742 2925 16776
rect 2891 16668 2925 16702
rect 2891 16594 2925 16628
rect 2891 16520 2925 16554
rect 2891 16446 2925 16480
rect 2891 16372 2925 16406
rect 2891 16298 2925 16332
rect 2891 16224 2925 16258
rect 2891 16150 2925 16184
rect 2891 16076 2925 16110
rect 2891 16002 2925 16036
rect 2891 15928 2925 15962
rect 2891 15854 2925 15888
rect 2891 15780 2925 15814
rect 2891 15706 2925 15740
rect 3036 17622 3070 17650
rect 3036 17616 3070 17622
rect 3036 17554 3070 17578
rect 3036 17544 3070 17554
rect 3036 17486 3070 17506
rect 3036 17472 3070 17486
rect 3036 17418 3070 17434
rect 3036 17400 3070 17418
rect 3036 17350 3070 17362
rect 3036 17328 3070 17350
rect 3036 17282 3070 17290
rect 3036 17256 3070 17282
rect 3036 17214 3070 17218
rect 3036 17184 3070 17214
rect 3036 17112 3070 17146
rect 3036 17044 3070 17074
rect 3036 17040 3070 17044
rect 3036 16976 3070 17002
rect 3036 16968 3070 16976
rect 3036 16908 3070 16930
rect 3036 16896 3070 16908
rect 3036 16840 3070 16858
rect 3036 16824 3070 16840
rect 3036 16772 3070 16786
rect 3036 16752 3070 16772
rect 3036 16704 3070 16714
rect 3036 16680 3070 16704
rect 3036 16636 3070 16642
rect 3036 16608 3070 16636
rect 3036 16568 3070 16570
rect 3036 16536 3070 16568
rect 3036 16466 3070 16498
rect 3036 16464 3070 16466
rect 3036 16398 3070 16426
rect 3036 16392 3070 16398
rect 3036 16330 3070 16354
rect 3036 16320 3070 16330
rect 3036 16262 3070 16282
rect 3036 16248 3070 16262
rect 3036 16194 3070 16210
rect 3036 16176 3070 16194
rect 3036 16126 3070 16138
rect 3036 16104 3070 16126
rect 3036 16058 3070 16066
rect 3036 16032 3070 16058
rect 3036 15990 3070 15994
rect 3036 15960 3070 15990
rect 3036 15888 3070 15922
rect 3036 15820 3070 15850
rect 3036 15816 3070 15820
rect 3036 15752 3070 15778
rect 3036 15744 3070 15752
rect 386 15663 420 15687
rect 386 15653 420 15663
rect 3036 15684 3070 15706
rect 3036 15672 3070 15684
rect 386 15595 420 15615
rect 386 15581 420 15595
rect 625 15590 626 15624
rect 626 15590 659 15624
rect 700 15590 732 15624
rect 732 15590 734 15624
rect 775 15590 802 15624
rect 802 15590 809 15624
rect 850 15590 872 15624
rect 872 15590 884 15624
rect 925 15590 942 15624
rect 942 15590 959 15624
rect 1000 15590 1012 15624
rect 1012 15590 1034 15624
rect 1075 15590 1082 15624
rect 1082 15590 1109 15624
rect 1150 15590 1152 15624
rect 1152 15590 1184 15624
rect 1225 15590 1256 15624
rect 1256 15590 1259 15624
rect 1300 15590 1326 15624
rect 1326 15590 1334 15624
rect 1375 15590 1396 15624
rect 1396 15590 1409 15624
rect 1450 15590 1466 15624
rect 1466 15590 1484 15624
rect 1525 15590 1536 15624
rect 1536 15590 1559 15624
rect 1600 15590 1606 15624
rect 1606 15590 1634 15624
rect 1674 15590 1676 15624
rect 1676 15590 1708 15624
rect 1748 15590 1782 15624
rect 1822 15590 1852 15624
rect 1852 15590 1856 15624
rect 1896 15590 1922 15624
rect 1922 15590 1930 15624
rect 1970 15590 1992 15624
rect 1992 15590 2004 15624
rect 2044 15590 2062 15624
rect 2062 15590 2078 15624
rect 2118 15590 2132 15624
rect 2132 15590 2152 15624
rect 2192 15590 2202 15624
rect 2202 15590 2226 15624
rect 2266 15590 2272 15624
rect 2272 15590 2300 15624
rect 2340 15590 2342 15624
rect 2342 15590 2374 15624
rect 2414 15590 2446 15624
rect 2446 15590 2448 15624
rect 2488 15590 2516 15624
rect 2516 15590 2522 15624
rect 2562 15590 2586 15624
rect 2586 15590 2596 15624
rect 2636 15590 2656 15624
rect 2656 15590 2670 15624
rect 2710 15590 2726 15624
rect 2726 15590 2744 15624
rect 2784 15590 2795 15624
rect 2795 15590 2818 15624
rect 3036 15616 3070 15634
rect 3036 15600 3070 15616
rect 386 15527 420 15543
rect 386 15509 420 15527
rect 3036 15548 3070 15562
rect 3036 15528 3070 15548
rect 386 15459 420 15471
rect 386 15437 420 15459
rect 386 15391 420 15399
rect 386 15365 420 15391
rect 386 15323 420 15327
rect 386 15293 420 15323
rect 386 15221 420 15255
rect 386 15153 420 15183
rect 386 15149 420 15153
rect 386 15085 420 15111
rect 386 15077 420 15085
rect 386 15017 420 15039
rect 386 15005 420 15017
rect 386 14949 420 14967
rect 386 14933 420 14949
rect 386 14881 420 14895
rect 386 14861 420 14881
rect 386 14813 420 14823
rect 386 14789 420 14813
rect 386 14745 420 14751
rect 386 14717 420 14745
rect 386 14677 420 14679
rect 386 14645 420 14677
rect 386 14575 420 14607
rect 386 14573 420 14575
rect 386 14507 420 14535
rect 386 14501 420 14507
rect 386 14439 420 14463
rect 386 14429 420 14439
rect 386 14371 420 14391
rect 386 14357 420 14371
rect 386 14303 420 14319
rect 386 14285 420 14303
rect 386 14235 420 14247
rect 386 14213 420 14235
rect 386 14167 420 14175
rect 386 14141 420 14167
rect 386 14099 420 14103
rect 386 14069 420 14099
rect 386 13997 420 14031
rect 386 13929 420 13959
rect 386 13925 420 13929
rect 386 13861 420 13887
rect 386 13853 420 13861
rect 386 13793 420 13815
rect 386 13781 420 13793
rect 386 13725 420 13743
rect 386 13709 420 13725
rect 386 13657 420 13671
rect 386 13637 420 13657
rect 386 13589 420 13599
rect 386 13565 420 13589
rect 531 15474 565 15508
rect 531 15401 565 15435
rect 531 15328 565 15362
rect 531 15255 565 15289
rect 531 15182 565 15216
rect 531 15109 565 15143
rect 531 15036 565 15070
rect 531 14963 565 14997
rect 531 14890 565 14924
rect 531 14817 565 14851
rect 531 14744 565 14778
rect 531 14671 565 14705
rect 531 14598 565 14632
rect 531 14524 565 14558
rect 531 14450 565 14484
rect 531 14376 565 14410
rect 531 14302 565 14336
rect 531 14228 565 14262
rect 531 14154 565 14188
rect 531 14080 565 14114
rect 531 14006 565 14040
rect 531 13932 565 13966
rect 531 13858 565 13892
rect 531 13784 565 13818
rect 531 13710 565 13744
rect 531 13636 565 13670
rect 531 13562 565 13596
rect 767 15474 801 15508
rect 767 15401 801 15435
rect 767 15328 801 15362
rect 767 15255 801 15289
rect 767 15182 801 15216
rect 767 15109 801 15143
rect 767 15036 801 15070
rect 767 14963 801 14997
rect 767 14890 801 14924
rect 767 14817 801 14851
rect 767 14744 801 14778
rect 767 14671 801 14705
rect 767 14598 801 14632
rect 767 14524 801 14558
rect 767 14450 801 14484
rect 767 14376 801 14410
rect 767 14302 801 14336
rect 767 14228 801 14262
rect 767 14154 801 14188
rect 767 14080 801 14114
rect 767 14006 801 14040
rect 767 13932 801 13966
rect 767 13858 801 13892
rect 767 13784 801 13818
rect 767 13710 801 13744
rect 767 13636 801 13670
rect 767 13562 801 13596
rect 1003 15474 1037 15508
rect 1003 15401 1037 15435
rect 1003 15328 1037 15362
rect 1003 15255 1037 15289
rect 1003 15182 1037 15216
rect 1003 15109 1037 15143
rect 1003 15036 1037 15070
rect 1003 14963 1037 14997
rect 1003 14890 1037 14924
rect 1003 14817 1037 14851
rect 1003 14744 1037 14778
rect 1003 14671 1037 14705
rect 1003 14598 1037 14632
rect 1003 14524 1037 14558
rect 1003 14450 1037 14484
rect 1003 14376 1037 14410
rect 1003 14302 1037 14336
rect 1003 14228 1037 14262
rect 1003 14154 1037 14188
rect 1003 14080 1037 14114
rect 1003 14006 1037 14040
rect 1003 13932 1037 13966
rect 1003 13858 1037 13892
rect 1003 13784 1037 13818
rect 1003 13710 1037 13744
rect 1003 13636 1037 13670
rect 1003 13562 1037 13596
rect 1239 15474 1273 15508
rect 1239 15401 1273 15435
rect 1239 15328 1273 15362
rect 1239 15255 1273 15289
rect 1239 15182 1273 15216
rect 1239 15109 1273 15143
rect 1239 15036 1273 15070
rect 1239 14963 1273 14997
rect 1239 14890 1273 14924
rect 1239 14817 1273 14851
rect 1239 14744 1273 14778
rect 1239 14671 1273 14705
rect 1239 14598 1273 14632
rect 1239 14524 1273 14558
rect 1239 14450 1273 14484
rect 1239 14376 1273 14410
rect 1239 14302 1273 14336
rect 1239 14228 1273 14262
rect 1239 14154 1273 14188
rect 1239 14080 1273 14114
rect 1239 14006 1273 14040
rect 1239 13932 1273 13966
rect 1239 13858 1273 13892
rect 1239 13784 1273 13818
rect 1239 13710 1273 13744
rect 1239 13636 1273 13670
rect 1239 13562 1273 13596
rect 1475 15474 1509 15508
rect 1475 15401 1509 15435
rect 1475 15328 1509 15362
rect 1475 15255 1509 15289
rect 1475 15182 1509 15216
rect 1475 15109 1509 15143
rect 1475 15036 1509 15070
rect 1475 14963 1509 14997
rect 1475 14890 1509 14924
rect 1475 14817 1509 14851
rect 1475 14744 1509 14778
rect 1475 14671 1509 14705
rect 1475 14598 1509 14632
rect 1475 14524 1509 14558
rect 1475 14450 1509 14484
rect 1475 14376 1509 14410
rect 1475 14302 1509 14336
rect 1475 14228 1509 14262
rect 1475 14154 1509 14188
rect 1475 14080 1509 14114
rect 1475 14006 1509 14040
rect 1475 13932 1509 13966
rect 1475 13858 1509 13892
rect 1475 13784 1509 13818
rect 1475 13710 1509 13744
rect 1475 13636 1509 13670
rect 1475 13562 1509 13596
rect 1711 15474 1745 15508
rect 1711 15401 1745 15435
rect 1711 15328 1745 15362
rect 1711 15255 1745 15289
rect 1711 15182 1745 15216
rect 1711 15109 1745 15143
rect 1711 15036 1745 15070
rect 1711 14963 1745 14997
rect 1711 14890 1745 14924
rect 1711 14817 1745 14851
rect 1711 14744 1745 14778
rect 1711 14671 1745 14705
rect 1711 14598 1745 14632
rect 1711 14524 1745 14558
rect 1711 14450 1745 14484
rect 1711 14376 1745 14410
rect 1711 14302 1745 14336
rect 1711 14228 1745 14262
rect 1711 14154 1745 14188
rect 1711 14080 1745 14114
rect 1711 14006 1745 14040
rect 1711 13932 1745 13966
rect 1711 13858 1745 13892
rect 1711 13784 1745 13818
rect 1711 13710 1745 13744
rect 1711 13636 1745 13670
rect 1711 13562 1745 13596
rect 1947 15474 1981 15508
rect 1947 15401 1981 15435
rect 1947 15328 1981 15362
rect 1947 15255 1981 15289
rect 1947 15182 1981 15216
rect 1947 15109 1981 15143
rect 1947 15036 1981 15070
rect 1947 14963 1981 14997
rect 1947 14890 1981 14924
rect 1947 14817 1981 14851
rect 1947 14744 1981 14778
rect 1947 14671 1981 14705
rect 1947 14598 1981 14632
rect 1947 14524 1981 14558
rect 1947 14450 1981 14484
rect 1947 14376 1981 14410
rect 1947 14302 1981 14336
rect 1947 14228 1981 14262
rect 1947 14154 1981 14188
rect 1947 14080 1981 14114
rect 1947 14006 1981 14040
rect 1947 13932 1981 13966
rect 1947 13858 1981 13892
rect 1947 13784 1981 13818
rect 1947 13710 1981 13744
rect 1947 13636 1981 13670
rect 1947 13562 1981 13596
rect 2183 15474 2217 15508
rect 2183 15401 2217 15435
rect 2183 15328 2217 15362
rect 2183 15255 2217 15289
rect 2183 15182 2217 15216
rect 2183 15109 2217 15143
rect 2183 15036 2217 15070
rect 2183 14963 2217 14997
rect 2183 14890 2217 14924
rect 2183 14817 2217 14851
rect 2183 14744 2217 14778
rect 2183 14671 2217 14705
rect 2183 14598 2217 14632
rect 2183 14524 2217 14558
rect 2183 14450 2217 14484
rect 2183 14376 2217 14410
rect 2183 14302 2217 14336
rect 2183 14228 2217 14262
rect 2183 14154 2217 14188
rect 2183 14080 2217 14114
rect 2183 14006 2217 14040
rect 2183 13932 2217 13966
rect 2183 13858 2217 13892
rect 2183 13784 2217 13818
rect 2183 13710 2217 13744
rect 2183 13636 2217 13670
rect 2183 13562 2217 13596
rect 2419 15474 2453 15508
rect 2419 15401 2453 15435
rect 2419 15328 2453 15362
rect 2419 15255 2453 15289
rect 2419 15182 2453 15216
rect 2419 15109 2453 15143
rect 2419 15036 2453 15070
rect 2419 14963 2453 14997
rect 2419 14890 2453 14924
rect 2419 14817 2453 14851
rect 2419 14744 2453 14778
rect 2419 14671 2453 14705
rect 2419 14598 2453 14632
rect 2419 14524 2453 14558
rect 2419 14450 2453 14484
rect 2419 14376 2453 14410
rect 2419 14302 2453 14336
rect 2419 14228 2453 14262
rect 2419 14154 2453 14188
rect 2419 14080 2453 14114
rect 2419 14006 2453 14040
rect 2419 13932 2453 13966
rect 2419 13858 2453 13892
rect 2419 13784 2453 13818
rect 2419 13710 2453 13744
rect 2419 13636 2453 13670
rect 2419 13562 2453 13596
rect 2655 15474 2689 15508
rect 2655 15401 2689 15435
rect 2655 15328 2689 15362
rect 2655 15255 2689 15289
rect 2655 15182 2689 15216
rect 2655 15109 2689 15143
rect 2655 15036 2689 15070
rect 2655 14963 2689 14997
rect 2655 14890 2689 14924
rect 2655 14817 2689 14851
rect 2655 14744 2689 14778
rect 2655 14671 2689 14705
rect 2655 14598 2689 14632
rect 2655 14524 2689 14558
rect 2655 14450 2689 14484
rect 2655 14376 2689 14410
rect 2655 14302 2689 14336
rect 2655 14228 2689 14262
rect 2655 14154 2689 14188
rect 2655 14080 2689 14114
rect 2655 14006 2689 14040
rect 2655 13932 2689 13966
rect 2655 13858 2689 13892
rect 2655 13784 2689 13818
rect 2655 13710 2689 13744
rect 2655 13636 2689 13670
rect 2655 13562 2689 13596
rect 2891 15474 2925 15508
rect 2891 15401 2925 15435
rect 2891 15328 2925 15362
rect 2891 15255 2925 15289
rect 2891 15182 2925 15216
rect 2891 15109 2925 15143
rect 2891 15036 2925 15070
rect 2891 14963 2925 14997
rect 2891 14890 2925 14924
rect 2891 14817 2925 14851
rect 2891 14744 2925 14778
rect 2891 14671 2925 14705
rect 2891 14598 2925 14632
rect 2891 14524 2925 14558
rect 2891 14450 2925 14484
rect 2891 14376 2925 14410
rect 2891 14302 2925 14336
rect 2891 14228 2925 14262
rect 2891 14154 2925 14188
rect 2891 14080 2925 14114
rect 2891 14006 2925 14040
rect 2891 13932 2925 13966
rect 2891 13858 2925 13892
rect 2891 13784 2925 13818
rect 2891 13710 2925 13744
rect 2891 13636 2925 13670
rect 2891 13562 2925 13596
rect 3036 15480 3070 15490
rect 3036 15456 3070 15480
rect 3036 15412 3070 15418
rect 3036 15384 3070 15412
rect 3036 15344 3070 15346
rect 3036 15312 3070 15344
rect 3036 15242 3070 15274
rect 3036 15240 3070 15242
rect 3036 15174 3070 15202
rect 3036 15168 3070 15174
rect 3036 15106 3070 15130
rect 3036 15096 3070 15106
rect 3036 15038 3070 15058
rect 3036 15024 3070 15038
rect 3036 14970 3070 14986
rect 3036 14952 3070 14970
rect 3036 14902 3070 14914
rect 3036 14880 3070 14902
rect 3036 14834 3070 14842
rect 3036 14808 3070 14834
rect 3036 14766 3070 14770
rect 3036 14736 3070 14766
rect 3036 14664 3070 14698
rect 3036 14596 3070 14626
rect 3036 14592 3070 14596
rect 3036 14528 3070 14554
rect 3036 14520 3070 14528
rect 3036 14460 3070 14482
rect 3036 14448 3070 14460
rect 3036 14392 3070 14410
rect 3036 14376 3070 14392
rect 3036 14324 3070 14338
rect 3036 14304 3070 14324
rect 3036 14256 3070 14266
rect 3036 14232 3070 14256
rect 3036 14188 3070 14194
rect 3036 14160 3070 14188
rect 3036 14120 3070 14122
rect 3036 14088 3070 14120
rect 3036 14018 3070 14050
rect 3036 14016 3070 14018
rect 3036 13950 3070 13978
rect 3036 13944 3070 13950
rect 3036 13882 3070 13906
rect 3036 13872 3070 13882
rect 3036 13814 3070 13834
rect 3036 13800 3070 13814
rect 3036 13746 3070 13762
rect 3036 13728 3070 13746
rect 3036 13678 3070 13690
rect 3036 13656 3070 13678
rect 3036 13610 3070 13618
rect 3036 13584 3070 13610
rect 386 13521 420 13527
rect 386 13493 420 13521
rect 3036 13542 3070 13546
rect 3036 13512 3070 13542
rect 386 13453 420 13455
rect 386 13421 420 13453
rect 625 13460 626 13494
rect 626 13460 659 13494
rect 700 13460 732 13494
rect 732 13460 734 13494
rect 775 13460 802 13494
rect 802 13460 809 13494
rect 850 13460 872 13494
rect 872 13460 884 13494
rect 925 13460 942 13494
rect 942 13460 959 13494
rect 1000 13460 1012 13494
rect 1012 13460 1034 13494
rect 1075 13460 1082 13494
rect 1082 13460 1109 13494
rect 1150 13460 1152 13494
rect 1152 13460 1184 13494
rect 1225 13460 1256 13494
rect 1256 13460 1259 13494
rect 1300 13460 1326 13494
rect 1326 13460 1334 13494
rect 1375 13460 1396 13494
rect 1396 13460 1409 13494
rect 1450 13460 1466 13494
rect 1466 13460 1484 13494
rect 1525 13460 1536 13494
rect 1536 13460 1559 13494
rect 1600 13460 1606 13494
rect 1606 13460 1634 13494
rect 1674 13460 1676 13494
rect 1676 13460 1708 13494
rect 1748 13460 1782 13494
rect 1822 13460 1852 13494
rect 1852 13460 1856 13494
rect 1896 13460 1922 13494
rect 1922 13460 1930 13494
rect 1970 13460 1992 13494
rect 1992 13460 2004 13494
rect 2044 13460 2062 13494
rect 2062 13460 2078 13494
rect 2118 13460 2132 13494
rect 2132 13460 2152 13494
rect 2192 13460 2202 13494
rect 2202 13460 2226 13494
rect 2266 13460 2272 13494
rect 2272 13460 2300 13494
rect 2340 13460 2342 13494
rect 2342 13460 2374 13494
rect 2414 13460 2446 13494
rect 2446 13460 2448 13494
rect 2488 13460 2516 13494
rect 2516 13460 2522 13494
rect 2562 13460 2586 13494
rect 2586 13460 2596 13494
rect 2636 13460 2656 13494
rect 2656 13460 2670 13494
rect 2710 13460 2726 13494
rect 2726 13460 2744 13494
rect 2784 13460 2795 13494
rect 2795 13460 2818 13494
rect 3036 13440 3070 13474
rect 386 13351 420 13383
rect 386 13349 420 13351
rect 386 13283 420 13311
rect 386 13277 420 13283
rect 386 13215 420 13239
rect 386 13205 420 13215
rect 386 13147 420 13167
rect 386 13133 420 13147
rect 386 13079 420 13095
rect 386 13061 420 13079
rect 386 13011 420 13023
rect 386 12989 420 13011
rect 386 12943 420 12951
rect 386 12917 420 12943
rect 386 12875 420 12879
rect 386 12845 420 12875
rect 386 12773 420 12807
rect 386 12705 420 12735
rect 386 12701 420 12705
rect 386 12637 420 12663
rect 386 12629 420 12637
rect 386 12569 420 12591
rect 386 12557 420 12569
rect 386 12501 420 12519
rect 386 12485 420 12501
rect 386 12433 420 12447
rect 386 12413 420 12433
rect 386 12365 420 12375
rect 386 12341 420 12365
rect 386 12297 420 12303
rect 386 12269 420 12297
rect 386 12229 420 12231
rect 386 12197 420 12229
rect 386 12127 420 12159
rect 386 12125 420 12127
rect 386 12059 420 12087
rect 386 12053 420 12059
rect 386 11991 420 12015
rect 386 11981 420 11991
rect 386 11923 420 11943
rect 386 11909 420 11923
rect 386 11855 420 11871
rect 386 11837 420 11855
rect 386 11787 420 11799
rect 386 11765 420 11787
rect 386 11719 420 11727
rect 386 11693 420 11719
rect 386 11651 420 11655
rect 386 11621 420 11651
rect 386 11549 420 11583
rect 386 11481 420 11511
rect 386 11477 420 11481
rect 386 11413 420 11439
rect 386 11405 420 11413
rect 531 13358 565 13392
rect 531 13285 565 13319
rect 531 13212 565 13246
rect 531 13139 565 13173
rect 531 13066 565 13100
rect 531 12993 565 13027
rect 531 12920 565 12954
rect 531 12847 565 12881
rect 531 12774 565 12808
rect 531 12701 565 12735
rect 531 12628 565 12662
rect 531 12555 565 12589
rect 531 12482 565 12516
rect 531 12408 565 12442
rect 531 12334 565 12368
rect 531 12260 565 12294
rect 531 12186 565 12220
rect 531 12112 565 12146
rect 531 12038 565 12072
rect 531 11964 565 11998
rect 531 11890 565 11924
rect 531 11816 565 11850
rect 531 11742 565 11776
rect 531 11668 565 11702
rect 531 11594 565 11628
rect 531 11520 565 11554
rect 531 11446 565 11480
rect 767 13358 801 13392
rect 767 13285 801 13319
rect 767 13212 801 13246
rect 767 13139 801 13173
rect 767 13066 801 13100
rect 767 12993 801 13027
rect 767 12920 801 12954
rect 767 12847 801 12881
rect 767 12774 801 12808
rect 767 12701 801 12735
rect 767 12628 801 12662
rect 767 12555 801 12589
rect 767 12482 801 12516
rect 767 12408 801 12442
rect 767 12334 801 12368
rect 767 12260 801 12294
rect 767 12186 801 12220
rect 767 12112 801 12146
rect 767 12038 801 12072
rect 767 11964 801 11998
rect 767 11890 801 11924
rect 767 11816 801 11850
rect 767 11742 801 11776
rect 767 11668 801 11702
rect 767 11594 801 11628
rect 767 11520 801 11554
rect 767 11446 801 11480
rect 1003 13358 1037 13392
rect 1003 13285 1037 13319
rect 1003 13212 1037 13246
rect 1003 13139 1037 13173
rect 1003 13066 1037 13100
rect 1003 12993 1037 13027
rect 1003 12920 1037 12954
rect 1003 12847 1037 12881
rect 1003 12774 1037 12808
rect 1003 12701 1037 12735
rect 1003 12628 1037 12662
rect 1003 12555 1037 12589
rect 1003 12482 1037 12516
rect 1003 12408 1037 12442
rect 1003 12334 1037 12368
rect 1003 12260 1037 12294
rect 1003 12186 1037 12220
rect 1003 12112 1037 12146
rect 1003 12038 1037 12072
rect 1003 11964 1037 11998
rect 1003 11890 1037 11924
rect 1003 11816 1037 11850
rect 1003 11742 1037 11776
rect 1003 11668 1037 11702
rect 1003 11594 1037 11628
rect 1003 11520 1037 11554
rect 1003 11446 1037 11480
rect 1239 13358 1273 13392
rect 1239 13285 1273 13319
rect 1239 13212 1273 13246
rect 1239 13139 1273 13173
rect 1239 13066 1273 13100
rect 1239 12993 1273 13027
rect 1239 12920 1273 12954
rect 1239 12847 1273 12881
rect 1239 12774 1273 12808
rect 1239 12701 1273 12735
rect 1239 12628 1273 12662
rect 1239 12555 1273 12589
rect 1239 12482 1273 12516
rect 1239 12408 1273 12442
rect 1239 12334 1273 12368
rect 1239 12260 1273 12294
rect 1239 12186 1273 12220
rect 1239 12112 1273 12146
rect 1239 12038 1273 12072
rect 1239 11964 1273 11998
rect 1239 11890 1273 11924
rect 1239 11816 1273 11850
rect 1239 11742 1273 11776
rect 1239 11668 1273 11702
rect 1239 11594 1273 11628
rect 1239 11520 1273 11554
rect 1239 11446 1273 11480
rect 1475 13358 1509 13392
rect 1475 13285 1509 13319
rect 1475 13212 1509 13246
rect 1475 13139 1509 13173
rect 1475 13066 1509 13100
rect 1475 12993 1509 13027
rect 1475 12920 1509 12954
rect 1475 12847 1509 12881
rect 1475 12774 1509 12808
rect 1475 12701 1509 12735
rect 1475 12628 1509 12662
rect 1475 12555 1509 12589
rect 1475 12482 1509 12516
rect 1475 12408 1509 12442
rect 1475 12334 1509 12368
rect 1475 12260 1509 12294
rect 1475 12186 1509 12220
rect 1475 12112 1509 12146
rect 1475 12038 1509 12072
rect 1475 11964 1509 11998
rect 1475 11890 1509 11924
rect 1475 11816 1509 11850
rect 1475 11742 1509 11776
rect 1475 11668 1509 11702
rect 1475 11594 1509 11628
rect 1475 11520 1509 11554
rect 1475 11446 1509 11480
rect 1711 13358 1745 13392
rect 1711 13285 1745 13319
rect 1711 13212 1745 13246
rect 1711 13139 1745 13173
rect 1711 13066 1745 13100
rect 1711 12993 1745 13027
rect 1711 12920 1745 12954
rect 1711 12847 1745 12881
rect 1711 12774 1745 12808
rect 1711 12701 1745 12735
rect 1711 12628 1745 12662
rect 1711 12555 1745 12589
rect 1711 12482 1745 12516
rect 1711 12408 1745 12442
rect 1711 12334 1745 12368
rect 1711 12260 1745 12294
rect 1711 12186 1745 12220
rect 1711 12112 1745 12146
rect 1711 12038 1745 12072
rect 1711 11964 1745 11998
rect 1711 11890 1745 11924
rect 1711 11816 1745 11850
rect 1711 11742 1745 11776
rect 1711 11668 1745 11702
rect 1711 11594 1745 11628
rect 1711 11520 1745 11554
rect 1711 11446 1745 11480
rect 1947 13358 1981 13392
rect 1947 13285 1981 13319
rect 1947 13212 1981 13246
rect 1947 13139 1981 13173
rect 1947 13066 1981 13100
rect 1947 12993 1981 13027
rect 1947 12920 1981 12954
rect 1947 12847 1981 12881
rect 1947 12774 1981 12808
rect 1947 12701 1981 12735
rect 1947 12628 1981 12662
rect 1947 12555 1981 12589
rect 1947 12482 1981 12516
rect 1947 12408 1981 12442
rect 1947 12334 1981 12368
rect 1947 12260 1981 12294
rect 1947 12186 1981 12220
rect 1947 12112 1981 12146
rect 1947 12038 1981 12072
rect 1947 11964 1981 11998
rect 1947 11890 1981 11924
rect 1947 11816 1981 11850
rect 1947 11742 1981 11776
rect 1947 11668 1981 11702
rect 1947 11594 1981 11628
rect 1947 11520 1981 11554
rect 1947 11446 1981 11480
rect 2183 13358 2217 13392
rect 2183 13285 2217 13319
rect 2183 13212 2217 13246
rect 2183 13139 2217 13173
rect 2183 13066 2217 13100
rect 2183 12993 2217 13027
rect 2183 12920 2217 12954
rect 2183 12847 2217 12881
rect 2183 12774 2217 12808
rect 2183 12701 2217 12735
rect 2183 12628 2217 12662
rect 2183 12555 2217 12589
rect 2183 12482 2217 12516
rect 2183 12408 2217 12442
rect 2183 12334 2217 12368
rect 2183 12260 2217 12294
rect 2183 12186 2217 12220
rect 2183 12112 2217 12146
rect 2183 12038 2217 12072
rect 2183 11964 2217 11998
rect 2183 11890 2217 11924
rect 2183 11816 2217 11850
rect 2183 11742 2217 11776
rect 2183 11668 2217 11702
rect 2183 11594 2217 11628
rect 2183 11520 2217 11554
rect 2183 11446 2217 11480
rect 2419 13358 2453 13392
rect 2419 13285 2453 13319
rect 2419 13212 2453 13246
rect 2419 13139 2453 13173
rect 2419 13066 2453 13100
rect 2419 12993 2453 13027
rect 2419 12920 2453 12954
rect 2419 12847 2453 12881
rect 2419 12774 2453 12808
rect 2419 12701 2453 12735
rect 2419 12628 2453 12662
rect 2419 12555 2453 12589
rect 2419 12482 2453 12516
rect 2419 12408 2453 12442
rect 2419 12334 2453 12368
rect 2419 12260 2453 12294
rect 2419 12186 2453 12220
rect 2419 12112 2453 12146
rect 2419 12038 2453 12072
rect 2419 11964 2453 11998
rect 2419 11890 2453 11924
rect 2419 11816 2453 11850
rect 2419 11742 2453 11776
rect 2419 11668 2453 11702
rect 2419 11594 2453 11628
rect 2419 11520 2453 11554
rect 2419 11446 2453 11480
rect 2655 13358 2689 13392
rect 2655 13285 2689 13319
rect 2655 13212 2689 13246
rect 2655 13139 2689 13173
rect 2655 13066 2689 13100
rect 2655 12993 2689 13027
rect 2655 12920 2689 12954
rect 2655 12847 2689 12881
rect 2655 12774 2689 12808
rect 2655 12701 2689 12735
rect 2655 12628 2689 12662
rect 2655 12555 2689 12589
rect 2655 12482 2689 12516
rect 2655 12408 2689 12442
rect 2655 12334 2689 12368
rect 2655 12260 2689 12294
rect 2655 12186 2689 12220
rect 2655 12112 2689 12146
rect 2655 12038 2689 12072
rect 2655 11964 2689 11998
rect 2655 11890 2689 11924
rect 2655 11816 2689 11850
rect 2655 11742 2689 11776
rect 2655 11668 2689 11702
rect 2655 11594 2689 11628
rect 2655 11520 2689 11554
rect 2655 11446 2689 11480
rect 2891 13358 2925 13392
rect 2891 13285 2925 13319
rect 2891 13212 2925 13246
rect 2891 13139 2925 13173
rect 2891 13066 2925 13100
rect 2891 12993 2925 13027
rect 2891 12920 2925 12954
rect 2891 12847 2925 12881
rect 2891 12774 2925 12808
rect 2891 12701 2925 12735
rect 2891 12628 2925 12662
rect 2891 12555 2925 12589
rect 2891 12482 2925 12516
rect 2891 12408 2925 12442
rect 2891 12334 2925 12368
rect 2891 12260 2925 12294
rect 2891 12186 2925 12220
rect 2891 12112 2925 12146
rect 2891 12038 2925 12072
rect 2891 11964 2925 11998
rect 2891 11890 2925 11924
rect 2891 11816 2925 11850
rect 2891 11742 2925 11776
rect 2891 11668 2925 11702
rect 2891 11594 2925 11628
rect 2891 11520 2925 11554
rect 2891 11446 2925 11480
rect 3036 13372 3070 13402
rect 3036 13368 3070 13372
rect 3036 13304 3070 13330
rect 3036 13296 3070 13304
rect 3036 13236 3070 13258
rect 3036 13224 3070 13236
rect 3036 13168 3070 13186
rect 3036 13152 3070 13168
rect 3036 13100 3070 13114
rect 3036 13080 3070 13100
rect 3036 13032 3070 13042
rect 3036 13008 3070 13032
rect 3036 12964 3070 12970
rect 3036 12936 3070 12964
rect 3036 12896 3070 12898
rect 3036 12864 3070 12896
rect 3036 12794 3070 12826
rect 3036 12792 3070 12794
rect 3036 12726 3070 12754
rect 3036 12720 3070 12726
rect 3036 12658 3070 12682
rect 3036 12648 3070 12658
rect 3036 12590 3070 12610
rect 3036 12576 3070 12590
rect 3036 12522 3070 12538
rect 3036 12504 3070 12522
rect 3036 12454 3070 12466
rect 3036 12432 3070 12454
rect 3036 12386 3070 12394
rect 3036 12360 3070 12386
rect 3036 12318 3070 12322
rect 3036 12288 3070 12318
rect 3036 12216 3070 12250
rect 3036 12148 3070 12178
rect 3036 12144 3070 12148
rect 3036 12080 3070 12106
rect 3036 12072 3070 12080
rect 3036 12012 3070 12034
rect 3036 12000 3070 12012
rect 3036 11944 3070 11962
rect 3036 11928 3070 11944
rect 3036 11876 3070 11890
rect 3036 11856 3070 11876
rect 3036 11808 3070 11818
rect 3036 11784 3070 11808
rect 3036 11740 3070 11746
rect 3036 11712 3070 11740
rect 3036 11672 3070 11674
rect 3036 11640 3070 11672
rect 3036 11570 3070 11602
rect 3036 11568 3070 11570
rect 3036 11502 3070 11530
rect 3036 11496 3070 11502
rect 386 11345 420 11367
rect 386 11333 420 11345
rect 3036 11434 3070 11458
rect 3036 11424 3070 11434
rect 625 11330 626 11364
rect 626 11330 659 11364
rect 700 11330 732 11364
rect 732 11330 734 11364
rect 775 11330 802 11364
rect 802 11330 809 11364
rect 850 11330 872 11364
rect 872 11330 884 11364
rect 925 11330 942 11364
rect 942 11330 959 11364
rect 1000 11330 1012 11364
rect 1012 11330 1034 11364
rect 1075 11330 1082 11364
rect 1082 11330 1109 11364
rect 1150 11330 1152 11364
rect 1152 11330 1184 11364
rect 1225 11330 1256 11364
rect 1256 11330 1259 11364
rect 1300 11330 1326 11364
rect 1326 11330 1334 11364
rect 1375 11330 1396 11364
rect 1396 11330 1409 11364
rect 1450 11330 1466 11364
rect 1466 11330 1484 11364
rect 1525 11330 1536 11364
rect 1536 11330 1559 11364
rect 1600 11330 1606 11364
rect 1606 11330 1634 11364
rect 1674 11330 1676 11364
rect 1676 11330 1708 11364
rect 1748 11330 1782 11364
rect 1822 11330 1852 11364
rect 1852 11330 1856 11364
rect 1896 11330 1922 11364
rect 1922 11330 1930 11364
rect 1970 11330 1992 11364
rect 1992 11330 2004 11364
rect 2044 11330 2062 11364
rect 2062 11330 2078 11364
rect 2118 11330 2132 11364
rect 2132 11330 2152 11364
rect 2192 11330 2202 11364
rect 2202 11330 2226 11364
rect 2266 11330 2272 11364
rect 2272 11330 2300 11364
rect 2340 11330 2342 11364
rect 2342 11330 2374 11364
rect 2414 11330 2446 11364
rect 2446 11330 2448 11364
rect 2488 11330 2516 11364
rect 2516 11330 2522 11364
rect 2562 11330 2586 11364
rect 2586 11330 2596 11364
rect 2636 11330 2656 11364
rect 2656 11330 2670 11364
rect 2710 11330 2726 11364
rect 2726 11330 2744 11364
rect 2784 11330 2795 11364
rect 2795 11330 2818 11364
rect 3036 11366 3070 11386
rect 3036 11352 3070 11366
rect 386 11277 420 11295
rect 386 11261 420 11277
rect 3036 11298 3070 11314
rect 3036 11280 3070 11298
rect 386 11209 420 11223
rect 386 11189 420 11209
rect 386 11141 420 11151
rect 386 11117 420 11141
rect 386 11073 420 11079
rect 386 11045 420 11073
rect 386 11005 420 11007
rect 386 10973 420 11005
rect 386 10903 420 10935
rect 386 10901 420 10903
rect 386 10835 420 10863
rect 386 10829 420 10835
rect 386 10767 420 10791
rect 386 10757 420 10767
rect 386 10699 420 10719
rect 386 10685 420 10699
rect 386 10631 420 10647
rect 386 10613 420 10631
rect 386 10563 420 10575
rect 386 10541 420 10563
rect 386 10495 420 10503
rect 386 10469 420 10495
rect 386 10427 420 10431
rect 386 10397 420 10427
rect 386 10325 420 10359
rect 386 10257 420 10287
rect 386 10253 420 10257
rect 386 10189 420 10215
rect 386 10181 420 10189
rect 386 10121 420 10143
rect 386 10109 420 10121
rect 386 10053 420 10071
rect 386 10037 420 10053
rect 386 9985 420 9999
rect 386 9965 420 9985
rect 386 9917 420 9927
rect 386 9893 420 9917
rect 386 9849 420 9855
rect 386 9821 420 9849
rect 386 9781 420 9783
rect 386 9749 420 9781
rect 386 9679 420 9711
rect 386 9677 420 9679
rect 386 9611 420 9639
rect 386 9605 420 9611
rect 386 9543 420 9567
rect 386 9533 420 9543
rect 386 9475 420 9495
rect 386 9461 420 9475
rect 386 9407 420 9423
rect 386 9389 420 9407
rect 386 9339 420 9351
rect 386 9317 420 9339
rect 531 11214 565 11248
rect 531 11141 565 11175
rect 531 11068 565 11102
rect 531 10995 565 11029
rect 531 10922 565 10956
rect 531 10849 565 10883
rect 531 10776 565 10810
rect 531 10703 565 10737
rect 531 10630 565 10664
rect 531 10557 565 10591
rect 531 10484 565 10518
rect 531 10411 565 10445
rect 531 10338 565 10372
rect 531 10264 565 10298
rect 531 10190 565 10224
rect 531 10116 565 10150
rect 531 10042 565 10076
rect 531 9968 565 10002
rect 531 9894 565 9928
rect 531 9820 565 9854
rect 531 9746 565 9780
rect 531 9672 565 9706
rect 531 9598 565 9632
rect 531 9524 565 9558
rect 531 9450 565 9484
rect 531 9376 565 9410
rect 531 9302 565 9336
rect 767 11214 801 11248
rect 767 11141 801 11175
rect 767 11068 801 11102
rect 767 10995 801 11029
rect 767 10922 801 10956
rect 767 10849 801 10883
rect 767 10776 801 10810
rect 767 10703 801 10737
rect 767 10630 801 10664
rect 767 10557 801 10591
rect 767 10484 801 10518
rect 767 10411 801 10445
rect 767 10338 801 10372
rect 767 10264 801 10298
rect 767 10190 801 10224
rect 767 10116 801 10150
rect 767 10042 801 10076
rect 767 9968 801 10002
rect 767 9894 801 9928
rect 767 9820 801 9854
rect 767 9746 801 9780
rect 767 9672 801 9706
rect 767 9598 801 9632
rect 767 9524 801 9558
rect 767 9450 801 9484
rect 767 9376 801 9410
rect 767 9302 801 9336
rect 1003 11214 1037 11248
rect 1003 11141 1037 11175
rect 1003 11068 1037 11102
rect 1003 10995 1037 11029
rect 1003 10922 1037 10956
rect 1003 10849 1037 10883
rect 1003 10776 1037 10810
rect 1003 10703 1037 10737
rect 1003 10630 1037 10664
rect 1003 10557 1037 10591
rect 1003 10484 1037 10518
rect 1003 10411 1037 10445
rect 1003 10338 1037 10372
rect 1003 10264 1037 10298
rect 1003 10190 1037 10224
rect 1003 10116 1037 10150
rect 1003 10042 1037 10076
rect 1003 9968 1037 10002
rect 1003 9894 1037 9928
rect 1003 9820 1037 9854
rect 1003 9746 1037 9780
rect 1003 9672 1037 9706
rect 1003 9598 1037 9632
rect 1003 9524 1037 9558
rect 1003 9450 1037 9484
rect 1003 9376 1037 9410
rect 1003 9302 1037 9336
rect 1239 11214 1273 11248
rect 1239 11141 1273 11175
rect 1239 11068 1273 11102
rect 1239 10995 1273 11029
rect 1239 10922 1273 10956
rect 1239 10849 1273 10883
rect 1239 10776 1273 10810
rect 1239 10703 1273 10737
rect 1239 10630 1273 10664
rect 1239 10557 1273 10591
rect 1239 10484 1273 10518
rect 1239 10411 1273 10445
rect 1239 10338 1273 10372
rect 1239 10264 1273 10298
rect 1239 10190 1273 10224
rect 1239 10116 1273 10150
rect 1239 10042 1273 10076
rect 1239 9968 1273 10002
rect 1239 9894 1273 9928
rect 1239 9820 1273 9854
rect 1239 9746 1273 9780
rect 1239 9672 1273 9706
rect 1239 9598 1273 9632
rect 1239 9524 1273 9558
rect 1239 9450 1273 9484
rect 1239 9376 1273 9410
rect 1239 9302 1273 9336
rect 1475 11214 1509 11248
rect 1475 11141 1509 11175
rect 1475 11068 1509 11102
rect 1475 10995 1509 11029
rect 1475 10922 1509 10956
rect 1475 10849 1509 10883
rect 1475 10776 1509 10810
rect 1475 10703 1509 10737
rect 1475 10630 1509 10664
rect 1475 10557 1509 10591
rect 1475 10484 1509 10518
rect 1475 10411 1509 10445
rect 1475 10338 1509 10372
rect 1475 10264 1509 10298
rect 1475 10190 1509 10224
rect 1475 10116 1509 10150
rect 1475 10042 1509 10076
rect 1475 9968 1509 10002
rect 1475 9894 1509 9928
rect 1475 9820 1509 9854
rect 1475 9746 1509 9780
rect 1475 9672 1509 9706
rect 1475 9598 1509 9632
rect 1475 9524 1509 9558
rect 1475 9450 1509 9484
rect 1475 9376 1509 9410
rect 1475 9302 1509 9336
rect 1711 11214 1745 11248
rect 1711 11141 1745 11175
rect 1711 11068 1745 11102
rect 1711 10995 1745 11029
rect 1711 10922 1745 10956
rect 1711 10849 1745 10883
rect 1711 10776 1745 10810
rect 1711 10703 1745 10737
rect 1711 10630 1745 10664
rect 1711 10557 1745 10591
rect 1711 10484 1745 10518
rect 1711 10411 1745 10445
rect 1711 10338 1745 10372
rect 1711 10264 1745 10298
rect 1711 10190 1745 10224
rect 1711 10116 1745 10150
rect 1711 10042 1745 10076
rect 1711 9968 1745 10002
rect 1711 9894 1745 9928
rect 1711 9820 1745 9854
rect 1711 9746 1745 9780
rect 1711 9672 1745 9706
rect 1711 9598 1745 9632
rect 1711 9524 1745 9558
rect 1711 9450 1745 9484
rect 1711 9376 1745 9410
rect 1711 9302 1745 9336
rect 1947 11214 1981 11248
rect 1947 11141 1981 11175
rect 1947 11068 1981 11102
rect 1947 10995 1981 11029
rect 1947 10922 1981 10956
rect 1947 10849 1981 10883
rect 1947 10776 1981 10810
rect 1947 10703 1981 10737
rect 1947 10630 1981 10664
rect 1947 10557 1981 10591
rect 1947 10484 1981 10518
rect 1947 10411 1981 10445
rect 1947 10338 1981 10372
rect 1947 10264 1981 10298
rect 1947 10190 1981 10224
rect 1947 10116 1981 10150
rect 1947 10042 1981 10076
rect 1947 9968 1981 10002
rect 1947 9894 1981 9928
rect 1947 9820 1981 9854
rect 1947 9746 1981 9780
rect 1947 9672 1981 9706
rect 1947 9598 1981 9632
rect 1947 9524 1981 9558
rect 1947 9450 1981 9484
rect 1947 9376 1981 9410
rect 1947 9302 1981 9336
rect 2183 11214 2217 11248
rect 2183 11141 2217 11175
rect 2183 11068 2217 11102
rect 2183 10995 2217 11029
rect 2183 10922 2217 10956
rect 2183 10849 2217 10883
rect 2183 10776 2217 10810
rect 2183 10703 2217 10737
rect 2183 10630 2217 10664
rect 2183 10557 2217 10591
rect 2183 10484 2217 10518
rect 2183 10411 2217 10445
rect 2183 10338 2217 10372
rect 2183 10264 2217 10298
rect 2183 10190 2217 10224
rect 2183 10116 2217 10150
rect 2183 10042 2217 10076
rect 2183 9968 2217 10002
rect 2183 9894 2217 9928
rect 2183 9820 2217 9854
rect 2183 9746 2217 9780
rect 2183 9672 2217 9706
rect 2183 9598 2217 9632
rect 2183 9524 2217 9558
rect 2183 9450 2217 9484
rect 2183 9376 2217 9410
rect 2183 9302 2217 9336
rect 2419 11214 2453 11248
rect 2419 11141 2453 11175
rect 2419 11068 2453 11102
rect 2419 10995 2453 11029
rect 2419 10922 2453 10956
rect 2419 10849 2453 10883
rect 2419 10776 2453 10810
rect 2419 10703 2453 10737
rect 2419 10630 2453 10664
rect 2419 10557 2453 10591
rect 2419 10484 2453 10518
rect 2419 10411 2453 10445
rect 2419 10338 2453 10372
rect 2419 10264 2453 10298
rect 2419 10190 2453 10224
rect 2419 10116 2453 10150
rect 2419 10042 2453 10076
rect 2419 9968 2453 10002
rect 2419 9894 2453 9928
rect 2419 9820 2453 9854
rect 2419 9746 2453 9780
rect 2419 9672 2453 9706
rect 2419 9598 2453 9632
rect 2419 9524 2453 9558
rect 2419 9450 2453 9484
rect 2419 9376 2453 9410
rect 2419 9302 2453 9336
rect 2655 11214 2689 11248
rect 2655 11141 2689 11175
rect 2655 11068 2689 11102
rect 2655 10995 2689 11029
rect 2655 10922 2689 10956
rect 2655 10849 2689 10883
rect 2655 10776 2689 10810
rect 2655 10703 2689 10737
rect 2655 10630 2689 10664
rect 2655 10557 2689 10591
rect 2655 10484 2689 10518
rect 2655 10411 2689 10445
rect 2655 10338 2689 10372
rect 2655 10264 2689 10298
rect 2655 10190 2689 10224
rect 2655 10116 2689 10150
rect 2655 10042 2689 10076
rect 2655 9968 2689 10002
rect 2655 9894 2689 9928
rect 2655 9820 2689 9854
rect 2655 9746 2689 9780
rect 2655 9672 2689 9706
rect 2655 9598 2689 9632
rect 2655 9524 2689 9558
rect 2655 9450 2689 9484
rect 2655 9376 2689 9410
rect 2655 9302 2689 9336
rect 2891 11214 2925 11248
rect 2891 11141 2925 11175
rect 2891 11068 2925 11102
rect 2891 10995 2925 11029
rect 2891 10922 2925 10956
rect 2891 10849 2925 10883
rect 2891 10776 2925 10810
rect 2891 10703 2925 10737
rect 2891 10630 2925 10664
rect 2891 10557 2925 10591
rect 2891 10484 2925 10518
rect 2891 10411 2925 10445
rect 2891 10338 2925 10372
rect 2891 10264 2925 10298
rect 2891 10190 2925 10224
rect 2891 10116 2925 10150
rect 2891 10042 2925 10076
rect 2891 9968 2925 10002
rect 2891 9894 2925 9928
rect 2891 9820 2925 9854
rect 2891 9746 2925 9780
rect 2891 9672 2925 9706
rect 2891 9598 2925 9632
rect 2891 9524 2925 9558
rect 2891 9450 2925 9484
rect 2891 9376 2925 9410
rect 2891 9302 2925 9336
rect 3036 11230 3070 11242
rect 3036 11208 3070 11230
rect 3036 11162 3070 11170
rect 3036 11136 3070 11162
rect 3036 11094 3070 11098
rect 3036 11064 3070 11094
rect 3036 10992 3070 11026
rect 3036 10924 3070 10954
rect 3036 10920 3070 10924
rect 3036 10856 3070 10882
rect 3036 10848 3070 10856
rect 3036 10788 3070 10810
rect 3036 10776 3070 10788
rect 3036 10720 3070 10738
rect 3036 10704 3070 10720
rect 3036 10652 3070 10666
rect 3036 10632 3070 10652
rect 3036 10584 3070 10594
rect 3036 10560 3070 10584
rect 3036 10516 3070 10522
rect 3036 10488 3070 10516
rect 3036 10448 3070 10450
rect 3036 10416 3070 10448
rect 3036 10346 3070 10378
rect 3036 10344 3070 10346
rect 3036 10278 3070 10306
rect 3036 10272 3070 10278
rect 3036 10210 3070 10234
rect 3036 10200 3070 10210
rect 3036 10142 3070 10162
rect 3036 10128 3070 10142
rect 3036 10074 3070 10090
rect 3036 10056 3070 10074
rect 3036 10006 3070 10018
rect 3036 9984 3070 10006
rect 3036 9938 3070 9946
rect 3036 9912 3070 9938
rect 3036 9870 3070 9874
rect 3036 9840 3070 9870
rect 3036 9768 3070 9802
rect 3036 9700 3070 9730
rect 3036 9696 3070 9700
rect 3036 9632 3070 9658
rect 3036 9624 3070 9632
rect 3036 9564 3070 9586
rect 3036 9552 3070 9564
rect 3036 9496 3070 9514
rect 3036 9480 3070 9496
rect 3036 9428 3070 9442
rect 3036 9408 3070 9428
rect 3036 9360 3070 9370
rect 3036 9336 3070 9360
rect 386 9271 420 9279
rect 386 9245 420 9271
rect 3036 9292 3070 9298
rect 3036 9264 3070 9292
rect 386 9203 420 9207
rect 386 9173 420 9203
rect 625 9200 626 9234
rect 626 9200 659 9234
rect 700 9200 732 9234
rect 732 9200 734 9234
rect 775 9200 802 9234
rect 802 9200 809 9234
rect 850 9200 872 9234
rect 872 9200 884 9234
rect 925 9200 942 9234
rect 942 9200 959 9234
rect 1000 9200 1012 9234
rect 1012 9200 1034 9234
rect 1075 9200 1082 9234
rect 1082 9200 1109 9234
rect 1150 9200 1152 9234
rect 1152 9200 1184 9234
rect 1225 9200 1256 9234
rect 1256 9200 1259 9234
rect 1300 9200 1326 9234
rect 1326 9200 1334 9234
rect 1375 9200 1396 9234
rect 1396 9200 1409 9234
rect 1450 9200 1466 9234
rect 1466 9200 1484 9234
rect 1525 9200 1536 9234
rect 1536 9200 1559 9234
rect 1600 9200 1606 9234
rect 1606 9200 1634 9234
rect 1674 9200 1676 9234
rect 1676 9200 1708 9234
rect 1748 9200 1782 9234
rect 1822 9200 1852 9234
rect 1852 9200 1856 9234
rect 1896 9200 1922 9234
rect 1922 9200 1930 9234
rect 1970 9200 1992 9234
rect 1992 9200 2004 9234
rect 2044 9200 2062 9234
rect 2062 9200 2078 9234
rect 2118 9200 2132 9234
rect 2132 9200 2152 9234
rect 2192 9200 2202 9234
rect 2202 9200 2226 9234
rect 2266 9200 2272 9234
rect 2272 9200 2300 9234
rect 2340 9200 2342 9234
rect 2342 9200 2374 9234
rect 2414 9200 2446 9234
rect 2446 9200 2448 9234
rect 2488 9200 2516 9234
rect 2516 9200 2522 9234
rect 2562 9200 2586 9234
rect 2586 9200 2596 9234
rect 2636 9200 2656 9234
rect 2656 9200 2670 9234
rect 2710 9200 2726 9234
rect 2726 9200 2744 9234
rect 2784 9200 2795 9234
rect 2795 9200 2818 9234
rect 386 9101 420 9135
rect 3036 9224 3070 9226
rect 3036 9192 3070 9224
rect 386 9033 420 9063
rect 386 9029 420 9033
rect 386 8965 420 8991
rect 386 8957 420 8965
rect 386 8897 420 8919
rect 386 8885 420 8897
rect 386 8829 420 8847
rect 386 8813 420 8829
rect 386 8761 420 8775
rect 386 8741 420 8761
rect 386 8693 420 8703
rect 386 8669 420 8693
rect 386 8625 420 8631
rect 386 8597 420 8625
rect 386 8557 420 8559
rect 386 8525 420 8557
rect 386 8455 420 8487
rect 386 8453 420 8455
rect 386 8387 420 8415
rect 386 8381 420 8387
rect 386 8319 420 8343
rect 386 8309 420 8319
rect 386 8251 420 8271
rect 386 8237 420 8251
rect 386 8183 420 8199
rect 386 8165 420 8183
rect 386 8115 420 8127
rect 386 8093 420 8115
rect 386 8047 420 8055
rect 386 8021 420 8047
rect 386 7979 420 7983
rect 386 7949 420 7979
rect 386 7877 420 7911
rect 386 7809 420 7839
rect 386 7805 420 7809
rect 386 7741 420 7767
rect 386 7733 420 7741
rect 386 7673 420 7695
rect 386 7661 420 7673
rect 386 7605 420 7623
rect 386 7589 420 7605
rect 386 7537 420 7551
rect 386 7517 420 7537
rect 386 7469 420 7479
rect 386 7445 420 7469
rect 386 7401 420 7407
rect 386 7373 420 7401
rect 386 7333 420 7335
rect 386 7301 420 7333
rect 386 7231 420 7263
rect 386 7229 420 7231
rect 386 7163 420 7191
rect 386 7157 420 7163
rect 531 9098 565 9132
rect 531 9025 565 9059
rect 531 8952 565 8986
rect 531 8879 565 8913
rect 531 8806 565 8840
rect 531 8733 565 8767
rect 531 8660 565 8694
rect 531 8587 565 8621
rect 531 8514 565 8548
rect 531 8441 565 8475
rect 531 8368 565 8402
rect 531 8295 565 8329
rect 531 8222 565 8256
rect 531 8148 565 8182
rect 531 8074 565 8108
rect 531 8000 565 8034
rect 531 7926 565 7960
rect 531 7852 565 7886
rect 531 7778 565 7812
rect 531 7704 565 7738
rect 531 7630 565 7664
rect 531 7556 565 7590
rect 531 7482 565 7516
rect 531 7408 565 7442
rect 531 7334 565 7368
rect 531 7260 565 7294
rect 531 7186 565 7220
rect 767 9098 801 9132
rect 767 9025 801 9059
rect 767 8952 801 8986
rect 767 8879 801 8913
rect 767 8806 801 8840
rect 767 8733 801 8767
rect 767 8660 801 8694
rect 767 8587 801 8621
rect 767 8514 801 8548
rect 767 8441 801 8475
rect 767 8368 801 8402
rect 767 8295 801 8329
rect 767 8222 801 8256
rect 767 8148 801 8182
rect 767 8074 801 8108
rect 767 8000 801 8034
rect 767 7926 801 7960
rect 767 7852 801 7886
rect 767 7778 801 7812
rect 767 7704 801 7738
rect 767 7630 801 7664
rect 767 7556 801 7590
rect 767 7482 801 7516
rect 767 7408 801 7442
rect 767 7334 801 7368
rect 767 7260 801 7294
rect 767 7186 801 7220
rect 1003 9098 1037 9132
rect 1003 9025 1037 9059
rect 1003 8952 1037 8986
rect 1003 8879 1037 8913
rect 1003 8806 1037 8840
rect 1003 8733 1037 8767
rect 1003 8660 1037 8694
rect 1003 8587 1037 8621
rect 1003 8514 1037 8548
rect 1003 8441 1037 8475
rect 1003 8368 1037 8402
rect 1003 8295 1037 8329
rect 1003 8222 1037 8256
rect 1003 8148 1037 8182
rect 1003 8074 1037 8108
rect 1003 8000 1037 8034
rect 1003 7926 1037 7960
rect 1003 7852 1037 7886
rect 1003 7778 1037 7812
rect 1003 7704 1037 7738
rect 1003 7630 1037 7664
rect 1003 7556 1037 7590
rect 1003 7482 1037 7516
rect 1003 7408 1037 7442
rect 1003 7334 1037 7368
rect 1003 7260 1037 7294
rect 1003 7186 1037 7220
rect 1239 9098 1273 9132
rect 1239 9025 1273 9059
rect 1239 8952 1273 8986
rect 1239 8879 1273 8913
rect 1239 8806 1273 8840
rect 1239 8733 1273 8767
rect 1239 8660 1273 8694
rect 1239 8587 1273 8621
rect 1239 8514 1273 8548
rect 1239 8441 1273 8475
rect 1239 8368 1273 8402
rect 1239 8295 1273 8329
rect 1239 8222 1273 8256
rect 1239 8148 1273 8182
rect 1239 8074 1273 8108
rect 1239 8000 1273 8034
rect 1239 7926 1273 7960
rect 1239 7852 1273 7886
rect 1239 7778 1273 7812
rect 1239 7704 1273 7738
rect 1239 7630 1273 7664
rect 1239 7556 1273 7590
rect 1239 7482 1273 7516
rect 1239 7408 1273 7442
rect 1239 7334 1273 7368
rect 1239 7260 1273 7294
rect 1239 7186 1273 7220
rect 1475 9098 1509 9132
rect 1475 9025 1509 9059
rect 1475 8952 1509 8986
rect 1475 8879 1509 8913
rect 1475 8806 1509 8840
rect 1475 8733 1509 8767
rect 1475 8660 1509 8694
rect 1475 8587 1509 8621
rect 1475 8514 1509 8548
rect 1475 8441 1509 8475
rect 1475 8368 1509 8402
rect 1475 8295 1509 8329
rect 1475 8222 1509 8256
rect 1475 8148 1509 8182
rect 1475 8074 1509 8108
rect 1475 8000 1509 8034
rect 1475 7926 1509 7960
rect 1475 7852 1509 7886
rect 1475 7778 1509 7812
rect 1475 7704 1509 7738
rect 1475 7630 1509 7664
rect 1475 7556 1509 7590
rect 1475 7482 1509 7516
rect 1475 7408 1509 7442
rect 1475 7334 1509 7368
rect 1475 7260 1509 7294
rect 1475 7186 1509 7220
rect 1711 9098 1745 9132
rect 1711 9025 1745 9059
rect 1711 8952 1745 8986
rect 1711 8879 1745 8913
rect 1711 8806 1745 8840
rect 1711 8733 1745 8767
rect 1711 8660 1745 8694
rect 1711 8587 1745 8621
rect 1711 8514 1745 8548
rect 1711 8441 1745 8475
rect 1711 8368 1745 8402
rect 1711 8295 1745 8329
rect 1711 8222 1745 8256
rect 1711 8148 1745 8182
rect 1711 8074 1745 8108
rect 1711 8000 1745 8034
rect 1711 7926 1745 7960
rect 1711 7852 1745 7886
rect 1711 7778 1745 7812
rect 1711 7704 1745 7738
rect 1711 7630 1745 7664
rect 1711 7556 1745 7590
rect 1711 7482 1745 7516
rect 1711 7408 1745 7442
rect 1711 7334 1745 7368
rect 1711 7260 1745 7294
rect 1711 7186 1745 7220
rect 1947 9098 1981 9132
rect 1947 9025 1981 9059
rect 1947 8952 1981 8986
rect 1947 8879 1981 8913
rect 1947 8806 1981 8840
rect 1947 8733 1981 8767
rect 1947 8660 1981 8694
rect 1947 8587 1981 8621
rect 1947 8514 1981 8548
rect 1947 8441 1981 8475
rect 1947 8368 1981 8402
rect 1947 8295 1981 8329
rect 1947 8222 1981 8256
rect 1947 8148 1981 8182
rect 1947 8074 1981 8108
rect 1947 8000 1981 8034
rect 1947 7926 1981 7960
rect 1947 7852 1981 7886
rect 1947 7778 1981 7812
rect 1947 7704 1981 7738
rect 1947 7630 1981 7664
rect 1947 7556 1981 7590
rect 1947 7482 1981 7516
rect 1947 7408 1981 7442
rect 1947 7334 1981 7368
rect 1947 7260 1981 7294
rect 1947 7186 1981 7220
rect 2183 9098 2217 9132
rect 2183 9025 2217 9059
rect 2183 8952 2217 8986
rect 2183 8879 2217 8913
rect 2183 8806 2217 8840
rect 2183 8733 2217 8767
rect 2183 8660 2217 8694
rect 2183 8587 2217 8621
rect 2183 8514 2217 8548
rect 2183 8441 2217 8475
rect 2183 8368 2217 8402
rect 2183 8295 2217 8329
rect 2183 8222 2217 8256
rect 2183 8148 2217 8182
rect 2183 8074 2217 8108
rect 2183 8000 2217 8034
rect 2183 7926 2217 7960
rect 2183 7852 2217 7886
rect 2183 7778 2217 7812
rect 2183 7704 2217 7738
rect 2183 7630 2217 7664
rect 2183 7556 2217 7590
rect 2183 7482 2217 7516
rect 2183 7408 2217 7442
rect 2183 7334 2217 7368
rect 2183 7260 2217 7294
rect 2183 7186 2217 7220
rect 2419 9098 2453 9132
rect 2419 9025 2453 9059
rect 2419 8952 2453 8986
rect 2419 8879 2453 8913
rect 2419 8806 2453 8840
rect 2419 8733 2453 8767
rect 2419 8660 2453 8694
rect 2419 8587 2453 8621
rect 2419 8514 2453 8548
rect 2419 8441 2453 8475
rect 2419 8368 2453 8402
rect 2419 8295 2453 8329
rect 2419 8222 2453 8256
rect 2419 8148 2453 8182
rect 2419 8074 2453 8108
rect 2419 8000 2453 8034
rect 2419 7926 2453 7960
rect 2419 7852 2453 7886
rect 2419 7778 2453 7812
rect 2419 7704 2453 7738
rect 2419 7630 2453 7664
rect 2419 7556 2453 7590
rect 2419 7482 2453 7516
rect 2419 7408 2453 7442
rect 2419 7334 2453 7368
rect 2419 7260 2453 7294
rect 2419 7186 2453 7220
rect 2655 9098 2689 9132
rect 2655 9025 2689 9059
rect 2655 8952 2689 8986
rect 2655 8879 2689 8913
rect 2655 8806 2689 8840
rect 2655 8733 2689 8767
rect 2655 8660 2689 8694
rect 2655 8587 2689 8621
rect 2655 8514 2689 8548
rect 2655 8441 2689 8475
rect 2655 8368 2689 8402
rect 2655 8295 2689 8329
rect 2655 8222 2689 8256
rect 2655 8148 2689 8182
rect 2655 8074 2689 8108
rect 2655 8000 2689 8034
rect 2655 7926 2689 7960
rect 2655 7852 2689 7886
rect 2655 7778 2689 7812
rect 2655 7704 2689 7738
rect 2655 7630 2689 7664
rect 2655 7556 2689 7590
rect 2655 7482 2689 7516
rect 2655 7408 2689 7442
rect 2655 7334 2689 7368
rect 2655 7260 2689 7294
rect 2655 7186 2689 7220
rect 2891 9098 2925 9132
rect 2891 9025 2925 9059
rect 2891 8952 2925 8986
rect 2891 8879 2925 8913
rect 2891 8806 2925 8840
rect 2891 8733 2925 8767
rect 2891 8660 2925 8694
rect 2891 8587 2925 8621
rect 2891 8514 2925 8548
rect 2891 8441 2925 8475
rect 2891 8368 2925 8402
rect 2891 8295 2925 8329
rect 2891 8222 2925 8256
rect 2891 8148 2925 8182
rect 2891 8074 2925 8108
rect 2891 8000 2925 8034
rect 2891 7926 2925 7960
rect 2891 7852 2925 7886
rect 2891 7778 2925 7812
rect 2891 7704 2925 7738
rect 2891 7630 2925 7664
rect 2891 7556 2925 7590
rect 2891 7482 2925 7516
rect 2891 7408 2925 7442
rect 2891 7334 2925 7368
rect 2891 7260 2925 7294
rect 2891 7186 2925 7220
rect 3036 9122 3070 9154
rect 3036 9120 3070 9122
rect 3036 9054 3070 9082
rect 3036 9048 3070 9054
rect 3036 8986 3070 9010
rect 3036 8976 3070 8986
rect 3036 8918 3070 8938
rect 3036 8904 3070 8918
rect 3036 8850 3070 8866
rect 3036 8832 3070 8850
rect 3036 8782 3070 8794
rect 3036 8760 3070 8782
rect 3036 8714 3070 8722
rect 3036 8688 3070 8714
rect 3036 8646 3070 8650
rect 3036 8616 3070 8646
rect 3036 8544 3070 8578
rect 3036 8476 3070 8506
rect 3036 8472 3070 8476
rect 3036 8408 3070 8434
rect 3036 8400 3070 8408
rect 3036 8340 3070 8362
rect 3036 8328 3070 8340
rect 3036 8272 3070 8290
rect 3036 8256 3070 8272
rect 3036 8204 3070 8218
rect 3036 8184 3070 8204
rect 3036 8136 3070 8146
rect 3036 8112 3070 8136
rect 3036 8068 3070 8074
rect 3036 8040 3070 8068
rect 3036 8000 3070 8002
rect 3036 7968 3070 8000
rect 3036 7898 3070 7930
rect 3036 7896 3070 7898
rect 3036 7830 3070 7858
rect 3036 7824 3070 7830
rect 3036 7762 3070 7786
rect 3036 7752 3070 7762
rect 3036 7694 3070 7714
rect 3036 7680 3070 7694
rect 3036 7626 3070 7642
rect 3036 7608 3070 7626
rect 3036 7558 3070 7570
rect 3036 7536 3070 7558
rect 3036 7490 3070 7498
rect 3036 7464 3070 7490
rect 3036 7422 3070 7426
rect 3036 7392 3070 7422
rect 3036 7320 3070 7354
rect 3036 7252 3070 7282
rect 3036 7248 3070 7252
rect 386 7095 420 7119
rect 386 7085 420 7095
rect 3036 7184 3070 7210
rect 3036 7176 3070 7184
rect 3036 7116 3070 7138
rect 3036 7104 3070 7116
rect 625 7070 626 7104
rect 626 7070 659 7104
rect 700 7070 732 7104
rect 732 7070 734 7104
rect 775 7070 802 7104
rect 802 7070 809 7104
rect 850 7070 872 7104
rect 872 7070 884 7104
rect 925 7070 942 7104
rect 942 7070 959 7104
rect 1000 7070 1012 7104
rect 1012 7070 1034 7104
rect 1075 7070 1082 7104
rect 1082 7070 1109 7104
rect 1150 7070 1152 7104
rect 1152 7070 1184 7104
rect 1225 7070 1256 7104
rect 1256 7070 1259 7104
rect 1300 7070 1326 7104
rect 1326 7070 1334 7104
rect 1375 7070 1396 7104
rect 1396 7070 1409 7104
rect 1450 7070 1466 7104
rect 1466 7070 1484 7104
rect 1525 7070 1536 7104
rect 1536 7070 1559 7104
rect 1600 7070 1606 7104
rect 1606 7070 1634 7104
rect 1674 7070 1676 7104
rect 1676 7070 1708 7104
rect 1748 7070 1782 7104
rect 1822 7070 1852 7104
rect 1852 7070 1856 7104
rect 1896 7070 1922 7104
rect 1922 7070 1930 7104
rect 1970 7070 1992 7104
rect 1992 7070 2004 7104
rect 2044 7070 2062 7104
rect 2062 7070 2078 7104
rect 2118 7070 2132 7104
rect 2132 7070 2152 7104
rect 2192 7070 2202 7104
rect 2202 7070 2226 7104
rect 2266 7070 2272 7104
rect 2272 7070 2300 7104
rect 2340 7070 2342 7104
rect 2342 7070 2374 7104
rect 2414 7070 2446 7104
rect 2446 7070 2448 7104
rect 2488 7070 2516 7104
rect 2516 7070 2522 7104
rect 2562 7070 2586 7104
rect 2586 7070 2596 7104
rect 2636 7070 2656 7104
rect 2656 7070 2670 7104
rect 2710 7070 2726 7104
rect 2726 7070 2744 7104
rect 2784 7070 2795 7104
rect 2795 7070 2818 7104
rect 386 7027 420 7047
rect 386 7013 420 7027
rect 3036 7048 3070 7066
rect 3036 7032 3070 7048
rect 386 6959 420 6975
rect 386 6941 420 6959
rect 386 6891 420 6903
rect 386 6869 420 6891
rect 386 6823 420 6831
rect 386 6797 420 6823
rect 386 6755 420 6759
rect 386 6725 420 6755
rect 386 6653 420 6687
rect 386 6585 420 6615
rect 386 6581 420 6585
rect 386 6517 420 6543
rect 386 6509 420 6517
rect 386 6449 420 6471
rect 386 6437 420 6449
rect 386 6381 420 6399
rect 386 6365 420 6381
rect 386 6313 420 6327
rect 386 6293 420 6313
rect 386 6245 420 6255
rect 386 6221 420 6245
rect 386 6177 420 6183
rect 386 6149 420 6177
rect 386 6109 420 6111
rect 386 6077 420 6109
rect 386 6007 420 6039
rect 386 6005 420 6007
rect 386 5939 420 5967
rect 386 5933 420 5939
rect 386 5871 420 5895
rect 386 5861 420 5871
rect 386 5803 420 5823
rect 386 5789 420 5803
rect 386 5735 420 5751
rect 386 5717 420 5735
rect 386 5667 420 5679
rect 386 5645 420 5667
rect 386 5599 420 5607
rect 386 5573 420 5599
rect 386 5531 420 5535
rect 386 5501 420 5531
rect 386 5429 420 5463
rect 386 5361 420 5391
rect 386 5357 420 5361
rect 386 5293 420 5319
rect 386 5285 420 5293
rect 386 5225 420 5247
rect 386 5213 420 5225
rect 386 5157 420 5175
rect 386 5141 420 5157
rect 386 5089 420 5103
rect 386 5069 420 5089
rect 386 5021 420 5031
rect 386 4997 420 5021
rect 531 6954 565 6988
rect 531 6881 565 6915
rect 531 6808 565 6842
rect 531 6735 565 6769
rect 531 6662 565 6696
rect 531 6589 565 6623
rect 531 6516 565 6550
rect 531 6443 565 6477
rect 531 6370 565 6404
rect 531 6297 565 6331
rect 531 6224 565 6258
rect 531 6151 565 6185
rect 531 6078 565 6112
rect 531 6004 565 6038
rect 531 5930 565 5964
rect 531 5856 565 5890
rect 531 5782 565 5816
rect 531 5708 565 5742
rect 531 5634 565 5668
rect 531 5560 565 5594
rect 531 5486 565 5520
rect 531 5412 565 5446
rect 531 5338 565 5372
rect 531 5264 565 5298
rect 531 5190 565 5224
rect 531 5116 565 5150
rect 531 5042 565 5076
rect 767 6954 801 6988
rect 767 6881 801 6915
rect 767 6808 801 6842
rect 767 6735 801 6769
rect 767 6662 801 6696
rect 767 6589 801 6623
rect 767 6516 801 6550
rect 767 6443 801 6477
rect 767 6370 801 6404
rect 767 6297 801 6331
rect 767 6224 801 6258
rect 767 6151 801 6185
rect 767 6078 801 6112
rect 767 6004 801 6038
rect 767 5930 801 5964
rect 767 5856 801 5890
rect 767 5782 801 5816
rect 767 5708 801 5742
rect 767 5634 801 5668
rect 767 5560 801 5594
rect 767 5486 801 5520
rect 767 5412 801 5446
rect 767 5338 801 5372
rect 767 5264 801 5298
rect 767 5190 801 5224
rect 767 5116 801 5150
rect 767 5042 801 5076
rect 1003 6954 1037 6988
rect 1003 6881 1037 6915
rect 1003 6808 1037 6842
rect 1003 6735 1037 6769
rect 1003 6662 1037 6696
rect 1003 6589 1037 6623
rect 1003 6516 1037 6550
rect 1003 6443 1037 6477
rect 1003 6370 1037 6404
rect 1003 6297 1037 6331
rect 1003 6224 1037 6258
rect 1003 6151 1037 6185
rect 1003 6078 1037 6112
rect 1003 6004 1037 6038
rect 1003 5930 1037 5964
rect 1003 5856 1037 5890
rect 1003 5782 1037 5816
rect 1003 5708 1037 5742
rect 1003 5634 1037 5668
rect 1003 5560 1037 5594
rect 1003 5486 1037 5520
rect 1003 5412 1037 5446
rect 1003 5338 1037 5372
rect 1003 5264 1037 5298
rect 1003 5190 1037 5224
rect 1003 5116 1037 5150
rect 1003 5042 1037 5076
rect 1239 6954 1273 6988
rect 1239 6881 1273 6915
rect 1239 6808 1273 6842
rect 1239 6735 1273 6769
rect 1239 6662 1273 6696
rect 1239 6589 1273 6623
rect 1239 6516 1273 6550
rect 1239 6443 1273 6477
rect 1239 6370 1273 6404
rect 1239 6297 1273 6331
rect 1239 6224 1273 6258
rect 1239 6151 1273 6185
rect 1239 6078 1273 6112
rect 1239 6004 1273 6038
rect 1239 5930 1273 5964
rect 1239 5856 1273 5890
rect 1239 5782 1273 5816
rect 1239 5708 1273 5742
rect 1239 5634 1273 5668
rect 1239 5560 1273 5594
rect 1239 5486 1273 5520
rect 1239 5412 1273 5446
rect 1239 5338 1273 5372
rect 1239 5264 1273 5298
rect 1239 5190 1273 5224
rect 1239 5116 1273 5150
rect 1239 5042 1273 5076
rect 1475 6954 1509 6988
rect 1475 6881 1509 6915
rect 1475 6808 1509 6842
rect 1475 6735 1509 6769
rect 1475 6662 1509 6696
rect 1475 6589 1509 6623
rect 1475 6516 1509 6550
rect 1475 6443 1509 6477
rect 1475 6370 1509 6404
rect 1475 6297 1509 6331
rect 1475 6224 1509 6258
rect 1475 6151 1509 6185
rect 1475 6078 1509 6112
rect 1475 6004 1509 6038
rect 1475 5930 1509 5964
rect 1475 5856 1509 5890
rect 1475 5782 1509 5816
rect 1475 5708 1509 5742
rect 1475 5634 1509 5668
rect 1475 5560 1509 5594
rect 1475 5486 1509 5520
rect 1475 5412 1509 5446
rect 1475 5338 1509 5372
rect 1475 5264 1509 5298
rect 1475 5190 1509 5224
rect 1475 5116 1509 5150
rect 1475 5042 1509 5076
rect 1711 6954 1745 6988
rect 1711 6881 1745 6915
rect 1711 6808 1745 6842
rect 1711 6735 1745 6769
rect 1711 6662 1745 6696
rect 1711 6589 1745 6623
rect 1711 6516 1745 6550
rect 1711 6443 1745 6477
rect 1711 6370 1745 6404
rect 1711 6297 1745 6331
rect 1711 6224 1745 6258
rect 1711 6151 1745 6185
rect 1711 6078 1745 6112
rect 1711 6004 1745 6038
rect 1711 5930 1745 5964
rect 1711 5856 1745 5890
rect 1711 5782 1745 5816
rect 1711 5708 1745 5742
rect 1711 5634 1745 5668
rect 1711 5560 1745 5594
rect 1711 5486 1745 5520
rect 1711 5412 1745 5446
rect 1711 5338 1745 5372
rect 1711 5264 1745 5298
rect 1711 5190 1745 5224
rect 1711 5116 1745 5150
rect 1711 5042 1745 5076
rect 1947 6954 1981 6988
rect 1947 6881 1981 6915
rect 1947 6808 1981 6842
rect 1947 6735 1981 6769
rect 1947 6662 1981 6696
rect 1947 6589 1981 6623
rect 1947 6516 1981 6550
rect 1947 6443 1981 6477
rect 1947 6370 1981 6404
rect 1947 6297 1981 6331
rect 1947 6224 1981 6258
rect 1947 6151 1981 6185
rect 1947 6078 1981 6112
rect 1947 6004 1981 6038
rect 1947 5930 1981 5964
rect 1947 5856 1981 5890
rect 1947 5782 1981 5816
rect 1947 5708 1981 5742
rect 1947 5634 1981 5668
rect 1947 5560 1981 5594
rect 1947 5486 1981 5520
rect 1947 5412 1981 5446
rect 1947 5338 1981 5372
rect 1947 5264 1981 5298
rect 1947 5190 1981 5224
rect 1947 5116 1981 5150
rect 1947 5042 1981 5076
rect 2183 6954 2217 6988
rect 2183 6881 2217 6915
rect 2183 6808 2217 6842
rect 2183 6735 2217 6769
rect 2183 6662 2217 6696
rect 2183 6589 2217 6623
rect 2183 6516 2217 6550
rect 2183 6443 2217 6477
rect 2183 6370 2217 6404
rect 2183 6297 2217 6331
rect 2183 6224 2217 6258
rect 2183 6151 2217 6185
rect 2183 6078 2217 6112
rect 2183 6004 2217 6038
rect 2183 5930 2217 5964
rect 2183 5856 2217 5890
rect 2183 5782 2217 5816
rect 2183 5708 2217 5742
rect 2183 5634 2217 5668
rect 2183 5560 2217 5594
rect 2183 5486 2217 5520
rect 2183 5412 2217 5446
rect 2183 5338 2217 5372
rect 2183 5264 2217 5298
rect 2183 5190 2217 5224
rect 2183 5116 2217 5150
rect 2183 5042 2217 5076
rect 2419 6954 2453 6988
rect 2419 6881 2453 6915
rect 2419 6808 2453 6842
rect 2419 6735 2453 6769
rect 2419 6662 2453 6696
rect 2419 6589 2453 6623
rect 2419 6516 2453 6550
rect 2419 6443 2453 6477
rect 2419 6370 2453 6404
rect 2419 6297 2453 6331
rect 2419 6224 2453 6258
rect 2419 6151 2453 6185
rect 2419 6078 2453 6112
rect 2419 6004 2453 6038
rect 2419 5930 2453 5964
rect 2419 5856 2453 5890
rect 2419 5782 2453 5816
rect 2419 5708 2453 5742
rect 2419 5634 2453 5668
rect 2419 5560 2453 5594
rect 2419 5486 2453 5520
rect 2419 5412 2453 5446
rect 2419 5338 2453 5372
rect 2419 5264 2453 5298
rect 2419 5190 2453 5224
rect 2419 5116 2453 5150
rect 2419 5042 2453 5076
rect 2655 6954 2689 6988
rect 2655 6881 2689 6915
rect 2655 6808 2689 6842
rect 2655 6735 2689 6769
rect 2655 6662 2689 6696
rect 2655 6589 2689 6623
rect 2655 6516 2689 6550
rect 2655 6443 2689 6477
rect 2655 6370 2689 6404
rect 2655 6297 2689 6331
rect 2655 6224 2689 6258
rect 2655 6151 2689 6185
rect 2655 6078 2689 6112
rect 2655 6004 2689 6038
rect 2655 5930 2689 5964
rect 2655 5856 2689 5890
rect 2655 5782 2689 5816
rect 2655 5708 2689 5742
rect 2655 5634 2689 5668
rect 2655 5560 2689 5594
rect 2655 5486 2689 5520
rect 2655 5412 2689 5446
rect 2655 5338 2689 5372
rect 2655 5264 2689 5298
rect 2655 5190 2689 5224
rect 2655 5116 2689 5150
rect 2655 5042 2689 5076
rect 2891 6954 2925 6988
rect 2891 6881 2925 6915
rect 2891 6808 2925 6842
rect 2891 6735 2925 6769
rect 2891 6662 2925 6696
rect 2891 6589 2925 6623
rect 2891 6516 2925 6550
rect 2891 6443 2925 6477
rect 2891 6370 2925 6404
rect 2891 6297 2925 6331
rect 2891 6224 2925 6258
rect 2891 6151 2925 6185
rect 2891 6078 2925 6112
rect 2891 6004 2925 6038
rect 2891 5930 2925 5964
rect 2891 5856 2925 5890
rect 2891 5782 2925 5816
rect 2891 5708 2925 5742
rect 2891 5634 2925 5668
rect 2891 5560 2925 5594
rect 2891 5486 2925 5520
rect 2891 5412 2925 5446
rect 2891 5338 2925 5372
rect 2891 5264 2925 5298
rect 2891 5190 2925 5224
rect 2891 5116 2925 5150
rect 2891 5042 2925 5076
rect 3036 6980 3070 6994
rect 3036 6960 3070 6980
rect 3036 6912 3070 6922
rect 3036 6888 3070 6912
rect 3036 6844 3070 6850
rect 3036 6816 3070 6844
rect 3036 6776 3070 6778
rect 3036 6744 3070 6776
rect 3036 6674 3070 6706
rect 3036 6672 3070 6674
rect 3036 6606 3070 6634
rect 3036 6600 3070 6606
rect 3036 6538 3070 6562
rect 3036 6528 3070 6538
rect 3036 6470 3070 6490
rect 3036 6456 3070 6470
rect 3036 6402 3070 6418
rect 3036 6384 3070 6402
rect 3036 6334 3070 6346
rect 3036 6312 3070 6334
rect 3036 6266 3070 6274
rect 3036 6240 3070 6266
rect 3036 6198 3070 6202
rect 3036 6168 3070 6198
rect 3036 6096 3070 6130
rect 3036 6028 3070 6058
rect 3036 6024 3070 6028
rect 3036 5960 3070 5986
rect 3036 5952 3070 5960
rect 3036 5892 3070 5914
rect 3036 5880 3070 5892
rect 3036 5824 3070 5842
rect 3036 5808 3070 5824
rect 3036 5756 3070 5770
rect 3036 5736 3070 5756
rect 3036 5688 3070 5698
rect 3036 5664 3070 5688
rect 3036 5620 3070 5626
rect 3036 5592 3070 5620
rect 3036 5552 3070 5554
rect 3036 5520 3070 5552
rect 3036 5450 3070 5482
rect 3036 5448 3070 5450
rect 3036 5382 3070 5410
rect 3036 5376 3070 5382
rect 3036 5314 3070 5338
rect 3036 5304 3070 5314
rect 3036 5246 3070 5266
rect 3036 5232 3070 5246
rect 3036 5178 3070 5194
rect 3036 5160 3070 5178
rect 3036 5110 3070 5122
rect 3036 5088 3070 5110
rect 386 4953 420 4959
rect 386 4925 420 4953
rect 3036 5042 3070 5050
rect 3036 5016 3070 5042
rect 625 4940 626 4974
rect 626 4940 659 4974
rect 700 4940 732 4974
rect 732 4940 734 4974
rect 775 4940 802 4974
rect 802 4940 809 4974
rect 850 4940 872 4974
rect 872 4940 884 4974
rect 925 4940 942 4974
rect 942 4940 959 4974
rect 1000 4940 1012 4974
rect 1012 4940 1034 4974
rect 1075 4940 1082 4974
rect 1082 4940 1109 4974
rect 1150 4940 1152 4974
rect 1152 4940 1184 4974
rect 1225 4940 1256 4974
rect 1256 4940 1259 4974
rect 1300 4940 1326 4974
rect 1326 4940 1334 4974
rect 1375 4940 1396 4974
rect 1396 4940 1409 4974
rect 1450 4940 1466 4974
rect 1466 4940 1484 4974
rect 1525 4940 1536 4974
rect 1536 4940 1559 4974
rect 1600 4940 1606 4974
rect 1606 4940 1634 4974
rect 1674 4940 1676 4974
rect 1676 4940 1708 4974
rect 1748 4940 1782 4974
rect 1822 4940 1852 4974
rect 1852 4940 1856 4974
rect 1896 4940 1922 4974
rect 1922 4940 1930 4974
rect 1970 4940 1992 4974
rect 1992 4940 2004 4974
rect 2044 4940 2062 4974
rect 2062 4940 2078 4974
rect 2118 4940 2132 4974
rect 2132 4940 2152 4974
rect 2192 4940 2202 4974
rect 2202 4940 2226 4974
rect 2266 4940 2272 4974
rect 2272 4940 2300 4974
rect 2340 4940 2342 4974
rect 2342 4940 2374 4974
rect 2414 4940 2446 4974
rect 2446 4940 2448 4974
rect 2488 4940 2516 4974
rect 2516 4940 2522 4974
rect 2562 4940 2586 4974
rect 2586 4940 2596 4974
rect 2636 4940 2656 4974
rect 2656 4940 2670 4974
rect 2710 4940 2726 4974
rect 2726 4940 2744 4974
rect 2784 4940 2795 4974
rect 2795 4940 2818 4974
rect 3036 4974 3070 4978
rect 3036 4944 3070 4974
rect 386 4885 420 4887
rect 386 4853 420 4885
rect 3036 4872 3070 4906
rect 386 4783 420 4815
rect 386 4781 420 4783
rect 386 4715 420 4743
rect 386 4709 420 4715
rect 386 4647 420 4671
rect 386 4637 420 4647
rect 386 4579 420 4599
rect 386 4565 420 4579
rect 386 4511 420 4527
rect 386 4493 420 4511
rect 386 4443 420 4455
rect 386 4421 420 4443
rect 386 4375 420 4383
rect 386 4349 420 4375
rect 386 4307 420 4311
rect 386 4277 420 4307
rect 386 4205 420 4239
rect 386 4137 420 4167
rect 386 4133 420 4137
rect 386 4069 420 4095
rect 386 4061 420 4069
rect 386 4001 420 4023
rect 386 3989 420 4001
rect 386 3933 420 3951
rect 386 3917 420 3933
rect 386 3865 420 3879
rect 386 3845 420 3865
rect 386 3797 420 3807
rect 386 3773 420 3797
rect 386 3729 420 3735
rect 386 3701 420 3729
rect 386 3661 420 3663
rect 386 3629 420 3661
rect 386 3559 420 3591
rect 386 3557 420 3559
rect 386 3491 420 3519
rect 386 3485 420 3491
rect 386 3423 420 3447
rect 386 3413 420 3423
rect 386 3355 420 3375
rect 386 3341 420 3355
rect 386 3287 420 3303
rect 386 3269 420 3287
rect 386 3219 420 3231
rect 386 3197 420 3219
rect 386 3151 420 3159
rect 386 3125 420 3151
rect 386 3083 420 3087
rect 386 3053 420 3083
rect 386 2981 420 3015
rect 386 2913 420 2943
rect 386 2909 420 2913
rect 531 4838 565 4872
rect 531 4765 565 4799
rect 531 4692 565 4726
rect 531 4619 565 4653
rect 531 4546 565 4580
rect 531 4473 565 4507
rect 531 4400 565 4434
rect 531 4327 565 4361
rect 531 4254 565 4288
rect 531 4181 565 4215
rect 531 4108 565 4142
rect 531 4035 565 4069
rect 531 3962 565 3996
rect 531 3888 565 3922
rect 531 3814 565 3848
rect 531 3740 565 3774
rect 531 3666 565 3700
rect 531 3592 565 3626
rect 531 3518 565 3552
rect 531 3444 565 3478
rect 531 3370 565 3404
rect 531 3296 565 3330
rect 531 3222 565 3256
rect 531 3148 565 3182
rect 531 3074 565 3108
rect 531 3000 565 3034
rect 531 2926 565 2960
rect 767 4838 801 4872
rect 767 4765 801 4799
rect 767 4692 801 4726
rect 767 4619 801 4653
rect 767 4546 801 4580
rect 767 4473 801 4507
rect 767 4400 801 4434
rect 767 4327 801 4361
rect 767 4254 801 4288
rect 767 4181 801 4215
rect 767 4108 801 4142
rect 767 4035 801 4069
rect 767 3962 801 3996
rect 767 3888 801 3922
rect 767 3814 801 3848
rect 767 3740 801 3774
rect 767 3666 801 3700
rect 767 3592 801 3626
rect 767 3518 801 3552
rect 767 3444 801 3478
rect 767 3370 801 3404
rect 767 3296 801 3330
rect 767 3222 801 3256
rect 767 3148 801 3182
rect 767 3074 801 3108
rect 767 3000 801 3034
rect 767 2926 801 2960
rect 1003 4838 1037 4872
rect 1003 4765 1037 4799
rect 1003 4692 1037 4726
rect 1003 4619 1037 4653
rect 1003 4546 1037 4580
rect 1003 4473 1037 4507
rect 1003 4400 1037 4434
rect 1003 4327 1037 4361
rect 1003 4254 1037 4288
rect 1003 4181 1037 4215
rect 1003 4108 1037 4142
rect 1003 4035 1037 4069
rect 1003 3962 1037 3996
rect 1003 3888 1037 3922
rect 1003 3814 1037 3848
rect 1003 3740 1037 3774
rect 1003 3666 1037 3700
rect 1003 3592 1037 3626
rect 1003 3518 1037 3552
rect 1003 3444 1037 3478
rect 1003 3370 1037 3404
rect 1003 3296 1037 3330
rect 1003 3222 1037 3256
rect 1003 3148 1037 3182
rect 1003 3074 1037 3108
rect 1003 3000 1037 3034
rect 1003 2926 1037 2960
rect 1239 4838 1273 4872
rect 1239 4765 1273 4799
rect 1239 4692 1273 4726
rect 1239 4619 1273 4653
rect 1239 4546 1273 4580
rect 1239 4473 1273 4507
rect 1239 4400 1273 4434
rect 1239 4327 1273 4361
rect 1239 4254 1273 4288
rect 1239 4181 1273 4215
rect 1239 4108 1273 4142
rect 1239 4035 1273 4069
rect 1239 3962 1273 3996
rect 1239 3888 1273 3922
rect 1239 3814 1273 3848
rect 1239 3740 1273 3774
rect 1239 3666 1273 3700
rect 1239 3592 1273 3626
rect 1239 3518 1273 3552
rect 1239 3444 1273 3478
rect 1239 3370 1273 3404
rect 1239 3296 1273 3330
rect 1239 3222 1273 3256
rect 1239 3148 1273 3182
rect 1239 3074 1273 3108
rect 1239 3000 1273 3034
rect 1239 2926 1273 2960
rect 1475 4838 1509 4872
rect 1475 4765 1509 4799
rect 1475 4692 1509 4726
rect 1475 4619 1509 4653
rect 1475 4546 1509 4580
rect 1475 4473 1509 4507
rect 1475 4400 1509 4434
rect 1475 4327 1509 4361
rect 1475 4254 1509 4288
rect 1475 4181 1509 4215
rect 1475 4108 1509 4142
rect 1475 4035 1509 4069
rect 1475 3962 1509 3996
rect 1475 3888 1509 3922
rect 1475 3814 1509 3848
rect 1475 3740 1509 3774
rect 1475 3666 1509 3700
rect 1475 3592 1509 3626
rect 1475 3518 1509 3552
rect 1475 3444 1509 3478
rect 1475 3370 1509 3404
rect 1475 3296 1509 3330
rect 1475 3222 1509 3256
rect 1475 3148 1509 3182
rect 1475 3074 1509 3108
rect 1475 3000 1509 3034
rect 1475 2926 1509 2960
rect 1711 4838 1745 4872
rect 1711 4765 1745 4799
rect 1711 4692 1745 4726
rect 1711 4619 1745 4653
rect 1711 4546 1745 4580
rect 1711 4473 1745 4507
rect 1711 4400 1745 4434
rect 1711 4327 1745 4361
rect 1711 4254 1745 4288
rect 1711 4181 1745 4215
rect 1711 4108 1745 4142
rect 1711 4035 1745 4069
rect 1711 3962 1745 3996
rect 1711 3888 1745 3922
rect 1711 3814 1745 3848
rect 1711 3740 1745 3774
rect 1711 3666 1745 3700
rect 1711 3592 1745 3626
rect 1711 3518 1745 3552
rect 1711 3444 1745 3478
rect 1711 3370 1745 3404
rect 1711 3296 1745 3330
rect 1711 3222 1745 3256
rect 1711 3148 1745 3182
rect 1711 3074 1745 3108
rect 1711 3000 1745 3034
rect 1711 2926 1745 2960
rect 1947 4838 1981 4872
rect 1947 4765 1981 4799
rect 1947 4692 1981 4726
rect 1947 4619 1981 4653
rect 1947 4546 1981 4580
rect 1947 4473 1981 4507
rect 1947 4400 1981 4434
rect 1947 4327 1981 4361
rect 1947 4254 1981 4288
rect 1947 4181 1981 4215
rect 1947 4108 1981 4142
rect 1947 4035 1981 4069
rect 1947 3962 1981 3996
rect 1947 3888 1981 3922
rect 1947 3814 1981 3848
rect 1947 3740 1981 3774
rect 1947 3666 1981 3700
rect 1947 3592 1981 3626
rect 1947 3518 1981 3552
rect 1947 3444 1981 3478
rect 1947 3370 1981 3404
rect 1947 3296 1981 3330
rect 1947 3222 1981 3256
rect 1947 3148 1981 3182
rect 1947 3074 1981 3108
rect 1947 3000 1981 3034
rect 1947 2926 1981 2960
rect 2183 4838 2217 4872
rect 2183 4765 2217 4799
rect 2183 4692 2217 4726
rect 2183 4619 2217 4653
rect 2183 4546 2217 4580
rect 2183 4473 2217 4507
rect 2183 4400 2217 4434
rect 2183 4327 2217 4361
rect 2183 4254 2217 4288
rect 2183 4181 2217 4215
rect 2183 4108 2217 4142
rect 2183 4035 2217 4069
rect 2183 3962 2217 3996
rect 2183 3888 2217 3922
rect 2183 3814 2217 3848
rect 2183 3740 2217 3774
rect 2183 3666 2217 3700
rect 2183 3592 2217 3626
rect 2183 3518 2217 3552
rect 2183 3444 2217 3478
rect 2183 3370 2217 3404
rect 2183 3296 2217 3330
rect 2183 3222 2217 3256
rect 2183 3148 2217 3182
rect 2183 3074 2217 3108
rect 2183 3000 2217 3034
rect 2183 2926 2217 2960
rect 2419 4838 2453 4872
rect 2419 4765 2453 4799
rect 2419 4692 2453 4726
rect 2419 4619 2453 4653
rect 2419 4546 2453 4580
rect 2419 4473 2453 4507
rect 2419 4400 2453 4434
rect 2419 4327 2453 4361
rect 2419 4254 2453 4288
rect 2419 4181 2453 4215
rect 2419 4108 2453 4142
rect 2419 4035 2453 4069
rect 2419 3962 2453 3996
rect 2419 3888 2453 3922
rect 2419 3814 2453 3848
rect 2419 3740 2453 3774
rect 2419 3666 2453 3700
rect 2419 3592 2453 3626
rect 2419 3518 2453 3552
rect 2419 3444 2453 3478
rect 2419 3370 2453 3404
rect 2419 3296 2453 3330
rect 2419 3222 2453 3256
rect 2419 3148 2453 3182
rect 2419 3074 2453 3108
rect 2419 3000 2453 3034
rect 2419 2926 2453 2960
rect 2655 4838 2689 4872
rect 2655 4765 2689 4799
rect 2655 4692 2689 4726
rect 2655 4619 2689 4653
rect 2655 4546 2689 4580
rect 2655 4473 2689 4507
rect 2655 4400 2689 4434
rect 2655 4327 2689 4361
rect 2655 4254 2689 4288
rect 2655 4181 2689 4215
rect 2655 4108 2689 4142
rect 2655 4035 2689 4069
rect 2655 3962 2689 3996
rect 2655 3888 2689 3922
rect 2655 3814 2689 3848
rect 2655 3740 2689 3774
rect 2655 3666 2689 3700
rect 2655 3592 2689 3626
rect 2655 3518 2689 3552
rect 2655 3444 2689 3478
rect 2655 3370 2689 3404
rect 2655 3296 2689 3330
rect 2655 3222 2689 3256
rect 2655 3148 2689 3182
rect 2655 3074 2689 3108
rect 2655 3000 2689 3034
rect 2655 2926 2689 2960
rect 2891 4838 2925 4872
rect 2891 4765 2925 4799
rect 2891 4692 2925 4726
rect 2891 4619 2925 4653
rect 2891 4546 2925 4580
rect 2891 4473 2925 4507
rect 2891 4400 2925 4434
rect 2891 4327 2925 4361
rect 2891 4254 2925 4288
rect 2891 4181 2925 4215
rect 2891 4108 2925 4142
rect 2891 4035 2925 4069
rect 2891 3962 2925 3996
rect 2891 3888 2925 3922
rect 2891 3814 2925 3848
rect 2891 3740 2925 3774
rect 2891 3666 2925 3700
rect 2891 3592 2925 3626
rect 2891 3518 2925 3552
rect 2891 3444 2925 3478
rect 2891 3370 2925 3404
rect 2891 3296 2925 3330
rect 2891 3222 2925 3256
rect 2891 3148 2925 3182
rect 2891 3074 2925 3108
rect 2891 3000 2925 3034
rect 2891 2926 2925 2960
rect 3036 4804 3070 4834
rect 3036 4800 3070 4804
rect 3036 4736 3070 4762
rect 3036 4728 3070 4736
rect 3036 4668 3070 4690
rect 3036 4656 3070 4668
rect 3036 4600 3070 4618
rect 3036 4584 3070 4600
rect 3036 4532 3070 4546
rect 3036 4512 3070 4532
rect 3036 4464 3070 4474
rect 3036 4440 3070 4464
rect 3036 4396 3070 4402
rect 3036 4368 3070 4396
rect 3036 4328 3070 4330
rect 3036 4296 3070 4328
rect 3036 4226 3070 4258
rect 3036 4224 3070 4226
rect 3036 4158 3070 4186
rect 3036 4152 3070 4158
rect 3036 4090 3070 4114
rect 3036 4080 3070 4090
rect 3036 4022 3070 4042
rect 3036 4008 3070 4022
rect 3036 3954 3070 3970
rect 3036 3936 3070 3954
rect 3036 3886 3070 3898
rect 3036 3864 3070 3886
rect 3036 3818 3070 3826
rect 3036 3792 3070 3818
rect 3036 3750 3070 3754
rect 3036 3720 3070 3750
rect 3036 3648 3070 3682
rect 3036 3580 3070 3610
rect 3036 3576 3070 3580
rect 3036 3512 3070 3538
rect 3036 3504 3070 3512
rect 3036 3444 3070 3466
rect 3036 3432 3070 3444
rect 3036 3376 3070 3394
rect 3036 3360 3070 3376
rect 3036 3308 3070 3322
rect 3036 3288 3070 3308
rect 3036 3240 3070 3250
rect 3036 3216 3070 3240
rect 3036 3172 3070 3178
rect 3036 3144 3070 3172
rect 3036 3104 3070 3106
rect 3036 3072 3070 3104
rect 3036 3002 3070 3034
rect 3036 3000 3070 3002
rect 386 2845 420 2871
rect 386 2837 420 2845
rect 3036 2934 3070 2962
rect 3036 2928 3070 2934
rect 386 2777 420 2799
rect 386 2765 420 2777
rect 625 2810 626 2844
rect 626 2810 659 2844
rect 700 2810 732 2844
rect 732 2810 734 2844
rect 775 2810 802 2844
rect 802 2810 809 2844
rect 850 2810 872 2844
rect 872 2810 884 2844
rect 925 2810 942 2844
rect 942 2810 959 2844
rect 1000 2810 1012 2844
rect 1012 2810 1034 2844
rect 1075 2810 1082 2844
rect 1082 2810 1109 2844
rect 1150 2810 1152 2844
rect 1152 2810 1184 2844
rect 1225 2810 1256 2844
rect 1256 2810 1259 2844
rect 1300 2810 1326 2844
rect 1326 2810 1334 2844
rect 1375 2810 1396 2844
rect 1396 2810 1409 2844
rect 1450 2810 1466 2844
rect 1466 2810 1484 2844
rect 1525 2810 1536 2844
rect 1536 2810 1559 2844
rect 1600 2810 1606 2844
rect 1606 2810 1634 2844
rect 1674 2810 1676 2844
rect 1676 2810 1708 2844
rect 1748 2810 1782 2844
rect 1822 2810 1852 2844
rect 1852 2810 1856 2844
rect 1896 2810 1922 2844
rect 1922 2810 1930 2844
rect 1970 2810 1992 2844
rect 1992 2810 2004 2844
rect 2044 2810 2062 2844
rect 2062 2810 2078 2844
rect 2118 2810 2132 2844
rect 2132 2810 2152 2844
rect 2192 2810 2202 2844
rect 2202 2810 2226 2844
rect 2266 2810 2272 2844
rect 2272 2810 2300 2844
rect 2340 2810 2342 2844
rect 2342 2810 2374 2844
rect 2414 2810 2446 2844
rect 2446 2810 2448 2844
rect 2488 2810 2516 2844
rect 2516 2810 2522 2844
rect 2562 2810 2586 2844
rect 2586 2810 2596 2844
rect 2636 2810 2656 2844
rect 2656 2810 2670 2844
rect 2710 2810 2726 2844
rect 2726 2810 2744 2844
rect 2784 2810 2795 2844
rect 2795 2810 2818 2844
rect 3036 2866 3070 2890
rect 3036 2856 3070 2866
rect 386 2709 420 2727
rect 386 2693 420 2709
rect 3036 2798 3070 2818
rect 3036 2784 3070 2798
rect 386 2641 420 2655
rect 386 2621 420 2641
rect 386 2573 420 2583
rect 386 2549 420 2573
rect 386 2505 420 2511
rect 386 2477 420 2505
rect 386 2437 420 2439
rect 386 2405 420 2437
rect 386 2335 420 2367
rect 386 2333 420 2335
rect 386 2267 420 2295
rect 386 2261 420 2267
rect 386 2199 420 2223
rect 386 2189 420 2199
rect 386 2131 420 2151
rect 386 2117 420 2131
rect 386 2063 420 2079
rect 386 2045 420 2063
rect 386 1995 420 2007
rect 386 1973 420 1995
rect 386 1927 420 1935
rect 386 1901 420 1927
rect 386 1859 420 1863
rect 386 1829 420 1859
rect 386 1757 420 1791
rect 386 1689 420 1719
rect 386 1685 420 1689
rect 386 1621 420 1647
rect 386 1613 420 1621
rect 386 1553 420 1575
rect 386 1541 420 1553
rect 386 1485 420 1503
rect 386 1469 420 1485
rect 386 1417 420 1431
rect 386 1397 420 1417
rect 386 1349 420 1359
rect 386 1325 420 1349
rect 386 1281 420 1287
rect 386 1253 420 1281
rect 386 1213 420 1215
rect 386 1181 420 1213
rect 386 1111 420 1143
rect 386 1109 420 1111
rect 386 1043 420 1071
rect 386 1037 420 1043
rect 386 975 420 999
rect 386 965 420 975
rect 386 907 420 927
rect 386 893 420 907
rect 386 839 420 855
rect 386 821 420 839
rect 386 771 420 783
rect 386 749 420 771
rect 531 2686 565 2720
rect 531 2613 565 2647
rect 531 2540 565 2574
rect 531 2467 565 2501
rect 531 2394 565 2428
rect 531 2321 565 2355
rect 531 2248 565 2282
rect 531 2175 565 2209
rect 531 2102 565 2136
rect 531 2029 565 2063
rect 531 1956 565 1990
rect 531 1883 565 1917
rect 531 1810 565 1844
rect 531 1736 565 1770
rect 531 1662 565 1696
rect 531 1588 565 1622
rect 531 1514 565 1548
rect 531 1440 565 1474
rect 531 1366 565 1400
rect 531 1292 565 1326
rect 531 1218 565 1252
rect 531 1144 565 1178
rect 531 1070 565 1104
rect 531 996 565 1030
rect 531 922 565 956
rect 531 848 565 882
rect 531 774 565 808
rect 767 2686 801 2720
rect 767 2613 801 2647
rect 767 2540 801 2574
rect 767 2467 801 2501
rect 767 2394 801 2428
rect 767 2321 801 2355
rect 767 2248 801 2282
rect 767 2175 801 2209
rect 767 2102 801 2136
rect 767 2029 801 2063
rect 767 1956 801 1990
rect 767 1883 801 1917
rect 767 1810 801 1844
rect 767 1736 801 1770
rect 767 1662 801 1696
rect 767 1588 801 1622
rect 767 1514 801 1548
rect 767 1440 801 1474
rect 767 1366 801 1400
rect 767 1292 801 1326
rect 767 1218 801 1252
rect 767 1144 801 1178
rect 767 1070 801 1104
rect 767 996 801 1030
rect 767 922 801 956
rect 767 848 801 882
rect 767 774 801 808
rect 1003 2686 1037 2720
rect 1003 2613 1037 2647
rect 1003 2540 1037 2574
rect 1003 2467 1037 2501
rect 1003 2394 1037 2428
rect 1003 2321 1037 2355
rect 1003 2248 1037 2282
rect 1003 2175 1037 2209
rect 1003 2102 1037 2136
rect 1003 2029 1037 2063
rect 1003 1956 1037 1990
rect 1003 1883 1037 1917
rect 1003 1810 1037 1844
rect 1003 1736 1037 1770
rect 1003 1662 1037 1696
rect 1003 1588 1037 1622
rect 1003 1514 1037 1548
rect 1003 1440 1037 1474
rect 1003 1366 1037 1400
rect 1003 1292 1037 1326
rect 1003 1218 1037 1252
rect 1003 1144 1037 1178
rect 1003 1070 1037 1104
rect 1003 996 1037 1030
rect 1003 922 1037 956
rect 1003 848 1037 882
rect 1003 774 1037 808
rect 1239 2686 1273 2720
rect 1239 2613 1273 2647
rect 1239 2540 1273 2574
rect 1239 2467 1273 2501
rect 1239 2394 1273 2428
rect 1239 2321 1273 2355
rect 1239 2248 1273 2282
rect 1239 2175 1273 2209
rect 1239 2102 1273 2136
rect 1239 2029 1273 2063
rect 1239 1956 1273 1990
rect 1239 1883 1273 1917
rect 1239 1810 1273 1844
rect 1239 1736 1273 1770
rect 1239 1662 1273 1696
rect 1239 1588 1273 1622
rect 1239 1514 1273 1548
rect 1239 1440 1273 1474
rect 1239 1366 1273 1400
rect 1239 1292 1273 1326
rect 1239 1218 1273 1252
rect 1239 1144 1273 1178
rect 1239 1070 1273 1104
rect 1239 996 1273 1030
rect 1239 922 1273 956
rect 1239 848 1273 882
rect 1239 774 1273 808
rect 1475 2686 1509 2720
rect 1475 2613 1509 2647
rect 1475 2540 1509 2574
rect 1475 2467 1509 2501
rect 1475 2394 1509 2428
rect 1475 2321 1509 2355
rect 1475 2248 1509 2282
rect 1475 2175 1509 2209
rect 1475 2102 1509 2136
rect 1475 2029 1509 2063
rect 1475 1956 1509 1990
rect 1475 1883 1509 1917
rect 1475 1810 1509 1844
rect 1475 1736 1509 1770
rect 1475 1662 1509 1696
rect 1475 1588 1509 1622
rect 1475 1514 1509 1548
rect 1475 1440 1509 1474
rect 1475 1366 1509 1400
rect 1475 1292 1509 1326
rect 1475 1218 1509 1252
rect 1475 1144 1509 1178
rect 1475 1070 1509 1104
rect 1475 996 1509 1030
rect 1475 922 1509 956
rect 1475 848 1509 882
rect 1475 774 1509 808
rect 1711 2686 1745 2720
rect 1711 2613 1745 2647
rect 1711 2540 1745 2574
rect 1711 2467 1745 2501
rect 1711 2394 1745 2428
rect 1711 2321 1745 2355
rect 1711 2248 1745 2282
rect 1711 2175 1745 2209
rect 1711 2102 1745 2136
rect 1711 2029 1745 2063
rect 1711 1956 1745 1990
rect 1711 1883 1745 1917
rect 1711 1810 1745 1844
rect 1711 1736 1745 1770
rect 1711 1662 1745 1696
rect 1711 1588 1745 1622
rect 1711 1514 1745 1548
rect 1711 1440 1745 1474
rect 1711 1366 1745 1400
rect 1711 1292 1745 1326
rect 1711 1218 1745 1252
rect 1711 1144 1745 1178
rect 1711 1070 1745 1104
rect 1711 996 1745 1030
rect 1711 922 1745 956
rect 1711 848 1745 882
rect 1711 774 1745 808
rect 1947 2686 1981 2720
rect 1947 2613 1981 2647
rect 1947 2540 1981 2574
rect 1947 2467 1981 2501
rect 1947 2394 1981 2428
rect 1947 2321 1981 2355
rect 1947 2248 1981 2282
rect 1947 2175 1981 2209
rect 1947 2102 1981 2136
rect 1947 2029 1981 2063
rect 1947 1956 1981 1990
rect 1947 1883 1981 1917
rect 1947 1810 1981 1844
rect 1947 1736 1981 1770
rect 1947 1662 1981 1696
rect 1947 1588 1981 1622
rect 1947 1514 1981 1548
rect 1947 1440 1981 1474
rect 1947 1366 1981 1400
rect 1947 1292 1981 1326
rect 1947 1218 1981 1252
rect 1947 1144 1981 1178
rect 1947 1070 1981 1104
rect 1947 996 1981 1030
rect 1947 922 1981 956
rect 1947 848 1981 882
rect 1947 774 1981 808
rect 2183 2686 2217 2720
rect 2183 2613 2217 2647
rect 2183 2540 2217 2574
rect 2183 2467 2217 2501
rect 2183 2394 2217 2428
rect 2183 2321 2217 2355
rect 2183 2248 2217 2282
rect 2183 2175 2217 2209
rect 2183 2102 2217 2136
rect 2183 2029 2217 2063
rect 2183 1956 2217 1990
rect 2183 1883 2217 1917
rect 2183 1810 2217 1844
rect 2183 1736 2217 1770
rect 2183 1662 2217 1696
rect 2183 1588 2217 1622
rect 2183 1514 2217 1548
rect 2183 1440 2217 1474
rect 2183 1366 2217 1400
rect 2183 1292 2217 1326
rect 2183 1218 2217 1252
rect 2183 1144 2217 1178
rect 2183 1070 2217 1104
rect 2183 996 2217 1030
rect 2183 922 2217 956
rect 2183 848 2217 882
rect 2183 774 2217 808
rect 2419 2686 2453 2720
rect 2419 2613 2453 2647
rect 2419 2540 2453 2574
rect 2419 2467 2453 2501
rect 2419 2394 2453 2428
rect 2419 2321 2453 2355
rect 2419 2248 2453 2282
rect 2419 2175 2453 2209
rect 2419 2102 2453 2136
rect 2419 2029 2453 2063
rect 2419 1956 2453 1990
rect 2419 1883 2453 1917
rect 2419 1810 2453 1844
rect 2419 1736 2453 1770
rect 2419 1662 2453 1696
rect 2419 1588 2453 1622
rect 2419 1514 2453 1548
rect 2419 1440 2453 1474
rect 2419 1366 2453 1400
rect 2419 1292 2453 1326
rect 2419 1218 2453 1252
rect 2419 1144 2453 1178
rect 2419 1070 2453 1104
rect 2419 996 2453 1030
rect 2419 922 2453 956
rect 2419 848 2453 882
rect 2419 774 2453 808
rect 2655 2686 2689 2720
rect 2655 2613 2689 2647
rect 2655 2540 2689 2574
rect 2655 2467 2689 2501
rect 2655 2394 2689 2428
rect 2655 2321 2689 2355
rect 2655 2248 2689 2282
rect 2655 2175 2689 2209
rect 2655 2102 2689 2136
rect 2655 2029 2689 2063
rect 2655 1956 2689 1990
rect 2655 1883 2689 1917
rect 2655 1810 2689 1844
rect 2655 1736 2689 1770
rect 2655 1662 2689 1696
rect 2655 1588 2689 1622
rect 2655 1514 2689 1548
rect 2655 1440 2689 1474
rect 2655 1366 2689 1400
rect 2655 1292 2689 1326
rect 2655 1218 2689 1252
rect 2655 1144 2689 1178
rect 2655 1070 2689 1104
rect 2655 996 2689 1030
rect 2655 922 2689 956
rect 2655 848 2689 882
rect 2655 774 2689 808
rect 2891 2678 2925 2712
rect 2891 2605 2925 2639
rect 2891 2532 2925 2566
rect 2891 2459 2925 2493
rect 2891 2386 2925 2420
rect 2891 2313 2925 2347
rect 2891 2240 2925 2274
rect 2891 2167 2925 2201
rect 2891 2094 2925 2128
rect 2891 2021 2925 2055
rect 2891 1948 2925 1982
rect 2891 1875 2925 1909
rect 2891 1802 2925 1836
rect 2891 1728 2925 1762
rect 2891 1654 2925 1688
rect 2891 1580 2925 1614
rect 2891 1506 2925 1540
rect 2891 1432 2925 1466
rect 2891 1358 2925 1392
rect 2891 1284 2925 1318
rect 2891 1210 2925 1244
rect 2891 1136 2925 1170
rect 2891 1062 2925 1096
rect 2891 988 2925 1022
rect 2891 914 2925 948
rect 2891 840 2925 874
rect 2891 766 2925 800
rect 3036 2730 3070 2746
rect 3036 2712 3070 2730
rect 3036 2662 3070 2674
rect 3036 2640 3070 2662
rect 3036 2594 3070 2602
rect 3036 2568 3070 2594
rect 3036 2526 3070 2530
rect 3036 2496 3070 2526
rect 3036 2424 3070 2458
rect 3036 2356 3070 2386
rect 3036 2352 3070 2356
rect 3036 2288 3070 2314
rect 3036 2280 3070 2288
rect 3036 2220 3070 2242
rect 3036 2208 3070 2220
rect 3036 2152 3070 2170
rect 3036 2136 3070 2152
rect 3036 2084 3070 2098
rect 3036 2064 3070 2084
rect 3036 2016 3070 2026
rect 3036 1992 3070 2016
rect 3036 1948 3070 1953
rect 3036 1919 3070 1948
rect 3036 1846 3070 1880
rect 3036 1778 3070 1807
rect 3036 1773 3070 1778
rect 3036 1710 3070 1734
rect 3036 1700 3070 1710
rect 3036 1642 3070 1661
rect 3036 1627 3070 1642
rect 3036 1574 3070 1588
rect 3036 1554 3070 1574
rect 3036 1506 3070 1515
rect 3036 1481 3070 1506
rect 3036 1438 3070 1442
rect 3036 1408 3070 1438
rect 3036 1336 3070 1369
rect 3036 1335 3070 1336
rect 3036 1268 3070 1296
rect 3036 1262 3070 1268
rect 3036 1200 3070 1223
rect 3036 1189 3070 1200
rect 3036 1132 3070 1150
rect 3036 1116 3070 1132
rect 3036 1064 3070 1077
rect 3036 1043 3070 1064
rect 3036 996 3070 1004
rect 3036 970 3070 996
rect 3036 928 3070 931
rect 3036 897 3070 928
rect 3036 826 3070 858
rect 3036 824 3070 826
rect 3036 758 3070 785
rect 3036 751 3070 758
rect 386 703 420 711
rect 386 677 420 703
rect 625 680 626 714
rect 626 680 659 714
rect 700 680 732 714
rect 732 680 734 714
rect 775 680 802 714
rect 802 680 809 714
rect 850 680 872 714
rect 872 680 884 714
rect 925 680 942 714
rect 942 680 959 714
rect 1000 680 1012 714
rect 1012 680 1034 714
rect 1075 680 1082 714
rect 1082 680 1109 714
rect 1150 680 1152 714
rect 1152 680 1184 714
rect 1225 680 1256 714
rect 1256 680 1259 714
rect 1300 680 1326 714
rect 1326 680 1334 714
rect 1375 680 1396 714
rect 1396 680 1409 714
rect 1450 680 1466 714
rect 1466 680 1484 714
rect 1525 680 1536 714
rect 1536 680 1559 714
rect 1600 680 1606 714
rect 1606 680 1634 714
rect 1674 680 1676 714
rect 1676 680 1708 714
rect 1748 680 1782 714
rect 1822 680 1852 714
rect 1852 680 1856 714
rect 1896 680 1922 714
rect 1922 680 1930 714
rect 1970 680 1992 714
rect 1992 680 2004 714
rect 2044 680 2062 714
rect 2062 680 2078 714
rect 2118 680 2132 714
rect 2132 680 2152 714
rect 2192 680 2202 714
rect 2202 680 2226 714
rect 2266 680 2272 714
rect 2272 680 2300 714
rect 2340 680 2342 714
rect 2342 680 2374 714
rect 2414 680 2446 714
rect 2446 680 2448 714
rect 2488 680 2516 714
rect 2516 680 2522 714
rect 2562 680 2586 714
rect 2586 680 2596 714
rect 2636 680 2656 714
rect 2656 680 2670 714
rect 2710 680 2726 714
rect 2726 680 2744 714
rect 2784 680 2795 714
rect 2795 680 2818 714
rect 386 605 420 639
rect 3036 690 3070 712
rect 3036 678 3070 690
rect 3036 622 3070 639
rect 3036 605 3070 622
rect 458 533 475 567
rect 475 533 492 567
rect 532 533 543 567
rect 543 533 566 567
rect 606 533 611 567
rect 611 533 640 567
rect 680 533 713 567
rect 713 533 714 567
rect 754 533 781 567
rect 781 533 788 567
rect 828 533 849 567
rect 849 533 862 567
rect 902 533 917 567
rect 917 533 936 567
rect 976 533 985 567
rect 985 533 1010 567
rect 1050 533 1053 567
rect 1053 533 1084 567
rect 1124 533 1155 567
rect 1155 533 1158 567
rect 1198 533 1223 567
rect 1223 533 1232 567
rect 1272 533 1291 567
rect 1291 533 1306 567
rect 1346 533 1359 567
rect 1359 533 1380 567
rect 1420 533 1427 567
rect 1427 533 1454 567
rect 1494 533 1495 567
rect 1495 533 1528 567
rect 1568 533 1597 567
rect 1597 533 1602 567
rect 1642 533 1665 567
rect 1665 533 1676 567
rect 1716 533 1733 567
rect 1733 533 1750 567
rect 1790 533 1801 567
rect 1801 533 1824 567
rect 1864 533 1869 567
rect 1869 533 1898 567
rect 1938 533 1971 567
rect 1971 533 1972 567
rect 2012 533 2039 567
rect 2039 533 2046 567
rect 2086 533 2107 567
rect 2107 533 2120 567
rect 2160 533 2175 567
rect 2175 533 2194 567
rect 2233 533 2243 567
rect 2243 533 2267 567
rect 2306 533 2311 567
rect 2311 533 2340 567
rect 2379 533 2413 567
rect 2452 533 2481 567
rect 2481 533 2486 567
rect 2525 533 2549 567
rect 2549 533 2559 567
rect 2598 533 2617 567
rect 2617 533 2632 567
rect 2671 533 2685 567
rect 2685 533 2705 567
rect 2744 533 2753 567
rect 2753 533 2778 567
rect 2817 533 2821 567
rect 2821 533 2851 567
rect 2890 533 2923 567
rect 2923 533 2924 567
rect 2963 533 2991 567
rect 2991 533 2997 567
rect 3296 39192 3330 39226
rect 3296 39124 3330 39154
rect 3296 39120 3330 39124
rect 3296 39056 3330 39082
rect 3296 39048 3330 39056
rect 3296 38988 3330 39010
rect 3296 38976 3330 38988
rect 3296 38920 3330 38938
rect 3296 38904 3330 38920
rect 3296 38852 3330 38866
rect 3296 38832 3330 38852
rect 3296 38784 3330 38794
rect 3296 38760 3330 38784
rect 3296 38716 3330 38722
rect 3296 38688 3330 38716
rect 3296 38648 3330 38650
rect 3296 38616 3330 38648
rect 3296 38546 3330 38578
rect 3296 38544 3330 38546
rect 3296 38478 3330 38506
rect 3296 38472 3330 38478
rect 3296 38410 3330 38434
rect 3296 38400 3330 38410
rect 3296 38342 3330 38362
rect 3296 38328 3330 38342
rect 3296 38274 3330 38290
rect 3296 38256 3330 38274
rect 3296 38206 3330 38218
rect 3296 38184 3330 38206
rect 3296 38138 3330 38146
rect 3296 38112 3330 38138
rect 3296 38070 3330 38074
rect 3296 38040 3330 38070
rect 3296 37968 3330 38002
rect 3296 37900 3330 37930
rect 3296 37896 3330 37900
rect 3296 37832 3330 37858
rect 3296 37824 3330 37832
rect 3296 37764 3330 37786
rect 3296 37752 3330 37764
rect 3296 37696 3330 37714
rect 3296 37680 3330 37696
rect 3296 37628 3330 37642
rect 3296 37608 3330 37628
rect 3296 37560 3330 37570
rect 3296 37536 3330 37560
rect 3296 37492 3330 37498
rect 3296 37464 3330 37492
rect 3296 37424 3330 37426
rect 3296 37392 3330 37424
rect 3296 37322 3330 37354
rect 3296 37320 3330 37322
rect 3296 37254 3330 37282
rect 3296 37248 3330 37254
rect 3296 37186 3330 37210
rect 3296 37176 3330 37186
rect 3296 37118 3330 37138
rect 3296 37104 3330 37118
rect 3296 37050 3330 37066
rect 3296 37032 3330 37050
rect 3296 36982 3330 36994
rect 3296 36960 3330 36982
rect 3296 36914 3330 36922
rect 3296 36888 3330 36914
rect 3296 36846 3330 36850
rect 3296 36816 3330 36846
rect 3296 36744 3330 36778
rect 3296 36676 3330 36706
rect 3296 36672 3330 36676
rect 3296 36608 3330 36634
rect 3296 36600 3330 36608
rect 3296 36540 3330 36562
rect 3296 36528 3330 36540
rect 3296 36472 3330 36490
rect 3296 36456 3330 36472
rect 3296 36404 3330 36418
rect 3296 36384 3330 36404
rect 3296 36336 3330 36346
rect 3296 36312 3330 36336
rect 3296 36268 3330 36274
rect 3296 36240 3330 36268
rect 3296 36200 3330 36202
rect 3296 36168 3330 36200
rect 3296 36098 3330 36130
rect 3296 36096 3330 36098
rect 3296 36030 3330 36058
rect 3296 36024 3330 36030
rect 3296 35962 3330 35986
rect 3296 35952 3330 35962
rect 3296 35894 3330 35914
rect 3296 35880 3330 35894
rect 3296 35826 3330 35842
rect 3296 35808 3330 35826
rect 3296 35758 3330 35770
rect 3296 35736 3330 35758
rect 3296 35690 3330 35698
rect 3296 35664 3330 35690
rect 3296 35622 3330 35626
rect 3296 35592 3330 35622
rect 3296 35520 3330 35554
rect 3296 35452 3330 35482
rect 3296 35448 3330 35452
rect 3296 35384 3330 35410
rect 3296 35376 3330 35384
rect 3296 35316 3330 35338
rect 3296 35304 3330 35316
rect 3296 35248 3330 35266
rect 3296 35232 3330 35248
rect 3296 35180 3330 35194
rect 3296 35160 3330 35180
rect 3296 35112 3330 35122
rect 3296 35088 3330 35112
rect 3296 35044 3330 35050
rect 3296 35016 3330 35044
rect 3296 34976 3330 34978
rect 3296 34944 3330 34976
rect 3296 34874 3330 34906
rect 3296 34872 3330 34874
rect 3296 34806 3330 34834
rect 3296 34800 3330 34806
rect 3296 34738 3330 34762
rect 3296 34728 3330 34738
rect 3296 34670 3330 34690
rect 3296 34656 3330 34670
rect 3296 34602 3330 34618
rect 3296 34584 3330 34602
rect 3296 34534 3330 34546
rect 3296 34512 3330 34534
rect 3296 34466 3330 34474
rect 3296 34440 3330 34466
rect 3296 34398 3330 34402
rect 3296 34368 3330 34398
rect 3296 34296 3330 34330
rect 3296 34228 3330 34258
rect 3296 34224 3330 34228
rect 3296 34160 3330 34186
rect 3296 34152 3330 34160
rect 3296 34092 3330 34114
rect 3296 34080 3330 34092
rect 3296 34024 3330 34042
rect 3296 34008 3330 34024
rect 3296 33956 3330 33970
rect 3296 33936 3330 33956
rect 3296 33888 3330 33898
rect 3296 33864 3330 33888
rect 3296 33820 3330 33826
rect 3296 33792 3330 33820
rect 3296 33752 3330 33754
rect 3296 33720 3330 33752
rect 3296 33650 3330 33682
rect 3296 33648 3330 33650
rect 3296 33582 3330 33610
rect 3296 33576 3330 33582
rect 3296 33514 3330 33538
rect 3296 33504 3330 33514
rect 3296 33446 3330 33466
rect 3296 33432 3330 33446
rect 3296 33378 3330 33394
rect 3296 33360 3330 33378
rect 3296 33310 3330 33322
rect 3296 33288 3330 33310
rect 3296 33242 3330 33250
rect 3296 33216 3330 33242
rect 3296 33174 3330 33178
rect 3296 33144 3330 33174
rect 3296 33072 3330 33106
rect 3296 33004 3330 33034
rect 3296 33000 3330 33004
rect 3296 32936 3330 32962
rect 3296 32928 3330 32936
rect 3296 32868 3330 32890
rect 3296 32856 3330 32868
rect 3296 32800 3330 32818
rect 3296 32784 3330 32800
rect 3296 32732 3330 32746
rect 3296 32712 3330 32732
rect 3296 32664 3330 32674
rect 3296 32640 3330 32664
rect 3296 32596 3330 32602
rect 3296 32568 3330 32596
rect 3296 32528 3330 32530
rect 3296 32496 3330 32528
rect 3296 32426 3330 32458
rect 3296 32424 3330 32426
rect 3296 32358 3330 32386
rect 3296 32352 3330 32358
rect 3296 32290 3330 32314
rect 3296 32280 3330 32290
rect 3296 32222 3330 32242
rect 3296 32208 3330 32222
rect 3296 32154 3330 32170
rect 3296 32136 3330 32154
rect 3296 32086 3330 32098
rect 3296 32064 3330 32086
rect 3296 32018 3330 32026
rect 3296 31992 3330 32018
rect 3296 31950 3330 31954
rect 3296 31920 3330 31950
rect 3296 31848 3330 31882
rect 3296 31780 3330 31810
rect 3296 31776 3330 31780
rect 3296 31712 3330 31738
rect 3296 31704 3330 31712
rect 3296 31644 3330 31666
rect 3296 31632 3330 31644
rect 3296 31576 3330 31594
rect 3296 31560 3330 31576
rect 3296 31508 3330 31522
rect 3296 31488 3330 31508
rect 3296 31440 3330 31450
rect 3296 31416 3330 31440
rect 3296 31372 3330 31378
rect 3296 31344 3330 31372
rect 3296 31304 3330 31306
rect 3296 31272 3330 31304
rect 3296 31202 3330 31234
rect 3296 31200 3330 31202
rect 3296 31134 3330 31162
rect 3296 31128 3330 31134
rect 3296 31066 3330 31090
rect 3296 31056 3330 31066
rect 3296 30998 3330 31018
rect 3296 30984 3330 30998
rect 3296 30930 3330 30946
rect 3296 30912 3330 30930
rect 3296 30862 3330 30874
rect 3296 30840 3330 30862
rect 3296 30794 3330 30802
rect 3296 30768 3330 30794
rect 3296 30726 3330 30730
rect 3296 30696 3330 30726
rect 3296 30624 3330 30658
rect 3296 30556 3330 30586
rect 3296 30552 3330 30556
rect 3296 30488 3330 30514
rect 3296 30480 3330 30488
rect 3296 30420 3330 30442
rect 3296 30408 3330 30420
rect 3296 30352 3330 30370
rect 3296 30336 3330 30352
rect 3296 30284 3330 30298
rect 3296 30264 3330 30284
rect 3296 30216 3330 30226
rect 3296 30192 3330 30216
rect 3296 30148 3330 30154
rect 3296 30120 3330 30148
rect 3296 30080 3330 30082
rect 3296 30048 3330 30080
rect 3296 29978 3330 30010
rect 3296 29976 3330 29978
rect 3296 29910 3330 29938
rect 3296 29904 3330 29910
rect 3296 29842 3330 29866
rect 3296 29832 3330 29842
rect 3296 29774 3330 29794
rect 3296 29760 3330 29774
rect 3296 29706 3330 29722
rect 3296 29688 3330 29706
rect 3296 29638 3330 29650
rect 3296 29616 3330 29638
rect 3296 29570 3330 29578
rect 3296 29544 3330 29570
rect 3296 29502 3330 29506
rect 3296 29472 3330 29502
rect 3296 29400 3330 29434
rect 3296 29332 3330 29362
rect 3296 29328 3330 29332
rect 3296 29264 3330 29290
rect 3296 29256 3330 29264
rect 3296 29196 3330 29218
rect 3296 29184 3330 29196
rect 3296 29128 3330 29146
rect 3296 29112 3330 29128
rect 3296 29060 3330 29074
rect 3296 29040 3330 29060
rect 3296 28992 3330 29002
rect 3296 28968 3330 28992
rect 3296 28924 3330 28930
rect 3296 28896 3330 28924
rect 3296 28856 3330 28858
rect 3296 28824 3330 28856
rect 3296 28754 3330 28786
rect 3296 28752 3330 28754
rect 3296 28686 3330 28714
rect 3296 28680 3330 28686
rect 3296 28618 3330 28642
rect 3296 28608 3330 28618
rect 3296 28550 3330 28570
rect 3296 28536 3330 28550
rect 3296 28482 3330 28498
rect 3296 28464 3330 28482
rect 3296 28414 3330 28426
rect 3296 28392 3330 28414
rect 3296 28346 3330 28354
rect 3296 28320 3330 28346
rect 3296 28278 3330 28282
rect 3296 28248 3330 28278
rect 3296 28176 3330 28210
rect 3296 28108 3330 28138
rect 3296 28104 3330 28108
rect 3296 28040 3330 28066
rect 3296 28032 3330 28040
rect 3296 27972 3330 27994
rect 3296 27960 3330 27972
rect 3296 27904 3330 27922
rect 3296 27888 3330 27904
rect 3296 27836 3330 27850
rect 3296 27816 3330 27836
rect 3296 27768 3330 27778
rect 3296 27744 3330 27768
rect 3296 27700 3330 27706
rect 3296 27672 3330 27700
rect 3296 27632 3330 27634
rect 3296 27600 3330 27632
rect 3296 27530 3330 27562
rect 3296 27528 3330 27530
rect 3296 27462 3330 27490
rect 3296 27456 3330 27462
rect 3296 27394 3330 27418
rect 3296 27384 3330 27394
rect 3296 27326 3330 27346
rect 3296 27312 3330 27326
rect 3296 27258 3330 27274
rect 3296 27240 3330 27258
rect 3296 27190 3330 27202
rect 3296 27168 3330 27190
rect 3296 27122 3330 27130
rect 3296 27096 3330 27122
rect 3296 27054 3330 27058
rect 3296 27024 3330 27054
rect 3296 26952 3330 26986
rect 3296 26884 3330 26914
rect 3296 26880 3330 26884
rect 3296 26816 3330 26842
rect 3296 26808 3330 26816
rect 3296 26748 3330 26770
rect 3296 26736 3330 26748
rect 3296 26680 3330 26698
rect 3296 26664 3330 26680
rect 3296 26612 3330 26626
rect 3296 26592 3330 26612
rect 3296 26544 3330 26554
rect 3296 26520 3330 26544
rect 3296 26476 3330 26482
rect 3296 26448 3330 26476
rect 3296 26408 3330 26410
rect 3296 26376 3330 26408
rect 3296 26306 3330 26338
rect 3296 26304 3330 26306
rect 3296 26238 3330 26266
rect 3296 26232 3330 26238
rect 3296 26170 3330 26194
rect 3296 26160 3330 26170
rect 3296 26102 3330 26122
rect 3296 26088 3330 26102
rect 3296 26034 3330 26050
rect 3296 26016 3330 26034
rect 3296 25966 3330 25978
rect 3296 25944 3330 25966
rect 3296 25898 3330 25906
rect 3296 25872 3330 25898
rect 3296 25830 3330 25834
rect 3296 25800 3330 25830
rect 3296 25728 3330 25762
rect 3296 25660 3330 25690
rect 3296 25656 3330 25660
rect 3296 25592 3330 25618
rect 3296 25584 3330 25592
rect 3296 25524 3330 25546
rect 3296 25512 3330 25524
rect 3296 25456 3330 25474
rect 3296 25440 3330 25456
rect 3296 25388 3330 25402
rect 3296 25368 3330 25388
rect 3296 25320 3330 25330
rect 3296 25296 3330 25320
rect 3296 25252 3330 25258
rect 3296 25224 3330 25252
rect 3296 25184 3330 25186
rect 3296 25152 3330 25184
rect 3296 25082 3330 25114
rect 3296 25080 3330 25082
rect 3296 25014 3330 25042
rect 3296 25008 3330 25014
rect 3296 24946 3330 24970
rect 3296 24936 3330 24946
rect 3296 24878 3330 24898
rect 3296 24864 3330 24878
rect 3296 24810 3330 24826
rect 3296 24792 3330 24810
rect 3296 24742 3330 24754
rect 3296 24720 3330 24742
rect 3296 24674 3330 24682
rect 3296 24648 3330 24674
rect 3296 24606 3330 24610
rect 3296 24576 3330 24606
rect 3296 24504 3330 24538
rect 3296 24436 3330 24466
rect 3296 24432 3330 24436
rect 3296 24368 3330 24394
rect 3296 24360 3330 24368
rect 3296 24300 3330 24322
rect 3296 24288 3330 24300
rect 3296 24232 3330 24250
rect 3296 24216 3330 24232
rect 3296 24164 3330 24178
rect 3296 24144 3330 24164
rect 3296 24096 3330 24106
rect 3296 24072 3330 24096
rect 3296 24028 3330 24034
rect 3296 24000 3330 24028
rect 3296 23960 3330 23962
rect 3296 23928 3330 23960
rect 3296 23858 3330 23890
rect 3296 23856 3330 23858
rect 3296 23790 3330 23818
rect 3296 23784 3330 23790
rect 3296 23722 3330 23746
rect 3296 23712 3330 23722
rect 3296 23654 3330 23674
rect 3296 23640 3330 23654
rect 3296 23586 3330 23602
rect 3296 23568 3330 23586
rect 3296 23518 3330 23530
rect 3296 23496 3330 23518
rect 3296 23450 3330 23458
rect 3296 23424 3330 23450
rect 3296 23382 3330 23386
rect 3296 23352 3330 23382
rect 3296 23280 3330 23314
rect 3296 23212 3330 23242
rect 3296 23208 3330 23212
rect 3296 23144 3330 23170
rect 3296 23136 3330 23144
rect 3296 23076 3330 23098
rect 3296 23064 3330 23076
rect 3296 23008 3330 23026
rect 3296 22992 3330 23008
rect 3296 22940 3330 22954
rect 3296 22920 3330 22940
rect 3296 22872 3330 22882
rect 3296 22848 3330 22872
rect 3296 22804 3330 22810
rect 3296 22776 3330 22804
rect 3296 22736 3330 22738
rect 3296 22704 3330 22736
rect 3296 22634 3330 22666
rect 3296 22632 3330 22634
rect 3296 22566 3330 22594
rect 3296 22560 3330 22566
rect 3296 22498 3330 22522
rect 3296 22488 3330 22498
rect 3296 22430 3330 22450
rect 3296 22416 3330 22430
rect 3296 22362 3330 22378
rect 3296 22344 3330 22362
rect 3296 22294 3330 22306
rect 3296 22272 3330 22294
rect 3296 22226 3330 22234
rect 3296 22200 3330 22226
rect 3296 22158 3330 22162
rect 3296 22128 3330 22158
rect 3296 22056 3330 22090
rect 3296 21988 3330 22018
rect 3296 21984 3330 21988
rect 3296 21920 3330 21946
rect 3296 21912 3330 21920
rect 3296 21852 3330 21874
rect 3296 21840 3330 21852
rect 3296 21784 3330 21802
rect 3296 21768 3330 21784
rect 3296 21716 3330 21730
rect 3296 21696 3330 21716
rect 3296 21648 3330 21658
rect 3296 21624 3330 21648
rect 3296 21580 3330 21586
rect 3296 21552 3330 21580
rect 3296 21512 3330 21514
rect 3296 21480 3330 21512
rect 3296 21410 3330 21442
rect 3296 21408 3330 21410
rect 3296 21342 3330 21370
rect 3296 21336 3330 21342
rect 3296 21274 3330 21298
rect 3296 21264 3330 21274
rect 3296 21206 3330 21226
rect 3296 21192 3330 21206
rect 3296 21138 3330 21154
rect 3296 21120 3330 21138
rect 3296 21070 3330 21082
rect 3296 21048 3330 21070
rect 3296 21002 3330 21010
rect 3296 20976 3330 21002
rect 3296 20934 3330 20938
rect 3296 20904 3330 20934
rect 3296 20832 3330 20866
rect 3296 20764 3330 20794
rect 3296 20760 3330 20764
rect 3296 20696 3330 20722
rect 3296 20688 3330 20696
rect 3296 20628 3330 20650
rect 3296 20616 3330 20628
rect 3296 20560 3330 20578
rect 3296 20544 3330 20560
rect 3296 20492 3330 20506
rect 3296 20472 3330 20492
rect 3296 20424 3330 20434
rect 3296 20400 3330 20424
rect 3296 20356 3330 20362
rect 3296 20328 3330 20356
rect 3296 20288 3330 20290
rect 3296 20256 3330 20288
rect 3296 20186 3330 20218
rect 3296 20184 3330 20186
rect 3296 20118 3330 20146
rect 3296 20112 3330 20118
rect 3296 20050 3330 20074
rect 3296 20040 3330 20050
rect 3296 19982 3330 20002
rect 3296 19968 3330 19982
rect 3296 19914 3330 19930
rect 3296 19896 3330 19914
rect 3296 19846 3330 19858
rect 3296 19824 3330 19846
rect 3296 19778 3330 19786
rect 3296 19752 3330 19778
rect 3296 19710 3330 19714
rect 3296 19680 3330 19710
rect 3296 19608 3330 19642
rect 3296 19540 3330 19570
rect 3296 19536 3330 19540
rect 3296 19472 3330 19498
rect 3296 19464 3330 19472
rect 3296 19404 3330 19426
rect 3296 19392 3330 19404
rect 3296 19336 3330 19354
rect 3296 19320 3330 19336
rect 3296 19268 3330 19282
rect 3296 19248 3330 19268
rect 3296 19200 3330 19210
rect 3296 19176 3330 19200
rect 3296 19132 3330 19138
rect 3296 19104 3330 19132
rect 3296 19064 3330 19066
rect 3296 19032 3330 19064
rect 3296 18962 3330 18994
rect 3296 18960 3330 18962
rect 3296 18894 3330 18922
rect 3296 18888 3330 18894
rect 3296 18826 3330 18850
rect 3296 18816 3330 18826
rect 3296 18758 3330 18778
rect 3296 18744 3330 18758
rect 3296 18690 3330 18706
rect 3296 18672 3330 18690
rect 3296 18622 3330 18634
rect 3296 18600 3330 18622
rect 3296 18554 3330 18562
rect 3296 18528 3330 18554
rect 3296 18486 3330 18490
rect 3296 18456 3330 18486
rect 3296 18384 3330 18418
rect 3296 18316 3330 18346
rect 3296 18312 3330 18316
rect 3296 18248 3330 18274
rect 3296 18240 3330 18248
rect 3296 18180 3330 18202
rect 3296 18168 3330 18180
rect 3296 18112 3330 18130
rect 3296 18096 3330 18112
rect 3296 18044 3330 18058
rect 3296 18024 3330 18044
rect 3296 17976 3330 17986
rect 3296 17952 3330 17976
rect 3296 17908 3330 17914
rect 3296 17880 3330 17908
rect 3296 17840 3330 17842
rect 3296 17808 3330 17840
rect 3296 17738 3330 17770
rect 3296 17736 3330 17738
rect 3296 17670 3330 17698
rect 3296 17664 3330 17670
rect 3296 17602 3330 17626
rect 3296 17592 3330 17602
rect 3296 17534 3330 17554
rect 3296 17520 3330 17534
rect 3296 17466 3330 17482
rect 3296 17448 3330 17466
rect 3296 17398 3330 17410
rect 3296 17376 3330 17398
rect 3296 17330 3330 17338
rect 3296 17304 3330 17330
rect 3296 17262 3330 17266
rect 3296 17232 3330 17262
rect 3296 17160 3330 17194
rect 3296 17092 3330 17122
rect 3296 17088 3330 17092
rect 3296 17024 3330 17050
rect 3296 17016 3330 17024
rect 3296 16956 3330 16978
rect 3296 16944 3330 16956
rect 3296 16888 3330 16906
rect 3296 16872 3330 16888
rect 3296 16820 3330 16834
rect 3296 16800 3330 16820
rect 3296 16752 3330 16762
rect 3296 16728 3330 16752
rect 3296 16684 3330 16690
rect 3296 16656 3330 16684
rect 3296 16616 3330 16618
rect 3296 16584 3330 16616
rect 3296 16514 3330 16546
rect 3296 16512 3330 16514
rect 3296 16446 3330 16474
rect 3296 16440 3330 16446
rect 3296 16378 3330 16402
rect 3296 16368 3330 16378
rect 3296 16310 3330 16330
rect 3296 16296 3330 16310
rect 3296 16242 3330 16258
rect 3296 16224 3330 16242
rect 3296 16174 3330 16186
rect 3296 16152 3330 16174
rect 3296 16106 3330 16114
rect 3296 16080 3330 16106
rect 3296 16038 3330 16042
rect 3296 16008 3330 16038
rect 3296 15936 3330 15970
rect 3296 15868 3330 15898
rect 3296 15864 3330 15868
rect 3296 15800 3330 15826
rect 3296 15792 3330 15800
rect 3296 15732 3330 15754
rect 3296 15720 3330 15732
rect 3296 15664 3330 15682
rect 3296 15648 3330 15664
rect 3296 15596 3330 15610
rect 3296 15576 3330 15596
rect 3296 15528 3330 15538
rect 3296 15504 3330 15528
rect 3296 15460 3330 15466
rect 3296 15432 3330 15460
rect 3296 15392 3330 15394
rect 3296 15360 3330 15392
rect 3296 15290 3330 15322
rect 3296 15288 3330 15290
rect 3296 15222 3330 15250
rect 3296 15216 3330 15222
rect 3296 15154 3330 15178
rect 3296 15144 3330 15154
rect 3296 15086 3330 15106
rect 3296 15072 3330 15086
rect 3296 15018 3330 15034
rect 3296 15000 3330 15018
rect 3296 14950 3330 14962
rect 3296 14928 3330 14950
rect 3296 14882 3330 14890
rect 3296 14856 3330 14882
rect 3296 14814 3330 14818
rect 3296 14784 3330 14814
rect 3296 14712 3330 14746
rect 3296 14644 3330 14674
rect 3296 14640 3330 14644
rect 3296 14576 3330 14602
rect 3296 14568 3330 14576
rect 3296 14508 3330 14530
rect 3296 14496 3330 14508
rect 3296 14440 3330 14458
rect 3296 14424 3330 14440
rect 3296 14372 3330 14386
rect 3296 14352 3330 14372
rect 3296 14304 3330 14314
rect 3296 14280 3330 14304
rect 3296 14236 3330 14242
rect 3296 14208 3330 14236
rect 3296 14168 3330 14170
rect 3296 14136 3330 14168
rect 3296 14066 3330 14098
rect 3296 14064 3330 14066
rect 3296 13998 3330 14026
rect 3296 13992 3330 13998
rect 3296 13930 3330 13954
rect 3296 13920 3330 13930
rect 3296 13862 3330 13882
rect 3296 13848 3330 13862
rect 3296 13794 3330 13810
rect 3296 13776 3330 13794
rect 3296 13726 3330 13738
rect 3296 13704 3330 13726
rect 3296 13658 3330 13666
rect 3296 13632 3330 13658
rect 3296 13590 3330 13594
rect 3296 13560 3330 13590
rect 3296 13488 3330 13522
rect 3296 13420 3330 13450
rect 3296 13416 3330 13420
rect 3296 13352 3330 13378
rect 3296 13344 3330 13352
rect 3296 13284 3330 13306
rect 3296 13272 3330 13284
rect 3296 13216 3330 13234
rect 3296 13200 3330 13216
rect 3296 13148 3330 13162
rect 3296 13128 3330 13148
rect 3296 13080 3330 13090
rect 3296 13056 3330 13080
rect 3296 13012 3330 13018
rect 3296 12984 3330 13012
rect 3296 12944 3330 12946
rect 3296 12912 3330 12944
rect 3296 12842 3330 12874
rect 3296 12840 3330 12842
rect 3296 12774 3330 12802
rect 3296 12768 3330 12774
rect 3296 12706 3330 12730
rect 3296 12696 3330 12706
rect 3296 12638 3330 12658
rect 3296 12624 3330 12638
rect 3296 12570 3330 12586
rect 3296 12552 3330 12570
rect 3296 12502 3330 12514
rect 3296 12480 3330 12502
rect 3296 12434 3330 12442
rect 3296 12408 3330 12434
rect 3296 12366 3330 12370
rect 3296 12336 3330 12366
rect 3296 12264 3330 12298
rect 3296 12196 3330 12226
rect 3296 12192 3330 12196
rect 3296 12128 3330 12154
rect 3296 12120 3330 12128
rect 3296 12060 3330 12082
rect 3296 12048 3330 12060
rect 3296 11992 3330 12010
rect 3296 11976 3330 11992
rect 3296 11924 3330 11938
rect 3296 11904 3330 11924
rect 3296 11856 3330 11866
rect 3296 11832 3330 11856
rect 3296 11788 3330 11794
rect 3296 11760 3330 11788
rect 3296 11720 3330 11722
rect 3296 11688 3330 11720
rect 3296 11618 3330 11650
rect 3296 11616 3330 11618
rect 3296 11550 3330 11578
rect 3296 11544 3330 11550
rect 3296 11482 3330 11506
rect 3296 11472 3330 11482
rect 3296 11414 3330 11434
rect 3296 11400 3330 11414
rect 3296 11346 3330 11362
rect 3296 11328 3330 11346
rect 3296 11278 3330 11290
rect 3296 11256 3330 11278
rect 3296 11210 3330 11218
rect 3296 11184 3330 11210
rect 3296 11142 3330 11146
rect 3296 11112 3330 11142
rect 3296 11040 3330 11074
rect 3296 10972 3330 11002
rect 3296 10968 3330 10972
rect 3296 10904 3330 10930
rect 3296 10896 3330 10904
rect 3296 10836 3330 10858
rect 3296 10824 3330 10836
rect 3296 10768 3330 10786
rect 3296 10752 3330 10768
rect 3296 10700 3330 10714
rect 3296 10680 3330 10700
rect 3296 10632 3330 10642
rect 3296 10608 3330 10632
rect 3296 10564 3330 10570
rect 3296 10536 3330 10564
rect 3296 10496 3330 10498
rect 3296 10464 3330 10496
rect 3296 10394 3330 10426
rect 3296 10392 3330 10394
rect 3296 10326 3330 10354
rect 3296 10320 3330 10326
rect 3296 10258 3330 10282
rect 3296 10248 3330 10258
rect 3296 10190 3330 10210
rect 3296 10176 3330 10190
rect 3296 10122 3330 10138
rect 3296 10104 3330 10122
rect 3296 10054 3330 10066
rect 3296 10032 3330 10054
rect 3296 9986 3330 9994
rect 3296 9960 3330 9986
rect 3296 9918 3330 9922
rect 3296 9888 3330 9918
rect 3296 9816 3330 9850
rect 3296 9748 3330 9778
rect 3296 9744 3330 9748
rect 3296 9680 3330 9706
rect 3296 9672 3330 9680
rect 3296 9612 3330 9634
rect 3296 9600 3330 9612
rect 3296 9544 3330 9562
rect 3296 9528 3330 9544
rect 3296 9476 3330 9490
rect 3296 9456 3330 9476
rect 3296 9408 3330 9418
rect 3296 9384 3330 9408
rect 3296 9340 3330 9346
rect 3296 9312 3330 9340
rect 3296 9272 3330 9274
rect 3296 9240 3330 9272
rect 3296 9170 3330 9202
rect 3296 9168 3330 9170
rect 3296 9102 3330 9130
rect 3296 9096 3330 9102
rect 3296 9034 3330 9058
rect 3296 9024 3330 9034
rect 3296 8966 3330 8986
rect 3296 8952 3330 8966
rect 3296 8898 3330 8914
rect 3296 8880 3330 8898
rect 3296 8830 3330 8842
rect 3296 8808 3330 8830
rect 3296 8762 3330 8770
rect 3296 8736 3330 8762
rect 3296 8694 3330 8698
rect 3296 8664 3330 8694
rect 3296 8592 3330 8626
rect 3296 8524 3330 8554
rect 3296 8520 3330 8524
rect 3296 8456 3330 8482
rect 3296 8448 3330 8456
rect 3296 8388 3330 8410
rect 3296 8376 3330 8388
rect 3296 8320 3330 8338
rect 3296 8304 3330 8320
rect 3296 8252 3330 8266
rect 3296 8232 3330 8252
rect 3296 8184 3330 8194
rect 3296 8160 3330 8184
rect 3296 8116 3330 8122
rect 3296 8088 3330 8116
rect 3296 8048 3330 8050
rect 3296 8016 3330 8048
rect 3296 7946 3330 7978
rect 3296 7944 3330 7946
rect 3296 7878 3330 7906
rect 3296 7872 3330 7878
rect 3296 7810 3330 7834
rect 3296 7800 3330 7810
rect 3296 7742 3330 7762
rect 3296 7728 3330 7742
rect 3296 7674 3330 7690
rect 3296 7656 3330 7674
rect 3296 7606 3330 7618
rect 3296 7584 3330 7606
rect 3296 7538 3330 7546
rect 3296 7512 3330 7538
rect 3296 7470 3330 7474
rect 3296 7440 3330 7470
rect 3296 7368 3330 7402
rect 3296 7300 3330 7330
rect 3296 7296 3330 7300
rect 3296 7232 3330 7258
rect 3296 7224 3330 7232
rect 3296 7164 3330 7186
rect 3296 7152 3330 7164
rect 3296 7096 3330 7114
rect 3296 7080 3330 7096
rect 3296 7028 3330 7042
rect 3296 7008 3330 7028
rect 3296 6960 3330 6970
rect 3296 6936 3330 6960
rect 3296 6892 3330 6898
rect 3296 6864 3330 6892
rect 3296 6824 3330 6826
rect 3296 6792 3330 6824
rect 3296 6722 3330 6754
rect 3296 6720 3330 6722
rect 3296 6654 3330 6682
rect 3296 6648 3330 6654
rect 3296 6586 3330 6610
rect 3296 6576 3330 6586
rect 3296 6518 3330 6538
rect 3296 6504 3330 6518
rect 3296 6450 3330 6466
rect 3296 6432 3330 6450
rect 3296 6382 3330 6394
rect 3296 6360 3330 6382
rect 3296 6314 3330 6322
rect 3296 6288 3330 6314
rect 3296 6246 3330 6250
rect 3296 6216 3330 6246
rect 3296 6144 3330 6178
rect 3296 6076 3330 6106
rect 3296 6072 3330 6076
rect 3296 6008 3330 6034
rect 3296 6000 3330 6008
rect 3296 5940 3330 5962
rect 3296 5928 3330 5940
rect 3296 5872 3330 5890
rect 3296 5856 3330 5872
rect 3296 5804 3330 5818
rect 3296 5784 3330 5804
rect 3296 5736 3330 5746
rect 3296 5712 3330 5736
rect 3296 5668 3330 5674
rect 3296 5640 3330 5668
rect 3296 5600 3330 5602
rect 3296 5568 3330 5600
rect 3296 5498 3330 5530
rect 3296 5496 3330 5498
rect 3296 5430 3330 5458
rect 3296 5424 3330 5430
rect 3296 5362 3330 5386
rect 3296 5352 3330 5362
rect 3296 5294 3330 5314
rect 3296 5280 3330 5294
rect 3296 5226 3330 5242
rect 3296 5208 3330 5226
rect 3296 5158 3330 5170
rect 3296 5136 3330 5158
rect 3296 5090 3330 5098
rect 3296 5064 3330 5090
rect 3296 5022 3330 5026
rect 3296 4992 3330 5022
rect 3296 4920 3330 4954
rect 3296 4852 3330 4882
rect 3296 4848 3330 4852
rect 3296 4784 3330 4810
rect 3296 4776 3330 4784
rect 3296 4716 3330 4738
rect 3296 4704 3330 4716
rect 3296 4648 3330 4666
rect 3296 4632 3330 4648
rect 3296 4580 3330 4594
rect 3296 4560 3330 4580
rect 3296 4512 3330 4522
rect 3296 4488 3330 4512
rect 3296 4444 3330 4450
rect 3296 4416 3330 4444
rect 3296 4376 3330 4378
rect 3296 4344 3330 4376
rect 3296 4274 3330 4306
rect 3296 4272 3330 4274
rect 3296 4206 3330 4234
rect 3296 4200 3330 4206
rect 3296 4138 3330 4162
rect 3296 4128 3330 4138
rect 3296 4070 3330 4090
rect 3296 4056 3330 4070
rect 3296 4002 3330 4018
rect 3296 3984 3330 4002
rect 3296 3934 3330 3946
rect 3296 3912 3330 3934
rect 3296 3866 3330 3874
rect 3296 3840 3330 3866
rect 3296 3798 3330 3802
rect 3296 3768 3330 3798
rect 3296 3696 3330 3730
rect 3296 3628 3330 3658
rect 3296 3624 3330 3628
rect 3296 3560 3330 3586
rect 3296 3552 3330 3560
rect 3296 3492 3330 3514
rect 3296 3480 3330 3492
rect 3296 3424 3330 3442
rect 3296 3408 3330 3424
rect 3296 3356 3330 3370
rect 3296 3336 3330 3356
rect 3296 3288 3330 3298
rect 3296 3264 3330 3288
rect 3296 3220 3330 3225
rect 3296 3191 3330 3220
rect 3296 3118 3330 3152
rect 3296 3050 3330 3079
rect 3296 3045 3330 3050
rect 3296 2982 3330 3006
rect 3296 2972 3330 2982
rect 3296 2914 3330 2933
rect 3296 2899 3330 2914
rect 3296 2846 3330 2860
rect 3296 2826 3330 2846
rect 3296 2778 3330 2787
rect 3296 2753 3330 2778
rect 3296 2710 3330 2714
rect 3296 2680 3330 2710
rect 3296 2608 3330 2641
rect 3296 2607 3330 2608
rect 3296 2540 3330 2568
rect 3296 2534 3330 2540
rect 3296 2472 3330 2495
rect 3296 2461 3330 2472
rect 3296 2404 3330 2422
rect 3296 2388 3330 2404
rect 3296 2336 3330 2349
rect 3296 2315 3330 2336
rect 3296 2268 3330 2276
rect 3296 2242 3330 2268
rect 3296 2200 3330 2203
rect 3296 2169 3330 2200
rect 3296 2098 3330 2130
rect 3296 2096 3330 2098
rect 3296 2030 3330 2057
rect 3296 2023 3330 2030
rect 3296 1962 3330 1984
rect 3296 1950 3330 1962
rect 3296 1894 3330 1911
rect 3296 1877 3330 1894
rect 3296 1826 3330 1838
rect 3296 1804 3330 1826
rect 3296 1758 3330 1765
rect 3296 1731 3330 1758
rect 3296 1690 3330 1692
rect 3296 1658 3330 1690
rect 3296 1588 3330 1619
rect 3296 1585 3330 1588
rect 3296 1520 3330 1546
rect 3296 1512 3330 1520
rect 3296 1452 3330 1473
rect 3296 1439 3330 1452
rect 3296 1384 3330 1400
rect 3296 1366 3330 1384
rect 3296 1316 3330 1327
rect 3296 1293 3330 1316
rect 3296 1248 3330 1254
rect 3296 1220 3330 1248
rect 3296 1180 3330 1181
rect 3296 1147 3330 1180
rect 3296 1078 3330 1108
rect 3296 1074 3330 1078
rect 3296 1010 3330 1035
rect 3296 1001 3330 1010
rect 3296 942 3330 962
rect 3296 928 3330 942
rect 3296 874 3330 889
rect 3296 855 3330 874
rect 3296 806 3330 816
rect 3296 782 3330 806
rect 3296 738 3330 743
rect 3296 709 3330 738
rect 3296 636 3330 670
rect 3296 568 3330 597
rect 3296 563 3330 568
rect 126 502 160 520
rect 126 486 160 502
rect 126 434 160 448
rect 126 414 160 434
rect 126 366 160 376
rect 126 342 160 366
rect 126 270 160 304
rect 126 218 160 232
rect 126 198 160 218
rect 3296 500 3330 524
rect 3296 490 3330 500
rect 3296 432 3330 451
rect 3296 417 3330 432
rect 3296 364 3330 378
rect 3296 344 3330 364
rect 3296 296 3330 305
rect 3296 271 3330 296
rect 3296 228 3330 232
rect 3296 198 3330 228
rect 198 126 228 160
rect 228 126 232 160
rect 271 126 296 160
rect 296 126 305 160
rect 344 126 364 160
rect 364 126 378 160
rect 416 126 432 160
rect 432 126 450 160
rect 488 126 500 160
rect 500 126 522 160
rect 560 126 568 160
rect 568 126 594 160
rect 632 126 636 160
rect 636 126 666 160
rect 704 126 738 160
rect 776 126 806 160
rect 806 126 810 160
rect 848 126 874 160
rect 874 126 882 160
rect 920 126 942 160
rect 942 126 954 160
rect 992 126 1010 160
rect 1010 126 1026 160
rect 1064 126 1078 160
rect 1078 126 1098 160
rect 1136 126 1146 160
rect 1146 126 1170 160
rect 1208 126 1214 160
rect 1214 126 1242 160
rect 1280 126 1282 160
rect 1282 126 1314 160
rect 1352 126 1384 160
rect 1384 126 1386 160
rect 1424 126 1452 160
rect 1452 126 1458 160
rect 1496 126 1520 160
rect 1520 126 1530 160
rect 1568 126 1588 160
rect 1588 126 1602 160
rect 1640 126 1656 160
rect 1656 126 1674 160
rect 1712 126 1724 160
rect 1724 126 1746 160
rect 1784 126 1792 160
rect 1792 126 1818 160
rect 1856 126 1860 160
rect 1860 126 1890 160
rect 1928 126 1962 160
rect 2000 126 2030 160
rect 2030 126 2034 160
rect 2072 126 2098 160
rect 2098 126 2106 160
rect 2144 126 2166 160
rect 2166 126 2178 160
rect 2216 126 2234 160
rect 2234 126 2250 160
rect 2288 126 2302 160
rect 2302 126 2322 160
rect 2360 126 2370 160
rect 2370 126 2394 160
rect 2432 126 2438 160
rect 2438 126 2466 160
rect 2504 126 2506 160
rect 2506 126 2538 160
rect 2576 126 2608 160
rect 2608 126 2610 160
rect 2648 126 2676 160
rect 2676 126 2682 160
rect 2720 126 2744 160
rect 2744 126 2754 160
rect 2792 126 2812 160
rect 2812 126 2826 160
rect 2864 126 2880 160
rect 2880 126 2898 160
rect 2936 126 2948 160
rect 2948 126 2970 160
rect 3008 126 3016 160
rect 3016 126 3042 160
rect 3080 126 3084 160
rect 3084 126 3114 160
rect 3152 126 3186 160
rect 3224 126 3258 160
<< metal1 >>
rect 117 39874 3339 39880
rect 117 39840 206 39874
rect 240 39840 286 39874
rect 320 39840 366 39874
rect 400 39840 447 39874
rect 481 39840 528 39874
rect 562 39840 609 39874
rect 643 39840 690 39874
rect 724 39840 800 39874
rect 834 39840 873 39874
rect 907 39840 946 39874
rect 980 39840 1019 39874
rect 1053 39840 1092 39874
rect 1126 39840 1165 39874
rect 1199 39840 1238 39874
rect 1272 39840 1311 39874
rect 1345 39840 1384 39874
rect 1418 39840 1457 39874
rect 1491 39840 1530 39874
rect 1564 39840 1603 39874
rect 1637 39840 1676 39874
rect 1710 39840 1749 39874
rect 1783 39840 1822 39874
rect 1856 39840 1895 39874
rect 1929 39840 1968 39874
rect 2002 39840 2041 39874
rect 2075 39840 2114 39874
rect 2148 39840 2188 39874
rect 2222 39840 2262 39874
rect 2296 39840 2336 39874
rect 2370 39840 2410 39874
rect 2444 39840 2484 39874
rect 2518 39840 2558 39874
rect 2592 39840 2632 39874
rect 2666 39840 2706 39874
rect 2740 39840 2780 39874
rect 2814 39840 2854 39874
rect 2888 39840 2928 39874
rect 2962 39840 3002 39874
rect 3036 39840 3076 39874
rect 3110 39840 3150 39874
rect 3184 39840 3224 39874
rect 3258 39840 3339 39874
rect 117 39834 3339 39840
rect 117 39802 171 39834
tri 171 39802 203 39834 nw
tri 3253 39802 3285 39834 ne
rect 3285 39802 3339 39834
rect 117 39768 126 39802
rect 160 39768 169 39802
tri 169 39800 171 39802 nw
tri 3285 39800 3287 39802 ne
rect 117 39729 169 39768
rect 117 39695 126 39729
rect 160 39695 169 39729
rect 117 39656 169 39695
rect 117 39622 126 39656
rect 160 39622 169 39656
rect 117 39583 169 39622
rect 117 39549 126 39583
rect 160 39549 169 39583
rect 117 39510 169 39549
rect 117 39476 126 39510
rect 160 39476 169 39510
rect 117 39437 169 39476
rect 117 39403 126 39437
rect 160 39403 169 39437
rect 117 39364 169 39403
rect 117 39330 126 39364
rect 160 39330 169 39364
rect 117 39291 169 39330
rect 117 39257 126 39291
rect 160 39257 169 39291
rect 117 39218 169 39257
rect 117 39184 126 39218
rect 160 39184 169 39218
rect 3287 39768 3296 39802
rect 3330 39768 3339 39802
rect 3287 39730 3339 39768
rect 3287 39696 3296 39730
rect 3330 39696 3339 39730
rect 3287 39658 3339 39696
rect 3287 39624 3296 39658
rect 3330 39624 3339 39658
rect 3287 39586 3339 39624
rect 3287 39552 3296 39586
rect 3330 39552 3339 39586
rect 3287 39514 3339 39552
rect 3287 39480 3296 39514
rect 3330 39480 3339 39514
rect 3287 39442 3339 39480
rect 3287 39408 3296 39442
rect 3330 39408 3339 39442
rect 3287 39370 3339 39408
rect 3287 39336 3296 39370
rect 3330 39336 3339 39370
rect 3287 39298 3339 39336
rect 3287 39264 3296 39298
rect 3330 39264 3339 39298
rect 3287 39226 3339 39264
rect 3287 39192 3296 39226
rect 3330 39192 3339 39226
rect 117 39145 169 39184
rect 117 39111 126 39145
rect 160 39111 169 39145
rect 117 39072 169 39111
rect 117 39038 126 39072
rect 160 39038 169 39072
rect 117 38999 169 39038
rect 117 38965 126 38999
rect 160 38965 169 38999
rect 117 38926 169 38965
rect 117 38892 126 38926
rect 160 38892 169 38926
rect 117 38853 169 38892
rect 117 38819 126 38853
rect 160 38819 169 38853
rect 117 38780 169 38819
rect 117 38746 126 38780
rect 160 38746 169 38780
rect 117 38707 169 38746
rect 117 38673 126 38707
rect 160 38673 169 38707
rect 117 38634 169 38673
rect 117 38600 126 38634
rect 160 38600 169 38634
rect 117 38561 169 38600
rect 117 38527 126 38561
rect 160 38527 169 38561
rect 117 38488 169 38527
rect 117 38454 126 38488
rect 160 38454 169 38488
rect 117 38415 169 38454
rect 117 38381 126 38415
rect 160 38381 169 38415
rect 117 38342 169 38381
rect 117 38308 126 38342
rect 160 38308 169 38342
rect 117 38269 169 38308
rect 117 38235 126 38269
rect 160 38235 169 38269
rect 117 38196 169 38235
rect 117 38162 126 38196
rect 160 38162 169 38196
rect 117 38123 169 38162
rect 117 38089 126 38123
rect 160 38089 169 38123
rect 117 38050 169 38089
rect 117 38016 126 38050
rect 160 38016 169 38050
rect 117 37977 169 38016
rect 117 37943 126 37977
rect 160 37943 169 37977
rect 117 37904 169 37943
rect 117 37870 126 37904
rect 160 37870 169 37904
rect 117 37831 169 37870
rect 117 37797 126 37831
rect 160 37797 169 37831
rect 117 37758 169 37797
rect 117 37724 126 37758
rect 160 37724 169 37758
rect 117 37685 169 37724
rect 117 37651 126 37685
rect 160 37651 169 37685
rect 117 37612 169 37651
rect 117 37578 126 37612
rect 160 37578 169 37612
rect 117 37539 169 37578
rect 117 37505 126 37539
rect 160 37505 169 37539
rect 117 37466 169 37505
rect 117 37432 126 37466
rect 160 37432 169 37466
rect 117 37393 169 37432
rect 117 37359 126 37393
rect 160 37359 169 37393
rect 117 37320 169 37359
rect 117 37286 126 37320
rect 160 37286 169 37320
rect 117 37247 169 37286
rect 117 37213 126 37247
rect 160 37213 169 37247
rect 117 37174 169 37213
rect 117 37140 126 37174
rect 160 37140 169 37174
rect 117 37101 169 37140
rect 117 37067 126 37101
rect 160 37067 169 37101
rect 117 37028 169 37067
rect 117 36994 126 37028
rect 160 36994 169 37028
rect 117 36955 169 36994
rect 117 36921 126 36955
rect 160 36921 169 36955
rect 117 36882 169 36921
rect 117 36848 126 36882
rect 160 36848 169 36882
rect 117 36809 169 36848
rect 117 36775 126 36809
rect 160 36775 169 36809
rect 117 36736 169 36775
rect 117 36702 126 36736
rect 160 36702 169 36736
rect 117 36664 169 36702
rect 117 36630 126 36664
rect 160 36630 169 36664
rect 117 36592 169 36630
rect 117 36558 126 36592
rect 160 36558 169 36592
rect 117 36520 169 36558
rect 117 36486 126 36520
rect 160 36486 169 36520
rect 117 36448 169 36486
rect 117 36414 126 36448
rect 160 36414 169 36448
rect 117 36376 169 36414
rect 117 36342 126 36376
rect 160 36342 169 36376
rect 117 36304 169 36342
rect 117 36270 126 36304
rect 160 36270 169 36304
rect 117 36232 169 36270
rect 117 36198 126 36232
rect 160 36198 169 36232
rect 117 36160 169 36198
rect 117 36126 126 36160
rect 160 36126 169 36160
rect 117 36088 169 36126
rect 117 36054 126 36088
rect 160 36054 169 36088
rect 117 36016 169 36054
rect 117 35982 126 36016
rect 160 35982 169 36016
rect 117 35944 169 35982
rect 117 35910 126 35944
rect 160 35910 169 35944
rect 117 35872 169 35910
rect 117 35838 126 35872
rect 160 35838 169 35872
rect 117 35800 169 35838
rect 117 35766 126 35800
rect 160 35766 169 35800
rect 117 35728 169 35766
rect 117 35694 126 35728
rect 160 35694 169 35728
rect 117 35656 169 35694
rect 117 35622 126 35656
rect 160 35622 169 35656
rect 117 35584 169 35622
rect 117 35550 126 35584
rect 160 35550 169 35584
rect 117 35512 169 35550
rect 117 35478 126 35512
rect 160 35478 169 35512
rect 117 35440 169 35478
rect 117 35406 126 35440
rect 160 35406 169 35440
rect 117 35368 169 35406
rect 117 35334 126 35368
rect 160 35334 169 35368
rect 117 35296 169 35334
rect 117 35262 126 35296
rect 160 35262 169 35296
rect 117 35224 169 35262
rect 117 35190 126 35224
rect 160 35190 169 35224
rect 117 35152 169 35190
rect 117 35118 126 35152
rect 160 35118 169 35152
rect 117 35080 169 35118
rect 117 35046 126 35080
rect 160 35046 169 35080
rect 117 35008 169 35046
rect 117 34974 126 35008
rect 160 34974 169 35008
rect 117 34936 169 34974
rect 117 34902 126 34936
rect 160 34902 169 34936
rect 117 34864 169 34902
rect 117 34830 126 34864
rect 160 34830 169 34864
rect 117 34792 169 34830
rect 117 34758 126 34792
rect 160 34758 169 34792
rect 117 34720 169 34758
rect 117 34686 126 34720
rect 160 34686 169 34720
rect 117 34648 169 34686
rect 117 34614 126 34648
rect 160 34614 169 34648
rect 117 34576 169 34614
rect 117 34542 126 34576
rect 160 34542 169 34576
rect 117 34504 169 34542
rect 117 34470 126 34504
rect 160 34470 169 34504
rect 117 34432 169 34470
rect 117 34398 126 34432
rect 160 34398 169 34432
rect 117 34360 169 34398
rect 117 34326 126 34360
rect 160 34326 169 34360
rect 117 34288 169 34326
rect 117 34254 126 34288
rect 160 34254 169 34288
rect 117 34216 169 34254
rect 117 34182 126 34216
rect 160 34182 169 34216
rect 117 34144 169 34182
rect 117 34110 126 34144
rect 160 34110 169 34144
rect 117 34072 169 34110
rect 117 34038 126 34072
rect 160 34038 169 34072
rect 117 34000 169 34038
rect 117 33966 126 34000
rect 160 33966 169 34000
rect 117 33928 169 33966
rect 117 33894 126 33928
rect 160 33894 169 33928
rect 117 33856 169 33894
rect 117 33822 126 33856
rect 160 33822 169 33856
rect 117 33784 169 33822
rect 117 33750 126 33784
rect 160 33750 169 33784
rect 117 33712 169 33750
rect 117 33678 126 33712
rect 160 33678 169 33712
rect 117 33640 169 33678
rect 117 33606 126 33640
rect 160 33606 169 33640
rect 117 33568 169 33606
rect 117 33534 126 33568
rect 160 33534 169 33568
rect 117 33496 169 33534
rect 117 33462 126 33496
rect 160 33462 169 33496
rect 117 33424 169 33462
rect 117 33390 126 33424
rect 160 33390 169 33424
rect 117 33352 169 33390
rect 117 33318 126 33352
rect 160 33318 169 33352
rect 117 33280 169 33318
rect 117 33246 126 33280
rect 160 33246 169 33280
rect 117 33208 169 33246
rect 117 33174 126 33208
rect 160 33174 169 33208
rect 117 33136 169 33174
rect 117 33102 126 33136
rect 160 33102 169 33136
rect 117 33064 169 33102
rect 117 33030 126 33064
rect 160 33030 169 33064
rect 117 32992 169 33030
rect 117 32958 126 32992
rect 160 32958 169 32992
rect 117 32920 169 32958
rect 117 32886 126 32920
rect 160 32886 169 32920
rect 117 32848 169 32886
rect 117 32814 126 32848
rect 160 32814 169 32848
rect 117 32776 169 32814
rect 117 32742 126 32776
rect 160 32742 169 32776
rect 117 32704 169 32742
rect 117 32670 126 32704
rect 160 32670 169 32704
rect 117 32632 169 32670
rect 117 32598 126 32632
rect 160 32598 169 32632
rect 117 32560 169 32598
rect 117 32526 126 32560
rect 160 32526 169 32560
rect 117 32488 169 32526
rect 117 32454 126 32488
rect 160 32454 169 32488
rect 117 32416 169 32454
rect 117 32382 126 32416
rect 160 32382 169 32416
rect 117 32344 169 32382
rect 117 32310 126 32344
rect 160 32310 169 32344
rect 117 32272 169 32310
rect 117 32238 126 32272
rect 160 32238 169 32272
rect 117 32200 169 32238
rect 117 32166 126 32200
rect 160 32166 169 32200
rect 117 32128 169 32166
rect 117 32094 126 32128
rect 160 32094 169 32128
rect 117 32056 169 32094
rect 117 32022 126 32056
rect 160 32022 169 32056
rect 117 31984 169 32022
rect 117 31950 126 31984
rect 160 31950 169 31984
rect 117 31912 169 31950
rect 117 31878 126 31912
rect 160 31878 169 31912
rect 117 31840 169 31878
rect 117 31806 126 31840
rect 160 31806 169 31840
rect 117 31768 169 31806
rect 117 31734 126 31768
rect 160 31734 169 31768
rect 117 31696 169 31734
rect 117 31662 126 31696
rect 160 31662 169 31696
rect 117 31624 169 31662
rect 117 31590 126 31624
rect 160 31590 169 31624
rect 117 31552 169 31590
rect 117 31518 126 31552
rect 160 31518 169 31552
rect 117 31480 169 31518
rect 117 31446 126 31480
rect 160 31446 169 31480
rect 117 31408 169 31446
rect 117 31374 126 31408
rect 160 31374 169 31408
rect 117 31336 169 31374
rect 117 31302 126 31336
rect 160 31302 169 31336
rect 117 31264 169 31302
rect 117 31230 126 31264
rect 160 31230 169 31264
rect 117 31192 169 31230
rect 117 31158 126 31192
rect 160 31158 169 31192
rect 117 31120 169 31158
rect 117 31086 126 31120
rect 160 31086 169 31120
rect 117 31048 169 31086
rect 117 31014 126 31048
rect 160 31014 169 31048
rect 117 30976 169 31014
rect 117 30942 126 30976
rect 160 30942 169 30976
rect 117 30904 169 30942
rect 117 30870 126 30904
rect 160 30870 169 30904
rect 117 30832 169 30870
rect 117 30798 126 30832
rect 160 30798 169 30832
rect 117 30760 169 30798
rect 117 30726 126 30760
rect 160 30726 169 30760
rect 117 30688 169 30726
rect 117 30654 126 30688
rect 160 30654 169 30688
rect 117 30616 169 30654
rect 117 30582 126 30616
rect 160 30582 169 30616
rect 117 30544 169 30582
rect 117 30510 126 30544
rect 160 30510 169 30544
rect 117 30472 169 30510
rect 117 30438 126 30472
rect 160 30438 169 30472
rect 117 30400 169 30438
rect 117 30366 126 30400
rect 160 30366 169 30400
rect 117 30328 169 30366
rect 117 30294 126 30328
rect 160 30294 169 30328
rect 117 30256 169 30294
rect 117 30222 126 30256
rect 160 30222 169 30256
rect 117 30184 169 30222
rect 117 30150 126 30184
rect 160 30150 169 30184
rect 117 30112 169 30150
rect 117 30078 126 30112
rect 160 30078 169 30112
rect 117 30040 169 30078
rect 117 30006 126 30040
rect 160 30006 169 30040
rect 117 29968 169 30006
rect 117 29934 126 29968
rect 160 29934 169 29968
rect 117 29896 169 29934
rect 117 29862 126 29896
rect 160 29862 169 29896
rect 117 29824 169 29862
rect 117 29790 126 29824
rect 160 29790 169 29824
rect 117 29752 169 29790
rect 117 29718 126 29752
rect 160 29718 169 29752
rect 117 29680 169 29718
rect 117 29646 126 29680
rect 160 29646 169 29680
rect 117 29608 169 29646
rect 117 29574 126 29608
rect 160 29574 169 29608
rect 117 29536 169 29574
rect 117 29502 126 29536
rect 160 29502 169 29536
rect 117 29464 169 29502
rect 117 29430 126 29464
rect 160 29430 169 29464
rect 117 29392 169 29430
rect 117 29358 126 29392
rect 160 29358 169 29392
rect 117 29320 169 29358
rect 117 29286 126 29320
rect 160 29286 169 29320
rect 117 29248 169 29286
rect 117 29214 126 29248
rect 160 29214 169 29248
rect 117 29176 169 29214
rect 117 29142 126 29176
rect 160 29142 169 29176
rect 117 29104 169 29142
rect 117 29070 126 29104
rect 160 29070 169 29104
rect 117 29032 169 29070
rect 117 28998 126 29032
rect 160 28998 169 29032
rect 117 28960 169 28998
rect 117 28926 126 28960
rect 160 28926 169 28960
rect 117 28888 169 28926
rect 117 28854 126 28888
rect 160 28854 169 28888
rect 117 28816 169 28854
rect 117 28782 126 28816
rect 160 28782 169 28816
rect 117 28744 169 28782
rect 117 28710 126 28744
rect 160 28710 169 28744
rect 117 28672 169 28710
rect 117 28638 126 28672
rect 160 28638 169 28672
rect 117 28600 169 28638
rect 117 28566 126 28600
rect 160 28566 169 28600
rect 117 28528 169 28566
rect 117 28494 126 28528
rect 160 28494 169 28528
rect 117 28456 169 28494
rect 117 28422 126 28456
rect 160 28422 169 28456
rect 117 28384 169 28422
rect 117 28350 126 28384
rect 160 28350 169 28384
rect 117 28312 169 28350
rect 117 28278 126 28312
rect 160 28278 169 28312
rect 117 28240 169 28278
rect 117 28206 126 28240
rect 160 28206 169 28240
rect 117 28168 169 28206
rect 117 28134 126 28168
rect 160 28134 169 28168
rect 117 28096 169 28134
rect 117 28062 126 28096
rect 160 28062 169 28096
rect 117 28024 169 28062
rect 117 27990 126 28024
rect 160 27990 169 28024
rect 117 27952 169 27990
rect 117 27918 126 27952
rect 160 27918 169 27952
rect 117 27880 169 27918
rect 117 27846 126 27880
rect 160 27846 169 27880
rect 117 27808 169 27846
rect 117 27774 126 27808
rect 160 27774 169 27808
rect 117 27736 169 27774
rect 117 27702 126 27736
rect 160 27702 169 27736
rect 117 27664 169 27702
rect 117 27630 126 27664
rect 160 27630 169 27664
rect 117 27592 169 27630
rect 117 27558 126 27592
rect 160 27558 169 27592
rect 117 27520 169 27558
rect 117 27486 126 27520
rect 160 27486 169 27520
rect 117 27448 169 27486
rect 117 27414 126 27448
rect 160 27414 169 27448
rect 117 27376 169 27414
rect 117 27342 126 27376
rect 160 27342 169 27376
rect 117 27304 169 27342
rect 117 27270 126 27304
rect 160 27270 169 27304
rect 117 27232 169 27270
rect 117 27198 126 27232
rect 160 27198 169 27232
rect 117 27160 169 27198
rect 117 27126 126 27160
rect 160 27126 169 27160
rect 117 27088 169 27126
rect 117 27054 126 27088
rect 160 27054 169 27088
rect 117 27016 169 27054
rect 117 26982 126 27016
rect 160 26982 169 27016
rect 117 26944 169 26982
rect 117 26910 126 26944
rect 160 26910 169 26944
rect 117 26872 169 26910
rect 117 26838 126 26872
rect 160 26838 169 26872
rect 117 26800 169 26838
rect 117 26766 126 26800
rect 160 26766 169 26800
rect 117 26728 169 26766
rect 117 26694 126 26728
rect 160 26694 169 26728
rect 117 26656 169 26694
rect 117 26622 126 26656
rect 160 26622 169 26656
rect 117 26584 169 26622
rect 117 26550 126 26584
rect 160 26550 169 26584
rect 117 26512 169 26550
rect 117 26478 126 26512
rect 160 26478 169 26512
rect 117 26440 169 26478
rect 117 26406 126 26440
rect 160 26406 169 26440
rect 117 26368 169 26406
rect 117 26334 126 26368
rect 160 26334 169 26368
rect 117 26296 169 26334
rect 117 26262 126 26296
rect 160 26262 169 26296
rect 117 26224 169 26262
rect 117 26190 126 26224
rect 160 26190 169 26224
rect 117 26152 169 26190
rect 117 26118 126 26152
rect 160 26118 169 26152
rect 117 26080 169 26118
rect 117 26046 126 26080
rect 160 26046 169 26080
rect 117 26008 169 26046
rect 117 25974 126 26008
rect 160 25974 169 26008
rect 117 25936 169 25974
rect 117 25902 126 25936
rect 160 25902 169 25936
rect 117 25864 169 25902
rect 117 25830 126 25864
rect 160 25830 169 25864
rect 117 25792 169 25830
rect 117 25758 126 25792
rect 160 25758 169 25792
rect 117 25720 169 25758
rect 117 25686 126 25720
rect 160 25686 169 25720
rect 117 25648 169 25686
rect 117 25614 126 25648
rect 160 25614 169 25648
rect 117 25576 169 25614
rect 117 25542 126 25576
rect 160 25542 169 25576
rect 117 25504 169 25542
rect 117 25470 126 25504
rect 160 25470 169 25504
rect 117 25432 169 25470
rect 117 25398 126 25432
rect 160 25398 169 25432
rect 117 25360 169 25398
rect 117 25326 126 25360
rect 160 25326 169 25360
rect 117 25288 169 25326
rect 117 25254 126 25288
rect 160 25254 169 25288
rect 117 25216 169 25254
rect 117 25182 126 25216
rect 160 25182 169 25216
rect 117 25144 169 25182
rect 117 25110 126 25144
rect 160 25110 169 25144
rect 117 25072 169 25110
rect 117 25038 126 25072
rect 160 25038 169 25072
rect 117 25000 169 25038
rect 117 24966 126 25000
rect 160 24966 169 25000
rect 117 24928 169 24966
rect 117 24894 126 24928
rect 160 24894 169 24928
rect 117 24856 169 24894
rect 117 24822 126 24856
rect 160 24822 169 24856
rect 117 24784 169 24822
rect 117 24750 126 24784
rect 160 24750 169 24784
rect 117 24712 169 24750
rect 117 24678 126 24712
rect 160 24678 169 24712
rect 117 24640 169 24678
rect 117 24606 126 24640
rect 160 24606 169 24640
rect 117 24568 169 24606
rect 117 24534 126 24568
rect 160 24534 169 24568
rect 117 24496 169 24534
rect 117 24462 126 24496
rect 160 24462 169 24496
rect 117 24424 169 24462
rect 117 24390 126 24424
rect 160 24390 169 24424
rect 117 24352 169 24390
rect 117 24318 126 24352
rect 160 24318 169 24352
rect 117 24280 169 24318
rect 117 24246 126 24280
rect 160 24246 169 24280
rect 117 24208 169 24246
rect 117 24174 126 24208
rect 160 24174 169 24208
rect 117 24136 169 24174
rect 117 24102 126 24136
rect 160 24102 169 24136
rect 117 24064 169 24102
rect 117 24030 126 24064
rect 160 24030 169 24064
rect 117 23992 169 24030
rect 117 23958 126 23992
rect 160 23958 169 23992
rect 117 23920 169 23958
rect 117 23886 126 23920
rect 160 23886 169 23920
rect 117 23848 169 23886
rect 117 23814 126 23848
rect 160 23814 169 23848
rect 117 23776 169 23814
rect 117 23742 126 23776
rect 160 23742 169 23776
rect 117 23704 169 23742
rect 117 23670 126 23704
rect 160 23670 169 23704
rect 117 23632 169 23670
rect 117 23598 126 23632
rect 160 23598 169 23632
rect 117 23560 169 23598
rect 117 23526 126 23560
rect 160 23526 169 23560
rect 117 23488 169 23526
rect 117 23454 126 23488
rect 160 23454 169 23488
rect 117 23416 169 23454
rect 117 23382 126 23416
rect 160 23382 169 23416
rect 117 23344 169 23382
rect 117 23310 126 23344
rect 160 23310 169 23344
rect 117 23272 169 23310
rect 117 23238 126 23272
rect 160 23238 169 23272
rect 117 23200 169 23238
rect 117 23166 126 23200
rect 160 23166 169 23200
rect 117 23128 169 23166
rect 117 23094 126 23128
rect 160 23094 169 23128
rect 117 23056 169 23094
rect 117 23022 126 23056
rect 160 23022 169 23056
rect 117 22984 169 23022
rect 117 22950 126 22984
rect 160 22950 169 22984
rect 117 22912 169 22950
rect 117 22878 126 22912
rect 160 22878 169 22912
rect 117 22840 169 22878
rect 117 22806 126 22840
rect 160 22806 169 22840
rect 117 22768 169 22806
rect 117 22734 126 22768
rect 160 22734 169 22768
rect 117 22696 169 22734
rect 117 22662 126 22696
rect 160 22662 169 22696
rect 117 22624 169 22662
rect 117 22590 126 22624
rect 160 22590 169 22624
rect 117 22552 169 22590
rect 117 22518 126 22552
rect 160 22518 169 22552
rect 117 22480 169 22518
rect 117 22446 126 22480
rect 160 22446 169 22480
rect 117 22408 169 22446
rect 117 22374 126 22408
rect 160 22374 169 22408
rect 117 22336 169 22374
rect 117 22302 126 22336
rect 160 22302 169 22336
rect 117 22264 169 22302
rect 117 22230 126 22264
rect 160 22230 169 22264
rect 117 22192 169 22230
rect 117 22158 126 22192
rect 160 22158 169 22192
rect 117 22120 169 22158
rect 117 22086 126 22120
rect 160 22086 169 22120
rect 117 22048 169 22086
rect 117 22014 126 22048
rect 160 22014 169 22048
rect 117 21976 169 22014
rect 117 21942 126 21976
rect 160 21942 169 21976
rect 117 21904 169 21942
rect 117 21870 126 21904
rect 160 21870 169 21904
rect 117 21832 169 21870
rect 117 21798 126 21832
rect 160 21798 169 21832
rect 117 21760 169 21798
rect 117 21726 126 21760
rect 160 21726 169 21760
rect 117 21688 169 21726
rect 117 21654 126 21688
rect 160 21654 169 21688
rect 117 21616 169 21654
rect 117 21582 126 21616
rect 160 21582 169 21616
rect 117 21544 169 21582
rect 117 21510 126 21544
rect 160 21510 169 21544
rect 117 21472 169 21510
rect 117 21438 126 21472
rect 160 21438 169 21472
rect 117 21400 169 21438
rect 117 21366 126 21400
rect 160 21366 169 21400
rect 117 21328 169 21366
rect 117 21294 126 21328
rect 160 21294 169 21328
rect 117 21256 169 21294
rect 117 21222 126 21256
rect 160 21222 169 21256
rect 117 21184 169 21222
rect 117 21150 126 21184
rect 160 21150 169 21184
rect 117 21112 169 21150
rect 117 21078 126 21112
rect 160 21078 169 21112
rect 117 21040 169 21078
rect 117 21006 126 21040
rect 160 21006 169 21040
rect 117 20968 169 21006
rect 117 20934 126 20968
rect 160 20934 169 20968
rect 117 20896 169 20934
rect 117 20862 126 20896
rect 160 20862 169 20896
rect 117 20824 169 20862
rect 117 20790 126 20824
rect 160 20790 169 20824
rect 117 20752 169 20790
rect 117 20718 126 20752
rect 160 20718 169 20752
rect 117 20680 169 20718
rect 117 20646 126 20680
rect 160 20646 169 20680
rect 117 20608 169 20646
rect 117 20574 126 20608
rect 160 20574 169 20608
rect 117 20536 169 20574
rect 117 20502 126 20536
rect 160 20502 169 20536
rect 117 20464 169 20502
rect 117 20430 126 20464
rect 160 20430 169 20464
rect 117 20392 169 20430
rect 117 20358 126 20392
rect 160 20358 169 20392
rect 117 20320 169 20358
rect 117 20286 126 20320
rect 160 20286 169 20320
rect 117 20248 169 20286
rect 117 20214 126 20248
rect 160 20214 169 20248
rect 117 20176 169 20214
rect 117 20142 126 20176
rect 160 20142 169 20176
rect 117 20104 169 20142
rect 117 20070 126 20104
rect 160 20070 169 20104
rect 117 20032 169 20070
rect 117 19998 126 20032
rect 160 19998 169 20032
rect 117 19960 169 19998
rect 117 19926 126 19960
rect 160 19926 169 19960
rect 117 19888 169 19926
rect 117 19854 126 19888
rect 160 19854 169 19888
rect 117 19816 169 19854
rect 117 19782 126 19816
rect 160 19782 169 19816
rect 117 19744 169 19782
rect 117 19710 126 19744
rect 160 19710 169 19744
rect 117 19672 169 19710
rect 117 19638 126 19672
rect 160 19638 169 19672
rect 117 19600 169 19638
rect 117 19566 126 19600
rect 160 19566 169 19600
rect 117 19528 169 19566
rect 117 19494 126 19528
rect 160 19494 169 19528
rect 117 19456 169 19494
rect 117 19422 126 19456
rect 160 19422 169 19456
rect 117 19384 169 19422
rect 117 19350 126 19384
rect 160 19350 169 19384
rect 117 19312 169 19350
rect 117 19278 126 19312
rect 160 19278 169 19312
rect 117 19240 169 19278
rect 117 19206 126 19240
rect 160 19206 169 19240
rect 117 19168 169 19206
rect 117 19134 126 19168
rect 160 19134 169 19168
rect 117 19096 169 19134
rect 117 19062 126 19096
rect 160 19062 169 19096
rect 117 19024 169 19062
rect 117 18990 126 19024
rect 160 18990 169 19024
rect 117 18952 169 18990
rect 117 18918 126 18952
rect 160 18918 169 18952
rect 117 18880 169 18918
rect 117 18846 126 18880
rect 160 18846 169 18880
rect 117 18808 169 18846
rect 117 18774 126 18808
rect 160 18774 169 18808
rect 117 18736 169 18774
rect 117 18702 126 18736
rect 160 18702 169 18736
rect 117 18664 169 18702
rect 117 18630 126 18664
rect 160 18630 169 18664
rect 117 18592 169 18630
rect 117 18558 126 18592
rect 160 18558 169 18592
rect 117 18520 169 18558
rect 117 18486 126 18520
rect 160 18486 169 18520
rect 117 18448 169 18486
rect 117 18414 126 18448
rect 160 18414 169 18448
rect 117 18376 169 18414
rect 117 18342 126 18376
rect 160 18342 169 18376
rect 117 18304 169 18342
rect 117 18270 126 18304
rect 160 18270 169 18304
rect 117 18232 169 18270
rect 117 18198 126 18232
rect 160 18198 169 18232
rect 117 18160 169 18198
rect 117 18126 126 18160
rect 160 18126 169 18160
rect 117 18088 169 18126
rect 117 18054 126 18088
rect 160 18054 169 18088
rect 117 18016 169 18054
rect 117 17982 126 18016
rect 160 17982 169 18016
rect 117 17944 169 17982
rect 117 17910 126 17944
rect 160 17910 169 17944
rect 117 17872 169 17910
rect 117 17838 126 17872
rect 160 17838 169 17872
rect 117 17800 169 17838
rect 117 17766 126 17800
rect 160 17766 169 17800
rect 117 17728 169 17766
rect 117 17694 126 17728
rect 160 17694 169 17728
rect 117 17656 169 17694
rect 117 17622 126 17656
rect 160 17622 169 17656
rect 117 17584 169 17622
rect 117 17550 126 17584
rect 160 17550 169 17584
rect 117 17512 169 17550
rect 117 17478 126 17512
rect 160 17478 169 17512
rect 117 17440 169 17478
rect 117 17406 126 17440
rect 160 17406 169 17440
rect 117 17368 169 17406
rect 117 17334 126 17368
rect 160 17334 169 17368
rect 117 17296 169 17334
rect 117 17262 126 17296
rect 160 17262 169 17296
rect 117 17224 169 17262
rect 117 17190 126 17224
rect 160 17190 169 17224
rect 117 17152 169 17190
rect 117 17118 126 17152
rect 160 17118 169 17152
rect 117 17080 169 17118
rect 117 17046 126 17080
rect 160 17046 169 17080
rect 117 17008 169 17046
rect 117 16974 126 17008
rect 160 16974 169 17008
rect 117 16936 169 16974
rect 117 16902 126 16936
rect 160 16902 169 16936
rect 117 16864 169 16902
rect 117 16830 126 16864
rect 160 16830 169 16864
rect 117 16792 169 16830
rect 117 16758 126 16792
rect 160 16758 169 16792
rect 117 16720 169 16758
rect 117 16686 126 16720
rect 160 16686 169 16720
rect 117 16648 169 16686
rect 117 16614 126 16648
rect 160 16614 169 16648
rect 117 16576 169 16614
rect 117 16542 126 16576
rect 160 16542 169 16576
rect 117 16504 169 16542
rect 117 16470 126 16504
rect 160 16470 169 16504
rect 117 16432 169 16470
rect 117 16398 126 16432
rect 160 16398 169 16432
rect 117 16360 169 16398
rect 117 16326 126 16360
rect 160 16326 169 16360
rect 117 16288 169 16326
rect 117 16254 126 16288
rect 160 16254 169 16288
rect 117 16216 169 16254
rect 117 16182 126 16216
rect 160 16182 169 16216
rect 117 16144 169 16182
rect 117 16110 126 16144
rect 160 16110 169 16144
rect 117 16072 169 16110
rect 117 16038 126 16072
rect 160 16038 169 16072
rect 117 16000 169 16038
rect 117 15966 126 16000
rect 160 15966 169 16000
rect 117 15928 169 15966
rect 117 15894 126 15928
rect 160 15894 169 15928
rect 117 15856 169 15894
rect 117 15822 126 15856
rect 160 15822 169 15856
rect 117 15784 169 15822
rect 117 15750 126 15784
rect 160 15750 169 15784
rect 117 15712 169 15750
rect 117 15678 126 15712
rect 160 15678 169 15712
rect 117 15640 169 15678
rect 117 15606 126 15640
rect 160 15606 169 15640
rect 117 15568 169 15606
rect 117 15534 126 15568
rect 160 15534 169 15568
rect 117 15496 169 15534
rect 117 15462 126 15496
rect 160 15462 169 15496
rect 117 15424 169 15462
rect 117 15390 126 15424
rect 160 15390 169 15424
rect 117 15352 169 15390
rect 117 15318 126 15352
rect 160 15318 169 15352
rect 117 15280 169 15318
rect 117 15246 126 15280
rect 160 15246 169 15280
rect 117 15208 169 15246
rect 117 15174 126 15208
rect 160 15174 169 15208
rect 117 15136 169 15174
rect 117 15102 126 15136
rect 160 15102 169 15136
rect 117 15064 169 15102
rect 117 15030 126 15064
rect 160 15030 169 15064
rect 117 14992 169 15030
rect 117 14958 126 14992
rect 160 14958 169 14992
rect 117 14920 169 14958
rect 117 14886 126 14920
rect 160 14886 169 14920
rect 117 14848 169 14886
rect 117 14814 126 14848
rect 160 14814 169 14848
rect 117 14776 169 14814
rect 117 14742 126 14776
rect 160 14742 169 14776
rect 117 14704 169 14742
rect 117 14670 126 14704
rect 160 14670 169 14704
rect 117 14632 169 14670
rect 117 14598 126 14632
rect 160 14598 169 14632
rect 117 14560 169 14598
rect 117 14526 126 14560
rect 160 14526 169 14560
rect 117 14488 169 14526
rect 117 14454 126 14488
rect 160 14454 169 14488
rect 117 14416 169 14454
rect 117 14382 126 14416
rect 160 14382 169 14416
rect 117 14344 169 14382
rect 117 14310 126 14344
rect 160 14310 169 14344
rect 117 14272 169 14310
rect 117 14238 126 14272
rect 160 14238 169 14272
rect 117 14200 169 14238
rect 117 14166 126 14200
rect 160 14166 169 14200
rect 117 14128 169 14166
rect 117 14094 126 14128
rect 160 14094 169 14128
rect 117 14056 169 14094
rect 117 14022 126 14056
rect 160 14022 169 14056
rect 117 13984 169 14022
rect 117 13950 126 13984
rect 160 13950 169 13984
rect 117 13912 169 13950
rect 117 13878 126 13912
rect 160 13878 169 13912
rect 117 13840 169 13878
rect 117 13806 126 13840
rect 160 13806 169 13840
rect 117 13768 169 13806
rect 117 13734 126 13768
rect 160 13734 169 13768
rect 117 13701 169 13734
rect 117 13633 169 13649
rect 117 13565 169 13581
rect 117 13496 169 13513
rect 117 13427 169 13444
rect 117 13374 126 13375
rect 160 13374 169 13375
rect 117 13358 169 13374
rect 117 13302 126 13306
rect 160 13302 169 13306
rect 117 13289 169 13302
rect 117 13230 126 13237
rect 160 13230 169 13237
rect 117 13220 169 13230
rect 117 13158 126 13168
rect 160 13158 169 13168
rect 117 13151 169 13158
rect 117 13086 126 13099
rect 160 13086 169 13099
rect 117 13082 169 13086
rect 117 13014 126 13030
rect 160 13014 169 13030
rect 117 13013 169 13014
rect 117 12944 126 12961
rect 160 12944 169 12961
rect 117 12875 126 12892
rect 160 12875 169 12892
rect 117 12798 126 12823
rect 160 12798 169 12823
rect 117 12760 169 12798
rect 117 12726 126 12760
rect 160 12726 169 12760
rect 117 12688 169 12726
rect 117 12654 126 12688
rect 160 12654 169 12688
rect 117 12616 169 12654
rect 117 12582 126 12616
rect 160 12582 169 12616
rect 117 12544 169 12582
rect 117 12510 126 12544
rect 160 12510 169 12544
rect 117 12472 169 12510
rect 117 12438 126 12472
rect 160 12438 169 12472
rect 117 12400 169 12438
rect 117 12366 126 12400
rect 160 12366 169 12400
rect 117 12328 169 12366
rect 117 12294 126 12328
rect 160 12294 169 12328
rect 117 12256 169 12294
rect 117 12222 126 12256
rect 160 12222 169 12256
rect 117 12184 169 12222
rect 117 12150 126 12184
rect 160 12150 169 12184
rect 117 12112 169 12150
rect 117 12078 126 12112
rect 160 12078 169 12112
rect 117 12040 169 12078
rect 117 12006 126 12040
rect 160 12006 169 12040
rect 117 11968 169 12006
rect 117 11934 126 11968
rect 160 11934 169 11968
rect 117 11896 169 11934
rect 117 11862 126 11896
rect 160 11862 169 11896
rect 117 11824 169 11862
rect 117 11790 126 11824
rect 160 11790 169 11824
rect 117 11752 169 11790
rect 117 11718 126 11752
rect 160 11718 169 11752
rect 117 11680 169 11718
rect 117 11646 126 11680
rect 160 11646 169 11680
rect 117 11608 169 11646
rect 117 11574 126 11608
rect 160 11574 169 11608
rect 117 11536 169 11574
rect 117 11502 126 11536
rect 160 11502 169 11536
rect 117 11464 169 11502
rect 117 11430 126 11464
rect 160 11430 169 11464
rect 117 11392 169 11430
rect 117 11358 126 11392
rect 160 11358 169 11392
rect 117 11320 169 11358
rect 117 11286 126 11320
rect 160 11286 169 11320
rect 117 11248 169 11286
rect 117 11214 126 11248
rect 160 11214 169 11248
rect 117 11176 169 11214
rect 117 11142 126 11176
rect 160 11142 169 11176
rect 117 11104 169 11142
rect 117 11070 126 11104
rect 160 11070 169 11104
rect 117 11032 169 11070
rect 117 10998 126 11032
rect 160 10998 169 11032
rect 117 10960 169 10998
rect 117 10926 126 10960
rect 160 10926 169 10960
rect 117 10888 169 10926
rect 117 10854 126 10888
rect 160 10854 169 10888
rect 117 10816 169 10854
rect 117 10782 126 10816
rect 160 10782 169 10816
rect 117 10744 169 10782
rect 117 10710 126 10744
rect 160 10710 169 10744
rect 117 10672 169 10710
rect 117 10638 126 10672
rect 160 10638 169 10672
rect 117 10600 169 10638
rect 117 10566 126 10600
rect 160 10566 169 10600
rect 117 10528 169 10566
rect 117 10494 126 10528
rect 160 10494 169 10528
rect 117 10456 169 10494
rect 117 10422 126 10456
rect 160 10422 169 10456
rect 117 10384 169 10422
rect 117 10350 126 10384
rect 160 10350 169 10384
rect 117 10312 169 10350
rect 117 10278 126 10312
rect 160 10278 169 10312
rect 117 10240 169 10278
rect 117 10206 126 10240
rect 160 10206 169 10240
rect 117 10168 169 10206
rect 117 10134 126 10168
rect 160 10134 169 10168
rect 117 10096 169 10134
rect 117 10062 126 10096
rect 160 10062 169 10096
rect 117 10024 169 10062
rect 117 9990 126 10024
rect 160 9990 169 10024
rect 117 9952 169 9990
rect 117 9918 126 9952
rect 160 9918 169 9952
rect 117 9880 169 9918
rect 117 9846 126 9880
rect 160 9846 169 9880
rect 117 9808 169 9846
rect 117 9774 126 9808
rect 160 9774 169 9808
rect 117 9736 169 9774
rect 117 9702 126 9736
rect 160 9702 169 9736
rect 117 9664 169 9702
rect 117 9630 126 9664
rect 160 9630 169 9664
rect 117 9592 169 9630
rect 117 9558 126 9592
rect 160 9558 169 9592
rect 117 9520 169 9558
rect 117 9486 126 9520
rect 160 9486 169 9520
rect 117 9448 169 9486
rect 117 9414 126 9448
rect 160 9414 169 9448
rect 117 9376 169 9414
rect 117 9342 126 9376
rect 160 9342 169 9376
rect 117 9304 169 9342
rect 117 9270 126 9304
rect 160 9270 169 9304
rect 117 9232 169 9270
rect 117 9198 126 9232
rect 160 9198 169 9232
rect 117 9160 169 9198
rect 117 9126 126 9160
rect 160 9126 169 9160
rect 117 9088 169 9126
rect 117 9054 126 9088
rect 160 9054 169 9088
rect 117 9016 169 9054
rect 117 8982 126 9016
rect 160 8982 169 9016
rect 117 8944 169 8982
rect 117 8910 126 8944
rect 160 8910 169 8944
rect 117 8872 169 8910
rect 117 8838 126 8872
rect 160 8838 169 8872
rect 117 8800 169 8838
rect 117 8766 126 8800
rect 160 8766 169 8800
rect 117 8728 169 8766
rect 117 8694 126 8728
rect 160 8694 169 8728
rect 117 8656 169 8694
rect 117 8622 126 8656
rect 160 8622 169 8656
rect 117 8584 169 8622
rect 117 8550 126 8584
rect 160 8550 169 8584
rect 117 8512 169 8550
rect 117 8478 126 8512
rect 160 8478 169 8512
rect 117 8440 169 8478
rect 117 8406 126 8440
rect 160 8406 169 8440
rect 117 8368 169 8406
rect 117 8334 126 8368
rect 160 8334 169 8368
rect 117 8296 169 8334
rect 117 8262 126 8296
rect 160 8262 169 8296
rect 117 8224 169 8262
rect 117 8190 126 8224
rect 160 8190 169 8224
rect 117 8152 169 8190
rect 117 8118 126 8152
rect 160 8118 169 8152
rect 117 8080 169 8118
rect 117 8046 126 8080
rect 160 8046 169 8080
rect 117 8008 169 8046
rect 117 7974 126 8008
rect 160 7974 169 8008
rect 117 7936 169 7974
rect 117 7902 126 7936
rect 160 7902 169 7936
rect 117 7864 169 7902
rect 117 7830 126 7864
rect 160 7830 169 7864
rect 117 7792 169 7830
rect 117 7758 126 7792
rect 160 7758 169 7792
rect 117 7720 169 7758
rect 117 7686 126 7720
rect 160 7686 169 7720
rect 117 7648 169 7686
rect 117 7614 126 7648
rect 160 7614 169 7648
rect 117 7576 169 7614
rect 117 7542 126 7576
rect 160 7542 169 7576
rect 117 7504 169 7542
rect 117 7470 126 7504
rect 160 7470 169 7504
rect 117 7432 169 7470
rect 117 7398 126 7432
rect 160 7398 169 7432
rect 117 7360 169 7398
rect 117 7326 126 7360
rect 160 7326 169 7360
rect 117 7288 169 7326
rect 117 7254 126 7288
rect 160 7254 169 7288
rect 117 7216 169 7254
rect 117 7182 126 7216
rect 160 7182 169 7216
rect 117 7144 169 7182
rect 117 7110 126 7144
rect 160 7110 169 7144
rect 117 7072 169 7110
rect 117 7038 126 7072
rect 160 7038 169 7072
rect 117 7000 169 7038
rect 117 6966 126 7000
rect 160 6966 169 7000
rect 117 6928 169 6966
rect 117 6894 126 6928
rect 160 6894 169 6928
rect 117 6856 169 6894
rect 117 6822 126 6856
rect 160 6822 169 6856
rect 117 6784 169 6822
rect 117 6750 126 6784
rect 160 6750 169 6784
rect 117 6712 169 6750
rect 117 6678 126 6712
rect 160 6678 169 6712
rect 117 6640 169 6678
rect 117 6606 126 6640
rect 160 6606 169 6640
rect 117 6568 169 6606
rect 117 6534 126 6568
rect 160 6534 169 6568
rect 117 6496 169 6534
rect 117 6462 126 6496
rect 160 6462 169 6496
rect 117 6424 169 6462
rect 117 6390 126 6424
rect 160 6390 169 6424
rect 117 6352 169 6390
rect 117 6318 126 6352
rect 160 6318 169 6352
rect 117 6280 169 6318
rect 117 6246 126 6280
rect 160 6246 169 6280
rect 117 6208 169 6246
rect 117 6174 126 6208
rect 160 6174 169 6208
rect 117 6136 169 6174
rect 117 6102 126 6136
rect 160 6102 169 6136
rect 117 6064 169 6102
rect 117 6030 126 6064
rect 160 6030 169 6064
rect 117 5992 169 6030
rect 117 5958 126 5992
rect 160 5958 169 5992
rect 117 5920 169 5958
rect 117 5886 126 5920
rect 160 5886 169 5920
rect 117 5848 169 5886
rect 117 5814 126 5848
rect 160 5814 169 5848
rect 117 5776 169 5814
rect 117 5742 126 5776
rect 160 5742 169 5776
rect 117 5704 169 5742
rect 117 5670 126 5704
rect 160 5670 169 5704
rect 117 5632 169 5670
rect 117 5598 126 5632
rect 160 5598 169 5632
rect 117 5560 169 5598
rect 117 5526 126 5560
rect 160 5526 169 5560
rect 117 5488 169 5526
rect 117 5454 126 5488
rect 160 5454 169 5488
rect 117 5416 169 5454
rect 117 5382 126 5416
rect 160 5382 169 5416
rect 117 5344 169 5382
rect 117 5310 126 5344
rect 160 5310 169 5344
rect 117 5272 169 5310
rect 117 5238 126 5272
rect 160 5238 169 5272
rect 117 5200 169 5238
rect 117 5166 126 5200
rect 160 5166 169 5200
rect 117 5128 169 5166
rect 117 5094 126 5128
rect 160 5094 169 5128
rect 117 5056 169 5094
rect 117 5022 126 5056
rect 160 5022 169 5056
rect 117 4984 169 5022
rect 117 4950 126 4984
rect 160 4950 169 4984
rect 117 4912 169 4950
rect 117 4878 126 4912
rect 160 4878 169 4912
rect 117 4840 169 4878
rect 117 4806 126 4840
rect 160 4806 169 4840
rect 117 4768 169 4806
rect 117 4734 126 4768
rect 160 4734 169 4768
rect 117 4696 169 4734
rect 117 4662 126 4696
rect 160 4662 169 4696
rect 117 4624 169 4662
rect 117 4590 126 4624
rect 160 4590 169 4624
rect 117 4552 169 4590
rect 117 4518 126 4552
rect 160 4518 169 4552
rect 117 4480 169 4518
rect 117 4446 126 4480
rect 160 4446 169 4480
rect 117 4408 169 4446
rect 117 4374 126 4408
rect 160 4374 169 4408
rect 117 4336 169 4374
rect 117 4302 126 4336
rect 160 4302 169 4336
rect 117 4264 169 4302
rect 117 4230 126 4264
rect 160 4230 169 4264
rect 117 4192 169 4230
rect 117 4158 126 4192
rect 160 4158 169 4192
rect 117 4120 169 4158
rect 117 4086 126 4120
rect 160 4086 169 4120
rect 117 4048 169 4086
rect 117 4014 126 4048
rect 160 4014 169 4048
rect 117 3976 169 4014
rect 117 3942 126 3976
rect 160 3942 169 3976
rect 117 3904 169 3942
rect 117 3870 126 3904
rect 160 3870 169 3904
rect 117 3832 169 3870
rect 117 3798 126 3832
rect 160 3798 169 3832
rect 117 3760 169 3798
rect 117 3726 126 3760
rect 160 3726 169 3760
rect 117 3688 169 3726
rect 117 3654 126 3688
rect 160 3654 169 3688
rect 117 3616 169 3654
rect 117 3582 126 3616
rect 160 3582 169 3616
rect 117 3544 169 3582
rect 117 3510 126 3544
rect 160 3510 169 3544
rect 117 3472 169 3510
rect 117 3438 126 3472
rect 160 3438 169 3472
rect 117 3400 169 3438
rect 117 3366 126 3400
rect 160 3366 169 3400
rect 117 3328 169 3366
rect 117 3294 126 3328
rect 160 3294 169 3328
rect 117 3256 169 3294
rect 117 3222 126 3256
rect 160 3222 169 3256
rect 117 3184 169 3222
rect 117 3150 126 3184
rect 160 3150 169 3184
rect 117 3112 169 3150
rect 117 3078 126 3112
rect 160 3078 169 3112
rect 117 3040 169 3078
rect 117 3006 126 3040
rect 160 3006 169 3040
rect 117 2968 169 3006
rect 117 2934 126 2968
rect 160 2934 169 2968
rect 117 2896 169 2934
rect 117 2862 126 2896
rect 160 2862 169 2896
rect 117 2824 169 2862
rect 117 2790 126 2824
rect 160 2790 169 2824
rect 117 2752 169 2790
rect 117 2718 126 2752
rect 160 2718 169 2752
rect 117 2680 169 2718
rect 117 2646 126 2680
rect 160 2646 169 2680
rect 117 2608 169 2646
rect 117 2574 126 2608
rect 160 2574 169 2608
rect 117 2536 169 2574
rect 117 2502 126 2536
rect 160 2502 169 2536
rect 117 2464 169 2502
rect 117 2430 126 2464
rect 160 2430 169 2464
rect 117 2392 169 2430
rect 117 2358 126 2392
rect 160 2358 169 2392
rect 117 2320 169 2358
rect 117 2286 126 2320
rect 160 2286 169 2320
rect 117 2248 169 2286
rect 117 2214 126 2248
rect 160 2214 169 2248
rect 117 2176 169 2214
rect 117 2142 126 2176
rect 160 2142 169 2176
rect 117 2104 169 2142
rect 117 2070 126 2104
rect 160 2070 169 2104
rect 117 2032 169 2070
rect 117 1998 126 2032
rect 160 1998 169 2032
rect 117 1960 169 1998
rect 117 1926 126 1960
rect 160 1926 169 1960
rect 117 1888 169 1926
rect 117 1854 126 1888
rect 160 1854 169 1888
rect 117 1816 169 1854
rect 117 1782 126 1816
rect 160 1782 169 1816
rect 117 1744 169 1782
rect 117 1710 126 1744
rect 160 1710 169 1744
rect 117 1672 169 1710
rect 117 1638 126 1672
rect 160 1638 169 1672
rect 117 1600 169 1638
rect 117 1566 126 1600
rect 160 1566 169 1600
rect 117 1528 169 1566
rect 117 1494 126 1528
rect 160 1494 169 1528
rect 117 1456 169 1494
rect 117 1422 126 1456
rect 160 1422 169 1456
rect 117 1384 169 1422
rect 117 1350 126 1384
rect 160 1350 169 1384
rect 117 1312 169 1350
rect 117 1278 126 1312
rect 160 1278 169 1312
rect 117 1240 169 1278
rect 117 1206 126 1240
rect 160 1206 169 1240
rect 117 1168 169 1206
rect 117 1134 126 1168
rect 160 1134 169 1168
rect 117 1096 169 1134
rect 117 1062 126 1096
rect 160 1062 169 1096
rect 117 1024 169 1062
rect 117 990 126 1024
rect 160 990 169 1024
rect 117 952 169 990
rect 117 918 126 952
rect 160 918 169 952
rect 117 880 169 918
rect 117 846 126 880
rect 160 846 169 880
rect 117 808 169 846
rect 117 774 126 808
rect 160 774 169 808
rect 117 736 169 774
rect 117 702 126 736
rect 160 702 169 736
rect 117 664 169 702
rect 117 630 126 664
rect 160 630 169 664
rect 117 592 169 630
rect 117 558 126 592
rect 160 558 169 592
rect 117 520 169 558
rect 380 39178 3076 39184
rect 380 39144 462 39178
rect 496 39144 538 39178
rect 572 39144 648 39178
rect 682 39144 720 39178
rect 754 39144 792 39178
rect 826 39144 864 39178
rect 898 39144 936 39178
rect 970 39144 1008 39178
rect 1042 39144 1080 39178
rect 1114 39144 1152 39178
rect 1186 39144 1224 39178
rect 1258 39144 1296 39178
rect 1330 39144 1368 39178
rect 1402 39144 1440 39178
rect 1474 39144 1512 39178
rect 1546 39144 1584 39178
rect 1618 39144 1656 39178
rect 1690 39144 1728 39178
rect 1762 39144 1800 39178
rect 1834 39144 1872 39178
rect 1906 39144 1944 39178
rect 1978 39144 2016 39178
rect 2050 39144 2088 39178
rect 2122 39144 2161 39178
rect 2195 39144 2234 39178
rect 2268 39144 2307 39178
rect 2341 39144 2380 39178
rect 2414 39144 2453 39178
rect 2487 39144 2526 39178
rect 2560 39144 2599 39178
rect 2633 39144 2672 39178
rect 2706 39144 2745 39178
rect 2779 39144 2818 39178
rect 2852 39144 2891 39178
rect 2925 39144 2964 39178
rect 2998 39144 3076 39178
rect 380 39138 3076 39144
rect 380 39120 587 39138
tri 587 39120 605 39138 nw
tri 2851 39120 2869 39138 ne
rect 2869 39120 3076 39138
rect 380 39106 573 39120
tri 573 39106 587 39120 nw
tri 2869 39106 2883 39120 ne
rect 2883 39106 3076 39120
rect 380 39072 386 39106
rect 420 39072 571 39106
tri 571 39104 573 39106 nw
tri 2883 39104 2885 39106 ne
rect 380 39033 571 39072
rect 2885 39072 3036 39106
rect 3070 39072 3076 39106
rect 380 38999 386 39033
rect 420 38999 571 39033
rect 613 39011 1501 39063
rect 1553 39011 1569 39063
rect 1621 39011 1636 39063
rect 1688 39011 1703 39063
rect 1755 39011 1770 39063
rect 1822 39011 1837 39063
rect 1889 39011 2830 39063
rect 2885 39034 3076 39072
rect 380 38964 571 38999
rect 2885 39000 3036 39034
rect 3070 39000 3076 39034
rect 380 38960 531 38964
rect 380 38926 386 38960
rect 420 38930 531 38960
rect 565 38930 571 38964
rect 420 38926 571 38930
rect 380 38891 571 38926
rect 380 38887 531 38891
rect 380 38853 386 38887
rect 420 38857 531 38887
rect 565 38857 571 38891
rect 420 38853 571 38857
rect 380 38818 571 38853
rect 380 38814 531 38818
rect 380 38780 386 38814
rect 420 38784 531 38814
rect 565 38784 571 38818
rect 420 38780 571 38784
rect 380 38745 571 38780
rect 380 38741 531 38745
rect 380 38707 386 38741
rect 420 38711 531 38741
rect 565 38711 571 38745
rect 420 38707 571 38711
rect 380 38672 571 38707
rect 380 38668 531 38672
rect 380 38634 386 38668
rect 420 38638 531 38668
rect 565 38638 571 38672
rect 420 38634 571 38638
rect 380 38599 571 38634
rect 380 38595 531 38599
rect 380 38561 386 38595
rect 420 38565 531 38595
rect 565 38565 571 38599
rect 420 38561 571 38565
rect 380 38526 571 38561
rect 380 38522 531 38526
rect 380 38488 386 38522
rect 420 38492 531 38522
rect 565 38492 571 38526
rect 420 38488 571 38492
rect 761 38964 807 38976
rect 761 38930 767 38964
rect 801 38930 807 38964
rect 761 38891 807 38930
rect 761 38857 767 38891
rect 801 38857 807 38891
rect 761 38818 807 38857
rect 761 38784 767 38818
rect 801 38784 807 38818
rect 761 38745 807 38784
rect 761 38711 767 38745
rect 801 38711 807 38745
rect 761 38672 807 38711
rect 761 38638 767 38672
rect 801 38638 807 38672
rect 761 38599 807 38638
rect 761 38565 767 38599
rect 801 38565 807 38599
rect 761 38526 807 38565
rect 761 38492 767 38526
rect 801 38492 807 38526
rect 380 38472 571 38488
tri 571 38472 587 38488 sw
tri 745 38472 761 38488 se
rect 761 38472 807 38492
rect 997 38964 1043 38976
rect 997 38930 1003 38964
rect 1037 38930 1043 38964
rect 997 38891 1043 38930
rect 997 38857 1003 38891
rect 1037 38857 1043 38891
rect 997 38818 1043 38857
rect 997 38784 1003 38818
rect 1037 38784 1043 38818
rect 997 38745 1043 38784
rect 997 38711 1003 38745
rect 1037 38711 1043 38745
rect 997 38672 1043 38711
rect 997 38638 1003 38672
rect 1037 38638 1043 38672
rect 997 38599 1043 38638
rect 997 38565 1003 38599
rect 1037 38565 1043 38599
rect 997 38526 1043 38565
rect 997 38492 1003 38526
rect 1037 38492 1043 38526
tri 807 38472 823 38488 sw
tri 981 38472 997 38488 se
rect 997 38472 1043 38492
rect 1233 38964 1279 38976
rect 1233 38930 1239 38964
rect 1273 38930 1279 38964
rect 1233 38891 1279 38930
rect 1233 38857 1239 38891
rect 1273 38857 1279 38891
rect 1233 38818 1279 38857
rect 1233 38784 1239 38818
rect 1273 38784 1279 38818
rect 1233 38745 1279 38784
rect 1233 38711 1239 38745
rect 1273 38711 1279 38745
rect 1233 38672 1279 38711
rect 1233 38638 1239 38672
rect 1273 38638 1279 38672
rect 1233 38599 1279 38638
rect 1233 38565 1239 38599
rect 1273 38565 1279 38599
rect 1233 38526 1279 38565
rect 1233 38492 1239 38526
rect 1273 38492 1279 38526
tri 1043 38472 1059 38488 sw
tri 1217 38472 1233 38488 se
rect 1233 38472 1279 38492
rect 1469 38964 1515 38976
rect 1469 38930 1475 38964
rect 1509 38930 1515 38964
rect 1469 38891 1515 38930
rect 1469 38857 1475 38891
rect 1509 38857 1515 38891
rect 1469 38818 1515 38857
rect 1469 38784 1475 38818
rect 1509 38784 1515 38818
rect 1469 38745 1515 38784
rect 1469 38711 1475 38745
rect 1509 38711 1515 38745
rect 1469 38672 1515 38711
rect 1469 38638 1475 38672
rect 1509 38638 1515 38672
rect 1469 38599 1515 38638
rect 1469 38565 1475 38599
rect 1509 38565 1515 38599
rect 1469 38526 1515 38565
rect 1469 38492 1475 38526
rect 1509 38492 1515 38526
tri 1279 38472 1295 38488 sw
tri 1453 38472 1469 38488 se
rect 1469 38472 1515 38492
rect 1705 38964 1751 38976
rect 1705 38930 1711 38964
rect 1745 38930 1751 38964
rect 1705 38891 1751 38930
rect 1705 38857 1711 38891
rect 1745 38857 1751 38891
rect 1705 38818 1751 38857
rect 1705 38784 1711 38818
rect 1745 38784 1751 38818
rect 1705 38745 1751 38784
rect 1705 38711 1711 38745
rect 1745 38711 1751 38745
rect 1705 38672 1751 38711
rect 1705 38638 1711 38672
rect 1745 38638 1751 38672
rect 1705 38599 1751 38638
rect 1705 38565 1711 38599
rect 1745 38565 1751 38599
rect 1705 38526 1751 38565
rect 1705 38492 1711 38526
rect 1745 38492 1751 38526
tri 1515 38472 1531 38488 sw
tri 1689 38472 1705 38488 se
rect 1705 38472 1751 38492
rect 1941 38964 1987 38976
rect 1941 38930 1947 38964
rect 1981 38930 1987 38964
rect 1941 38891 1987 38930
rect 1941 38857 1947 38891
rect 1981 38857 1987 38891
rect 1941 38818 1987 38857
rect 1941 38784 1947 38818
rect 1981 38784 1987 38818
rect 1941 38745 1987 38784
rect 1941 38711 1947 38745
rect 1981 38711 1987 38745
rect 1941 38672 1987 38711
rect 1941 38638 1947 38672
rect 1981 38638 1987 38672
rect 1941 38599 1987 38638
rect 1941 38565 1947 38599
rect 1981 38565 1987 38599
rect 1941 38526 1987 38565
rect 1941 38492 1947 38526
rect 1981 38492 1987 38526
tri 1751 38472 1767 38488 sw
tri 1925 38472 1941 38488 se
rect 1941 38472 1987 38492
rect 2177 38964 2223 38976
rect 2177 38930 2183 38964
rect 2217 38930 2223 38964
rect 2177 38891 2223 38930
rect 2177 38857 2183 38891
rect 2217 38857 2223 38891
rect 2177 38818 2223 38857
rect 2177 38784 2183 38818
rect 2217 38784 2223 38818
rect 2177 38745 2223 38784
rect 2177 38711 2183 38745
rect 2217 38711 2223 38745
rect 2177 38672 2223 38711
rect 2177 38638 2183 38672
rect 2217 38638 2223 38672
rect 2177 38599 2223 38638
rect 2177 38565 2183 38599
rect 2217 38565 2223 38599
rect 2177 38526 2223 38565
rect 2177 38492 2183 38526
rect 2217 38492 2223 38526
tri 1987 38472 2003 38488 sw
tri 2161 38472 2177 38488 se
rect 2177 38472 2223 38492
rect 2413 38964 2459 38976
rect 2413 38930 2419 38964
rect 2453 38930 2459 38964
rect 2413 38891 2459 38930
rect 2413 38857 2419 38891
rect 2453 38857 2459 38891
rect 2413 38818 2459 38857
rect 2413 38784 2419 38818
rect 2453 38784 2459 38818
rect 2413 38745 2459 38784
rect 2413 38711 2419 38745
rect 2453 38711 2459 38745
rect 2413 38672 2459 38711
rect 2413 38638 2419 38672
rect 2453 38638 2459 38672
rect 2413 38599 2459 38638
rect 2413 38565 2419 38599
rect 2453 38565 2459 38599
rect 2413 38526 2459 38565
rect 2413 38492 2419 38526
rect 2453 38492 2459 38526
tri 2223 38472 2239 38488 sw
tri 2397 38472 2413 38488 se
rect 2413 38472 2459 38492
rect 2649 38964 2695 38976
rect 2649 38930 2655 38964
rect 2689 38930 2695 38964
rect 2649 38891 2695 38930
rect 2649 38857 2655 38891
rect 2689 38857 2695 38891
rect 2649 38818 2695 38857
rect 2649 38784 2655 38818
rect 2689 38784 2695 38818
rect 2649 38745 2695 38784
rect 2649 38711 2655 38745
rect 2689 38711 2695 38745
rect 2649 38672 2695 38711
rect 2649 38638 2655 38672
rect 2689 38638 2695 38672
rect 2649 38599 2695 38638
rect 2649 38565 2655 38599
rect 2689 38565 2695 38599
rect 2649 38526 2695 38565
rect 2649 38492 2655 38526
rect 2689 38492 2695 38526
tri 2459 38472 2475 38488 sw
tri 2633 38472 2649 38488 se
rect 2649 38472 2695 38492
rect 2885 38964 3076 39000
rect 2885 38930 2891 38964
rect 2925 38962 3076 38964
rect 2925 38930 3036 38962
rect 2885 38928 3036 38930
rect 3070 38928 3076 38962
rect 2885 38891 3076 38928
rect 2885 38857 2891 38891
rect 2925 38890 3076 38891
rect 2925 38857 3036 38890
rect 2885 38856 3036 38857
rect 3070 38856 3076 38890
rect 2885 38818 3076 38856
rect 2885 38784 2891 38818
rect 2925 38784 3036 38818
rect 3070 38784 3076 38818
rect 2885 38746 3076 38784
rect 2885 38745 3036 38746
rect 2885 38711 2891 38745
rect 2925 38712 3036 38745
rect 3070 38712 3076 38746
rect 2925 38711 3076 38712
rect 2885 38674 3076 38711
rect 2885 38672 3036 38674
rect 2885 38638 2891 38672
rect 2925 38640 3036 38672
rect 3070 38640 3076 38674
rect 2925 38638 3076 38640
rect 2885 38602 3076 38638
rect 2885 38599 3036 38602
rect 2885 38565 2891 38599
rect 2925 38568 3036 38599
rect 3070 38568 3076 38602
rect 2925 38565 3076 38568
rect 2885 38530 3076 38565
rect 2885 38526 3036 38530
rect 2885 38492 2891 38526
rect 2925 38496 3036 38526
rect 3070 38496 3076 38530
rect 2925 38492 3076 38496
tri 2695 38472 2711 38488 sw
tri 2869 38472 2885 38488 se
rect 2885 38472 3076 38492
rect 380 38458 587 38472
tri 587 38458 601 38472 sw
tri 731 38458 745 38472 se
rect 745 38458 823 38472
tri 823 38458 837 38472 sw
tri 967 38458 981 38472 se
rect 981 38458 1059 38472
tri 1059 38458 1073 38472 sw
tri 1203 38458 1217 38472 se
rect 1217 38458 1295 38472
tri 1295 38458 1309 38472 sw
tri 1439 38458 1453 38472 se
rect 1453 38458 1531 38472
tri 1531 38458 1545 38472 sw
tri 1675 38458 1689 38472 se
rect 1689 38458 1767 38472
tri 1767 38458 1781 38472 sw
tri 1911 38458 1925 38472 se
rect 1925 38458 2003 38472
tri 2003 38458 2017 38472 sw
tri 2147 38458 2161 38472 se
rect 2161 38458 2239 38472
tri 2239 38458 2253 38472 sw
tri 2383 38458 2397 38472 se
rect 2397 38458 2475 38472
tri 2475 38458 2489 38472 sw
tri 2619 38458 2633 38472 se
rect 2633 38458 2711 38472
tri 2711 38458 2725 38472 sw
tri 2855 38458 2869 38472 se
rect 2869 38458 3076 38472
rect 380 38454 601 38458
tri 601 38454 605 38458 sw
tri 727 38454 731 38458 se
rect 731 38454 837 38458
tri 837 38454 841 38458 sw
tri 963 38454 967 38458 se
rect 967 38454 1073 38458
tri 1073 38454 1077 38458 sw
tri 1199 38454 1203 38458 se
rect 1203 38454 1309 38458
tri 1309 38454 1313 38458 sw
tri 1435 38454 1439 38458 se
rect 1439 38454 1545 38458
tri 1545 38454 1549 38458 sw
tri 1671 38454 1675 38458 se
rect 1675 38454 1781 38458
tri 1781 38454 1785 38458 sw
tri 1907 38454 1911 38458 se
rect 1911 38454 2017 38458
tri 2017 38454 2021 38458 sw
tri 2143 38454 2147 38458 se
rect 2147 38454 2253 38458
tri 2253 38454 2257 38458 sw
tri 2379 38454 2383 38458 se
rect 2383 38454 2489 38458
tri 2489 38454 2493 38458 sw
tri 2615 38454 2619 38458 se
rect 2619 38454 2725 38458
tri 2725 38454 2729 38458 sw
tri 2851 38454 2855 38458 se
rect 2855 38454 3036 38458
rect 380 38453 3036 38454
rect 380 38449 531 38453
rect 380 38415 386 38449
rect 420 38419 531 38449
rect 565 38423 767 38453
rect 801 38423 1003 38453
rect 1037 38423 1239 38453
rect 1273 38423 1475 38453
rect 565 38419 697 38423
rect 420 38415 697 38419
rect 380 38380 697 38415
rect 380 38376 531 38380
rect 380 38342 386 38376
rect 420 38346 531 38376
rect 565 38371 697 38380
rect 749 38371 765 38423
rect 817 38371 833 38423
rect 885 38371 901 38423
rect 953 38371 969 38423
rect 1021 38380 1037 38419
rect 1089 38371 1105 38423
rect 1157 38371 1173 38423
rect 1225 38419 1239 38423
rect 1293 38419 1475 38423
rect 1509 38419 1711 38453
rect 1745 38419 1947 38453
rect 1981 38423 2183 38453
rect 2217 38423 2419 38453
rect 2453 38423 2655 38453
rect 2689 38423 2891 38453
rect 1981 38419 2097 38423
rect 1225 38380 1241 38419
rect 1293 38380 2097 38419
rect 1225 38371 1239 38380
rect 1293 38371 1475 38380
rect 565 38359 767 38371
rect 801 38359 1003 38371
rect 1037 38359 1239 38371
rect 1273 38359 1475 38371
rect 565 38346 697 38359
rect 420 38342 697 38346
rect 380 38307 697 38342
rect 749 38307 765 38359
rect 817 38307 833 38359
rect 885 38307 901 38359
rect 953 38307 969 38359
rect 1021 38307 1037 38346
rect 1089 38307 1105 38359
rect 1157 38307 1173 38359
rect 1225 38346 1239 38359
rect 1293 38346 1475 38359
rect 1509 38346 1711 38380
rect 1745 38346 1947 38380
rect 1981 38371 2097 38380
rect 2149 38371 2165 38423
rect 2217 38371 2233 38423
rect 2285 38371 2301 38423
rect 2353 38371 2369 38423
rect 2421 38380 2437 38419
rect 2489 38371 2505 38423
rect 2557 38371 2573 38423
rect 2625 38371 2641 38423
rect 2693 38419 2891 38423
rect 2925 38424 3036 38453
rect 3070 38424 3076 38458
rect 2925 38419 3076 38424
rect 2693 38386 3076 38419
rect 2693 38380 3036 38386
rect 2693 38371 2891 38380
rect 1981 38359 2183 38371
rect 2217 38359 2419 38371
rect 2453 38359 2655 38371
rect 2689 38359 2891 38371
rect 1981 38346 2097 38359
rect 1225 38307 1241 38346
rect 1293 38307 2097 38346
rect 2149 38307 2165 38359
rect 2217 38307 2233 38359
rect 2285 38307 2301 38359
rect 2353 38307 2369 38359
rect 2421 38307 2437 38346
rect 2489 38307 2505 38359
rect 2557 38307 2573 38359
rect 2625 38307 2641 38359
rect 2693 38346 2891 38359
rect 2925 38352 3036 38380
rect 3070 38352 3076 38386
rect 2925 38346 3076 38352
rect 2693 38314 3076 38346
rect 2693 38307 3036 38314
rect 380 38303 531 38307
rect 380 38269 386 38303
rect 420 38273 531 38303
rect 565 38295 767 38307
rect 801 38295 1003 38307
rect 1037 38295 1239 38307
rect 1273 38295 1475 38307
rect 565 38273 697 38295
rect 420 38269 697 38273
rect 380 38243 697 38269
rect 749 38243 765 38295
rect 817 38243 833 38295
rect 885 38243 901 38295
rect 953 38243 969 38295
rect 1021 38243 1037 38273
rect 1089 38243 1105 38295
rect 1157 38243 1173 38295
rect 1225 38273 1239 38295
rect 1293 38273 1475 38295
rect 1509 38273 1711 38307
rect 1745 38273 1947 38307
rect 1981 38295 2183 38307
rect 2217 38295 2419 38307
rect 2453 38295 2655 38307
rect 2689 38295 2891 38307
rect 1981 38273 2097 38295
rect 1225 38243 1241 38273
rect 1293 38243 2097 38273
rect 2149 38243 2165 38295
rect 2217 38243 2233 38295
rect 2285 38243 2301 38295
rect 2353 38243 2369 38295
rect 2421 38243 2437 38273
rect 2489 38243 2505 38295
rect 2557 38243 2573 38295
rect 2625 38243 2641 38295
rect 2693 38273 2891 38295
rect 2925 38280 3036 38307
rect 3070 38280 3076 38314
rect 2925 38273 3076 38280
rect 2693 38243 3076 38273
rect 380 38242 3076 38243
rect 380 38234 3036 38242
rect 380 38230 531 38234
rect 380 38196 386 38230
rect 420 38200 531 38230
rect 565 38231 767 38234
rect 801 38231 1003 38234
rect 1037 38231 1239 38234
rect 1273 38231 1475 38234
rect 565 38200 697 38231
rect 420 38196 697 38200
rect 380 38179 697 38196
rect 749 38179 765 38231
rect 817 38179 833 38231
rect 885 38179 901 38231
rect 953 38179 969 38231
rect 1021 38179 1037 38200
rect 1089 38179 1105 38231
rect 1157 38179 1173 38231
rect 1225 38200 1239 38231
rect 1293 38200 1475 38231
rect 1509 38200 1711 38234
rect 1745 38200 1947 38234
rect 1981 38231 2183 38234
rect 2217 38231 2419 38234
rect 2453 38231 2655 38234
rect 2689 38231 2891 38234
rect 1981 38200 2097 38231
rect 1225 38179 1241 38200
rect 1293 38179 2097 38200
rect 2149 38179 2165 38231
rect 2217 38179 2233 38231
rect 2285 38179 2301 38231
rect 2353 38179 2369 38231
rect 2421 38179 2437 38200
rect 2489 38179 2505 38231
rect 2557 38179 2573 38231
rect 2625 38179 2641 38231
rect 2693 38200 2891 38231
rect 2925 38208 3036 38234
rect 3070 38208 3076 38242
rect 2925 38200 3076 38208
rect 2693 38179 3076 38200
rect 380 38170 3076 38179
rect 380 38167 3036 38170
rect 380 38161 697 38167
rect 380 38157 531 38161
rect 380 38123 386 38157
rect 420 38127 531 38157
rect 565 38127 697 38161
rect 420 38123 697 38127
rect 380 38115 697 38123
rect 749 38115 765 38167
rect 817 38115 833 38167
rect 885 38115 901 38167
rect 953 38115 969 38167
rect 1021 38161 1037 38167
rect 1021 38115 1037 38127
rect 1089 38115 1105 38167
rect 1157 38115 1173 38167
rect 1225 38161 1241 38167
rect 1293 38161 2097 38167
rect 1225 38127 1239 38161
rect 1293 38127 1475 38161
rect 1509 38127 1711 38161
rect 1745 38127 1947 38161
rect 1981 38127 2097 38161
rect 1225 38115 1241 38127
rect 1293 38115 2097 38127
rect 2149 38115 2165 38167
rect 2217 38115 2233 38167
rect 2285 38115 2301 38167
rect 2353 38115 2369 38167
rect 2421 38161 2437 38167
rect 2421 38115 2437 38127
rect 2489 38115 2505 38167
rect 2557 38115 2573 38167
rect 2625 38115 2641 38167
rect 2693 38161 3036 38167
rect 2693 38127 2891 38161
rect 2925 38136 3036 38161
rect 3070 38136 3076 38170
rect 2925 38127 3076 38136
rect 2693 38115 3076 38127
rect 380 38103 3076 38115
rect 380 38088 697 38103
rect 380 38084 531 38088
rect 380 38050 386 38084
rect 420 38054 531 38084
rect 565 38054 697 38088
rect 420 38051 697 38054
rect 749 38051 765 38103
rect 817 38051 833 38103
rect 885 38051 901 38103
rect 953 38051 969 38103
rect 1021 38088 1037 38103
rect 1021 38051 1037 38054
rect 1089 38051 1105 38103
rect 1157 38051 1173 38103
rect 1225 38088 1241 38103
rect 1293 38088 2097 38103
rect 1225 38054 1239 38088
rect 1293 38054 1475 38088
rect 1509 38054 1711 38088
rect 1745 38054 1947 38088
rect 1981 38054 2097 38088
rect 1225 38051 1241 38054
rect 1293 38051 2097 38054
rect 2149 38051 2165 38103
rect 2217 38051 2233 38103
rect 2285 38051 2301 38103
rect 2353 38051 2369 38103
rect 2421 38088 2437 38103
rect 2421 38051 2437 38054
rect 2489 38051 2505 38103
rect 2557 38051 2573 38103
rect 2625 38051 2641 38103
rect 2693 38098 3076 38103
rect 2693 38088 3036 38098
rect 2693 38054 2891 38088
rect 2925 38064 3036 38088
rect 3070 38064 3076 38098
rect 2925 38054 3076 38064
rect 2693 38051 3076 38054
rect 420 38050 3076 38051
rect 380 38039 3076 38050
rect 380 38014 697 38039
rect 380 38011 531 38014
rect 380 37977 386 38011
rect 420 37980 531 38011
rect 565 37987 697 38014
rect 749 37987 765 38039
rect 817 37987 833 38039
rect 885 37987 901 38039
rect 953 37987 969 38039
rect 1021 38014 1037 38039
rect 1089 37987 1105 38039
rect 1157 37987 1173 38039
rect 1225 38014 1241 38039
rect 1293 38014 2097 38039
rect 1225 37987 1239 38014
rect 1293 37987 1475 38014
rect 565 37980 767 37987
rect 801 37980 1003 37987
rect 1037 37980 1239 37987
rect 1273 37980 1475 37987
rect 1509 37980 1711 38014
rect 1745 37980 1947 38014
rect 1981 37987 2097 38014
rect 2149 37987 2165 38039
rect 2217 37987 2233 38039
rect 2285 37987 2301 38039
rect 2353 37987 2369 38039
rect 2421 38014 2437 38039
rect 2489 37987 2505 38039
rect 2557 37987 2573 38039
rect 2625 37987 2641 38039
rect 2693 38026 3076 38039
rect 2693 38014 3036 38026
rect 2693 37987 2891 38014
rect 1981 37980 2183 37987
rect 2217 37980 2419 37987
rect 2453 37980 2655 37987
rect 2689 37980 2891 37987
rect 2925 37992 3036 38014
rect 3070 37992 3076 38026
rect 2925 37980 3076 37992
rect 420 37977 3076 37980
rect 380 37975 3076 37977
rect 380 37940 697 37975
rect 380 37938 531 37940
rect 380 37904 386 37938
rect 420 37906 531 37938
rect 565 37923 697 37940
rect 749 37923 765 37975
rect 817 37923 833 37975
rect 885 37923 901 37975
rect 953 37923 969 37975
rect 1021 37940 1037 37975
rect 1089 37923 1105 37975
rect 1157 37923 1173 37975
rect 1225 37940 1241 37975
rect 1293 37940 2097 37975
rect 1225 37923 1239 37940
rect 1293 37923 1475 37940
rect 565 37911 767 37923
rect 801 37911 1003 37923
rect 1037 37911 1239 37923
rect 1273 37911 1475 37923
rect 565 37906 697 37911
rect 420 37904 697 37906
rect 380 37866 697 37904
rect 380 37865 531 37866
rect 380 37831 386 37865
rect 420 37832 531 37865
rect 565 37859 697 37866
rect 749 37859 765 37911
rect 817 37859 833 37911
rect 885 37859 901 37911
rect 953 37859 969 37911
rect 1021 37866 1037 37906
rect 1089 37859 1105 37911
rect 1157 37859 1173 37911
rect 1225 37906 1239 37911
rect 1293 37906 1475 37911
rect 1509 37906 1711 37940
rect 1745 37906 1947 37940
rect 1981 37923 2097 37940
rect 2149 37923 2165 37975
rect 2217 37923 2233 37975
rect 2285 37923 2301 37975
rect 2353 37923 2369 37975
rect 2421 37940 2437 37975
rect 2489 37923 2505 37975
rect 2557 37923 2573 37975
rect 2625 37923 2641 37975
rect 2693 37954 3076 37975
rect 2693 37940 3036 37954
rect 2693 37923 2891 37940
rect 1981 37911 2183 37923
rect 2217 37911 2419 37923
rect 2453 37911 2655 37923
rect 2689 37911 2891 37923
rect 1981 37906 2097 37911
rect 1225 37866 1241 37906
rect 1293 37866 2097 37906
rect 1225 37859 1239 37866
rect 1293 37859 1475 37866
rect 565 37847 767 37859
rect 801 37847 1003 37859
rect 1037 37847 1239 37859
rect 1273 37847 1475 37859
rect 565 37832 697 37847
rect 420 37831 697 37832
rect 380 37795 697 37831
rect 749 37795 765 37847
rect 817 37795 833 37847
rect 885 37795 901 37847
rect 953 37795 969 37847
rect 1021 37795 1037 37832
rect 1089 37795 1105 37847
rect 1157 37795 1173 37847
rect 1225 37832 1239 37847
rect 1293 37832 1475 37847
rect 1509 37832 1711 37866
rect 1745 37832 1947 37866
rect 1981 37859 2097 37866
rect 2149 37859 2165 37911
rect 2217 37859 2233 37911
rect 2285 37859 2301 37911
rect 2353 37859 2369 37911
rect 2421 37866 2437 37906
rect 2489 37859 2505 37911
rect 2557 37859 2573 37911
rect 2625 37859 2641 37911
rect 2693 37906 2891 37911
rect 2925 37920 3036 37940
rect 3070 37920 3076 37954
rect 2925 37906 3076 37920
rect 2693 37882 3076 37906
rect 2693 37866 3036 37882
rect 2693 37859 2891 37866
rect 1981 37847 2183 37859
rect 2217 37847 2419 37859
rect 2453 37847 2655 37859
rect 2689 37847 2891 37859
rect 1981 37832 2097 37847
rect 1225 37795 1241 37832
rect 1293 37795 2097 37832
rect 2149 37795 2165 37847
rect 2217 37795 2233 37847
rect 2285 37795 2301 37847
rect 2353 37795 2369 37847
rect 2421 37795 2437 37832
rect 2489 37795 2505 37847
rect 2557 37795 2573 37847
rect 2625 37795 2641 37847
rect 2693 37832 2891 37847
rect 2925 37848 3036 37866
rect 3070 37848 3076 37882
rect 2925 37832 3076 37848
rect 2693 37810 3076 37832
rect 2693 37795 3036 37810
rect 380 37792 3036 37795
rect 380 37758 386 37792
rect 420 37758 531 37792
rect 565 37783 767 37792
rect 801 37783 1003 37792
rect 1037 37783 1239 37792
rect 1273 37783 1475 37792
rect 565 37758 697 37783
rect 380 37731 697 37758
rect 749 37731 765 37783
rect 817 37731 833 37783
rect 885 37731 901 37783
rect 953 37731 969 37783
rect 1021 37731 1037 37758
rect 1089 37731 1105 37783
rect 1157 37731 1173 37783
rect 1225 37758 1239 37783
rect 1293 37758 1475 37783
rect 1509 37758 1711 37792
rect 1745 37758 1947 37792
rect 1981 37783 2183 37792
rect 2217 37783 2419 37792
rect 2453 37783 2655 37792
rect 2689 37783 2891 37792
rect 1981 37758 2097 37783
rect 1225 37731 1241 37758
rect 1293 37731 2097 37758
rect 2149 37731 2165 37783
rect 2217 37731 2233 37783
rect 2285 37731 2301 37783
rect 2353 37731 2369 37783
rect 2421 37731 2437 37758
rect 2489 37731 2505 37783
rect 2557 37731 2573 37783
rect 2625 37731 2641 37783
rect 2693 37758 2891 37783
rect 2925 37776 3036 37792
rect 3070 37776 3076 37810
rect 2925 37758 3076 37776
rect 2693 37738 3076 37758
rect 2693 37731 3036 37738
rect 380 37719 3036 37731
rect 380 37685 386 37719
rect 420 37718 697 37719
rect 420 37685 531 37718
rect 380 37684 531 37685
rect 565 37684 697 37718
rect 380 37667 697 37684
rect 749 37667 765 37719
rect 817 37667 833 37719
rect 885 37667 901 37719
rect 953 37667 969 37719
rect 1021 37718 1037 37719
rect 1021 37667 1037 37684
rect 1089 37667 1105 37719
rect 1157 37667 1173 37719
rect 1225 37718 1241 37719
rect 1293 37718 2097 37719
rect 1225 37684 1239 37718
rect 1293 37684 1475 37718
rect 1509 37684 1711 37718
rect 1745 37684 1947 37718
rect 1981 37684 2097 37718
rect 1225 37667 1241 37684
rect 1293 37667 2097 37684
rect 2149 37667 2165 37719
rect 2217 37667 2233 37719
rect 2285 37667 2301 37719
rect 2353 37667 2369 37719
rect 2421 37718 2437 37719
rect 2421 37667 2437 37684
rect 2489 37667 2505 37719
rect 2557 37667 2573 37719
rect 2625 37667 2641 37719
rect 2693 37718 3036 37719
rect 2693 37684 2891 37718
rect 2925 37704 3036 37718
rect 3070 37704 3076 37738
rect 2925 37684 3076 37704
rect 2693 37667 3076 37684
rect 380 37666 3076 37667
rect 380 37655 3036 37666
rect 380 37647 697 37655
rect 380 37613 386 37647
rect 420 37644 697 37647
rect 420 37613 531 37644
rect 380 37610 531 37613
rect 565 37610 697 37644
rect 380 37603 697 37610
rect 749 37603 765 37655
rect 817 37603 833 37655
rect 885 37603 901 37655
rect 953 37603 969 37655
rect 1021 37644 1037 37655
rect 1021 37603 1037 37610
rect 1089 37603 1105 37655
rect 1157 37603 1173 37655
rect 1225 37644 1241 37655
rect 1293 37644 2097 37655
rect 1225 37610 1239 37644
rect 1293 37610 1475 37644
rect 1509 37610 1711 37644
rect 1745 37610 1947 37644
rect 1981 37610 2097 37644
rect 1225 37603 1241 37610
rect 1293 37603 2097 37610
rect 2149 37603 2165 37655
rect 2217 37603 2233 37655
rect 2285 37603 2301 37655
rect 2353 37603 2369 37655
rect 2421 37644 2437 37655
rect 2421 37603 2437 37610
rect 2489 37603 2505 37655
rect 2557 37603 2573 37655
rect 2625 37603 2641 37655
rect 2693 37644 3036 37655
rect 2693 37610 2891 37644
rect 2925 37632 3036 37644
rect 3070 37632 3076 37666
rect 2925 37610 3076 37632
rect 2693 37603 3076 37610
rect 380 37594 3076 37603
rect 380 37591 3036 37594
rect 380 37575 697 37591
rect 380 37541 386 37575
rect 420 37570 697 37575
rect 420 37541 531 37570
rect 380 37536 531 37541
rect 565 37539 697 37570
rect 749 37539 765 37591
rect 817 37539 833 37591
rect 885 37539 901 37591
rect 953 37539 969 37591
rect 1021 37570 1037 37591
rect 1089 37539 1105 37591
rect 1157 37539 1173 37591
rect 1225 37570 1241 37591
rect 1293 37570 2097 37591
rect 1225 37539 1239 37570
rect 1293 37539 1475 37570
rect 565 37536 767 37539
rect 801 37536 1003 37539
rect 1037 37536 1239 37539
rect 1273 37536 1475 37539
rect 1509 37536 1711 37570
rect 1745 37536 1947 37570
rect 1981 37539 2097 37570
rect 2149 37539 2165 37591
rect 2217 37539 2233 37591
rect 2285 37539 2301 37591
rect 2353 37539 2369 37591
rect 2421 37570 2437 37591
rect 2489 37539 2505 37591
rect 2557 37539 2573 37591
rect 2625 37539 2641 37591
rect 2693 37570 3036 37591
rect 2693 37539 2891 37570
rect 1981 37536 2183 37539
rect 2217 37536 2419 37539
rect 2453 37536 2655 37539
rect 2689 37536 2891 37539
rect 2925 37560 3036 37570
rect 3070 37560 3076 37594
rect 2925 37536 3076 37560
rect 380 37527 3076 37536
rect 380 37503 697 37527
rect 380 37469 386 37503
rect 420 37496 697 37503
rect 420 37469 531 37496
rect 380 37462 531 37469
rect 565 37475 697 37496
rect 749 37475 765 37527
rect 817 37475 833 37527
rect 885 37475 901 37527
rect 953 37475 969 37527
rect 1021 37496 1037 37527
rect 1089 37475 1105 37527
rect 1157 37475 1173 37527
rect 1225 37496 1241 37527
rect 1293 37496 2097 37527
rect 1225 37475 1239 37496
rect 1293 37475 1475 37496
rect 565 37462 767 37475
rect 801 37462 1003 37475
rect 1037 37462 1239 37475
rect 1273 37462 1475 37475
rect 1509 37462 1711 37496
rect 1745 37462 1947 37496
rect 1981 37475 2097 37496
rect 2149 37475 2165 37527
rect 2217 37475 2233 37527
rect 2285 37475 2301 37527
rect 2353 37475 2369 37527
rect 2421 37496 2437 37527
rect 2489 37475 2505 37527
rect 2557 37475 2573 37527
rect 2625 37475 2641 37527
rect 2693 37522 3076 37527
rect 2693 37496 3036 37522
rect 2693 37475 2891 37496
rect 1981 37462 2183 37475
rect 2217 37462 2419 37475
rect 2453 37462 2655 37475
rect 2689 37462 2891 37475
rect 2925 37488 3036 37496
rect 3070 37488 3076 37522
rect 2925 37462 3076 37488
rect 380 37454 3076 37462
rect 380 37450 601 37454
tri 601 37450 605 37454 nw
tri 727 37450 731 37454 ne
rect 731 37450 837 37454
tri 837 37450 841 37454 nw
tri 963 37450 967 37454 ne
rect 967 37450 1073 37454
tri 1073 37450 1077 37454 nw
tri 1199 37450 1203 37454 ne
rect 1203 37450 1309 37454
tri 1309 37450 1313 37454 nw
tri 1435 37450 1439 37454 ne
rect 1439 37450 1545 37454
tri 1545 37450 1549 37454 nw
tri 1671 37450 1675 37454 ne
rect 1675 37450 1781 37454
tri 1781 37450 1785 37454 nw
tri 1907 37450 1911 37454 ne
rect 1911 37450 2017 37454
tri 2017 37450 2021 37454 nw
tri 2143 37450 2147 37454 ne
rect 2147 37450 2253 37454
tri 2253 37450 2257 37454 nw
tri 2379 37450 2383 37454 ne
rect 2383 37450 2489 37454
tri 2489 37450 2493 37454 nw
tri 2615 37450 2619 37454 ne
rect 2619 37450 2725 37454
tri 2725 37450 2729 37454 nw
tri 2851 37450 2855 37454 ne
rect 2855 37450 3076 37454
rect 380 37431 573 37450
rect 380 37397 386 37431
rect 420 37422 573 37431
tri 573 37422 601 37450 nw
tri 731 37422 759 37450 ne
rect 759 37422 809 37450
tri 809 37422 837 37450 nw
tri 967 37422 995 37450 ne
rect 995 37422 1045 37450
tri 1045 37422 1073 37450 nw
tri 1203 37422 1231 37450 ne
rect 1231 37422 1281 37450
tri 1281 37422 1309 37450 nw
tri 1439 37422 1467 37450 ne
rect 1467 37422 1517 37450
tri 1517 37422 1545 37450 nw
tri 1675 37422 1703 37450 ne
rect 1703 37422 1753 37450
tri 1753 37422 1781 37450 nw
tri 1911 37422 1939 37450 ne
rect 1939 37422 1989 37450
tri 1989 37422 2017 37450 nw
tri 2147 37422 2175 37450 ne
rect 2175 37422 2225 37450
tri 2225 37422 2253 37450 nw
tri 2383 37422 2411 37450 ne
rect 2411 37422 2461 37450
tri 2461 37422 2489 37450 nw
tri 2619 37422 2647 37450 ne
rect 2647 37422 2697 37450
tri 2697 37422 2725 37450 nw
tri 2855 37422 2883 37450 ne
rect 2883 37422 3036 37450
rect 420 37397 531 37422
rect 380 37388 531 37397
rect 565 37388 571 37422
tri 571 37420 573 37422 nw
tri 759 37420 761 37422 ne
rect 380 37359 571 37388
rect 380 37325 386 37359
rect 420 37348 571 37359
rect 420 37325 531 37348
rect 380 37314 531 37325
rect 565 37314 571 37348
rect 380 37287 571 37314
rect 380 37253 386 37287
rect 420 37274 571 37287
rect 420 37253 531 37274
rect 380 37240 531 37253
rect 565 37240 571 37274
rect 380 37215 571 37240
rect 380 37181 386 37215
rect 420 37200 571 37215
rect 420 37181 531 37200
rect 380 37166 531 37181
rect 565 37166 571 37200
rect 380 37143 571 37166
rect 380 37109 386 37143
rect 420 37126 571 37143
rect 420 37109 531 37126
rect 380 37092 531 37109
rect 565 37092 571 37126
rect 380 37071 571 37092
rect 380 37037 386 37071
rect 420 37052 571 37071
rect 420 37037 531 37052
rect 380 37018 531 37037
rect 565 37018 571 37052
rect 380 36999 571 37018
rect 761 37388 767 37422
rect 801 37388 807 37422
tri 807 37420 809 37422 nw
tri 995 37420 997 37422 ne
rect 761 37348 807 37388
rect 761 37314 767 37348
rect 801 37314 807 37348
rect 761 37274 807 37314
rect 761 37240 767 37274
rect 801 37240 807 37274
rect 761 37200 807 37240
rect 761 37166 767 37200
rect 801 37166 807 37200
rect 761 37126 807 37166
rect 761 37092 767 37126
rect 801 37092 807 37126
rect 761 37052 807 37092
rect 761 37018 767 37052
rect 801 37018 807 37052
rect 761 37006 807 37018
rect 997 37388 1003 37422
rect 1037 37388 1043 37422
tri 1043 37420 1045 37422 nw
tri 1231 37420 1233 37422 ne
rect 997 37348 1043 37388
rect 997 37314 1003 37348
rect 1037 37314 1043 37348
rect 997 37274 1043 37314
rect 997 37240 1003 37274
rect 1037 37240 1043 37274
rect 997 37200 1043 37240
rect 997 37166 1003 37200
rect 1037 37166 1043 37200
rect 997 37126 1043 37166
rect 997 37092 1003 37126
rect 1037 37092 1043 37126
rect 997 37052 1043 37092
rect 997 37018 1003 37052
rect 1037 37018 1043 37052
rect 997 37006 1043 37018
rect 1233 37388 1239 37422
rect 1273 37388 1279 37422
tri 1279 37420 1281 37422 nw
tri 1467 37420 1469 37422 ne
rect 1233 37348 1279 37388
rect 1233 37314 1239 37348
rect 1273 37314 1279 37348
rect 1233 37274 1279 37314
rect 1233 37240 1239 37274
rect 1273 37240 1279 37274
rect 1233 37200 1279 37240
rect 1233 37166 1239 37200
rect 1273 37166 1279 37200
rect 1233 37126 1279 37166
rect 1233 37092 1239 37126
rect 1273 37092 1279 37126
rect 1233 37052 1279 37092
rect 1233 37018 1239 37052
rect 1273 37018 1279 37052
rect 1233 37006 1279 37018
rect 1469 37388 1475 37422
rect 1509 37388 1515 37422
tri 1515 37420 1517 37422 nw
tri 1703 37420 1705 37422 ne
rect 1469 37348 1515 37388
rect 1469 37314 1475 37348
rect 1509 37314 1515 37348
rect 1469 37274 1515 37314
rect 1469 37240 1475 37274
rect 1509 37240 1515 37274
rect 1469 37200 1515 37240
rect 1469 37166 1475 37200
rect 1509 37166 1515 37200
rect 1469 37126 1515 37166
rect 1469 37092 1475 37126
rect 1509 37092 1515 37126
rect 1469 37052 1515 37092
rect 1469 37018 1475 37052
rect 1509 37018 1515 37052
rect 1469 37006 1515 37018
rect 1705 37388 1711 37422
rect 1745 37388 1751 37422
tri 1751 37420 1753 37422 nw
tri 1939 37420 1941 37422 ne
rect 1705 37348 1751 37388
rect 1705 37314 1711 37348
rect 1745 37314 1751 37348
rect 1705 37274 1751 37314
rect 1705 37240 1711 37274
rect 1745 37240 1751 37274
rect 1705 37200 1751 37240
rect 1705 37166 1711 37200
rect 1745 37166 1751 37200
rect 1705 37126 1751 37166
rect 1705 37092 1711 37126
rect 1745 37092 1751 37126
rect 1705 37052 1751 37092
rect 1705 37018 1711 37052
rect 1745 37018 1751 37052
rect 1705 37006 1751 37018
rect 1941 37388 1947 37422
rect 1981 37388 1987 37422
tri 1987 37420 1989 37422 nw
tri 2175 37420 2177 37422 ne
rect 1941 37348 1987 37388
rect 1941 37314 1947 37348
rect 1981 37314 1987 37348
rect 1941 37274 1987 37314
rect 1941 37240 1947 37274
rect 1981 37240 1987 37274
rect 1941 37200 1987 37240
rect 1941 37166 1947 37200
rect 1981 37166 1987 37200
rect 1941 37126 1987 37166
rect 1941 37092 1947 37126
rect 1981 37092 1987 37126
rect 1941 37052 1987 37092
rect 1941 37018 1947 37052
rect 1981 37018 1987 37052
rect 1941 37006 1987 37018
rect 2177 37388 2183 37422
rect 2217 37388 2223 37422
tri 2223 37420 2225 37422 nw
tri 2411 37420 2413 37422 ne
rect 2177 37348 2223 37388
rect 2177 37314 2183 37348
rect 2217 37314 2223 37348
rect 2177 37274 2223 37314
rect 2177 37240 2183 37274
rect 2217 37240 2223 37274
rect 2177 37200 2223 37240
rect 2177 37166 2183 37200
rect 2217 37166 2223 37200
rect 2177 37126 2223 37166
rect 2177 37092 2183 37126
rect 2217 37092 2223 37126
rect 2177 37052 2223 37092
rect 2177 37018 2183 37052
rect 2217 37018 2223 37052
rect 2177 37006 2223 37018
rect 2413 37388 2419 37422
rect 2453 37388 2459 37422
tri 2459 37420 2461 37422 nw
tri 2647 37420 2649 37422 ne
rect 2413 37348 2459 37388
rect 2413 37314 2419 37348
rect 2453 37314 2459 37348
rect 2413 37274 2459 37314
rect 2413 37240 2419 37274
rect 2453 37240 2459 37274
rect 2413 37200 2459 37240
rect 2413 37166 2419 37200
rect 2453 37166 2459 37200
rect 2413 37126 2459 37166
rect 2413 37092 2419 37126
rect 2453 37092 2459 37126
rect 2413 37052 2459 37092
rect 2413 37018 2419 37052
rect 2453 37018 2459 37052
rect 2413 37006 2459 37018
rect 2649 37388 2655 37422
rect 2689 37388 2695 37422
tri 2695 37420 2697 37422 nw
tri 2883 37420 2885 37422 ne
rect 2649 37348 2695 37388
rect 2649 37314 2655 37348
rect 2689 37314 2695 37348
rect 2649 37274 2695 37314
rect 2649 37240 2655 37274
rect 2689 37240 2695 37274
rect 2649 37200 2695 37240
rect 2649 37166 2655 37200
rect 2689 37166 2695 37200
rect 2649 37126 2695 37166
rect 2649 37092 2655 37126
rect 2689 37092 2695 37126
rect 2649 37052 2695 37092
rect 2649 37018 2655 37052
rect 2689 37018 2695 37052
rect 2649 37006 2695 37018
rect 2885 37388 2891 37422
rect 2925 37416 3036 37422
rect 3070 37416 3076 37450
rect 2925 37388 3076 37416
rect 2885 37378 3076 37388
rect 2885 37348 3036 37378
rect 2885 37314 2891 37348
rect 2925 37344 3036 37348
rect 3070 37344 3076 37378
rect 2925 37314 3076 37344
rect 2885 37306 3076 37314
rect 2885 37274 3036 37306
rect 2885 37240 2891 37274
rect 2925 37272 3036 37274
rect 3070 37272 3076 37306
rect 2925 37240 3076 37272
rect 2885 37234 3076 37240
rect 2885 37200 3036 37234
rect 3070 37200 3076 37234
rect 2885 37166 2891 37200
rect 2925 37166 3076 37200
rect 2885 37162 3076 37166
rect 2885 37128 3036 37162
rect 3070 37128 3076 37162
rect 2885 37126 3076 37128
rect 2885 37092 2891 37126
rect 2925 37092 3076 37126
rect 2885 37090 3076 37092
rect 2885 37056 3036 37090
rect 3070 37056 3076 37090
rect 2885 37052 3076 37056
rect 2885 37018 2891 37052
rect 2925 37018 3076 37052
rect 380 36965 386 36999
rect 420 36965 571 36999
rect 380 36927 571 36965
rect 2885 36984 3036 37018
rect 3070 36984 3076 37018
rect 2885 36946 3076 36984
rect 380 36893 386 36927
rect 420 36893 571 36927
rect 380 36855 571 36893
rect 613 36924 1501 36933
rect 1553 36924 1569 36933
rect 1621 36924 1636 36933
rect 1688 36924 1703 36933
rect 1755 36924 1770 36933
rect 1822 36924 1837 36933
rect 1889 36924 2830 36933
rect 613 36890 625 36924
rect 659 36890 700 36924
rect 734 36890 775 36924
rect 809 36890 850 36924
rect 884 36890 925 36924
rect 959 36890 1000 36924
rect 1034 36890 1075 36924
rect 1109 36890 1150 36924
rect 1184 36890 1225 36924
rect 1259 36890 1300 36924
rect 1334 36890 1375 36924
rect 1409 36890 1450 36924
rect 1484 36890 1501 36924
rect 1559 36890 1569 36924
rect 1634 36890 1636 36924
rect 1889 36890 1896 36924
rect 1930 36890 1970 36924
rect 2004 36890 2044 36924
rect 2078 36890 2118 36924
rect 2152 36890 2192 36924
rect 2226 36890 2266 36924
rect 2300 36890 2340 36924
rect 2374 36890 2414 36924
rect 2448 36890 2488 36924
rect 2522 36890 2562 36924
rect 2596 36890 2636 36924
rect 2670 36890 2710 36924
rect 2744 36890 2784 36924
rect 2818 36890 2830 36924
rect 613 36881 1501 36890
rect 1553 36881 1569 36890
rect 1621 36881 1636 36890
rect 1688 36881 1703 36890
rect 1755 36881 1770 36890
rect 1822 36881 1837 36890
rect 1889 36881 2830 36890
rect 2885 36912 3036 36946
rect 3070 36912 3076 36946
rect 380 36821 386 36855
rect 420 36822 571 36855
rect 2885 36874 3076 36912
rect 2885 36840 3036 36874
rect 3070 36840 3076 36874
rect 420 36821 531 36822
rect 380 36788 531 36821
rect 565 36788 571 36822
rect 380 36783 571 36788
rect 380 36749 386 36783
rect 420 36749 571 36783
rect 380 36715 531 36749
rect 565 36715 571 36749
rect 380 36711 571 36715
rect 380 36677 386 36711
rect 420 36677 571 36711
rect 380 36676 571 36677
rect 380 36642 531 36676
rect 565 36642 571 36676
rect 380 36639 571 36642
rect 380 36605 386 36639
rect 420 36605 571 36639
rect 380 36603 571 36605
rect 380 36569 531 36603
rect 565 36569 571 36603
rect 380 36567 571 36569
rect 380 36533 386 36567
rect 420 36533 571 36567
rect 380 36530 571 36533
rect 380 36496 531 36530
rect 565 36496 571 36530
rect 380 36495 571 36496
rect 380 36461 386 36495
rect 420 36461 571 36495
rect 380 36457 571 36461
rect 380 36423 531 36457
rect 565 36423 571 36457
rect 761 36822 807 36834
rect 761 36788 767 36822
rect 801 36788 807 36822
rect 761 36749 807 36788
rect 761 36715 767 36749
rect 801 36715 807 36749
rect 761 36676 807 36715
rect 761 36642 767 36676
rect 801 36642 807 36676
rect 761 36603 807 36642
rect 761 36569 767 36603
rect 801 36569 807 36603
rect 761 36530 807 36569
rect 761 36496 767 36530
rect 801 36496 807 36530
rect 761 36457 807 36496
tri 571 36423 575 36427 sw
tri 757 36423 761 36427 se
rect 761 36423 767 36457
rect 801 36423 807 36457
rect 997 36822 1043 36834
rect 997 36788 1003 36822
rect 1037 36788 1043 36822
rect 997 36749 1043 36788
rect 997 36715 1003 36749
rect 1037 36715 1043 36749
rect 997 36676 1043 36715
rect 997 36642 1003 36676
rect 1037 36642 1043 36676
rect 997 36603 1043 36642
rect 997 36569 1003 36603
rect 1037 36569 1043 36603
rect 997 36530 1043 36569
rect 997 36496 1003 36530
rect 1037 36496 1043 36530
rect 997 36457 1043 36496
tri 807 36423 811 36427 sw
tri 993 36423 997 36427 se
rect 997 36423 1003 36457
rect 1037 36423 1043 36457
rect 1233 36822 1279 36834
rect 1233 36788 1239 36822
rect 1273 36788 1279 36822
rect 1233 36749 1279 36788
rect 1233 36715 1239 36749
rect 1273 36715 1279 36749
rect 1233 36676 1279 36715
rect 1233 36642 1239 36676
rect 1273 36642 1279 36676
rect 1233 36603 1279 36642
rect 1233 36569 1239 36603
rect 1273 36569 1279 36603
rect 1233 36530 1279 36569
rect 1233 36496 1239 36530
rect 1273 36496 1279 36530
rect 1233 36457 1279 36496
tri 1043 36423 1047 36427 sw
tri 1229 36423 1233 36427 se
rect 1233 36423 1239 36457
rect 1273 36423 1279 36457
rect 1469 36822 1515 36834
rect 1469 36788 1475 36822
rect 1509 36788 1515 36822
rect 1469 36749 1515 36788
rect 1469 36715 1475 36749
rect 1509 36715 1515 36749
rect 1469 36676 1515 36715
rect 1469 36642 1475 36676
rect 1509 36642 1515 36676
rect 1469 36603 1515 36642
rect 1469 36569 1475 36603
rect 1509 36569 1515 36603
rect 1469 36530 1515 36569
rect 1469 36496 1475 36530
rect 1509 36496 1515 36530
rect 1469 36457 1515 36496
tri 1279 36423 1283 36427 sw
tri 1465 36423 1469 36427 se
rect 1469 36423 1475 36457
rect 1509 36423 1515 36457
rect 1705 36822 1751 36834
rect 1705 36788 1711 36822
rect 1745 36788 1751 36822
rect 1705 36749 1751 36788
rect 1705 36715 1711 36749
rect 1745 36715 1751 36749
rect 1705 36676 1751 36715
rect 1705 36642 1711 36676
rect 1745 36642 1751 36676
rect 1705 36603 1751 36642
rect 1705 36569 1711 36603
rect 1745 36569 1751 36603
rect 1705 36530 1751 36569
rect 1705 36496 1711 36530
rect 1745 36496 1751 36530
rect 1705 36457 1751 36496
tri 1515 36423 1519 36427 sw
tri 1701 36423 1705 36427 se
rect 1705 36423 1711 36457
rect 1745 36423 1751 36457
rect 1941 36822 1987 36834
rect 1941 36788 1947 36822
rect 1981 36788 1987 36822
rect 1941 36749 1987 36788
rect 1941 36715 1947 36749
rect 1981 36715 1987 36749
rect 1941 36676 1987 36715
rect 1941 36642 1947 36676
rect 1981 36642 1987 36676
rect 1941 36603 1987 36642
rect 1941 36569 1947 36603
rect 1981 36569 1987 36603
rect 1941 36530 1987 36569
rect 1941 36496 1947 36530
rect 1981 36496 1987 36530
rect 1941 36457 1987 36496
tri 1751 36423 1755 36427 sw
tri 1937 36423 1941 36427 se
rect 1941 36423 1947 36457
rect 1981 36423 1987 36457
rect 2177 36822 2223 36834
rect 2177 36788 2183 36822
rect 2217 36788 2223 36822
rect 2177 36749 2223 36788
rect 2177 36715 2183 36749
rect 2217 36715 2223 36749
rect 2177 36676 2223 36715
rect 2177 36642 2183 36676
rect 2217 36642 2223 36676
rect 2177 36603 2223 36642
rect 2177 36569 2183 36603
rect 2217 36569 2223 36603
rect 2177 36530 2223 36569
rect 2177 36496 2183 36530
rect 2217 36496 2223 36530
rect 2177 36457 2223 36496
tri 1987 36423 1991 36427 sw
tri 2173 36423 2177 36427 se
rect 2177 36423 2183 36457
rect 2217 36423 2223 36457
rect 2413 36822 2459 36834
rect 2413 36788 2419 36822
rect 2453 36788 2459 36822
rect 2413 36749 2459 36788
rect 2413 36715 2419 36749
rect 2453 36715 2459 36749
rect 2413 36676 2459 36715
rect 2413 36642 2419 36676
rect 2453 36642 2459 36676
rect 2413 36603 2459 36642
rect 2413 36569 2419 36603
rect 2453 36569 2459 36603
rect 2413 36530 2459 36569
rect 2413 36496 2419 36530
rect 2453 36496 2459 36530
rect 2413 36457 2459 36496
tri 2223 36423 2227 36427 sw
tri 2409 36423 2413 36427 se
rect 2413 36423 2419 36457
rect 2453 36423 2459 36457
rect 2649 36822 2695 36834
rect 2649 36788 2655 36822
rect 2689 36788 2695 36822
rect 2649 36749 2695 36788
rect 2649 36715 2655 36749
rect 2689 36715 2695 36749
rect 2649 36676 2695 36715
rect 2649 36642 2655 36676
rect 2689 36642 2695 36676
rect 2649 36603 2695 36642
rect 2649 36569 2655 36603
rect 2689 36569 2695 36603
rect 2649 36530 2695 36569
rect 2649 36496 2655 36530
rect 2689 36496 2695 36530
rect 2649 36457 2695 36496
tri 2459 36423 2463 36427 sw
tri 2645 36423 2649 36427 se
rect 2649 36423 2655 36457
rect 2689 36423 2695 36457
rect 2885 36822 3076 36840
rect 2885 36788 2891 36822
rect 2925 36802 3076 36822
rect 2925 36788 3036 36802
rect 2885 36768 3036 36788
rect 3070 36768 3076 36802
rect 2885 36749 3076 36768
rect 2885 36715 2891 36749
rect 2925 36730 3076 36749
rect 2925 36715 3036 36730
rect 2885 36696 3036 36715
rect 3070 36696 3076 36730
rect 2885 36676 3076 36696
rect 2885 36642 2891 36676
rect 2925 36658 3076 36676
rect 2925 36642 3036 36658
rect 2885 36624 3036 36642
rect 3070 36624 3076 36658
rect 2885 36603 3076 36624
rect 2885 36569 2891 36603
rect 2925 36586 3076 36603
rect 2925 36569 3036 36586
rect 2885 36552 3036 36569
rect 3070 36552 3076 36586
rect 2885 36530 3076 36552
rect 2885 36496 2891 36530
rect 2925 36514 3076 36530
rect 2925 36496 3036 36514
rect 2885 36480 3036 36496
rect 3070 36480 3076 36514
rect 2885 36457 3076 36480
tri 2695 36423 2699 36427 sw
tri 2881 36423 2885 36427 se
rect 2885 36423 2891 36457
rect 2925 36442 3076 36457
rect 2925 36423 3036 36442
rect 380 36389 386 36423
rect 420 36408 575 36423
tri 575 36408 590 36423 sw
tri 742 36408 757 36423 se
rect 757 36408 811 36423
tri 811 36408 826 36423 sw
tri 978 36408 993 36423 se
rect 993 36408 1047 36423
tri 1047 36408 1062 36423 sw
tri 1214 36408 1229 36423 se
rect 1229 36408 1283 36423
tri 1283 36408 1298 36423 sw
tri 1450 36408 1465 36423 se
rect 1465 36408 1519 36423
tri 1519 36408 1534 36423 sw
tri 1686 36408 1701 36423 se
rect 1701 36408 1755 36423
tri 1755 36408 1770 36423 sw
tri 1922 36408 1937 36423 se
rect 1937 36408 1991 36423
tri 1991 36408 2006 36423 sw
tri 2158 36408 2173 36423 se
rect 2173 36408 2227 36423
tri 2227 36408 2242 36423 sw
tri 2394 36408 2409 36423 se
rect 2409 36408 2463 36423
tri 2463 36408 2478 36423 sw
tri 2630 36408 2645 36423 se
rect 2645 36408 2699 36423
tri 2699 36408 2714 36423 sw
tri 2866 36408 2881 36423 se
rect 2881 36408 3036 36423
rect 3070 36408 3076 36442
rect 420 36393 590 36408
tri 590 36393 605 36408 sw
tri 727 36393 742 36408 se
rect 742 36393 826 36408
tri 826 36393 841 36408 sw
tri 963 36393 978 36408 se
rect 978 36393 1062 36408
tri 1062 36393 1077 36408 sw
tri 1199 36393 1214 36408 se
rect 1214 36393 1298 36408
tri 1298 36393 1313 36408 sw
tri 1435 36393 1450 36408 se
rect 1450 36393 1534 36408
tri 1534 36393 1549 36408 sw
tri 1671 36393 1686 36408 se
rect 1686 36393 1770 36408
tri 1770 36393 1785 36408 sw
tri 1907 36393 1922 36408 se
rect 1922 36393 2006 36408
tri 2006 36393 2021 36408 sw
tri 2143 36393 2158 36408 se
rect 2158 36393 2242 36408
tri 2242 36393 2257 36408 sw
tri 2379 36393 2394 36408 se
rect 2394 36393 2478 36408
tri 2478 36393 2493 36408 sw
tri 2615 36393 2630 36408 se
rect 2630 36393 2714 36408
tri 2714 36393 2729 36408 sw
tri 2851 36393 2866 36408 se
rect 2866 36393 3076 36408
rect 420 36389 3076 36393
rect 380 36384 3076 36389
rect 380 36351 531 36384
rect 380 36317 386 36351
rect 420 36350 531 36351
rect 565 36369 767 36384
rect 801 36369 1003 36384
rect 1037 36369 1239 36384
rect 1273 36369 1475 36384
rect 565 36350 697 36369
rect 420 36317 697 36350
rect 749 36317 765 36369
rect 817 36317 833 36369
rect 885 36317 901 36369
rect 953 36317 969 36369
rect 1021 36317 1037 36350
rect 1089 36317 1105 36369
rect 1157 36317 1173 36369
rect 1225 36350 1239 36369
rect 1293 36350 1475 36369
rect 1509 36350 1711 36384
rect 1745 36350 1947 36384
rect 1981 36369 2183 36384
rect 2217 36369 2419 36384
rect 2453 36369 2655 36384
rect 2689 36369 2891 36384
rect 1981 36350 2097 36369
rect 1225 36317 1241 36350
rect 1293 36317 2097 36350
rect 2149 36317 2165 36369
rect 2217 36317 2233 36369
rect 2285 36317 2301 36369
rect 2353 36317 2369 36369
rect 2421 36317 2437 36350
rect 2489 36317 2505 36369
rect 2557 36317 2573 36369
rect 2625 36317 2641 36369
rect 2693 36350 2891 36369
rect 2925 36370 3076 36384
rect 2925 36350 3036 36370
rect 2693 36336 3036 36350
rect 3070 36336 3076 36370
rect 2693 36317 3076 36336
rect 380 36311 3076 36317
rect 380 36279 531 36311
rect 380 36245 386 36279
rect 420 36277 531 36279
rect 565 36305 767 36311
rect 801 36305 1003 36311
rect 1037 36305 1239 36311
rect 1273 36305 1475 36311
rect 565 36277 697 36305
rect 420 36253 697 36277
rect 749 36253 765 36305
rect 817 36253 833 36305
rect 885 36253 901 36305
rect 953 36253 969 36305
rect 1021 36253 1037 36277
rect 1089 36253 1105 36305
rect 1157 36253 1173 36305
rect 1225 36277 1239 36305
rect 1293 36277 1475 36305
rect 1509 36277 1711 36311
rect 1745 36277 1947 36311
rect 1981 36305 2183 36311
rect 2217 36305 2419 36311
rect 2453 36305 2655 36311
rect 2689 36305 2891 36311
rect 1981 36277 2097 36305
rect 1225 36253 1241 36277
rect 1293 36253 2097 36277
rect 2149 36253 2165 36305
rect 2217 36253 2233 36305
rect 2285 36253 2301 36305
rect 2353 36253 2369 36305
rect 2421 36253 2437 36277
rect 2489 36253 2505 36305
rect 2557 36253 2573 36305
rect 2625 36253 2641 36305
rect 2693 36277 2891 36305
rect 2925 36298 3076 36311
rect 2925 36277 3036 36298
rect 2693 36264 3036 36277
rect 3070 36264 3076 36298
rect 2693 36253 3076 36264
rect 420 36245 3076 36253
rect 380 36241 3076 36245
rect 380 36238 697 36241
rect 380 36207 531 36238
rect 380 36173 386 36207
rect 420 36204 531 36207
rect 565 36204 697 36238
rect 420 36189 697 36204
rect 749 36189 765 36241
rect 817 36189 833 36241
rect 885 36189 901 36241
rect 953 36189 969 36241
rect 1021 36238 1037 36241
rect 1021 36189 1037 36204
rect 1089 36189 1105 36241
rect 1157 36189 1173 36241
rect 1225 36238 1241 36241
rect 1293 36238 2097 36241
rect 1225 36204 1239 36238
rect 1293 36204 1475 36238
rect 1509 36204 1711 36238
rect 1745 36204 1947 36238
rect 1981 36204 2097 36238
rect 1225 36189 1241 36204
rect 1293 36189 2097 36204
rect 2149 36189 2165 36241
rect 2217 36189 2233 36241
rect 2285 36189 2301 36241
rect 2353 36189 2369 36241
rect 2421 36238 2437 36241
rect 2421 36189 2437 36204
rect 2489 36189 2505 36241
rect 2557 36189 2573 36241
rect 2625 36189 2641 36241
rect 2693 36238 3076 36241
rect 2693 36204 2891 36238
rect 2925 36226 3076 36238
rect 2925 36204 3036 36226
rect 2693 36192 3036 36204
rect 3070 36192 3076 36226
rect 2693 36189 3076 36192
rect 420 36177 3076 36189
rect 420 36173 697 36177
rect 380 36165 697 36173
rect 380 36135 531 36165
rect 380 36101 386 36135
rect 420 36131 531 36135
rect 565 36131 697 36165
rect 420 36125 697 36131
rect 749 36125 765 36177
rect 817 36125 833 36177
rect 885 36125 901 36177
rect 953 36125 969 36177
rect 1021 36165 1037 36177
rect 1021 36125 1037 36131
rect 1089 36125 1105 36177
rect 1157 36125 1173 36177
rect 1225 36165 1241 36177
rect 1293 36165 2097 36177
rect 1225 36131 1239 36165
rect 1293 36131 1475 36165
rect 1509 36131 1711 36165
rect 1745 36131 1947 36165
rect 1981 36131 2097 36165
rect 1225 36125 1241 36131
rect 1293 36125 2097 36131
rect 2149 36125 2165 36177
rect 2217 36125 2233 36177
rect 2285 36125 2301 36177
rect 2353 36125 2369 36177
rect 2421 36165 2437 36177
rect 2421 36125 2437 36131
rect 2489 36125 2505 36177
rect 2557 36125 2573 36177
rect 2625 36125 2641 36177
rect 2693 36165 3076 36177
rect 2693 36131 2891 36165
rect 2925 36154 3076 36165
rect 2925 36131 3036 36154
rect 2693 36125 3036 36131
rect 420 36120 3036 36125
rect 3070 36120 3076 36154
rect 420 36113 3076 36120
rect 420 36101 697 36113
rect 380 36092 697 36101
rect 380 36063 531 36092
rect 380 36029 386 36063
rect 420 36058 531 36063
rect 565 36061 697 36092
rect 749 36061 765 36113
rect 817 36061 833 36113
rect 885 36061 901 36113
rect 953 36061 969 36113
rect 1021 36092 1037 36113
rect 1089 36061 1105 36113
rect 1157 36061 1173 36113
rect 1225 36092 1241 36113
rect 1293 36092 2097 36113
rect 1225 36061 1239 36092
rect 1293 36061 1475 36092
rect 565 36058 767 36061
rect 801 36058 1003 36061
rect 1037 36058 1239 36061
rect 1273 36058 1475 36061
rect 1509 36058 1711 36092
rect 1745 36058 1947 36092
rect 1981 36061 2097 36092
rect 2149 36061 2165 36113
rect 2217 36061 2233 36113
rect 2285 36061 2301 36113
rect 2353 36061 2369 36113
rect 2421 36092 2437 36113
rect 2489 36061 2505 36113
rect 2557 36061 2573 36113
rect 2625 36061 2641 36113
rect 2693 36092 3076 36113
rect 2693 36061 2891 36092
rect 1981 36058 2183 36061
rect 2217 36058 2419 36061
rect 2453 36058 2655 36061
rect 2689 36058 2891 36061
rect 2925 36082 3076 36092
rect 2925 36058 3036 36082
rect 420 36049 3036 36058
rect 420 36029 697 36049
rect 380 36019 697 36029
rect 380 35991 531 36019
rect 380 35957 386 35991
rect 420 35985 531 35991
rect 565 35997 697 36019
rect 749 35997 765 36049
rect 817 35997 833 36049
rect 885 35997 901 36049
rect 953 35997 969 36049
rect 1021 36019 1037 36049
rect 1089 35997 1105 36049
rect 1157 35997 1173 36049
rect 1225 36019 1241 36049
rect 1293 36019 2097 36049
rect 1225 35997 1239 36019
rect 1293 35997 1475 36019
rect 565 35985 767 35997
rect 801 35985 1003 35997
rect 1037 35985 1239 35997
rect 1273 35985 1475 35997
rect 1509 35985 1711 36019
rect 1745 35985 1947 36019
rect 1981 35997 2097 36019
rect 2149 35997 2165 36049
rect 2217 35997 2233 36049
rect 2285 35997 2301 36049
rect 2353 35997 2369 36049
rect 2421 36019 2437 36049
rect 2489 35997 2505 36049
rect 2557 35997 2573 36049
rect 2625 35997 2641 36049
rect 2693 36048 3036 36049
rect 3070 36048 3076 36082
rect 2693 36019 3076 36048
rect 2693 35997 2891 36019
rect 1981 35985 2183 35997
rect 2217 35985 2419 35997
rect 2453 35985 2655 35997
rect 2689 35985 2891 35997
rect 2925 36010 3076 36019
rect 2925 35985 3036 36010
rect 420 35957 697 35985
rect 380 35946 697 35957
rect 380 35919 531 35946
rect 380 35885 386 35919
rect 420 35912 531 35919
rect 565 35933 697 35946
rect 749 35933 765 35985
rect 817 35933 833 35985
rect 885 35933 901 35985
rect 953 35933 969 35985
rect 1021 35946 1037 35985
rect 1089 35933 1105 35985
rect 1157 35933 1173 35985
rect 1225 35946 1241 35985
rect 1293 35946 2097 35985
rect 1225 35933 1239 35946
rect 1293 35933 1475 35946
rect 565 35921 767 35933
rect 801 35921 1003 35933
rect 1037 35921 1239 35933
rect 1273 35921 1475 35933
rect 565 35912 697 35921
rect 420 35885 697 35912
rect 380 35872 697 35885
rect 380 35847 531 35872
rect 380 35813 386 35847
rect 420 35838 531 35847
rect 565 35869 697 35872
rect 749 35869 765 35921
rect 817 35869 833 35921
rect 885 35869 901 35921
rect 953 35869 969 35921
rect 1021 35872 1037 35912
rect 1089 35869 1105 35921
rect 1157 35869 1173 35921
rect 1225 35912 1239 35921
rect 1293 35912 1475 35921
rect 1509 35912 1711 35946
rect 1745 35912 1947 35946
rect 1981 35933 2097 35946
rect 2149 35933 2165 35985
rect 2217 35933 2233 35985
rect 2285 35933 2301 35985
rect 2353 35933 2369 35985
rect 2421 35946 2437 35985
rect 2489 35933 2505 35985
rect 2557 35933 2573 35985
rect 2625 35933 2641 35985
rect 2693 35976 3036 35985
rect 3070 35976 3076 36010
rect 2693 35946 3076 35976
rect 2693 35933 2891 35946
rect 1981 35921 2183 35933
rect 2217 35921 2419 35933
rect 2453 35921 2655 35933
rect 2689 35921 2891 35933
rect 1981 35912 2097 35921
rect 1225 35872 1241 35912
rect 1293 35872 2097 35912
rect 1225 35869 1239 35872
rect 1293 35869 1475 35872
rect 565 35857 767 35869
rect 801 35857 1003 35869
rect 1037 35857 1239 35869
rect 1273 35857 1475 35869
rect 565 35838 697 35857
rect 420 35813 697 35838
rect 380 35805 697 35813
rect 749 35805 765 35857
rect 817 35805 833 35857
rect 885 35805 901 35857
rect 953 35805 969 35857
rect 1021 35805 1037 35838
rect 1089 35805 1105 35857
rect 1157 35805 1173 35857
rect 1225 35838 1239 35857
rect 1293 35838 1475 35857
rect 1509 35838 1711 35872
rect 1745 35838 1947 35872
rect 1981 35869 2097 35872
rect 2149 35869 2165 35921
rect 2217 35869 2233 35921
rect 2285 35869 2301 35921
rect 2353 35869 2369 35921
rect 2421 35872 2437 35912
rect 2489 35869 2505 35921
rect 2557 35869 2573 35921
rect 2625 35869 2641 35921
rect 2693 35912 2891 35921
rect 2925 35938 3076 35946
rect 2925 35912 3036 35938
rect 2693 35904 3036 35912
rect 3070 35904 3076 35938
rect 2693 35872 3076 35904
rect 2693 35869 2891 35872
rect 1981 35857 2183 35869
rect 2217 35857 2419 35869
rect 2453 35857 2655 35869
rect 2689 35857 2891 35869
rect 1981 35838 2097 35857
rect 1225 35805 1241 35838
rect 1293 35805 2097 35838
rect 2149 35805 2165 35857
rect 2217 35805 2233 35857
rect 2285 35805 2301 35857
rect 2353 35805 2369 35857
rect 2421 35805 2437 35838
rect 2489 35805 2505 35857
rect 2557 35805 2573 35857
rect 2625 35805 2641 35857
rect 2693 35838 2891 35857
rect 2925 35866 3076 35872
rect 2925 35838 3036 35866
rect 2693 35832 3036 35838
rect 3070 35832 3076 35866
rect 2693 35805 3076 35832
rect 380 35798 3076 35805
rect 380 35775 531 35798
rect 380 35741 386 35775
rect 420 35764 531 35775
rect 565 35793 767 35798
rect 801 35793 1003 35798
rect 1037 35793 1239 35798
rect 1273 35793 1475 35798
rect 565 35764 697 35793
rect 420 35741 697 35764
rect 749 35741 765 35793
rect 817 35741 833 35793
rect 885 35741 901 35793
rect 953 35741 969 35793
rect 1021 35741 1037 35764
rect 1089 35741 1105 35793
rect 1157 35741 1173 35793
rect 1225 35764 1239 35793
rect 1293 35764 1475 35793
rect 1509 35764 1711 35798
rect 1745 35764 1947 35798
rect 1981 35793 2183 35798
rect 2217 35793 2419 35798
rect 2453 35793 2655 35798
rect 2689 35793 2891 35798
rect 1981 35764 2097 35793
rect 1225 35741 1241 35764
rect 1293 35741 2097 35764
rect 2149 35741 2165 35793
rect 2217 35741 2233 35793
rect 2285 35741 2301 35793
rect 2353 35741 2369 35793
rect 2421 35741 2437 35764
rect 2489 35741 2505 35793
rect 2557 35741 2573 35793
rect 2625 35741 2641 35793
rect 2693 35764 2891 35793
rect 2925 35794 3076 35798
rect 2925 35764 3036 35794
rect 2693 35760 3036 35764
rect 3070 35760 3076 35794
rect 2693 35741 3076 35760
rect 380 35729 3076 35741
rect 380 35724 697 35729
rect 380 35703 531 35724
rect 380 35669 386 35703
rect 420 35690 531 35703
rect 565 35690 697 35724
rect 420 35677 697 35690
rect 749 35677 765 35729
rect 817 35677 833 35729
rect 885 35677 901 35729
rect 953 35677 969 35729
rect 1021 35724 1037 35729
rect 1021 35677 1037 35690
rect 1089 35677 1105 35729
rect 1157 35677 1173 35729
rect 1225 35724 1241 35729
rect 1293 35724 2097 35729
rect 1225 35690 1239 35724
rect 1293 35690 1475 35724
rect 1509 35690 1711 35724
rect 1745 35690 1947 35724
rect 1981 35690 2097 35724
rect 1225 35677 1241 35690
rect 1293 35677 2097 35690
rect 2149 35677 2165 35729
rect 2217 35677 2233 35729
rect 2285 35677 2301 35729
rect 2353 35677 2369 35729
rect 2421 35724 2437 35729
rect 2421 35677 2437 35690
rect 2489 35677 2505 35729
rect 2557 35677 2573 35729
rect 2625 35677 2641 35729
rect 2693 35724 3076 35729
rect 2693 35690 2891 35724
rect 2925 35722 3076 35724
rect 2925 35690 3036 35722
rect 2693 35688 3036 35690
rect 3070 35688 3076 35722
rect 2693 35677 3076 35688
rect 420 35669 3076 35677
rect 380 35665 3076 35669
rect 380 35650 697 35665
rect 380 35631 531 35650
rect 380 35597 386 35631
rect 420 35616 531 35631
rect 565 35616 697 35650
rect 420 35613 697 35616
rect 749 35613 765 35665
rect 817 35613 833 35665
rect 885 35613 901 35665
rect 953 35613 969 35665
rect 1021 35650 1037 35665
rect 1021 35613 1037 35616
rect 1089 35613 1105 35665
rect 1157 35613 1173 35665
rect 1225 35650 1241 35665
rect 1293 35650 2097 35665
rect 1225 35616 1239 35650
rect 1293 35616 1475 35650
rect 1509 35616 1711 35650
rect 1745 35616 1947 35650
rect 1981 35616 2097 35650
rect 1225 35613 1241 35616
rect 1293 35613 2097 35616
rect 2149 35613 2165 35665
rect 2217 35613 2233 35665
rect 2285 35613 2301 35665
rect 2353 35613 2369 35665
rect 2421 35650 2437 35665
rect 2421 35613 2437 35616
rect 2489 35613 2505 35665
rect 2557 35613 2573 35665
rect 2625 35613 2641 35665
rect 2693 35650 3076 35665
rect 2693 35616 2891 35650
rect 2925 35616 3036 35650
rect 3070 35616 3076 35650
rect 2693 35613 3076 35616
rect 420 35601 3076 35613
rect 420 35597 697 35601
rect 380 35576 697 35597
rect 380 35559 531 35576
rect 380 35525 386 35559
rect 420 35542 531 35559
rect 565 35549 697 35576
rect 749 35549 765 35601
rect 817 35549 833 35601
rect 885 35549 901 35601
rect 953 35549 969 35601
rect 1021 35576 1037 35601
rect 1089 35549 1105 35601
rect 1157 35549 1173 35601
rect 1225 35576 1241 35601
rect 1293 35576 2097 35601
rect 1225 35549 1239 35576
rect 1293 35549 1475 35576
rect 565 35542 767 35549
rect 801 35542 1003 35549
rect 1037 35542 1239 35549
rect 1273 35542 1475 35549
rect 1509 35542 1711 35576
rect 1745 35542 1947 35576
rect 1981 35549 2097 35576
rect 2149 35549 2165 35601
rect 2217 35549 2233 35601
rect 2285 35549 2301 35601
rect 2353 35549 2369 35601
rect 2421 35576 2437 35601
rect 2489 35549 2505 35601
rect 2557 35549 2573 35601
rect 2625 35549 2641 35601
rect 2693 35578 3076 35601
rect 2693 35576 3036 35578
rect 2693 35549 2891 35576
rect 1981 35542 2183 35549
rect 2217 35542 2419 35549
rect 2453 35542 2655 35549
rect 2689 35542 2891 35549
rect 2925 35544 3036 35576
rect 3070 35544 3076 35578
rect 2925 35542 3076 35544
rect 420 35537 3076 35542
rect 420 35525 697 35537
rect 380 35502 697 35525
rect 380 35487 531 35502
rect 380 35453 386 35487
rect 420 35468 531 35487
rect 565 35485 697 35502
rect 749 35485 765 35537
rect 817 35485 833 35537
rect 885 35485 901 35537
rect 953 35485 969 35537
rect 1021 35502 1037 35537
rect 1089 35485 1105 35537
rect 1157 35485 1173 35537
rect 1225 35502 1241 35537
rect 1293 35502 2097 35537
rect 1225 35485 1239 35502
rect 1293 35485 1475 35502
rect 565 35473 767 35485
rect 801 35473 1003 35485
rect 1037 35473 1239 35485
rect 1273 35473 1475 35485
rect 565 35468 697 35473
rect 420 35453 697 35468
rect 380 35428 697 35453
rect 380 35415 531 35428
rect 380 35381 386 35415
rect 420 35394 531 35415
rect 565 35421 697 35428
rect 749 35421 765 35473
rect 817 35421 833 35473
rect 885 35421 901 35473
rect 953 35421 969 35473
rect 1021 35428 1037 35468
rect 1089 35421 1105 35473
rect 1157 35421 1173 35473
rect 1225 35468 1239 35473
rect 1293 35468 1475 35473
rect 1509 35468 1711 35502
rect 1745 35468 1947 35502
rect 1981 35485 2097 35502
rect 2149 35485 2165 35537
rect 2217 35485 2233 35537
rect 2285 35485 2301 35537
rect 2353 35485 2369 35537
rect 2421 35502 2437 35537
rect 2489 35485 2505 35537
rect 2557 35485 2573 35537
rect 2625 35485 2641 35537
rect 2693 35506 3076 35537
rect 2693 35502 3036 35506
rect 2693 35485 2891 35502
rect 1981 35473 2183 35485
rect 2217 35473 2419 35485
rect 2453 35473 2655 35485
rect 2689 35473 2891 35485
rect 1981 35468 2097 35473
rect 1225 35428 1241 35468
rect 1293 35428 2097 35468
rect 1225 35421 1239 35428
rect 1293 35421 1475 35428
rect 565 35394 767 35421
rect 801 35394 1003 35421
rect 1037 35394 1239 35421
rect 1273 35394 1475 35421
rect 1509 35394 1711 35428
rect 1745 35394 1947 35428
rect 1981 35421 2097 35428
rect 2149 35421 2165 35473
rect 2217 35421 2233 35473
rect 2285 35421 2301 35473
rect 2353 35421 2369 35473
rect 2421 35428 2437 35468
rect 2489 35421 2505 35473
rect 2557 35421 2573 35473
rect 2625 35421 2641 35473
rect 2693 35468 2891 35473
rect 2925 35472 3036 35502
rect 3070 35472 3076 35506
rect 2925 35468 3076 35472
rect 2693 35434 3076 35468
rect 2693 35428 3036 35434
rect 2693 35421 2891 35428
rect 1981 35394 2183 35421
rect 2217 35394 2419 35421
rect 2453 35394 2655 35421
rect 2689 35394 2891 35421
rect 2925 35400 3036 35428
rect 3070 35400 3076 35434
rect 2925 35394 3076 35400
rect 420 35393 3076 35394
rect 420 35381 588 35393
rect 380 35376 588 35381
tri 588 35376 605 35393 nw
tri 727 35376 744 35393 ne
rect 744 35376 824 35393
tri 824 35376 841 35393 nw
tri 963 35376 980 35393 ne
rect 980 35376 1060 35393
tri 1060 35376 1077 35393 nw
tri 1199 35376 1216 35393 ne
rect 1216 35376 1296 35393
tri 1296 35376 1313 35393 nw
tri 1435 35376 1452 35393 ne
rect 1452 35376 1532 35393
tri 1532 35376 1549 35393 nw
tri 1671 35376 1688 35393 ne
rect 1688 35376 1768 35393
tri 1768 35376 1785 35393 nw
tri 1907 35376 1924 35393 ne
rect 1924 35376 2004 35393
tri 2004 35376 2021 35393 nw
tri 2143 35376 2160 35393 ne
rect 2160 35376 2240 35393
tri 2240 35376 2257 35393 nw
tri 2379 35376 2396 35393 ne
rect 2396 35376 2476 35393
tri 2476 35376 2493 35393 nw
tri 2615 35376 2632 35393 ne
rect 2632 35376 2712 35393
tri 2712 35376 2729 35393 nw
tri 2851 35376 2868 35393 ne
rect 2868 35376 3076 35393
rect 380 35362 574 35376
tri 574 35362 588 35376 nw
tri 744 35362 758 35376 ne
rect 758 35362 810 35376
tri 810 35362 824 35376 nw
tri 980 35362 994 35376 ne
rect 994 35362 1046 35376
tri 1046 35362 1060 35376 nw
tri 1216 35362 1230 35376 ne
rect 1230 35362 1282 35376
tri 1282 35362 1296 35376 nw
tri 1452 35362 1466 35376 ne
rect 1466 35362 1518 35376
tri 1518 35362 1532 35376 nw
tri 1688 35362 1702 35376 ne
rect 1702 35362 1754 35376
tri 1754 35362 1768 35376 nw
tri 1924 35362 1938 35376 ne
rect 1938 35362 1990 35376
tri 1990 35362 2004 35376 nw
tri 2160 35362 2174 35376 ne
rect 2174 35362 2226 35376
tri 2226 35362 2240 35376 nw
tri 2396 35362 2410 35376 ne
rect 2410 35362 2462 35376
tri 2462 35362 2476 35376 nw
tri 2632 35362 2646 35376 ne
rect 2646 35362 2698 35376
tri 2698 35362 2712 35376 nw
tri 2868 35362 2882 35376 ne
rect 2882 35362 3076 35376
rect 380 35354 571 35362
tri 571 35359 574 35362 nw
tri 758 35359 761 35362 ne
rect 380 35343 531 35354
rect 380 35309 386 35343
rect 420 35320 531 35343
rect 565 35320 571 35354
rect 420 35309 571 35320
rect 380 35280 571 35309
rect 380 35271 531 35280
rect 380 35237 386 35271
rect 420 35246 531 35271
rect 565 35246 571 35280
rect 420 35237 571 35246
rect 380 35206 571 35237
rect 380 35199 531 35206
rect 380 35165 386 35199
rect 420 35172 531 35199
rect 565 35172 571 35206
rect 420 35165 571 35172
rect 380 35132 571 35165
rect 380 35127 531 35132
rect 380 35093 386 35127
rect 420 35098 531 35127
rect 565 35098 571 35132
rect 420 35093 571 35098
rect 380 35058 571 35093
rect 380 35055 531 35058
rect 380 35021 386 35055
rect 420 35024 531 35055
rect 565 35024 571 35058
rect 420 35021 571 35024
rect 380 34984 571 35021
rect 380 34983 531 34984
rect 380 34949 386 34983
rect 420 34950 531 34983
rect 565 34950 571 34984
rect 420 34949 571 34950
rect 380 34911 571 34949
rect 380 34877 386 34911
rect 420 34910 571 34911
rect 420 34877 531 34910
rect 380 34876 531 34877
rect 565 34876 571 34910
rect 380 34839 571 34876
rect 761 35354 807 35362
tri 807 35359 810 35362 nw
tri 994 35359 997 35362 ne
rect 761 35320 767 35354
rect 801 35320 807 35354
rect 761 35280 807 35320
rect 761 35246 767 35280
rect 801 35246 807 35280
rect 761 35206 807 35246
rect 761 35172 767 35206
rect 801 35172 807 35206
rect 761 35132 807 35172
rect 761 35098 767 35132
rect 801 35098 807 35132
rect 761 35058 807 35098
rect 761 35024 767 35058
rect 801 35024 807 35058
rect 761 34984 807 35024
rect 761 34950 767 34984
rect 801 34950 807 34984
rect 761 34910 807 34950
rect 761 34876 767 34910
rect 801 34876 807 34910
rect 761 34864 807 34876
rect 997 35354 1043 35362
tri 1043 35359 1046 35362 nw
tri 1230 35359 1233 35362 ne
rect 997 35320 1003 35354
rect 1037 35320 1043 35354
rect 997 35280 1043 35320
rect 997 35246 1003 35280
rect 1037 35246 1043 35280
rect 997 35206 1043 35246
rect 997 35172 1003 35206
rect 1037 35172 1043 35206
rect 997 35132 1043 35172
rect 997 35098 1003 35132
rect 1037 35098 1043 35132
rect 997 35058 1043 35098
rect 997 35024 1003 35058
rect 1037 35024 1043 35058
rect 997 34984 1043 35024
rect 997 34950 1003 34984
rect 1037 34950 1043 34984
rect 997 34910 1043 34950
rect 997 34876 1003 34910
rect 1037 34876 1043 34910
rect 997 34864 1043 34876
rect 1233 35354 1279 35362
tri 1279 35359 1282 35362 nw
tri 1466 35359 1469 35362 ne
rect 1233 35320 1239 35354
rect 1273 35320 1279 35354
rect 1233 35280 1279 35320
rect 1233 35246 1239 35280
rect 1273 35246 1279 35280
rect 1233 35206 1279 35246
rect 1233 35172 1239 35206
rect 1273 35172 1279 35206
rect 1233 35132 1279 35172
rect 1233 35098 1239 35132
rect 1273 35098 1279 35132
rect 1233 35058 1279 35098
rect 1233 35024 1239 35058
rect 1273 35024 1279 35058
rect 1233 34984 1279 35024
rect 1233 34950 1239 34984
rect 1273 34950 1279 34984
rect 1233 34910 1279 34950
rect 1233 34876 1239 34910
rect 1273 34876 1279 34910
rect 1233 34864 1279 34876
rect 1469 35354 1515 35362
tri 1515 35359 1518 35362 nw
tri 1702 35359 1705 35362 ne
rect 1469 35320 1475 35354
rect 1509 35320 1515 35354
rect 1469 35280 1515 35320
rect 1469 35246 1475 35280
rect 1509 35246 1515 35280
rect 1469 35206 1515 35246
rect 1469 35172 1475 35206
rect 1509 35172 1515 35206
rect 1469 35132 1515 35172
rect 1469 35098 1475 35132
rect 1509 35098 1515 35132
rect 1469 35058 1515 35098
rect 1469 35024 1475 35058
rect 1509 35024 1515 35058
rect 1469 34984 1515 35024
rect 1469 34950 1475 34984
rect 1509 34950 1515 34984
rect 1469 34910 1515 34950
rect 1469 34876 1475 34910
rect 1509 34876 1515 34910
rect 1469 34864 1515 34876
rect 1705 35354 1751 35362
tri 1751 35359 1754 35362 nw
tri 1938 35359 1941 35362 ne
rect 1705 35320 1711 35354
rect 1745 35320 1751 35354
rect 1705 35280 1751 35320
rect 1705 35246 1711 35280
rect 1745 35246 1751 35280
rect 1705 35206 1751 35246
rect 1705 35172 1711 35206
rect 1745 35172 1751 35206
rect 1705 35132 1751 35172
rect 1705 35098 1711 35132
rect 1745 35098 1751 35132
rect 1705 35058 1751 35098
rect 1705 35024 1711 35058
rect 1745 35024 1751 35058
rect 1705 34984 1751 35024
rect 1705 34950 1711 34984
rect 1745 34950 1751 34984
rect 1705 34910 1751 34950
rect 1705 34876 1711 34910
rect 1745 34876 1751 34910
rect 1705 34864 1751 34876
rect 1941 35354 1987 35362
tri 1987 35359 1990 35362 nw
tri 2174 35359 2177 35362 ne
rect 1941 35320 1947 35354
rect 1981 35320 1987 35354
rect 1941 35280 1987 35320
rect 1941 35246 1947 35280
rect 1981 35246 1987 35280
rect 1941 35206 1987 35246
rect 1941 35172 1947 35206
rect 1981 35172 1987 35206
rect 1941 35132 1987 35172
rect 1941 35098 1947 35132
rect 1981 35098 1987 35132
rect 1941 35058 1987 35098
rect 1941 35024 1947 35058
rect 1981 35024 1987 35058
rect 1941 34984 1987 35024
rect 1941 34950 1947 34984
rect 1981 34950 1987 34984
rect 1941 34910 1987 34950
rect 1941 34876 1947 34910
rect 1981 34876 1987 34910
rect 1941 34864 1987 34876
rect 2177 35354 2223 35362
tri 2223 35359 2226 35362 nw
tri 2410 35359 2413 35362 ne
rect 2177 35320 2183 35354
rect 2217 35320 2223 35354
rect 2177 35280 2223 35320
rect 2177 35246 2183 35280
rect 2217 35246 2223 35280
rect 2177 35206 2223 35246
rect 2177 35172 2183 35206
rect 2217 35172 2223 35206
rect 2177 35132 2223 35172
rect 2177 35098 2183 35132
rect 2217 35098 2223 35132
rect 2177 35058 2223 35098
rect 2177 35024 2183 35058
rect 2217 35024 2223 35058
rect 2177 34984 2223 35024
rect 2177 34950 2183 34984
rect 2217 34950 2223 34984
rect 2177 34910 2223 34950
rect 2177 34876 2183 34910
rect 2217 34876 2223 34910
rect 2177 34864 2223 34876
rect 2413 35354 2459 35362
tri 2459 35359 2462 35362 nw
tri 2646 35359 2649 35362 ne
rect 2413 35320 2419 35354
rect 2453 35320 2459 35354
rect 2413 35280 2459 35320
rect 2413 35246 2419 35280
rect 2453 35246 2459 35280
rect 2413 35206 2459 35246
rect 2413 35172 2419 35206
rect 2453 35172 2459 35206
rect 2413 35132 2459 35172
rect 2413 35098 2419 35132
rect 2453 35098 2459 35132
rect 2413 35058 2459 35098
rect 2413 35024 2419 35058
rect 2453 35024 2459 35058
rect 2413 34984 2459 35024
rect 2413 34950 2419 34984
rect 2453 34950 2459 34984
rect 2413 34910 2459 34950
rect 2413 34876 2419 34910
rect 2453 34876 2459 34910
rect 2413 34864 2459 34876
rect 2649 35354 2695 35362
tri 2695 35359 2698 35362 nw
tri 2882 35359 2885 35362 ne
rect 2649 35320 2655 35354
rect 2689 35320 2695 35354
rect 2649 35280 2695 35320
rect 2649 35246 2655 35280
rect 2689 35246 2695 35280
rect 2649 35206 2695 35246
rect 2649 35172 2655 35206
rect 2689 35172 2695 35206
rect 2649 35132 2695 35172
rect 2649 35098 2655 35132
rect 2689 35098 2695 35132
rect 2649 35058 2695 35098
rect 2649 35024 2655 35058
rect 2689 35024 2695 35058
rect 2649 34984 2695 35024
rect 2649 34950 2655 34984
rect 2689 34950 2695 34984
rect 2649 34910 2695 34950
rect 2649 34876 2655 34910
rect 2689 34876 2695 34910
rect 2649 34864 2695 34876
rect 2885 35354 3036 35362
rect 2885 35320 2891 35354
rect 2925 35328 3036 35354
rect 3070 35328 3076 35362
rect 2925 35320 3076 35328
rect 2885 35290 3076 35320
rect 2885 35280 3036 35290
rect 2885 35246 2891 35280
rect 2925 35256 3036 35280
rect 3070 35256 3076 35290
rect 2925 35246 3076 35256
rect 2885 35218 3076 35246
rect 2885 35206 3036 35218
rect 2885 35172 2891 35206
rect 2925 35184 3036 35206
rect 3070 35184 3076 35218
rect 2925 35172 3076 35184
rect 2885 35146 3076 35172
rect 2885 35132 3036 35146
rect 2885 35098 2891 35132
rect 2925 35112 3036 35132
rect 3070 35112 3076 35146
rect 2925 35098 3076 35112
rect 2885 35074 3076 35098
rect 2885 35058 3036 35074
rect 2885 35024 2891 35058
rect 2925 35040 3036 35058
rect 3070 35040 3076 35074
rect 2925 35024 3076 35040
rect 2885 35002 3076 35024
rect 2885 34984 3036 35002
rect 2885 34950 2891 34984
rect 2925 34968 3036 34984
rect 3070 34968 3076 35002
rect 2925 34950 3076 34968
rect 2885 34930 3076 34950
rect 2885 34910 3036 34930
rect 2885 34876 2891 34910
rect 2925 34896 3036 34910
rect 3070 34896 3076 34930
rect 2925 34876 3076 34896
rect 380 34805 386 34839
rect 420 34805 571 34839
rect 380 34767 571 34805
rect 2885 34858 3076 34876
rect 2885 34824 3036 34858
rect 3070 34824 3076 34858
rect 380 34733 386 34767
rect 420 34733 571 34767
rect 613 34794 1501 34803
rect 1553 34794 1569 34803
rect 1621 34794 1636 34803
rect 1688 34794 1703 34803
rect 1755 34794 1770 34803
rect 1822 34794 1837 34803
rect 1889 34794 2830 34803
rect 613 34760 625 34794
rect 659 34760 700 34794
rect 734 34760 775 34794
rect 809 34760 850 34794
rect 884 34760 925 34794
rect 959 34760 1000 34794
rect 1034 34760 1075 34794
rect 1109 34760 1150 34794
rect 1184 34760 1225 34794
rect 1259 34760 1300 34794
rect 1334 34760 1375 34794
rect 1409 34760 1450 34794
rect 1484 34760 1501 34794
rect 1559 34760 1569 34794
rect 1634 34760 1636 34794
rect 1889 34760 1896 34794
rect 1930 34760 1970 34794
rect 2004 34760 2044 34794
rect 2078 34760 2118 34794
rect 2152 34760 2192 34794
rect 2226 34760 2266 34794
rect 2300 34760 2340 34794
rect 2374 34760 2414 34794
rect 2448 34760 2488 34794
rect 2522 34760 2562 34794
rect 2596 34760 2636 34794
rect 2670 34760 2710 34794
rect 2744 34760 2784 34794
rect 2818 34760 2830 34794
rect 613 34751 1501 34760
rect 1553 34751 1569 34760
rect 1621 34751 1636 34760
rect 1688 34751 1703 34760
rect 1755 34751 1770 34760
rect 1822 34751 1837 34760
rect 1889 34751 2830 34760
rect 2885 34786 3076 34824
rect 2885 34752 3036 34786
rect 3070 34752 3076 34786
rect 380 34695 571 34733
rect 2885 34714 3076 34752
rect 380 34661 386 34695
rect 420 34692 571 34695
rect 420 34661 531 34692
rect 380 34658 531 34661
rect 565 34658 571 34692
rect 380 34623 571 34658
rect 380 34589 386 34623
rect 420 34619 571 34623
rect 420 34589 531 34619
rect 380 34585 531 34589
rect 565 34585 571 34619
rect 380 34551 571 34585
rect 380 34517 386 34551
rect 420 34546 571 34551
rect 420 34517 531 34546
rect 380 34512 531 34517
rect 565 34512 571 34546
rect 380 34479 571 34512
rect 380 34445 386 34479
rect 420 34473 571 34479
rect 420 34445 531 34473
rect 380 34439 531 34445
rect 565 34439 571 34473
rect 380 34407 571 34439
rect 380 34373 386 34407
rect 420 34400 571 34407
rect 420 34373 531 34400
rect 380 34366 531 34373
rect 565 34366 571 34400
rect 380 34335 571 34366
rect 380 34301 386 34335
rect 420 34327 571 34335
rect 420 34301 531 34327
rect 380 34293 531 34301
rect 565 34293 571 34327
rect 380 34263 571 34293
rect 380 34229 386 34263
rect 420 34254 571 34263
rect 420 34229 531 34254
rect 380 34220 531 34229
rect 565 34220 571 34254
rect 380 34191 571 34220
rect 761 34692 807 34704
rect 761 34658 767 34692
rect 801 34658 807 34692
rect 761 34619 807 34658
rect 761 34585 767 34619
rect 801 34585 807 34619
rect 761 34546 807 34585
rect 761 34512 767 34546
rect 801 34512 807 34546
rect 761 34473 807 34512
rect 761 34439 767 34473
rect 801 34439 807 34473
rect 761 34400 807 34439
rect 761 34366 767 34400
rect 801 34366 807 34400
rect 761 34327 807 34366
rect 761 34293 767 34327
rect 801 34293 807 34327
rect 761 34254 807 34293
rect 761 34220 767 34254
rect 801 34220 807 34254
rect 380 34157 386 34191
rect 420 34181 571 34191
tri 571 34181 600 34210 sw
tri 732 34181 761 34210 se
rect 761 34181 807 34220
rect 997 34692 1043 34704
rect 997 34658 1003 34692
rect 1037 34658 1043 34692
rect 997 34619 1043 34658
rect 997 34585 1003 34619
rect 1037 34585 1043 34619
rect 997 34546 1043 34585
rect 997 34512 1003 34546
rect 1037 34512 1043 34546
rect 997 34473 1043 34512
rect 997 34439 1003 34473
rect 1037 34439 1043 34473
rect 997 34400 1043 34439
rect 997 34366 1003 34400
rect 1037 34366 1043 34400
rect 997 34327 1043 34366
rect 997 34293 1003 34327
rect 1037 34293 1043 34327
rect 997 34254 1043 34293
rect 997 34220 1003 34254
rect 1037 34220 1043 34254
tri 807 34181 836 34210 sw
tri 968 34181 997 34210 se
rect 997 34181 1043 34220
rect 1233 34692 1279 34704
rect 1233 34658 1239 34692
rect 1273 34658 1279 34692
rect 1233 34619 1279 34658
rect 1233 34585 1239 34619
rect 1273 34585 1279 34619
rect 1233 34546 1279 34585
rect 1233 34512 1239 34546
rect 1273 34512 1279 34546
rect 1233 34473 1279 34512
rect 1233 34439 1239 34473
rect 1273 34439 1279 34473
rect 1233 34400 1279 34439
rect 1233 34366 1239 34400
rect 1273 34366 1279 34400
rect 1233 34327 1279 34366
rect 1233 34293 1239 34327
rect 1273 34293 1279 34327
rect 1233 34254 1279 34293
rect 1233 34220 1239 34254
rect 1273 34220 1279 34254
tri 1043 34181 1072 34210 sw
tri 1204 34181 1233 34210 se
rect 1233 34181 1279 34220
rect 1469 34692 1515 34704
rect 1469 34658 1475 34692
rect 1509 34658 1515 34692
rect 1469 34619 1515 34658
rect 1469 34585 1475 34619
rect 1509 34585 1515 34619
rect 1469 34546 1515 34585
rect 1469 34512 1475 34546
rect 1509 34512 1515 34546
rect 1469 34473 1515 34512
rect 1469 34439 1475 34473
rect 1509 34439 1515 34473
rect 1469 34400 1515 34439
rect 1469 34366 1475 34400
rect 1509 34366 1515 34400
rect 1469 34327 1515 34366
rect 1469 34293 1475 34327
rect 1509 34293 1515 34327
rect 1469 34254 1515 34293
rect 1469 34220 1475 34254
rect 1509 34220 1515 34254
tri 1279 34181 1308 34210 sw
tri 1440 34181 1469 34210 se
rect 1469 34181 1515 34220
rect 1705 34692 1751 34704
rect 1705 34658 1711 34692
rect 1745 34658 1751 34692
rect 1705 34619 1751 34658
rect 1705 34585 1711 34619
rect 1745 34585 1751 34619
rect 1705 34546 1751 34585
rect 1705 34512 1711 34546
rect 1745 34512 1751 34546
rect 1705 34473 1751 34512
rect 1705 34439 1711 34473
rect 1745 34439 1751 34473
rect 1705 34400 1751 34439
rect 1705 34366 1711 34400
rect 1745 34366 1751 34400
rect 1705 34327 1751 34366
rect 1705 34293 1711 34327
rect 1745 34293 1751 34327
rect 1705 34254 1751 34293
rect 1705 34220 1711 34254
rect 1745 34220 1751 34254
tri 1515 34181 1544 34210 sw
tri 1676 34181 1705 34210 se
rect 1705 34181 1751 34220
rect 1941 34692 1987 34704
rect 1941 34658 1947 34692
rect 1981 34658 1987 34692
rect 1941 34619 1987 34658
rect 1941 34585 1947 34619
rect 1981 34585 1987 34619
rect 1941 34546 1987 34585
rect 1941 34512 1947 34546
rect 1981 34512 1987 34546
rect 1941 34473 1987 34512
rect 1941 34439 1947 34473
rect 1981 34439 1987 34473
rect 1941 34400 1987 34439
rect 1941 34366 1947 34400
rect 1981 34366 1987 34400
rect 1941 34327 1987 34366
rect 1941 34293 1947 34327
rect 1981 34293 1987 34327
rect 1941 34254 1987 34293
rect 1941 34220 1947 34254
rect 1981 34220 1987 34254
tri 1751 34181 1780 34210 sw
tri 1912 34181 1941 34210 se
rect 1941 34181 1987 34220
rect 2177 34692 2223 34704
rect 2177 34658 2183 34692
rect 2217 34658 2223 34692
rect 2177 34619 2223 34658
rect 2177 34585 2183 34619
rect 2217 34585 2223 34619
rect 2177 34546 2223 34585
rect 2177 34512 2183 34546
rect 2217 34512 2223 34546
rect 2177 34473 2223 34512
rect 2177 34439 2183 34473
rect 2217 34439 2223 34473
rect 2177 34400 2223 34439
rect 2177 34366 2183 34400
rect 2217 34366 2223 34400
rect 2177 34327 2223 34366
rect 2177 34293 2183 34327
rect 2217 34293 2223 34327
rect 2177 34254 2223 34293
rect 2177 34220 2183 34254
rect 2217 34220 2223 34254
tri 1987 34181 2016 34210 sw
tri 2148 34181 2177 34210 se
rect 2177 34181 2223 34220
rect 2413 34692 2459 34704
rect 2413 34658 2419 34692
rect 2453 34658 2459 34692
rect 2413 34619 2459 34658
rect 2413 34585 2419 34619
rect 2453 34585 2459 34619
rect 2413 34546 2459 34585
rect 2413 34512 2419 34546
rect 2453 34512 2459 34546
rect 2413 34473 2459 34512
rect 2413 34439 2419 34473
rect 2453 34439 2459 34473
rect 2413 34400 2459 34439
rect 2413 34366 2419 34400
rect 2453 34366 2459 34400
rect 2413 34327 2459 34366
rect 2413 34293 2419 34327
rect 2453 34293 2459 34327
rect 2413 34254 2459 34293
rect 2413 34220 2419 34254
rect 2453 34220 2459 34254
tri 2223 34181 2252 34210 sw
tri 2384 34181 2413 34210 se
rect 2413 34181 2459 34220
rect 2649 34692 2695 34704
rect 2649 34658 2655 34692
rect 2689 34658 2695 34692
rect 2649 34619 2695 34658
rect 2649 34585 2655 34619
rect 2689 34585 2695 34619
rect 2649 34546 2695 34585
rect 2649 34512 2655 34546
rect 2689 34512 2695 34546
rect 2649 34473 2695 34512
rect 2649 34439 2655 34473
rect 2689 34439 2695 34473
rect 2649 34400 2695 34439
rect 2649 34366 2655 34400
rect 2689 34366 2695 34400
rect 2649 34327 2695 34366
rect 2649 34293 2655 34327
rect 2689 34293 2695 34327
rect 2649 34254 2695 34293
rect 2649 34220 2655 34254
rect 2689 34220 2695 34254
tri 2459 34181 2488 34210 sw
tri 2620 34181 2649 34210 se
rect 2649 34181 2695 34220
rect 2885 34692 3036 34714
rect 2885 34658 2891 34692
rect 2925 34680 3036 34692
rect 3070 34680 3076 34714
rect 2925 34658 3076 34680
rect 2885 34642 3076 34658
rect 2885 34619 3036 34642
rect 2885 34585 2891 34619
rect 2925 34608 3036 34619
rect 3070 34608 3076 34642
rect 2925 34585 3076 34608
rect 2885 34570 3076 34585
rect 2885 34546 3036 34570
rect 2885 34512 2891 34546
rect 2925 34536 3036 34546
rect 3070 34536 3076 34570
rect 2925 34512 3076 34536
rect 2885 34498 3076 34512
rect 2885 34473 3036 34498
rect 2885 34439 2891 34473
rect 2925 34464 3036 34473
rect 3070 34464 3076 34498
rect 2925 34439 3076 34464
rect 2885 34426 3076 34439
rect 2885 34400 3036 34426
rect 2885 34366 2891 34400
rect 2925 34392 3036 34400
rect 3070 34392 3076 34426
rect 2925 34366 3076 34392
rect 2885 34354 3076 34366
rect 2885 34327 3036 34354
rect 2885 34293 2891 34327
rect 2925 34320 3036 34327
rect 3070 34320 3076 34354
rect 2925 34293 3076 34320
rect 2885 34282 3076 34293
rect 2885 34254 3036 34282
rect 2885 34220 2891 34254
rect 2925 34248 3036 34254
rect 3070 34248 3076 34282
rect 2925 34220 3076 34248
rect 2885 34210 3076 34220
tri 2695 34181 2724 34210 sw
tri 2856 34181 2885 34210 se
rect 2885 34181 3036 34210
rect 420 34157 531 34181
rect 380 34147 531 34157
rect 565 34176 600 34181
tri 600 34176 605 34181 sw
tri 727 34176 732 34181 se
rect 732 34176 767 34181
rect 565 34150 767 34176
rect 801 34176 836 34181
tri 836 34176 841 34181 sw
tri 963 34176 968 34181 se
rect 968 34176 1003 34181
rect 801 34150 1003 34176
rect 1037 34176 1072 34181
tri 1072 34176 1077 34181 sw
tri 1199 34176 1204 34181 se
rect 1204 34176 1239 34181
rect 1037 34150 1239 34176
rect 1273 34176 1308 34181
tri 1308 34176 1313 34181 sw
tri 1435 34176 1440 34181 se
rect 1440 34176 1475 34181
rect 1273 34150 1475 34176
rect 565 34147 697 34150
rect 380 34119 697 34147
rect 380 34085 386 34119
rect 420 34108 697 34119
rect 420 34085 531 34108
rect 380 34074 531 34085
rect 565 34098 697 34108
rect 749 34098 765 34150
rect 817 34098 833 34150
rect 885 34098 901 34150
rect 953 34098 969 34150
rect 1021 34108 1037 34147
rect 1089 34098 1105 34150
rect 1157 34098 1173 34150
rect 1225 34147 1239 34150
rect 1293 34147 1475 34150
rect 1509 34176 1544 34181
tri 1544 34176 1549 34181 sw
tri 1671 34176 1676 34181 se
rect 1676 34176 1711 34181
rect 1509 34147 1711 34176
rect 1745 34176 1780 34181
tri 1780 34176 1785 34181 sw
tri 1907 34176 1912 34181 se
rect 1912 34176 1947 34181
rect 1745 34147 1947 34176
rect 1981 34176 2016 34181
tri 2016 34176 2021 34181 sw
tri 2143 34176 2148 34181 se
rect 2148 34176 2183 34181
rect 1981 34150 2183 34176
rect 2217 34176 2252 34181
tri 2252 34176 2257 34181 sw
tri 2379 34176 2384 34181 se
rect 2384 34176 2419 34181
rect 2217 34150 2419 34176
rect 2453 34176 2488 34181
tri 2488 34176 2493 34181 sw
tri 2615 34176 2620 34181 se
rect 2620 34176 2655 34181
rect 2453 34150 2655 34176
rect 2689 34176 2724 34181
tri 2724 34176 2729 34181 sw
tri 2851 34176 2856 34181 se
rect 2856 34176 2891 34181
rect 2689 34150 2891 34176
rect 1981 34147 2097 34150
rect 1225 34108 1241 34147
rect 1293 34108 2097 34147
rect 1225 34098 1239 34108
rect 1293 34098 1475 34108
rect 565 34086 767 34098
rect 801 34086 1003 34098
rect 1037 34086 1239 34098
rect 1273 34086 1475 34098
rect 565 34074 697 34086
rect 380 34047 697 34074
rect 380 34013 386 34047
rect 420 34035 697 34047
rect 420 34013 531 34035
rect 380 34001 531 34013
rect 565 34034 697 34035
rect 749 34034 765 34086
rect 817 34034 833 34086
rect 885 34034 901 34086
rect 953 34034 969 34086
rect 1021 34035 1037 34074
rect 1089 34034 1105 34086
rect 1157 34034 1173 34086
rect 1225 34074 1239 34086
rect 1293 34074 1475 34086
rect 1509 34074 1711 34108
rect 1745 34074 1947 34108
rect 1981 34098 2097 34108
rect 2149 34098 2165 34150
rect 2217 34098 2233 34150
rect 2285 34098 2301 34150
rect 2353 34098 2369 34150
rect 2421 34108 2437 34147
rect 2489 34098 2505 34150
rect 2557 34098 2573 34150
rect 2625 34098 2641 34150
rect 2693 34147 2891 34150
rect 2925 34176 3036 34181
rect 3070 34176 3076 34210
rect 2925 34147 3076 34176
rect 2693 34138 3076 34147
rect 2693 34108 3036 34138
rect 2693 34098 2891 34108
rect 1981 34086 2183 34098
rect 2217 34086 2419 34098
rect 2453 34086 2655 34098
rect 2689 34086 2891 34098
rect 1981 34074 2097 34086
rect 1225 34035 1241 34074
rect 1293 34035 2097 34074
rect 1225 34034 1239 34035
rect 1293 34034 1475 34035
rect 565 34022 767 34034
rect 801 34022 1003 34034
rect 1037 34022 1239 34034
rect 1273 34022 1475 34034
rect 565 34001 697 34022
rect 380 33975 697 34001
rect 380 33941 386 33975
rect 420 33970 697 33975
rect 749 33970 765 34022
rect 817 33970 833 34022
rect 885 33970 901 34022
rect 953 33970 969 34022
rect 1021 33970 1037 34001
rect 1089 33970 1105 34022
rect 1157 33970 1173 34022
rect 1225 34001 1239 34022
rect 1293 34001 1475 34022
rect 1509 34001 1711 34035
rect 1745 34001 1947 34035
rect 1981 34034 2097 34035
rect 2149 34034 2165 34086
rect 2217 34034 2233 34086
rect 2285 34034 2301 34086
rect 2353 34034 2369 34086
rect 2421 34035 2437 34074
rect 2489 34034 2505 34086
rect 2557 34034 2573 34086
rect 2625 34034 2641 34086
rect 2693 34074 2891 34086
rect 2925 34104 3036 34108
rect 3070 34104 3076 34138
rect 2925 34074 3076 34104
rect 2693 34066 3076 34074
rect 2693 34035 3036 34066
rect 2693 34034 2891 34035
rect 1981 34022 2183 34034
rect 2217 34022 2419 34034
rect 2453 34022 2655 34034
rect 2689 34022 2891 34034
rect 1981 34001 2097 34022
rect 1225 33970 1241 34001
rect 1293 33970 2097 34001
rect 2149 33970 2165 34022
rect 2217 33970 2233 34022
rect 2285 33970 2301 34022
rect 2353 33970 2369 34022
rect 2421 33970 2437 34001
rect 2489 33970 2505 34022
rect 2557 33970 2573 34022
rect 2625 33970 2641 34022
rect 2693 34001 2891 34022
rect 2925 34032 3036 34035
rect 3070 34032 3076 34066
rect 2925 34001 3076 34032
rect 2693 33994 3076 34001
rect 2693 33970 3036 33994
rect 420 33962 3036 33970
rect 420 33941 531 33962
rect 380 33928 531 33941
rect 565 33958 767 33962
rect 801 33958 1003 33962
rect 1037 33958 1239 33962
rect 1273 33958 1475 33962
rect 565 33928 697 33958
rect 380 33906 697 33928
rect 749 33906 765 33958
rect 817 33906 833 33958
rect 885 33906 901 33958
rect 953 33906 969 33958
rect 1021 33906 1037 33928
rect 1089 33906 1105 33958
rect 1157 33906 1173 33958
rect 1225 33928 1239 33958
rect 1293 33928 1475 33958
rect 1509 33928 1711 33962
rect 1745 33928 1947 33962
rect 1981 33958 2183 33962
rect 2217 33958 2419 33962
rect 2453 33958 2655 33962
rect 2689 33958 2891 33962
rect 1981 33928 2097 33958
rect 1225 33906 1241 33928
rect 1293 33906 2097 33928
rect 2149 33906 2165 33958
rect 2217 33906 2233 33958
rect 2285 33906 2301 33958
rect 2353 33906 2369 33958
rect 2421 33906 2437 33928
rect 2489 33906 2505 33958
rect 2557 33906 2573 33958
rect 2625 33906 2641 33958
rect 2693 33928 2891 33958
rect 2925 33960 3036 33962
rect 3070 33960 3076 33994
rect 2925 33928 3076 33960
rect 2693 33922 3076 33928
rect 2693 33906 3036 33922
rect 380 33903 3036 33906
rect 380 33869 386 33903
rect 420 33894 3036 33903
rect 420 33889 697 33894
rect 420 33869 531 33889
rect 380 33855 531 33869
rect 565 33855 697 33889
rect 380 33842 697 33855
rect 749 33842 765 33894
rect 817 33842 833 33894
rect 885 33842 901 33894
rect 953 33842 969 33894
rect 1021 33889 1037 33894
rect 1021 33842 1037 33855
rect 1089 33842 1105 33894
rect 1157 33842 1173 33894
rect 1225 33889 1241 33894
rect 1293 33889 2097 33894
rect 1225 33855 1239 33889
rect 1293 33855 1475 33889
rect 1509 33855 1711 33889
rect 1745 33855 1947 33889
rect 1981 33855 2097 33889
rect 1225 33842 1241 33855
rect 1293 33842 2097 33855
rect 2149 33842 2165 33894
rect 2217 33842 2233 33894
rect 2285 33842 2301 33894
rect 2353 33842 2369 33894
rect 2421 33889 2437 33894
rect 2421 33842 2437 33855
rect 2489 33842 2505 33894
rect 2557 33842 2573 33894
rect 2625 33842 2641 33894
rect 2693 33889 3036 33894
rect 2693 33855 2891 33889
rect 2925 33888 3036 33889
rect 3070 33888 3076 33922
rect 2925 33855 3076 33888
rect 2693 33850 3076 33855
rect 2693 33842 3036 33850
rect 380 33831 3036 33842
rect 380 33797 386 33831
rect 420 33830 3036 33831
rect 420 33816 697 33830
rect 420 33797 531 33816
rect 380 33782 531 33797
rect 565 33782 697 33816
rect 380 33778 697 33782
rect 749 33778 765 33830
rect 817 33778 833 33830
rect 885 33778 901 33830
rect 953 33778 969 33830
rect 1021 33816 1037 33830
rect 1021 33778 1037 33782
rect 1089 33778 1105 33830
rect 1157 33778 1173 33830
rect 1225 33816 1241 33830
rect 1293 33816 2097 33830
rect 1225 33782 1239 33816
rect 1293 33782 1475 33816
rect 1509 33782 1711 33816
rect 1745 33782 1947 33816
rect 1981 33782 2097 33816
rect 1225 33778 1241 33782
rect 1293 33778 2097 33782
rect 2149 33778 2165 33830
rect 2217 33778 2233 33830
rect 2285 33778 2301 33830
rect 2353 33778 2369 33830
rect 2421 33816 2437 33830
rect 2421 33778 2437 33782
rect 2489 33778 2505 33830
rect 2557 33778 2573 33830
rect 2625 33778 2641 33830
rect 2693 33816 3036 33830
rect 3070 33816 3076 33850
rect 2693 33782 2891 33816
rect 2925 33782 3076 33816
rect 2693 33778 3076 33782
rect 380 33766 3036 33778
rect 380 33759 697 33766
rect 380 33725 386 33759
rect 420 33742 697 33759
rect 420 33725 531 33742
rect 380 33708 531 33725
rect 565 33714 697 33742
rect 749 33714 765 33766
rect 817 33714 833 33766
rect 885 33714 901 33766
rect 953 33714 969 33766
rect 1021 33742 1037 33766
rect 1089 33714 1105 33766
rect 1157 33714 1173 33766
rect 1225 33742 1241 33766
rect 1293 33742 2097 33766
rect 1225 33714 1239 33742
rect 1293 33714 1475 33742
rect 565 33708 767 33714
rect 801 33708 1003 33714
rect 1037 33708 1239 33714
rect 1273 33708 1475 33714
rect 1509 33708 1711 33742
rect 1745 33708 1947 33742
rect 1981 33714 2097 33742
rect 2149 33714 2165 33766
rect 2217 33714 2233 33766
rect 2285 33714 2301 33766
rect 2353 33714 2369 33766
rect 2421 33742 2437 33766
rect 2489 33714 2505 33766
rect 2557 33714 2573 33766
rect 2625 33714 2641 33766
rect 2693 33744 3036 33766
rect 3070 33744 3076 33778
rect 2693 33742 3076 33744
rect 2693 33714 2891 33742
rect 1981 33708 2183 33714
rect 2217 33708 2419 33714
rect 2453 33708 2655 33714
rect 2689 33708 2891 33714
rect 2925 33708 3076 33742
rect 380 33706 3076 33708
rect 380 33702 3036 33706
rect 380 33687 697 33702
rect 380 33653 386 33687
rect 420 33668 697 33687
rect 420 33653 531 33668
rect 380 33634 531 33653
rect 565 33650 697 33668
rect 749 33650 765 33702
rect 817 33650 833 33702
rect 885 33650 901 33702
rect 953 33650 969 33702
rect 1021 33668 1037 33702
rect 1089 33650 1105 33702
rect 1157 33650 1173 33702
rect 1225 33668 1241 33702
rect 1293 33668 2097 33702
rect 1225 33650 1239 33668
rect 1293 33650 1475 33668
rect 565 33638 767 33650
rect 801 33638 1003 33650
rect 1037 33638 1239 33650
rect 1273 33638 1475 33650
rect 565 33634 697 33638
rect 380 33615 697 33634
rect 380 33581 386 33615
rect 420 33594 697 33615
rect 420 33581 531 33594
rect 380 33560 531 33581
rect 565 33586 697 33594
rect 749 33586 765 33638
rect 817 33586 833 33638
rect 885 33586 901 33638
rect 953 33586 969 33638
rect 1021 33594 1037 33634
rect 1089 33586 1105 33638
rect 1157 33586 1173 33638
rect 1225 33634 1239 33638
rect 1293 33634 1475 33638
rect 1509 33634 1711 33668
rect 1745 33634 1947 33668
rect 1981 33650 2097 33668
rect 2149 33650 2165 33702
rect 2217 33650 2233 33702
rect 2285 33650 2301 33702
rect 2353 33650 2369 33702
rect 2421 33668 2437 33702
rect 2489 33650 2505 33702
rect 2557 33650 2573 33702
rect 2625 33650 2641 33702
rect 2693 33672 3036 33702
rect 3070 33672 3076 33706
rect 2693 33668 3076 33672
rect 2693 33650 2891 33668
rect 1981 33638 2183 33650
rect 2217 33638 2419 33650
rect 2453 33638 2655 33650
rect 2689 33638 2891 33650
rect 1981 33634 2097 33638
rect 1225 33594 1241 33634
rect 1293 33594 2097 33634
rect 1225 33586 1239 33594
rect 1293 33586 1475 33594
rect 565 33574 767 33586
rect 801 33574 1003 33586
rect 1037 33574 1239 33586
rect 1273 33574 1475 33586
rect 565 33560 697 33574
rect 380 33543 697 33560
rect 380 33509 386 33543
rect 420 33522 697 33543
rect 749 33522 765 33574
rect 817 33522 833 33574
rect 885 33522 901 33574
rect 953 33522 969 33574
rect 1021 33522 1037 33560
rect 1089 33522 1105 33574
rect 1157 33522 1173 33574
rect 1225 33560 1239 33574
rect 1293 33560 1475 33574
rect 1509 33560 1711 33594
rect 1745 33560 1947 33594
rect 1981 33586 2097 33594
rect 2149 33586 2165 33638
rect 2217 33586 2233 33638
rect 2285 33586 2301 33638
rect 2353 33586 2369 33638
rect 2421 33594 2437 33634
rect 2489 33586 2505 33638
rect 2557 33586 2573 33638
rect 2625 33586 2641 33638
rect 2693 33634 2891 33638
rect 2925 33634 3076 33668
rect 2693 33600 3036 33634
rect 3070 33600 3076 33634
rect 2693 33594 3076 33600
rect 2693 33586 2891 33594
rect 1981 33574 2183 33586
rect 2217 33574 2419 33586
rect 2453 33574 2655 33586
rect 2689 33574 2891 33586
rect 1981 33560 2097 33574
rect 1225 33522 1241 33560
rect 1293 33522 2097 33560
rect 2149 33522 2165 33574
rect 2217 33522 2233 33574
rect 2285 33522 2301 33574
rect 2353 33522 2369 33574
rect 2421 33522 2437 33560
rect 2489 33522 2505 33574
rect 2557 33522 2573 33574
rect 2625 33522 2641 33574
rect 2693 33560 2891 33574
rect 2925 33562 3076 33594
rect 2925 33560 3036 33562
rect 2693 33528 3036 33560
rect 3070 33528 3076 33562
rect 2693 33522 3076 33528
rect 420 33520 3076 33522
rect 420 33509 531 33520
rect 380 33486 531 33509
rect 565 33510 767 33520
rect 801 33510 1003 33520
rect 1037 33510 1239 33520
rect 1273 33510 1475 33520
rect 565 33486 697 33510
rect 380 33471 697 33486
rect 380 33437 386 33471
rect 420 33458 697 33471
rect 749 33458 765 33510
rect 817 33458 833 33510
rect 885 33458 901 33510
rect 953 33458 969 33510
rect 1021 33458 1037 33486
rect 1089 33458 1105 33510
rect 1157 33458 1173 33510
rect 1225 33486 1239 33510
rect 1293 33486 1475 33510
rect 1509 33486 1711 33520
rect 1745 33486 1947 33520
rect 1981 33510 2183 33520
rect 2217 33510 2419 33520
rect 2453 33510 2655 33520
rect 2689 33510 2891 33520
rect 1981 33486 2097 33510
rect 1225 33458 1241 33486
rect 1293 33458 2097 33486
rect 2149 33458 2165 33510
rect 2217 33458 2233 33510
rect 2285 33458 2301 33510
rect 2353 33458 2369 33510
rect 2421 33458 2437 33486
rect 2489 33458 2505 33510
rect 2557 33458 2573 33510
rect 2625 33458 2641 33510
rect 2693 33486 2891 33510
rect 2925 33490 3076 33520
rect 2925 33486 3036 33490
rect 2693 33458 3036 33486
rect 420 33456 3036 33458
rect 3070 33456 3076 33490
rect 420 33446 3076 33456
rect 420 33437 531 33446
rect 380 33412 531 33437
rect 565 33412 697 33446
rect 380 33399 697 33412
rect 380 33365 386 33399
rect 420 33394 697 33399
rect 749 33394 765 33446
rect 817 33394 833 33446
rect 885 33394 901 33446
rect 953 33394 969 33446
rect 1021 33394 1037 33412
rect 1089 33394 1105 33446
rect 1157 33394 1173 33446
rect 1225 33412 1239 33446
rect 1293 33412 1475 33446
rect 1509 33412 1711 33446
rect 1745 33412 1947 33446
rect 1981 33412 2097 33446
rect 1225 33394 1241 33412
rect 1293 33394 2097 33412
rect 2149 33394 2165 33446
rect 2217 33394 2233 33446
rect 2285 33394 2301 33446
rect 2353 33394 2369 33446
rect 2421 33394 2437 33412
rect 2489 33394 2505 33446
rect 2557 33394 2573 33446
rect 2625 33394 2641 33446
rect 2693 33412 2891 33446
rect 2925 33418 3076 33446
rect 2925 33412 3036 33418
rect 2693 33394 3036 33412
rect 420 33384 3036 33394
rect 3070 33384 3076 33418
rect 420 33382 3076 33384
rect 420 33372 697 33382
rect 420 33365 531 33372
rect 380 33338 531 33365
rect 565 33338 697 33372
rect 380 33330 697 33338
rect 749 33330 765 33382
rect 817 33330 833 33382
rect 885 33330 901 33382
rect 953 33330 969 33382
rect 1021 33372 1037 33382
rect 1021 33330 1037 33338
rect 1089 33330 1105 33382
rect 1157 33330 1173 33382
rect 1225 33372 1241 33382
rect 1293 33372 2097 33382
rect 1225 33338 1239 33372
rect 1293 33338 1475 33372
rect 1509 33338 1711 33372
rect 1745 33338 1947 33372
rect 1981 33338 2097 33372
rect 1225 33330 1241 33338
rect 1293 33330 2097 33338
rect 2149 33330 2165 33382
rect 2217 33330 2233 33382
rect 2285 33330 2301 33382
rect 2353 33330 2369 33382
rect 2421 33372 2437 33382
rect 2421 33330 2437 33338
rect 2489 33330 2505 33382
rect 2557 33330 2573 33382
rect 2625 33330 2641 33382
rect 2693 33372 3076 33382
rect 2693 33338 2891 33372
rect 2925 33346 3076 33372
rect 2925 33338 3036 33346
rect 2693 33330 3036 33338
rect 380 33327 3036 33330
rect 380 33293 386 33327
rect 420 33318 3036 33327
rect 420 33298 697 33318
rect 420 33293 531 33298
rect 380 33264 531 33293
rect 565 33266 697 33298
rect 749 33266 765 33318
rect 817 33266 833 33318
rect 885 33266 901 33318
rect 953 33266 969 33318
rect 1021 33298 1037 33318
rect 1089 33266 1105 33318
rect 1157 33266 1173 33318
rect 1225 33298 1241 33318
rect 1293 33298 2097 33318
rect 1225 33266 1239 33298
rect 1293 33266 1475 33298
rect 565 33264 767 33266
rect 801 33264 1003 33266
rect 1037 33264 1239 33266
rect 1273 33264 1475 33266
rect 1509 33264 1711 33298
rect 1745 33264 1947 33298
rect 1981 33266 2097 33298
rect 2149 33266 2165 33318
rect 2217 33266 2233 33318
rect 2285 33266 2301 33318
rect 2353 33266 2369 33318
rect 2421 33298 2437 33318
rect 2489 33266 2505 33318
rect 2557 33266 2573 33318
rect 2625 33266 2641 33318
rect 2693 33312 3036 33318
rect 3070 33312 3076 33346
rect 2693 33298 3076 33312
rect 2693 33266 2891 33298
rect 1981 33264 2183 33266
rect 2217 33264 2419 33266
rect 2453 33264 2655 33266
rect 2689 33264 2891 33266
rect 2925 33274 3076 33298
rect 2925 33264 3036 33274
rect 380 33255 3036 33264
rect 380 33221 386 33255
rect 420 33254 3036 33255
rect 420 33224 697 33254
rect 420 33221 531 33224
rect 380 33190 531 33221
rect 565 33202 697 33224
rect 749 33202 765 33254
rect 817 33202 833 33254
rect 885 33202 901 33254
rect 953 33202 969 33254
rect 1021 33224 1037 33254
rect 1089 33202 1105 33254
rect 1157 33202 1173 33254
rect 1225 33224 1241 33254
rect 1293 33224 2097 33254
rect 1225 33202 1239 33224
rect 1293 33202 1475 33224
rect 565 33190 767 33202
rect 801 33190 1003 33202
rect 1037 33190 1239 33202
rect 1273 33190 1475 33202
rect 1509 33190 1711 33224
rect 1745 33190 1947 33224
rect 1981 33202 2097 33224
rect 2149 33202 2165 33254
rect 2217 33202 2233 33254
rect 2285 33202 2301 33254
rect 2353 33202 2369 33254
rect 2421 33224 2437 33254
rect 2489 33202 2505 33254
rect 2557 33202 2573 33254
rect 2625 33202 2641 33254
rect 2693 33240 3036 33254
rect 3070 33240 3076 33274
rect 2693 33224 3076 33240
rect 2693 33202 2891 33224
rect 1981 33190 2183 33202
rect 2217 33190 2419 33202
rect 2453 33190 2655 33202
rect 2689 33190 2891 33202
rect 2925 33202 3076 33224
rect 2925 33190 3036 33202
rect 380 33183 3036 33190
rect 380 33149 386 33183
rect 420 33176 3036 33183
rect 420 33168 597 33176
tri 597 33168 605 33176 nw
tri 727 33168 735 33176 ne
rect 735 33168 833 33176
tri 833 33168 841 33176 nw
tri 963 33168 971 33176 ne
rect 971 33168 1069 33176
tri 1069 33168 1077 33176 nw
tri 1199 33168 1207 33176 ne
rect 1207 33168 1305 33176
tri 1305 33168 1313 33176 nw
tri 1435 33168 1443 33176 ne
rect 1443 33168 1541 33176
tri 1541 33168 1549 33176 nw
tri 1671 33168 1679 33176 ne
rect 1679 33168 1777 33176
tri 1777 33168 1785 33176 nw
tri 1907 33168 1915 33176 ne
rect 1915 33168 2013 33176
tri 2013 33168 2021 33176 nw
tri 2143 33168 2151 33176 ne
rect 2151 33168 2249 33176
tri 2249 33168 2257 33176 nw
tri 2379 33168 2387 33176 ne
rect 2387 33168 2485 33176
tri 2485 33168 2493 33176 nw
tri 2615 33168 2623 33176 ne
rect 2623 33168 2721 33176
tri 2721 33168 2729 33176 nw
tri 2851 33168 2859 33176 ne
rect 2859 33168 3036 33176
rect 3070 33168 3076 33202
rect 420 33150 579 33168
tri 579 33150 597 33168 nw
tri 735 33150 753 33168 ne
rect 753 33150 815 33168
tri 815 33150 833 33168 nw
tri 971 33150 989 33168 ne
rect 989 33150 1051 33168
tri 1051 33150 1069 33168 nw
tri 1207 33150 1225 33168 ne
rect 1225 33150 1287 33168
tri 1287 33150 1305 33168 nw
tri 1443 33150 1461 33168 ne
rect 1461 33150 1523 33168
tri 1523 33150 1541 33168 nw
tri 1679 33150 1697 33168 ne
rect 1697 33150 1759 33168
tri 1759 33150 1777 33168 nw
tri 1915 33150 1933 33168 ne
rect 1933 33150 1995 33168
tri 1995 33150 2013 33168 nw
tri 2151 33150 2169 33168 ne
rect 2169 33150 2231 33168
tri 2231 33150 2249 33168 nw
tri 2387 33150 2405 33168 ne
rect 2405 33150 2467 33168
tri 2467 33150 2485 33168 nw
tri 2623 33150 2641 33168 ne
rect 2641 33150 2703 33168
tri 2703 33150 2721 33168 nw
tri 2859 33150 2877 33168 ne
rect 2877 33150 3076 33168
rect 420 33149 531 33150
rect 380 33116 531 33149
rect 565 33116 571 33150
tri 571 33142 579 33150 nw
tri 753 33142 761 33150 ne
rect 380 33111 571 33116
rect 380 33077 386 33111
rect 420 33077 571 33111
rect 380 33076 571 33077
rect 380 33042 531 33076
rect 565 33042 571 33076
rect 380 33039 571 33042
rect 380 33005 386 33039
rect 420 33005 571 33039
rect 380 33002 571 33005
rect 380 32968 531 33002
rect 565 32968 571 33002
rect 380 32967 571 32968
rect 380 32933 386 32967
rect 420 32933 571 32967
rect 380 32928 571 32933
rect 380 32895 531 32928
rect 380 32861 386 32895
rect 420 32894 531 32895
rect 565 32894 571 32928
rect 420 32861 571 32894
rect 380 32854 571 32861
rect 380 32823 531 32854
rect 380 32789 386 32823
rect 420 32820 531 32823
rect 565 32820 571 32854
rect 420 32789 571 32820
rect 380 32780 571 32789
rect 380 32751 531 32780
rect 380 32717 386 32751
rect 420 32746 531 32751
rect 565 32746 571 32780
rect 420 32717 571 32746
rect 761 33116 767 33150
rect 801 33116 807 33150
tri 807 33142 815 33150 nw
tri 989 33142 997 33150 ne
rect 761 33076 807 33116
rect 761 33042 767 33076
rect 801 33042 807 33076
rect 761 33002 807 33042
rect 761 32968 767 33002
rect 801 32968 807 33002
rect 761 32928 807 32968
rect 761 32894 767 32928
rect 801 32894 807 32928
rect 761 32854 807 32894
rect 761 32820 767 32854
rect 801 32820 807 32854
rect 761 32780 807 32820
rect 761 32746 767 32780
rect 801 32746 807 32780
rect 761 32734 807 32746
rect 997 33116 1003 33150
rect 1037 33116 1043 33150
tri 1043 33142 1051 33150 nw
tri 1225 33142 1233 33150 ne
rect 997 33076 1043 33116
rect 997 33042 1003 33076
rect 1037 33042 1043 33076
rect 997 33002 1043 33042
rect 997 32968 1003 33002
rect 1037 32968 1043 33002
rect 997 32928 1043 32968
rect 997 32894 1003 32928
rect 1037 32894 1043 32928
rect 997 32854 1043 32894
rect 997 32820 1003 32854
rect 1037 32820 1043 32854
rect 997 32780 1043 32820
rect 997 32746 1003 32780
rect 1037 32746 1043 32780
rect 997 32734 1043 32746
rect 1233 33116 1239 33150
rect 1273 33116 1279 33150
tri 1279 33142 1287 33150 nw
tri 1461 33142 1469 33150 ne
rect 1233 33076 1279 33116
rect 1233 33042 1239 33076
rect 1273 33042 1279 33076
rect 1233 33002 1279 33042
rect 1233 32968 1239 33002
rect 1273 32968 1279 33002
rect 1233 32928 1279 32968
rect 1233 32894 1239 32928
rect 1273 32894 1279 32928
rect 1233 32854 1279 32894
rect 1233 32820 1239 32854
rect 1273 32820 1279 32854
rect 1233 32780 1279 32820
rect 1233 32746 1239 32780
rect 1273 32746 1279 32780
rect 1233 32734 1279 32746
rect 1469 33116 1475 33150
rect 1509 33116 1515 33150
tri 1515 33142 1523 33150 nw
tri 1697 33142 1705 33150 ne
rect 1469 33076 1515 33116
rect 1469 33042 1475 33076
rect 1509 33042 1515 33076
rect 1469 33002 1515 33042
rect 1469 32968 1475 33002
rect 1509 32968 1515 33002
rect 1469 32928 1515 32968
rect 1469 32894 1475 32928
rect 1509 32894 1515 32928
rect 1469 32854 1515 32894
rect 1469 32820 1475 32854
rect 1509 32820 1515 32854
rect 1469 32780 1515 32820
rect 1469 32746 1475 32780
rect 1509 32746 1515 32780
rect 1469 32734 1515 32746
rect 1705 33116 1711 33150
rect 1745 33116 1751 33150
tri 1751 33142 1759 33150 nw
tri 1933 33142 1941 33150 ne
rect 1705 33076 1751 33116
rect 1705 33042 1711 33076
rect 1745 33042 1751 33076
rect 1705 33002 1751 33042
rect 1705 32968 1711 33002
rect 1745 32968 1751 33002
rect 1705 32928 1751 32968
rect 1705 32894 1711 32928
rect 1745 32894 1751 32928
rect 1705 32854 1751 32894
rect 1705 32820 1711 32854
rect 1745 32820 1751 32854
rect 1705 32780 1751 32820
rect 1705 32746 1711 32780
rect 1745 32746 1751 32780
rect 1705 32734 1751 32746
rect 1941 33116 1947 33150
rect 1981 33116 1987 33150
tri 1987 33142 1995 33150 nw
tri 2169 33142 2177 33150 ne
rect 1941 33076 1987 33116
rect 1941 33042 1947 33076
rect 1981 33042 1987 33076
rect 1941 33002 1987 33042
rect 1941 32968 1947 33002
rect 1981 32968 1987 33002
rect 1941 32928 1987 32968
rect 1941 32894 1947 32928
rect 1981 32894 1987 32928
rect 1941 32854 1987 32894
rect 1941 32820 1947 32854
rect 1981 32820 1987 32854
rect 1941 32780 1987 32820
rect 1941 32746 1947 32780
rect 1981 32746 1987 32780
rect 1941 32734 1987 32746
rect 2177 33116 2183 33150
rect 2217 33116 2223 33150
tri 2223 33142 2231 33150 nw
tri 2405 33142 2413 33150 ne
rect 2177 33076 2223 33116
rect 2177 33042 2183 33076
rect 2217 33042 2223 33076
rect 2177 33002 2223 33042
rect 2177 32968 2183 33002
rect 2217 32968 2223 33002
rect 2177 32928 2223 32968
rect 2177 32894 2183 32928
rect 2217 32894 2223 32928
rect 2177 32854 2223 32894
rect 2177 32820 2183 32854
rect 2217 32820 2223 32854
rect 2177 32780 2223 32820
rect 2177 32746 2183 32780
rect 2217 32746 2223 32780
rect 2177 32734 2223 32746
rect 2413 33116 2419 33150
rect 2453 33116 2459 33150
tri 2459 33142 2467 33150 nw
tri 2641 33142 2649 33150 ne
rect 2413 33076 2459 33116
rect 2413 33042 2419 33076
rect 2453 33042 2459 33076
rect 2413 33002 2459 33042
rect 2413 32968 2419 33002
rect 2453 32968 2459 33002
rect 2413 32928 2459 32968
rect 2413 32894 2419 32928
rect 2453 32894 2459 32928
rect 2413 32854 2459 32894
rect 2413 32820 2419 32854
rect 2453 32820 2459 32854
rect 2413 32780 2459 32820
rect 2413 32746 2419 32780
rect 2453 32746 2459 32780
rect 2413 32734 2459 32746
rect 2649 33116 2655 33150
rect 2689 33116 2695 33150
tri 2695 33142 2703 33150 nw
tri 2877 33142 2885 33150 ne
rect 2649 33076 2695 33116
rect 2649 33042 2655 33076
rect 2689 33042 2695 33076
rect 2649 33002 2695 33042
rect 2649 32968 2655 33002
rect 2689 32968 2695 33002
rect 2649 32928 2695 32968
rect 2649 32894 2655 32928
rect 2689 32894 2695 32928
rect 2649 32854 2695 32894
rect 2649 32820 2655 32854
rect 2689 32820 2695 32854
rect 2649 32780 2695 32820
rect 2649 32746 2655 32780
rect 2689 32746 2695 32780
rect 2649 32734 2695 32746
rect 2885 33116 2891 33150
rect 2925 33130 3076 33150
rect 2925 33116 3036 33130
rect 2885 33096 3036 33116
rect 3070 33096 3076 33130
rect 2885 33076 3076 33096
rect 2885 33042 2891 33076
rect 2925 33058 3076 33076
rect 2925 33042 3036 33058
rect 2885 33024 3036 33042
rect 3070 33024 3076 33058
rect 2885 33002 3076 33024
rect 2885 32968 2891 33002
rect 2925 32986 3076 33002
rect 2925 32968 3036 32986
rect 2885 32952 3036 32968
rect 3070 32952 3076 32986
rect 2885 32928 3076 32952
rect 2885 32894 2891 32928
rect 2925 32914 3076 32928
rect 2925 32894 3036 32914
rect 2885 32880 3036 32894
rect 3070 32880 3076 32914
rect 2885 32854 3076 32880
rect 2885 32820 2891 32854
rect 2925 32842 3076 32854
rect 2925 32820 3036 32842
rect 2885 32808 3036 32820
rect 3070 32808 3076 32842
rect 2885 32780 3076 32808
rect 2885 32746 2891 32780
rect 2925 32770 3076 32780
rect 2925 32746 3036 32770
rect 2885 32736 3036 32746
rect 3070 32736 3076 32770
rect 380 32679 571 32717
rect 380 32645 386 32679
rect 420 32645 571 32679
rect 2885 32698 3076 32736
rect 380 32607 571 32645
rect 613 32664 1501 32673
rect 1553 32664 1569 32673
rect 1621 32664 1636 32673
rect 1688 32664 1703 32673
rect 1755 32664 1770 32673
rect 1822 32664 1837 32673
rect 1889 32664 2830 32673
rect 613 32630 625 32664
rect 659 32630 700 32664
rect 734 32630 775 32664
rect 809 32630 850 32664
rect 884 32630 925 32664
rect 959 32630 1000 32664
rect 1034 32630 1075 32664
rect 1109 32630 1150 32664
rect 1184 32630 1225 32664
rect 1259 32630 1300 32664
rect 1334 32630 1375 32664
rect 1409 32630 1450 32664
rect 1484 32630 1501 32664
rect 1559 32630 1569 32664
rect 1634 32630 1636 32664
rect 1889 32630 1896 32664
rect 1930 32630 1970 32664
rect 2004 32630 2044 32664
rect 2078 32630 2118 32664
rect 2152 32630 2192 32664
rect 2226 32630 2266 32664
rect 2300 32630 2340 32664
rect 2374 32630 2414 32664
rect 2448 32630 2488 32664
rect 2522 32630 2562 32664
rect 2596 32630 2636 32664
rect 2670 32630 2710 32664
rect 2744 32630 2784 32664
rect 2818 32630 2830 32664
rect 613 32621 1501 32630
rect 1553 32621 1569 32630
rect 1621 32621 1636 32630
rect 1688 32621 1703 32630
rect 1755 32621 1770 32630
rect 1822 32621 1837 32630
rect 1889 32621 2830 32630
rect 2885 32664 3036 32698
rect 3070 32664 3076 32698
rect 2885 32626 3076 32664
rect 380 32573 386 32607
rect 420 32573 571 32607
rect 380 32548 571 32573
rect 2885 32592 3036 32626
rect 3070 32592 3076 32626
rect 380 32535 531 32548
rect 380 32501 386 32535
rect 420 32514 531 32535
rect 565 32514 571 32548
rect 420 32501 571 32514
rect 380 32475 571 32501
rect 380 32463 531 32475
rect 380 32429 386 32463
rect 420 32441 531 32463
rect 565 32441 571 32475
rect 420 32429 571 32441
rect 380 32402 571 32429
rect 380 32391 531 32402
rect 380 32357 386 32391
rect 420 32368 531 32391
rect 565 32368 571 32402
rect 420 32357 571 32368
rect 380 32329 571 32357
rect 380 32319 531 32329
rect 380 32285 386 32319
rect 420 32295 531 32319
rect 565 32295 571 32329
rect 420 32285 571 32295
rect 380 32256 571 32285
rect 380 32247 531 32256
rect 380 32213 386 32247
rect 420 32222 531 32247
rect 565 32222 571 32256
rect 420 32213 571 32222
rect 380 32183 571 32213
rect 380 32175 531 32183
rect 380 32141 386 32175
rect 420 32149 531 32175
rect 565 32149 571 32183
rect 420 32141 571 32149
rect 380 32110 571 32141
rect 380 32103 531 32110
rect 380 32069 386 32103
rect 420 32076 531 32103
rect 565 32076 571 32110
rect 761 32548 807 32560
rect 761 32514 767 32548
rect 801 32514 807 32548
rect 761 32475 807 32514
rect 761 32441 767 32475
rect 801 32441 807 32475
rect 761 32402 807 32441
rect 761 32368 767 32402
rect 801 32368 807 32402
rect 761 32329 807 32368
rect 761 32295 767 32329
rect 801 32295 807 32329
rect 761 32256 807 32295
rect 761 32222 767 32256
rect 801 32222 807 32256
rect 761 32183 807 32222
rect 761 32149 767 32183
rect 801 32149 807 32183
rect 761 32110 807 32149
tri 571 32076 576 32081 sw
tri 756 32076 761 32081 se
rect 761 32076 767 32110
rect 801 32076 807 32110
rect 997 32548 1043 32560
rect 997 32514 1003 32548
rect 1037 32514 1043 32548
rect 997 32475 1043 32514
rect 997 32441 1003 32475
rect 1037 32441 1043 32475
rect 997 32402 1043 32441
rect 997 32368 1003 32402
rect 1037 32368 1043 32402
rect 997 32329 1043 32368
rect 997 32295 1003 32329
rect 1037 32295 1043 32329
rect 997 32256 1043 32295
rect 997 32222 1003 32256
rect 1037 32222 1043 32256
rect 997 32183 1043 32222
rect 997 32149 1003 32183
rect 1037 32149 1043 32183
rect 997 32110 1043 32149
tri 807 32076 812 32081 sw
tri 992 32076 997 32081 se
rect 997 32076 1003 32110
rect 1037 32076 1043 32110
rect 1233 32548 1279 32560
rect 1233 32514 1239 32548
rect 1273 32514 1279 32548
rect 1233 32475 1279 32514
rect 1233 32441 1239 32475
rect 1273 32441 1279 32475
rect 1233 32402 1279 32441
rect 1233 32368 1239 32402
rect 1273 32368 1279 32402
rect 1233 32329 1279 32368
rect 1233 32295 1239 32329
rect 1273 32295 1279 32329
rect 1233 32256 1279 32295
rect 1233 32222 1239 32256
rect 1273 32222 1279 32256
rect 1233 32183 1279 32222
rect 1233 32149 1239 32183
rect 1273 32149 1279 32183
rect 1233 32110 1279 32149
tri 1043 32076 1048 32081 sw
tri 1228 32076 1233 32081 se
rect 1233 32076 1239 32110
rect 1273 32076 1279 32110
rect 1469 32548 1515 32560
rect 1469 32514 1475 32548
rect 1509 32514 1515 32548
rect 1469 32475 1515 32514
rect 1469 32441 1475 32475
rect 1509 32441 1515 32475
rect 1469 32402 1515 32441
rect 1469 32368 1475 32402
rect 1509 32368 1515 32402
rect 1469 32329 1515 32368
rect 1469 32295 1475 32329
rect 1509 32295 1515 32329
rect 1469 32256 1515 32295
rect 1469 32222 1475 32256
rect 1509 32222 1515 32256
rect 1469 32183 1515 32222
rect 1469 32149 1475 32183
rect 1509 32149 1515 32183
rect 1469 32110 1515 32149
tri 1279 32076 1284 32081 sw
tri 1464 32076 1469 32081 se
rect 1469 32076 1475 32110
rect 1509 32076 1515 32110
rect 1705 32548 1751 32560
rect 1705 32514 1711 32548
rect 1745 32514 1751 32548
rect 1705 32475 1751 32514
rect 1705 32441 1711 32475
rect 1745 32441 1751 32475
rect 1705 32402 1751 32441
rect 1705 32368 1711 32402
rect 1745 32368 1751 32402
rect 1705 32329 1751 32368
rect 1705 32295 1711 32329
rect 1745 32295 1751 32329
rect 1705 32256 1751 32295
rect 1705 32222 1711 32256
rect 1745 32222 1751 32256
rect 1705 32183 1751 32222
rect 1705 32149 1711 32183
rect 1745 32149 1751 32183
rect 1705 32110 1751 32149
tri 1515 32076 1520 32081 sw
tri 1700 32076 1705 32081 se
rect 1705 32076 1711 32110
rect 1745 32076 1751 32110
rect 1941 32548 1987 32560
rect 1941 32514 1947 32548
rect 1981 32514 1987 32548
rect 1941 32475 1987 32514
rect 1941 32441 1947 32475
rect 1981 32441 1987 32475
rect 1941 32402 1987 32441
rect 1941 32368 1947 32402
rect 1981 32368 1987 32402
rect 1941 32329 1987 32368
rect 1941 32295 1947 32329
rect 1981 32295 1987 32329
rect 1941 32256 1987 32295
rect 1941 32222 1947 32256
rect 1981 32222 1987 32256
rect 1941 32183 1987 32222
rect 1941 32149 1947 32183
rect 1981 32149 1987 32183
rect 1941 32110 1987 32149
tri 1751 32076 1756 32081 sw
tri 1936 32076 1941 32081 se
rect 1941 32076 1947 32110
rect 1981 32076 1987 32110
rect 2177 32548 2223 32560
rect 2177 32514 2183 32548
rect 2217 32514 2223 32548
rect 2177 32475 2223 32514
rect 2177 32441 2183 32475
rect 2217 32441 2223 32475
rect 2177 32402 2223 32441
rect 2177 32368 2183 32402
rect 2217 32368 2223 32402
rect 2177 32329 2223 32368
rect 2177 32295 2183 32329
rect 2217 32295 2223 32329
rect 2177 32256 2223 32295
rect 2177 32222 2183 32256
rect 2217 32222 2223 32256
rect 2177 32183 2223 32222
rect 2177 32149 2183 32183
rect 2217 32149 2223 32183
rect 2177 32110 2223 32149
tri 1987 32076 1992 32081 sw
tri 2172 32076 2177 32081 se
rect 2177 32076 2183 32110
rect 2217 32076 2223 32110
rect 2413 32548 2459 32560
rect 2413 32514 2419 32548
rect 2453 32514 2459 32548
rect 2413 32475 2459 32514
rect 2413 32441 2419 32475
rect 2453 32441 2459 32475
rect 2413 32402 2459 32441
rect 2413 32368 2419 32402
rect 2453 32368 2459 32402
rect 2413 32329 2459 32368
rect 2413 32295 2419 32329
rect 2453 32295 2459 32329
rect 2413 32256 2459 32295
rect 2413 32222 2419 32256
rect 2453 32222 2459 32256
rect 2413 32183 2459 32222
rect 2413 32149 2419 32183
rect 2453 32149 2459 32183
rect 2413 32110 2459 32149
tri 2223 32076 2228 32081 sw
tri 2408 32076 2413 32081 se
rect 2413 32076 2419 32110
rect 2453 32076 2459 32110
rect 2649 32548 2695 32560
rect 2649 32514 2655 32548
rect 2689 32514 2695 32548
rect 2649 32475 2695 32514
rect 2649 32441 2655 32475
rect 2689 32441 2695 32475
rect 2649 32402 2695 32441
rect 2649 32368 2655 32402
rect 2689 32368 2695 32402
rect 2649 32329 2695 32368
rect 2649 32295 2655 32329
rect 2689 32295 2695 32329
rect 2649 32256 2695 32295
rect 2649 32222 2655 32256
rect 2689 32222 2695 32256
rect 2649 32183 2695 32222
rect 2649 32149 2655 32183
rect 2689 32149 2695 32183
rect 2649 32110 2695 32149
tri 2459 32076 2464 32081 sw
tri 2644 32076 2649 32081 se
rect 2649 32076 2655 32110
rect 2689 32076 2695 32110
rect 2885 32554 3076 32592
rect 2885 32548 3036 32554
rect 2885 32514 2891 32548
rect 2925 32520 3036 32548
rect 3070 32520 3076 32554
rect 2925 32514 3076 32520
rect 2885 32482 3076 32514
rect 2885 32475 3036 32482
rect 2885 32441 2891 32475
rect 2925 32448 3036 32475
rect 3070 32448 3076 32482
rect 2925 32441 3076 32448
rect 2885 32410 3076 32441
rect 2885 32402 3036 32410
rect 2885 32368 2891 32402
rect 2925 32376 3036 32402
rect 3070 32376 3076 32410
rect 2925 32368 3076 32376
rect 2885 32338 3076 32368
rect 2885 32329 3036 32338
rect 2885 32295 2891 32329
rect 2925 32304 3036 32329
rect 3070 32304 3076 32338
rect 2925 32295 3076 32304
rect 2885 32266 3076 32295
rect 2885 32256 3036 32266
rect 2885 32222 2891 32256
rect 2925 32232 3036 32256
rect 3070 32232 3076 32266
rect 2925 32222 3076 32232
rect 2885 32194 3076 32222
rect 2885 32183 3036 32194
rect 2885 32149 2891 32183
rect 2925 32160 3036 32183
rect 3070 32160 3076 32194
rect 2925 32149 3076 32160
rect 2885 32122 3076 32149
rect 2885 32110 3036 32122
tri 2695 32076 2700 32081 sw
tri 2880 32076 2885 32081 se
rect 2885 32076 2891 32110
rect 2925 32088 3036 32110
rect 3070 32088 3076 32122
rect 2925 32076 3076 32088
rect 420 32069 576 32076
rect 380 32064 576 32069
tri 576 32064 588 32076 sw
tri 744 32064 756 32076 se
rect 756 32064 812 32076
tri 812 32064 824 32076 sw
tri 980 32064 992 32076 se
rect 992 32064 1048 32076
tri 1048 32064 1060 32076 sw
tri 1216 32064 1228 32076 se
rect 1228 32064 1284 32076
tri 1284 32064 1296 32076 sw
tri 1452 32064 1464 32076 se
rect 1464 32064 1520 32076
tri 1520 32064 1532 32076 sw
tri 1688 32064 1700 32076 se
rect 1700 32064 1756 32076
tri 1756 32064 1768 32076 sw
tri 1924 32064 1936 32076 se
rect 1936 32064 1992 32076
tri 1992 32064 2004 32076 sw
tri 2160 32064 2172 32076 se
rect 2172 32064 2228 32076
tri 2228 32064 2240 32076 sw
tri 2396 32064 2408 32076 se
rect 2408 32064 2464 32076
tri 2464 32064 2476 32076 sw
tri 2632 32064 2644 32076 se
rect 2644 32064 2700 32076
tri 2700 32064 2712 32076 sw
tri 2868 32064 2880 32076 se
rect 2880 32064 3076 32076
rect 380 32050 588 32064
tri 588 32050 602 32064 sw
tri 730 32050 744 32064 se
rect 744 32050 824 32064
tri 824 32050 838 32064 sw
tri 966 32050 980 32064 se
rect 980 32050 1060 32064
tri 1060 32050 1074 32064 sw
tri 1202 32050 1216 32064 se
rect 1216 32050 1296 32064
tri 1296 32050 1310 32064 sw
tri 1438 32050 1452 32064 se
rect 1452 32050 1532 32064
tri 1532 32050 1546 32064 sw
tri 1674 32050 1688 32064 se
rect 1688 32050 1768 32064
tri 1768 32050 1782 32064 sw
tri 1910 32050 1924 32064 se
rect 1924 32050 2004 32064
tri 2004 32050 2018 32064 sw
tri 2146 32050 2160 32064 se
rect 2160 32050 2240 32064
tri 2240 32050 2254 32064 sw
tri 2382 32050 2396 32064 se
rect 2396 32050 2476 32064
tri 2476 32050 2490 32064 sw
tri 2618 32050 2632 32064 se
rect 2632 32050 2712 32064
tri 2712 32050 2726 32064 sw
tri 2854 32050 2868 32064 se
rect 2868 32050 3076 32064
rect 380 32047 602 32050
tri 602 32047 605 32050 sw
tri 727 32047 730 32050 se
rect 730 32047 838 32050
tri 838 32047 841 32050 sw
tri 963 32047 966 32050 se
rect 966 32047 1074 32050
tri 1074 32047 1077 32050 sw
tri 1199 32047 1202 32050 se
rect 1202 32047 1310 32050
tri 1310 32047 1313 32050 sw
tri 1435 32047 1438 32050 se
rect 1438 32047 1546 32050
tri 1546 32047 1549 32050 sw
tri 1671 32047 1674 32050 se
rect 1674 32047 1782 32050
tri 1782 32047 1785 32050 sw
tri 1907 32047 1910 32050 se
rect 1910 32047 2018 32050
tri 2018 32047 2021 32050 sw
tri 2143 32047 2146 32050 se
rect 2146 32047 2254 32050
tri 2254 32047 2257 32050 sw
tri 2379 32047 2382 32050 se
rect 2382 32047 2490 32050
tri 2490 32047 2493 32050 sw
tri 2615 32047 2618 32050 se
rect 2618 32047 2726 32050
tri 2726 32047 2729 32050 sw
tri 2851 32047 2854 32050 se
rect 2854 32047 3036 32050
rect 380 32037 3036 32047
rect 380 32031 531 32037
rect 380 31997 386 32031
rect 420 32003 531 32031
rect 565 32021 767 32037
rect 801 32021 1003 32037
rect 1037 32021 1239 32037
rect 1273 32021 1475 32037
rect 565 32003 697 32021
rect 420 31997 697 32003
rect 380 31969 697 31997
rect 749 31969 765 32021
rect 817 31969 833 32021
rect 885 31969 901 32021
rect 953 31969 969 32021
rect 1021 31969 1037 32003
rect 1089 31969 1105 32021
rect 1157 31969 1173 32021
rect 1225 32003 1239 32021
rect 1293 32003 1475 32021
rect 1509 32003 1711 32037
rect 1745 32003 1947 32037
rect 1981 32021 2183 32037
rect 2217 32021 2419 32037
rect 2453 32021 2655 32037
rect 2689 32021 2891 32037
rect 1981 32003 2097 32021
rect 1225 31969 1241 32003
rect 1293 31969 2097 32003
rect 2149 31969 2165 32021
rect 2217 31969 2233 32021
rect 2285 31969 2301 32021
rect 2353 31969 2369 32021
rect 2421 31969 2437 32003
rect 2489 31969 2505 32021
rect 2557 31969 2573 32021
rect 2625 31969 2641 32021
rect 2693 32003 2891 32021
rect 2925 32016 3036 32037
rect 3070 32016 3076 32050
rect 2925 32003 3076 32016
rect 2693 31978 3076 32003
rect 2693 31969 3036 31978
rect 380 31964 3036 31969
rect 380 31959 531 31964
rect 380 31925 386 31959
rect 420 31930 531 31959
rect 565 31957 767 31964
rect 801 31957 1003 31964
rect 1037 31957 1239 31964
rect 1273 31957 1475 31964
rect 565 31930 697 31957
rect 420 31925 697 31930
rect 380 31905 697 31925
rect 749 31905 765 31957
rect 817 31905 833 31957
rect 885 31905 901 31957
rect 953 31905 969 31957
rect 1021 31905 1037 31930
rect 1089 31905 1105 31957
rect 1157 31905 1173 31957
rect 1225 31930 1239 31957
rect 1293 31930 1475 31957
rect 1509 31930 1711 31964
rect 1745 31930 1947 31964
rect 1981 31957 2183 31964
rect 2217 31957 2419 31964
rect 2453 31957 2655 31964
rect 2689 31957 2891 31964
rect 1981 31930 2097 31957
rect 1225 31905 1241 31930
rect 1293 31905 2097 31930
rect 2149 31905 2165 31957
rect 2217 31905 2233 31957
rect 2285 31905 2301 31957
rect 2353 31905 2369 31957
rect 2421 31905 2437 31930
rect 2489 31905 2505 31957
rect 2557 31905 2573 31957
rect 2625 31905 2641 31957
rect 2693 31930 2891 31957
rect 2925 31944 3036 31964
rect 3070 31944 3076 31978
rect 2925 31930 3076 31944
rect 2693 31906 3076 31930
rect 2693 31905 3036 31906
rect 380 31893 3036 31905
rect 380 31891 697 31893
rect 380 31887 531 31891
rect 380 31853 386 31887
rect 420 31857 531 31887
rect 565 31857 697 31891
rect 420 31853 697 31857
rect 380 31841 697 31853
rect 749 31841 765 31893
rect 817 31841 833 31893
rect 885 31841 901 31893
rect 953 31841 969 31893
rect 1021 31891 1037 31893
rect 1021 31841 1037 31857
rect 1089 31841 1105 31893
rect 1157 31841 1173 31893
rect 1225 31891 1241 31893
rect 1293 31891 2097 31893
rect 1225 31857 1239 31891
rect 1293 31857 1475 31891
rect 1509 31857 1711 31891
rect 1745 31857 1947 31891
rect 1981 31857 2097 31891
rect 1225 31841 1241 31857
rect 1293 31841 2097 31857
rect 2149 31841 2165 31893
rect 2217 31841 2233 31893
rect 2285 31841 2301 31893
rect 2353 31841 2369 31893
rect 2421 31891 2437 31893
rect 2421 31841 2437 31857
rect 2489 31841 2505 31893
rect 2557 31841 2573 31893
rect 2625 31841 2641 31893
rect 2693 31891 3036 31893
rect 2693 31857 2891 31891
rect 2925 31872 3036 31891
rect 3070 31872 3076 31906
rect 2925 31857 3076 31872
rect 2693 31841 3076 31857
rect 380 31834 3076 31841
rect 380 31829 3036 31834
rect 380 31818 697 31829
rect 380 31815 531 31818
rect 380 31781 386 31815
rect 420 31784 531 31815
rect 565 31784 697 31818
rect 420 31781 697 31784
rect 380 31777 697 31781
rect 749 31777 765 31829
rect 817 31777 833 31829
rect 885 31777 901 31829
rect 953 31777 969 31829
rect 1021 31818 1037 31829
rect 1021 31777 1037 31784
rect 1089 31777 1105 31829
rect 1157 31777 1173 31829
rect 1225 31818 1241 31829
rect 1293 31818 2097 31829
rect 1225 31784 1239 31818
rect 1293 31784 1475 31818
rect 1509 31784 1711 31818
rect 1745 31784 1947 31818
rect 1981 31784 2097 31818
rect 1225 31777 1241 31784
rect 1293 31777 2097 31784
rect 2149 31777 2165 31829
rect 2217 31777 2233 31829
rect 2285 31777 2301 31829
rect 2353 31777 2369 31829
rect 2421 31818 2437 31829
rect 2421 31777 2437 31784
rect 2489 31777 2505 31829
rect 2557 31777 2573 31829
rect 2625 31777 2641 31829
rect 2693 31818 3036 31829
rect 2693 31784 2891 31818
rect 2925 31800 3036 31818
rect 3070 31800 3076 31834
rect 2925 31784 3076 31800
rect 2693 31777 3076 31784
rect 380 31765 3076 31777
rect 380 31745 697 31765
rect 380 31743 531 31745
rect 380 31709 386 31743
rect 420 31711 531 31743
rect 565 31713 697 31745
rect 749 31713 765 31765
rect 817 31713 833 31765
rect 885 31713 901 31765
rect 953 31713 969 31765
rect 1021 31745 1037 31765
rect 1089 31713 1105 31765
rect 1157 31713 1173 31765
rect 1225 31745 1241 31765
rect 1293 31745 2097 31765
rect 1225 31713 1239 31745
rect 1293 31713 1475 31745
rect 565 31711 767 31713
rect 801 31711 1003 31713
rect 1037 31711 1239 31713
rect 1273 31711 1475 31713
rect 1509 31711 1711 31745
rect 1745 31711 1947 31745
rect 1981 31713 2097 31745
rect 2149 31713 2165 31765
rect 2217 31713 2233 31765
rect 2285 31713 2301 31765
rect 2353 31713 2369 31765
rect 2421 31745 2437 31765
rect 2489 31713 2505 31765
rect 2557 31713 2573 31765
rect 2625 31713 2641 31765
rect 2693 31762 3076 31765
rect 2693 31745 3036 31762
rect 2693 31713 2891 31745
rect 1981 31711 2183 31713
rect 2217 31711 2419 31713
rect 2453 31711 2655 31713
rect 2689 31711 2891 31713
rect 2925 31728 3036 31745
rect 3070 31728 3076 31762
rect 2925 31711 3076 31728
rect 420 31709 3076 31711
rect 380 31701 3076 31709
rect 380 31672 697 31701
rect 380 31671 531 31672
rect 380 31637 386 31671
rect 420 31638 531 31671
rect 565 31649 697 31672
rect 749 31649 765 31701
rect 817 31649 833 31701
rect 885 31649 901 31701
rect 953 31649 969 31701
rect 1021 31672 1037 31701
rect 1089 31649 1105 31701
rect 1157 31649 1173 31701
rect 1225 31672 1241 31701
rect 1293 31672 2097 31701
rect 1225 31649 1239 31672
rect 1293 31649 1475 31672
rect 565 31638 767 31649
rect 801 31638 1003 31649
rect 1037 31638 1239 31649
rect 1273 31638 1475 31649
rect 1509 31638 1711 31672
rect 1745 31638 1947 31672
rect 1981 31649 2097 31672
rect 2149 31649 2165 31701
rect 2217 31649 2233 31701
rect 2285 31649 2301 31701
rect 2353 31649 2369 31701
rect 2421 31672 2437 31701
rect 2489 31649 2505 31701
rect 2557 31649 2573 31701
rect 2625 31649 2641 31701
rect 2693 31690 3076 31701
rect 2693 31672 3036 31690
rect 2693 31649 2891 31672
rect 1981 31638 2183 31649
rect 2217 31638 2419 31649
rect 2453 31638 2655 31649
rect 2689 31638 2891 31649
rect 2925 31656 3036 31672
rect 3070 31656 3076 31690
rect 2925 31638 3076 31656
rect 420 31637 3076 31638
rect 380 31599 697 31637
rect 380 31565 386 31599
rect 420 31598 697 31599
rect 420 31565 531 31598
rect 380 31564 531 31565
rect 565 31585 697 31598
rect 749 31585 765 31637
rect 817 31585 833 31637
rect 885 31585 901 31637
rect 953 31585 969 31637
rect 1021 31598 1037 31637
rect 1089 31585 1105 31637
rect 1157 31585 1173 31637
rect 1225 31598 1241 31637
rect 1293 31598 2097 31637
rect 1225 31585 1239 31598
rect 1293 31585 1475 31598
rect 565 31573 767 31585
rect 801 31573 1003 31585
rect 1037 31573 1239 31585
rect 1273 31573 1475 31585
rect 565 31564 697 31573
rect 380 31527 697 31564
rect 380 31493 386 31527
rect 420 31524 697 31527
rect 420 31493 531 31524
rect 380 31490 531 31493
rect 565 31521 697 31524
rect 749 31521 765 31573
rect 817 31521 833 31573
rect 885 31521 901 31573
rect 953 31521 969 31573
rect 1021 31524 1037 31564
rect 1089 31521 1105 31573
rect 1157 31521 1173 31573
rect 1225 31564 1239 31573
rect 1293 31564 1475 31573
rect 1509 31564 1711 31598
rect 1745 31564 1947 31598
rect 1981 31585 2097 31598
rect 2149 31585 2165 31637
rect 2217 31585 2233 31637
rect 2285 31585 2301 31637
rect 2353 31585 2369 31637
rect 2421 31598 2437 31637
rect 2489 31585 2505 31637
rect 2557 31585 2573 31637
rect 2625 31585 2641 31637
rect 2693 31618 3076 31637
rect 2693 31598 3036 31618
rect 2693 31585 2891 31598
rect 1981 31573 2183 31585
rect 2217 31573 2419 31585
rect 2453 31573 2655 31585
rect 2689 31573 2891 31585
rect 1981 31564 2097 31573
rect 1225 31524 1241 31564
rect 1293 31524 2097 31564
rect 1225 31521 1239 31524
rect 1293 31521 1475 31524
rect 565 31509 767 31521
rect 801 31509 1003 31521
rect 1037 31509 1239 31521
rect 1273 31509 1475 31521
rect 565 31490 697 31509
rect 380 31457 697 31490
rect 749 31457 765 31509
rect 817 31457 833 31509
rect 885 31457 901 31509
rect 953 31457 969 31509
rect 1021 31457 1037 31490
rect 1089 31457 1105 31509
rect 1157 31457 1173 31509
rect 1225 31490 1239 31509
rect 1293 31490 1475 31509
rect 1509 31490 1711 31524
rect 1745 31490 1947 31524
rect 1981 31521 2097 31524
rect 2149 31521 2165 31573
rect 2217 31521 2233 31573
rect 2285 31521 2301 31573
rect 2353 31521 2369 31573
rect 2421 31524 2437 31564
rect 2489 31521 2505 31573
rect 2557 31521 2573 31573
rect 2625 31521 2641 31573
rect 2693 31564 2891 31573
rect 2925 31584 3036 31598
rect 3070 31584 3076 31618
rect 2925 31564 3076 31584
rect 2693 31546 3076 31564
rect 2693 31524 3036 31546
rect 2693 31521 2891 31524
rect 1981 31509 2183 31521
rect 2217 31509 2419 31521
rect 2453 31509 2655 31521
rect 2689 31509 2891 31521
rect 1981 31490 2097 31509
rect 1225 31457 1241 31490
rect 1293 31457 2097 31490
rect 2149 31457 2165 31509
rect 2217 31457 2233 31509
rect 2285 31457 2301 31509
rect 2353 31457 2369 31509
rect 2421 31457 2437 31490
rect 2489 31457 2505 31509
rect 2557 31457 2573 31509
rect 2625 31457 2641 31509
rect 2693 31490 2891 31509
rect 2925 31512 3036 31524
rect 3070 31512 3076 31546
rect 2925 31490 3076 31512
rect 2693 31474 3076 31490
rect 2693 31457 3036 31474
rect 380 31455 3036 31457
rect 380 31421 386 31455
rect 420 31450 3036 31455
rect 420 31421 531 31450
rect 380 31416 531 31421
rect 565 31445 767 31450
rect 801 31445 1003 31450
rect 1037 31445 1239 31450
rect 1273 31445 1475 31450
rect 565 31416 697 31445
rect 380 31393 697 31416
rect 749 31393 765 31445
rect 817 31393 833 31445
rect 885 31393 901 31445
rect 953 31393 969 31445
rect 1021 31393 1037 31416
rect 1089 31393 1105 31445
rect 1157 31393 1173 31445
rect 1225 31416 1239 31445
rect 1293 31416 1475 31445
rect 1509 31416 1711 31450
rect 1745 31416 1947 31450
rect 1981 31445 2183 31450
rect 2217 31445 2419 31450
rect 2453 31445 2655 31450
rect 2689 31445 2891 31450
rect 1981 31416 2097 31445
rect 1225 31393 1241 31416
rect 1293 31393 2097 31416
rect 2149 31393 2165 31445
rect 2217 31393 2233 31445
rect 2285 31393 2301 31445
rect 2353 31393 2369 31445
rect 2421 31393 2437 31416
rect 2489 31393 2505 31445
rect 2557 31393 2573 31445
rect 2625 31393 2641 31445
rect 2693 31416 2891 31445
rect 2925 31440 3036 31450
rect 3070 31440 3076 31474
rect 2925 31416 3076 31440
rect 2693 31402 3076 31416
rect 2693 31393 3036 31402
rect 380 31383 3036 31393
rect 380 31349 386 31383
rect 420 31381 3036 31383
rect 420 31376 697 31381
rect 420 31349 531 31376
rect 380 31342 531 31349
rect 565 31342 697 31376
rect 380 31329 697 31342
rect 749 31329 765 31381
rect 817 31329 833 31381
rect 885 31329 901 31381
rect 953 31329 969 31381
rect 1021 31376 1037 31381
rect 1021 31329 1037 31342
rect 1089 31329 1105 31381
rect 1157 31329 1173 31381
rect 1225 31376 1241 31381
rect 1293 31376 2097 31381
rect 1225 31342 1239 31376
rect 1293 31342 1475 31376
rect 1509 31342 1711 31376
rect 1745 31342 1947 31376
rect 1981 31342 2097 31376
rect 1225 31329 1241 31342
rect 1293 31329 2097 31342
rect 2149 31329 2165 31381
rect 2217 31329 2233 31381
rect 2285 31329 2301 31381
rect 2353 31329 2369 31381
rect 2421 31376 2437 31381
rect 2421 31329 2437 31342
rect 2489 31329 2505 31381
rect 2557 31329 2573 31381
rect 2625 31329 2641 31381
rect 2693 31376 3036 31381
rect 2693 31342 2891 31376
rect 2925 31368 3036 31376
rect 3070 31368 3076 31402
rect 2925 31342 3076 31368
rect 2693 31330 3076 31342
rect 2693 31329 3036 31330
rect 380 31317 3036 31329
rect 380 31311 697 31317
rect 380 31277 386 31311
rect 420 31302 697 31311
rect 420 31277 531 31302
rect 380 31268 531 31277
rect 565 31268 697 31302
rect 380 31265 697 31268
rect 749 31265 765 31317
rect 817 31265 833 31317
rect 885 31265 901 31317
rect 953 31265 969 31317
rect 1021 31302 1037 31317
rect 1021 31265 1037 31268
rect 1089 31265 1105 31317
rect 1157 31265 1173 31317
rect 1225 31302 1241 31317
rect 1293 31302 2097 31317
rect 1225 31268 1239 31302
rect 1293 31268 1475 31302
rect 1509 31268 1711 31302
rect 1745 31268 1947 31302
rect 1981 31268 2097 31302
rect 1225 31265 1241 31268
rect 1293 31265 2097 31268
rect 2149 31265 2165 31317
rect 2217 31265 2233 31317
rect 2285 31265 2301 31317
rect 2353 31265 2369 31317
rect 2421 31302 2437 31317
rect 2421 31265 2437 31268
rect 2489 31265 2505 31317
rect 2557 31265 2573 31317
rect 2625 31265 2641 31317
rect 2693 31302 3036 31317
rect 2693 31268 2891 31302
rect 2925 31296 3036 31302
rect 3070 31296 3076 31330
rect 2925 31268 3076 31296
rect 2693 31265 3076 31268
rect 380 31258 3076 31265
rect 380 31253 3036 31258
rect 380 31239 697 31253
rect 380 31205 386 31239
rect 420 31228 697 31239
rect 420 31205 531 31228
rect 380 31194 531 31205
rect 565 31201 697 31228
rect 749 31201 765 31253
rect 817 31201 833 31253
rect 885 31201 901 31253
rect 953 31201 969 31253
rect 1021 31228 1037 31253
rect 1089 31201 1105 31253
rect 1157 31201 1173 31253
rect 1225 31228 1241 31253
rect 1293 31228 2097 31253
rect 1225 31201 1239 31228
rect 1293 31201 1475 31228
rect 565 31194 767 31201
rect 801 31194 1003 31201
rect 1037 31194 1239 31201
rect 1273 31194 1475 31201
rect 1509 31194 1711 31228
rect 1745 31194 1947 31228
rect 1981 31201 2097 31228
rect 2149 31201 2165 31253
rect 2217 31201 2233 31253
rect 2285 31201 2301 31253
rect 2353 31201 2369 31253
rect 2421 31228 2437 31253
rect 2489 31201 2505 31253
rect 2557 31201 2573 31253
rect 2625 31201 2641 31253
rect 2693 31228 3036 31253
rect 2693 31201 2891 31228
rect 1981 31194 2183 31201
rect 2217 31194 2419 31201
rect 2453 31194 2655 31201
rect 2689 31194 2891 31201
rect 2925 31224 3036 31228
rect 3070 31224 3076 31258
rect 2925 31194 3076 31224
rect 380 31189 3076 31194
rect 380 31167 697 31189
rect 380 31133 386 31167
rect 420 31154 697 31167
rect 420 31133 531 31154
rect 380 31120 531 31133
rect 565 31137 697 31154
rect 749 31137 765 31189
rect 817 31137 833 31189
rect 885 31137 901 31189
rect 953 31137 969 31189
rect 1021 31154 1037 31189
rect 1089 31137 1105 31189
rect 1157 31137 1173 31189
rect 1225 31154 1241 31189
rect 1293 31154 2097 31189
rect 1225 31137 1239 31154
rect 1293 31137 1475 31154
rect 565 31125 767 31137
rect 801 31125 1003 31137
rect 1037 31125 1239 31137
rect 1273 31125 1475 31137
rect 565 31120 697 31125
rect 380 31095 697 31120
rect 380 31061 386 31095
rect 420 31080 697 31095
rect 420 31061 531 31080
rect 380 31046 531 31061
rect 565 31073 697 31080
rect 749 31073 765 31125
rect 817 31073 833 31125
rect 885 31073 901 31125
rect 953 31073 969 31125
rect 1021 31080 1037 31120
rect 1089 31073 1105 31125
rect 1157 31073 1173 31125
rect 1225 31120 1239 31125
rect 1293 31120 1475 31125
rect 1509 31120 1711 31154
rect 1745 31120 1947 31154
rect 1981 31137 2097 31154
rect 2149 31137 2165 31189
rect 2217 31137 2233 31189
rect 2285 31137 2301 31189
rect 2353 31137 2369 31189
rect 2421 31154 2437 31189
rect 2489 31137 2505 31189
rect 2557 31137 2573 31189
rect 2625 31137 2641 31189
rect 2693 31186 3076 31189
rect 2693 31154 3036 31186
rect 2693 31137 2891 31154
rect 1981 31125 2183 31137
rect 2217 31125 2419 31137
rect 2453 31125 2655 31137
rect 2689 31125 2891 31137
rect 1981 31120 2097 31125
rect 1225 31080 1241 31120
rect 1293 31080 2097 31120
rect 1225 31073 1239 31080
rect 1293 31073 1475 31080
rect 565 31047 767 31073
rect 565 31046 604 31047
tri 604 31046 605 31047 nw
tri 727 31046 728 31047 ne
rect 728 31046 767 31047
rect 801 31047 1003 31073
rect 801 31046 840 31047
tri 840 31046 841 31047 nw
tri 963 31046 964 31047 ne
rect 964 31046 1003 31047
rect 1037 31047 1239 31073
rect 1037 31046 1076 31047
tri 1076 31046 1077 31047 nw
tri 1199 31046 1200 31047 ne
rect 1200 31046 1239 31047
rect 1273 31047 1475 31073
rect 1273 31046 1312 31047
tri 1312 31046 1313 31047 nw
tri 1435 31046 1436 31047 ne
rect 1436 31046 1475 31047
rect 1509 31047 1711 31080
rect 1509 31046 1548 31047
tri 1548 31046 1549 31047 nw
tri 1671 31046 1672 31047 ne
rect 1672 31046 1711 31047
rect 1745 31047 1947 31080
rect 1745 31046 1784 31047
tri 1784 31046 1785 31047 nw
tri 1907 31046 1908 31047 ne
rect 1908 31046 1947 31047
rect 1981 31073 2097 31080
rect 2149 31073 2165 31125
rect 2217 31073 2233 31125
rect 2285 31073 2301 31125
rect 2353 31073 2369 31125
rect 2421 31080 2437 31120
rect 2489 31073 2505 31125
rect 2557 31073 2573 31125
rect 2625 31073 2641 31125
rect 2693 31120 2891 31125
rect 2925 31152 3036 31154
rect 3070 31152 3076 31186
rect 2925 31120 3076 31152
rect 2693 31114 3076 31120
rect 2693 31080 3036 31114
rect 3070 31080 3076 31114
rect 2693 31073 2891 31080
rect 1981 31047 2183 31073
rect 1981 31046 2020 31047
tri 2020 31046 2021 31047 nw
tri 2143 31046 2144 31047 ne
rect 2144 31046 2183 31047
rect 2217 31047 2419 31073
rect 2217 31046 2256 31047
tri 2256 31046 2257 31047 nw
tri 2379 31046 2380 31047 ne
rect 2380 31046 2419 31047
rect 2453 31047 2655 31073
rect 2453 31046 2492 31047
tri 2492 31046 2493 31047 nw
tri 2615 31046 2616 31047 ne
rect 2616 31046 2655 31047
rect 2689 31047 2891 31073
rect 2689 31046 2728 31047
tri 2728 31046 2729 31047 nw
tri 2851 31046 2852 31047 ne
rect 2852 31046 2891 31047
rect 2925 31046 3076 31080
rect 380 31042 600 31046
tri 600 31042 604 31046 nw
tri 728 31042 732 31046 ne
rect 732 31042 836 31046
tri 836 31042 840 31046 nw
tri 964 31042 968 31046 ne
rect 968 31042 1072 31046
tri 1072 31042 1076 31046 nw
tri 1200 31042 1204 31046 ne
rect 1204 31042 1308 31046
tri 1308 31042 1312 31046 nw
tri 1436 31042 1440 31046 ne
rect 1440 31042 1544 31046
tri 1544 31042 1548 31046 nw
tri 1672 31042 1676 31046 ne
rect 1676 31042 1780 31046
tri 1780 31042 1784 31046 nw
tri 1908 31042 1912 31046 ne
rect 1912 31042 2016 31046
tri 2016 31042 2020 31046 nw
tri 2144 31042 2148 31046 ne
rect 2148 31042 2252 31046
tri 2252 31042 2256 31046 nw
tri 2380 31042 2384 31046 ne
rect 2384 31042 2488 31046
tri 2488 31042 2492 31046 nw
tri 2616 31042 2620 31046 ne
rect 2620 31042 2724 31046
tri 2724 31042 2728 31046 nw
tri 2852 31042 2856 31046 ne
rect 2856 31042 3076 31046
rect 380 31023 571 31042
rect 380 30989 386 31023
rect 420 31006 571 31023
tri 571 31013 600 31042 nw
tri 732 31013 761 31042 ne
rect 420 30989 531 31006
rect 380 30972 531 30989
rect 565 30972 571 31006
rect 380 30951 571 30972
rect 380 30917 386 30951
rect 420 30932 571 30951
rect 420 30917 531 30932
rect 380 30898 531 30917
rect 565 30898 571 30932
rect 380 30879 571 30898
rect 380 30845 386 30879
rect 420 30858 571 30879
rect 420 30845 531 30858
rect 380 30824 531 30845
rect 565 30824 571 30858
rect 380 30807 571 30824
rect 380 30773 386 30807
rect 420 30784 571 30807
rect 420 30773 531 30784
rect 380 30750 531 30773
rect 565 30750 571 30784
rect 380 30735 571 30750
rect 380 30701 386 30735
rect 420 30710 571 30735
rect 420 30701 531 30710
rect 380 30676 531 30701
rect 565 30676 571 30710
rect 380 30663 571 30676
rect 380 30629 386 30663
rect 420 30636 571 30663
rect 420 30629 531 30636
rect 380 30602 531 30629
rect 565 30602 571 30636
rect 380 30591 571 30602
rect 380 30557 386 30591
rect 420 30557 571 30591
rect 761 31006 807 31042
tri 807 31013 836 31042 nw
tri 968 31013 997 31042 ne
rect 761 30972 767 31006
rect 801 30972 807 31006
rect 761 30932 807 30972
rect 761 30898 767 30932
rect 801 30898 807 30932
rect 761 30858 807 30898
rect 761 30824 767 30858
rect 801 30824 807 30858
rect 761 30784 807 30824
rect 761 30750 767 30784
rect 801 30750 807 30784
rect 761 30710 807 30750
rect 761 30676 767 30710
rect 801 30676 807 30710
rect 761 30636 807 30676
rect 761 30602 767 30636
rect 801 30602 807 30636
rect 761 30590 807 30602
rect 997 31006 1043 31042
tri 1043 31013 1072 31042 nw
tri 1204 31013 1233 31042 ne
rect 997 30972 1003 31006
rect 1037 30972 1043 31006
rect 997 30932 1043 30972
rect 997 30898 1003 30932
rect 1037 30898 1043 30932
rect 997 30858 1043 30898
rect 997 30824 1003 30858
rect 1037 30824 1043 30858
rect 997 30784 1043 30824
rect 997 30750 1003 30784
rect 1037 30750 1043 30784
rect 997 30710 1043 30750
rect 997 30676 1003 30710
rect 1037 30676 1043 30710
rect 997 30636 1043 30676
rect 997 30602 1003 30636
rect 1037 30602 1043 30636
rect 997 30590 1043 30602
rect 1233 31006 1279 31042
tri 1279 31013 1308 31042 nw
tri 1440 31013 1469 31042 ne
rect 1233 30972 1239 31006
rect 1273 30972 1279 31006
rect 1233 30932 1279 30972
rect 1233 30898 1239 30932
rect 1273 30898 1279 30932
rect 1233 30858 1279 30898
rect 1233 30824 1239 30858
rect 1273 30824 1279 30858
rect 1233 30784 1279 30824
rect 1233 30750 1239 30784
rect 1273 30750 1279 30784
rect 1233 30710 1279 30750
rect 1233 30676 1239 30710
rect 1273 30676 1279 30710
rect 1233 30636 1279 30676
rect 1233 30602 1239 30636
rect 1273 30602 1279 30636
rect 1233 30590 1279 30602
rect 1469 31006 1515 31042
tri 1515 31013 1544 31042 nw
tri 1676 31013 1705 31042 ne
rect 1469 30972 1475 31006
rect 1509 30972 1515 31006
rect 1469 30932 1515 30972
rect 1469 30898 1475 30932
rect 1509 30898 1515 30932
rect 1469 30858 1515 30898
rect 1469 30824 1475 30858
rect 1509 30824 1515 30858
rect 1469 30784 1515 30824
rect 1469 30750 1475 30784
rect 1509 30750 1515 30784
rect 1469 30710 1515 30750
rect 1469 30676 1475 30710
rect 1509 30676 1515 30710
rect 1469 30636 1515 30676
rect 1469 30602 1475 30636
rect 1509 30602 1515 30636
rect 1469 30590 1515 30602
rect 1705 31006 1751 31042
tri 1751 31013 1780 31042 nw
tri 1912 31013 1941 31042 ne
rect 1705 30972 1711 31006
rect 1745 30972 1751 31006
rect 1705 30932 1751 30972
rect 1705 30898 1711 30932
rect 1745 30898 1751 30932
rect 1705 30858 1751 30898
rect 1705 30824 1711 30858
rect 1745 30824 1751 30858
rect 1705 30784 1751 30824
rect 1705 30750 1711 30784
rect 1745 30750 1751 30784
rect 1705 30710 1751 30750
rect 1705 30676 1711 30710
rect 1745 30676 1751 30710
rect 1705 30636 1751 30676
rect 1705 30602 1711 30636
rect 1745 30602 1751 30636
rect 1705 30590 1751 30602
rect 1941 31006 1987 31042
tri 1987 31013 2016 31042 nw
tri 2148 31013 2177 31042 ne
rect 1941 30972 1947 31006
rect 1981 30972 1987 31006
rect 1941 30932 1987 30972
rect 1941 30898 1947 30932
rect 1981 30898 1987 30932
rect 1941 30858 1987 30898
rect 1941 30824 1947 30858
rect 1981 30824 1987 30858
rect 1941 30784 1987 30824
rect 1941 30750 1947 30784
rect 1981 30750 1987 30784
rect 1941 30710 1987 30750
rect 1941 30676 1947 30710
rect 1981 30676 1987 30710
rect 1941 30636 1987 30676
rect 1941 30602 1947 30636
rect 1981 30602 1987 30636
rect 1941 30590 1987 30602
rect 2177 31006 2223 31042
tri 2223 31013 2252 31042 nw
tri 2384 31013 2413 31042 ne
rect 2177 30972 2183 31006
rect 2217 30972 2223 31006
rect 2177 30932 2223 30972
rect 2177 30898 2183 30932
rect 2217 30898 2223 30932
rect 2177 30858 2223 30898
rect 2177 30824 2183 30858
rect 2217 30824 2223 30858
rect 2177 30784 2223 30824
rect 2177 30750 2183 30784
rect 2217 30750 2223 30784
rect 2177 30710 2223 30750
rect 2177 30676 2183 30710
rect 2217 30676 2223 30710
rect 2177 30636 2223 30676
rect 2177 30602 2183 30636
rect 2217 30602 2223 30636
rect 2177 30590 2223 30602
rect 2413 31006 2459 31042
tri 2459 31013 2488 31042 nw
tri 2620 31013 2649 31042 ne
rect 2413 30972 2419 31006
rect 2453 30972 2459 31006
rect 2413 30932 2459 30972
rect 2413 30898 2419 30932
rect 2453 30898 2459 30932
rect 2413 30858 2459 30898
rect 2413 30824 2419 30858
rect 2453 30824 2459 30858
rect 2413 30784 2459 30824
rect 2413 30750 2419 30784
rect 2453 30750 2459 30784
rect 2413 30710 2459 30750
rect 2413 30676 2419 30710
rect 2453 30676 2459 30710
rect 2413 30636 2459 30676
rect 2413 30602 2419 30636
rect 2453 30602 2459 30636
rect 2413 30590 2459 30602
rect 2649 31006 2695 31042
tri 2695 31013 2724 31042 nw
tri 2856 31013 2885 31042 ne
rect 2649 30972 2655 31006
rect 2689 30972 2695 31006
rect 2649 30932 2695 30972
rect 2649 30898 2655 30932
rect 2689 30898 2695 30932
rect 2649 30858 2695 30898
rect 2649 30824 2655 30858
rect 2689 30824 2695 30858
rect 2649 30784 2695 30824
rect 2649 30750 2655 30784
rect 2689 30750 2695 30784
rect 2649 30710 2695 30750
rect 2649 30676 2655 30710
rect 2689 30676 2695 30710
rect 2649 30636 2695 30676
rect 2649 30602 2655 30636
rect 2689 30602 2695 30636
rect 2649 30590 2695 30602
rect 2885 31008 3036 31042
rect 3070 31008 3076 31042
rect 2885 31006 3076 31008
rect 2885 30972 2891 31006
rect 2925 30972 3076 31006
rect 2885 30970 3076 30972
rect 2885 30936 3036 30970
rect 3070 30936 3076 30970
rect 2885 30932 3076 30936
rect 2885 30898 2891 30932
rect 2925 30898 3076 30932
rect 2885 30864 3036 30898
rect 3070 30864 3076 30898
rect 2885 30858 3076 30864
rect 2885 30824 2891 30858
rect 2925 30826 3076 30858
rect 2925 30824 3036 30826
rect 2885 30792 3036 30824
rect 3070 30792 3076 30826
rect 2885 30784 3076 30792
rect 2885 30750 2891 30784
rect 2925 30754 3076 30784
rect 2925 30750 3036 30754
rect 2885 30720 3036 30750
rect 3070 30720 3076 30754
rect 2885 30710 3076 30720
rect 2885 30676 2891 30710
rect 2925 30682 3076 30710
rect 2925 30676 3036 30682
rect 2885 30648 3036 30676
rect 3070 30648 3076 30682
rect 2885 30636 3076 30648
rect 2885 30602 2891 30636
rect 2925 30610 3076 30636
rect 2925 30602 3036 30610
rect 380 30519 571 30557
rect 2885 30576 3036 30602
rect 3070 30576 3076 30610
rect 380 30485 386 30519
rect 420 30485 571 30519
rect 613 30534 1501 30543
rect 1553 30534 1569 30543
rect 1621 30534 1636 30543
rect 1688 30534 1703 30543
rect 1755 30534 1770 30543
rect 1822 30534 1837 30543
rect 1889 30534 2830 30543
rect 613 30500 625 30534
rect 659 30500 700 30534
rect 734 30500 775 30534
rect 809 30500 850 30534
rect 884 30500 925 30534
rect 959 30500 1000 30534
rect 1034 30500 1075 30534
rect 1109 30500 1150 30534
rect 1184 30500 1225 30534
rect 1259 30500 1300 30534
rect 1334 30500 1375 30534
rect 1409 30500 1450 30534
rect 1484 30500 1501 30534
rect 1559 30500 1569 30534
rect 1634 30500 1636 30534
rect 1889 30500 1896 30534
rect 1930 30500 1970 30534
rect 2004 30500 2044 30534
rect 2078 30500 2118 30534
rect 2152 30500 2192 30534
rect 2226 30500 2266 30534
rect 2300 30500 2340 30534
rect 2374 30500 2414 30534
rect 2448 30500 2488 30534
rect 2522 30500 2562 30534
rect 2596 30500 2636 30534
rect 2670 30500 2710 30534
rect 2744 30500 2784 30534
rect 2818 30500 2830 30534
rect 613 30491 1501 30500
rect 1553 30491 1569 30500
rect 1621 30491 1636 30500
rect 1688 30491 1703 30500
rect 1755 30491 1770 30500
rect 1822 30491 1837 30500
rect 1889 30491 2830 30500
rect 2885 30538 3076 30576
rect 2885 30504 3036 30538
rect 3070 30504 3076 30538
rect 380 30447 571 30485
rect 380 30413 386 30447
rect 420 30432 571 30447
rect 2885 30466 3076 30504
rect 420 30413 531 30432
rect 380 30398 531 30413
rect 565 30398 571 30432
rect 380 30375 571 30398
rect 380 30341 386 30375
rect 420 30359 571 30375
rect 420 30341 531 30359
rect 380 30325 531 30341
rect 565 30325 571 30359
rect 380 30303 571 30325
rect 380 30269 386 30303
rect 420 30286 571 30303
rect 420 30269 531 30286
rect 380 30252 531 30269
rect 565 30252 571 30286
rect 380 30231 571 30252
rect 380 30197 386 30231
rect 420 30213 571 30231
rect 420 30197 531 30213
rect 380 30179 531 30197
rect 565 30179 571 30213
rect 380 30159 571 30179
rect 380 30125 386 30159
rect 420 30140 571 30159
rect 420 30125 531 30140
rect 380 30106 531 30125
rect 565 30106 571 30140
rect 380 30087 571 30106
rect 380 30053 386 30087
rect 420 30067 571 30087
rect 420 30053 531 30067
rect 380 30033 531 30053
rect 565 30033 571 30067
rect 380 30015 571 30033
rect 380 29981 386 30015
rect 420 29994 571 30015
rect 420 29981 531 29994
rect 380 29960 531 29981
rect 565 29960 571 29994
rect 380 29943 571 29960
rect 380 29909 386 29943
rect 420 29928 571 29943
rect 761 30432 807 30444
rect 761 30398 767 30432
rect 801 30398 807 30432
rect 761 30359 807 30398
rect 761 30325 767 30359
rect 801 30325 807 30359
rect 761 30286 807 30325
rect 761 30252 767 30286
rect 801 30252 807 30286
rect 761 30213 807 30252
rect 761 30179 767 30213
rect 801 30179 807 30213
rect 761 30140 807 30179
rect 761 30106 767 30140
rect 801 30106 807 30140
rect 761 30067 807 30106
rect 761 30033 767 30067
rect 801 30033 807 30067
rect 761 29994 807 30033
rect 761 29960 767 29994
rect 801 29960 807 29994
tri 571 29928 577 29934 sw
tri 755 29928 761 29934 se
rect 761 29928 807 29960
rect 997 30432 1043 30444
rect 997 30398 1003 30432
rect 1037 30398 1043 30432
rect 997 30359 1043 30398
rect 997 30325 1003 30359
rect 1037 30325 1043 30359
rect 997 30286 1043 30325
rect 997 30252 1003 30286
rect 1037 30252 1043 30286
rect 997 30213 1043 30252
rect 997 30179 1003 30213
rect 1037 30179 1043 30213
rect 997 30140 1043 30179
rect 997 30106 1003 30140
rect 1037 30106 1043 30140
rect 997 30067 1043 30106
rect 997 30033 1003 30067
rect 1037 30033 1043 30067
rect 997 29994 1043 30033
rect 997 29960 1003 29994
rect 1037 29960 1043 29994
tri 807 29928 813 29934 sw
tri 991 29928 997 29934 se
rect 997 29928 1043 29960
rect 1233 30432 1279 30444
rect 1233 30398 1239 30432
rect 1273 30398 1279 30432
rect 1233 30359 1279 30398
rect 1233 30325 1239 30359
rect 1273 30325 1279 30359
rect 1233 30286 1279 30325
rect 1233 30252 1239 30286
rect 1273 30252 1279 30286
rect 1233 30213 1279 30252
rect 1233 30179 1239 30213
rect 1273 30179 1279 30213
rect 1233 30140 1279 30179
rect 1233 30106 1239 30140
rect 1273 30106 1279 30140
rect 1233 30067 1279 30106
rect 1233 30033 1239 30067
rect 1273 30033 1279 30067
rect 1233 29994 1279 30033
rect 1233 29960 1239 29994
rect 1273 29960 1279 29994
tri 1043 29928 1049 29934 sw
tri 1227 29928 1233 29934 se
rect 1233 29928 1279 29960
rect 1469 30432 1515 30444
rect 1469 30398 1475 30432
rect 1509 30398 1515 30432
rect 1469 30359 1515 30398
rect 1469 30325 1475 30359
rect 1509 30325 1515 30359
rect 1469 30286 1515 30325
rect 1469 30252 1475 30286
rect 1509 30252 1515 30286
rect 1469 30213 1515 30252
rect 1469 30179 1475 30213
rect 1509 30179 1515 30213
rect 1469 30140 1515 30179
rect 1469 30106 1475 30140
rect 1509 30106 1515 30140
rect 1469 30067 1515 30106
rect 1469 30033 1475 30067
rect 1509 30033 1515 30067
rect 1469 29994 1515 30033
rect 1469 29960 1475 29994
rect 1509 29960 1515 29994
tri 1279 29928 1285 29934 sw
tri 1463 29928 1469 29934 se
rect 1469 29928 1515 29960
rect 1705 30432 1751 30444
rect 1705 30398 1711 30432
rect 1745 30398 1751 30432
rect 1705 30359 1751 30398
rect 1705 30325 1711 30359
rect 1745 30325 1751 30359
rect 1705 30286 1751 30325
rect 1705 30252 1711 30286
rect 1745 30252 1751 30286
rect 1705 30213 1751 30252
rect 1705 30179 1711 30213
rect 1745 30179 1751 30213
rect 1705 30140 1751 30179
rect 1705 30106 1711 30140
rect 1745 30106 1751 30140
rect 1705 30067 1751 30106
rect 1705 30033 1711 30067
rect 1745 30033 1751 30067
rect 1705 29994 1751 30033
rect 1705 29960 1711 29994
rect 1745 29960 1751 29994
tri 1515 29928 1521 29934 sw
tri 1699 29928 1705 29934 se
rect 1705 29928 1751 29960
rect 1941 30432 1987 30444
rect 1941 30398 1947 30432
rect 1981 30398 1987 30432
rect 1941 30359 1987 30398
rect 1941 30325 1947 30359
rect 1981 30325 1987 30359
rect 1941 30286 1987 30325
rect 1941 30252 1947 30286
rect 1981 30252 1987 30286
rect 1941 30213 1987 30252
rect 1941 30179 1947 30213
rect 1981 30179 1987 30213
rect 1941 30140 1987 30179
rect 1941 30106 1947 30140
rect 1981 30106 1987 30140
rect 1941 30067 1987 30106
rect 1941 30033 1947 30067
rect 1981 30033 1987 30067
rect 1941 29994 1987 30033
rect 1941 29960 1947 29994
rect 1981 29960 1987 29994
tri 1751 29928 1757 29934 sw
tri 1935 29928 1941 29934 se
rect 1941 29928 1987 29960
rect 2177 30432 2223 30444
rect 2177 30398 2183 30432
rect 2217 30398 2223 30432
rect 2177 30359 2223 30398
rect 2177 30325 2183 30359
rect 2217 30325 2223 30359
rect 2177 30286 2223 30325
rect 2177 30252 2183 30286
rect 2217 30252 2223 30286
rect 2177 30213 2223 30252
rect 2177 30179 2183 30213
rect 2217 30179 2223 30213
rect 2177 30140 2223 30179
rect 2177 30106 2183 30140
rect 2217 30106 2223 30140
rect 2177 30067 2223 30106
rect 2177 30033 2183 30067
rect 2217 30033 2223 30067
rect 2177 29994 2223 30033
rect 2177 29960 2183 29994
rect 2217 29960 2223 29994
tri 1987 29928 1993 29934 sw
tri 2171 29928 2177 29934 se
rect 2177 29928 2223 29960
rect 2413 30432 2459 30444
rect 2413 30398 2419 30432
rect 2453 30398 2459 30432
rect 2413 30359 2459 30398
rect 2413 30325 2419 30359
rect 2453 30325 2459 30359
rect 2413 30286 2459 30325
rect 2413 30252 2419 30286
rect 2453 30252 2459 30286
rect 2413 30213 2459 30252
rect 2413 30179 2419 30213
rect 2453 30179 2459 30213
rect 2413 30140 2459 30179
rect 2413 30106 2419 30140
rect 2453 30106 2459 30140
rect 2413 30067 2459 30106
rect 2413 30033 2419 30067
rect 2453 30033 2459 30067
rect 2413 29994 2459 30033
rect 2413 29960 2419 29994
rect 2453 29960 2459 29994
tri 2223 29928 2229 29934 sw
tri 2407 29928 2413 29934 se
rect 2413 29928 2459 29960
rect 2649 30432 2695 30444
rect 2649 30398 2655 30432
rect 2689 30398 2695 30432
rect 2649 30359 2695 30398
rect 2649 30325 2655 30359
rect 2689 30325 2695 30359
rect 2649 30286 2695 30325
rect 2649 30252 2655 30286
rect 2689 30252 2695 30286
rect 2649 30213 2695 30252
rect 2649 30179 2655 30213
rect 2689 30179 2695 30213
rect 2649 30140 2695 30179
rect 2649 30106 2655 30140
rect 2689 30106 2695 30140
rect 2649 30067 2695 30106
rect 2649 30033 2655 30067
rect 2689 30033 2695 30067
rect 2649 29994 2695 30033
rect 2649 29960 2655 29994
rect 2689 29960 2695 29994
tri 2459 29928 2465 29934 sw
tri 2643 29928 2649 29934 se
rect 2649 29928 2695 29960
rect 2885 30432 3036 30466
rect 3070 30432 3076 30466
rect 2885 30398 2891 30432
rect 2925 30398 3076 30432
rect 2885 30394 3076 30398
rect 2885 30360 3036 30394
rect 3070 30360 3076 30394
rect 2885 30359 3076 30360
rect 2885 30325 2891 30359
rect 2925 30325 3076 30359
rect 2885 30322 3076 30325
rect 2885 30288 3036 30322
rect 3070 30288 3076 30322
rect 2885 30286 3076 30288
rect 2885 30252 2891 30286
rect 2925 30252 3076 30286
rect 2885 30250 3076 30252
rect 2885 30216 3036 30250
rect 3070 30216 3076 30250
rect 2885 30213 3076 30216
rect 2885 30179 2891 30213
rect 2925 30179 3076 30213
rect 2885 30178 3076 30179
rect 2885 30144 3036 30178
rect 3070 30144 3076 30178
rect 2885 30140 3076 30144
rect 2885 30106 2891 30140
rect 2925 30106 3076 30140
rect 2885 30072 3036 30106
rect 3070 30072 3076 30106
rect 2885 30067 3076 30072
rect 2885 30033 2891 30067
rect 2925 30034 3076 30067
rect 2925 30033 3036 30034
rect 2885 30000 3036 30033
rect 3070 30000 3076 30034
rect 2885 29994 3076 30000
rect 2885 29960 2891 29994
rect 2925 29962 3076 29994
rect 2925 29960 3036 29962
tri 2695 29928 2701 29934 sw
tri 2879 29928 2885 29934 se
rect 2885 29928 3036 29960
rect 3070 29928 3076 29962
rect 420 29921 577 29928
tri 577 29921 584 29928 sw
tri 748 29921 755 29928 se
rect 755 29921 813 29928
tri 813 29921 820 29928 sw
tri 984 29921 991 29928 se
rect 991 29921 1049 29928
tri 1049 29921 1056 29928 sw
tri 1220 29921 1227 29928 se
rect 1227 29921 1285 29928
tri 1285 29921 1292 29928 sw
tri 1456 29921 1463 29928 se
rect 1463 29921 1521 29928
tri 1521 29921 1528 29928 sw
tri 1692 29921 1699 29928 se
rect 1699 29921 1757 29928
tri 1757 29921 1764 29928 sw
tri 1928 29921 1935 29928 se
rect 1935 29921 1993 29928
tri 1993 29921 2000 29928 sw
tri 2164 29921 2171 29928 se
rect 2171 29921 2229 29928
tri 2229 29921 2236 29928 sw
tri 2400 29921 2407 29928 se
rect 2407 29921 2465 29928
tri 2465 29921 2472 29928 sw
tri 2636 29921 2643 29928 se
rect 2643 29921 2701 29928
tri 2701 29921 2708 29928 sw
tri 2872 29921 2879 29928 se
rect 2879 29921 3076 29928
rect 420 29909 531 29921
rect 380 29887 531 29909
rect 565 29900 584 29921
tri 584 29900 605 29921 sw
tri 727 29900 748 29921 se
rect 748 29900 767 29921
rect 565 29887 767 29900
rect 801 29900 820 29921
tri 820 29900 841 29921 sw
tri 963 29900 984 29921 se
rect 984 29900 1003 29921
rect 801 29887 1003 29900
rect 1037 29900 1056 29921
tri 1056 29900 1077 29921 sw
tri 1199 29900 1220 29921 se
rect 1220 29900 1239 29921
rect 1037 29887 1239 29900
rect 1273 29900 1292 29921
tri 1292 29900 1313 29921 sw
tri 1435 29900 1456 29921 se
rect 1456 29900 1475 29921
rect 1273 29887 1475 29900
rect 1509 29900 1528 29921
tri 1528 29900 1549 29921 sw
tri 1671 29900 1692 29921 se
rect 1692 29900 1711 29921
rect 1509 29887 1711 29900
rect 1745 29900 1764 29921
tri 1764 29900 1785 29921 sw
tri 1907 29900 1928 29921 se
rect 1928 29900 1947 29921
rect 1745 29887 1947 29900
rect 1981 29900 2000 29921
tri 2000 29900 2021 29921 sw
tri 2143 29900 2164 29921 se
rect 2164 29900 2183 29921
rect 1981 29887 2183 29900
rect 2217 29900 2236 29921
tri 2236 29900 2257 29921 sw
tri 2379 29900 2400 29921 se
rect 2400 29900 2419 29921
rect 2217 29887 2419 29900
rect 2453 29900 2472 29921
tri 2472 29900 2493 29921 sw
tri 2615 29900 2636 29921 se
rect 2636 29900 2655 29921
rect 2453 29887 2655 29900
rect 2689 29900 2708 29921
tri 2708 29900 2729 29921 sw
tri 2851 29900 2872 29921 se
rect 2872 29900 2891 29921
rect 2689 29887 2891 29900
rect 2925 29890 3076 29921
rect 2925 29887 3036 29890
rect 380 29872 3036 29887
rect 380 29871 697 29872
rect 380 29837 386 29871
rect 420 29848 697 29871
rect 420 29837 531 29848
rect 380 29814 531 29837
rect 565 29820 697 29848
rect 749 29820 765 29872
rect 817 29820 833 29872
rect 885 29820 901 29872
rect 953 29820 969 29872
rect 1021 29848 1037 29872
rect 1089 29820 1105 29872
rect 1157 29820 1173 29872
rect 1225 29848 1241 29872
rect 1293 29848 2097 29872
rect 1225 29820 1239 29848
rect 1293 29820 1475 29848
rect 565 29814 767 29820
rect 801 29814 1003 29820
rect 1037 29814 1239 29820
rect 1273 29814 1475 29820
rect 1509 29814 1711 29848
rect 1745 29814 1947 29848
rect 1981 29820 2097 29848
rect 2149 29820 2165 29872
rect 2217 29820 2233 29872
rect 2285 29820 2301 29872
rect 2353 29820 2369 29872
rect 2421 29848 2437 29872
rect 2489 29820 2505 29872
rect 2557 29820 2573 29872
rect 2625 29820 2641 29872
rect 2693 29856 3036 29872
rect 3070 29856 3076 29890
rect 2693 29848 3076 29856
rect 2693 29820 2891 29848
rect 1981 29814 2183 29820
rect 2217 29814 2419 29820
rect 2453 29814 2655 29820
rect 2689 29814 2891 29820
rect 2925 29818 3076 29848
rect 2925 29814 3036 29818
rect 380 29808 3036 29814
rect 380 29799 697 29808
rect 380 29765 386 29799
rect 420 29775 697 29799
rect 420 29765 531 29775
rect 380 29741 531 29765
rect 565 29756 697 29775
rect 749 29756 765 29808
rect 817 29756 833 29808
rect 885 29756 901 29808
rect 953 29756 969 29808
rect 1021 29775 1037 29808
rect 1089 29756 1105 29808
rect 1157 29756 1173 29808
rect 1225 29775 1241 29808
rect 1293 29775 2097 29808
rect 1225 29756 1239 29775
rect 1293 29756 1475 29775
rect 565 29744 767 29756
rect 801 29744 1003 29756
rect 1037 29744 1239 29756
rect 1273 29744 1475 29756
rect 565 29741 697 29744
rect 380 29727 697 29741
rect 380 29693 386 29727
rect 420 29702 697 29727
rect 420 29693 531 29702
rect 380 29668 531 29693
rect 565 29692 697 29702
rect 749 29692 765 29744
rect 817 29692 833 29744
rect 885 29692 901 29744
rect 953 29692 969 29744
rect 1021 29702 1037 29741
rect 1089 29692 1105 29744
rect 1157 29692 1173 29744
rect 1225 29741 1239 29744
rect 1293 29741 1475 29744
rect 1509 29741 1711 29775
rect 1745 29741 1947 29775
rect 1981 29756 2097 29775
rect 2149 29756 2165 29808
rect 2217 29756 2233 29808
rect 2285 29756 2301 29808
rect 2353 29756 2369 29808
rect 2421 29775 2437 29808
rect 2489 29756 2505 29808
rect 2557 29756 2573 29808
rect 2625 29756 2641 29808
rect 2693 29784 3036 29808
rect 3070 29784 3076 29818
rect 2693 29775 3076 29784
rect 2693 29756 2891 29775
rect 1981 29744 2183 29756
rect 2217 29744 2419 29756
rect 2453 29744 2655 29756
rect 2689 29744 2891 29756
rect 1981 29741 2097 29744
rect 1225 29702 1241 29741
rect 1293 29702 2097 29741
rect 1225 29692 1239 29702
rect 1293 29692 1475 29702
rect 565 29680 767 29692
rect 801 29680 1003 29692
rect 1037 29680 1239 29692
rect 1273 29680 1475 29692
rect 565 29668 697 29680
rect 380 29655 697 29668
rect 380 29621 386 29655
rect 420 29629 697 29655
rect 420 29621 531 29629
rect 380 29595 531 29621
rect 565 29628 697 29629
rect 749 29628 765 29680
rect 817 29628 833 29680
rect 885 29628 901 29680
rect 953 29628 969 29680
rect 1021 29629 1037 29668
rect 1089 29628 1105 29680
rect 1157 29628 1173 29680
rect 1225 29668 1239 29680
rect 1293 29668 1475 29680
rect 1509 29668 1711 29702
rect 1745 29668 1947 29702
rect 1981 29692 2097 29702
rect 2149 29692 2165 29744
rect 2217 29692 2233 29744
rect 2285 29692 2301 29744
rect 2353 29692 2369 29744
rect 2421 29702 2437 29741
rect 2489 29692 2505 29744
rect 2557 29692 2573 29744
rect 2625 29692 2641 29744
rect 2693 29741 2891 29744
rect 2925 29746 3076 29775
rect 2925 29741 3036 29746
rect 2693 29712 3036 29741
rect 3070 29712 3076 29746
rect 2693 29702 3076 29712
rect 2693 29692 2891 29702
rect 1981 29680 2183 29692
rect 2217 29680 2419 29692
rect 2453 29680 2655 29692
rect 2689 29680 2891 29692
rect 1981 29668 2097 29680
rect 1225 29629 1241 29668
rect 1293 29629 2097 29668
rect 1225 29628 1239 29629
rect 1293 29628 1475 29629
rect 565 29616 767 29628
rect 801 29616 1003 29628
rect 1037 29616 1239 29628
rect 1273 29616 1475 29628
rect 565 29595 697 29616
rect 380 29583 697 29595
rect 380 29549 386 29583
rect 420 29564 697 29583
rect 749 29564 765 29616
rect 817 29564 833 29616
rect 885 29564 901 29616
rect 953 29564 969 29616
rect 1021 29564 1037 29595
rect 1089 29564 1105 29616
rect 1157 29564 1173 29616
rect 1225 29595 1239 29616
rect 1293 29595 1475 29616
rect 1509 29595 1711 29629
rect 1745 29595 1947 29629
rect 1981 29628 2097 29629
rect 2149 29628 2165 29680
rect 2217 29628 2233 29680
rect 2285 29628 2301 29680
rect 2353 29628 2369 29680
rect 2421 29629 2437 29668
rect 2489 29628 2505 29680
rect 2557 29628 2573 29680
rect 2625 29628 2641 29680
rect 2693 29668 2891 29680
rect 2925 29674 3076 29702
rect 2925 29668 3036 29674
rect 2693 29640 3036 29668
rect 3070 29640 3076 29674
rect 2693 29629 3076 29640
rect 2693 29628 2891 29629
rect 1981 29616 2183 29628
rect 2217 29616 2419 29628
rect 2453 29616 2655 29628
rect 2689 29616 2891 29628
rect 1981 29595 2097 29616
rect 1225 29564 1241 29595
rect 1293 29564 2097 29595
rect 2149 29564 2165 29616
rect 2217 29564 2233 29616
rect 2285 29564 2301 29616
rect 2353 29564 2369 29616
rect 2421 29564 2437 29595
rect 2489 29564 2505 29616
rect 2557 29564 2573 29616
rect 2625 29564 2641 29616
rect 2693 29595 2891 29616
rect 2925 29602 3076 29629
rect 2925 29595 3036 29602
rect 2693 29568 3036 29595
rect 3070 29568 3076 29602
rect 2693 29564 3076 29568
rect 420 29556 3076 29564
rect 420 29549 531 29556
rect 380 29522 531 29549
rect 565 29552 767 29556
rect 801 29552 1003 29556
rect 1037 29552 1239 29556
rect 1273 29552 1475 29556
rect 565 29522 697 29552
rect 380 29511 697 29522
rect 380 29477 386 29511
rect 420 29500 697 29511
rect 749 29500 765 29552
rect 817 29500 833 29552
rect 885 29500 901 29552
rect 953 29500 969 29552
rect 1021 29500 1037 29522
rect 1089 29500 1105 29552
rect 1157 29500 1173 29552
rect 1225 29522 1239 29552
rect 1293 29522 1475 29552
rect 1509 29522 1711 29556
rect 1745 29522 1947 29556
rect 1981 29552 2183 29556
rect 2217 29552 2419 29556
rect 2453 29552 2655 29556
rect 2689 29552 2891 29556
rect 1981 29522 2097 29552
rect 1225 29500 1241 29522
rect 1293 29500 2097 29522
rect 2149 29500 2165 29552
rect 2217 29500 2233 29552
rect 2285 29500 2301 29552
rect 2353 29500 2369 29552
rect 2421 29500 2437 29522
rect 2489 29500 2505 29552
rect 2557 29500 2573 29552
rect 2625 29500 2641 29552
rect 2693 29522 2891 29552
rect 2925 29530 3076 29556
rect 2925 29522 3036 29530
rect 2693 29500 3036 29522
rect 420 29496 3036 29500
rect 3070 29496 3076 29530
rect 420 29488 3076 29496
rect 420 29482 697 29488
rect 420 29477 531 29482
rect 380 29448 531 29477
rect 565 29448 697 29482
rect 380 29439 697 29448
rect 380 29405 386 29439
rect 420 29436 697 29439
rect 749 29436 765 29488
rect 817 29436 833 29488
rect 885 29436 901 29488
rect 953 29436 969 29488
rect 1021 29482 1037 29488
rect 1021 29436 1037 29448
rect 1089 29436 1105 29488
rect 1157 29436 1173 29488
rect 1225 29482 1241 29488
rect 1293 29482 2097 29488
rect 1225 29448 1239 29482
rect 1293 29448 1475 29482
rect 1509 29448 1711 29482
rect 1745 29448 1947 29482
rect 1981 29448 2097 29482
rect 1225 29436 1241 29448
rect 1293 29436 2097 29448
rect 2149 29436 2165 29488
rect 2217 29436 2233 29488
rect 2285 29436 2301 29488
rect 2353 29436 2369 29488
rect 2421 29482 2437 29488
rect 2421 29436 2437 29448
rect 2489 29436 2505 29488
rect 2557 29436 2573 29488
rect 2625 29436 2641 29488
rect 2693 29482 3076 29488
rect 2693 29448 2891 29482
rect 2925 29458 3076 29482
rect 2925 29448 3036 29458
rect 2693 29436 3036 29448
rect 420 29424 3036 29436
rect 3070 29424 3076 29458
rect 420 29408 697 29424
rect 420 29405 531 29408
rect 380 29374 531 29405
rect 565 29374 697 29408
rect 380 29372 697 29374
rect 749 29372 765 29424
rect 817 29372 833 29424
rect 885 29372 901 29424
rect 953 29372 969 29424
rect 1021 29408 1037 29424
rect 1021 29372 1037 29374
rect 1089 29372 1105 29424
rect 1157 29372 1173 29424
rect 1225 29408 1241 29424
rect 1293 29408 2097 29424
rect 1225 29374 1239 29408
rect 1293 29374 1475 29408
rect 1509 29374 1711 29408
rect 1745 29374 1947 29408
rect 1981 29374 2097 29408
rect 1225 29372 1241 29374
rect 1293 29372 2097 29374
rect 2149 29372 2165 29424
rect 2217 29372 2233 29424
rect 2285 29372 2301 29424
rect 2353 29372 2369 29424
rect 2421 29408 2437 29424
rect 2421 29372 2437 29374
rect 2489 29372 2505 29424
rect 2557 29372 2573 29424
rect 2625 29372 2641 29424
rect 2693 29408 3076 29424
rect 2693 29374 2891 29408
rect 2925 29386 3076 29408
rect 2925 29374 3036 29386
rect 2693 29372 3036 29374
rect 380 29367 3036 29372
rect 380 29333 386 29367
rect 420 29360 3036 29367
rect 420 29334 697 29360
rect 420 29333 531 29334
rect 380 29300 531 29333
rect 565 29308 697 29334
rect 749 29308 765 29360
rect 817 29308 833 29360
rect 885 29308 901 29360
rect 953 29308 969 29360
rect 1021 29334 1037 29360
rect 1089 29308 1105 29360
rect 1157 29308 1173 29360
rect 1225 29334 1241 29360
rect 1293 29334 2097 29360
rect 1225 29308 1239 29334
rect 1293 29308 1475 29334
rect 565 29300 767 29308
rect 801 29300 1003 29308
rect 1037 29300 1239 29308
rect 1273 29300 1475 29308
rect 1509 29300 1711 29334
rect 1745 29300 1947 29334
rect 1981 29308 2097 29334
rect 2149 29308 2165 29360
rect 2217 29308 2233 29360
rect 2285 29308 2301 29360
rect 2353 29308 2369 29360
rect 2421 29334 2437 29360
rect 2489 29308 2505 29360
rect 2557 29308 2573 29360
rect 2625 29308 2641 29360
rect 2693 29352 3036 29360
rect 3070 29352 3076 29386
rect 2693 29334 3076 29352
rect 2693 29308 2891 29334
rect 1981 29300 2183 29308
rect 2217 29300 2419 29308
rect 2453 29300 2655 29308
rect 2689 29300 2891 29308
rect 2925 29314 3076 29334
rect 2925 29300 3036 29314
rect 380 29296 3036 29300
rect 380 29295 697 29296
rect 380 29261 386 29295
rect 420 29261 697 29295
rect 380 29260 697 29261
rect 380 29226 531 29260
rect 565 29244 697 29260
rect 749 29244 765 29296
rect 817 29244 833 29296
rect 885 29244 901 29296
rect 953 29244 969 29296
rect 1021 29260 1037 29296
rect 1089 29244 1105 29296
rect 1157 29244 1173 29296
rect 1225 29260 1241 29296
rect 1293 29260 2097 29296
rect 1225 29244 1239 29260
rect 1293 29244 1475 29260
rect 565 29232 767 29244
rect 801 29232 1003 29244
rect 1037 29232 1239 29244
rect 1273 29232 1475 29244
rect 565 29226 697 29232
rect 380 29223 697 29226
rect 380 29189 386 29223
rect 420 29189 697 29223
rect 380 29186 697 29189
rect 380 29152 531 29186
rect 565 29180 697 29186
rect 749 29180 765 29232
rect 817 29180 833 29232
rect 885 29180 901 29232
rect 953 29180 969 29232
rect 1021 29186 1037 29226
rect 1089 29180 1105 29232
rect 1157 29180 1173 29232
rect 1225 29226 1239 29232
rect 1293 29226 1475 29232
rect 1509 29226 1711 29260
rect 1745 29226 1947 29260
rect 1981 29244 2097 29260
rect 2149 29244 2165 29296
rect 2217 29244 2233 29296
rect 2285 29244 2301 29296
rect 2353 29244 2369 29296
rect 2421 29260 2437 29296
rect 2489 29244 2505 29296
rect 2557 29244 2573 29296
rect 2625 29244 2641 29296
rect 2693 29280 3036 29296
rect 3070 29280 3076 29314
rect 2693 29260 3076 29280
rect 2693 29244 2891 29260
rect 1981 29232 2183 29244
rect 2217 29232 2419 29244
rect 2453 29232 2655 29244
rect 2689 29232 2891 29244
rect 1981 29226 2097 29232
rect 1225 29186 1241 29226
rect 1293 29186 2097 29226
rect 1225 29180 1239 29186
rect 1293 29180 1475 29186
rect 565 29168 767 29180
rect 801 29168 1003 29180
rect 1037 29168 1239 29180
rect 1273 29168 1475 29180
rect 565 29152 697 29168
rect 380 29151 697 29152
rect 380 29117 386 29151
rect 420 29117 697 29151
rect 380 29116 697 29117
rect 749 29116 765 29168
rect 817 29116 833 29168
rect 885 29116 901 29168
rect 953 29116 969 29168
rect 1021 29116 1037 29152
rect 1089 29116 1105 29168
rect 1157 29116 1173 29168
rect 1225 29152 1239 29168
rect 1293 29152 1475 29168
rect 1509 29152 1711 29186
rect 1745 29152 1947 29186
rect 1981 29180 2097 29186
rect 2149 29180 2165 29232
rect 2217 29180 2233 29232
rect 2285 29180 2301 29232
rect 2353 29180 2369 29232
rect 2421 29186 2437 29226
rect 2489 29180 2505 29232
rect 2557 29180 2573 29232
rect 2625 29180 2641 29232
rect 2693 29226 2891 29232
rect 2925 29242 3076 29260
rect 2925 29226 3036 29242
rect 2693 29208 3036 29226
rect 3070 29208 3076 29242
rect 2693 29186 3076 29208
rect 2693 29180 2891 29186
rect 1981 29168 2183 29180
rect 2217 29168 2419 29180
rect 2453 29168 2655 29180
rect 2689 29168 2891 29180
rect 1981 29152 2097 29168
rect 1225 29116 1241 29152
rect 1293 29116 2097 29152
rect 2149 29116 2165 29168
rect 2217 29116 2233 29168
rect 2285 29116 2301 29168
rect 2353 29116 2369 29168
rect 2421 29116 2437 29152
rect 2489 29116 2505 29168
rect 2557 29116 2573 29168
rect 2625 29116 2641 29168
rect 2693 29152 2891 29168
rect 2925 29170 3076 29186
rect 2925 29152 3036 29170
rect 2693 29136 3036 29152
rect 3070 29136 3076 29170
rect 2693 29116 3076 29136
rect 380 29112 3076 29116
rect 380 29079 531 29112
rect 380 29045 386 29079
rect 420 29078 531 29079
rect 565 29104 767 29112
rect 801 29104 1003 29112
rect 1037 29104 1239 29112
rect 1273 29104 1475 29112
rect 565 29078 697 29104
rect 420 29052 697 29078
rect 749 29052 765 29104
rect 817 29052 833 29104
rect 885 29052 901 29104
rect 953 29052 969 29104
rect 1021 29052 1037 29078
rect 1089 29052 1105 29104
rect 1157 29052 1173 29104
rect 1225 29078 1239 29104
rect 1293 29078 1475 29104
rect 1509 29078 1711 29112
rect 1745 29078 1947 29112
rect 1981 29104 2183 29112
rect 2217 29104 2419 29112
rect 2453 29104 2655 29112
rect 2689 29104 2891 29112
rect 1981 29078 2097 29104
rect 1225 29052 1241 29078
rect 1293 29052 2097 29078
rect 2149 29052 2165 29104
rect 2217 29052 2233 29104
rect 2285 29052 2301 29104
rect 2353 29052 2369 29104
rect 2421 29052 2437 29078
rect 2489 29052 2505 29104
rect 2557 29052 2573 29104
rect 2625 29052 2641 29104
rect 2693 29078 2891 29104
rect 2925 29098 3076 29112
rect 2925 29078 3036 29098
rect 2693 29064 3036 29078
rect 3070 29064 3076 29098
rect 2693 29052 3076 29064
rect 420 29045 3076 29052
rect 380 29040 3076 29045
rect 380 29038 697 29040
rect 380 29007 531 29038
rect 380 28973 386 29007
rect 420 29004 531 29007
rect 565 29004 697 29038
rect 420 28988 697 29004
rect 749 28988 765 29040
rect 817 28988 833 29040
rect 885 28988 901 29040
rect 953 28988 969 29040
rect 1021 29038 1037 29040
rect 1021 28988 1037 29004
rect 1089 28988 1105 29040
rect 1157 28988 1173 29040
rect 1225 29038 1241 29040
rect 1293 29038 2097 29040
rect 1225 29004 1239 29038
rect 1293 29004 1475 29038
rect 1509 29004 1711 29038
rect 1745 29004 1947 29038
rect 1981 29004 2097 29038
rect 1225 28988 1241 29004
rect 1293 28988 2097 29004
rect 2149 28988 2165 29040
rect 2217 28988 2233 29040
rect 2285 28988 2301 29040
rect 2353 28988 2369 29040
rect 2421 29038 2437 29040
rect 2421 28988 2437 29004
rect 2489 28988 2505 29040
rect 2557 28988 2573 29040
rect 2625 28988 2641 29040
rect 2693 29038 3076 29040
rect 2693 29004 2891 29038
rect 2925 29026 3076 29038
rect 2925 29004 3036 29026
rect 2693 28992 3036 29004
rect 3070 28992 3076 29026
rect 2693 28988 3076 28992
rect 420 28976 3076 28988
rect 420 28973 697 28976
rect 380 28964 697 28973
rect 380 28935 531 28964
rect 380 28901 386 28935
rect 420 28930 531 28935
rect 565 28930 697 28964
rect 420 28924 697 28930
rect 749 28924 765 28976
rect 817 28924 833 28976
rect 885 28924 901 28976
rect 953 28924 969 28976
rect 1021 28964 1037 28976
rect 1021 28924 1037 28930
rect 1089 28924 1105 28976
rect 1157 28924 1173 28976
rect 1225 28964 1241 28976
rect 1293 28964 2097 28976
rect 1225 28930 1239 28964
rect 1293 28930 1475 28964
rect 1509 28930 1711 28964
rect 1745 28930 1947 28964
rect 1981 28930 2097 28964
rect 1225 28924 1241 28930
rect 1293 28924 2097 28930
rect 2149 28924 2165 28976
rect 2217 28924 2233 28976
rect 2285 28924 2301 28976
rect 2353 28924 2369 28976
rect 2421 28964 2437 28976
rect 2421 28924 2437 28930
rect 2489 28924 2505 28976
rect 2557 28924 2573 28976
rect 2625 28924 2641 28976
rect 2693 28964 3076 28976
rect 2693 28930 2891 28964
rect 2925 28954 3076 28964
rect 2925 28930 3036 28954
rect 2693 28924 3036 28930
rect 420 28920 3036 28924
rect 3070 28920 3076 28954
rect 420 28901 3076 28920
rect 380 28900 3076 28901
rect 380 28896 601 28900
tri 601 28896 605 28900 nw
tri 727 28896 731 28900 ne
rect 731 28896 837 28900
tri 837 28896 841 28900 nw
tri 963 28896 967 28900 ne
rect 967 28896 1073 28900
tri 1073 28896 1077 28900 nw
tri 1199 28896 1203 28900 ne
rect 1203 28896 1309 28900
tri 1309 28896 1313 28900 nw
tri 1435 28896 1439 28900 ne
rect 1439 28896 1545 28900
tri 1545 28896 1549 28900 nw
tri 1671 28896 1675 28900 ne
rect 1675 28896 1781 28900
tri 1781 28896 1785 28900 nw
tri 1907 28896 1911 28900 ne
rect 1911 28896 2017 28900
tri 2017 28896 2021 28900 nw
tri 2143 28896 2147 28900 ne
rect 2147 28896 2253 28900
tri 2253 28896 2257 28900 nw
tri 2379 28896 2383 28900 ne
rect 2383 28896 2489 28900
tri 2489 28896 2493 28900 nw
tri 2615 28896 2619 28900 ne
rect 2619 28896 2725 28900
tri 2725 28896 2729 28900 nw
tri 2851 28896 2855 28900 ne
rect 2855 28896 3076 28900
rect 380 28890 595 28896
tri 595 28890 601 28896 nw
tri 731 28890 737 28896 ne
rect 737 28890 831 28896
tri 831 28890 837 28896 nw
tri 967 28890 973 28896 ne
rect 973 28890 1067 28896
tri 1067 28890 1073 28896 nw
tri 1203 28890 1209 28896 ne
rect 1209 28890 1303 28896
tri 1303 28890 1309 28896 nw
tri 1439 28890 1445 28896 ne
rect 1445 28890 1539 28896
tri 1539 28890 1545 28896 nw
tri 1675 28890 1681 28896 ne
rect 1681 28890 1775 28896
tri 1775 28890 1781 28896 nw
tri 1911 28890 1917 28896 ne
rect 1917 28890 2011 28896
tri 2011 28890 2017 28896 nw
tri 2147 28890 2153 28896 ne
rect 2153 28890 2247 28896
tri 2247 28890 2253 28896 nw
tri 2383 28890 2389 28896 ne
rect 2389 28890 2483 28896
tri 2483 28890 2489 28896 nw
tri 2619 28890 2625 28896 ne
rect 2625 28890 2719 28896
tri 2719 28890 2725 28896 nw
tri 2855 28890 2861 28896 ne
rect 2861 28890 3076 28896
rect 380 28863 531 28890
rect 380 28829 386 28863
rect 420 28856 531 28863
rect 565 28856 571 28890
tri 571 28866 595 28890 nw
tri 737 28866 761 28890 ne
rect 420 28829 571 28856
rect 380 28816 571 28829
rect 380 28791 531 28816
rect 380 28757 386 28791
rect 420 28782 531 28791
rect 565 28782 571 28816
rect 420 28757 571 28782
rect 380 28742 571 28757
rect 380 28719 531 28742
rect 380 28685 386 28719
rect 420 28708 531 28719
rect 565 28708 571 28742
rect 420 28685 571 28708
rect 380 28668 571 28685
rect 380 28647 531 28668
rect 380 28613 386 28647
rect 420 28634 531 28647
rect 565 28634 571 28668
rect 420 28613 571 28634
rect 380 28594 571 28613
rect 380 28575 531 28594
rect 380 28541 386 28575
rect 420 28560 531 28575
rect 565 28560 571 28594
rect 420 28541 571 28560
rect 380 28520 571 28541
rect 380 28503 531 28520
rect 380 28469 386 28503
rect 420 28486 531 28503
rect 565 28486 571 28520
rect 420 28469 571 28486
rect 761 28856 767 28890
rect 801 28856 807 28890
tri 807 28866 831 28890 nw
tri 973 28866 997 28890 ne
rect 761 28816 807 28856
rect 761 28782 767 28816
rect 801 28782 807 28816
rect 761 28742 807 28782
rect 761 28708 767 28742
rect 801 28708 807 28742
rect 761 28668 807 28708
rect 761 28634 767 28668
rect 801 28634 807 28668
rect 761 28594 807 28634
rect 761 28560 767 28594
rect 801 28560 807 28594
rect 761 28520 807 28560
rect 761 28486 767 28520
rect 801 28486 807 28520
rect 761 28474 807 28486
rect 997 28856 1003 28890
rect 1037 28856 1043 28890
tri 1043 28866 1067 28890 nw
tri 1209 28866 1233 28890 ne
rect 997 28816 1043 28856
rect 997 28782 1003 28816
rect 1037 28782 1043 28816
rect 997 28742 1043 28782
rect 997 28708 1003 28742
rect 1037 28708 1043 28742
rect 997 28668 1043 28708
rect 997 28634 1003 28668
rect 1037 28634 1043 28668
rect 997 28594 1043 28634
rect 997 28560 1003 28594
rect 1037 28560 1043 28594
rect 997 28520 1043 28560
rect 997 28486 1003 28520
rect 1037 28486 1043 28520
rect 997 28474 1043 28486
rect 1233 28856 1239 28890
rect 1273 28856 1279 28890
tri 1279 28866 1303 28890 nw
tri 1445 28866 1469 28890 ne
rect 1233 28816 1279 28856
rect 1233 28782 1239 28816
rect 1273 28782 1279 28816
rect 1233 28742 1279 28782
rect 1233 28708 1239 28742
rect 1273 28708 1279 28742
rect 1233 28668 1279 28708
rect 1233 28634 1239 28668
rect 1273 28634 1279 28668
rect 1233 28594 1279 28634
rect 1233 28560 1239 28594
rect 1273 28560 1279 28594
rect 1233 28520 1279 28560
rect 1233 28486 1239 28520
rect 1273 28486 1279 28520
rect 1233 28474 1279 28486
rect 1469 28856 1475 28890
rect 1509 28856 1515 28890
tri 1515 28866 1539 28890 nw
tri 1681 28866 1705 28890 ne
rect 1469 28816 1515 28856
rect 1469 28782 1475 28816
rect 1509 28782 1515 28816
rect 1469 28742 1515 28782
rect 1469 28708 1475 28742
rect 1509 28708 1515 28742
rect 1469 28668 1515 28708
rect 1469 28634 1475 28668
rect 1509 28634 1515 28668
rect 1469 28594 1515 28634
rect 1469 28560 1475 28594
rect 1509 28560 1515 28594
rect 1469 28520 1515 28560
rect 1469 28486 1475 28520
rect 1509 28486 1515 28520
rect 1469 28474 1515 28486
rect 1705 28856 1711 28890
rect 1745 28856 1751 28890
tri 1751 28866 1775 28890 nw
tri 1917 28866 1941 28890 ne
rect 1705 28816 1751 28856
rect 1705 28782 1711 28816
rect 1745 28782 1751 28816
rect 1705 28742 1751 28782
rect 1705 28708 1711 28742
rect 1745 28708 1751 28742
rect 1705 28668 1751 28708
rect 1705 28634 1711 28668
rect 1745 28634 1751 28668
rect 1705 28594 1751 28634
rect 1705 28560 1711 28594
rect 1745 28560 1751 28594
rect 1705 28520 1751 28560
rect 1705 28486 1711 28520
rect 1745 28486 1751 28520
rect 1705 28474 1751 28486
rect 1941 28856 1947 28890
rect 1981 28856 1987 28890
tri 1987 28866 2011 28890 nw
tri 2153 28866 2177 28890 ne
rect 1941 28816 1987 28856
rect 1941 28782 1947 28816
rect 1981 28782 1987 28816
rect 1941 28742 1987 28782
rect 1941 28708 1947 28742
rect 1981 28708 1987 28742
rect 1941 28668 1987 28708
rect 1941 28634 1947 28668
rect 1981 28634 1987 28668
rect 1941 28594 1987 28634
rect 1941 28560 1947 28594
rect 1981 28560 1987 28594
rect 1941 28520 1987 28560
rect 1941 28486 1947 28520
rect 1981 28486 1987 28520
rect 1941 28474 1987 28486
rect 2177 28856 2183 28890
rect 2217 28856 2223 28890
tri 2223 28866 2247 28890 nw
tri 2389 28866 2413 28890 ne
rect 2177 28816 2223 28856
rect 2177 28782 2183 28816
rect 2217 28782 2223 28816
rect 2177 28742 2223 28782
rect 2177 28708 2183 28742
rect 2217 28708 2223 28742
rect 2177 28668 2223 28708
rect 2177 28634 2183 28668
rect 2217 28634 2223 28668
rect 2177 28594 2223 28634
rect 2177 28560 2183 28594
rect 2217 28560 2223 28594
rect 2177 28520 2223 28560
rect 2177 28486 2183 28520
rect 2217 28486 2223 28520
rect 2177 28474 2223 28486
rect 2413 28856 2419 28890
rect 2453 28856 2459 28890
tri 2459 28866 2483 28890 nw
tri 2625 28866 2649 28890 ne
rect 2413 28816 2459 28856
rect 2413 28782 2419 28816
rect 2453 28782 2459 28816
rect 2413 28742 2459 28782
rect 2413 28708 2419 28742
rect 2453 28708 2459 28742
rect 2413 28668 2459 28708
rect 2413 28634 2419 28668
rect 2453 28634 2459 28668
rect 2413 28594 2459 28634
rect 2413 28560 2419 28594
rect 2453 28560 2459 28594
rect 2413 28520 2459 28560
rect 2413 28486 2419 28520
rect 2453 28486 2459 28520
rect 2413 28474 2459 28486
rect 2649 28856 2655 28890
rect 2689 28856 2695 28890
tri 2695 28866 2719 28890 nw
tri 2861 28866 2885 28890 ne
rect 2649 28816 2695 28856
rect 2649 28782 2655 28816
rect 2689 28782 2695 28816
rect 2649 28742 2695 28782
rect 2649 28708 2655 28742
rect 2689 28708 2695 28742
rect 2649 28668 2695 28708
rect 2649 28634 2655 28668
rect 2689 28634 2695 28668
rect 2649 28594 2695 28634
rect 2649 28560 2655 28594
rect 2689 28560 2695 28594
rect 2649 28520 2695 28560
rect 2649 28486 2655 28520
rect 2689 28486 2695 28520
rect 2649 28474 2695 28486
rect 2885 28856 2891 28890
rect 2925 28882 3076 28890
rect 2925 28856 3036 28882
rect 2885 28848 3036 28856
rect 3070 28848 3076 28882
rect 2885 28816 3076 28848
rect 2885 28782 2891 28816
rect 2925 28810 3076 28816
rect 2925 28782 3036 28810
rect 2885 28776 3036 28782
rect 3070 28776 3076 28810
rect 2885 28742 3076 28776
rect 2885 28708 2891 28742
rect 2925 28738 3076 28742
rect 2925 28708 3036 28738
rect 2885 28704 3036 28708
rect 3070 28704 3076 28738
rect 2885 28668 3076 28704
rect 2885 28634 2891 28668
rect 2925 28666 3076 28668
rect 2925 28634 3036 28666
rect 2885 28632 3036 28634
rect 3070 28632 3076 28666
rect 2885 28594 3076 28632
rect 2885 28560 2891 28594
rect 2925 28560 3036 28594
rect 3070 28560 3076 28594
rect 2885 28522 3076 28560
rect 2885 28520 3036 28522
rect 2885 28486 2891 28520
rect 2925 28488 3036 28520
rect 3070 28488 3076 28522
rect 2925 28486 3076 28488
rect 380 28431 571 28469
rect 380 28397 386 28431
rect 420 28397 571 28431
rect 2885 28450 3076 28486
rect 2885 28416 3036 28450
rect 3070 28416 3076 28450
rect 380 28359 571 28397
rect 613 28404 1501 28413
rect 1553 28404 1569 28413
rect 1621 28404 1636 28413
rect 1688 28404 1703 28413
rect 1755 28404 1770 28413
rect 1822 28404 1837 28413
rect 1889 28404 2830 28413
rect 613 28370 625 28404
rect 659 28370 700 28404
rect 734 28370 775 28404
rect 809 28370 850 28404
rect 884 28370 925 28404
rect 959 28370 1000 28404
rect 1034 28370 1075 28404
rect 1109 28370 1150 28404
rect 1184 28370 1225 28404
rect 1259 28370 1300 28404
rect 1334 28370 1375 28404
rect 1409 28370 1450 28404
rect 1484 28370 1501 28404
rect 1559 28370 1569 28404
rect 1634 28370 1636 28404
rect 1889 28370 1896 28404
rect 1930 28370 1970 28404
rect 2004 28370 2044 28404
rect 2078 28370 2118 28404
rect 2152 28370 2192 28404
rect 2226 28370 2266 28404
rect 2300 28370 2340 28404
rect 2374 28370 2414 28404
rect 2448 28370 2488 28404
rect 2522 28370 2562 28404
rect 2596 28370 2636 28404
rect 2670 28370 2710 28404
rect 2744 28370 2784 28404
rect 2818 28370 2830 28404
rect 613 28361 1501 28370
rect 1553 28361 1569 28370
rect 1621 28361 1636 28370
rect 1688 28361 1703 28370
rect 1755 28361 1770 28370
rect 1822 28361 1837 28370
rect 1889 28361 2830 28370
rect 2885 28378 3076 28416
rect 380 28325 386 28359
rect 420 28325 571 28359
rect 380 28288 571 28325
rect 2885 28344 3036 28378
rect 3070 28344 3076 28378
rect 2885 28306 3076 28344
rect 380 28287 531 28288
rect 380 28253 386 28287
rect 420 28254 531 28287
rect 565 28254 571 28288
rect 420 28253 571 28254
rect 380 28215 571 28253
rect 380 28181 386 28215
rect 420 28181 531 28215
rect 565 28181 571 28215
rect 380 28143 571 28181
rect 380 28109 386 28143
rect 420 28142 571 28143
rect 420 28109 531 28142
rect 380 28108 531 28109
rect 565 28108 571 28142
rect 380 28071 571 28108
rect 380 28037 386 28071
rect 420 28069 571 28071
rect 420 28037 531 28069
rect 380 28035 531 28037
rect 565 28035 571 28069
rect 380 27999 571 28035
rect 380 27965 386 27999
rect 420 27996 571 27999
rect 420 27965 531 27996
rect 380 27962 531 27965
rect 565 27962 571 27996
rect 380 27927 571 27962
rect 380 27893 386 27927
rect 420 27923 571 27927
rect 420 27893 531 27923
rect 380 27889 531 27893
rect 565 27889 571 27923
rect 761 28288 807 28300
rect 761 28254 767 28288
rect 801 28254 807 28288
rect 761 28215 807 28254
rect 761 28181 767 28215
rect 801 28181 807 28215
rect 761 28142 807 28181
rect 761 28108 767 28142
rect 801 28108 807 28142
rect 761 28069 807 28108
rect 761 28035 767 28069
rect 801 28035 807 28069
rect 761 27996 807 28035
rect 761 27962 767 27996
rect 801 27962 807 27996
rect 761 27923 807 27962
tri 571 27889 598 27916 sw
tri 734 27889 761 27916 se
rect 761 27889 767 27923
rect 801 27889 807 27923
rect 997 28288 1043 28300
rect 997 28254 1003 28288
rect 1037 28254 1043 28288
rect 997 28215 1043 28254
rect 997 28181 1003 28215
rect 1037 28181 1043 28215
rect 997 28142 1043 28181
rect 997 28108 1003 28142
rect 1037 28108 1043 28142
rect 997 28069 1043 28108
rect 997 28035 1003 28069
rect 1037 28035 1043 28069
rect 997 27996 1043 28035
rect 997 27962 1003 27996
rect 1037 27962 1043 27996
rect 997 27923 1043 27962
tri 807 27889 834 27916 sw
tri 970 27889 997 27916 se
rect 997 27889 1003 27923
rect 1037 27889 1043 27923
rect 1233 28288 1279 28300
rect 1233 28254 1239 28288
rect 1273 28254 1279 28288
rect 1233 28215 1279 28254
rect 1233 28181 1239 28215
rect 1273 28181 1279 28215
rect 1233 28142 1279 28181
rect 1233 28108 1239 28142
rect 1273 28108 1279 28142
rect 1233 28069 1279 28108
rect 1233 28035 1239 28069
rect 1273 28035 1279 28069
rect 1233 27996 1279 28035
rect 1233 27962 1239 27996
rect 1273 27962 1279 27996
rect 1233 27923 1279 27962
tri 1043 27889 1070 27916 sw
tri 1206 27889 1233 27916 se
rect 1233 27889 1239 27923
rect 1273 27889 1279 27923
rect 1469 28288 1515 28300
rect 1469 28254 1475 28288
rect 1509 28254 1515 28288
rect 1469 28215 1515 28254
rect 1469 28181 1475 28215
rect 1509 28181 1515 28215
rect 1469 28142 1515 28181
rect 1469 28108 1475 28142
rect 1509 28108 1515 28142
rect 1469 28069 1515 28108
rect 1469 28035 1475 28069
rect 1509 28035 1515 28069
rect 1469 27996 1515 28035
rect 1469 27962 1475 27996
rect 1509 27962 1515 27996
rect 1469 27923 1515 27962
tri 1279 27889 1306 27916 sw
tri 1442 27889 1469 27916 se
rect 1469 27889 1475 27923
rect 1509 27889 1515 27923
rect 1705 28288 1751 28300
rect 1705 28254 1711 28288
rect 1745 28254 1751 28288
rect 1705 28215 1751 28254
rect 1705 28181 1711 28215
rect 1745 28181 1751 28215
rect 1705 28142 1751 28181
rect 1705 28108 1711 28142
rect 1745 28108 1751 28142
rect 1705 28069 1751 28108
rect 1705 28035 1711 28069
rect 1745 28035 1751 28069
rect 1705 27996 1751 28035
rect 1705 27962 1711 27996
rect 1745 27962 1751 27996
rect 1705 27923 1751 27962
tri 1515 27889 1542 27916 sw
tri 1678 27889 1705 27916 se
rect 1705 27889 1711 27923
rect 1745 27889 1751 27923
rect 1941 28288 1987 28300
rect 1941 28254 1947 28288
rect 1981 28254 1987 28288
rect 1941 28215 1987 28254
rect 1941 28181 1947 28215
rect 1981 28181 1987 28215
rect 1941 28142 1987 28181
rect 1941 28108 1947 28142
rect 1981 28108 1987 28142
rect 1941 28069 1987 28108
rect 1941 28035 1947 28069
rect 1981 28035 1987 28069
rect 1941 27996 1987 28035
rect 1941 27962 1947 27996
rect 1981 27962 1987 27996
rect 1941 27923 1987 27962
tri 1751 27889 1778 27916 sw
tri 1914 27889 1941 27916 se
rect 1941 27889 1947 27923
rect 1981 27889 1987 27923
rect 2177 28288 2223 28300
rect 2177 28254 2183 28288
rect 2217 28254 2223 28288
rect 2177 28215 2223 28254
rect 2177 28181 2183 28215
rect 2217 28181 2223 28215
rect 2177 28142 2223 28181
rect 2177 28108 2183 28142
rect 2217 28108 2223 28142
rect 2177 28069 2223 28108
rect 2177 28035 2183 28069
rect 2217 28035 2223 28069
rect 2177 27996 2223 28035
rect 2177 27962 2183 27996
rect 2217 27962 2223 27996
rect 2177 27923 2223 27962
tri 1987 27889 2014 27916 sw
tri 2150 27889 2177 27916 se
rect 2177 27889 2183 27923
rect 2217 27889 2223 27923
rect 2413 28288 2459 28300
rect 2413 28254 2419 28288
rect 2453 28254 2459 28288
rect 2413 28215 2459 28254
rect 2413 28181 2419 28215
rect 2453 28181 2459 28215
rect 2413 28142 2459 28181
rect 2413 28108 2419 28142
rect 2453 28108 2459 28142
rect 2413 28069 2459 28108
rect 2413 28035 2419 28069
rect 2453 28035 2459 28069
rect 2413 27996 2459 28035
rect 2413 27962 2419 27996
rect 2453 27962 2459 27996
rect 2413 27923 2459 27962
tri 2223 27889 2250 27916 sw
tri 2386 27889 2413 27916 se
rect 2413 27889 2419 27923
rect 2453 27889 2459 27923
rect 2649 28288 2695 28300
rect 2649 28254 2655 28288
rect 2689 28254 2695 28288
rect 2649 28215 2695 28254
rect 2649 28181 2655 28215
rect 2689 28181 2695 28215
rect 2649 28142 2695 28181
rect 2649 28108 2655 28142
rect 2689 28108 2695 28142
rect 2649 28069 2695 28108
rect 2649 28035 2655 28069
rect 2689 28035 2695 28069
rect 2649 27996 2695 28035
rect 2649 27962 2655 27996
rect 2689 27962 2695 27996
rect 2649 27923 2695 27962
tri 2459 27889 2486 27916 sw
tri 2622 27889 2649 27916 se
rect 2649 27889 2655 27923
rect 2689 27889 2695 27923
rect 2885 28288 3036 28306
rect 2885 28254 2891 28288
rect 2925 28272 3036 28288
rect 3070 28272 3076 28306
rect 2925 28254 3076 28272
rect 2885 28234 3076 28254
rect 2885 28215 3036 28234
rect 2885 28181 2891 28215
rect 2925 28200 3036 28215
rect 3070 28200 3076 28234
rect 2925 28181 3076 28200
rect 2885 28162 3076 28181
rect 2885 28142 3036 28162
rect 2885 28108 2891 28142
rect 2925 28128 3036 28142
rect 3070 28128 3076 28162
rect 2925 28108 3076 28128
rect 2885 28090 3076 28108
rect 2885 28069 3036 28090
rect 2885 28035 2891 28069
rect 2925 28056 3036 28069
rect 3070 28056 3076 28090
rect 2925 28035 3076 28056
rect 2885 28018 3076 28035
rect 2885 27996 3036 28018
rect 2885 27962 2891 27996
rect 2925 27984 3036 27996
rect 3070 27984 3076 28018
rect 2925 27962 3076 27984
rect 2885 27946 3076 27962
rect 2885 27923 3036 27946
tri 2695 27889 2722 27916 sw
tri 2858 27889 2885 27916 se
rect 2885 27889 2891 27923
rect 2925 27912 3036 27923
rect 3070 27912 3076 27946
rect 2925 27889 3076 27912
rect 380 27888 598 27889
tri 598 27888 599 27889 sw
tri 733 27888 734 27889 se
rect 734 27888 834 27889
tri 834 27888 835 27889 sw
tri 969 27888 970 27889 se
rect 970 27888 1070 27889
tri 1070 27888 1071 27889 sw
tri 1205 27888 1206 27889 se
rect 1206 27888 1306 27889
tri 1306 27888 1307 27889 sw
tri 1441 27888 1442 27889 se
rect 1442 27888 1542 27889
tri 1542 27888 1543 27889 sw
tri 1677 27888 1678 27889 se
rect 1678 27888 1778 27889
tri 1778 27888 1779 27889 sw
tri 1913 27888 1914 27889 se
rect 1914 27888 2014 27889
tri 2014 27888 2015 27889 sw
tri 2149 27888 2150 27889 se
rect 2150 27888 2250 27889
tri 2250 27888 2251 27889 sw
tri 2385 27888 2386 27889 se
rect 2386 27888 2486 27889
tri 2486 27888 2487 27889 sw
tri 2621 27888 2622 27889 se
rect 2622 27888 2722 27889
tri 2722 27888 2723 27889 sw
tri 2857 27888 2858 27889 se
rect 2858 27888 3076 27889
rect 380 27882 599 27888
tri 599 27882 605 27888 sw
tri 727 27882 733 27888 se
rect 733 27882 835 27888
tri 835 27882 841 27888 sw
tri 963 27882 969 27888 se
rect 969 27882 1071 27888
tri 1071 27882 1077 27888 sw
tri 1199 27882 1205 27888 se
rect 1205 27882 1307 27888
tri 1307 27882 1313 27888 sw
tri 1435 27882 1441 27888 se
rect 1441 27882 1543 27888
tri 1543 27882 1549 27888 sw
tri 1671 27882 1677 27888 se
rect 1677 27882 1779 27888
tri 1779 27882 1785 27888 sw
tri 1907 27882 1913 27888 se
rect 1913 27882 2015 27888
tri 2015 27882 2021 27888 sw
tri 2143 27882 2149 27888 se
rect 2149 27882 2251 27888
tri 2251 27882 2257 27888 sw
tri 2379 27882 2385 27888 se
rect 2385 27882 2487 27888
tri 2487 27882 2493 27888 sw
tri 2615 27882 2621 27888 se
rect 2621 27882 2723 27888
tri 2723 27882 2729 27888 sw
tri 2851 27882 2857 27888 se
rect 2857 27882 3076 27888
rect 380 27874 3076 27882
rect 380 27865 3036 27874
rect 380 27855 697 27865
rect 380 27821 386 27855
rect 420 27850 697 27855
rect 420 27821 531 27850
rect 380 27816 531 27821
rect 565 27816 697 27850
rect 380 27813 697 27816
rect 749 27813 765 27865
rect 817 27813 833 27865
rect 885 27813 901 27865
rect 953 27813 969 27865
rect 1021 27850 1037 27865
rect 1021 27813 1037 27816
rect 1089 27813 1105 27865
rect 1157 27813 1173 27865
rect 1225 27850 1241 27865
rect 1293 27850 2097 27865
rect 1225 27816 1239 27850
rect 1293 27816 1475 27850
rect 1509 27816 1711 27850
rect 1745 27816 1947 27850
rect 1981 27816 2097 27850
rect 1225 27813 1241 27816
rect 1293 27813 2097 27816
rect 2149 27813 2165 27865
rect 2217 27813 2233 27865
rect 2285 27813 2301 27865
rect 2353 27813 2369 27865
rect 2421 27850 2437 27865
rect 2421 27813 2437 27816
rect 2489 27813 2505 27865
rect 2557 27813 2573 27865
rect 2625 27813 2641 27865
rect 2693 27850 3036 27865
rect 2693 27816 2891 27850
rect 2925 27840 3036 27850
rect 3070 27840 3076 27874
rect 2925 27816 3076 27840
rect 2693 27813 3076 27816
rect 380 27802 3076 27813
rect 380 27801 3036 27802
rect 380 27783 697 27801
rect 380 27749 386 27783
rect 420 27777 697 27783
rect 420 27749 531 27777
rect 380 27743 531 27749
rect 565 27749 697 27777
rect 749 27749 765 27801
rect 817 27749 833 27801
rect 885 27749 901 27801
rect 953 27749 969 27801
rect 1021 27777 1037 27801
rect 1089 27749 1105 27801
rect 1157 27749 1173 27801
rect 1225 27777 1241 27801
rect 1293 27777 2097 27801
rect 1225 27749 1239 27777
rect 1293 27749 1475 27777
rect 565 27743 767 27749
rect 801 27743 1003 27749
rect 1037 27743 1239 27749
rect 1273 27743 1475 27749
rect 1509 27743 1711 27777
rect 1745 27743 1947 27777
rect 1981 27749 2097 27777
rect 2149 27749 2165 27801
rect 2217 27749 2233 27801
rect 2285 27749 2301 27801
rect 2353 27749 2369 27801
rect 2421 27777 2437 27801
rect 2489 27749 2505 27801
rect 2557 27749 2573 27801
rect 2625 27749 2641 27801
rect 2693 27777 3036 27801
rect 2693 27749 2891 27777
rect 1981 27743 2183 27749
rect 2217 27743 2419 27749
rect 2453 27743 2655 27749
rect 2689 27743 2891 27749
rect 2925 27768 3036 27777
rect 3070 27768 3076 27802
rect 2925 27743 3076 27768
rect 380 27737 3076 27743
rect 380 27711 697 27737
rect 380 27677 386 27711
rect 420 27704 697 27711
rect 420 27677 531 27704
rect 380 27670 531 27677
rect 565 27685 697 27704
rect 749 27685 765 27737
rect 817 27685 833 27737
rect 885 27685 901 27737
rect 953 27685 969 27737
rect 1021 27704 1037 27737
rect 1089 27685 1105 27737
rect 1157 27685 1173 27737
rect 1225 27704 1241 27737
rect 1293 27704 2097 27737
rect 1225 27685 1239 27704
rect 1293 27685 1475 27704
rect 565 27673 767 27685
rect 801 27673 1003 27685
rect 1037 27673 1239 27685
rect 1273 27673 1475 27685
rect 565 27670 697 27673
rect 380 27639 697 27670
rect 380 27605 386 27639
rect 420 27631 697 27639
rect 420 27605 531 27631
rect 380 27597 531 27605
rect 565 27621 697 27631
rect 749 27621 765 27673
rect 817 27621 833 27673
rect 885 27621 901 27673
rect 953 27621 969 27673
rect 1021 27631 1037 27670
rect 1089 27621 1105 27673
rect 1157 27621 1173 27673
rect 1225 27670 1239 27673
rect 1293 27670 1475 27673
rect 1509 27670 1711 27704
rect 1745 27670 1947 27704
rect 1981 27685 2097 27704
rect 2149 27685 2165 27737
rect 2217 27685 2233 27737
rect 2285 27685 2301 27737
rect 2353 27685 2369 27737
rect 2421 27704 2437 27737
rect 2489 27685 2505 27737
rect 2557 27685 2573 27737
rect 2625 27685 2641 27737
rect 2693 27730 3076 27737
rect 2693 27704 3036 27730
rect 2693 27685 2891 27704
rect 1981 27673 2183 27685
rect 2217 27673 2419 27685
rect 2453 27673 2655 27685
rect 2689 27673 2891 27685
rect 1981 27670 2097 27673
rect 1225 27631 1241 27670
rect 1293 27631 2097 27670
rect 1225 27621 1239 27631
rect 1293 27621 1475 27631
rect 565 27609 767 27621
rect 801 27609 1003 27621
rect 1037 27609 1239 27621
rect 1273 27609 1475 27621
rect 565 27597 697 27609
rect 380 27567 697 27597
rect 380 27533 386 27567
rect 420 27558 697 27567
rect 420 27533 531 27558
rect 380 27524 531 27533
rect 565 27557 697 27558
rect 749 27557 765 27609
rect 817 27557 833 27609
rect 885 27557 901 27609
rect 953 27557 969 27609
rect 1021 27558 1037 27597
rect 1089 27557 1105 27609
rect 1157 27557 1173 27609
rect 1225 27597 1239 27609
rect 1293 27597 1475 27609
rect 1509 27597 1711 27631
rect 1745 27597 1947 27631
rect 1981 27621 2097 27631
rect 2149 27621 2165 27673
rect 2217 27621 2233 27673
rect 2285 27621 2301 27673
rect 2353 27621 2369 27673
rect 2421 27631 2437 27670
rect 2489 27621 2505 27673
rect 2557 27621 2573 27673
rect 2625 27621 2641 27673
rect 2693 27670 2891 27673
rect 2925 27696 3036 27704
rect 3070 27696 3076 27730
rect 2925 27670 3076 27696
rect 2693 27658 3076 27670
rect 2693 27631 3036 27658
rect 2693 27621 2891 27631
rect 1981 27609 2183 27621
rect 2217 27609 2419 27621
rect 2453 27609 2655 27621
rect 2689 27609 2891 27621
rect 1981 27597 2097 27609
rect 1225 27558 1241 27597
rect 1293 27558 2097 27597
rect 1225 27557 1239 27558
rect 1293 27557 1475 27558
rect 565 27545 767 27557
rect 801 27545 1003 27557
rect 1037 27545 1239 27557
rect 1273 27545 1475 27557
rect 565 27524 697 27545
rect 380 27495 697 27524
rect 380 27461 386 27495
rect 420 27493 697 27495
rect 749 27493 765 27545
rect 817 27493 833 27545
rect 885 27493 901 27545
rect 953 27493 969 27545
rect 1021 27493 1037 27524
rect 1089 27493 1105 27545
rect 1157 27493 1173 27545
rect 1225 27524 1239 27545
rect 1293 27524 1475 27545
rect 1509 27524 1711 27558
rect 1745 27524 1947 27558
rect 1981 27557 2097 27558
rect 2149 27557 2165 27609
rect 2217 27557 2233 27609
rect 2285 27557 2301 27609
rect 2353 27557 2369 27609
rect 2421 27558 2437 27597
rect 2489 27557 2505 27609
rect 2557 27557 2573 27609
rect 2625 27557 2641 27609
rect 2693 27597 2891 27609
rect 2925 27624 3036 27631
rect 3070 27624 3076 27658
rect 2925 27597 3076 27624
rect 2693 27586 3076 27597
rect 2693 27558 3036 27586
rect 2693 27557 2891 27558
rect 1981 27545 2183 27557
rect 2217 27545 2419 27557
rect 2453 27545 2655 27557
rect 2689 27545 2891 27557
rect 1981 27524 2097 27545
rect 1225 27493 1241 27524
rect 1293 27493 2097 27524
rect 2149 27493 2165 27545
rect 2217 27493 2233 27545
rect 2285 27493 2301 27545
rect 2353 27493 2369 27545
rect 2421 27493 2437 27524
rect 2489 27493 2505 27545
rect 2557 27493 2573 27545
rect 2625 27493 2641 27545
rect 2693 27524 2891 27545
rect 2925 27552 3036 27558
rect 3070 27552 3076 27586
rect 2925 27524 3076 27552
rect 2693 27514 3076 27524
rect 2693 27493 3036 27514
rect 420 27485 3036 27493
rect 420 27461 531 27485
rect 380 27451 531 27461
rect 565 27481 767 27485
rect 801 27481 1003 27485
rect 1037 27481 1239 27485
rect 1273 27481 1475 27485
rect 565 27451 697 27481
rect 380 27429 697 27451
rect 749 27429 765 27481
rect 817 27429 833 27481
rect 885 27429 901 27481
rect 953 27429 969 27481
rect 1021 27429 1037 27451
rect 1089 27429 1105 27481
rect 1157 27429 1173 27481
rect 1225 27451 1239 27481
rect 1293 27451 1475 27481
rect 1509 27451 1711 27485
rect 1745 27451 1947 27485
rect 1981 27481 2183 27485
rect 2217 27481 2419 27485
rect 2453 27481 2655 27485
rect 2689 27481 2891 27485
rect 1981 27451 2097 27481
rect 1225 27429 1241 27451
rect 1293 27429 2097 27451
rect 2149 27429 2165 27481
rect 2217 27429 2233 27481
rect 2285 27429 2301 27481
rect 2353 27429 2369 27481
rect 2421 27429 2437 27451
rect 2489 27429 2505 27481
rect 2557 27429 2573 27481
rect 2625 27429 2641 27481
rect 2693 27451 2891 27481
rect 2925 27480 3036 27485
rect 3070 27480 3076 27514
rect 2925 27451 3076 27480
rect 2693 27442 3076 27451
rect 2693 27429 3036 27442
rect 380 27423 3036 27429
rect 380 27389 386 27423
rect 420 27417 3036 27423
rect 420 27412 697 27417
rect 420 27389 531 27412
rect 380 27378 531 27389
rect 565 27378 697 27412
rect 380 27365 697 27378
rect 749 27365 765 27417
rect 817 27365 833 27417
rect 885 27365 901 27417
rect 953 27365 969 27417
rect 1021 27412 1037 27417
rect 1021 27365 1037 27378
rect 1089 27365 1105 27417
rect 1157 27365 1173 27417
rect 1225 27412 1241 27417
rect 1293 27412 2097 27417
rect 1225 27378 1239 27412
rect 1293 27378 1475 27412
rect 1509 27378 1711 27412
rect 1745 27378 1947 27412
rect 1981 27378 2097 27412
rect 1225 27365 1241 27378
rect 1293 27365 2097 27378
rect 2149 27365 2165 27417
rect 2217 27365 2233 27417
rect 2285 27365 2301 27417
rect 2353 27365 2369 27417
rect 2421 27412 2437 27417
rect 2421 27365 2437 27378
rect 2489 27365 2505 27417
rect 2557 27365 2573 27417
rect 2625 27365 2641 27417
rect 2693 27412 3036 27417
rect 2693 27378 2891 27412
rect 2925 27408 3036 27412
rect 3070 27408 3076 27442
rect 2925 27378 3076 27408
rect 2693 27370 3076 27378
rect 2693 27365 3036 27370
rect 380 27353 3036 27365
rect 380 27351 697 27353
rect 380 27317 386 27351
rect 420 27338 697 27351
rect 420 27317 531 27338
rect 380 27304 531 27317
rect 565 27304 697 27338
rect 380 27301 697 27304
rect 749 27301 765 27353
rect 817 27301 833 27353
rect 885 27301 901 27353
rect 953 27301 969 27353
rect 1021 27338 1037 27353
rect 1021 27301 1037 27304
rect 1089 27301 1105 27353
rect 1157 27301 1173 27353
rect 1225 27338 1241 27353
rect 1293 27338 2097 27353
rect 1225 27304 1239 27338
rect 1293 27304 1475 27338
rect 1509 27304 1711 27338
rect 1745 27304 1947 27338
rect 1981 27304 2097 27338
rect 1225 27301 1241 27304
rect 1293 27301 2097 27304
rect 2149 27301 2165 27353
rect 2217 27301 2233 27353
rect 2285 27301 2301 27353
rect 2353 27301 2369 27353
rect 2421 27338 2437 27353
rect 2421 27301 2437 27304
rect 2489 27301 2505 27353
rect 2557 27301 2573 27353
rect 2625 27301 2641 27353
rect 2693 27338 3036 27353
rect 2693 27304 2891 27338
rect 2925 27336 3036 27338
rect 3070 27336 3076 27370
rect 2925 27304 3076 27336
rect 2693 27301 3076 27304
rect 380 27298 3076 27301
rect 380 27289 3036 27298
rect 380 27279 697 27289
rect 380 27245 386 27279
rect 420 27264 697 27279
rect 420 27245 531 27264
rect 380 27230 531 27245
rect 565 27237 697 27264
rect 749 27237 765 27289
rect 817 27237 833 27289
rect 885 27237 901 27289
rect 953 27237 969 27289
rect 1021 27264 1037 27289
rect 1089 27237 1105 27289
rect 1157 27237 1173 27289
rect 1225 27264 1241 27289
rect 1293 27264 2097 27289
rect 1225 27237 1239 27264
rect 1293 27237 1475 27264
rect 565 27230 767 27237
rect 801 27230 1003 27237
rect 1037 27230 1239 27237
rect 1273 27230 1475 27237
rect 1509 27230 1711 27264
rect 1745 27230 1947 27264
rect 1981 27237 2097 27264
rect 2149 27237 2165 27289
rect 2217 27237 2233 27289
rect 2285 27237 2301 27289
rect 2353 27237 2369 27289
rect 2421 27264 2437 27289
rect 2489 27237 2505 27289
rect 2557 27237 2573 27289
rect 2625 27237 2641 27289
rect 2693 27264 3036 27289
rect 3070 27264 3076 27298
rect 2693 27237 2891 27264
rect 1981 27230 2183 27237
rect 2217 27230 2419 27237
rect 2453 27230 2655 27237
rect 2689 27230 2891 27237
rect 2925 27230 3076 27264
rect 380 27226 3076 27230
rect 380 27225 3036 27226
rect 380 27207 697 27225
rect 380 27173 386 27207
rect 420 27190 697 27207
rect 420 27173 531 27190
rect 380 27156 531 27173
rect 565 27173 697 27190
rect 749 27173 765 27225
rect 817 27173 833 27225
rect 885 27173 901 27225
rect 953 27173 969 27225
rect 1021 27190 1037 27225
rect 1089 27173 1105 27225
rect 1157 27173 1173 27225
rect 1225 27190 1241 27225
rect 1293 27190 2097 27225
rect 1225 27173 1239 27190
rect 1293 27173 1475 27190
rect 565 27161 767 27173
rect 801 27161 1003 27173
rect 1037 27161 1239 27173
rect 1273 27161 1475 27173
rect 565 27156 697 27161
rect 380 27135 697 27156
rect 380 27101 386 27135
rect 420 27116 697 27135
rect 420 27101 531 27116
rect 380 27082 531 27101
rect 565 27109 697 27116
rect 749 27109 765 27161
rect 817 27109 833 27161
rect 885 27109 901 27161
rect 953 27109 969 27161
rect 1021 27116 1037 27156
rect 1089 27109 1105 27161
rect 1157 27109 1173 27161
rect 1225 27156 1239 27161
rect 1293 27156 1475 27161
rect 1509 27156 1711 27190
rect 1745 27156 1947 27190
rect 1981 27173 2097 27190
rect 2149 27173 2165 27225
rect 2217 27173 2233 27225
rect 2285 27173 2301 27225
rect 2353 27173 2369 27225
rect 2421 27190 2437 27225
rect 2489 27173 2505 27225
rect 2557 27173 2573 27225
rect 2625 27173 2641 27225
rect 2693 27192 3036 27225
rect 3070 27192 3076 27226
rect 2693 27190 3076 27192
rect 2693 27173 2891 27190
rect 1981 27161 2183 27173
rect 2217 27161 2419 27173
rect 2453 27161 2655 27173
rect 2689 27161 2891 27173
rect 1981 27156 2097 27161
rect 1225 27116 1241 27156
rect 1293 27116 2097 27156
rect 1225 27109 1239 27116
rect 1293 27109 1475 27116
rect 565 27097 767 27109
rect 801 27097 1003 27109
rect 1037 27097 1239 27109
rect 1273 27097 1475 27109
rect 565 27082 697 27097
rect 380 27063 697 27082
rect 380 27029 386 27063
rect 420 27045 697 27063
rect 749 27045 765 27097
rect 817 27045 833 27097
rect 885 27045 901 27097
rect 953 27045 969 27097
rect 1021 27045 1037 27082
rect 1089 27045 1105 27097
rect 1157 27045 1173 27097
rect 1225 27082 1239 27097
rect 1293 27082 1475 27097
rect 1509 27082 1711 27116
rect 1745 27082 1947 27116
rect 1981 27109 2097 27116
rect 2149 27109 2165 27161
rect 2217 27109 2233 27161
rect 2285 27109 2301 27161
rect 2353 27109 2369 27161
rect 2421 27116 2437 27156
rect 2489 27109 2505 27161
rect 2557 27109 2573 27161
rect 2625 27109 2641 27161
rect 2693 27156 2891 27161
rect 2925 27156 3076 27190
rect 2693 27154 3076 27156
rect 2693 27120 3036 27154
rect 3070 27120 3076 27154
rect 2693 27116 3076 27120
rect 2693 27109 2891 27116
rect 1981 27097 2183 27109
rect 2217 27097 2419 27109
rect 2453 27097 2655 27109
rect 2689 27097 2891 27109
rect 1981 27082 2097 27097
rect 1225 27045 1241 27082
rect 1293 27045 2097 27082
rect 2149 27045 2165 27097
rect 2217 27045 2233 27097
rect 2285 27045 2301 27097
rect 2353 27045 2369 27097
rect 2421 27045 2437 27082
rect 2489 27045 2505 27097
rect 2557 27045 2573 27097
rect 2625 27045 2641 27097
rect 2693 27082 2891 27097
rect 2925 27082 3076 27116
rect 2693 27048 3036 27082
rect 3070 27048 3076 27082
rect 2693 27045 3076 27048
rect 420 27042 3076 27045
rect 420 27029 531 27042
rect 380 27008 531 27029
rect 565 27033 767 27042
rect 801 27033 1003 27042
rect 1037 27033 1239 27042
rect 1273 27033 1475 27042
rect 565 27008 697 27033
rect 380 26991 697 27008
rect 380 26957 386 26991
rect 420 26981 697 26991
rect 749 26981 765 27033
rect 817 26981 833 27033
rect 885 26981 901 27033
rect 953 26981 969 27033
rect 1021 26981 1037 27008
rect 1089 26981 1105 27033
rect 1157 26981 1173 27033
rect 1225 27008 1239 27033
rect 1293 27008 1475 27033
rect 1509 27008 1711 27042
rect 1745 27008 1947 27042
rect 1981 27033 2183 27042
rect 2217 27033 2419 27042
rect 2453 27033 2655 27042
rect 2689 27033 2891 27042
rect 1981 27008 2097 27033
rect 1225 26981 1241 27008
rect 1293 26981 2097 27008
rect 2149 26981 2165 27033
rect 2217 26981 2233 27033
rect 2285 26981 2301 27033
rect 2353 26981 2369 27033
rect 2421 26981 2437 27008
rect 2489 26981 2505 27033
rect 2557 26981 2573 27033
rect 2625 26981 2641 27033
rect 2693 27008 2891 27033
rect 2925 27010 3076 27042
rect 2925 27008 3036 27010
rect 2693 26981 3036 27008
rect 420 26976 3036 26981
rect 3070 26976 3076 27010
rect 420 26969 3076 26976
rect 420 26968 697 26969
rect 420 26957 531 26968
rect 380 26934 531 26957
rect 565 26934 697 26968
rect 380 26919 697 26934
rect 380 26885 386 26919
rect 420 26917 697 26919
rect 749 26917 765 26969
rect 817 26917 833 26969
rect 885 26917 901 26969
rect 953 26917 969 26969
rect 1021 26968 1037 26969
rect 1021 26917 1037 26934
rect 1089 26917 1105 26969
rect 1157 26917 1173 26969
rect 1225 26968 1241 26969
rect 1293 26968 2097 26969
rect 1225 26934 1239 26968
rect 1293 26934 1475 26968
rect 1509 26934 1711 26968
rect 1745 26934 1947 26968
rect 1981 26934 2097 26968
rect 1225 26917 1241 26934
rect 1293 26917 2097 26934
rect 2149 26917 2165 26969
rect 2217 26917 2233 26969
rect 2285 26917 2301 26969
rect 2353 26917 2369 26969
rect 2421 26968 2437 26969
rect 2421 26917 2437 26934
rect 2489 26917 2505 26969
rect 2557 26917 2573 26969
rect 2625 26917 2641 26969
rect 2693 26968 3076 26969
rect 2693 26934 2891 26968
rect 2925 26938 3076 26968
rect 2925 26934 3036 26938
rect 2693 26917 3036 26934
rect 420 26904 3036 26917
rect 3070 26904 3076 26938
rect 420 26894 3076 26904
rect 420 26885 531 26894
rect 380 26860 531 26885
rect 565 26882 767 26894
rect 565 26860 583 26882
tri 583 26860 605 26882 nw
tri 727 26860 749 26882 ne
rect 749 26860 767 26882
rect 801 26882 1003 26894
rect 801 26860 819 26882
tri 819 26860 841 26882 nw
tri 963 26860 985 26882 ne
rect 985 26860 1003 26882
rect 1037 26882 1239 26894
rect 1037 26860 1055 26882
tri 1055 26860 1077 26882 nw
tri 1199 26860 1221 26882 ne
rect 1221 26860 1239 26882
rect 1273 26882 1475 26894
rect 1273 26860 1291 26882
tri 1291 26860 1313 26882 nw
tri 1435 26860 1457 26882 ne
rect 1457 26860 1475 26882
rect 1509 26882 1711 26894
rect 1509 26860 1527 26882
tri 1527 26860 1549 26882 nw
tri 1671 26860 1693 26882 ne
rect 1693 26860 1711 26882
rect 1745 26882 1947 26894
rect 1745 26860 1763 26882
tri 1763 26860 1785 26882 nw
tri 1907 26860 1929 26882 ne
rect 1929 26860 1947 26882
rect 1981 26882 2183 26894
rect 1981 26860 1999 26882
tri 1999 26860 2021 26882 nw
tri 2143 26860 2165 26882 ne
rect 2165 26860 2183 26882
rect 2217 26882 2419 26894
rect 2217 26860 2235 26882
tri 2235 26860 2257 26882 nw
tri 2379 26860 2401 26882 ne
rect 2401 26860 2419 26882
rect 2453 26882 2655 26894
rect 2453 26860 2471 26882
tri 2471 26860 2493 26882 nw
tri 2615 26860 2637 26882 ne
rect 2637 26860 2655 26882
rect 2689 26882 2891 26894
rect 2689 26860 2707 26882
tri 2707 26860 2729 26882 nw
tri 2851 26860 2873 26882 ne
rect 2873 26860 2891 26882
rect 2925 26866 3076 26894
rect 2925 26860 3036 26866
rect 380 26847 571 26860
tri 571 26848 583 26860 nw
tri 749 26848 761 26860 ne
rect 380 26813 386 26847
rect 420 26820 571 26847
rect 420 26813 531 26820
rect 380 26786 531 26813
rect 565 26786 571 26820
rect 380 26775 571 26786
rect 380 26741 386 26775
rect 420 26746 571 26775
rect 420 26741 531 26746
rect 380 26712 531 26741
rect 565 26712 571 26746
rect 380 26703 571 26712
rect 380 26669 386 26703
rect 420 26672 571 26703
rect 420 26669 531 26672
rect 380 26638 531 26669
rect 565 26638 571 26672
rect 380 26631 571 26638
rect 380 26597 386 26631
rect 420 26598 571 26631
rect 420 26597 531 26598
rect 380 26564 531 26597
rect 565 26564 571 26598
rect 380 26559 571 26564
rect 380 26525 386 26559
rect 420 26525 571 26559
rect 380 26524 571 26525
rect 380 26490 531 26524
rect 565 26490 571 26524
rect 380 26487 571 26490
rect 380 26453 386 26487
rect 420 26453 571 26487
rect 380 26450 571 26453
rect 380 26416 531 26450
rect 565 26416 571 26450
rect 380 26415 571 26416
rect 380 26381 386 26415
rect 420 26381 571 26415
rect 380 26376 571 26381
rect 380 26343 531 26376
rect 380 26309 386 26343
rect 420 26342 531 26343
rect 565 26342 571 26376
rect 420 26309 571 26342
rect 761 26820 807 26860
tri 807 26848 819 26860 nw
tri 985 26848 997 26860 ne
rect 761 26786 767 26820
rect 801 26786 807 26820
rect 761 26746 807 26786
rect 761 26712 767 26746
rect 801 26712 807 26746
rect 761 26672 807 26712
rect 761 26638 767 26672
rect 801 26638 807 26672
rect 761 26598 807 26638
rect 761 26564 767 26598
rect 801 26564 807 26598
rect 761 26524 807 26564
rect 761 26490 767 26524
rect 801 26490 807 26524
rect 761 26450 807 26490
rect 761 26416 767 26450
rect 801 26416 807 26450
rect 761 26376 807 26416
rect 761 26342 767 26376
rect 801 26342 807 26376
rect 761 26330 807 26342
rect 997 26820 1043 26860
tri 1043 26848 1055 26860 nw
tri 1221 26848 1233 26860 ne
rect 997 26786 1003 26820
rect 1037 26786 1043 26820
rect 997 26746 1043 26786
rect 997 26712 1003 26746
rect 1037 26712 1043 26746
rect 997 26672 1043 26712
rect 997 26638 1003 26672
rect 1037 26638 1043 26672
rect 997 26598 1043 26638
rect 997 26564 1003 26598
rect 1037 26564 1043 26598
rect 997 26524 1043 26564
rect 997 26490 1003 26524
rect 1037 26490 1043 26524
rect 997 26450 1043 26490
rect 997 26416 1003 26450
rect 1037 26416 1043 26450
rect 997 26376 1043 26416
rect 997 26342 1003 26376
rect 1037 26342 1043 26376
rect 997 26330 1043 26342
rect 1233 26820 1279 26860
tri 1279 26848 1291 26860 nw
tri 1457 26848 1469 26860 ne
rect 1233 26786 1239 26820
rect 1273 26786 1279 26820
rect 1233 26746 1279 26786
rect 1233 26712 1239 26746
rect 1273 26712 1279 26746
rect 1233 26672 1279 26712
rect 1233 26638 1239 26672
rect 1273 26638 1279 26672
rect 1233 26598 1279 26638
rect 1233 26564 1239 26598
rect 1273 26564 1279 26598
rect 1233 26524 1279 26564
rect 1233 26490 1239 26524
rect 1273 26490 1279 26524
rect 1233 26450 1279 26490
rect 1233 26416 1239 26450
rect 1273 26416 1279 26450
rect 1233 26376 1279 26416
rect 1233 26342 1239 26376
rect 1273 26342 1279 26376
rect 1233 26330 1279 26342
rect 1469 26820 1515 26860
tri 1515 26848 1527 26860 nw
tri 1693 26848 1705 26860 ne
rect 1469 26786 1475 26820
rect 1509 26786 1515 26820
rect 1469 26746 1515 26786
rect 1469 26712 1475 26746
rect 1509 26712 1515 26746
rect 1469 26672 1515 26712
rect 1469 26638 1475 26672
rect 1509 26638 1515 26672
rect 1469 26598 1515 26638
rect 1469 26564 1475 26598
rect 1509 26564 1515 26598
rect 1469 26524 1515 26564
rect 1469 26490 1475 26524
rect 1509 26490 1515 26524
rect 1469 26450 1515 26490
rect 1469 26416 1475 26450
rect 1509 26416 1515 26450
rect 1469 26376 1515 26416
rect 1469 26342 1475 26376
rect 1509 26342 1515 26376
rect 1469 26330 1515 26342
rect 1705 26820 1751 26860
tri 1751 26848 1763 26860 nw
tri 1929 26848 1941 26860 ne
rect 1705 26786 1711 26820
rect 1745 26786 1751 26820
rect 1705 26746 1751 26786
rect 1705 26712 1711 26746
rect 1745 26712 1751 26746
rect 1705 26672 1751 26712
rect 1705 26638 1711 26672
rect 1745 26638 1751 26672
rect 1705 26598 1751 26638
rect 1705 26564 1711 26598
rect 1745 26564 1751 26598
rect 1705 26524 1751 26564
rect 1705 26490 1711 26524
rect 1745 26490 1751 26524
rect 1705 26450 1751 26490
rect 1705 26416 1711 26450
rect 1745 26416 1751 26450
rect 1705 26376 1751 26416
rect 1705 26342 1711 26376
rect 1745 26342 1751 26376
rect 1705 26330 1751 26342
rect 1941 26820 1987 26860
tri 1987 26848 1999 26860 nw
tri 2165 26848 2177 26860 ne
rect 1941 26786 1947 26820
rect 1981 26786 1987 26820
rect 1941 26746 1987 26786
rect 1941 26712 1947 26746
rect 1981 26712 1987 26746
rect 1941 26672 1987 26712
rect 1941 26638 1947 26672
rect 1981 26638 1987 26672
rect 1941 26598 1987 26638
rect 1941 26564 1947 26598
rect 1981 26564 1987 26598
rect 1941 26524 1987 26564
rect 1941 26490 1947 26524
rect 1981 26490 1987 26524
rect 1941 26450 1987 26490
rect 1941 26416 1947 26450
rect 1981 26416 1987 26450
rect 1941 26376 1987 26416
rect 1941 26342 1947 26376
rect 1981 26342 1987 26376
rect 1941 26330 1987 26342
rect 2177 26820 2223 26860
tri 2223 26848 2235 26860 nw
tri 2401 26848 2413 26860 ne
rect 2177 26786 2183 26820
rect 2217 26786 2223 26820
rect 2177 26746 2223 26786
rect 2177 26712 2183 26746
rect 2217 26712 2223 26746
rect 2177 26672 2223 26712
rect 2177 26638 2183 26672
rect 2217 26638 2223 26672
rect 2177 26598 2223 26638
rect 2177 26564 2183 26598
rect 2217 26564 2223 26598
rect 2177 26524 2223 26564
rect 2177 26490 2183 26524
rect 2217 26490 2223 26524
rect 2177 26450 2223 26490
rect 2177 26416 2183 26450
rect 2217 26416 2223 26450
rect 2177 26376 2223 26416
rect 2177 26342 2183 26376
rect 2217 26342 2223 26376
rect 2177 26330 2223 26342
rect 2413 26820 2459 26860
tri 2459 26848 2471 26860 nw
tri 2637 26848 2649 26860 ne
rect 2413 26786 2419 26820
rect 2453 26786 2459 26820
rect 2413 26746 2459 26786
rect 2413 26712 2419 26746
rect 2453 26712 2459 26746
rect 2413 26672 2459 26712
rect 2413 26638 2419 26672
rect 2453 26638 2459 26672
rect 2413 26598 2459 26638
rect 2413 26564 2419 26598
rect 2453 26564 2459 26598
rect 2413 26524 2459 26564
rect 2413 26490 2419 26524
rect 2453 26490 2459 26524
rect 2413 26450 2459 26490
rect 2413 26416 2419 26450
rect 2453 26416 2459 26450
rect 2413 26376 2459 26416
rect 2413 26342 2419 26376
rect 2453 26342 2459 26376
rect 2413 26330 2459 26342
rect 2649 26820 2695 26860
tri 2695 26848 2707 26860 nw
tri 2873 26848 2885 26860 ne
rect 2649 26786 2655 26820
rect 2689 26786 2695 26820
rect 2649 26746 2695 26786
rect 2649 26712 2655 26746
rect 2689 26712 2695 26746
rect 2649 26672 2695 26712
rect 2649 26638 2655 26672
rect 2689 26638 2695 26672
rect 2649 26598 2695 26638
rect 2649 26564 2655 26598
rect 2689 26564 2695 26598
rect 2649 26524 2695 26564
rect 2649 26490 2655 26524
rect 2689 26490 2695 26524
rect 2649 26450 2695 26490
rect 2649 26416 2655 26450
rect 2689 26416 2695 26450
rect 2649 26376 2695 26416
rect 2649 26342 2655 26376
rect 2689 26342 2695 26376
rect 2649 26330 2695 26342
rect 2885 26832 3036 26860
rect 3070 26832 3076 26866
rect 2885 26820 3076 26832
rect 2885 26786 2891 26820
rect 2925 26794 3076 26820
rect 2925 26786 3036 26794
rect 2885 26760 3036 26786
rect 3070 26760 3076 26794
rect 2885 26746 3076 26760
rect 2885 26712 2891 26746
rect 2925 26722 3076 26746
rect 2925 26712 3036 26722
rect 2885 26688 3036 26712
rect 3070 26688 3076 26722
rect 2885 26672 3076 26688
rect 2885 26638 2891 26672
rect 2925 26650 3076 26672
rect 2925 26638 3036 26650
rect 2885 26616 3036 26638
rect 3070 26616 3076 26650
rect 2885 26598 3076 26616
rect 2885 26564 2891 26598
rect 2925 26578 3076 26598
rect 2925 26564 3036 26578
rect 2885 26544 3036 26564
rect 3070 26544 3076 26578
rect 2885 26524 3076 26544
rect 2885 26490 2891 26524
rect 2925 26506 3076 26524
rect 2925 26490 3036 26506
rect 2885 26472 3036 26490
rect 3070 26472 3076 26506
rect 2885 26450 3076 26472
rect 2885 26416 2891 26450
rect 2925 26434 3076 26450
rect 2925 26416 3036 26434
rect 2885 26400 3036 26416
rect 3070 26400 3076 26434
rect 2885 26376 3076 26400
rect 2885 26342 2891 26376
rect 2925 26362 3076 26376
rect 2925 26342 3036 26362
rect 380 26271 571 26309
rect 2885 26328 3036 26342
rect 3070 26328 3076 26362
rect 2885 26290 3076 26328
rect 380 26237 386 26271
rect 420 26237 571 26271
rect 380 26199 571 26237
rect 613 26274 1501 26283
rect 1553 26274 1569 26283
rect 1621 26274 1636 26283
rect 1688 26274 1703 26283
rect 1755 26274 1770 26283
rect 1822 26274 1837 26283
rect 1889 26274 2830 26283
rect 613 26240 625 26274
rect 659 26240 700 26274
rect 734 26240 775 26274
rect 809 26240 850 26274
rect 884 26240 925 26274
rect 959 26240 1000 26274
rect 1034 26240 1075 26274
rect 1109 26240 1150 26274
rect 1184 26240 1225 26274
rect 1259 26240 1300 26274
rect 1334 26240 1375 26274
rect 1409 26240 1450 26274
rect 1484 26240 1501 26274
rect 1559 26240 1569 26274
rect 1634 26240 1636 26274
rect 1889 26240 1896 26274
rect 1930 26240 1970 26274
rect 2004 26240 2044 26274
rect 2078 26240 2118 26274
rect 2152 26240 2192 26274
rect 2226 26240 2266 26274
rect 2300 26240 2340 26274
rect 2374 26240 2414 26274
rect 2448 26240 2488 26274
rect 2522 26240 2562 26274
rect 2596 26240 2636 26274
rect 2670 26240 2710 26274
rect 2744 26240 2784 26274
rect 2818 26240 2830 26274
rect 613 26231 1501 26240
rect 1553 26231 1569 26240
rect 1621 26231 1636 26240
rect 1688 26231 1703 26240
rect 1755 26231 1770 26240
rect 1822 26231 1837 26240
rect 1889 26231 2830 26240
rect 2885 26256 3036 26290
rect 3070 26256 3076 26290
rect 380 26165 386 26199
rect 420 26172 571 26199
rect 2885 26218 3076 26256
rect 2885 26184 3036 26218
rect 3070 26184 3076 26218
rect 420 26165 531 26172
rect 380 26138 531 26165
rect 565 26138 571 26172
rect 380 26127 571 26138
rect 380 26093 386 26127
rect 420 26099 571 26127
rect 420 26093 531 26099
rect 380 26065 531 26093
rect 565 26065 571 26099
rect 380 26055 571 26065
rect 380 26021 386 26055
rect 420 26026 571 26055
rect 420 26021 531 26026
rect 380 25992 531 26021
rect 565 25992 571 26026
rect 380 25983 571 25992
rect 380 25949 386 25983
rect 420 25953 571 25983
rect 420 25949 531 25953
rect 380 25919 531 25949
rect 565 25919 571 25953
rect 380 25911 571 25919
rect 380 25877 386 25911
rect 420 25880 571 25911
rect 420 25877 531 25880
rect 380 25846 531 25877
rect 565 25846 571 25880
rect 380 25839 571 25846
rect 380 25805 386 25839
rect 420 25807 571 25839
rect 420 25805 531 25807
rect 380 25773 531 25805
rect 565 25773 571 25807
rect 380 25767 571 25773
rect 380 25733 386 25767
rect 420 25734 571 25767
rect 761 26172 807 26184
rect 761 26138 767 26172
rect 801 26138 807 26172
rect 761 26099 807 26138
rect 761 26065 767 26099
rect 801 26065 807 26099
rect 761 26026 807 26065
rect 761 25992 767 26026
rect 801 25992 807 26026
rect 761 25953 807 25992
rect 761 25919 767 25953
rect 801 25919 807 25953
rect 761 25880 807 25919
rect 761 25846 767 25880
rect 801 25846 807 25880
rect 761 25807 807 25846
rect 761 25773 767 25807
rect 801 25773 807 25807
tri 571 25734 573 25736 sw
tri 759 25734 761 25736 se
rect 761 25734 807 25773
rect 997 26172 1043 26184
rect 997 26138 1003 26172
rect 1037 26138 1043 26172
rect 997 26099 1043 26138
rect 997 26065 1003 26099
rect 1037 26065 1043 26099
rect 997 26026 1043 26065
rect 997 25992 1003 26026
rect 1037 25992 1043 26026
rect 997 25953 1043 25992
rect 997 25919 1003 25953
rect 1037 25919 1043 25953
rect 997 25880 1043 25919
rect 997 25846 1003 25880
rect 1037 25846 1043 25880
rect 997 25807 1043 25846
rect 997 25773 1003 25807
rect 1037 25773 1043 25807
tri 807 25734 809 25736 sw
tri 995 25734 997 25736 se
rect 997 25734 1043 25773
rect 1233 26172 1279 26184
rect 1233 26138 1239 26172
rect 1273 26138 1279 26172
rect 1233 26099 1279 26138
rect 1233 26065 1239 26099
rect 1273 26065 1279 26099
rect 1233 26026 1279 26065
rect 1233 25992 1239 26026
rect 1273 25992 1279 26026
rect 1233 25953 1279 25992
rect 1233 25919 1239 25953
rect 1273 25919 1279 25953
rect 1233 25880 1279 25919
rect 1233 25846 1239 25880
rect 1273 25846 1279 25880
rect 1233 25807 1279 25846
rect 1233 25773 1239 25807
rect 1273 25773 1279 25807
tri 1043 25734 1045 25736 sw
tri 1231 25734 1233 25736 se
rect 1233 25734 1279 25773
rect 1469 26172 1515 26184
rect 1469 26138 1475 26172
rect 1509 26138 1515 26172
rect 1469 26099 1515 26138
rect 1469 26065 1475 26099
rect 1509 26065 1515 26099
rect 1469 26026 1515 26065
rect 1469 25992 1475 26026
rect 1509 25992 1515 26026
rect 1469 25953 1515 25992
rect 1469 25919 1475 25953
rect 1509 25919 1515 25953
rect 1469 25880 1515 25919
rect 1469 25846 1475 25880
rect 1509 25846 1515 25880
rect 1469 25807 1515 25846
rect 1469 25773 1475 25807
rect 1509 25773 1515 25807
tri 1279 25734 1281 25736 sw
tri 1467 25734 1469 25736 se
rect 1469 25734 1515 25773
rect 1705 26172 1751 26184
rect 1705 26138 1711 26172
rect 1745 26138 1751 26172
rect 1705 26099 1751 26138
rect 1705 26065 1711 26099
rect 1745 26065 1751 26099
rect 1705 26026 1751 26065
rect 1705 25992 1711 26026
rect 1745 25992 1751 26026
rect 1705 25953 1751 25992
rect 1705 25919 1711 25953
rect 1745 25919 1751 25953
rect 1705 25880 1751 25919
rect 1705 25846 1711 25880
rect 1745 25846 1751 25880
rect 1705 25807 1751 25846
rect 1705 25773 1711 25807
rect 1745 25773 1751 25807
tri 1515 25734 1517 25736 sw
tri 1703 25734 1705 25736 se
rect 1705 25734 1751 25773
rect 1941 26172 1987 26184
rect 1941 26138 1947 26172
rect 1981 26138 1987 26172
rect 1941 26099 1987 26138
rect 1941 26065 1947 26099
rect 1981 26065 1987 26099
rect 1941 26026 1987 26065
rect 1941 25992 1947 26026
rect 1981 25992 1987 26026
rect 1941 25953 1987 25992
rect 1941 25919 1947 25953
rect 1981 25919 1987 25953
rect 1941 25880 1987 25919
rect 1941 25846 1947 25880
rect 1981 25846 1987 25880
rect 1941 25807 1987 25846
rect 1941 25773 1947 25807
rect 1981 25773 1987 25807
tri 1751 25734 1753 25736 sw
tri 1939 25734 1941 25736 se
rect 1941 25734 1987 25773
rect 2177 26172 2223 26184
rect 2177 26138 2183 26172
rect 2217 26138 2223 26172
rect 2177 26099 2223 26138
rect 2177 26065 2183 26099
rect 2217 26065 2223 26099
rect 2177 26026 2223 26065
rect 2177 25992 2183 26026
rect 2217 25992 2223 26026
rect 2177 25953 2223 25992
rect 2177 25919 2183 25953
rect 2217 25919 2223 25953
rect 2177 25880 2223 25919
rect 2177 25846 2183 25880
rect 2217 25846 2223 25880
rect 2177 25807 2223 25846
rect 2177 25773 2183 25807
rect 2217 25773 2223 25807
tri 1987 25734 1989 25736 sw
tri 2175 25734 2177 25736 se
rect 2177 25734 2223 25773
rect 2413 26172 2459 26184
rect 2413 26138 2419 26172
rect 2453 26138 2459 26172
rect 2413 26099 2459 26138
rect 2413 26065 2419 26099
rect 2453 26065 2459 26099
rect 2413 26026 2459 26065
rect 2413 25992 2419 26026
rect 2453 25992 2459 26026
rect 2413 25953 2459 25992
rect 2413 25919 2419 25953
rect 2453 25919 2459 25953
rect 2413 25880 2459 25919
rect 2413 25846 2419 25880
rect 2453 25846 2459 25880
rect 2413 25807 2459 25846
rect 2413 25773 2419 25807
rect 2453 25773 2459 25807
tri 2223 25734 2225 25736 sw
tri 2411 25734 2413 25736 se
rect 2413 25734 2459 25773
rect 2649 26172 2695 26184
rect 2649 26138 2655 26172
rect 2689 26138 2695 26172
rect 2649 26099 2695 26138
rect 2649 26065 2655 26099
rect 2689 26065 2695 26099
rect 2649 26026 2695 26065
rect 2649 25992 2655 26026
rect 2689 25992 2695 26026
rect 2649 25953 2695 25992
rect 2649 25919 2655 25953
rect 2689 25919 2695 25953
rect 2649 25880 2695 25919
rect 2649 25846 2655 25880
rect 2689 25846 2695 25880
rect 2649 25807 2695 25846
rect 2649 25773 2655 25807
rect 2689 25773 2695 25807
tri 2459 25734 2461 25736 sw
tri 2647 25734 2649 25736 se
rect 2649 25734 2695 25773
rect 2885 26172 3076 26184
rect 2885 26138 2891 26172
rect 2925 26146 3076 26172
rect 2925 26138 3036 26146
rect 2885 26112 3036 26138
rect 3070 26112 3076 26146
rect 2885 26099 3076 26112
rect 2885 26065 2891 26099
rect 2925 26074 3076 26099
rect 2925 26065 3036 26074
rect 2885 26040 3036 26065
rect 3070 26040 3076 26074
rect 2885 26026 3076 26040
rect 2885 25992 2891 26026
rect 2925 26002 3076 26026
rect 2925 25992 3036 26002
rect 2885 25968 3036 25992
rect 3070 25968 3076 26002
rect 2885 25953 3076 25968
rect 2885 25919 2891 25953
rect 2925 25930 3076 25953
rect 2925 25919 3036 25930
rect 2885 25896 3036 25919
rect 3070 25896 3076 25930
rect 2885 25880 3076 25896
rect 2885 25846 2891 25880
rect 2925 25858 3076 25880
rect 2925 25846 3036 25858
rect 2885 25824 3036 25846
rect 3070 25824 3076 25858
rect 2885 25807 3076 25824
rect 2885 25773 2891 25807
rect 2925 25786 3076 25807
rect 2925 25773 3036 25786
rect 2885 25752 3036 25773
rect 3070 25752 3076 25786
tri 2695 25734 2697 25736 sw
tri 2883 25734 2885 25736 se
rect 2885 25734 3076 25752
rect 420 25733 531 25734
rect 380 25700 531 25733
rect 565 25702 573 25734
tri 573 25702 605 25734 sw
tri 727 25702 759 25734 se
rect 759 25702 767 25734
rect 565 25700 767 25702
rect 801 25702 809 25734
tri 809 25702 841 25734 sw
tri 963 25702 995 25734 se
rect 995 25702 1003 25734
rect 801 25700 1003 25702
rect 1037 25702 1045 25734
tri 1045 25702 1077 25734 sw
tri 1199 25702 1231 25734 se
rect 1231 25702 1239 25734
rect 1037 25700 1239 25702
rect 1273 25702 1281 25734
tri 1281 25702 1313 25734 sw
tri 1435 25702 1467 25734 se
rect 1467 25702 1475 25734
rect 1273 25700 1475 25702
rect 1509 25702 1517 25734
tri 1517 25702 1549 25734 sw
tri 1671 25702 1703 25734 se
rect 1703 25702 1711 25734
rect 1509 25700 1711 25702
rect 1745 25702 1753 25734
tri 1753 25702 1785 25734 sw
tri 1907 25702 1939 25734 se
rect 1939 25702 1947 25734
rect 1745 25700 1947 25702
rect 1981 25702 1989 25734
tri 1989 25702 2021 25734 sw
tri 2143 25702 2175 25734 se
rect 2175 25702 2183 25734
rect 1981 25700 2183 25702
rect 2217 25702 2225 25734
tri 2225 25702 2257 25734 sw
tri 2379 25702 2411 25734 se
rect 2411 25702 2419 25734
rect 2217 25700 2419 25702
rect 2453 25702 2461 25734
tri 2461 25702 2493 25734 sw
tri 2615 25702 2647 25734 se
rect 2647 25702 2655 25734
rect 2453 25700 2655 25702
rect 2689 25702 2697 25734
tri 2697 25702 2729 25734 sw
tri 2851 25702 2883 25734 se
rect 2883 25702 2891 25734
rect 2689 25700 2891 25702
rect 2925 25714 3076 25734
rect 2925 25700 3036 25714
rect 380 25695 3036 25700
rect 380 25661 386 25695
rect 420 25680 3036 25695
rect 3070 25680 3076 25714
rect 420 25679 3076 25680
rect 420 25661 697 25679
rect 380 25627 531 25661
rect 565 25627 697 25661
rect 749 25627 765 25679
rect 817 25627 833 25679
rect 885 25627 901 25679
rect 953 25627 969 25679
rect 1021 25661 1037 25679
rect 1089 25627 1105 25679
rect 1157 25627 1173 25679
rect 1225 25661 1241 25679
rect 1293 25661 2097 25679
rect 1225 25627 1239 25661
rect 1293 25627 1475 25661
rect 1509 25627 1711 25661
rect 1745 25627 1947 25661
rect 1981 25627 2097 25661
rect 2149 25627 2165 25679
rect 2217 25627 2233 25679
rect 2285 25627 2301 25679
rect 2353 25627 2369 25679
rect 2421 25661 2437 25679
rect 2489 25627 2505 25679
rect 2557 25627 2573 25679
rect 2625 25627 2641 25679
rect 2693 25661 3076 25679
rect 2693 25627 2891 25661
rect 2925 25642 3076 25661
rect 2925 25627 3036 25642
rect 380 25623 3036 25627
rect 380 25589 386 25623
rect 420 25615 3036 25623
rect 420 25589 697 25615
rect 380 25588 697 25589
rect 380 25554 531 25588
rect 565 25563 697 25588
rect 749 25563 765 25615
rect 817 25563 833 25615
rect 885 25563 901 25615
rect 953 25563 969 25615
rect 1021 25588 1037 25615
rect 1089 25563 1105 25615
rect 1157 25563 1173 25615
rect 1225 25588 1241 25615
rect 1293 25588 2097 25615
rect 1225 25563 1239 25588
rect 1293 25563 1475 25588
rect 565 25554 767 25563
rect 801 25554 1003 25563
rect 1037 25554 1239 25563
rect 1273 25554 1475 25563
rect 1509 25554 1711 25588
rect 1745 25554 1947 25588
rect 1981 25563 2097 25588
rect 2149 25563 2165 25615
rect 2217 25563 2233 25615
rect 2285 25563 2301 25615
rect 2353 25563 2369 25615
rect 2421 25588 2437 25615
rect 2489 25563 2505 25615
rect 2557 25563 2573 25615
rect 2625 25563 2641 25615
rect 2693 25608 3036 25615
rect 3070 25608 3076 25642
rect 2693 25588 3076 25608
rect 2693 25563 2891 25588
rect 1981 25554 2183 25563
rect 2217 25554 2419 25563
rect 2453 25554 2655 25563
rect 2689 25554 2891 25563
rect 2925 25570 3076 25588
rect 2925 25554 3036 25570
rect 380 25551 3036 25554
rect 380 25517 386 25551
rect 420 25517 697 25551
rect 380 25515 697 25517
rect 380 25481 531 25515
rect 565 25499 697 25515
rect 749 25499 765 25551
rect 817 25499 833 25551
rect 885 25499 901 25551
rect 953 25499 969 25551
rect 1021 25515 1037 25551
rect 1089 25499 1105 25551
rect 1157 25499 1173 25551
rect 1225 25515 1241 25551
rect 1293 25515 2097 25551
rect 1225 25499 1239 25515
rect 1293 25499 1475 25515
rect 565 25487 767 25499
rect 801 25487 1003 25499
rect 1037 25487 1239 25499
rect 1273 25487 1475 25499
rect 565 25481 697 25487
rect 380 25479 697 25481
rect 380 25445 386 25479
rect 420 25445 697 25479
rect 380 25442 697 25445
rect 380 25408 531 25442
rect 565 25435 697 25442
rect 749 25435 765 25487
rect 817 25435 833 25487
rect 885 25435 901 25487
rect 953 25435 969 25487
rect 1021 25442 1037 25481
rect 1089 25435 1105 25487
rect 1157 25435 1173 25487
rect 1225 25481 1239 25487
rect 1293 25481 1475 25487
rect 1509 25481 1711 25515
rect 1745 25481 1947 25515
rect 1981 25499 2097 25515
rect 2149 25499 2165 25551
rect 2217 25499 2233 25551
rect 2285 25499 2301 25551
rect 2353 25499 2369 25551
rect 2421 25515 2437 25551
rect 2489 25499 2505 25551
rect 2557 25499 2573 25551
rect 2625 25499 2641 25551
rect 2693 25536 3036 25551
rect 3070 25536 3076 25570
rect 2693 25515 3076 25536
rect 2693 25499 2891 25515
rect 1981 25487 2183 25499
rect 2217 25487 2419 25499
rect 2453 25487 2655 25499
rect 2689 25487 2891 25499
rect 1981 25481 2097 25487
rect 1225 25442 1241 25481
rect 1293 25442 2097 25481
rect 1225 25435 1239 25442
rect 1293 25435 1475 25442
rect 565 25423 767 25435
rect 801 25423 1003 25435
rect 1037 25423 1239 25435
rect 1273 25423 1475 25435
rect 565 25408 697 25423
rect 380 25407 697 25408
rect 380 25373 386 25407
rect 420 25373 697 25407
rect 380 25371 697 25373
rect 749 25371 765 25423
rect 817 25371 833 25423
rect 885 25371 901 25423
rect 953 25371 969 25423
rect 1021 25371 1037 25408
rect 1089 25371 1105 25423
rect 1157 25371 1173 25423
rect 1225 25408 1239 25423
rect 1293 25408 1475 25423
rect 1509 25408 1711 25442
rect 1745 25408 1947 25442
rect 1981 25435 2097 25442
rect 2149 25435 2165 25487
rect 2217 25435 2233 25487
rect 2285 25435 2301 25487
rect 2353 25435 2369 25487
rect 2421 25442 2437 25481
rect 2489 25435 2505 25487
rect 2557 25435 2573 25487
rect 2625 25435 2641 25487
rect 2693 25481 2891 25487
rect 2925 25498 3076 25515
rect 2925 25481 3036 25498
rect 2693 25464 3036 25481
rect 3070 25464 3076 25498
rect 2693 25442 3076 25464
rect 2693 25435 2891 25442
rect 1981 25423 2183 25435
rect 2217 25423 2419 25435
rect 2453 25423 2655 25435
rect 2689 25423 2891 25435
rect 1981 25408 2097 25423
rect 1225 25371 1241 25408
rect 1293 25371 2097 25408
rect 2149 25371 2165 25423
rect 2217 25371 2233 25423
rect 2285 25371 2301 25423
rect 2353 25371 2369 25423
rect 2421 25371 2437 25408
rect 2489 25371 2505 25423
rect 2557 25371 2573 25423
rect 2625 25371 2641 25423
rect 2693 25408 2891 25423
rect 2925 25426 3076 25442
rect 2925 25408 3036 25426
rect 2693 25392 3036 25408
rect 3070 25392 3076 25426
rect 2693 25371 3076 25392
rect 380 25369 3076 25371
rect 380 25335 531 25369
rect 565 25359 767 25369
rect 801 25359 1003 25369
rect 1037 25359 1239 25369
rect 1273 25359 1475 25369
rect 565 25335 697 25359
rect 380 25301 386 25335
rect 420 25307 697 25335
rect 749 25307 765 25359
rect 817 25307 833 25359
rect 885 25307 901 25359
rect 953 25307 969 25359
rect 1021 25307 1037 25335
rect 1089 25307 1105 25359
rect 1157 25307 1173 25359
rect 1225 25335 1239 25359
rect 1293 25335 1475 25359
rect 1509 25335 1711 25369
rect 1745 25335 1947 25369
rect 1981 25359 2183 25369
rect 2217 25359 2419 25369
rect 2453 25359 2655 25369
rect 2689 25359 2891 25369
rect 1981 25335 2097 25359
rect 1225 25307 1241 25335
rect 1293 25307 2097 25335
rect 2149 25307 2165 25359
rect 2217 25307 2233 25359
rect 2285 25307 2301 25359
rect 2353 25307 2369 25359
rect 2421 25307 2437 25335
rect 2489 25307 2505 25359
rect 2557 25307 2573 25359
rect 2625 25307 2641 25359
rect 2693 25335 2891 25359
rect 2925 25354 3076 25369
rect 2925 25335 3036 25354
rect 2693 25320 3036 25335
rect 3070 25320 3076 25354
rect 2693 25307 3076 25320
rect 420 25301 3076 25307
rect 380 25296 3076 25301
rect 380 25263 531 25296
rect 380 25229 386 25263
rect 420 25262 531 25263
rect 565 25295 767 25296
rect 801 25295 1003 25296
rect 1037 25295 1239 25296
rect 1273 25295 1475 25296
rect 565 25262 697 25295
rect 420 25243 697 25262
rect 749 25243 765 25295
rect 817 25243 833 25295
rect 885 25243 901 25295
rect 953 25243 969 25295
rect 1021 25243 1037 25262
rect 1089 25243 1105 25295
rect 1157 25243 1173 25295
rect 1225 25262 1239 25295
rect 1293 25262 1475 25295
rect 1509 25262 1711 25296
rect 1745 25262 1947 25296
rect 1981 25295 2183 25296
rect 2217 25295 2419 25296
rect 2453 25295 2655 25296
rect 2689 25295 2891 25296
rect 1981 25262 2097 25295
rect 1225 25243 1241 25262
rect 1293 25243 2097 25262
rect 2149 25243 2165 25295
rect 2217 25243 2233 25295
rect 2285 25243 2301 25295
rect 2353 25243 2369 25295
rect 2421 25243 2437 25262
rect 2489 25243 2505 25295
rect 2557 25243 2573 25295
rect 2625 25243 2641 25295
rect 2693 25262 2891 25295
rect 2925 25282 3076 25296
rect 2925 25262 3036 25282
rect 2693 25248 3036 25262
rect 3070 25248 3076 25282
rect 2693 25243 3076 25248
rect 420 25231 3076 25243
rect 420 25229 697 25231
rect 380 25222 697 25229
rect 380 25191 531 25222
rect 380 25157 386 25191
rect 420 25188 531 25191
rect 565 25188 697 25222
rect 420 25179 697 25188
rect 749 25179 765 25231
rect 817 25179 833 25231
rect 885 25179 901 25231
rect 953 25179 969 25231
rect 1021 25222 1037 25231
rect 1021 25179 1037 25188
rect 1089 25179 1105 25231
rect 1157 25179 1173 25231
rect 1225 25222 1241 25231
rect 1293 25222 2097 25231
rect 1225 25188 1239 25222
rect 1293 25188 1475 25222
rect 1509 25188 1711 25222
rect 1745 25188 1947 25222
rect 1981 25188 2097 25222
rect 1225 25179 1241 25188
rect 1293 25179 2097 25188
rect 2149 25179 2165 25231
rect 2217 25179 2233 25231
rect 2285 25179 2301 25231
rect 2353 25179 2369 25231
rect 2421 25222 2437 25231
rect 2421 25179 2437 25188
rect 2489 25179 2505 25231
rect 2557 25179 2573 25231
rect 2625 25179 2641 25231
rect 2693 25222 3076 25231
rect 2693 25188 2891 25222
rect 2925 25210 3076 25222
rect 2925 25188 3036 25210
rect 2693 25179 3036 25188
rect 420 25176 3036 25179
rect 3070 25176 3076 25210
rect 420 25167 3076 25176
rect 420 25157 697 25167
rect 380 25148 697 25157
rect 380 25119 531 25148
rect 380 25085 386 25119
rect 420 25114 531 25119
rect 565 25115 697 25148
rect 749 25115 765 25167
rect 817 25115 833 25167
rect 885 25115 901 25167
rect 953 25115 969 25167
rect 1021 25148 1037 25167
rect 1089 25115 1105 25167
rect 1157 25115 1173 25167
rect 1225 25148 1241 25167
rect 1293 25148 2097 25167
rect 1225 25115 1239 25148
rect 1293 25115 1475 25148
rect 565 25114 767 25115
rect 801 25114 1003 25115
rect 1037 25114 1239 25115
rect 1273 25114 1475 25115
rect 1509 25114 1711 25148
rect 1745 25114 1947 25148
rect 1981 25115 2097 25148
rect 2149 25115 2165 25167
rect 2217 25115 2233 25167
rect 2285 25115 2301 25167
rect 2353 25115 2369 25167
rect 2421 25148 2437 25167
rect 2489 25115 2505 25167
rect 2557 25115 2573 25167
rect 2625 25115 2641 25167
rect 2693 25148 3076 25167
rect 2693 25115 2891 25148
rect 1981 25114 2183 25115
rect 2217 25114 2419 25115
rect 2453 25114 2655 25115
rect 2689 25114 2891 25115
rect 2925 25138 3076 25148
rect 2925 25114 3036 25138
rect 420 25104 3036 25114
rect 3070 25104 3076 25138
rect 420 25103 3076 25104
rect 420 25085 697 25103
rect 380 25074 697 25085
rect 380 25047 531 25074
rect 380 25013 386 25047
rect 420 25040 531 25047
rect 565 25051 697 25074
rect 749 25051 765 25103
rect 817 25051 833 25103
rect 885 25051 901 25103
rect 953 25051 969 25103
rect 1021 25074 1037 25103
rect 1089 25051 1105 25103
rect 1157 25051 1173 25103
rect 1225 25074 1241 25103
rect 1293 25074 2097 25103
rect 1225 25051 1239 25074
rect 1293 25051 1475 25074
rect 565 25040 767 25051
rect 801 25040 1003 25051
rect 1037 25040 1239 25051
rect 1273 25040 1475 25051
rect 1509 25040 1711 25074
rect 1745 25040 1947 25074
rect 1981 25051 2097 25074
rect 2149 25051 2165 25103
rect 2217 25051 2233 25103
rect 2285 25051 2301 25103
rect 2353 25051 2369 25103
rect 2421 25074 2437 25103
rect 2489 25051 2505 25103
rect 2557 25051 2573 25103
rect 2625 25051 2641 25103
rect 2693 25074 3076 25103
rect 2693 25051 2891 25074
rect 1981 25040 2183 25051
rect 2217 25040 2419 25051
rect 2453 25040 2655 25051
rect 2689 25040 2891 25051
rect 2925 25066 3076 25074
rect 2925 25040 3036 25066
rect 420 25039 3036 25040
rect 420 25013 697 25039
rect 380 25000 697 25013
rect 380 24975 531 25000
rect 380 24941 386 24975
rect 420 24966 531 24975
rect 565 24987 697 25000
rect 749 24987 765 25039
rect 817 24987 833 25039
rect 885 24987 901 25039
rect 953 24987 969 25039
rect 1021 25000 1037 25039
rect 1089 24987 1105 25039
rect 1157 24987 1173 25039
rect 1225 25000 1241 25039
rect 1293 25000 2097 25039
rect 1225 24987 1239 25000
rect 1293 24987 1475 25000
rect 565 24975 767 24987
rect 801 24975 1003 24987
rect 1037 24975 1239 24987
rect 1273 24975 1475 24987
rect 565 24966 697 24975
rect 420 24941 697 24966
rect 380 24926 697 24941
rect 380 24903 531 24926
rect 380 24869 386 24903
rect 420 24892 531 24903
rect 565 24923 697 24926
rect 749 24923 765 24975
rect 817 24923 833 24975
rect 885 24923 901 24975
rect 953 24923 969 24975
rect 1021 24926 1037 24966
rect 1089 24923 1105 24975
rect 1157 24923 1173 24975
rect 1225 24966 1239 24975
rect 1293 24966 1475 24975
rect 1509 24966 1711 25000
rect 1745 24966 1947 25000
rect 1981 24987 2097 25000
rect 2149 24987 2165 25039
rect 2217 24987 2233 25039
rect 2285 24987 2301 25039
rect 2353 24987 2369 25039
rect 2421 25000 2437 25039
rect 2489 24987 2505 25039
rect 2557 24987 2573 25039
rect 2625 24987 2641 25039
rect 2693 25032 3036 25039
rect 3070 25032 3076 25066
rect 2693 25000 3076 25032
rect 2693 24987 2891 25000
rect 1981 24975 2183 24987
rect 2217 24975 2419 24987
rect 2453 24975 2655 24987
rect 2689 24975 2891 24987
rect 1981 24966 2097 24975
rect 1225 24926 1241 24966
rect 1293 24926 2097 24966
rect 1225 24923 1239 24926
rect 1293 24923 1475 24926
rect 565 24911 767 24923
rect 801 24911 1003 24923
rect 1037 24911 1239 24923
rect 1273 24911 1475 24923
rect 565 24892 697 24911
rect 420 24869 697 24892
rect 380 24859 697 24869
rect 749 24859 765 24911
rect 817 24859 833 24911
rect 885 24859 901 24911
rect 953 24859 969 24911
rect 1021 24859 1037 24892
rect 1089 24859 1105 24911
rect 1157 24859 1173 24911
rect 1225 24892 1239 24911
rect 1293 24892 1475 24911
rect 1509 24892 1711 24926
rect 1745 24892 1947 24926
rect 1981 24923 2097 24926
rect 2149 24923 2165 24975
rect 2217 24923 2233 24975
rect 2285 24923 2301 24975
rect 2353 24923 2369 24975
rect 2421 24926 2437 24966
rect 2489 24923 2505 24975
rect 2557 24923 2573 24975
rect 2625 24923 2641 24975
rect 2693 24966 2891 24975
rect 2925 24994 3076 25000
rect 2925 24966 3036 24994
rect 2693 24960 3036 24966
rect 3070 24960 3076 24994
rect 2693 24926 3076 24960
rect 2693 24923 2891 24926
rect 1981 24911 2183 24923
rect 2217 24911 2419 24923
rect 2453 24911 2655 24923
rect 2689 24911 2891 24923
rect 1981 24892 2097 24911
rect 1225 24859 1241 24892
rect 1293 24859 2097 24892
rect 2149 24859 2165 24911
rect 2217 24859 2233 24911
rect 2285 24859 2301 24911
rect 2353 24859 2369 24911
rect 2421 24859 2437 24892
rect 2489 24859 2505 24911
rect 2557 24859 2573 24911
rect 2625 24859 2641 24911
rect 2693 24892 2891 24911
rect 2925 24922 3076 24926
rect 2925 24892 3036 24922
rect 2693 24888 3036 24892
rect 3070 24888 3076 24922
rect 2693 24859 3076 24888
rect 380 24852 3076 24859
rect 380 24831 531 24852
rect 380 24797 386 24831
rect 420 24818 531 24831
rect 565 24847 767 24852
rect 801 24847 1003 24852
rect 1037 24847 1239 24852
rect 1273 24847 1475 24852
rect 565 24818 697 24847
rect 420 24797 697 24818
rect 380 24795 697 24797
rect 749 24795 765 24847
rect 817 24795 833 24847
rect 885 24795 901 24847
rect 953 24795 969 24847
rect 1021 24795 1037 24818
rect 1089 24795 1105 24847
rect 1157 24795 1173 24847
rect 1225 24818 1239 24847
rect 1293 24818 1475 24847
rect 1509 24818 1711 24852
rect 1745 24818 1947 24852
rect 1981 24847 2183 24852
rect 2217 24847 2419 24852
rect 2453 24847 2655 24852
rect 2689 24847 2891 24852
rect 1981 24818 2097 24847
rect 1225 24795 1241 24818
rect 1293 24795 2097 24818
rect 2149 24795 2165 24847
rect 2217 24795 2233 24847
rect 2285 24795 2301 24847
rect 2353 24795 2369 24847
rect 2421 24795 2437 24818
rect 2489 24795 2505 24847
rect 2557 24795 2573 24847
rect 2625 24795 2641 24847
rect 2693 24818 2891 24847
rect 2925 24850 3076 24852
rect 2925 24818 3036 24850
rect 2693 24816 3036 24818
rect 3070 24816 3076 24850
rect 2693 24795 3076 24816
rect 380 24783 3076 24795
rect 380 24778 697 24783
rect 380 24759 531 24778
rect 380 24725 386 24759
rect 420 24744 531 24759
rect 565 24744 697 24778
rect 420 24731 697 24744
rect 749 24731 765 24783
rect 817 24731 833 24783
rect 885 24731 901 24783
rect 953 24731 969 24783
rect 1021 24778 1037 24783
rect 1021 24731 1037 24744
rect 1089 24731 1105 24783
rect 1157 24731 1173 24783
rect 1225 24778 1241 24783
rect 1293 24778 2097 24783
rect 1225 24744 1239 24778
rect 1293 24744 1475 24778
rect 1509 24744 1711 24778
rect 1745 24744 1947 24778
rect 1981 24744 2097 24778
rect 1225 24731 1241 24744
rect 1293 24731 2097 24744
rect 2149 24731 2165 24783
rect 2217 24731 2233 24783
rect 2285 24731 2301 24783
rect 2353 24731 2369 24783
rect 2421 24778 2437 24783
rect 2421 24731 2437 24744
rect 2489 24731 2505 24783
rect 2557 24731 2573 24783
rect 2625 24731 2641 24783
rect 2693 24778 3076 24783
rect 2693 24744 2891 24778
rect 2925 24744 3036 24778
rect 3070 24744 3076 24778
rect 2693 24731 3076 24744
rect 420 24725 3076 24731
rect 380 24706 3076 24725
rect 380 24704 3036 24706
rect 380 24687 531 24704
rect 380 24653 386 24687
rect 420 24670 531 24687
rect 565 24702 767 24704
rect 565 24687 590 24702
tri 590 24687 605 24702 nw
tri 727 24687 742 24702 ne
rect 742 24687 767 24702
rect 565 24670 573 24687
tri 573 24670 590 24687 nw
tri 742 24670 759 24687 ne
rect 759 24670 767 24687
rect 801 24702 1003 24704
rect 801 24687 826 24702
tri 826 24687 841 24702 nw
tri 963 24687 978 24702 ne
rect 978 24687 1003 24702
rect 801 24670 809 24687
tri 809 24670 826 24687 nw
tri 978 24670 995 24687 ne
rect 995 24670 1003 24687
rect 1037 24702 1239 24704
rect 1037 24687 1062 24702
tri 1062 24687 1077 24702 nw
tri 1199 24687 1214 24702 ne
rect 1214 24687 1239 24702
rect 1037 24670 1045 24687
tri 1045 24670 1062 24687 nw
tri 1214 24670 1231 24687 ne
rect 1231 24670 1239 24687
rect 1273 24702 1475 24704
rect 1273 24687 1298 24702
tri 1298 24687 1313 24702 nw
tri 1435 24687 1450 24702 ne
rect 1450 24687 1475 24702
rect 1273 24670 1281 24687
tri 1281 24670 1298 24687 nw
tri 1450 24670 1467 24687 ne
rect 1467 24670 1475 24687
rect 1509 24702 1711 24704
rect 1509 24687 1534 24702
tri 1534 24687 1549 24702 nw
tri 1671 24687 1686 24702 ne
rect 1686 24687 1711 24702
rect 1509 24670 1517 24687
tri 1517 24670 1534 24687 nw
tri 1686 24670 1703 24687 ne
rect 1703 24670 1711 24687
rect 1745 24702 1947 24704
rect 1745 24687 1770 24702
tri 1770 24687 1785 24702 nw
tri 1907 24687 1922 24702 ne
rect 1922 24687 1947 24702
rect 1745 24670 1753 24687
tri 1753 24670 1770 24687 nw
tri 1922 24670 1939 24687 ne
rect 1939 24670 1947 24687
rect 1981 24702 2183 24704
rect 1981 24687 2006 24702
tri 2006 24687 2021 24702 nw
tri 2143 24687 2158 24702 ne
rect 2158 24687 2183 24702
rect 1981 24670 1989 24687
tri 1989 24670 2006 24687 nw
tri 2158 24670 2175 24687 ne
rect 2175 24670 2183 24687
rect 2217 24702 2419 24704
rect 2217 24687 2242 24702
tri 2242 24687 2257 24702 nw
tri 2379 24687 2394 24702 ne
rect 2394 24687 2419 24702
rect 2217 24670 2225 24687
tri 2225 24670 2242 24687 nw
tri 2394 24670 2411 24687 ne
rect 2411 24670 2419 24687
rect 2453 24702 2655 24704
rect 2453 24687 2478 24702
tri 2478 24687 2493 24702 nw
tri 2615 24687 2630 24702 ne
rect 2630 24687 2655 24702
rect 2453 24670 2461 24687
tri 2461 24670 2478 24687 nw
tri 2630 24670 2647 24687 ne
rect 2647 24670 2655 24687
rect 2689 24702 2891 24704
rect 2689 24687 2714 24702
tri 2714 24687 2729 24702 nw
tri 2851 24687 2866 24702 ne
rect 2866 24687 2891 24702
rect 2689 24670 2697 24687
tri 2697 24670 2714 24687 nw
tri 2866 24670 2883 24687 ne
rect 2883 24670 2891 24687
rect 2925 24672 3036 24704
rect 3070 24672 3076 24706
rect 2925 24670 3076 24672
rect 420 24653 571 24670
tri 571 24668 573 24670 nw
tri 759 24668 761 24670 ne
rect 380 24630 571 24653
rect 380 24615 531 24630
rect 380 24581 386 24615
rect 420 24596 531 24615
rect 565 24596 571 24630
rect 420 24581 571 24596
rect 380 24556 571 24581
rect 380 24543 531 24556
rect 380 24509 386 24543
rect 420 24522 531 24543
rect 565 24522 571 24556
rect 420 24509 571 24522
rect 380 24482 571 24509
rect 380 24471 531 24482
rect 380 24437 386 24471
rect 420 24448 531 24471
rect 565 24448 571 24482
rect 420 24437 571 24448
rect 380 24408 571 24437
rect 380 24399 531 24408
rect 380 24365 386 24399
rect 420 24374 531 24399
rect 565 24374 571 24408
rect 420 24365 571 24374
rect 380 24334 571 24365
rect 380 24327 531 24334
rect 380 24293 386 24327
rect 420 24300 531 24327
rect 565 24300 571 24334
rect 420 24293 571 24300
rect 380 24260 571 24293
rect 380 24255 531 24260
rect 380 24221 386 24255
rect 420 24226 531 24255
rect 565 24226 571 24260
rect 420 24221 571 24226
rect 380 24183 571 24221
rect 761 24630 807 24670
tri 807 24668 809 24670 nw
tri 995 24668 997 24670 ne
rect 761 24596 767 24630
rect 801 24596 807 24630
rect 761 24556 807 24596
rect 761 24522 767 24556
rect 801 24522 807 24556
rect 761 24482 807 24522
rect 761 24448 767 24482
rect 801 24448 807 24482
rect 761 24408 807 24448
rect 761 24374 767 24408
rect 801 24374 807 24408
rect 761 24334 807 24374
rect 761 24300 767 24334
rect 801 24300 807 24334
rect 761 24260 807 24300
rect 761 24226 767 24260
rect 801 24226 807 24260
rect 761 24214 807 24226
rect 997 24630 1043 24670
tri 1043 24668 1045 24670 nw
tri 1231 24668 1233 24670 ne
rect 997 24596 1003 24630
rect 1037 24596 1043 24630
rect 997 24556 1043 24596
rect 997 24522 1003 24556
rect 1037 24522 1043 24556
rect 997 24482 1043 24522
rect 997 24448 1003 24482
rect 1037 24448 1043 24482
rect 997 24408 1043 24448
rect 997 24374 1003 24408
rect 1037 24374 1043 24408
rect 997 24334 1043 24374
rect 997 24300 1003 24334
rect 1037 24300 1043 24334
rect 997 24260 1043 24300
rect 997 24226 1003 24260
rect 1037 24226 1043 24260
rect 997 24214 1043 24226
rect 1233 24630 1279 24670
tri 1279 24668 1281 24670 nw
tri 1467 24668 1469 24670 ne
rect 1233 24596 1239 24630
rect 1273 24596 1279 24630
rect 1233 24556 1279 24596
rect 1233 24522 1239 24556
rect 1273 24522 1279 24556
rect 1233 24482 1279 24522
rect 1233 24448 1239 24482
rect 1273 24448 1279 24482
rect 1233 24408 1279 24448
rect 1233 24374 1239 24408
rect 1273 24374 1279 24408
rect 1233 24334 1279 24374
rect 1233 24300 1239 24334
rect 1273 24300 1279 24334
rect 1233 24260 1279 24300
rect 1233 24226 1239 24260
rect 1273 24226 1279 24260
rect 1233 24214 1279 24226
rect 1469 24630 1515 24670
tri 1515 24668 1517 24670 nw
tri 1703 24668 1705 24670 ne
rect 1469 24596 1475 24630
rect 1509 24596 1515 24630
rect 1469 24556 1515 24596
rect 1469 24522 1475 24556
rect 1509 24522 1515 24556
rect 1469 24482 1515 24522
rect 1469 24448 1475 24482
rect 1509 24448 1515 24482
rect 1469 24408 1515 24448
rect 1469 24374 1475 24408
rect 1509 24374 1515 24408
rect 1469 24334 1515 24374
rect 1469 24300 1475 24334
rect 1509 24300 1515 24334
rect 1469 24260 1515 24300
rect 1469 24226 1475 24260
rect 1509 24226 1515 24260
rect 1469 24214 1515 24226
rect 1705 24630 1751 24670
tri 1751 24668 1753 24670 nw
tri 1939 24668 1941 24670 ne
rect 1705 24596 1711 24630
rect 1745 24596 1751 24630
rect 1705 24556 1751 24596
rect 1705 24522 1711 24556
rect 1745 24522 1751 24556
rect 1705 24482 1751 24522
rect 1705 24448 1711 24482
rect 1745 24448 1751 24482
rect 1705 24408 1751 24448
rect 1705 24374 1711 24408
rect 1745 24374 1751 24408
rect 1705 24334 1751 24374
rect 1705 24300 1711 24334
rect 1745 24300 1751 24334
rect 1705 24260 1751 24300
rect 1705 24226 1711 24260
rect 1745 24226 1751 24260
rect 1705 24214 1751 24226
rect 1941 24630 1987 24670
tri 1987 24668 1989 24670 nw
tri 2175 24668 2177 24670 ne
rect 1941 24596 1947 24630
rect 1981 24596 1987 24630
rect 1941 24556 1987 24596
rect 1941 24522 1947 24556
rect 1981 24522 1987 24556
rect 1941 24482 1987 24522
rect 1941 24448 1947 24482
rect 1981 24448 1987 24482
rect 1941 24408 1987 24448
rect 1941 24374 1947 24408
rect 1981 24374 1987 24408
rect 1941 24334 1987 24374
rect 1941 24300 1947 24334
rect 1981 24300 1987 24334
rect 1941 24260 1987 24300
rect 1941 24226 1947 24260
rect 1981 24226 1987 24260
rect 1941 24214 1987 24226
rect 2177 24630 2223 24670
tri 2223 24668 2225 24670 nw
tri 2411 24668 2413 24670 ne
rect 2177 24596 2183 24630
rect 2217 24596 2223 24630
rect 2177 24556 2223 24596
rect 2177 24522 2183 24556
rect 2217 24522 2223 24556
rect 2177 24482 2223 24522
rect 2177 24448 2183 24482
rect 2217 24448 2223 24482
rect 2177 24408 2223 24448
rect 2177 24374 2183 24408
rect 2217 24374 2223 24408
rect 2177 24334 2223 24374
rect 2177 24300 2183 24334
rect 2217 24300 2223 24334
rect 2177 24260 2223 24300
rect 2177 24226 2183 24260
rect 2217 24226 2223 24260
rect 2177 24214 2223 24226
rect 2413 24630 2459 24670
tri 2459 24668 2461 24670 nw
tri 2647 24668 2649 24670 ne
rect 2413 24596 2419 24630
rect 2453 24596 2459 24630
rect 2413 24556 2459 24596
rect 2413 24522 2419 24556
rect 2453 24522 2459 24556
rect 2413 24482 2459 24522
rect 2413 24448 2419 24482
rect 2453 24448 2459 24482
rect 2413 24408 2459 24448
rect 2413 24374 2419 24408
rect 2453 24374 2459 24408
rect 2413 24334 2459 24374
rect 2413 24300 2419 24334
rect 2453 24300 2459 24334
rect 2413 24260 2459 24300
rect 2413 24226 2419 24260
rect 2453 24226 2459 24260
rect 2413 24214 2459 24226
rect 2649 24630 2695 24670
tri 2695 24668 2697 24670 nw
tri 2883 24668 2885 24670 ne
rect 2649 24596 2655 24630
rect 2689 24596 2695 24630
rect 2649 24556 2695 24596
rect 2649 24522 2655 24556
rect 2689 24522 2695 24556
rect 2649 24482 2695 24522
rect 2649 24448 2655 24482
rect 2689 24448 2695 24482
rect 2649 24408 2695 24448
rect 2649 24374 2655 24408
rect 2689 24374 2695 24408
rect 2649 24334 2695 24374
rect 2649 24300 2655 24334
rect 2689 24300 2695 24334
rect 2649 24260 2695 24300
rect 2649 24226 2655 24260
rect 2689 24226 2695 24260
rect 2649 24214 2695 24226
rect 2885 24634 3076 24670
rect 2885 24630 3036 24634
rect 2885 24596 2891 24630
rect 2925 24600 3036 24630
rect 3070 24600 3076 24634
rect 2925 24596 3076 24600
rect 2885 24562 3076 24596
rect 2885 24556 3036 24562
rect 2885 24522 2891 24556
rect 2925 24528 3036 24556
rect 3070 24528 3076 24562
rect 2925 24522 3076 24528
rect 2885 24490 3076 24522
rect 2885 24482 3036 24490
rect 2885 24448 2891 24482
rect 2925 24456 3036 24482
rect 3070 24456 3076 24490
rect 2925 24448 3076 24456
rect 2885 24418 3076 24448
rect 2885 24408 3036 24418
rect 2885 24374 2891 24408
rect 2925 24384 3036 24408
rect 3070 24384 3076 24418
rect 2925 24374 3076 24384
rect 2885 24346 3076 24374
rect 2885 24334 3036 24346
rect 2885 24300 2891 24334
rect 2925 24312 3036 24334
rect 3070 24312 3076 24346
rect 2925 24300 3076 24312
rect 2885 24274 3076 24300
rect 2885 24260 3036 24274
rect 2885 24226 2891 24260
rect 2925 24240 3036 24260
rect 3070 24240 3076 24274
rect 2925 24226 3076 24240
rect 380 24149 386 24183
rect 420 24149 571 24183
rect 2885 24202 3076 24226
rect 2885 24168 3036 24202
rect 3070 24168 3076 24202
rect 380 24111 571 24149
rect 380 24077 386 24111
rect 420 24077 571 24111
rect 613 24144 1501 24153
rect 1553 24144 1569 24153
rect 1621 24144 1636 24153
rect 1688 24144 1703 24153
rect 1755 24144 1770 24153
rect 1822 24144 1837 24153
rect 1889 24144 2830 24153
rect 613 24110 625 24144
rect 659 24110 700 24144
rect 734 24110 775 24144
rect 809 24110 850 24144
rect 884 24110 925 24144
rect 959 24110 1000 24144
rect 1034 24110 1075 24144
rect 1109 24110 1150 24144
rect 1184 24110 1225 24144
rect 1259 24110 1300 24144
rect 1334 24110 1375 24144
rect 1409 24110 1450 24144
rect 1484 24110 1501 24144
rect 1559 24110 1569 24144
rect 1634 24110 1636 24144
rect 1889 24110 1896 24144
rect 1930 24110 1970 24144
rect 2004 24110 2044 24144
rect 2078 24110 2118 24144
rect 2152 24110 2192 24144
rect 2226 24110 2266 24144
rect 2300 24110 2340 24144
rect 2374 24110 2414 24144
rect 2448 24110 2488 24144
rect 2522 24110 2562 24144
rect 2596 24110 2636 24144
rect 2670 24110 2710 24144
rect 2744 24110 2784 24144
rect 2818 24110 2830 24144
rect 613 24101 1501 24110
rect 1553 24101 1569 24110
rect 1621 24101 1636 24110
rect 1688 24101 1703 24110
rect 1755 24101 1770 24110
rect 1822 24101 1837 24110
rect 1889 24101 2830 24110
rect 2885 24130 3076 24168
rect 380 24039 571 24077
rect 2885 24096 3036 24130
rect 3070 24096 3076 24130
rect 2885 24058 3076 24096
rect 380 24005 386 24039
rect 420 24028 571 24039
rect 420 24005 531 24028
rect 380 23994 531 24005
rect 565 23994 571 24028
rect 380 23967 571 23994
rect 380 23933 386 23967
rect 420 23955 571 23967
rect 420 23933 531 23955
rect 380 23921 531 23933
rect 565 23921 571 23955
rect 380 23895 571 23921
rect 380 23861 386 23895
rect 420 23882 571 23895
rect 420 23861 531 23882
rect 380 23848 531 23861
rect 565 23848 571 23882
rect 380 23823 571 23848
rect 380 23789 386 23823
rect 420 23809 571 23823
rect 420 23789 531 23809
rect 380 23775 531 23789
rect 565 23775 571 23809
rect 380 23751 571 23775
rect 380 23717 386 23751
rect 420 23736 571 23751
rect 420 23717 531 23736
rect 380 23702 531 23717
rect 565 23702 571 23736
rect 380 23679 571 23702
rect 380 23645 386 23679
rect 420 23663 571 23679
rect 420 23645 531 23663
rect 380 23629 531 23645
rect 565 23629 571 23663
rect 380 23607 571 23629
rect 380 23573 386 23607
rect 420 23590 571 23607
rect 761 24028 807 24040
rect 761 23994 767 24028
rect 801 23994 807 24028
rect 761 23955 807 23994
rect 761 23921 767 23955
rect 801 23921 807 23955
rect 761 23882 807 23921
rect 761 23848 767 23882
rect 801 23848 807 23882
rect 761 23809 807 23848
rect 761 23775 767 23809
rect 801 23775 807 23809
rect 761 23736 807 23775
rect 761 23702 767 23736
rect 801 23702 807 23736
rect 761 23663 807 23702
rect 761 23629 767 23663
rect 801 23629 807 23663
rect 761 23590 807 23629
rect 997 24028 1043 24040
rect 997 23994 1003 24028
rect 1037 23994 1043 24028
rect 997 23955 1043 23994
rect 997 23921 1003 23955
rect 1037 23921 1043 23955
rect 997 23882 1043 23921
rect 997 23848 1003 23882
rect 1037 23848 1043 23882
rect 997 23809 1043 23848
rect 997 23775 1003 23809
rect 1037 23775 1043 23809
rect 997 23736 1043 23775
rect 997 23702 1003 23736
rect 1037 23702 1043 23736
rect 997 23663 1043 23702
rect 997 23629 1003 23663
rect 1037 23629 1043 23663
rect 997 23590 1043 23629
rect 1233 24028 1279 24040
rect 1233 23994 1239 24028
rect 1273 23994 1279 24028
rect 1233 23955 1279 23994
rect 1233 23921 1239 23955
rect 1273 23921 1279 23955
rect 1233 23882 1279 23921
rect 1233 23848 1239 23882
rect 1273 23848 1279 23882
rect 1233 23809 1279 23848
rect 1233 23775 1239 23809
rect 1273 23775 1279 23809
rect 1233 23736 1279 23775
rect 1233 23702 1239 23736
rect 1273 23702 1279 23736
rect 1233 23663 1279 23702
rect 1233 23629 1239 23663
rect 1273 23629 1279 23663
rect 1233 23590 1279 23629
rect 1469 24028 1515 24040
rect 1469 23994 1475 24028
rect 1509 23994 1515 24028
rect 1469 23955 1515 23994
rect 1469 23921 1475 23955
rect 1509 23921 1515 23955
rect 1469 23882 1515 23921
rect 1469 23848 1475 23882
rect 1509 23848 1515 23882
rect 1469 23809 1515 23848
rect 1469 23775 1475 23809
rect 1509 23775 1515 23809
rect 1469 23736 1515 23775
rect 1469 23702 1475 23736
rect 1509 23702 1515 23736
rect 1469 23663 1515 23702
rect 1469 23629 1475 23663
rect 1509 23629 1515 23663
rect 1469 23590 1515 23629
rect 1705 24028 1751 24040
rect 1705 23994 1711 24028
rect 1745 23994 1751 24028
rect 1705 23955 1751 23994
rect 1705 23921 1711 23955
rect 1745 23921 1751 23955
rect 1705 23882 1751 23921
rect 1705 23848 1711 23882
rect 1745 23848 1751 23882
rect 1705 23809 1751 23848
rect 1705 23775 1711 23809
rect 1745 23775 1751 23809
rect 1705 23736 1751 23775
rect 1705 23702 1711 23736
rect 1745 23702 1751 23736
rect 1705 23663 1751 23702
rect 1705 23629 1711 23663
rect 1745 23629 1751 23663
rect 1705 23590 1751 23629
rect 1941 24028 1987 24040
rect 1941 23994 1947 24028
rect 1981 23994 1987 24028
rect 1941 23955 1987 23994
rect 1941 23921 1947 23955
rect 1981 23921 1987 23955
rect 1941 23882 1987 23921
rect 1941 23848 1947 23882
rect 1981 23848 1987 23882
rect 1941 23809 1987 23848
rect 1941 23775 1947 23809
rect 1981 23775 1987 23809
rect 1941 23736 1987 23775
rect 1941 23702 1947 23736
rect 1981 23702 1987 23736
rect 1941 23663 1987 23702
rect 1941 23629 1947 23663
rect 1981 23629 1987 23663
rect 1941 23590 1987 23629
rect 2177 24028 2223 24040
rect 2177 23994 2183 24028
rect 2217 23994 2223 24028
rect 2177 23955 2223 23994
rect 2177 23921 2183 23955
rect 2217 23921 2223 23955
rect 2177 23882 2223 23921
rect 2177 23848 2183 23882
rect 2217 23848 2223 23882
rect 2177 23809 2223 23848
rect 2177 23775 2183 23809
rect 2217 23775 2223 23809
rect 2177 23736 2223 23775
rect 2177 23702 2183 23736
rect 2217 23702 2223 23736
rect 2177 23663 2223 23702
rect 2177 23629 2183 23663
rect 2217 23629 2223 23663
rect 2177 23590 2223 23629
rect 2413 24028 2459 24040
rect 2413 23994 2419 24028
rect 2453 23994 2459 24028
rect 2413 23955 2459 23994
rect 2413 23921 2419 23955
rect 2453 23921 2459 23955
rect 2413 23882 2459 23921
rect 2413 23848 2419 23882
rect 2453 23848 2459 23882
rect 2413 23809 2459 23848
rect 2413 23775 2419 23809
rect 2453 23775 2459 23809
rect 2413 23736 2459 23775
rect 2413 23702 2419 23736
rect 2453 23702 2459 23736
rect 2413 23663 2459 23702
rect 2413 23629 2419 23663
rect 2453 23629 2459 23663
rect 2413 23590 2459 23629
rect 2649 24028 2695 24040
rect 2649 23994 2655 24028
rect 2689 23994 2695 24028
rect 2649 23955 2695 23994
rect 2649 23921 2655 23955
rect 2689 23921 2695 23955
rect 2649 23882 2695 23921
rect 2649 23848 2655 23882
rect 2689 23848 2695 23882
rect 2649 23809 2695 23848
rect 2649 23775 2655 23809
rect 2689 23775 2695 23809
rect 2649 23736 2695 23775
rect 2649 23702 2655 23736
rect 2689 23702 2695 23736
rect 2649 23663 2695 23702
rect 2649 23629 2655 23663
rect 2689 23629 2695 23663
rect 2649 23590 2695 23629
rect 2885 24028 3036 24058
rect 2885 23994 2891 24028
rect 2925 24024 3036 24028
rect 3070 24024 3076 24058
rect 2925 23994 3076 24024
rect 2885 23986 3076 23994
rect 2885 23955 3036 23986
rect 2885 23921 2891 23955
rect 2925 23952 3036 23955
rect 3070 23952 3076 23986
rect 2925 23921 3076 23952
rect 2885 23914 3076 23921
rect 2885 23882 3036 23914
rect 2885 23848 2891 23882
rect 2925 23880 3036 23882
rect 3070 23880 3076 23914
rect 2925 23848 3076 23880
rect 2885 23842 3076 23848
rect 2885 23809 3036 23842
rect 2885 23775 2891 23809
rect 2925 23808 3036 23809
rect 3070 23808 3076 23842
rect 2925 23775 3076 23808
rect 2885 23770 3076 23775
rect 2885 23736 3036 23770
rect 3070 23736 3076 23770
rect 2885 23702 2891 23736
rect 2925 23702 3076 23736
rect 2885 23698 3076 23702
rect 2885 23664 3036 23698
rect 3070 23664 3076 23698
rect 2885 23663 3076 23664
rect 2885 23629 2891 23663
rect 2925 23629 3076 23663
rect 2885 23626 3076 23629
rect 2885 23592 3036 23626
rect 3070 23592 3076 23626
rect 2885 23590 3076 23592
rect 420 23573 531 23590
rect 380 23556 531 23573
rect 565 23556 571 23590
tri 571 23556 605 23590 sw
tri 727 23556 761 23590 se
rect 761 23556 767 23590
rect 801 23556 807 23590
tri 807 23556 841 23590 sw
tri 963 23556 997 23590 se
rect 997 23556 1003 23590
rect 1037 23556 1043 23590
tri 1043 23556 1077 23590 sw
tri 1199 23556 1233 23590 se
rect 1233 23556 1239 23590
rect 1273 23556 1279 23590
tri 1279 23556 1313 23590 sw
tri 1435 23556 1469 23590 se
rect 1469 23556 1475 23590
rect 1509 23556 1515 23590
tri 1515 23556 1549 23590 sw
tri 1671 23556 1705 23590 se
rect 1705 23556 1711 23590
rect 1745 23556 1751 23590
tri 1751 23556 1785 23590 sw
tri 1907 23556 1941 23590 se
rect 1941 23556 1947 23590
rect 1981 23556 1987 23590
tri 1987 23556 2021 23590 sw
tri 2143 23556 2177 23590 se
rect 2177 23556 2183 23590
rect 2217 23556 2223 23590
tri 2223 23556 2257 23590 sw
tri 2379 23556 2413 23590 se
rect 2413 23556 2419 23590
rect 2453 23556 2459 23590
tri 2459 23556 2493 23590 sw
tri 2615 23556 2649 23590 se
rect 2649 23556 2655 23590
rect 2689 23556 2695 23590
tri 2695 23556 2729 23590 sw
tri 2851 23556 2885 23590 se
rect 2885 23556 2891 23590
rect 2925 23556 3076 23590
rect 380 23554 3076 23556
rect 380 23535 3036 23554
rect 380 23501 386 23535
rect 420 23531 3036 23535
rect 420 23517 697 23531
rect 420 23501 531 23517
rect 380 23483 531 23501
rect 565 23483 697 23517
rect 380 23479 697 23483
rect 749 23479 765 23531
rect 817 23479 833 23531
rect 885 23479 901 23531
rect 953 23479 969 23531
rect 1021 23517 1037 23531
rect 1021 23479 1037 23483
rect 1089 23479 1105 23531
rect 1157 23479 1173 23531
rect 1225 23517 1241 23531
rect 1293 23517 2097 23531
rect 1225 23483 1239 23517
rect 1293 23483 1475 23517
rect 1509 23483 1711 23517
rect 1745 23483 1947 23517
rect 1981 23483 2097 23517
rect 1225 23479 1241 23483
rect 1293 23479 2097 23483
rect 2149 23479 2165 23531
rect 2217 23479 2233 23531
rect 2285 23479 2301 23531
rect 2353 23479 2369 23531
rect 2421 23517 2437 23531
rect 2421 23479 2437 23483
rect 2489 23479 2505 23531
rect 2557 23479 2573 23531
rect 2625 23479 2641 23531
rect 2693 23520 3036 23531
rect 3070 23520 3076 23554
rect 2693 23517 3076 23520
rect 2693 23483 2891 23517
rect 2925 23483 3076 23517
rect 2693 23482 3076 23483
rect 2693 23479 3036 23482
rect 380 23467 3036 23479
rect 380 23463 697 23467
rect 380 23429 386 23463
rect 420 23444 697 23463
rect 420 23429 531 23444
rect 380 23410 531 23429
rect 565 23415 697 23444
rect 749 23415 765 23467
rect 817 23415 833 23467
rect 885 23415 901 23467
rect 953 23415 969 23467
rect 1021 23444 1037 23467
rect 1089 23415 1105 23467
rect 1157 23415 1173 23467
rect 1225 23444 1241 23467
rect 1293 23444 2097 23467
rect 1225 23415 1239 23444
rect 1293 23415 1475 23444
rect 565 23410 767 23415
rect 801 23410 1003 23415
rect 1037 23410 1239 23415
rect 1273 23410 1475 23415
rect 1509 23410 1711 23444
rect 1745 23410 1947 23444
rect 1981 23415 2097 23444
rect 2149 23415 2165 23467
rect 2217 23415 2233 23467
rect 2285 23415 2301 23467
rect 2353 23415 2369 23467
rect 2421 23444 2437 23467
rect 2489 23415 2505 23467
rect 2557 23415 2573 23467
rect 2625 23415 2641 23467
rect 2693 23448 3036 23467
rect 3070 23448 3076 23482
rect 2693 23444 3076 23448
rect 2693 23415 2891 23444
rect 1981 23410 2183 23415
rect 2217 23410 2419 23415
rect 2453 23410 2655 23415
rect 2689 23410 2891 23415
rect 2925 23410 3076 23444
rect 380 23403 3036 23410
rect 380 23391 697 23403
rect 380 23357 386 23391
rect 420 23371 697 23391
rect 420 23357 531 23371
rect 380 23337 531 23357
rect 565 23351 697 23371
rect 749 23351 765 23403
rect 817 23351 833 23403
rect 885 23351 901 23403
rect 953 23351 969 23403
rect 1021 23371 1037 23403
rect 1089 23351 1105 23403
rect 1157 23351 1173 23403
rect 1225 23371 1241 23403
rect 1293 23371 2097 23403
rect 1225 23351 1239 23371
rect 1293 23351 1475 23371
rect 565 23339 767 23351
rect 801 23339 1003 23351
rect 1037 23339 1239 23351
rect 1273 23339 1475 23351
rect 565 23337 697 23339
rect 380 23319 697 23337
rect 380 23285 386 23319
rect 420 23298 697 23319
rect 420 23285 531 23298
rect 380 23264 531 23285
rect 565 23287 697 23298
rect 749 23287 765 23339
rect 817 23287 833 23339
rect 885 23287 901 23339
rect 953 23287 969 23339
rect 1021 23298 1037 23337
rect 1089 23287 1105 23339
rect 1157 23287 1173 23339
rect 1225 23337 1239 23339
rect 1293 23337 1475 23339
rect 1509 23337 1711 23371
rect 1745 23337 1947 23371
rect 1981 23351 2097 23371
rect 2149 23351 2165 23403
rect 2217 23351 2233 23403
rect 2285 23351 2301 23403
rect 2353 23351 2369 23403
rect 2421 23371 2437 23403
rect 2489 23351 2505 23403
rect 2557 23351 2573 23403
rect 2625 23351 2641 23403
rect 2693 23376 3036 23403
rect 3070 23376 3076 23410
rect 2693 23371 3076 23376
rect 2693 23351 2891 23371
rect 1981 23339 2183 23351
rect 2217 23339 2419 23351
rect 2453 23339 2655 23351
rect 2689 23339 2891 23351
rect 1981 23337 2097 23339
rect 1225 23298 1241 23337
rect 1293 23298 2097 23337
rect 1225 23287 1239 23298
rect 1293 23287 1475 23298
rect 565 23275 767 23287
rect 801 23275 1003 23287
rect 1037 23275 1239 23287
rect 1273 23275 1475 23287
rect 565 23264 697 23275
rect 380 23247 697 23264
rect 380 23213 386 23247
rect 420 23225 697 23247
rect 420 23213 531 23225
rect 380 23191 531 23213
rect 565 23223 697 23225
rect 749 23223 765 23275
rect 817 23223 833 23275
rect 885 23223 901 23275
rect 953 23223 969 23275
rect 1021 23225 1037 23264
rect 1089 23223 1105 23275
rect 1157 23223 1173 23275
rect 1225 23264 1239 23275
rect 1293 23264 1475 23275
rect 1509 23264 1711 23298
rect 1745 23264 1947 23298
rect 1981 23287 2097 23298
rect 2149 23287 2165 23339
rect 2217 23287 2233 23339
rect 2285 23287 2301 23339
rect 2353 23287 2369 23339
rect 2421 23298 2437 23337
rect 2489 23287 2505 23339
rect 2557 23287 2573 23339
rect 2625 23287 2641 23339
rect 2693 23337 2891 23339
rect 2925 23338 3076 23371
rect 2925 23337 3036 23338
rect 2693 23304 3036 23337
rect 3070 23304 3076 23338
rect 2693 23298 3076 23304
rect 2693 23287 2891 23298
rect 1981 23275 2183 23287
rect 2217 23275 2419 23287
rect 2453 23275 2655 23287
rect 2689 23275 2891 23287
rect 1981 23264 2097 23275
rect 1225 23225 1241 23264
rect 1293 23225 2097 23264
rect 1225 23223 1239 23225
rect 1293 23223 1475 23225
rect 565 23211 767 23223
rect 801 23211 1003 23223
rect 1037 23211 1239 23223
rect 1273 23211 1475 23223
rect 565 23191 697 23211
rect 380 23175 697 23191
rect 380 23141 386 23175
rect 420 23159 697 23175
rect 749 23159 765 23211
rect 817 23159 833 23211
rect 885 23159 901 23211
rect 953 23159 969 23211
rect 1021 23159 1037 23191
rect 1089 23159 1105 23211
rect 1157 23159 1173 23211
rect 1225 23191 1239 23211
rect 1293 23191 1475 23211
rect 1509 23191 1711 23225
rect 1745 23191 1947 23225
rect 1981 23223 2097 23225
rect 2149 23223 2165 23275
rect 2217 23223 2233 23275
rect 2285 23223 2301 23275
rect 2353 23223 2369 23275
rect 2421 23225 2437 23264
rect 2489 23223 2505 23275
rect 2557 23223 2573 23275
rect 2625 23223 2641 23275
rect 2693 23264 2891 23275
rect 2925 23266 3076 23298
rect 2925 23264 3036 23266
rect 2693 23232 3036 23264
rect 3070 23232 3076 23266
rect 2693 23225 3076 23232
rect 2693 23223 2891 23225
rect 1981 23211 2183 23223
rect 2217 23211 2419 23223
rect 2453 23211 2655 23223
rect 2689 23211 2891 23223
rect 1981 23191 2097 23211
rect 1225 23159 1241 23191
rect 1293 23159 2097 23191
rect 2149 23159 2165 23211
rect 2217 23159 2233 23211
rect 2285 23159 2301 23211
rect 2353 23159 2369 23211
rect 2421 23159 2437 23191
rect 2489 23159 2505 23211
rect 2557 23159 2573 23211
rect 2625 23159 2641 23211
rect 2693 23191 2891 23211
rect 2925 23194 3076 23225
rect 2925 23191 3036 23194
rect 2693 23160 3036 23191
rect 3070 23160 3076 23194
rect 2693 23159 3076 23160
rect 420 23152 3076 23159
rect 420 23141 531 23152
rect 380 23118 531 23141
rect 565 23147 767 23152
rect 801 23147 1003 23152
rect 1037 23147 1239 23152
rect 1273 23147 1475 23152
rect 565 23118 697 23147
rect 380 23103 697 23118
rect 380 23069 386 23103
rect 420 23095 697 23103
rect 749 23095 765 23147
rect 817 23095 833 23147
rect 885 23095 901 23147
rect 953 23095 969 23147
rect 1021 23095 1037 23118
rect 1089 23095 1105 23147
rect 1157 23095 1173 23147
rect 1225 23118 1239 23147
rect 1293 23118 1475 23147
rect 1509 23118 1711 23152
rect 1745 23118 1947 23152
rect 1981 23147 2183 23152
rect 2217 23147 2419 23152
rect 2453 23147 2655 23152
rect 2689 23147 2891 23152
rect 1981 23118 2097 23147
rect 1225 23095 1241 23118
rect 1293 23095 2097 23118
rect 2149 23095 2165 23147
rect 2217 23095 2233 23147
rect 2285 23095 2301 23147
rect 2353 23095 2369 23147
rect 2421 23095 2437 23118
rect 2489 23095 2505 23147
rect 2557 23095 2573 23147
rect 2625 23095 2641 23147
rect 2693 23118 2891 23147
rect 2925 23122 3076 23152
rect 2925 23118 3036 23122
rect 2693 23095 3036 23118
rect 420 23088 3036 23095
rect 3070 23088 3076 23122
rect 420 23083 3076 23088
rect 420 23078 697 23083
rect 420 23069 531 23078
rect 380 23044 531 23069
rect 565 23044 697 23078
rect 380 23031 697 23044
rect 749 23031 765 23083
rect 817 23031 833 23083
rect 885 23031 901 23083
rect 953 23031 969 23083
rect 1021 23078 1037 23083
rect 1021 23031 1037 23044
rect 1089 23031 1105 23083
rect 1157 23031 1173 23083
rect 1225 23078 1241 23083
rect 1293 23078 2097 23083
rect 1225 23044 1239 23078
rect 1293 23044 1475 23078
rect 1509 23044 1711 23078
rect 1745 23044 1947 23078
rect 1981 23044 2097 23078
rect 1225 23031 1241 23044
rect 1293 23031 2097 23044
rect 2149 23031 2165 23083
rect 2217 23031 2233 23083
rect 2285 23031 2301 23083
rect 2353 23031 2369 23083
rect 2421 23078 2437 23083
rect 2421 23031 2437 23044
rect 2489 23031 2505 23083
rect 2557 23031 2573 23083
rect 2625 23031 2641 23083
rect 2693 23078 3076 23083
rect 2693 23044 2891 23078
rect 2925 23050 3076 23078
rect 2925 23044 3036 23050
rect 2693 23031 3036 23044
rect 380 22997 386 23031
rect 420 23019 3036 23031
rect 420 23004 697 23019
rect 420 22997 531 23004
rect 380 22970 531 22997
rect 565 22970 697 23004
rect 380 22967 697 22970
rect 749 22967 765 23019
rect 817 22967 833 23019
rect 885 22967 901 23019
rect 953 22967 969 23019
rect 1021 23004 1037 23019
rect 1021 22967 1037 22970
rect 1089 22967 1105 23019
rect 1157 22967 1173 23019
rect 1225 23004 1241 23019
rect 1293 23004 2097 23019
rect 1225 22970 1239 23004
rect 1293 22970 1475 23004
rect 1509 22970 1711 23004
rect 1745 22970 1947 23004
rect 1981 22970 2097 23004
rect 1225 22967 1241 22970
rect 1293 22967 2097 22970
rect 2149 22967 2165 23019
rect 2217 22967 2233 23019
rect 2285 22967 2301 23019
rect 2353 22967 2369 23019
rect 2421 23004 2437 23019
rect 2421 22967 2437 22970
rect 2489 22967 2505 23019
rect 2557 22967 2573 23019
rect 2625 22967 2641 23019
rect 2693 23016 3036 23019
rect 3070 23016 3076 23050
rect 2693 23004 3076 23016
rect 2693 22970 2891 23004
rect 2925 22978 3076 23004
rect 2925 22970 3036 22978
rect 2693 22967 3036 22970
rect 380 22959 3036 22967
rect 380 22925 386 22959
rect 420 22955 3036 22959
rect 420 22930 697 22955
rect 420 22925 531 22930
rect 380 22896 531 22925
rect 565 22903 697 22930
rect 749 22903 765 22955
rect 817 22903 833 22955
rect 885 22903 901 22955
rect 953 22903 969 22955
rect 1021 22930 1037 22955
rect 1089 22903 1105 22955
rect 1157 22903 1173 22955
rect 1225 22930 1241 22955
rect 1293 22930 2097 22955
rect 1225 22903 1239 22930
rect 1293 22903 1475 22930
rect 565 22896 767 22903
rect 801 22896 1003 22903
rect 1037 22896 1239 22903
rect 1273 22896 1475 22903
rect 1509 22896 1711 22930
rect 1745 22896 1947 22930
rect 1981 22903 2097 22930
rect 2149 22903 2165 22955
rect 2217 22903 2233 22955
rect 2285 22903 2301 22955
rect 2353 22903 2369 22955
rect 2421 22930 2437 22955
rect 2489 22903 2505 22955
rect 2557 22903 2573 22955
rect 2625 22903 2641 22955
rect 2693 22944 3036 22955
rect 3070 22944 3076 22978
rect 2693 22930 3076 22944
rect 2693 22903 2891 22930
rect 1981 22896 2183 22903
rect 2217 22896 2419 22903
rect 2453 22896 2655 22903
rect 2689 22896 2891 22903
rect 2925 22906 3076 22930
rect 2925 22896 3036 22906
rect 380 22891 3036 22896
rect 380 22887 697 22891
rect 380 22853 386 22887
rect 420 22856 697 22887
rect 420 22853 531 22856
rect 380 22822 531 22853
rect 565 22839 697 22856
rect 749 22839 765 22891
rect 817 22839 833 22891
rect 885 22839 901 22891
rect 953 22839 969 22891
rect 1021 22856 1037 22891
rect 1089 22839 1105 22891
rect 1157 22839 1173 22891
rect 1225 22856 1241 22891
rect 1293 22856 2097 22891
rect 1225 22839 1239 22856
rect 1293 22839 1475 22856
rect 565 22827 767 22839
rect 801 22827 1003 22839
rect 1037 22827 1239 22839
rect 1273 22827 1475 22839
rect 565 22822 697 22827
rect 380 22815 697 22822
rect 380 22781 386 22815
rect 420 22782 697 22815
rect 420 22781 531 22782
rect 380 22748 531 22781
rect 565 22775 697 22782
rect 749 22775 765 22827
rect 817 22775 833 22827
rect 885 22775 901 22827
rect 953 22775 969 22827
rect 1021 22782 1037 22822
rect 1089 22775 1105 22827
rect 1157 22775 1173 22827
rect 1225 22822 1239 22827
rect 1293 22822 1475 22827
rect 1509 22822 1711 22856
rect 1745 22822 1947 22856
rect 1981 22839 2097 22856
rect 2149 22839 2165 22891
rect 2217 22839 2233 22891
rect 2285 22839 2301 22891
rect 2353 22839 2369 22891
rect 2421 22856 2437 22891
rect 2489 22839 2505 22891
rect 2557 22839 2573 22891
rect 2625 22839 2641 22891
rect 2693 22872 3036 22891
rect 3070 22872 3076 22906
rect 2693 22856 3076 22872
rect 2693 22839 2891 22856
rect 1981 22827 2183 22839
rect 2217 22827 2419 22839
rect 2453 22827 2655 22839
rect 2689 22827 2891 22839
rect 1981 22822 2097 22827
rect 1225 22782 1241 22822
rect 1293 22782 2097 22822
rect 1225 22775 1239 22782
rect 1293 22775 1475 22782
rect 565 22763 767 22775
rect 801 22763 1003 22775
rect 1037 22763 1239 22775
rect 1273 22763 1475 22775
rect 565 22748 697 22763
rect 380 22743 697 22748
rect 380 22709 386 22743
rect 420 22711 697 22743
rect 749 22711 765 22763
rect 817 22711 833 22763
rect 885 22711 901 22763
rect 953 22711 969 22763
rect 1021 22711 1037 22748
rect 1089 22711 1105 22763
rect 1157 22711 1173 22763
rect 1225 22748 1239 22763
rect 1293 22748 1475 22763
rect 1509 22748 1711 22782
rect 1745 22748 1947 22782
rect 1981 22775 2097 22782
rect 2149 22775 2165 22827
rect 2217 22775 2233 22827
rect 2285 22775 2301 22827
rect 2353 22775 2369 22827
rect 2421 22782 2437 22822
rect 2489 22775 2505 22827
rect 2557 22775 2573 22827
rect 2625 22775 2641 22827
rect 2693 22822 2891 22827
rect 2925 22834 3076 22856
rect 2925 22822 3036 22834
rect 2693 22800 3036 22822
rect 3070 22800 3076 22834
rect 2693 22782 3076 22800
rect 2693 22775 2891 22782
rect 1981 22763 2183 22775
rect 2217 22763 2419 22775
rect 2453 22763 2655 22775
rect 2689 22763 2891 22775
rect 1981 22748 2097 22763
rect 1225 22711 1241 22748
rect 1293 22711 2097 22748
rect 2149 22711 2165 22763
rect 2217 22711 2233 22763
rect 2285 22711 2301 22763
rect 2353 22711 2369 22763
rect 2421 22711 2437 22748
rect 2489 22711 2505 22763
rect 2557 22711 2573 22763
rect 2625 22711 2641 22763
rect 2693 22748 2891 22763
rect 2925 22762 3076 22782
rect 2925 22748 3036 22762
rect 2693 22728 3036 22748
rect 3070 22728 3076 22762
rect 2693 22711 3076 22728
rect 420 22709 3076 22711
rect 380 22708 3076 22709
rect 380 22674 531 22708
rect 565 22699 767 22708
rect 801 22699 1003 22708
rect 1037 22699 1239 22708
rect 1273 22699 1475 22708
rect 565 22674 697 22699
rect 380 22671 697 22674
rect 380 22637 386 22671
rect 420 22647 697 22671
rect 749 22647 765 22699
rect 817 22647 833 22699
rect 885 22647 901 22699
rect 953 22647 969 22699
rect 1021 22647 1037 22674
rect 1089 22647 1105 22699
rect 1157 22647 1173 22699
rect 1225 22674 1239 22699
rect 1293 22674 1475 22699
rect 1509 22674 1711 22708
rect 1745 22674 1947 22708
rect 1981 22699 2183 22708
rect 2217 22699 2419 22708
rect 2453 22699 2655 22708
rect 2689 22699 2891 22708
rect 1981 22674 2097 22699
rect 1225 22647 1241 22674
rect 1293 22647 2097 22674
rect 2149 22647 2165 22699
rect 2217 22647 2233 22699
rect 2285 22647 2301 22699
rect 2353 22647 2369 22699
rect 2421 22647 2437 22674
rect 2489 22647 2505 22699
rect 2557 22647 2573 22699
rect 2625 22647 2641 22699
rect 2693 22674 2891 22699
rect 2925 22690 3076 22708
rect 2925 22674 3036 22690
rect 2693 22656 3036 22674
rect 3070 22656 3076 22690
rect 2693 22647 3076 22656
rect 420 22637 3076 22647
rect 380 22635 3076 22637
rect 380 22634 697 22635
rect 380 22600 531 22634
rect 565 22600 697 22634
rect 380 22599 697 22600
rect 380 22565 386 22599
rect 420 22583 697 22599
rect 749 22583 765 22635
rect 817 22583 833 22635
rect 885 22583 901 22635
rect 953 22583 969 22635
rect 1021 22634 1037 22635
rect 1021 22583 1037 22600
rect 1089 22583 1105 22635
rect 1157 22583 1173 22635
rect 1225 22634 1241 22635
rect 1293 22634 2097 22635
rect 1225 22600 1239 22634
rect 1293 22600 1475 22634
rect 1509 22600 1711 22634
rect 1745 22600 1947 22634
rect 1981 22600 2097 22634
rect 1225 22583 1241 22600
rect 1293 22583 2097 22600
rect 2149 22583 2165 22635
rect 2217 22583 2233 22635
rect 2285 22583 2301 22635
rect 2353 22583 2369 22635
rect 2421 22634 2437 22635
rect 2421 22583 2437 22600
rect 2489 22583 2505 22635
rect 2557 22583 2573 22635
rect 2625 22583 2641 22635
rect 2693 22634 3076 22635
rect 2693 22600 2891 22634
rect 2925 22618 3076 22634
rect 2925 22600 3036 22618
rect 2693 22584 3036 22600
rect 3070 22584 3076 22618
rect 2693 22583 3076 22584
rect 420 22565 3076 22583
rect 380 22560 3076 22565
rect 380 22527 531 22560
rect 380 22493 386 22527
rect 420 22526 531 22527
rect 565 22556 767 22560
rect 565 22526 575 22556
tri 575 22526 605 22556 nw
tri 727 22526 757 22556 ne
rect 757 22526 767 22556
rect 801 22556 1003 22560
rect 801 22526 811 22556
tri 811 22526 841 22556 nw
tri 963 22526 993 22556 ne
rect 993 22526 1003 22556
rect 1037 22556 1239 22560
rect 1037 22526 1047 22556
tri 1047 22526 1077 22556 nw
tri 1199 22526 1229 22556 ne
rect 1229 22526 1239 22556
rect 1273 22556 1475 22560
rect 1273 22526 1283 22556
tri 1283 22526 1313 22556 nw
tri 1435 22526 1465 22556 ne
rect 1465 22526 1475 22556
rect 1509 22556 1711 22560
rect 1509 22526 1519 22556
tri 1519 22526 1549 22556 nw
tri 1671 22526 1701 22556 ne
rect 1701 22526 1711 22556
rect 1745 22556 1947 22560
rect 1745 22526 1755 22556
tri 1755 22526 1785 22556 nw
tri 1907 22526 1937 22556 ne
rect 1937 22526 1947 22556
rect 1981 22556 2183 22560
rect 1981 22526 1991 22556
tri 1991 22526 2021 22556 nw
tri 2143 22526 2173 22556 ne
rect 2173 22526 2183 22556
rect 2217 22556 2419 22560
rect 2217 22526 2227 22556
tri 2227 22526 2257 22556 nw
tri 2379 22526 2409 22556 ne
rect 2409 22526 2419 22556
rect 2453 22556 2655 22560
rect 2453 22526 2463 22556
tri 2463 22526 2493 22556 nw
tri 2615 22526 2645 22556 ne
rect 2645 22526 2655 22556
rect 2689 22556 2891 22560
rect 2689 22526 2699 22556
tri 2699 22526 2729 22556 nw
tri 2851 22526 2881 22556 ne
rect 2881 22526 2891 22556
rect 2925 22546 3076 22560
rect 2925 22526 3036 22546
rect 420 22493 571 22526
tri 571 22522 575 22526 nw
tri 757 22522 761 22526 ne
rect 380 22486 571 22493
rect 380 22455 531 22486
rect 380 22421 386 22455
rect 420 22452 531 22455
rect 565 22452 571 22486
rect 420 22421 571 22452
rect 380 22412 571 22421
rect 380 22383 531 22412
rect 380 22349 386 22383
rect 420 22378 531 22383
rect 565 22378 571 22412
rect 420 22349 571 22378
rect 380 22338 571 22349
rect 380 22311 531 22338
rect 380 22277 386 22311
rect 420 22304 531 22311
rect 565 22304 571 22338
rect 420 22277 571 22304
rect 380 22264 571 22277
rect 380 22239 531 22264
rect 380 22205 386 22239
rect 420 22230 531 22239
rect 565 22230 571 22264
rect 420 22205 571 22230
rect 380 22190 571 22205
rect 380 22167 531 22190
rect 380 22133 386 22167
rect 420 22156 531 22167
rect 565 22156 571 22190
rect 420 22133 571 22156
rect 380 22116 571 22133
rect 380 22095 531 22116
rect 380 22061 386 22095
rect 420 22082 531 22095
rect 565 22082 571 22116
rect 420 22061 571 22082
rect 761 22486 807 22526
tri 807 22522 811 22526 nw
tri 993 22522 997 22526 ne
rect 761 22452 767 22486
rect 801 22452 807 22486
rect 761 22412 807 22452
rect 761 22378 767 22412
rect 801 22378 807 22412
rect 761 22338 807 22378
rect 761 22304 767 22338
rect 801 22304 807 22338
rect 761 22264 807 22304
rect 761 22230 767 22264
rect 801 22230 807 22264
rect 761 22190 807 22230
rect 761 22156 767 22190
rect 801 22156 807 22190
rect 761 22116 807 22156
rect 761 22082 767 22116
rect 801 22082 807 22116
rect 761 22070 807 22082
rect 997 22486 1043 22526
tri 1043 22522 1047 22526 nw
tri 1229 22522 1233 22526 ne
rect 997 22452 1003 22486
rect 1037 22452 1043 22486
rect 997 22412 1043 22452
rect 997 22378 1003 22412
rect 1037 22378 1043 22412
rect 997 22338 1043 22378
rect 997 22304 1003 22338
rect 1037 22304 1043 22338
rect 997 22264 1043 22304
rect 997 22230 1003 22264
rect 1037 22230 1043 22264
rect 997 22190 1043 22230
rect 997 22156 1003 22190
rect 1037 22156 1043 22190
rect 997 22116 1043 22156
rect 997 22082 1003 22116
rect 1037 22082 1043 22116
rect 997 22070 1043 22082
rect 1233 22486 1279 22526
tri 1279 22522 1283 22526 nw
tri 1465 22522 1469 22526 ne
rect 1233 22452 1239 22486
rect 1273 22452 1279 22486
rect 1233 22412 1279 22452
rect 1233 22378 1239 22412
rect 1273 22378 1279 22412
rect 1233 22338 1279 22378
rect 1233 22304 1239 22338
rect 1273 22304 1279 22338
rect 1233 22264 1279 22304
rect 1233 22230 1239 22264
rect 1273 22230 1279 22264
rect 1233 22190 1279 22230
rect 1233 22156 1239 22190
rect 1273 22156 1279 22190
rect 1233 22116 1279 22156
rect 1233 22082 1239 22116
rect 1273 22082 1279 22116
rect 1233 22070 1279 22082
rect 1469 22486 1515 22526
tri 1515 22522 1519 22526 nw
tri 1701 22522 1705 22526 ne
rect 1469 22452 1475 22486
rect 1509 22452 1515 22486
rect 1469 22412 1515 22452
rect 1469 22378 1475 22412
rect 1509 22378 1515 22412
rect 1469 22338 1515 22378
rect 1469 22304 1475 22338
rect 1509 22304 1515 22338
rect 1469 22264 1515 22304
rect 1469 22230 1475 22264
rect 1509 22230 1515 22264
rect 1469 22190 1515 22230
rect 1469 22156 1475 22190
rect 1509 22156 1515 22190
rect 1469 22116 1515 22156
rect 1469 22082 1475 22116
rect 1509 22082 1515 22116
rect 1469 22070 1515 22082
rect 1705 22486 1751 22526
tri 1751 22522 1755 22526 nw
tri 1937 22522 1941 22526 ne
rect 1705 22452 1711 22486
rect 1745 22452 1751 22486
rect 1705 22412 1751 22452
rect 1705 22378 1711 22412
rect 1745 22378 1751 22412
rect 1705 22338 1751 22378
rect 1705 22304 1711 22338
rect 1745 22304 1751 22338
rect 1705 22264 1751 22304
rect 1705 22230 1711 22264
rect 1745 22230 1751 22264
rect 1705 22190 1751 22230
rect 1705 22156 1711 22190
rect 1745 22156 1751 22190
rect 1705 22116 1751 22156
rect 1705 22082 1711 22116
rect 1745 22082 1751 22116
rect 1705 22070 1751 22082
rect 1941 22486 1987 22526
tri 1987 22522 1991 22526 nw
tri 2173 22522 2177 22526 ne
rect 1941 22452 1947 22486
rect 1981 22452 1987 22486
rect 1941 22412 1987 22452
rect 1941 22378 1947 22412
rect 1981 22378 1987 22412
rect 1941 22338 1987 22378
rect 1941 22304 1947 22338
rect 1981 22304 1987 22338
rect 1941 22264 1987 22304
rect 1941 22230 1947 22264
rect 1981 22230 1987 22264
rect 1941 22190 1987 22230
rect 1941 22156 1947 22190
rect 1981 22156 1987 22190
rect 1941 22116 1987 22156
rect 1941 22082 1947 22116
rect 1981 22082 1987 22116
rect 1941 22070 1987 22082
rect 2177 22486 2223 22526
tri 2223 22522 2227 22526 nw
tri 2409 22522 2413 22526 ne
rect 2177 22452 2183 22486
rect 2217 22452 2223 22486
rect 2177 22412 2223 22452
rect 2177 22378 2183 22412
rect 2217 22378 2223 22412
rect 2177 22338 2223 22378
rect 2177 22304 2183 22338
rect 2217 22304 2223 22338
rect 2177 22264 2223 22304
rect 2177 22230 2183 22264
rect 2217 22230 2223 22264
rect 2177 22190 2223 22230
rect 2177 22156 2183 22190
rect 2217 22156 2223 22190
rect 2177 22116 2223 22156
rect 2177 22082 2183 22116
rect 2217 22082 2223 22116
rect 2177 22070 2223 22082
rect 2413 22486 2459 22526
tri 2459 22522 2463 22526 nw
tri 2645 22522 2649 22526 ne
rect 2413 22452 2419 22486
rect 2453 22452 2459 22486
rect 2413 22412 2459 22452
rect 2413 22378 2419 22412
rect 2453 22378 2459 22412
rect 2413 22338 2459 22378
rect 2413 22304 2419 22338
rect 2453 22304 2459 22338
rect 2413 22264 2459 22304
rect 2413 22230 2419 22264
rect 2453 22230 2459 22264
rect 2413 22190 2459 22230
rect 2413 22156 2419 22190
rect 2453 22156 2459 22190
rect 2413 22116 2459 22156
rect 2413 22082 2419 22116
rect 2453 22082 2459 22116
rect 2413 22070 2459 22082
rect 2649 22486 2695 22526
tri 2695 22522 2699 22526 nw
tri 2881 22522 2885 22526 ne
rect 2649 22452 2655 22486
rect 2689 22452 2695 22486
rect 2649 22412 2695 22452
rect 2649 22378 2655 22412
rect 2689 22378 2695 22412
rect 2649 22338 2695 22378
rect 2649 22304 2655 22338
rect 2689 22304 2695 22338
rect 2649 22264 2695 22304
rect 2649 22230 2655 22264
rect 2689 22230 2695 22264
rect 2649 22190 2695 22230
rect 2649 22156 2655 22190
rect 2689 22156 2695 22190
rect 2649 22116 2695 22156
rect 2649 22082 2655 22116
rect 2689 22082 2695 22116
rect 2649 22070 2695 22082
rect 2885 22512 3036 22526
rect 3070 22512 3076 22546
rect 2885 22486 3076 22512
rect 2885 22452 2891 22486
rect 2925 22474 3076 22486
rect 2925 22452 3036 22474
rect 2885 22440 3036 22452
rect 3070 22440 3076 22474
rect 2885 22412 3076 22440
rect 2885 22378 2891 22412
rect 2925 22402 3076 22412
rect 2925 22378 3036 22402
rect 2885 22368 3036 22378
rect 3070 22368 3076 22402
rect 2885 22338 3076 22368
rect 2885 22304 2891 22338
rect 2925 22330 3076 22338
rect 2925 22304 3036 22330
rect 2885 22296 3036 22304
rect 3070 22296 3076 22330
rect 2885 22264 3076 22296
rect 2885 22230 2891 22264
rect 2925 22258 3076 22264
rect 2925 22230 3036 22258
rect 2885 22224 3036 22230
rect 3070 22224 3076 22258
rect 2885 22190 3076 22224
rect 2885 22156 2891 22190
rect 2925 22186 3076 22190
rect 2925 22156 3036 22186
rect 2885 22152 3036 22156
rect 3070 22152 3076 22186
rect 2885 22116 3076 22152
rect 2885 22082 2891 22116
rect 2925 22114 3076 22116
rect 2925 22082 3036 22114
rect 2885 22080 3036 22082
rect 3070 22080 3076 22114
rect 380 22023 571 22061
rect 2885 22042 3076 22080
rect 380 21989 386 22023
rect 420 21989 571 22023
rect 380 21951 571 21989
rect 613 22014 1501 22023
rect 1553 22014 1569 22023
rect 1621 22014 1636 22023
rect 1688 22014 1703 22023
rect 1755 22014 1770 22023
rect 1822 22014 1837 22023
rect 1889 22014 2830 22023
rect 613 21980 625 22014
rect 659 21980 700 22014
rect 734 21980 775 22014
rect 809 21980 850 22014
rect 884 21980 925 22014
rect 959 21980 1000 22014
rect 1034 21980 1075 22014
rect 1109 21980 1150 22014
rect 1184 21980 1225 22014
rect 1259 21980 1300 22014
rect 1334 21980 1375 22014
rect 1409 21980 1450 22014
rect 1484 21980 1501 22014
rect 1559 21980 1569 22014
rect 1634 21980 1636 22014
rect 1889 21980 1896 22014
rect 1930 21980 1970 22014
rect 2004 21980 2044 22014
rect 2078 21980 2118 22014
rect 2152 21980 2192 22014
rect 2226 21980 2266 22014
rect 2300 21980 2340 22014
rect 2374 21980 2414 22014
rect 2448 21980 2488 22014
rect 2522 21980 2562 22014
rect 2596 21980 2636 22014
rect 2670 21980 2710 22014
rect 2744 21980 2784 22014
rect 2818 21980 2830 22014
rect 613 21971 1501 21980
rect 1553 21971 1569 21980
rect 1621 21971 1636 21980
rect 1688 21971 1703 21980
rect 1755 21971 1770 21980
rect 1822 21971 1837 21980
rect 1889 21971 2830 21980
rect 2885 22008 3036 22042
rect 3070 22008 3076 22042
rect 380 21917 386 21951
rect 420 21917 571 21951
rect 2885 21970 3076 22008
rect 2885 21936 3036 21970
rect 3070 21936 3076 21970
rect 380 21912 571 21917
rect 380 21879 531 21912
rect 380 21845 386 21879
rect 420 21878 531 21879
rect 565 21878 571 21912
rect 420 21845 571 21878
rect 380 21839 571 21845
rect 380 21807 531 21839
rect 380 21773 386 21807
rect 420 21805 531 21807
rect 565 21805 571 21839
rect 420 21773 571 21805
rect 380 21766 571 21773
rect 380 21735 531 21766
rect 380 21701 386 21735
rect 420 21732 531 21735
rect 565 21732 571 21766
rect 420 21701 571 21732
rect 380 21693 571 21701
rect 380 21663 531 21693
rect 380 21629 386 21663
rect 420 21659 531 21663
rect 565 21659 571 21693
rect 420 21629 571 21659
rect 380 21620 571 21629
rect 380 21591 531 21620
rect 380 21557 386 21591
rect 420 21586 531 21591
rect 565 21586 571 21620
rect 420 21557 571 21586
rect 380 21547 571 21557
rect 380 21519 531 21547
rect 380 21485 386 21519
rect 420 21513 531 21519
rect 565 21513 571 21547
rect 420 21485 571 21513
rect 380 21474 571 21485
rect 380 21447 531 21474
rect 380 21413 386 21447
rect 420 21440 531 21447
rect 565 21440 571 21474
rect 420 21413 571 21440
rect 761 21912 807 21924
rect 761 21878 767 21912
rect 801 21878 807 21912
rect 761 21839 807 21878
rect 761 21805 767 21839
rect 801 21805 807 21839
rect 761 21766 807 21805
rect 761 21732 767 21766
rect 801 21732 807 21766
rect 761 21693 807 21732
rect 761 21659 767 21693
rect 801 21659 807 21693
rect 761 21620 807 21659
rect 761 21586 767 21620
rect 801 21586 807 21620
rect 761 21547 807 21586
rect 761 21513 767 21547
rect 801 21513 807 21547
rect 761 21474 807 21513
rect 761 21440 767 21474
rect 801 21440 807 21474
rect 380 21408 571 21413
tri 571 21408 583 21420 sw
tri 749 21408 761 21420 se
rect 761 21408 807 21440
rect 997 21912 1043 21924
rect 997 21878 1003 21912
rect 1037 21878 1043 21912
rect 997 21839 1043 21878
rect 997 21805 1003 21839
rect 1037 21805 1043 21839
rect 997 21766 1043 21805
rect 997 21732 1003 21766
rect 1037 21732 1043 21766
rect 997 21693 1043 21732
rect 997 21659 1003 21693
rect 1037 21659 1043 21693
rect 997 21620 1043 21659
rect 997 21586 1003 21620
rect 1037 21586 1043 21620
rect 997 21547 1043 21586
rect 997 21513 1003 21547
rect 1037 21513 1043 21547
rect 997 21474 1043 21513
rect 997 21440 1003 21474
rect 1037 21440 1043 21474
tri 807 21408 819 21420 sw
tri 985 21408 997 21420 se
rect 997 21408 1043 21440
rect 1233 21912 1279 21924
rect 1233 21878 1239 21912
rect 1273 21878 1279 21912
rect 1233 21839 1279 21878
rect 1233 21805 1239 21839
rect 1273 21805 1279 21839
rect 1233 21766 1279 21805
rect 1233 21732 1239 21766
rect 1273 21732 1279 21766
rect 1233 21693 1279 21732
rect 1233 21659 1239 21693
rect 1273 21659 1279 21693
rect 1233 21620 1279 21659
rect 1233 21586 1239 21620
rect 1273 21586 1279 21620
rect 1233 21547 1279 21586
rect 1233 21513 1239 21547
rect 1273 21513 1279 21547
rect 1233 21474 1279 21513
rect 1233 21440 1239 21474
rect 1273 21440 1279 21474
tri 1043 21408 1055 21420 sw
tri 1221 21408 1233 21420 se
rect 1233 21408 1279 21440
rect 1469 21912 1515 21924
rect 1469 21878 1475 21912
rect 1509 21878 1515 21912
rect 1469 21839 1515 21878
rect 1469 21805 1475 21839
rect 1509 21805 1515 21839
rect 1469 21766 1515 21805
rect 1469 21732 1475 21766
rect 1509 21732 1515 21766
rect 1469 21693 1515 21732
rect 1469 21659 1475 21693
rect 1509 21659 1515 21693
rect 1469 21620 1515 21659
rect 1469 21586 1475 21620
rect 1509 21586 1515 21620
rect 1469 21547 1515 21586
rect 1469 21513 1475 21547
rect 1509 21513 1515 21547
rect 1469 21474 1515 21513
rect 1469 21440 1475 21474
rect 1509 21440 1515 21474
tri 1279 21408 1291 21420 sw
tri 1457 21408 1469 21420 se
rect 1469 21408 1515 21440
rect 1705 21912 1751 21924
rect 1705 21878 1711 21912
rect 1745 21878 1751 21912
rect 1705 21839 1751 21878
rect 1705 21805 1711 21839
rect 1745 21805 1751 21839
rect 1705 21766 1751 21805
rect 1705 21732 1711 21766
rect 1745 21732 1751 21766
rect 1705 21693 1751 21732
rect 1705 21659 1711 21693
rect 1745 21659 1751 21693
rect 1705 21620 1751 21659
rect 1705 21586 1711 21620
rect 1745 21586 1751 21620
rect 1705 21547 1751 21586
rect 1705 21513 1711 21547
rect 1745 21513 1751 21547
rect 1705 21474 1751 21513
rect 1705 21440 1711 21474
rect 1745 21440 1751 21474
tri 1515 21408 1527 21420 sw
tri 1693 21408 1705 21420 se
rect 1705 21408 1751 21440
rect 1941 21912 1987 21924
rect 1941 21878 1947 21912
rect 1981 21878 1987 21912
rect 1941 21839 1987 21878
rect 1941 21805 1947 21839
rect 1981 21805 1987 21839
rect 1941 21766 1987 21805
rect 1941 21732 1947 21766
rect 1981 21732 1987 21766
rect 1941 21693 1987 21732
rect 1941 21659 1947 21693
rect 1981 21659 1987 21693
rect 1941 21620 1987 21659
rect 1941 21586 1947 21620
rect 1981 21586 1987 21620
rect 1941 21547 1987 21586
rect 1941 21513 1947 21547
rect 1981 21513 1987 21547
rect 1941 21474 1987 21513
rect 1941 21440 1947 21474
rect 1981 21440 1987 21474
tri 1751 21408 1763 21420 sw
tri 1929 21408 1941 21420 se
rect 1941 21408 1987 21440
rect 2177 21912 2223 21924
rect 2177 21878 2183 21912
rect 2217 21878 2223 21912
rect 2177 21839 2223 21878
rect 2177 21805 2183 21839
rect 2217 21805 2223 21839
rect 2177 21766 2223 21805
rect 2177 21732 2183 21766
rect 2217 21732 2223 21766
rect 2177 21693 2223 21732
rect 2177 21659 2183 21693
rect 2217 21659 2223 21693
rect 2177 21620 2223 21659
rect 2177 21586 2183 21620
rect 2217 21586 2223 21620
rect 2177 21547 2223 21586
rect 2177 21513 2183 21547
rect 2217 21513 2223 21547
rect 2177 21474 2223 21513
rect 2177 21440 2183 21474
rect 2217 21440 2223 21474
tri 1987 21408 1999 21420 sw
tri 2165 21408 2177 21420 se
rect 2177 21408 2223 21440
rect 2413 21912 2459 21924
rect 2413 21878 2419 21912
rect 2453 21878 2459 21912
rect 2413 21839 2459 21878
rect 2413 21805 2419 21839
rect 2453 21805 2459 21839
rect 2413 21766 2459 21805
rect 2413 21732 2419 21766
rect 2453 21732 2459 21766
rect 2413 21693 2459 21732
rect 2413 21659 2419 21693
rect 2453 21659 2459 21693
rect 2413 21620 2459 21659
rect 2413 21586 2419 21620
rect 2453 21586 2459 21620
rect 2413 21547 2459 21586
rect 2413 21513 2419 21547
rect 2453 21513 2459 21547
rect 2413 21474 2459 21513
rect 2413 21440 2419 21474
rect 2453 21440 2459 21474
tri 2223 21408 2235 21420 sw
tri 2401 21408 2413 21420 se
rect 2413 21408 2459 21440
rect 2649 21912 2695 21924
rect 2649 21878 2655 21912
rect 2689 21878 2695 21912
rect 2649 21839 2695 21878
rect 2649 21805 2655 21839
rect 2689 21805 2695 21839
rect 2649 21766 2695 21805
rect 2649 21732 2655 21766
rect 2689 21732 2695 21766
rect 2649 21693 2695 21732
rect 2649 21659 2655 21693
rect 2689 21659 2695 21693
rect 2649 21620 2695 21659
rect 2649 21586 2655 21620
rect 2689 21586 2695 21620
rect 2649 21547 2695 21586
rect 2649 21513 2655 21547
rect 2689 21513 2695 21547
rect 2649 21474 2695 21513
rect 2649 21440 2655 21474
rect 2689 21440 2695 21474
tri 2459 21408 2471 21420 sw
tri 2637 21408 2649 21420 se
rect 2649 21408 2695 21440
rect 2885 21912 3076 21936
rect 2885 21878 2891 21912
rect 2925 21898 3076 21912
rect 2925 21878 3036 21898
rect 2885 21864 3036 21878
rect 3070 21864 3076 21898
rect 2885 21839 3076 21864
rect 2885 21805 2891 21839
rect 2925 21826 3076 21839
rect 2925 21805 3036 21826
rect 2885 21792 3036 21805
rect 3070 21792 3076 21826
rect 2885 21766 3076 21792
rect 2885 21732 2891 21766
rect 2925 21754 3076 21766
rect 2925 21732 3036 21754
rect 2885 21720 3036 21732
rect 3070 21720 3076 21754
rect 2885 21693 3076 21720
rect 2885 21659 2891 21693
rect 2925 21682 3076 21693
rect 2925 21659 3036 21682
rect 2885 21648 3036 21659
rect 3070 21648 3076 21682
rect 2885 21620 3076 21648
rect 2885 21586 2891 21620
rect 2925 21610 3076 21620
rect 2925 21586 3036 21610
rect 2885 21576 3036 21586
rect 3070 21576 3076 21610
rect 2885 21547 3076 21576
rect 2885 21513 2891 21547
rect 2925 21538 3076 21547
rect 2925 21513 3036 21538
rect 2885 21504 3036 21513
rect 3070 21504 3076 21538
rect 2885 21474 3076 21504
rect 2885 21440 2891 21474
rect 2925 21466 3076 21474
rect 2925 21440 3036 21466
rect 2885 21432 3036 21440
rect 3070 21432 3076 21466
tri 2695 21408 2707 21420 sw
tri 2873 21408 2885 21420 se
rect 2885 21408 3076 21432
rect 380 21401 583 21408
tri 583 21401 590 21408 sw
tri 742 21401 749 21408 se
rect 749 21401 819 21408
tri 819 21401 826 21408 sw
tri 978 21401 985 21408 se
rect 985 21401 1055 21408
tri 1055 21401 1062 21408 sw
tri 1214 21401 1221 21408 se
rect 1221 21401 1291 21408
tri 1291 21401 1298 21408 sw
tri 1450 21401 1457 21408 se
rect 1457 21401 1527 21408
tri 1527 21401 1534 21408 sw
tri 1686 21401 1693 21408 se
rect 1693 21401 1763 21408
tri 1763 21401 1770 21408 sw
tri 1922 21401 1929 21408 se
rect 1929 21401 1999 21408
tri 1999 21401 2006 21408 sw
tri 2158 21401 2165 21408 se
rect 2165 21401 2235 21408
tri 2235 21401 2242 21408 sw
tri 2394 21401 2401 21408 se
rect 2401 21401 2471 21408
tri 2471 21401 2478 21408 sw
tri 2630 21401 2637 21408 se
rect 2637 21401 2707 21408
tri 2707 21401 2714 21408 sw
tri 2866 21401 2873 21408 se
rect 2873 21401 3076 21408
rect 380 21375 531 21401
rect 380 21341 386 21375
rect 420 21367 531 21375
rect 565 21386 590 21401
tri 590 21386 605 21401 sw
tri 727 21386 742 21401 se
rect 742 21386 767 21401
rect 565 21367 767 21386
rect 801 21386 826 21401
tri 826 21386 841 21401 sw
tri 963 21386 978 21401 se
rect 978 21386 1003 21401
rect 801 21367 1003 21386
rect 1037 21386 1062 21401
tri 1062 21386 1077 21401 sw
tri 1199 21386 1214 21401 se
rect 1214 21386 1239 21401
rect 1037 21367 1239 21386
rect 1273 21386 1298 21401
tri 1298 21386 1313 21401 sw
tri 1435 21386 1450 21401 se
rect 1450 21386 1475 21401
rect 1273 21367 1475 21386
rect 1509 21386 1534 21401
tri 1534 21386 1549 21401 sw
tri 1671 21386 1686 21401 se
rect 1686 21386 1711 21401
rect 1509 21367 1711 21386
rect 1745 21386 1770 21401
tri 1770 21386 1785 21401 sw
tri 1907 21386 1922 21401 se
rect 1922 21386 1947 21401
rect 1745 21367 1947 21386
rect 1981 21386 2006 21401
tri 2006 21386 2021 21401 sw
tri 2143 21386 2158 21401 se
rect 2158 21386 2183 21401
rect 1981 21367 2183 21386
rect 2217 21386 2242 21401
tri 2242 21386 2257 21401 sw
tri 2379 21386 2394 21401 se
rect 2394 21386 2419 21401
rect 2217 21367 2419 21386
rect 2453 21386 2478 21401
tri 2478 21386 2493 21401 sw
tri 2615 21386 2630 21401 se
rect 2630 21386 2655 21401
rect 2453 21367 2655 21386
rect 2689 21386 2714 21401
tri 2714 21386 2729 21401 sw
tri 2851 21386 2866 21401 se
rect 2866 21386 2891 21401
rect 2689 21367 2891 21386
rect 2925 21394 3076 21401
rect 2925 21367 3036 21394
rect 420 21361 3036 21367
rect 420 21341 697 21361
rect 380 21328 697 21341
rect 380 21303 531 21328
rect 380 21269 386 21303
rect 420 21294 531 21303
rect 565 21309 697 21328
rect 749 21309 765 21361
rect 817 21309 833 21361
rect 885 21309 901 21361
rect 953 21309 969 21361
rect 1021 21328 1037 21361
rect 1089 21309 1105 21361
rect 1157 21309 1173 21361
rect 1225 21328 1241 21361
rect 1293 21328 2097 21361
rect 1225 21309 1239 21328
rect 1293 21309 1475 21328
rect 565 21297 767 21309
rect 801 21297 1003 21309
rect 1037 21297 1239 21309
rect 1273 21297 1475 21309
rect 565 21294 697 21297
rect 420 21269 697 21294
rect 380 21255 697 21269
rect 380 21231 531 21255
rect 380 21197 386 21231
rect 420 21221 531 21231
rect 565 21245 697 21255
rect 749 21245 765 21297
rect 817 21245 833 21297
rect 885 21245 901 21297
rect 953 21245 969 21297
rect 1021 21255 1037 21294
rect 1089 21245 1105 21297
rect 1157 21245 1173 21297
rect 1225 21294 1239 21297
rect 1293 21294 1475 21297
rect 1509 21294 1711 21328
rect 1745 21294 1947 21328
rect 1981 21309 2097 21328
rect 2149 21309 2165 21361
rect 2217 21309 2233 21361
rect 2285 21309 2301 21361
rect 2353 21309 2369 21361
rect 2421 21328 2437 21361
rect 2489 21309 2505 21361
rect 2557 21309 2573 21361
rect 2625 21309 2641 21361
rect 2693 21360 3036 21361
rect 3070 21360 3076 21394
rect 2693 21328 3076 21360
rect 2693 21309 2891 21328
rect 1981 21297 2183 21309
rect 2217 21297 2419 21309
rect 2453 21297 2655 21309
rect 2689 21297 2891 21309
rect 1981 21294 2097 21297
rect 1225 21255 1241 21294
rect 1293 21255 2097 21294
rect 1225 21245 1239 21255
rect 1293 21245 1475 21255
rect 565 21233 767 21245
rect 801 21233 1003 21245
rect 1037 21233 1239 21245
rect 1273 21233 1475 21245
rect 565 21221 697 21233
rect 420 21197 697 21221
rect 380 21182 697 21197
rect 380 21159 531 21182
rect 380 21125 386 21159
rect 420 21148 531 21159
rect 565 21181 697 21182
rect 749 21181 765 21233
rect 817 21181 833 21233
rect 885 21181 901 21233
rect 953 21181 969 21233
rect 1021 21182 1037 21221
rect 1089 21181 1105 21233
rect 1157 21181 1173 21233
rect 1225 21221 1239 21233
rect 1293 21221 1475 21233
rect 1509 21221 1711 21255
rect 1745 21221 1947 21255
rect 1981 21245 2097 21255
rect 2149 21245 2165 21297
rect 2217 21245 2233 21297
rect 2285 21245 2301 21297
rect 2353 21245 2369 21297
rect 2421 21255 2437 21294
rect 2489 21245 2505 21297
rect 2557 21245 2573 21297
rect 2625 21245 2641 21297
rect 2693 21294 2891 21297
rect 2925 21322 3076 21328
rect 2925 21294 3036 21322
rect 2693 21288 3036 21294
rect 3070 21288 3076 21322
rect 2693 21255 3076 21288
rect 2693 21245 2891 21255
rect 1981 21233 2183 21245
rect 2217 21233 2419 21245
rect 2453 21233 2655 21245
rect 2689 21233 2891 21245
rect 1981 21221 2097 21233
rect 1225 21182 1241 21221
rect 1293 21182 2097 21221
rect 1225 21181 1239 21182
rect 1293 21181 1475 21182
rect 565 21169 767 21181
rect 801 21169 1003 21181
rect 1037 21169 1239 21181
rect 1273 21169 1475 21181
rect 565 21148 697 21169
rect 420 21125 697 21148
rect 380 21117 697 21125
rect 749 21117 765 21169
rect 817 21117 833 21169
rect 885 21117 901 21169
rect 953 21117 969 21169
rect 1021 21117 1037 21148
rect 1089 21117 1105 21169
rect 1157 21117 1173 21169
rect 1225 21148 1239 21169
rect 1293 21148 1475 21169
rect 1509 21148 1711 21182
rect 1745 21148 1947 21182
rect 1981 21181 2097 21182
rect 2149 21181 2165 21233
rect 2217 21181 2233 21233
rect 2285 21181 2301 21233
rect 2353 21181 2369 21233
rect 2421 21182 2437 21221
rect 2489 21181 2505 21233
rect 2557 21181 2573 21233
rect 2625 21181 2641 21233
rect 2693 21221 2891 21233
rect 2925 21250 3076 21255
rect 2925 21221 3036 21250
rect 2693 21216 3036 21221
rect 3070 21216 3076 21250
rect 2693 21182 3076 21216
rect 2693 21181 2891 21182
rect 1981 21169 2183 21181
rect 2217 21169 2419 21181
rect 2453 21169 2655 21181
rect 2689 21169 2891 21181
rect 1981 21148 2097 21169
rect 1225 21117 1241 21148
rect 1293 21117 2097 21148
rect 2149 21117 2165 21169
rect 2217 21117 2233 21169
rect 2285 21117 2301 21169
rect 2353 21117 2369 21169
rect 2421 21117 2437 21148
rect 2489 21117 2505 21169
rect 2557 21117 2573 21169
rect 2625 21117 2641 21169
rect 2693 21148 2891 21169
rect 2925 21178 3076 21182
rect 2925 21148 3036 21178
rect 2693 21144 3036 21148
rect 3070 21144 3076 21178
rect 2693 21117 3076 21144
rect 380 21109 3076 21117
rect 380 21087 531 21109
rect 380 21053 386 21087
rect 420 21075 531 21087
rect 565 21105 767 21109
rect 801 21105 1003 21109
rect 1037 21105 1239 21109
rect 1273 21105 1475 21109
rect 565 21075 697 21105
rect 420 21053 697 21075
rect 749 21053 765 21105
rect 817 21053 833 21105
rect 885 21053 901 21105
rect 953 21053 969 21105
rect 1021 21053 1037 21075
rect 1089 21053 1105 21105
rect 1157 21053 1173 21105
rect 1225 21075 1239 21105
rect 1293 21075 1475 21105
rect 1509 21075 1711 21109
rect 1745 21075 1947 21109
rect 1981 21105 2183 21109
rect 2217 21105 2419 21109
rect 2453 21105 2655 21109
rect 2689 21105 2891 21109
rect 1981 21075 2097 21105
rect 1225 21053 1241 21075
rect 1293 21053 2097 21075
rect 2149 21053 2165 21105
rect 2217 21053 2233 21105
rect 2285 21053 2301 21105
rect 2353 21053 2369 21105
rect 2421 21053 2437 21075
rect 2489 21053 2505 21105
rect 2557 21053 2573 21105
rect 2625 21053 2641 21105
rect 2693 21075 2891 21105
rect 2925 21106 3076 21109
rect 2925 21075 3036 21106
rect 2693 21072 3036 21075
rect 3070 21072 3076 21106
rect 2693 21053 3076 21072
rect 380 21041 3076 21053
rect 380 21036 697 21041
rect 380 21015 531 21036
rect 380 20981 386 21015
rect 420 21002 531 21015
rect 565 21002 697 21036
rect 420 20989 697 21002
rect 749 20989 765 21041
rect 817 20989 833 21041
rect 885 20989 901 21041
rect 953 20989 969 21041
rect 1021 21036 1037 21041
rect 1021 20989 1037 21002
rect 1089 20989 1105 21041
rect 1157 20989 1173 21041
rect 1225 21036 1241 21041
rect 1293 21036 2097 21041
rect 1225 21002 1239 21036
rect 1293 21002 1475 21036
rect 1509 21002 1711 21036
rect 1745 21002 1947 21036
rect 1981 21002 2097 21036
rect 1225 20989 1241 21002
rect 1293 20989 2097 21002
rect 2149 20989 2165 21041
rect 2217 20989 2233 21041
rect 2285 20989 2301 21041
rect 2353 20989 2369 21041
rect 2421 21036 2437 21041
rect 2421 20989 2437 21002
rect 2489 20989 2505 21041
rect 2557 20989 2573 21041
rect 2625 20989 2641 21041
rect 2693 21036 3076 21041
rect 2693 21002 2891 21036
rect 2925 21034 3076 21036
rect 2925 21002 3036 21034
rect 2693 21000 3036 21002
rect 3070 21000 3076 21034
rect 2693 20989 3076 21000
rect 420 20981 3076 20989
rect 380 20977 3076 20981
rect 380 20962 697 20977
rect 380 20943 531 20962
rect 380 20909 386 20943
rect 420 20928 531 20943
rect 565 20928 697 20962
rect 420 20925 697 20928
rect 749 20925 765 20977
rect 817 20925 833 20977
rect 885 20925 901 20977
rect 953 20925 969 20977
rect 1021 20962 1037 20977
rect 1021 20925 1037 20928
rect 1089 20925 1105 20977
rect 1157 20925 1173 20977
rect 1225 20962 1241 20977
rect 1293 20962 2097 20977
rect 1225 20928 1239 20962
rect 1293 20928 1475 20962
rect 1509 20928 1711 20962
rect 1745 20928 1947 20962
rect 1981 20928 2097 20962
rect 1225 20925 1241 20928
rect 1293 20925 2097 20928
rect 2149 20925 2165 20977
rect 2217 20925 2233 20977
rect 2285 20925 2301 20977
rect 2353 20925 2369 20977
rect 2421 20962 2437 20977
rect 2421 20925 2437 20928
rect 2489 20925 2505 20977
rect 2557 20925 2573 20977
rect 2625 20925 2641 20977
rect 2693 20962 3076 20977
rect 2693 20928 2891 20962
rect 2925 20928 3036 20962
rect 3070 20928 3076 20962
rect 2693 20925 3076 20928
rect 420 20913 3076 20925
rect 420 20909 697 20913
rect 380 20888 697 20909
rect 380 20871 531 20888
rect 380 20837 386 20871
rect 420 20854 531 20871
rect 565 20861 697 20888
rect 749 20861 765 20913
rect 817 20861 833 20913
rect 885 20861 901 20913
rect 953 20861 969 20913
rect 1021 20888 1037 20913
rect 1089 20861 1105 20913
rect 1157 20861 1173 20913
rect 1225 20888 1241 20913
rect 1293 20888 2097 20913
rect 1225 20861 1239 20888
rect 1293 20861 1475 20888
rect 565 20854 767 20861
rect 801 20854 1003 20861
rect 1037 20854 1239 20861
rect 1273 20854 1475 20861
rect 1509 20854 1711 20888
rect 1745 20854 1947 20888
rect 1981 20861 2097 20888
rect 2149 20861 2165 20913
rect 2217 20861 2233 20913
rect 2285 20861 2301 20913
rect 2353 20861 2369 20913
rect 2421 20888 2437 20913
rect 2489 20861 2505 20913
rect 2557 20861 2573 20913
rect 2625 20861 2641 20913
rect 2693 20890 3076 20913
rect 2693 20888 3036 20890
rect 2693 20861 2891 20888
rect 1981 20854 2183 20861
rect 2217 20854 2419 20861
rect 2453 20854 2655 20861
rect 2689 20854 2891 20861
rect 2925 20856 3036 20888
rect 3070 20856 3076 20890
rect 2925 20854 3076 20856
rect 420 20849 3076 20854
rect 420 20837 697 20849
rect 380 20814 697 20837
rect 380 20799 531 20814
rect 380 20765 386 20799
rect 420 20780 531 20799
rect 565 20797 697 20814
rect 749 20797 765 20849
rect 817 20797 833 20849
rect 885 20797 901 20849
rect 953 20797 969 20849
rect 1021 20814 1037 20849
rect 1089 20797 1105 20849
rect 1157 20797 1173 20849
rect 1225 20814 1241 20849
rect 1293 20814 2097 20849
rect 1225 20797 1239 20814
rect 1293 20797 1475 20814
rect 565 20785 767 20797
rect 801 20785 1003 20797
rect 1037 20785 1239 20797
rect 1273 20785 1475 20797
rect 565 20780 697 20785
rect 420 20765 697 20780
rect 380 20740 697 20765
rect 380 20727 531 20740
rect 380 20693 386 20727
rect 420 20706 531 20727
rect 565 20733 697 20740
rect 749 20733 765 20785
rect 817 20733 833 20785
rect 885 20733 901 20785
rect 953 20733 969 20785
rect 1021 20740 1037 20780
rect 1089 20733 1105 20785
rect 1157 20733 1173 20785
rect 1225 20780 1239 20785
rect 1293 20780 1475 20785
rect 1509 20780 1711 20814
rect 1745 20780 1947 20814
rect 1981 20797 2097 20814
rect 2149 20797 2165 20849
rect 2217 20797 2233 20849
rect 2285 20797 2301 20849
rect 2353 20797 2369 20849
rect 2421 20814 2437 20849
rect 2489 20797 2505 20849
rect 2557 20797 2573 20849
rect 2625 20797 2641 20849
rect 2693 20818 3076 20849
rect 2693 20814 3036 20818
rect 2693 20797 2891 20814
rect 1981 20785 2183 20797
rect 2217 20785 2419 20797
rect 2453 20785 2655 20797
rect 2689 20785 2891 20797
rect 1981 20780 2097 20785
rect 1225 20740 1241 20780
rect 1293 20740 2097 20780
rect 1225 20733 1239 20740
rect 1293 20733 1475 20740
rect 565 20721 767 20733
rect 801 20721 1003 20733
rect 1037 20721 1239 20733
rect 1273 20721 1475 20733
rect 565 20706 697 20721
rect 420 20693 697 20706
rect 380 20669 697 20693
rect 749 20669 765 20721
rect 817 20669 833 20721
rect 885 20669 901 20721
rect 953 20669 969 20721
rect 1021 20669 1037 20706
rect 1089 20669 1105 20721
rect 1157 20669 1173 20721
rect 1225 20706 1239 20721
rect 1293 20706 1475 20721
rect 1509 20706 1711 20740
rect 1745 20706 1947 20740
rect 1981 20733 2097 20740
rect 2149 20733 2165 20785
rect 2217 20733 2233 20785
rect 2285 20733 2301 20785
rect 2353 20733 2369 20785
rect 2421 20740 2437 20780
rect 2489 20733 2505 20785
rect 2557 20733 2573 20785
rect 2625 20733 2641 20785
rect 2693 20780 2891 20785
rect 2925 20784 3036 20814
rect 3070 20784 3076 20818
rect 2925 20780 3076 20784
rect 2693 20746 3076 20780
rect 2693 20740 3036 20746
rect 2693 20733 2891 20740
rect 1981 20721 2183 20733
rect 2217 20721 2419 20733
rect 2453 20721 2655 20733
rect 2689 20721 2891 20733
rect 1981 20706 2097 20721
rect 1225 20669 1241 20706
rect 1293 20669 2097 20706
rect 2149 20669 2165 20721
rect 2217 20669 2233 20721
rect 2285 20669 2301 20721
rect 2353 20669 2369 20721
rect 2421 20669 2437 20706
rect 2489 20669 2505 20721
rect 2557 20669 2573 20721
rect 2625 20669 2641 20721
rect 2693 20706 2891 20721
rect 2925 20712 3036 20740
rect 3070 20712 3076 20746
rect 2925 20706 3076 20712
rect 2693 20674 3076 20706
rect 2693 20669 3036 20674
rect 380 20666 3036 20669
rect 380 20655 531 20666
rect 380 20621 386 20655
rect 420 20632 531 20655
rect 565 20657 767 20666
rect 801 20657 1003 20666
rect 1037 20657 1239 20666
rect 1273 20657 1475 20666
rect 565 20632 697 20657
rect 420 20621 697 20632
rect 380 20605 697 20621
rect 749 20605 765 20657
rect 817 20605 833 20657
rect 885 20605 901 20657
rect 953 20605 969 20657
rect 1021 20605 1037 20632
rect 1089 20605 1105 20657
rect 1157 20605 1173 20657
rect 1225 20632 1239 20657
rect 1293 20632 1475 20657
rect 1509 20632 1711 20666
rect 1745 20632 1947 20666
rect 1981 20657 2183 20666
rect 2217 20657 2419 20666
rect 2453 20657 2655 20666
rect 2689 20657 2891 20666
rect 1981 20632 2097 20657
rect 1225 20605 1241 20632
rect 1293 20605 2097 20632
rect 2149 20605 2165 20657
rect 2217 20605 2233 20657
rect 2285 20605 2301 20657
rect 2353 20605 2369 20657
rect 2421 20605 2437 20632
rect 2489 20605 2505 20657
rect 2557 20605 2573 20657
rect 2625 20605 2641 20657
rect 2693 20632 2891 20657
rect 2925 20640 3036 20666
rect 3070 20640 3076 20674
rect 2925 20632 3076 20640
rect 2693 20605 3076 20632
rect 380 20602 3076 20605
rect 380 20593 3036 20602
rect 380 20592 697 20593
rect 380 20583 531 20592
rect 380 20549 386 20583
rect 420 20558 531 20583
rect 565 20558 697 20592
rect 420 20549 697 20558
rect 380 20541 697 20549
rect 749 20541 765 20593
rect 817 20541 833 20593
rect 885 20541 901 20593
rect 953 20541 969 20593
rect 1021 20592 1037 20593
rect 1021 20541 1037 20558
rect 1089 20541 1105 20593
rect 1157 20541 1173 20593
rect 1225 20592 1241 20593
rect 1293 20592 2097 20593
rect 1225 20558 1239 20592
rect 1293 20558 1475 20592
rect 1509 20558 1711 20592
rect 1745 20558 1947 20592
rect 1981 20558 2097 20592
rect 1225 20541 1241 20558
rect 1293 20541 2097 20558
rect 2149 20541 2165 20593
rect 2217 20541 2233 20593
rect 2285 20541 2301 20593
rect 2353 20541 2369 20593
rect 2421 20592 2437 20593
rect 2421 20541 2437 20558
rect 2489 20541 2505 20593
rect 2557 20541 2573 20593
rect 2625 20541 2641 20593
rect 2693 20592 3036 20593
rect 2693 20558 2891 20592
rect 2925 20568 3036 20592
rect 3070 20568 3076 20602
rect 2925 20558 3076 20568
rect 2693 20541 3076 20558
rect 380 20530 3076 20541
rect 380 20529 3036 20530
rect 380 20518 697 20529
rect 380 20511 531 20518
rect 380 20477 386 20511
rect 420 20484 531 20511
rect 565 20484 697 20518
rect 420 20477 697 20484
rect 749 20477 765 20529
rect 817 20477 833 20529
rect 885 20477 901 20529
rect 953 20477 969 20529
rect 1021 20518 1037 20529
rect 1021 20477 1037 20484
rect 1089 20477 1105 20529
rect 1157 20477 1173 20529
rect 1225 20518 1241 20529
rect 1293 20518 2097 20529
rect 1225 20484 1239 20518
rect 1293 20484 1475 20518
rect 1509 20484 1711 20518
rect 1745 20484 1947 20518
rect 1981 20484 2097 20518
rect 1225 20477 1241 20484
rect 1293 20477 2097 20484
rect 2149 20477 2165 20529
rect 2217 20477 2233 20529
rect 2285 20477 2301 20529
rect 2353 20477 2369 20529
rect 2421 20518 2437 20529
rect 2421 20477 2437 20484
rect 2489 20477 2505 20529
rect 2557 20477 2573 20529
rect 2625 20477 2641 20529
rect 2693 20518 3036 20529
rect 2693 20484 2891 20518
rect 2925 20496 3036 20518
rect 3070 20496 3076 20530
rect 2925 20484 3076 20496
rect 2693 20477 3076 20484
rect 380 20465 3076 20477
rect 380 20444 697 20465
rect 380 20439 531 20444
rect 380 20405 386 20439
rect 420 20410 531 20439
rect 565 20413 697 20444
rect 749 20413 765 20465
rect 817 20413 833 20465
rect 885 20413 901 20465
rect 953 20413 969 20465
rect 1021 20444 1037 20465
rect 1089 20413 1105 20465
rect 1157 20413 1173 20465
rect 1225 20444 1241 20465
rect 1293 20444 2097 20465
rect 1225 20413 1239 20444
rect 1293 20413 1475 20444
rect 565 20410 767 20413
rect 801 20410 1003 20413
rect 1037 20410 1239 20413
rect 1273 20410 1475 20413
rect 1509 20410 1711 20444
rect 1745 20410 1947 20444
rect 1981 20413 2097 20444
rect 2149 20413 2165 20465
rect 2217 20413 2233 20465
rect 2285 20413 2301 20465
rect 2353 20413 2369 20465
rect 2421 20444 2437 20465
rect 2489 20413 2505 20465
rect 2557 20413 2573 20465
rect 2625 20413 2641 20465
rect 2693 20458 3076 20465
rect 2693 20444 3036 20458
rect 2693 20413 2891 20444
rect 1981 20410 2183 20413
rect 2217 20410 2419 20413
rect 2453 20410 2655 20413
rect 2689 20410 2891 20413
rect 2925 20424 3036 20444
rect 3070 20424 3076 20458
rect 2925 20410 3076 20424
rect 420 20405 3076 20410
rect 380 20386 3076 20405
rect 380 20370 589 20386
tri 589 20370 605 20386 nw
tri 727 20370 743 20386 ne
rect 743 20370 825 20386
tri 825 20370 841 20386 nw
tri 963 20370 979 20386 ne
rect 979 20370 1061 20386
tri 1061 20370 1077 20386 nw
tri 1199 20370 1215 20386 ne
rect 1215 20370 1297 20386
tri 1297 20370 1313 20386 nw
tri 1435 20370 1451 20386 ne
rect 1451 20370 1533 20386
tri 1533 20370 1549 20386 nw
tri 1671 20370 1687 20386 ne
rect 1687 20370 1769 20386
tri 1769 20370 1785 20386 nw
tri 1907 20370 1923 20386 ne
rect 1923 20370 2005 20386
tri 2005 20370 2021 20386 nw
tri 2143 20370 2159 20386 ne
rect 2159 20370 2241 20386
tri 2241 20370 2257 20386 nw
tri 2379 20370 2395 20386 ne
rect 2395 20370 2477 20386
tri 2477 20370 2493 20386 nw
tri 2615 20370 2631 20386 ne
rect 2631 20370 2713 20386
tri 2713 20370 2729 20386 nw
tri 2851 20370 2867 20386 ne
rect 2867 20370 3036 20386
rect 380 20367 531 20370
rect 380 20333 386 20367
rect 420 20336 531 20367
rect 565 20336 571 20370
tri 571 20352 589 20370 nw
tri 743 20352 761 20370 ne
rect 420 20333 571 20336
rect 380 20296 571 20333
rect 380 20295 531 20296
rect 380 20261 386 20295
rect 420 20262 531 20295
rect 565 20262 571 20296
rect 420 20261 571 20262
rect 380 20223 571 20261
rect 380 20189 386 20223
rect 420 20222 571 20223
rect 420 20189 531 20222
rect 380 20188 531 20189
rect 565 20188 571 20222
rect 380 20151 571 20188
rect 380 20117 386 20151
rect 420 20148 571 20151
rect 420 20117 531 20148
rect 380 20114 531 20117
rect 565 20114 571 20148
rect 380 20079 571 20114
rect 380 20045 386 20079
rect 420 20074 571 20079
rect 420 20045 531 20074
rect 380 20040 531 20045
rect 565 20040 571 20074
rect 380 20007 571 20040
rect 380 19973 386 20007
rect 420 20000 571 20007
rect 420 19973 531 20000
rect 380 19966 531 19973
rect 565 19966 571 20000
rect 380 19935 571 19966
rect 761 20336 767 20370
rect 801 20336 807 20370
tri 807 20352 825 20370 nw
tri 979 20352 997 20370 ne
rect 761 20296 807 20336
rect 761 20262 767 20296
rect 801 20262 807 20296
rect 761 20222 807 20262
rect 761 20188 767 20222
rect 801 20188 807 20222
rect 761 20148 807 20188
rect 761 20114 767 20148
rect 801 20114 807 20148
rect 761 20074 807 20114
rect 761 20040 767 20074
rect 801 20040 807 20074
rect 761 20000 807 20040
rect 761 19966 767 20000
rect 801 19966 807 20000
rect 761 19954 807 19966
rect 997 20336 1003 20370
rect 1037 20336 1043 20370
tri 1043 20352 1061 20370 nw
tri 1215 20352 1233 20370 ne
rect 997 20296 1043 20336
rect 997 20262 1003 20296
rect 1037 20262 1043 20296
rect 997 20222 1043 20262
rect 997 20188 1003 20222
rect 1037 20188 1043 20222
rect 997 20148 1043 20188
rect 997 20114 1003 20148
rect 1037 20114 1043 20148
rect 997 20074 1043 20114
rect 997 20040 1003 20074
rect 1037 20040 1043 20074
rect 997 20000 1043 20040
rect 997 19966 1003 20000
rect 1037 19966 1043 20000
rect 997 19954 1043 19966
rect 1233 20336 1239 20370
rect 1273 20336 1279 20370
tri 1279 20352 1297 20370 nw
tri 1451 20352 1469 20370 ne
rect 1233 20296 1279 20336
rect 1233 20262 1239 20296
rect 1273 20262 1279 20296
rect 1233 20222 1279 20262
rect 1233 20188 1239 20222
rect 1273 20188 1279 20222
rect 1233 20148 1279 20188
rect 1233 20114 1239 20148
rect 1273 20114 1279 20148
rect 1233 20074 1279 20114
rect 1233 20040 1239 20074
rect 1273 20040 1279 20074
rect 1233 20000 1279 20040
rect 1233 19966 1239 20000
rect 1273 19966 1279 20000
rect 1233 19954 1279 19966
rect 1469 20336 1475 20370
rect 1509 20336 1515 20370
tri 1515 20352 1533 20370 nw
tri 1687 20352 1705 20370 ne
rect 1469 20296 1515 20336
rect 1469 20262 1475 20296
rect 1509 20262 1515 20296
rect 1469 20222 1515 20262
rect 1469 20188 1475 20222
rect 1509 20188 1515 20222
rect 1469 20148 1515 20188
rect 1469 20114 1475 20148
rect 1509 20114 1515 20148
rect 1469 20074 1515 20114
rect 1469 20040 1475 20074
rect 1509 20040 1515 20074
rect 1469 20000 1515 20040
rect 1469 19966 1475 20000
rect 1509 19966 1515 20000
rect 1469 19954 1515 19966
rect 1705 20336 1711 20370
rect 1745 20336 1751 20370
tri 1751 20352 1769 20370 nw
tri 1923 20352 1941 20370 ne
rect 1705 20296 1751 20336
rect 1705 20262 1711 20296
rect 1745 20262 1751 20296
rect 1705 20222 1751 20262
rect 1705 20188 1711 20222
rect 1745 20188 1751 20222
rect 1705 20148 1751 20188
rect 1705 20114 1711 20148
rect 1745 20114 1751 20148
rect 1705 20074 1751 20114
rect 1705 20040 1711 20074
rect 1745 20040 1751 20074
rect 1705 20000 1751 20040
rect 1705 19966 1711 20000
rect 1745 19966 1751 20000
rect 1705 19954 1751 19966
rect 1941 20336 1947 20370
rect 1981 20336 1987 20370
tri 1987 20352 2005 20370 nw
tri 2159 20352 2177 20370 ne
rect 1941 20296 1987 20336
rect 1941 20262 1947 20296
rect 1981 20262 1987 20296
rect 1941 20222 1987 20262
rect 1941 20188 1947 20222
rect 1981 20188 1987 20222
rect 1941 20148 1987 20188
rect 1941 20114 1947 20148
rect 1981 20114 1987 20148
rect 1941 20074 1987 20114
rect 1941 20040 1947 20074
rect 1981 20040 1987 20074
rect 1941 20000 1987 20040
rect 1941 19966 1947 20000
rect 1981 19966 1987 20000
rect 1941 19954 1987 19966
rect 2177 20336 2183 20370
rect 2217 20336 2223 20370
tri 2223 20352 2241 20370 nw
tri 2395 20352 2413 20370 ne
rect 2177 20296 2223 20336
rect 2177 20262 2183 20296
rect 2217 20262 2223 20296
rect 2177 20222 2223 20262
rect 2177 20188 2183 20222
rect 2217 20188 2223 20222
rect 2177 20148 2223 20188
rect 2177 20114 2183 20148
rect 2217 20114 2223 20148
rect 2177 20074 2223 20114
rect 2177 20040 2183 20074
rect 2217 20040 2223 20074
rect 2177 20000 2223 20040
rect 2177 19966 2183 20000
rect 2217 19966 2223 20000
rect 2177 19954 2223 19966
rect 2413 20336 2419 20370
rect 2453 20336 2459 20370
tri 2459 20352 2477 20370 nw
tri 2631 20352 2649 20370 ne
rect 2413 20296 2459 20336
rect 2413 20262 2419 20296
rect 2453 20262 2459 20296
rect 2413 20222 2459 20262
rect 2413 20188 2419 20222
rect 2453 20188 2459 20222
rect 2413 20148 2459 20188
rect 2413 20114 2419 20148
rect 2453 20114 2459 20148
rect 2413 20074 2459 20114
rect 2413 20040 2419 20074
rect 2453 20040 2459 20074
rect 2413 20000 2459 20040
rect 2413 19966 2419 20000
rect 2453 19966 2459 20000
rect 2413 19954 2459 19966
rect 2649 20336 2655 20370
rect 2689 20336 2695 20370
tri 2695 20352 2713 20370 nw
tri 2867 20352 2885 20370 ne
rect 2649 20296 2695 20336
rect 2649 20262 2655 20296
rect 2689 20262 2695 20296
rect 2649 20222 2695 20262
rect 2649 20188 2655 20222
rect 2689 20188 2695 20222
rect 2649 20148 2695 20188
rect 2649 20114 2655 20148
rect 2689 20114 2695 20148
rect 2649 20074 2695 20114
rect 2649 20040 2655 20074
rect 2689 20040 2695 20074
rect 2649 20000 2695 20040
rect 2649 19966 2655 20000
rect 2689 19966 2695 20000
rect 2649 19954 2695 19966
rect 2885 20336 2891 20370
rect 2925 20352 3036 20370
rect 3070 20352 3076 20386
rect 2925 20336 3076 20352
rect 2885 20314 3076 20336
rect 2885 20296 3036 20314
rect 2885 20262 2891 20296
rect 2925 20280 3036 20296
rect 3070 20280 3076 20314
rect 2925 20262 3076 20280
rect 2885 20242 3076 20262
rect 2885 20222 3036 20242
rect 2885 20188 2891 20222
rect 2925 20208 3036 20222
rect 3070 20208 3076 20242
rect 2925 20188 3076 20208
rect 2885 20170 3076 20188
rect 2885 20148 3036 20170
rect 2885 20114 2891 20148
rect 2925 20136 3036 20148
rect 3070 20136 3076 20170
rect 2925 20114 3076 20136
rect 2885 20098 3076 20114
rect 2885 20074 3036 20098
rect 2885 20040 2891 20074
rect 2925 20064 3036 20074
rect 3070 20064 3076 20098
rect 2925 20040 3076 20064
rect 2885 20026 3076 20040
rect 2885 20000 3036 20026
rect 2885 19966 2891 20000
rect 2925 19992 3036 20000
rect 3070 19992 3076 20026
rect 2925 19966 3076 19992
rect 2885 19954 3076 19966
rect 380 19901 386 19935
rect 420 19901 571 19935
rect 380 19863 571 19901
rect 2885 19920 3036 19954
rect 3070 19920 3076 19954
rect 380 19829 386 19863
rect 420 19829 571 19863
rect 613 19884 1501 19893
rect 1553 19884 1569 19893
rect 1621 19884 1636 19893
rect 1688 19884 1703 19893
rect 1755 19884 1770 19893
rect 1822 19884 1837 19893
rect 1889 19884 2830 19893
rect 613 19850 625 19884
rect 659 19850 700 19884
rect 734 19850 775 19884
rect 809 19850 850 19884
rect 884 19850 925 19884
rect 959 19850 1000 19884
rect 1034 19850 1075 19884
rect 1109 19850 1150 19884
rect 1184 19850 1225 19884
rect 1259 19850 1300 19884
rect 1334 19850 1375 19884
rect 1409 19850 1450 19884
rect 1484 19850 1501 19884
rect 1559 19850 1569 19884
rect 1634 19850 1636 19884
rect 1889 19850 1896 19884
rect 1930 19850 1970 19884
rect 2004 19850 2044 19884
rect 2078 19850 2118 19884
rect 2152 19850 2192 19884
rect 2226 19850 2266 19884
rect 2300 19850 2340 19884
rect 2374 19850 2414 19884
rect 2448 19850 2488 19884
rect 2522 19850 2562 19884
rect 2596 19850 2636 19884
rect 2670 19850 2710 19884
rect 2744 19850 2784 19884
rect 2818 19850 2830 19884
rect 613 19841 1501 19850
rect 1553 19841 1569 19850
rect 1621 19841 1636 19850
rect 1688 19841 1703 19850
rect 1755 19841 1770 19850
rect 1822 19841 1837 19850
rect 1889 19841 2830 19850
rect 2885 19882 3076 19920
rect 2885 19848 3036 19882
rect 3070 19848 3076 19882
rect 380 19791 571 19829
rect 380 19757 386 19791
rect 420 19768 571 19791
rect 2885 19810 3076 19848
rect 420 19757 531 19768
rect 380 19734 531 19757
rect 565 19734 571 19768
rect 380 19719 571 19734
rect 380 19685 386 19719
rect 420 19695 571 19719
rect 420 19685 531 19695
rect 380 19661 531 19685
rect 565 19661 571 19695
rect 380 19647 571 19661
rect 380 19613 386 19647
rect 420 19622 571 19647
rect 420 19613 531 19622
rect 380 19588 531 19613
rect 565 19588 571 19622
rect 380 19575 571 19588
rect 380 19541 386 19575
rect 420 19549 571 19575
rect 420 19541 531 19549
rect 380 19515 531 19541
rect 565 19515 571 19549
rect 380 19503 571 19515
rect 380 19469 386 19503
rect 420 19476 571 19503
rect 420 19469 531 19476
rect 380 19442 531 19469
rect 565 19442 571 19476
rect 380 19431 571 19442
rect 380 19397 386 19431
rect 420 19403 571 19431
rect 420 19397 531 19403
rect 380 19369 531 19397
rect 565 19369 571 19403
rect 380 19359 571 19369
rect 380 19325 386 19359
rect 420 19330 571 19359
rect 420 19325 531 19330
rect 380 19296 531 19325
rect 565 19296 571 19330
rect 761 19768 807 19780
rect 761 19734 767 19768
rect 801 19734 807 19768
rect 761 19695 807 19734
rect 761 19661 767 19695
rect 801 19661 807 19695
rect 761 19622 807 19661
rect 761 19588 767 19622
rect 801 19588 807 19622
rect 761 19549 807 19588
rect 761 19515 767 19549
rect 801 19515 807 19549
rect 761 19476 807 19515
rect 761 19442 767 19476
rect 801 19442 807 19476
rect 761 19403 807 19442
rect 761 19369 767 19403
rect 801 19369 807 19403
rect 761 19330 807 19369
tri 571 19296 593 19318 sw
tri 739 19296 761 19318 se
rect 761 19296 767 19330
rect 801 19296 807 19330
rect 997 19768 1043 19780
rect 997 19734 1003 19768
rect 1037 19734 1043 19768
rect 997 19695 1043 19734
rect 997 19661 1003 19695
rect 1037 19661 1043 19695
rect 997 19622 1043 19661
rect 997 19588 1003 19622
rect 1037 19588 1043 19622
rect 997 19549 1043 19588
rect 997 19515 1003 19549
rect 1037 19515 1043 19549
rect 997 19476 1043 19515
rect 997 19442 1003 19476
rect 1037 19442 1043 19476
rect 997 19403 1043 19442
rect 997 19369 1003 19403
rect 1037 19369 1043 19403
rect 997 19330 1043 19369
tri 807 19296 829 19318 sw
tri 975 19296 997 19318 se
rect 997 19296 1003 19330
rect 1037 19296 1043 19330
rect 1233 19768 1279 19780
rect 1233 19734 1239 19768
rect 1273 19734 1279 19768
rect 1233 19695 1279 19734
rect 1233 19661 1239 19695
rect 1273 19661 1279 19695
rect 1233 19622 1279 19661
rect 1233 19588 1239 19622
rect 1273 19588 1279 19622
rect 1233 19549 1279 19588
rect 1233 19515 1239 19549
rect 1273 19515 1279 19549
rect 1233 19476 1279 19515
rect 1233 19442 1239 19476
rect 1273 19442 1279 19476
rect 1233 19403 1279 19442
rect 1233 19369 1239 19403
rect 1273 19369 1279 19403
rect 1233 19330 1279 19369
tri 1043 19296 1065 19318 sw
tri 1211 19296 1233 19318 se
rect 1233 19296 1239 19330
rect 1273 19296 1279 19330
rect 1469 19768 1515 19780
rect 1469 19734 1475 19768
rect 1509 19734 1515 19768
rect 1469 19695 1515 19734
rect 1469 19661 1475 19695
rect 1509 19661 1515 19695
rect 1469 19622 1515 19661
rect 1469 19588 1475 19622
rect 1509 19588 1515 19622
rect 1469 19549 1515 19588
rect 1469 19515 1475 19549
rect 1509 19515 1515 19549
rect 1469 19476 1515 19515
rect 1469 19442 1475 19476
rect 1509 19442 1515 19476
rect 1469 19403 1515 19442
rect 1469 19369 1475 19403
rect 1509 19369 1515 19403
rect 1469 19330 1515 19369
tri 1279 19296 1301 19318 sw
tri 1447 19296 1469 19318 se
rect 1469 19296 1475 19330
rect 1509 19296 1515 19330
rect 1705 19768 1751 19780
rect 1705 19734 1711 19768
rect 1745 19734 1751 19768
rect 1705 19695 1751 19734
rect 1705 19661 1711 19695
rect 1745 19661 1751 19695
rect 1705 19622 1751 19661
rect 1705 19588 1711 19622
rect 1745 19588 1751 19622
rect 1705 19549 1751 19588
rect 1705 19515 1711 19549
rect 1745 19515 1751 19549
rect 1705 19476 1751 19515
rect 1705 19442 1711 19476
rect 1745 19442 1751 19476
rect 1705 19403 1751 19442
rect 1705 19369 1711 19403
rect 1745 19369 1751 19403
rect 1705 19330 1751 19369
tri 1515 19296 1537 19318 sw
tri 1683 19296 1705 19318 se
rect 1705 19296 1711 19330
rect 1745 19296 1751 19330
rect 1941 19768 1987 19780
rect 1941 19734 1947 19768
rect 1981 19734 1987 19768
rect 1941 19695 1987 19734
rect 1941 19661 1947 19695
rect 1981 19661 1987 19695
rect 1941 19622 1987 19661
rect 1941 19588 1947 19622
rect 1981 19588 1987 19622
rect 1941 19549 1987 19588
rect 1941 19515 1947 19549
rect 1981 19515 1987 19549
rect 1941 19476 1987 19515
rect 1941 19442 1947 19476
rect 1981 19442 1987 19476
rect 1941 19403 1987 19442
rect 1941 19369 1947 19403
rect 1981 19369 1987 19403
rect 1941 19330 1987 19369
tri 1751 19296 1773 19318 sw
tri 1919 19296 1941 19318 se
rect 1941 19296 1947 19330
rect 1981 19296 1987 19330
rect 2177 19768 2223 19780
rect 2177 19734 2183 19768
rect 2217 19734 2223 19768
rect 2177 19695 2223 19734
rect 2177 19661 2183 19695
rect 2217 19661 2223 19695
rect 2177 19622 2223 19661
rect 2177 19588 2183 19622
rect 2217 19588 2223 19622
rect 2177 19549 2223 19588
rect 2177 19515 2183 19549
rect 2217 19515 2223 19549
rect 2177 19476 2223 19515
rect 2177 19442 2183 19476
rect 2217 19442 2223 19476
rect 2177 19403 2223 19442
rect 2177 19369 2183 19403
rect 2217 19369 2223 19403
rect 2177 19330 2223 19369
tri 1987 19296 2009 19318 sw
tri 2155 19296 2177 19318 se
rect 2177 19296 2183 19330
rect 2217 19296 2223 19330
rect 2413 19768 2459 19780
rect 2413 19734 2419 19768
rect 2453 19734 2459 19768
rect 2413 19695 2459 19734
rect 2413 19661 2419 19695
rect 2453 19661 2459 19695
rect 2413 19622 2459 19661
rect 2413 19588 2419 19622
rect 2453 19588 2459 19622
rect 2413 19549 2459 19588
rect 2413 19515 2419 19549
rect 2453 19515 2459 19549
rect 2413 19476 2459 19515
rect 2413 19442 2419 19476
rect 2453 19442 2459 19476
rect 2413 19403 2459 19442
rect 2413 19369 2419 19403
rect 2453 19369 2459 19403
rect 2413 19330 2459 19369
tri 2223 19296 2245 19318 sw
tri 2391 19296 2413 19318 se
rect 2413 19296 2419 19330
rect 2453 19296 2459 19330
rect 2649 19768 2695 19780
rect 2649 19734 2655 19768
rect 2689 19734 2695 19768
rect 2649 19695 2695 19734
rect 2649 19661 2655 19695
rect 2689 19661 2695 19695
rect 2649 19622 2695 19661
rect 2649 19588 2655 19622
rect 2689 19588 2695 19622
rect 2649 19549 2695 19588
rect 2649 19515 2655 19549
rect 2689 19515 2695 19549
rect 2649 19476 2695 19515
rect 2649 19442 2655 19476
rect 2689 19442 2695 19476
rect 2649 19403 2695 19442
rect 2649 19369 2655 19403
rect 2689 19369 2695 19403
rect 2649 19330 2695 19369
tri 2459 19296 2481 19318 sw
tri 2627 19296 2649 19318 se
rect 2649 19296 2655 19330
rect 2689 19296 2695 19330
rect 2885 19776 3036 19810
rect 3070 19776 3076 19810
rect 2885 19768 3076 19776
rect 2885 19734 2891 19768
rect 2925 19738 3076 19768
rect 2925 19734 3036 19738
rect 2885 19704 3036 19734
rect 3070 19704 3076 19738
rect 2885 19695 3076 19704
rect 2885 19661 2891 19695
rect 2925 19666 3076 19695
rect 2925 19661 3036 19666
rect 2885 19632 3036 19661
rect 3070 19632 3076 19666
rect 2885 19622 3076 19632
rect 2885 19588 2891 19622
rect 2925 19594 3076 19622
rect 2925 19588 3036 19594
rect 2885 19560 3036 19588
rect 3070 19560 3076 19594
rect 2885 19549 3076 19560
rect 2885 19515 2891 19549
rect 2925 19522 3076 19549
rect 2925 19515 3036 19522
rect 2885 19488 3036 19515
rect 3070 19488 3076 19522
rect 2885 19476 3076 19488
rect 2885 19442 2891 19476
rect 2925 19450 3076 19476
rect 2925 19442 3036 19450
rect 2885 19416 3036 19442
rect 3070 19416 3076 19450
rect 2885 19403 3076 19416
rect 2885 19369 2891 19403
rect 2925 19378 3076 19403
rect 2925 19369 3036 19378
rect 2885 19344 3036 19369
rect 3070 19344 3076 19378
rect 2885 19330 3076 19344
tri 2695 19296 2717 19318 sw
tri 2863 19296 2885 19318 se
rect 2885 19296 2891 19330
rect 2925 19306 3076 19330
rect 2925 19296 3036 19306
rect 380 19287 593 19296
rect 380 19253 386 19287
rect 420 19284 593 19287
tri 593 19284 605 19296 sw
tri 727 19284 739 19296 se
rect 739 19284 829 19296
tri 829 19284 841 19296 sw
tri 963 19284 975 19296 se
rect 975 19284 1065 19296
tri 1065 19284 1077 19296 sw
tri 1199 19284 1211 19296 se
rect 1211 19284 1301 19296
tri 1301 19284 1313 19296 sw
tri 1435 19284 1447 19296 se
rect 1447 19284 1537 19296
tri 1537 19284 1549 19296 sw
tri 1671 19284 1683 19296 se
rect 1683 19284 1773 19296
tri 1773 19284 1785 19296 sw
tri 1907 19284 1919 19296 se
rect 1919 19284 2009 19296
tri 2009 19284 2021 19296 sw
tri 2143 19284 2155 19296 se
rect 2155 19284 2245 19296
tri 2245 19284 2257 19296 sw
tri 2379 19284 2391 19296 se
rect 2391 19284 2481 19296
tri 2481 19284 2493 19296 sw
tri 2615 19284 2627 19296 se
rect 2627 19284 2717 19296
tri 2717 19284 2729 19296 sw
tri 2851 19284 2863 19296 se
rect 2863 19284 3036 19296
rect 420 19272 3036 19284
rect 3070 19272 3076 19306
rect 420 19257 3076 19272
rect 420 19253 531 19257
rect 380 19223 531 19253
rect 565 19223 697 19257
rect 380 19215 697 19223
rect 380 19181 386 19215
rect 420 19205 697 19215
rect 749 19205 765 19257
rect 817 19205 833 19257
rect 885 19205 901 19257
rect 953 19205 969 19257
rect 1021 19205 1037 19223
rect 1089 19205 1105 19257
rect 1157 19205 1173 19257
rect 1225 19223 1239 19257
rect 1293 19223 1475 19257
rect 1509 19223 1711 19257
rect 1745 19223 1947 19257
rect 1981 19223 2097 19257
rect 1225 19205 1241 19223
rect 1293 19205 2097 19223
rect 2149 19205 2165 19257
rect 2217 19205 2233 19257
rect 2285 19205 2301 19257
rect 2353 19205 2369 19257
rect 2421 19205 2437 19223
rect 2489 19205 2505 19257
rect 2557 19205 2573 19257
rect 2625 19205 2641 19257
rect 2693 19223 2891 19257
rect 2925 19234 3076 19257
rect 2925 19223 3036 19234
rect 2693 19205 3036 19223
rect 420 19200 3036 19205
rect 3070 19200 3076 19234
rect 420 19193 3076 19200
rect 420 19184 697 19193
rect 420 19181 531 19184
rect 380 19150 531 19181
rect 565 19150 697 19184
rect 380 19143 697 19150
rect 380 19109 386 19143
rect 420 19141 697 19143
rect 749 19141 765 19193
rect 817 19141 833 19193
rect 885 19141 901 19193
rect 953 19141 969 19193
rect 1021 19184 1037 19193
rect 1021 19141 1037 19150
rect 1089 19141 1105 19193
rect 1157 19141 1173 19193
rect 1225 19184 1241 19193
rect 1293 19184 2097 19193
rect 1225 19150 1239 19184
rect 1293 19150 1475 19184
rect 1509 19150 1711 19184
rect 1745 19150 1947 19184
rect 1981 19150 2097 19184
rect 1225 19141 1241 19150
rect 1293 19141 2097 19150
rect 2149 19141 2165 19193
rect 2217 19141 2233 19193
rect 2285 19141 2301 19193
rect 2353 19141 2369 19193
rect 2421 19184 2437 19193
rect 2421 19141 2437 19150
rect 2489 19141 2505 19193
rect 2557 19141 2573 19193
rect 2625 19141 2641 19193
rect 2693 19184 3076 19193
rect 2693 19150 2891 19184
rect 2925 19162 3076 19184
rect 2925 19150 3036 19162
rect 2693 19141 3036 19150
rect 420 19129 3036 19141
rect 420 19111 697 19129
rect 420 19109 531 19111
rect 380 19077 531 19109
rect 565 19077 697 19111
rect 749 19077 765 19129
rect 817 19077 833 19129
rect 885 19077 901 19129
rect 953 19077 969 19129
rect 1021 19111 1037 19129
rect 1089 19077 1105 19129
rect 1157 19077 1173 19129
rect 1225 19111 1241 19129
rect 1293 19111 2097 19129
rect 1225 19077 1239 19111
rect 1293 19077 1475 19111
rect 1509 19077 1711 19111
rect 1745 19077 1947 19111
rect 1981 19077 2097 19111
rect 2149 19077 2165 19129
rect 2217 19077 2233 19129
rect 2285 19077 2301 19129
rect 2353 19077 2369 19129
rect 2421 19111 2437 19129
rect 2489 19077 2505 19129
rect 2557 19077 2573 19129
rect 2625 19077 2641 19129
rect 2693 19128 3036 19129
rect 3070 19128 3076 19162
rect 2693 19111 3076 19128
rect 2693 19077 2891 19111
rect 2925 19090 3076 19111
rect 2925 19077 3036 19090
rect 380 19071 3036 19077
rect 380 19037 386 19071
rect 420 19065 3036 19071
rect 420 19038 697 19065
rect 420 19037 531 19038
rect 380 19004 531 19037
rect 565 19013 697 19038
rect 749 19013 765 19065
rect 817 19013 833 19065
rect 885 19013 901 19065
rect 953 19013 969 19065
rect 1021 19038 1037 19065
rect 1089 19013 1105 19065
rect 1157 19013 1173 19065
rect 1225 19038 1241 19065
rect 1293 19038 2097 19065
rect 1225 19013 1239 19038
rect 1293 19013 1475 19038
rect 565 19004 767 19013
rect 801 19004 1003 19013
rect 1037 19004 1239 19013
rect 1273 19004 1475 19013
rect 1509 19004 1711 19038
rect 1745 19004 1947 19038
rect 1981 19013 2097 19038
rect 2149 19013 2165 19065
rect 2217 19013 2233 19065
rect 2285 19013 2301 19065
rect 2353 19013 2369 19065
rect 2421 19038 2437 19065
rect 2489 19013 2505 19065
rect 2557 19013 2573 19065
rect 2625 19013 2641 19065
rect 2693 19056 3036 19065
rect 3070 19056 3076 19090
rect 2693 19038 3076 19056
rect 2693 19013 2891 19038
rect 1981 19004 2183 19013
rect 2217 19004 2419 19013
rect 2453 19004 2655 19013
rect 2689 19004 2891 19013
rect 2925 19018 3076 19038
rect 2925 19004 3036 19018
rect 380 19001 3036 19004
rect 380 18999 697 19001
rect 380 18965 386 18999
rect 420 18965 697 18999
rect 380 18931 531 18965
rect 565 18949 697 18965
rect 749 18949 765 19001
rect 817 18949 833 19001
rect 885 18949 901 19001
rect 953 18949 969 19001
rect 1021 18965 1037 19001
rect 1089 18949 1105 19001
rect 1157 18949 1173 19001
rect 1225 18965 1241 19001
rect 1293 18965 2097 19001
rect 1225 18949 1239 18965
rect 1293 18949 1475 18965
rect 565 18937 767 18949
rect 801 18937 1003 18949
rect 1037 18937 1239 18949
rect 1273 18937 1475 18949
rect 565 18931 697 18937
rect 380 18927 697 18931
rect 380 18893 386 18927
rect 420 18893 697 18927
rect 380 18892 697 18893
rect 380 18858 531 18892
rect 565 18885 697 18892
rect 749 18885 765 18937
rect 817 18885 833 18937
rect 885 18885 901 18937
rect 953 18885 969 18937
rect 1021 18892 1037 18931
rect 1089 18885 1105 18937
rect 1157 18885 1173 18937
rect 1225 18931 1239 18937
rect 1293 18931 1475 18937
rect 1509 18931 1711 18965
rect 1745 18931 1947 18965
rect 1981 18949 2097 18965
rect 2149 18949 2165 19001
rect 2217 18949 2233 19001
rect 2285 18949 2301 19001
rect 2353 18949 2369 19001
rect 2421 18965 2437 19001
rect 2489 18949 2505 19001
rect 2557 18949 2573 19001
rect 2625 18949 2641 19001
rect 2693 18984 3036 19001
rect 3070 18984 3076 19018
rect 2693 18965 3076 18984
rect 2693 18949 2891 18965
rect 1981 18937 2183 18949
rect 2217 18937 2419 18949
rect 2453 18937 2655 18949
rect 2689 18937 2891 18949
rect 1981 18931 2097 18937
rect 1225 18892 1241 18931
rect 1293 18892 2097 18931
rect 1225 18885 1239 18892
rect 1293 18885 1475 18892
rect 565 18873 767 18885
rect 801 18873 1003 18885
rect 1037 18873 1239 18885
rect 1273 18873 1475 18885
rect 565 18858 697 18873
rect 380 18855 697 18858
rect 380 18821 386 18855
rect 420 18821 697 18855
rect 749 18821 765 18873
rect 817 18821 833 18873
rect 885 18821 901 18873
rect 953 18821 969 18873
rect 1021 18821 1037 18858
rect 1089 18821 1105 18873
rect 1157 18821 1173 18873
rect 1225 18858 1239 18873
rect 1293 18858 1475 18873
rect 1509 18858 1711 18892
rect 1745 18858 1947 18892
rect 1981 18885 2097 18892
rect 2149 18885 2165 18937
rect 2217 18885 2233 18937
rect 2285 18885 2301 18937
rect 2353 18885 2369 18937
rect 2421 18892 2437 18931
rect 2489 18885 2505 18937
rect 2557 18885 2573 18937
rect 2625 18885 2641 18937
rect 2693 18931 2891 18937
rect 2925 18946 3076 18965
rect 2925 18931 3036 18946
rect 2693 18912 3036 18931
rect 3070 18912 3076 18946
rect 2693 18892 3076 18912
rect 2693 18885 2891 18892
rect 1981 18873 2183 18885
rect 2217 18873 2419 18885
rect 2453 18873 2655 18885
rect 2689 18873 2891 18885
rect 1981 18858 2097 18873
rect 1225 18821 1241 18858
rect 1293 18821 2097 18858
rect 2149 18821 2165 18873
rect 2217 18821 2233 18873
rect 2285 18821 2301 18873
rect 2353 18821 2369 18873
rect 2421 18821 2437 18858
rect 2489 18821 2505 18873
rect 2557 18821 2573 18873
rect 2625 18821 2641 18873
rect 2693 18858 2891 18873
rect 2925 18874 3076 18892
rect 2925 18858 3036 18874
rect 2693 18840 3036 18858
rect 3070 18840 3076 18874
rect 2693 18821 3076 18840
rect 380 18818 3076 18821
rect 380 18784 531 18818
rect 565 18809 767 18818
rect 801 18809 1003 18818
rect 1037 18809 1239 18818
rect 1273 18809 1475 18818
rect 565 18784 697 18809
rect 380 18783 697 18784
rect 380 18749 386 18783
rect 420 18757 697 18783
rect 749 18757 765 18809
rect 817 18757 833 18809
rect 885 18757 901 18809
rect 953 18757 969 18809
rect 1021 18757 1037 18784
rect 1089 18757 1105 18809
rect 1157 18757 1173 18809
rect 1225 18784 1239 18809
rect 1293 18784 1475 18809
rect 1509 18784 1711 18818
rect 1745 18784 1947 18818
rect 1981 18809 2183 18818
rect 2217 18809 2419 18818
rect 2453 18809 2655 18818
rect 2689 18809 2891 18818
rect 1981 18784 2097 18809
rect 1225 18757 1241 18784
rect 1293 18757 2097 18784
rect 2149 18757 2165 18809
rect 2217 18757 2233 18809
rect 2285 18757 2301 18809
rect 2353 18757 2369 18809
rect 2421 18757 2437 18784
rect 2489 18757 2505 18809
rect 2557 18757 2573 18809
rect 2625 18757 2641 18809
rect 2693 18784 2891 18809
rect 2925 18802 3076 18818
rect 2925 18784 3036 18802
rect 2693 18768 3036 18784
rect 3070 18768 3076 18802
rect 2693 18757 3076 18768
rect 420 18749 3076 18757
rect 380 18745 3076 18749
rect 380 18744 697 18745
rect 380 18711 531 18744
rect 380 18677 386 18711
rect 420 18710 531 18711
rect 565 18710 697 18744
rect 420 18693 697 18710
rect 749 18693 765 18745
rect 817 18693 833 18745
rect 885 18693 901 18745
rect 953 18693 969 18745
rect 1021 18744 1037 18745
rect 1021 18693 1037 18710
rect 1089 18693 1105 18745
rect 1157 18693 1173 18745
rect 1225 18744 1241 18745
rect 1293 18744 2097 18745
rect 1225 18710 1239 18744
rect 1293 18710 1475 18744
rect 1509 18710 1711 18744
rect 1745 18710 1947 18744
rect 1981 18710 2097 18744
rect 1225 18693 1241 18710
rect 1293 18693 2097 18710
rect 2149 18693 2165 18745
rect 2217 18693 2233 18745
rect 2285 18693 2301 18745
rect 2353 18693 2369 18745
rect 2421 18744 2437 18745
rect 2421 18693 2437 18710
rect 2489 18693 2505 18745
rect 2557 18693 2573 18745
rect 2625 18693 2641 18745
rect 2693 18744 3076 18745
rect 2693 18710 2891 18744
rect 2925 18730 3076 18744
rect 2925 18710 3036 18730
rect 2693 18696 3036 18710
rect 3070 18696 3076 18730
rect 2693 18693 3076 18696
rect 420 18681 3076 18693
rect 420 18677 697 18681
rect 380 18670 697 18677
rect 380 18639 531 18670
rect 380 18605 386 18639
rect 420 18636 531 18639
rect 565 18636 697 18670
rect 420 18629 697 18636
rect 749 18629 765 18681
rect 817 18629 833 18681
rect 885 18629 901 18681
rect 953 18629 969 18681
rect 1021 18670 1037 18681
rect 1021 18629 1037 18636
rect 1089 18629 1105 18681
rect 1157 18629 1173 18681
rect 1225 18670 1241 18681
rect 1293 18670 2097 18681
rect 1225 18636 1239 18670
rect 1293 18636 1475 18670
rect 1509 18636 1711 18670
rect 1745 18636 1947 18670
rect 1981 18636 2097 18670
rect 1225 18629 1241 18636
rect 1293 18629 2097 18636
rect 2149 18629 2165 18681
rect 2217 18629 2233 18681
rect 2285 18629 2301 18681
rect 2353 18629 2369 18681
rect 2421 18670 2437 18681
rect 2421 18629 2437 18636
rect 2489 18629 2505 18681
rect 2557 18629 2573 18681
rect 2625 18629 2641 18681
rect 2693 18670 3076 18681
rect 2693 18636 2891 18670
rect 2925 18658 3076 18670
rect 2925 18636 3036 18658
rect 2693 18629 3036 18636
rect 420 18624 3036 18629
rect 3070 18624 3076 18658
rect 420 18617 3076 18624
rect 420 18605 697 18617
rect 380 18596 697 18605
rect 380 18567 531 18596
rect 380 18533 386 18567
rect 420 18562 531 18567
rect 565 18565 697 18596
rect 749 18565 765 18617
rect 817 18565 833 18617
rect 885 18565 901 18617
rect 953 18565 969 18617
rect 1021 18596 1037 18617
rect 1089 18565 1105 18617
rect 1157 18565 1173 18617
rect 1225 18596 1241 18617
rect 1293 18596 2097 18617
rect 1225 18565 1239 18596
rect 1293 18565 1475 18596
rect 565 18562 767 18565
rect 801 18562 1003 18565
rect 1037 18562 1239 18565
rect 1273 18562 1475 18565
rect 1509 18562 1711 18596
rect 1745 18562 1947 18596
rect 1981 18565 2097 18596
rect 2149 18565 2165 18617
rect 2217 18565 2233 18617
rect 2285 18565 2301 18617
rect 2353 18565 2369 18617
rect 2421 18596 2437 18617
rect 2489 18565 2505 18617
rect 2557 18565 2573 18617
rect 2625 18565 2641 18617
rect 2693 18596 3076 18617
rect 2693 18565 2891 18596
rect 1981 18562 2183 18565
rect 2217 18562 2419 18565
rect 2453 18562 2655 18565
rect 2689 18562 2891 18565
rect 2925 18586 3076 18596
rect 2925 18562 3036 18586
rect 420 18553 3036 18562
rect 420 18533 697 18553
rect 380 18522 697 18533
rect 380 18495 531 18522
rect 380 18461 386 18495
rect 420 18488 531 18495
rect 565 18501 697 18522
rect 749 18501 765 18553
rect 817 18501 833 18553
rect 885 18501 901 18553
rect 953 18501 969 18553
rect 1021 18522 1037 18553
rect 1089 18501 1105 18553
rect 1157 18501 1173 18553
rect 1225 18522 1241 18553
rect 1293 18522 2097 18553
rect 1225 18501 1239 18522
rect 1293 18501 1475 18522
rect 565 18489 767 18501
rect 801 18489 1003 18501
rect 1037 18489 1239 18501
rect 1273 18489 1475 18501
rect 565 18488 697 18489
rect 420 18461 697 18488
rect 380 18448 697 18461
rect 380 18423 531 18448
rect 380 18389 386 18423
rect 420 18414 531 18423
rect 565 18437 697 18448
rect 749 18437 765 18489
rect 817 18437 833 18489
rect 885 18437 901 18489
rect 953 18437 969 18489
rect 1021 18448 1037 18488
rect 1089 18437 1105 18489
rect 1157 18437 1173 18489
rect 1225 18488 1239 18489
rect 1293 18488 1475 18489
rect 1509 18488 1711 18522
rect 1745 18488 1947 18522
rect 1981 18501 2097 18522
rect 2149 18501 2165 18553
rect 2217 18501 2233 18553
rect 2285 18501 2301 18553
rect 2353 18501 2369 18553
rect 2421 18522 2437 18553
rect 2489 18501 2505 18553
rect 2557 18501 2573 18553
rect 2625 18501 2641 18553
rect 2693 18552 3036 18553
rect 3070 18552 3076 18586
rect 2693 18522 3076 18552
rect 2693 18501 2891 18522
rect 1981 18489 2183 18501
rect 2217 18489 2419 18501
rect 2453 18489 2655 18501
rect 2689 18489 2891 18501
rect 1981 18488 2097 18489
rect 1225 18448 1241 18488
rect 1293 18448 2097 18488
rect 1225 18437 1239 18448
rect 1293 18437 1475 18448
rect 565 18425 767 18437
rect 801 18425 1003 18437
rect 1037 18425 1239 18437
rect 1273 18425 1475 18437
rect 565 18414 697 18425
rect 420 18389 697 18414
rect 380 18374 697 18389
rect 380 18351 531 18374
rect 380 18317 386 18351
rect 420 18340 531 18351
rect 565 18373 697 18374
rect 749 18373 765 18425
rect 817 18373 833 18425
rect 885 18373 901 18425
rect 953 18373 969 18425
rect 1021 18374 1037 18414
rect 1089 18373 1105 18425
rect 1157 18373 1173 18425
rect 1225 18414 1239 18425
rect 1293 18414 1475 18425
rect 1509 18414 1711 18448
rect 1745 18414 1947 18448
rect 1981 18437 2097 18448
rect 2149 18437 2165 18489
rect 2217 18437 2233 18489
rect 2285 18437 2301 18489
rect 2353 18437 2369 18489
rect 2421 18448 2437 18488
rect 2489 18437 2505 18489
rect 2557 18437 2573 18489
rect 2625 18437 2641 18489
rect 2693 18488 2891 18489
rect 2925 18514 3076 18522
rect 2925 18488 3036 18514
rect 2693 18480 3036 18488
rect 3070 18480 3076 18514
rect 2693 18448 3076 18480
rect 2693 18437 2891 18448
rect 1981 18425 2183 18437
rect 2217 18425 2419 18437
rect 2453 18425 2655 18437
rect 2689 18425 2891 18437
rect 1981 18414 2097 18425
rect 1225 18374 1241 18414
rect 1293 18374 2097 18414
rect 1225 18373 1239 18374
rect 1293 18373 1475 18374
rect 565 18361 767 18373
rect 801 18361 1003 18373
rect 1037 18361 1239 18373
rect 1273 18361 1475 18373
rect 565 18340 697 18361
rect 420 18317 697 18340
rect 380 18309 697 18317
rect 749 18309 765 18361
rect 817 18309 833 18361
rect 885 18309 901 18361
rect 953 18309 969 18361
rect 1021 18309 1037 18340
rect 1089 18309 1105 18361
rect 1157 18309 1173 18361
rect 1225 18340 1239 18361
rect 1293 18340 1475 18361
rect 1509 18340 1711 18374
rect 1745 18340 1947 18374
rect 1981 18373 2097 18374
rect 2149 18373 2165 18425
rect 2217 18373 2233 18425
rect 2285 18373 2301 18425
rect 2353 18373 2369 18425
rect 2421 18374 2437 18414
rect 2489 18373 2505 18425
rect 2557 18373 2573 18425
rect 2625 18373 2641 18425
rect 2693 18414 2891 18425
rect 2925 18442 3076 18448
rect 2925 18414 3036 18442
rect 2693 18408 3036 18414
rect 3070 18408 3076 18442
rect 2693 18374 3076 18408
rect 2693 18373 2891 18374
rect 1981 18361 2183 18373
rect 2217 18361 2419 18373
rect 2453 18361 2655 18373
rect 2689 18361 2891 18373
rect 1981 18340 2097 18361
rect 1225 18309 1241 18340
rect 1293 18309 2097 18340
rect 2149 18309 2165 18361
rect 2217 18309 2233 18361
rect 2285 18309 2301 18361
rect 2353 18309 2369 18361
rect 2421 18309 2437 18340
rect 2489 18309 2505 18361
rect 2557 18309 2573 18361
rect 2625 18309 2641 18361
rect 2693 18340 2891 18361
rect 2925 18370 3076 18374
rect 2925 18340 3036 18370
rect 2693 18336 3036 18340
rect 3070 18336 3076 18370
rect 2693 18309 3076 18336
rect 380 18300 3076 18309
rect 380 18279 531 18300
rect 380 18245 386 18279
rect 420 18266 531 18279
rect 565 18284 767 18300
rect 565 18266 587 18284
tri 587 18266 605 18284 nw
tri 727 18266 745 18284 ne
rect 745 18266 767 18284
rect 801 18284 1003 18300
rect 801 18266 823 18284
tri 823 18266 841 18284 nw
tri 963 18266 981 18284 ne
rect 981 18266 1003 18284
rect 1037 18284 1239 18300
rect 1037 18266 1059 18284
tri 1059 18266 1077 18284 nw
tri 1199 18266 1217 18284 ne
rect 1217 18266 1239 18284
rect 1273 18284 1475 18300
rect 1273 18266 1295 18284
tri 1295 18266 1313 18284 nw
tri 1435 18266 1453 18284 ne
rect 1453 18266 1475 18284
rect 1509 18284 1711 18300
rect 1509 18266 1531 18284
tri 1531 18266 1549 18284 nw
tri 1671 18266 1689 18284 ne
rect 1689 18266 1711 18284
rect 1745 18284 1947 18300
rect 1745 18266 1767 18284
tri 1767 18266 1785 18284 nw
tri 1907 18266 1925 18284 ne
rect 1925 18266 1947 18284
rect 1981 18284 2183 18300
rect 1981 18266 2003 18284
tri 2003 18266 2021 18284 nw
tri 2143 18266 2161 18284 ne
rect 2161 18266 2183 18284
rect 2217 18284 2419 18300
rect 2217 18266 2239 18284
tri 2239 18266 2257 18284 nw
tri 2379 18266 2397 18284 ne
rect 2397 18266 2419 18284
rect 2453 18284 2655 18300
rect 2453 18266 2475 18284
tri 2475 18266 2493 18284 nw
tri 2615 18266 2633 18284 ne
rect 2633 18266 2655 18284
rect 2689 18284 2891 18300
rect 2689 18266 2711 18284
tri 2711 18266 2729 18284 nw
tri 2851 18266 2869 18284 ne
rect 2869 18266 2891 18284
rect 2925 18298 3076 18300
rect 2925 18266 3036 18298
rect 420 18264 585 18266
tri 585 18264 587 18266 nw
tri 745 18264 747 18266 ne
rect 747 18264 821 18266
tri 821 18264 823 18266 nw
tri 981 18264 983 18266 ne
rect 983 18264 1057 18266
tri 1057 18264 1059 18266 nw
tri 1217 18264 1219 18266 ne
rect 1219 18264 1293 18266
tri 1293 18264 1295 18266 nw
tri 1453 18264 1455 18266 ne
rect 1455 18264 1529 18266
tri 1529 18264 1531 18266 nw
tri 1689 18264 1691 18266 ne
rect 1691 18264 1765 18266
tri 1765 18264 1767 18266 nw
tri 1925 18264 1927 18266 ne
rect 1927 18264 2001 18266
tri 2001 18264 2003 18266 nw
tri 2161 18264 2163 18266 ne
rect 2163 18264 2237 18266
tri 2237 18264 2239 18266 nw
tri 2397 18264 2399 18266 ne
rect 2399 18264 2473 18266
tri 2473 18264 2475 18266 nw
tri 2633 18264 2635 18266 ne
rect 2635 18264 2709 18266
tri 2709 18264 2711 18266 nw
tri 2869 18264 2871 18266 ne
rect 2871 18264 3036 18266
rect 3070 18264 3076 18298
rect 420 18245 571 18264
tri 571 18250 585 18264 nw
tri 747 18250 761 18264 ne
rect 380 18226 571 18245
rect 380 18207 531 18226
rect 380 18173 386 18207
rect 420 18192 531 18207
rect 565 18192 571 18226
rect 420 18173 571 18192
rect 380 18152 571 18173
rect 380 18135 531 18152
rect 380 18101 386 18135
rect 420 18118 531 18135
rect 565 18118 571 18152
rect 420 18101 571 18118
rect 380 18078 571 18101
rect 380 18063 531 18078
rect 380 18029 386 18063
rect 420 18044 531 18063
rect 565 18044 571 18078
rect 420 18029 571 18044
rect 380 18004 571 18029
rect 380 17991 531 18004
rect 380 17957 386 17991
rect 420 17970 531 17991
rect 565 17970 571 18004
rect 420 17957 571 17970
rect 380 17930 571 17957
rect 380 17919 531 17930
rect 380 17885 386 17919
rect 420 17896 531 17919
rect 565 17896 571 17930
rect 420 17885 571 17896
rect 380 17856 571 17885
rect 380 17847 531 17856
rect 380 17813 386 17847
rect 420 17822 531 17847
rect 565 17822 571 17856
rect 420 17813 571 17822
rect 380 17775 571 17813
rect 761 18226 807 18264
tri 807 18250 821 18264 nw
tri 983 18250 997 18264 ne
rect 761 18192 767 18226
rect 801 18192 807 18226
rect 761 18152 807 18192
rect 761 18118 767 18152
rect 801 18118 807 18152
rect 761 18078 807 18118
rect 761 18044 767 18078
rect 801 18044 807 18078
rect 761 18004 807 18044
rect 761 17970 767 18004
rect 801 17970 807 18004
rect 761 17930 807 17970
rect 761 17896 767 17930
rect 801 17896 807 17930
rect 761 17856 807 17896
rect 761 17822 767 17856
rect 801 17822 807 17856
rect 761 17810 807 17822
rect 997 18226 1043 18264
tri 1043 18250 1057 18264 nw
tri 1219 18250 1233 18264 ne
rect 997 18192 1003 18226
rect 1037 18192 1043 18226
rect 997 18152 1043 18192
rect 997 18118 1003 18152
rect 1037 18118 1043 18152
rect 997 18078 1043 18118
rect 997 18044 1003 18078
rect 1037 18044 1043 18078
rect 997 18004 1043 18044
rect 997 17970 1003 18004
rect 1037 17970 1043 18004
rect 997 17930 1043 17970
rect 997 17896 1003 17930
rect 1037 17896 1043 17930
rect 997 17856 1043 17896
rect 997 17822 1003 17856
rect 1037 17822 1043 17856
rect 997 17810 1043 17822
rect 1233 18226 1279 18264
tri 1279 18250 1293 18264 nw
tri 1455 18250 1469 18264 ne
rect 1233 18192 1239 18226
rect 1273 18192 1279 18226
rect 1233 18152 1279 18192
rect 1233 18118 1239 18152
rect 1273 18118 1279 18152
rect 1233 18078 1279 18118
rect 1233 18044 1239 18078
rect 1273 18044 1279 18078
rect 1233 18004 1279 18044
rect 1233 17970 1239 18004
rect 1273 17970 1279 18004
rect 1233 17930 1279 17970
rect 1233 17896 1239 17930
rect 1273 17896 1279 17930
rect 1233 17856 1279 17896
rect 1233 17822 1239 17856
rect 1273 17822 1279 17856
rect 1233 17810 1279 17822
rect 1469 18226 1515 18264
tri 1515 18250 1529 18264 nw
tri 1691 18250 1705 18264 ne
rect 1469 18192 1475 18226
rect 1509 18192 1515 18226
rect 1469 18152 1515 18192
rect 1469 18118 1475 18152
rect 1509 18118 1515 18152
rect 1469 18078 1515 18118
rect 1469 18044 1475 18078
rect 1509 18044 1515 18078
rect 1469 18004 1515 18044
rect 1469 17970 1475 18004
rect 1509 17970 1515 18004
rect 1469 17930 1515 17970
rect 1469 17896 1475 17930
rect 1509 17896 1515 17930
rect 1469 17856 1515 17896
rect 1469 17822 1475 17856
rect 1509 17822 1515 17856
rect 1469 17810 1515 17822
rect 1705 18226 1751 18264
tri 1751 18250 1765 18264 nw
tri 1927 18250 1941 18264 ne
rect 1705 18192 1711 18226
rect 1745 18192 1751 18226
rect 1705 18152 1751 18192
rect 1705 18118 1711 18152
rect 1745 18118 1751 18152
rect 1705 18078 1751 18118
rect 1705 18044 1711 18078
rect 1745 18044 1751 18078
rect 1705 18004 1751 18044
rect 1705 17970 1711 18004
rect 1745 17970 1751 18004
rect 1705 17930 1751 17970
rect 1705 17896 1711 17930
rect 1745 17896 1751 17930
rect 1705 17856 1751 17896
rect 1705 17822 1711 17856
rect 1745 17822 1751 17856
rect 1705 17810 1751 17822
rect 1941 18226 1987 18264
tri 1987 18250 2001 18264 nw
tri 2163 18250 2177 18264 ne
rect 1941 18192 1947 18226
rect 1981 18192 1987 18226
rect 1941 18152 1987 18192
rect 1941 18118 1947 18152
rect 1981 18118 1987 18152
rect 1941 18078 1987 18118
rect 1941 18044 1947 18078
rect 1981 18044 1987 18078
rect 1941 18004 1987 18044
rect 1941 17970 1947 18004
rect 1981 17970 1987 18004
rect 1941 17930 1987 17970
rect 1941 17896 1947 17930
rect 1981 17896 1987 17930
rect 1941 17856 1987 17896
rect 1941 17822 1947 17856
rect 1981 17822 1987 17856
rect 1941 17810 1987 17822
rect 2177 18226 2223 18264
tri 2223 18250 2237 18264 nw
tri 2399 18250 2413 18264 ne
rect 2177 18192 2183 18226
rect 2217 18192 2223 18226
rect 2177 18152 2223 18192
rect 2177 18118 2183 18152
rect 2217 18118 2223 18152
rect 2177 18078 2223 18118
rect 2177 18044 2183 18078
rect 2217 18044 2223 18078
rect 2177 18004 2223 18044
rect 2177 17970 2183 18004
rect 2217 17970 2223 18004
rect 2177 17930 2223 17970
rect 2177 17896 2183 17930
rect 2217 17896 2223 17930
rect 2177 17856 2223 17896
rect 2177 17822 2183 17856
rect 2217 17822 2223 17856
rect 2177 17810 2223 17822
rect 2413 18226 2459 18264
tri 2459 18250 2473 18264 nw
tri 2635 18250 2649 18264 ne
rect 2413 18192 2419 18226
rect 2453 18192 2459 18226
rect 2413 18152 2459 18192
rect 2413 18118 2419 18152
rect 2453 18118 2459 18152
rect 2413 18078 2459 18118
rect 2413 18044 2419 18078
rect 2453 18044 2459 18078
rect 2413 18004 2459 18044
rect 2413 17970 2419 18004
rect 2453 17970 2459 18004
rect 2413 17930 2459 17970
rect 2413 17896 2419 17930
rect 2453 17896 2459 17930
rect 2413 17856 2459 17896
rect 2413 17822 2419 17856
rect 2453 17822 2459 17856
rect 2413 17810 2459 17822
rect 2649 18226 2695 18264
tri 2695 18250 2709 18264 nw
tri 2871 18250 2885 18264 ne
rect 2649 18192 2655 18226
rect 2689 18192 2695 18226
rect 2649 18152 2695 18192
rect 2649 18118 2655 18152
rect 2689 18118 2695 18152
rect 2649 18078 2695 18118
rect 2649 18044 2655 18078
rect 2689 18044 2695 18078
rect 2649 18004 2695 18044
rect 2649 17970 2655 18004
rect 2689 17970 2695 18004
rect 2649 17930 2695 17970
rect 2649 17896 2655 17930
rect 2689 17896 2695 17930
rect 2649 17856 2695 17896
rect 2649 17822 2655 17856
rect 2689 17822 2695 17856
rect 2649 17810 2695 17822
rect 2885 18226 3076 18264
rect 2885 18192 2891 18226
rect 2925 18192 3036 18226
rect 3070 18192 3076 18226
rect 2885 18154 3076 18192
rect 2885 18152 3036 18154
rect 2885 18118 2891 18152
rect 2925 18120 3036 18152
rect 3070 18120 3076 18154
rect 2925 18118 3076 18120
rect 2885 18082 3076 18118
rect 2885 18078 3036 18082
rect 2885 18044 2891 18078
rect 2925 18048 3036 18078
rect 3070 18048 3076 18082
rect 2925 18044 3076 18048
rect 2885 18010 3076 18044
rect 2885 18004 3036 18010
rect 2885 17970 2891 18004
rect 2925 17976 3036 18004
rect 3070 17976 3076 18010
rect 2925 17970 3076 17976
rect 2885 17938 3076 17970
rect 2885 17930 3036 17938
rect 2885 17896 2891 17930
rect 2925 17904 3036 17930
rect 3070 17904 3076 17938
rect 2925 17896 3076 17904
rect 2885 17866 3076 17896
rect 2885 17856 3036 17866
rect 2885 17822 2891 17856
rect 2925 17832 3036 17856
rect 3070 17832 3076 17866
rect 2925 17822 3076 17832
rect 380 17741 386 17775
rect 420 17741 571 17775
rect 2885 17794 3076 17822
rect 380 17703 571 17741
rect 613 17754 1501 17763
rect 1553 17754 1569 17763
rect 1621 17754 1636 17763
rect 1688 17754 1703 17763
rect 1755 17754 1770 17763
rect 1822 17754 1837 17763
rect 1889 17754 2830 17763
rect 613 17720 625 17754
rect 659 17720 700 17754
rect 734 17720 775 17754
rect 809 17720 850 17754
rect 884 17720 925 17754
rect 959 17720 1000 17754
rect 1034 17720 1075 17754
rect 1109 17720 1150 17754
rect 1184 17720 1225 17754
rect 1259 17720 1300 17754
rect 1334 17720 1375 17754
rect 1409 17720 1450 17754
rect 1484 17720 1501 17754
rect 1559 17720 1569 17754
rect 1634 17720 1636 17754
rect 1889 17720 1896 17754
rect 1930 17720 1970 17754
rect 2004 17720 2044 17754
rect 2078 17720 2118 17754
rect 2152 17720 2192 17754
rect 2226 17720 2266 17754
rect 2300 17720 2340 17754
rect 2374 17720 2414 17754
rect 2448 17720 2488 17754
rect 2522 17720 2562 17754
rect 2596 17720 2636 17754
rect 2670 17720 2710 17754
rect 2744 17720 2784 17754
rect 2818 17720 2830 17754
rect 613 17711 1501 17720
rect 1553 17711 1569 17720
rect 1621 17711 1636 17720
rect 1688 17711 1703 17720
rect 1755 17711 1770 17720
rect 1822 17711 1837 17720
rect 1889 17711 2830 17720
rect 2885 17760 3036 17794
rect 3070 17760 3076 17794
rect 2885 17722 3076 17760
rect 380 17669 386 17703
rect 420 17669 571 17703
rect 380 17652 571 17669
rect 2885 17688 3036 17722
rect 3070 17688 3076 17722
rect 380 17631 531 17652
rect 380 17597 386 17631
rect 420 17618 531 17631
rect 565 17618 571 17652
rect 420 17597 571 17618
rect 380 17579 571 17597
rect 380 17559 531 17579
rect 380 17525 386 17559
rect 420 17545 531 17559
rect 565 17545 571 17579
rect 420 17525 571 17545
rect 380 17506 571 17525
rect 380 17487 531 17506
rect 380 17453 386 17487
rect 420 17472 531 17487
rect 565 17472 571 17506
rect 420 17453 571 17472
rect 380 17433 571 17453
rect 380 17415 531 17433
rect 380 17381 386 17415
rect 420 17399 531 17415
rect 565 17399 571 17433
rect 420 17381 571 17399
rect 380 17360 571 17381
rect 380 17343 531 17360
rect 380 17309 386 17343
rect 420 17326 531 17343
rect 565 17326 571 17360
rect 420 17309 571 17326
rect 380 17287 571 17309
rect 380 17271 531 17287
rect 380 17237 386 17271
rect 420 17253 531 17271
rect 565 17253 571 17287
rect 420 17237 571 17253
rect 380 17214 571 17237
rect 380 17199 531 17214
rect 380 17165 386 17199
rect 420 17180 531 17199
rect 565 17180 571 17214
rect 761 17652 807 17664
rect 761 17618 767 17652
rect 801 17618 807 17652
rect 761 17579 807 17618
rect 761 17545 767 17579
rect 801 17545 807 17579
rect 761 17506 807 17545
rect 761 17472 767 17506
rect 801 17472 807 17506
rect 761 17433 807 17472
rect 761 17399 767 17433
rect 801 17399 807 17433
rect 761 17360 807 17399
rect 761 17326 767 17360
rect 801 17326 807 17360
rect 761 17287 807 17326
rect 761 17253 767 17287
rect 801 17253 807 17287
rect 761 17214 807 17253
tri 571 17180 604 17213 sw
tri 728 17180 761 17213 se
rect 761 17180 767 17214
rect 801 17180 807 17214
rect 997 17652 1043 17664
rect 997 17618 1003 17652
rect 1037 17618 1043 17652
rect 997 17579 1043 17618
rect 997 17545 1003 17579
rect 1037 17545 1043 17579
rect 997 17506 1043 17545
rect 997 17472 1003 17506
rect 1037 17472 1043 17506
rect 997 17433 1043 17472
rect 997 17399 1003 17433
rect 1037 17399 1043 17433
rect 997 17360 1043 17399
rect 997 17326 1003 17360
rect 1037 17326 1043 17360
rect 997 17287 1043 17326
rect 997 17253 1003 17287
rect 1037 17253 1043 17287
rect 997 17214 1043 17253
tri 807 17180 840 17213 sw
tri 964 17180 997 17213 se
rect 997 17180 1003 17214
rect 1037 17180 1043 17214
rect 1233 17652 1279 17664
rect 1233 17618 1239 17652
rect 1273 17618 1279 17652
rect 1233 17579 1279 17618
rect 1233 17545 1239 17579
rect 1273 17545 1279 17579
rect 1233 17506 1279 17545
rect 1233 17472 1239 17506
rect 1273 17472 1279 17506
rect 1233 17433 1279 17472
rect 1233 17399 1239 17433
rect 1273 17399 1279 17433
rect 1233 17360 1279 17399
rect 1233 17326 1239 17360
rect 1273 17326 1279 17360
rect 1233 17287 1279 17326
rect 1233 17253 1239 17287
rect 1273 17253 1279 17287
rect 1233 17214 1279 17253
tri 1043 17180 1076 17213 sw
tri 1200 17180 1233 17213 se
rect 1233 17180 1239 17214
rect 1273 17180 1279 17214
rect 1469 17652 1515 17664
rect 1469 17618 1475 17652
rect 1509 17618 1515 17652
rect 1469 17579 1515 17618
rect 1469 17545 1475 17579
rect 1509 17545 1515 17579
rect 1469 17506 1515 17545
rect 1469 17472 1475 17506
rect 1509 17472 1515 17506
rect 1469 17433 1515 17472
rect 1469 17399 1475 17433
rect 1509 17399 1515 17433
rect 1469 17360 1515 17399
rect 1469 17326 1475 17360
rect 1509 17326 1515 17360
rect 1469 17287 1515 17326
rect 1469 17253 1475 17287
rect 1509 17253 1515 17287
rect 1469 17214 1515 17253
tri 1279 17180 1312 17213 sw
tri 1436 17180 1469 17213 se
rect 1469 17180 1475 17214
rect 1509 17180 1515 17214
rect 1705 17652 1751 17664
rect 1705 17618 1711 17652
rect 1745 17618 1751 17652
rect 1705 17579 1751 17618
rect 1705 17545 1711 17579
rect 1745 17545 1751 17579
rect 1705 17506 1751 17545
rect 1705 17472 1711 17506
rect 1745 17472 1751 17506
rect 1705 17433 1751 17472
rect 1705 17399 1711 17433
rect 1745 17399 1751 17433
rect 1705 17360 1751 17399
rect 1705 17326 1711 17360
rect 1745 17326 1751 17360
rect 1705 17287 1751 17326
rect 1705 17253 1711 17287
rect 1745 17253 1751 17287
rect 1705 17214 1751 17253
tri 1515 17180 1548 17213 sw
tri 1672 17180 1705 17213 se
rect 1705 17180 1711 17214
rect 1745 17180 1751 17214
rect 1941 17652 1987 17664
rect 1941 17618 1947 17652
rect 1981 17618 1987 17652
rect 1941 17579 1987 17618
rect 1941 17545 1947 17579
rect 1981 17545 1987 17579
rect 1941 17506 1987 17545
rect 1941 17472 1947 17506
rect 1981 17472 1987 17506
rect 1941 17433 1987 17472
rect 1941 17399 1947 17433
rect 1981 17399 1987 17433
rect 1941 17360 1987 17399
rect 1941 17326 1947 17360
rect 1981 17326 1987 17360
rect 1941 17287 1987 17326
rect 1941 17253 1947 17287
rect 1981 17253 1987 17287
rect 1941 17214 1987 17253
tri 1751 17180 1784 17213 sw
tri 1908 17180 1941 17213 se
rect 1941 17180 1947 17214
rect 1981 17180 1987 17214
rect 2177 17652 2223 17664
rect 2177 17618 2183 17652
rect 2217 17618 2223 17652
rect 2177 17579 2223 17618
rect 2177 17545 2183 17579
rect 2217 17545 2223 17579
rect 2177 17506 2223 17545
rect 2177 17472 2183 17506
rect 2217 17472 2223 17506
rect 2177 17433 2223 17472
rect 2177 17399 2183 17433
rect 2217 17399 2223 17433
rect 2177 17360 2223 17399
rect 2177 17326 2183 17360
rect 2217 17326 2223 17360
rect 2177 17287 2223 17326
rect 2177 17253 2183 17287
rect 2217 17253 2223 17287
rect 2177 17214 2223 17253
tri 1987 17180 2020 17213 sw
tri 2144 17180 2177 17213 se
rect 2177 17180 2183 17214
rect 2217 17180 2223 17214
rect 2413 17652 2459 17664
rect 2413 17618 2419 17652
rect 2453 17618 2459 17652
rect 2413 17579 2459 17618
rect 2413 17545 2419 17579
rect 2453 17545 2459 17579
rect 2413 17506 2459 17545
rect 2413 17472 2419 17506
rect 2453 17472 2459 17506
rect 2413 17433 2459 17472
rect 2413 17399 2419 17433
rect 2453 17399 2459 17433
rect 2413 17360 2459 17399
rect 2413 17326 2419 17360
rect 2453 17326 2459 17360
rect 2413 17287 2459 17326
rect 2413 17253 2419 17287
rect 2453 17253 2459 17287
rect 2413 17214 2459 17253
tri 2223 17180 2256 17213 sw
tri 2380 17180 2413 17213 se
rect 2413 17180 2419 17214
rect 2453 17180 2459 17214
rect 2649 17652 2695 17664
rect 2649 17618 2655 17652
rect 2689 17618 2695 17652
rect 2649 17579 2695 17618
rect 2649 17545 2655 17579
rect 2689 17545 2695 17579
rect 2649 17506 2695 17545
rect 2649 17472 2655 17506
rect 2689 17472 2695 17506
rect 2649 17433 2695 17472
rect 2649 17399 2655 17433
rect 2689 17399 2695 17433
rect 2649 17360 2695 17399
rect 2649 17326 2655 17360
rect 2689 17326 2695 17360
rect 2649 17287 2695 17326
rect 2649 17253 2655 17287
rect 2689 17253 2695 17287
rect 2649 17214 2695 17253
tri 2459 17180 2492 17213 sw
tri 2616 17180 2649 17213 se
rect 2649 17180 2655 17214
rect 2689 17180 2695 17214
rect 2885 17652 3076 17688
rect 2885 17618 2891 17652
rect 2925 17650 3076 17652
rect 2925 17618 3036 17650
rect 2885 17616 3036 17618
rect 3070 17616 3076 17650
rect 2885 17579 3076 17616
rect 2885 17545 2891 17579
rect 2925 17578 3076 17579
rect 2925 17545 3036 17578
rect 2885 17544 3036 17545
rect 3070 17544 3076 17578
rect 2885 17506 3076 17544
rect 2885 17472 2891 17506
rect 2925 17472 3036 17506
rect 3070 17472 3076 17506
rect 2885 17434 3076 17472
rect 2885 17433 3036 17434
rect 2885 17399 2891 17433
rect 2925 17400 3036 17433
rect 3070 17400 3076 17434
rect 2925 17399 3076 17400
rect 2885 17362 3076 17399
rect 2885 17360 3036 17362
rect 2885 17326 2891 17360
rect 2925 17328 3036 17360
rect 3070 17328 3076 17362
rect 2925 17326 3076 17328
rect 2885 17290 3076 17326
rect 2885 17287 3036 17290
rect 2885 17253 2891 17287
rect 2925 17256 3036 17287
rect 3070 17256 3076 17290
rect 2925 17253 3076 17256
rect 2885 17218 3076 17253
rect 2885 17214 3036 17218
tri 2695 17180 2728 17213 sw
tri 2852 17180 2885 17213 se
rect 2885 17180 2891 17214
rect 2925 17184 3036 17214
rect 3070 17184 3076 17218
rect 2925 17180 3076 17184
rect 420 17179 604 17180
tri 604 17179 605 17180 sw
tri 727 17179 728 17180 se
rect 728 17179 840 17180
tri 840 17179 841 17180 sw
tri 963 17179 964 17180 se
rect 964 17179 1076 17180
tri 1076 17179 1077 17180 sw
tri 1199 17179 1200 17180 se
rect 1200 17179 1312 17180
tri 1312 17179 1313 17180 sw
tri 1435 17179 1436 17180 se
rect 1436 17179 1548 17180
tri 1548 17179 1549 17180 sw
tri 1671 17179 1672 17180 se
rect 1672 17179 1784 17180
tri 1784 17179 1785 17180 sw
tri 1907 17179 1908 17180 se
rect 1908 17179 2020 17180
tri 2020 17179 2021 17180 sw
tri 2143 17179 2144 17180 se
rect 2144 17179 2256 17180
tri 2256 17179 2257 17180 sw
tri 2379 17179 2380 17180 se
rect 2380 17179 2492 17180
tri 2492 17179 2493 17180 sw
tri 2615 17179 2616 17180 se
rect 2616 17179 2728 17180
tri 2728 17179 2729 17180 sw
tri 2851 17179 2852 17180 se
rect 2852 17179 3076 17180
rect 420 17165 3076 17179
rect 380 17146 3076 17165
rect 380 17141 697 17146
rect 380 17127 531 17141
rect 380 17093 386 17127
rect 420 17107 531 17127
rect 565 17107 697 17141
rect 420 17094 697 17107
rect 749 17094 765 17146
rect 817 17094 833 17146
rect 885 17094 901 17146
rect 953 17094 969 17146
rect 1021 17141 1037 17146
rect 1021 17094 1037 17107
rect 1089 17094 1105 17146
rect 1157 17094 1173 17146
rect 1225 17141 1241 17146
rect 1293 17141 2097 17146
rect 1225 17107 1239 17141
rect 1293 17107 1475 17141
rect 1509 17107 1711 17141
rect 1745 17107 1947 17141
rect 1981 17107 2097 17141
rect 1225 17094 1241 17107
rect 1293 17094 2097 17107
rect 2149 17094 2165 17146
rect 2217 17094 2233 17146
rect 2285 17094 2301 17146
rect 2353 17094 2369 17146
rect 2421 17141 2437 17146
rect 2421 17094 2437 17107
rect 2489 17094 2505 17146
rect 2557 17094 2573 17146
rect 2625 17094 2641 17146
rect 2693 17141 3036 17146
rect 2693 17107 2891 17141
rect 2925 17112 3036 17141
rect 3070 17112 3076 17146
rect 2925 17107 3076 17112
rect 2693 17094 3076 17107
rect 420 17093 3076 17094
rect 380 17082 3076 17093
rect 380 17068 697 17082
rect 380 17055 531 17068
rect 380 17021 386 17055
rect 420 17034 531 17055
rect 565 17034 697 17068
rect 420 17030 697 17034
rect 749 17030 765 17082
rect 817 17030 833 17082
rect 885 17030 901 17082
rect 953 17030 969 17082
rect 1021 17068 1037 17082
rect 1021 17030 1037 17034
rect 1089 17030 1105 17082
rect 1157 17030 1173 17082
rect 1225 17068 1241 17082
rect 1293 17068 2097 17082
rect 1225 17034 1239 17068
rect 1293 17034 1475 17068
rect 1509 17034 1711 17068
rect 1745 17034 1947 17068
rect 1981 17034 2097 17068
rect 1225 17030 1241 17034
rect 1293 17030 2097 17034
rect 2149 17030 2165 17082
rect 2217 17030 2233 17082
rect 2285 17030 2301 17082
rect 2353 17030 2369 17082
rect 2421 17068 2437 17082
rect 2421 17030 2437 17034
rect 2489 17030 2505 17082
rect 2557 17030 2573 17082
rect 2625 17030 2641 17082
rect 2693 17074 3076 17082
rect 2693 17068 3036 17074
rect 2693 17034 2891 17068
rect 2925 17040 3036 17068
rect 3070 17040 3076 17074
rect 2925 17034 3076 17040
rect 2693 17030 3076 17034
rect 420 17021 3076 17030
rect 380 17018 3076 17021
rect 380 16995 697 17018
rect 380 16983 531 16995
rect 380 16949 386 16983
rect 420 16961 531 16983
rect 565 16966 697 16995
rect 749 16966 765 17018
rect 817 16966 833 17018
rect 885 16966 901 17018
rect 953 16966 969 17018
rect 1021 16995 1037 17018
rect 1089 16966 1105 17018
rect 1157 16966 1173 17018
rect 1225 16995 1241 17018
rect 1293 16995 2097 17018
rect 1225 16966 1239 16995
rect 1293 16966 1475 16995
rect 565 16961 767 16966
rect 801 16961 1003 16966
rect 1037 16961 1239 16966
rect 1273 16961 1475 16966
rect 1509 16961 1711 16995
rect 1745 16961 1947 16995
rect 1981 16966 2097 16995
rect 2149 16966 2165 17018
rect 2217 16966 2233 17018
rect 2285 16966 2301 17018
rect 2353 16966 2369 17018
rect 2421 16995 2437 17018
rect 2489 16966 2505 17018
rect 2557 16966 2573 17018
rect 2625 16966 2641 17018
rect 2693 17002 3076 17018
rect 2693 16995 3036 17002
rect 2693 16966 2891 16995
rect 1981 16961 2183 16966
rect 2217 16961 2419 16966
rect 2453 16961 2655 16966
rect 2689 16961 2891 16966
rect 2925 16968 3036 16995
rect 3070 16968 3076 17002
rect 2925 16961 3076 16968
rect 420 16954 3076 16961
rect 420 16949 697 16954
rect 380 16922 697 16949
rect 380 16911 531 16922
rect 380 16877 386 16911
rect 420 16888 531 16911
rect 565 16902 697 16922
rect 749 16902 765 16954
rect 817 16902 833 16954
rect 885 16902 901 16954
rect 953 16902 969 16954
rect 1021 16922 1037 16954
rect 1089 16902 1105 16954
rect 1157 16902 1173 16954
rect 1225 16922 1241 16954
rect 1293 16922 2097 16954
rect 1225 16902 1239 16922
rect 1293 16902 1475 16922
rect 565 16890 767 16902
rect 801 16890 1003 16902
rect 1037 16890 1239 16902
rect 1273 16890 1475 16902
rect 565 16888 697 16890
rect 420 16877 697 16888
rect 380 16849 697 16877
rect 380 16839 531 16849
rect 380 16805 386 16839
rect 420 16815 531 16839
rect 565 16838 697 16849
rect 749 16838 765 16890
rect 817 16838 833 16890
rect 885 16838 901 16890
rect 953 16838 969 16890
rect 1021 16849 1037 16888
rect 1089 16838 1105 16890
rect 1157 16838 1173 16890
rect 1225 16888 1239 16890
rect 1293 16888 1475 16890
rect 1509 16888 1711 16922
rect 1745 16888 1947 16922
rect 1981 16902 2097 16922
rect 2149 16902 2165 16954
rect 2217 16902 2233 16954
rect 2285 16902 2301 16954
rect 2353 16902 2369 16954
rect 2421 16922 2437 16954
rect 2489 16902 2505 16954
rect 2557 16902 2573 16954
rect 2625 16902 2641 16954
rect 2693 16930 3076 16954
rect 2693 16922 3036 16930
rect 2693 16902 2891 16922
rect 1981 16890 2183 16902
rect 2217 16890 2419 16902
rect 2453 16890 2655 16902
rect 2689 16890 2891 16902
rect 1981 16888 2097 16890
rect 1225 16849 1241 16888
rect 1293 16849 2097 16888
rect 1225 16838 1239 16849
rect 1293 16838 1475 16849
rect 565 16826 767 16838
rect 801 16826 1003 16838
rect 1037 16826 1239 16838
rect 1273 16826 1475 16838
rect 565 16815 697 16826
rect 420 16805 697 16815
rect 380 16776 697 16805
rect 380 16767 531 16776
rect 380 16733 386 16767
rect 420 16742 531 16767
rect 565 16774 697 16776
rect 749 16774 765 16826
rect 817 16774 833 16826
rect 885 16774 901 16826
rect 953 16774 969 16826
rect 1021 16776 1037 16815
rect 1089 16774 1105 16826
rect 1157 16774 1173 16826
rect 1225 16815 1239 16826
rect 1293 16815 1475 16826
rect 1509 16815 1711 16849
rect 1745 16815 1947 16849
rect 1981 16838 2097 16849
rect 2149 16838 2165 16890
rect 2217 16838 2233 16890
rect 2285 16838 2301 16890
rect 2353 16838 2369 16890
rect 2421 16849 2437 16888
rect 2489 16838 2505 16890
rect 2557 16838 2573 16890
rect 2625 16838 2641 16890
rect 2693 16888 2891 16890
rect 2925 16896 3036 16922
rect 3070 16896 3076 16930
rect 2925 16888 3076 16896
rect 2693 16858 3076 16888
rect 2693 16849 3036 16858
rect 2693 16838 2891 16849
rect 1981 16826 2183 16838
rect 2217 16826 2419 16838
rect 2453 16826 2655 16838
rect 2689 16826 2891 16838
rect 1981 16815 2097 16826
rect 1225 16776 1241 16815
rect 1293 16776 2097 16815
rect 1225 16774 1239 16776
rect 1293 16774 1475 16776
rect 565 16762 767 16774
rect 801 16762 1003 16774
rect 1037 16762 1239 16774
rect 1273 16762 1475 16774
rect 565 16742 697 16762
rect 420 16733 697 16742
rect 380 16710 697 16733
rect 749 16710 765 16762
rect 817 16710 833 16762
rect 885 16710 901 16762
rect 953 16710 969 16762
rect 1021 16710 1037 16742
rect 1089 16710 1105 16762
rect 1157 16710 1173 16762
rect 1225 16742 1239 16762
rect 1293 16742 1475 16762
rect 1509 16742 1711 16776
rect 1745 16742 1947 16776
rect 1981 16774 2097 16776
rect 2149 16774 2165 16826
rect 2217 16774 2233 16826
rect 2285 16774 2301 16826
rect 2353 16774 2369 16826
rect 2421 16776 2437 16815
rect 2489 16774 2505 16826
rect 2557 16774 2573 16826
rect 2625 16774 2641 16826
rect 2693 16815 2891 16826
rect 2925 16824 3036 16849
rect 3070 16824 3076 16858
rect 2925 16815 3076 16824
rect 2693 16786 3076 16815
rect 2693 16776 3036 16786
rect 2693 16774 2891 16776
rect 1981 16762 2183 16774
rect 2217 16762 2419 16774
rect 2453 16762 2655 16774
rect 2689 16762 2891 16774
rect 1981 16742 2097 16762
rect 1225 16710 1241 16742
rect 1293 16710 2097 16742
rect 2149 16710 2165 16762
rect 2217 16710 2233 16762
rect 2285 16710 2301 16762
rect 2353 16710 2369 16762
rect 2421 16710 2437 16742
rect 2489 16710 2505 16762
rect 2557 16710 2573 16762
rect 2625 16710 2641 16762
rect 2693 16742 2891 16762
rect 2925 16752 3036 16776
rect 3070 16752 3076 16786
rect 2925 16742 3076 16752
rect 2693 16714 3076 16742
rect 2693 16710 3036 16714
rect 380 16702 3036 16710
rect 380 16695 531 16702
rect 380 16661 386 16695
rect 420 16668 531 16695
rect 565 16698 767 16702
rect 801 16698 1003 16702
rect 1037 16698 1239 16702
rect 1273 16698 1475 16702
rect 565 16668 697 16698
rect 420 16661 697 16668
rect 380 16646 697 16661
rect 749 16646 765 16698
rect 817 16646 833 16698
rect 885 16646 901 16698
rect 953 16646 969 16698
rect 1021 16646 1037 16668
rect 1089 16646 1105 16698
rect 1157 16646 1173 16698
rect 1225 16668 1239 16698
rect 1293 16668 1475 16698
rect 1509 16668 1711 16702
rect 1745 16668 1947 16702
rect 1981 16698 2183 16702
rect 2217 16698 2419 16702
rect 2453 16698 2655 16702
rect 2689 16698 2891 16702
rect 1981 16668 2097 16698
rect 1225 16646 1241 16668
rect 1293 16646 2097 16668
rect 2149 16646 2165 16698
rect 2217 16646 2233 16698
rect 2285 16646 2301 16698
rect 2353 16646 2369 16698
rect 2421 16646 2437 16668
rect 2489 16646 2505 16698
rect 2557 16646 2573 16698
rect 2625 16646 2641 16698
rect 2693 16668 2891 16698
rect 2925 16680 3036 16702
rect 3070 16680 3076 16714
rect 2925 16668 3076 16680
rect 2693 16646 3076 16668
rect 380 16642 3076 16646
rect 380 16634 3036 16642
rect 380 16628 697 16634
rect 380 16623 531 16628
rect 380 16589 386 16623
rect 420 16594 531 16623
rect 565 16594 697 16628
rect 420 16589 697 16594
rect 380 16582 697 16589
rect 749 16582 765 16634
rect 817 16582 833 16634
rect 885 16582 901 16634
rect 953 16582 969 16634
rect 1021 16628 1037 16634
rect 1021 16582 1037 16594
rect 1089 16582 1105 16634
rect 1157 16582 1173 16634
rect 1225 16628 1241 16634
rect 1293 16628 2097 16634
rect 1225 16594 1239 16628
rect 1293 16594 1475 16628
rect 1509 16594 1711 16628
rect 1745 16594 1947 16628
rect 1981 16594 2097 16628
rect 1225 16582 1241 16594
rect 1293 16582 2097 16594
rect 2149 16582 2165 16634
rect 2217 16582 2233 16634
rect 2285 16582 2301 16634
rect 2353 16582 2369 16634
rect 2421 16628 2437 16634
rect 2421 16582 2437 16594
rect 2489 16582 2505 16634
rect 2557 16582 2573 16634
rect 2625 16582 2641 16634
rect 2693 16628 3036 16634
rect 2693 16594 2891 16628
rect 2925 16608 3036 16628
rect 3070 16608 3076 16642
rect 2925 16594 3076 16608
rect 2693 16582 3076 16594
rect 380 16570 3076 16582
rect 380 16554 697 16570
rect 380 16551 531 16554
rect 380 16517 386 16551
rect 420 16520 531 16551
rect 565 16520 697 16554
rect 420 16518 697 16520
rect 749 16518 765 16570
rect 817 16518 833 16570
rect 885 16518 901 16570
rect 953 16518 969 16570
rect 1021 16554 1037 16570
rect 1021 16518 1037 16520
rect 1089 16518 1105 16570
rect 1157 16518 1173 16570
rect 1225 16554 1241 16570
rect 1293 16554 2097 16570
rect 1225 16520 1239 16554
rect 1293 16520 1475 16554
rect 1509 16520 1711 16554
rect 1745 16520 1947 16554
rect 1981 16520 2097 16554
rect 1225 16518 1241 16520
rect 1293 16518 2097 16520
rect 2149 16518 2165 16570
rect 2217 16518 2233 16570
rect 2285 16518 2301 16570
rect 2353 16518 2369 16570
rect 2421 16554 2437 16570
rect 2421 16518 2437 16520
rect 2489 16518 2505 16570
rect 2557 16518 2573 16570
rect 2625 16518 2641 16570
rect 2693 16554 3036 16570
rect 2693 16520 2891 16554
rect 2925 16536 3036 16554
rect 3070 16536 3076 16570
rect 2925 16520 3076 16536
rect 2693 16518 3076 16520
rect 420 16517 3076 16518
rect 380 16506 3076 16517
rect 380 16480 697 16506
rect 380 16479 531 16480
rect 380 16445 386 16479
rect 420 16446 531 16479
rect 565 16454 697 16480
rect 749 16454 765 16506
rect 817 16454 833 16506
rect 885 16454 901 16506
rect 953 16454 969 16506
rect 1021 16480 1037 16506
rect 1089 16454 1105 16506
rect 1157 16454 1173 16506
rect 1225 16480 1241 16506
rect 1293 16480 2097 16506
rect 1225 16454 1239 16480
rect 1293 16454 1475 16480
rect 565 16446 767 16454
rect 801 16446 1003 16454
rect 1037 16446 1239 16454
rect 1273 16446 1475 16454
rect 1509 16446 1711 16480
rect 1745 16446 1947 16480
rect 1981 16454 2097 16480
rect 2149 16454 2165 16506
rect 2217 16454 2233 16506
rect 2285 16454 2301 16506
rect 2353 16454 2369 16506
rect 2421 16480 2437 16506
rect 2489 16454 2505 16506
rect 2557 16454 2573 16506
rect 2625 16454 2641 16506
rect 2693 16498 3076 16506
rect 2693 16480 3036 16498
rect 2693 16454 2891 16480
rect 1981 16446 2183 16454
rect 2217 16446 2419 16454
rect 2453 16446 2655 16454
rect 2689 16446 2891 16454
rect 2925 16464 3036 16480
rect 3070 16464 3076 16498
rect 2925 16446 3076 16464
rect 420 16445 3076 16446
rect 380 16442 3076 16445
rect 380 16407 697 16442
rect 380 16373 386 16407
rect 420 16406 697 16407
rect 420 16373 531 16406
rect 380 16372 531 16373
rect 565 16390 697 16406
rect 749 16390 765 16442
rect 817 16390 833 16442
rect 885 16390 901 16442
rect 953 16390 969 16442
rect 1021 16406 1037 16442
rect 1089 16390 1105 16442
rect 1157 16390 1173 16442
rect 1225 16406 1241 16442
rect 1293 16406 2097 16442
rect 1225 16390 1239 16406
rect 1293 16390 1475 16406
rect 565 16378 767 16390
rect 801 16378 1003 16390
rect 1037 16378 1239 16390
rect 1273 16378 1475 16390
rect 565 16372 697 16378
rect 380 16335 697 16372
rect 380 16301 386 16335
rect 420 16332 697 16335
rect 420 16301 531 16332
rect 380 16298 531 16301
rect 565 16326 697 16332
rect 749 16326 765 16378
rect 817 16326 833 16378
rect 885 16326 901 16378
rect 953 16326 969 16378
rect 1021 16332 1037 16372
rect 1089 16326 1105 16378
rect 1157 16326 1173 16378
rect 1225 16372 1239 16378
rect 1293 16372 1475 16378
rect 1509 16372 1711 16406
rect 1745 16372 1947 16406
rect 1981 16390 2097 16406
rect 2149 16390 2165 16442
rect 2217 16390 2233 16442
rect 2285 16390 2301 16442
rect 2353 16390 2369 16442
rect 2421 16406 2437 16442
rect 2489 16390 2505 16442
rect 2557 16390 2573 16442
rect 2625 16390 2641 16442
rect 2693 16426 3076 16442
rect 2693 16406 3036 16426
rect 2693 16390 2891 16406
rect 1981 16378 2183 16390
rect 2217 16378 2419 16390
rect 2453 16378 2655 16390
rect 2689 16378 2891 16390
rect 1981 16372 2097 16378
rect 1225 16332 1241 16372
rect 1293 16332 2097 16372
rect 1225 16326 1239 16332
rect 1293 16326 1475 16332
rect 565 16314 767 16326
rect 801 16314 1003 16326
rect 1037 16314 1239 16326
rect 1273 16314 1475 16326
rect 565 16298 697 16314
rect 380 16263 697 16298
rect 380 16229 386 16263
rect 420 16262 697 16263
rect 749 16262 765 16314
rect 817 16262 833 16314
rect 885 16262 901 16314
rect 953 16262 969 16314
rect 1021 16262 1037 16298
rect 1089 16262 1105 16314
rect 1157 16262 1173 16314
rect 1225 16298 1239 16314
rect 1293 16298 1475 16314
rect 1509 16298 1711 16332
rect 1745 16298 1947 16332
rect 1981 16326 2097 16332
rect 2149 16326 2165 16378
rect 2217 16326 2233 16378
rect 2285 16326 2301 16378
rect 2353 16326 2369 16378
rect 2421 16332 2437 16372
rect 2489 16326 2505 16378
rect 2557 16326 2573 16378
rect 2625 16326 2641 16378
rect 2693 16372 2891 16378
rect 2925 16392 3036 16406
rect 3070 16392 3076 16426
rect 2925 16372 3076 16392
rect 2693 16354 3076 16372
rect 2693 16332 3036 16354
rect 2693 16326 2891 16332
rect 1981 16314 2183 16326
rect 2217 16314 2419 16326
rect 2453 16314 2655 16326
rect 2689 16314 2891 16326
rect 1981 16298 2097 16314
rect 1225 16262 1241 16298
rect 1293 16262 2097 16298
rect 2149 16262 2165 16314
rect 2217 16262 2233 16314
rect 2285 16262 2301 16314
rect 2353 16262 2369 16314
rect 2421 16262 2437 16298
rect 2489 16262 2505 16314
rect 2557 16262 2573 16314
rect 2625 16262 2641 16314
rect 2693 16298 2891 16314
rect 2925 16320 3036 16332
rect 3070 16320 3076 16354
rect 2925 16298 3076 16320
rect 2693 16282 3076 16298
rect 2693 16262 3036 16282
rect 420 16258 3036 16262
rect 420 16229 531 16258
rect 380 16224 531 16229
rect 565 16250 767 16258
rect 801 16250 1003 16258
rect 1037 16250 1239 16258
rect 1273 16250 1475 16258
rect 565 16224 697 16250
rect 380 16198 697 16224
rect 749 16198 765 16250
rect 817 16198 833 16250
rect 885 16198 901 16250
rect 953 16198 969 16250
rect 1021 16198 1037 16224
rect 1089 16198 1105 16250
rect 1157 16198 1173 16250
rect 1225 16224 1239 16250
rect 1293 16224 1475 16250
rect 1509 16224 1711 16258
rect 1745 16224 1947 16258
rect 1981 16250 2183 16258
rect 2217 16250 2419 16258
rect 2453 16250 2655 16258
rect 2689 16250 2891 16258
rect 1981 16224 2097 16250
rect 1225 16198 1241 16224
rect 1293 16198 2097 16224
rect 2149 16198 2165 16250
rect 2217 16198 2233 16250
rect 2285 16198 2301 16250
rect 2353 16198 2369 16250
rect 2421 16198 2437 16224
rect 2489 16198 2505 16250
rect 2557 16198 2573 16250
rect 2625 16198 2641 16250
rect 2693 16224 2891 16250
rect 2925 16248 3036 16258
rect 3070 16248 3076 16282
rect 2925 16224 3076 16248
rect 2693 16210 3076 16224
rect 2693 16198 3036 16210
rect 380 16191 3036 16198
rect 380 16157 386 16191
rect 420 16184 3036 16191
rect 420 16157 531 16184
rect 380 16150 531 16157
rect 565 16179 767 16184
rect 565 16150 576 16179
tri 576 16150 605 16179 nw
tri 727 16150 756 16179 ne
rect 756 16150 767 16179
rect 801 16179 1003 16184
rect 801 16150 812 16179
tri 812 16150 841 16179 nw
tri 963 16150 992 16179 ne
rect 992 16150 1003 16179
rect 1037 16179 1239 16184
rect 1037 16150 1048 16179
tri 1048 16150 1077 16179 nw
tri 1199 16150 1228 16179 ne
rect 1228 16150 1239 16179
rect 1273 16179 1475 16184
rect 1273 16150 1284 16179
tri 1284 16150 1313 16179 nw
tri 1435 16150 1464 16179 ne
rect 1464 16150 1475 16179
rect 1509 16179 1711 16184
rect 1509 16150 1520 16179
tri 1520 16150 1549 16179 nw
tri 1671 16150 1700 16179 ne
rect 1700 16150 1711 16179
rect 1745 16179 1947 16184
rect 1745 16150 1756 16179
tri 1756 16150 1785 16179 nw
tri 1907 16150 1936 16179 ne
rect 1936 16150 1947 16179
rect 1981 16179 2183 16184
rect 1981 16150 1992 16179
tri 1992 16150 2021 16179 nw
tri 2143 16150 2172 16179 ne
rect 2172 16150 2183 16179
rect 2217 16179 2419 16184
rect 2217 16150 2228 16179
tri 2228 16150 2257 16179 nw
tri 2379 16150 2408 16179 ne
rect 2408 16150 2419 16179
rect 2453 16179 2655 16184
rect 2453 16150 2464 16179
tri 2464 16150 2493 16179 nw
tri 2615 16150 2644 16179 ne
rect 2644 16150 2655 16179
rect 2689 16179 2891 16184
rect 2689 16150 2700 16179
tri 2700 16150 2729 16179 nw
tri 2851 16150 2880 16179 ne
rect 2880 16150 2891 16179
rect 2925 16176 3036 16184
rect 3070 16176 3076 16210
rect 2925 16150 3076 16176
rect 380 16119 571 16150
tri 571 16145 576 16150 nw
tri 756 16145 761 16150 ne
rect 380 16085 386 16119
rect 420 16110 571 16119
rect 420 16085 531 16110
rect 380 16076 531 16085
rect 565 16076 571 16110
rect 380 16047 571 16076
rect 380 16013 386 16047
rect 420 16036 571 16047
rect 420 16013 531 16036
rect 380 16002 531 16013
rect 565 16002 571 16036
rect 380 15975 571 16002
rect 380 15941 386 15975
rect 420 15962 571 15975
rect 420 15941 531 15962
rect 380 15928 531 15941
rect 565 15928 571 15962
rect 380 15903 571 15928
rect 380 15869 386 15903
rect 420 15888 571 15903
rect 420 15869 531 15888
rect 380 15854 531 15869
rect 565 15854 571 15888
rect 380 15831 571 15854
rect 380 15797 386 15831
rect 420 15814 571 15831
rect 420 15797 531 15814
rect 380 15780 531 15797
rect 565 15780 571 15814
rect 380 15759 571 15780
rect 380 15725 386 15759
rect 420 15740 571 15759
rect 420 15725 531 15740
rect 380 15706 531 15725
rect 565 15706 571 15740
rect 380 15687 571 15706
rect 761 16110 807 16150
tri 807 16145 812 16150 nw
tri 992 16145 997 16150 ne
rect 761 16076 767 16110
rect 801 16076 807 16110
rect 761 16036 807 16076
rect 761 16002 767 16036
rect 801 16002 807 16036
rect 761 15962 807 16002
rect 761 15928 767 15962
rect 801 15928 807 15962
rect 761 15888 807 15928
rect 761 15854 767 15888
rect 801 15854 807 15888
rect 761 15814 807 15854
rect 761 15780 767 15814
rect 801 15780 807 15814
rect 761 15740 807 15780
rect 761 15706 767 15740
rect 801 15706 807 15740
rect 761 15694 807 15706
rect 997 16110 1043 16150
tri 1043 16145 1048 16150 nw
tri 1228 16145 1233 16150 ne
rect 997 16076 1003 16110
rect 1037 16076 1043 16110
rect 997 16036 1043 16076
rect 997 16002 1003 16036
rect 1037 16002 1043 16036
rect 997 15962 1043 16002
rect 997 15928 1003 15962
rect 1037 15928 1043 15962
rect 997 15888 1043 15928
rect 997 15854 1003 15888
rect 1037 15854 1043 15888
rect 997 15814 1043 15854
rect 997 15780 1003 15814
rect 1037 15780 1043 15814
rect 997 15740 1043 15780
rect 997 15706 1003 15740
rect 1037 15706 1043 15740
rect 997 15694 1043 15706
rect 1233 16110 1279 16150
tri 1279 16145 1284 16150 nw
tri 1464 16145 1469 16150 ne
rect 1233 16076 1239 16110
rect 1273 16076 1279 16110
rect 1233 16036 1279 16076
rect 1233 16002 1239 16036
rect 1273 16002 1279 16036
rect 1233 15962 1279 16002
rect 1233 15928 1239 15962
rect 1273 15928 1279 15962
rect 1233 15888 1279 15928
rect 1233 15854 1239 15888
rect 1273 15854 1279 15888
rect 1233 15814 1279 15854
rect 1233 15780 1239 15814
rect 1273 15780 1279 15814
rect 1233 15740 1279 15780
rect 1233 15706 1239 15740
rect 1273 15706 1279 15740
rect 1233 15694 1279 15706
rect 1469 16110 1515 16150
tri 1515 16145 1520 16150 nw
tri 1700 16145 1705 16150 ne
rect 1469 16076 1475 16110
rect 1509 16076 1515 16110
rect 1469 16036 1515 16076
rect 1469 16002 1475 16036
rect 1509 16002 1515 16036
rect 1469 15962 1515 16002
rect 1469 15928 1475 15962
rect 1509 15928 1515 15962
rect 1469 15888 1515 15928
rect 1469 15854 1475 15888
rect 1509 15854 1515 15888
rect 1469 15814 1515 15854
rect 1469 15780 1475 15814
rect 1509 15780 1515 15814
rect 1469 15740 1515 15780
rect 1469 15706 1475 15740
rect 1509 15706 1515 15740
rect 1469 15694 1515 15706
rect 1705 16110 1751 16150
tri 1751 16145 1756 16150 nw
tri 1936 16145 1941 16150 ne
rect 1705 16076 1711 16110
rect 1745 16076 1751 16110
rect 1705 16036 1751 16076
rect 1705 16002 1711 16036
rect 1745 16002 1751 16036
rect 1705 15962 1751 16002
rect 1705 15928 1711 15962
rect 1745 15928 1751 15962
rect 1705 15888 1751 15928
rect 1705 15854 1711 15888
rect 1745 15854 1751 15888
rect 1705 15814 1751 15854
rect 1705 15780 1711 15814
rect 1745 15780 1751 15814
rect 1705 15740 1751 15780
rect 1705 15706 1711 15740
rect 1745 15706 1751 15740
rect 1705 15694 1751 15706
rect 1941 16110 1987 16150
tri 1987 16145 1992 16150 nw
tri 2172 16145 2177 16150 ne
rect 1941 16076 1947 16110
rect 1981 16076 1987 16110
rect 1941 16036 1987 16076
rect 1941 16002 1947 16036
rect 1981 16002 1987 16036
rect 1941 15962 1987 16002
rect 1941 15928 1947 15962
rect 1981 15928 1987 15962
rect 1941 15888 1987 15928
rect 1941 15854 1947 15888
rect 1981 15854 1987 15888
rect 1941 15814 1987 15854
rect 1941 15780 1947 15814
rect 1981 15780 1987 15814
rect 1941 15740 1987 15780
rect 1941 15706 1947 15740
rect 1981 15706 1987 15740
rect 1941 15694 1987 15706
rect 2177 16110 2223 16150
tri 2223 16145 2228 16150 nw
tri 2408 16145 2413 16150 ne
rect 2177 16076 2183 16110
rect 2217 16076 2223 16110
rect 2177 16036 2223 16076
rect 2177 16002 2183 16036
rect 2217 16002 2223 16036
rect 2177 15962 2223 16002
rect 2177 15928 2183 15962
rect 2217 15928 2223 15962
rect 2177 15888 2223 15928
rect 2177 15854 2183 15888
rect 2217 15854 2223 15888
rect 2177 15814 2223 15854
rect 2177 15780 2183 15814
rect 2217 15780 2223 15814
rect 2177 15740 2223 15780
rect 2177 15706 2183 15740
rect 2217 15706 2223 15740
rect 2177 15694 2223 15706
rect 2413 16110 2459 16150
tri 2459 16145 2464 16150 nw
tri 2644 16145 2649 16150 ne
rect 2413 16076 2419 16110
rect 2453 16076 2459 16110
rect 2413 16036 2459 16076
rect 2413 16002 2419 16036
rect 2453 16002 2459 16036
rect 2413 15962 2459 16002
rect 2413 15928 2419 15962
rect 2453 15928 2459 15962
rect 2413 15888 2459 15928
rect 2413 15854 2419 15888
rect 2453 15854 2459 15888
rect 2413 15814 2459 15854
rect 2413 15780 2419 15814
rect 2453 15780 2459 15814
rect 2413 15740 2459 15780
rect 2413 15706 2419 15740
rect 2453 15706 2459 15740
rect 2413 15694 2459 15706
rect 2649 16110 2695 16150
tri 2695 16145 2700 16150 nw
tri 2880 16145 2885 16150 ne
rect 2649 16076 2655 16110
rect 2689 16076 2695 16110
rect 2649 16036 2695 16076
rect 2649 16002 2655 16036
rect 2689 16002 2695 16036
rect 2649 15962 2695 16002
rect 2649 15928 2655 15962
rect 2689 15928 2695 15962
rect 2649 15888 2695 15928
rect 2649 15854 2655 15888
rect 2689 15854 2695 15888
rect 2649 15814 2695 15854
rect 2649 15780 2655 15814
rect 2689 15780 2695 15814
rect 2649 15740 2695 15780
rect 2649 15706 2655 15740
rect 2689 15706 2695 15740
rect 2649 15694 2695 15706
rect 2885 16138 3076 16150
rect 2885 16110 3036 16138
rect 2885 16076 2891 16110
rect 2925 16104 3036 16110
rect 3070 16104 3076 16138
rect 2925 16076 3076 16104
rect 2885 16066 3076 16076
rect 2885 16036 3036 16066
rect 2885 16002 2891 16036
rect 2925 16032 3036 16036
rect 3070 16032 3076 16066
rect 2925 16002 3076 16032
rect 2885 15994 3076 16002
rect 2885 15962 3036 15994
rect 2885 15928 2891 15962
rect 2925 15960 3036 15962
rect 3070 15960 3076 15994
rect 2925 15928 3076 15960
rect 2885 15922 3076 15928
rect 2885 15888 3036 15922
rect 3070 15888 3076 15922
rect 2885 15854 2891 15888
rect 2925 15854 3076 15888
rect 2885 15850 3076 15854
rect 2885 15816 3036 15850
rect 3070 15816 3076 15850
rect 2885 15814 3076 15816
rect 2885 15780 2891 15814
rect 2925 15780 3076 15814
rect 2885 15778 3076 15780
rect 2885 15744 3036 15778
rect 3070 15744 3076 15778
rect 2885 15740 3076 15744
rect 2885 15706 2891 15740
rect 2925 15706 3076 15740
rect 380 15653 386 15687
rect 420 15653 571 15687
rect 380 15615 571 15653
rect 2885 15672 3036 15706
rect 3070 15672 3076 15706
rect 2885 15634 3076 15672
rect 380 15581 386 15615
rect 420 15581 571 15615
rect 613 15624 1501 15633
rect 1553 15624 1569 15633
rect 1621 15624 1636 15633
rect 1688 15624 1703 15633
rect 1755 15624 1770 15633
rect 1822 15624 1837 15633
rect 1889 15624 2830 15633
rect 613 15590 625 15624
rect 659 15590 700 15624
rect 734 15590 775 15624
rect 809 15590 850 15624
rect 884 15590 925 15624
rect 959 15590 1000 15624
rect 1034 15590 1075 15624
rect 1109 15590 1150 15624
rect 1184 15590 1225 15624
rect 1259 15590 1300 15624
rect 1334 15590 1375 15624
rect 1409 15590 1450 15624
rect 1484 15590 1501 15624
rect 1559 15590 1569 15624
rect 1634 15590 1636 15624
rect 1889 15590 1896 15624
rect 1930 15590 1970 15624
rect 2004 15590 2044 15624
rect 2078 15590 2118 15624
rect 2152 15590 2192 15624
rect 2226 15590 2266 15624
rect 2300 15590 2340 15624
rect 2374 15590 2414 15624
rect 2448 15590 2488 15624
rect 2522 15590 2562 15624
rect 2596 15590 2636 15624
rect 2670 15590 2710 15624
rect 2744 15590 2784 15624
rect 2818 15590 2830 15624
rect 613 15581 1501 15590
rect 1553 15581 1569 15590
rect 1621 15581 1636 15590
rect 1688 15581 1703 15590
rect 1755 15581 1770 15590
rect 1822 15581 1837 15590
rect 1889 15581 2830 15590
rect 2885 15600 3036 15634
rect 3070 15600 3076 15634
rect 380 15543 571 15581
rect 380 15509 386 15543
rect 420 15509 571 15543
rect 2885 15562 3076 15600
rect 2885 15528 3036 15562
rect 3070 15528 3076 15562
rect 380 15508 571 15509
rect 380 15474 531 15508
rect 565 15474 571 15508
rect 380 15471 571 15474
rect 380 15437 386 15471
rect 420 15437 571 15471
rect 380 15435 571 15437
rect 380 15401 531 15435
rect 565 15401 571 15435
rect 380 15399 571 15401
rect 380 15365 386 15399
rect 420 15365 571 15399
rect 380 15362 571 15365
rect 380 15328 531 15362
rect 565 15328 571 15362
rect 380 15327 571 15328
rect 380 15293 386 15327
rect 420 15293 571 15327
rect 380 15289 571 15293
rect 380 15255 531 15289
rect 565 15255 571 15289
rect 380 15221 386 15255
rect 420 15221 571 15255
rect 380 15216 571 15221
rect 380 15183 531 15216
rect 380 15149 386 15183
rect 420 15182 531 15183
rect 565 15182 571 15216
rect 420 15149 571 15182
rect 380 15143 571 15149
rect 380 15111 531 15143
rect 380 15077 386 15111
rect 420 15109 531 15111
rect 565 15109 571 15143
rect 420 15077 571 15109
rect 380 15072 571 15077
rect 761 15508 807 15520
rect 761 15474 767 15508
rect 801 15474 807 15508
rect 761 15435 807 15474
rect 761 15401 767 15435
rect 801 15401 807 15435
rect 761 15362 807 15401
rect 761 15328 767 15362
rect 801 15328 807 15362
rect 761 15289 807 15328
rect 761 15255 767 15289
rect 801 15255 807 15289
rect 761 15216 807 15255
rect 761 15182 767 15216
rect 801 15182 807 15216
rect 761 15143 807 15182
rect 761 15109 767 15143
rect 801 15109 807 15143
tri 571 15072 574 15075 sw
tri 758 15072 761 15075 se
rect 761 15072 807 15109
rect 997 15508 1043 15520
rect 997 15474 1003 15508
rect 1037 15474 1043 15508
rect 997 15435 1043 15474
rect 997 15401 1003 15435
rect 1037 15401 1043 15435
rect 997 15362 1043 15401
rect 997 15328 1003 15362
rect 1037 15328 1043 15362
rect 997 15289 1043 15328
rect 997 15255 1003 15289
rect 1037 15255 1043 15289
rect 997 15216 1043 15255
rect 997 15182 1003 15216
rect 1037 15182 1043 15216
rect 997 15143 1043 15182
rect 997 15109 1003 15143
rect 1037 15109 1043 15143
tri 807 15072 810 15075 sw
tri 994 15072 997 15075 se
rect 997 15072 1043 15109
rect 1233 15508 1279 15520
rect 1233 15474 1239 15508
rect 1273 15474 1279 15508
rect 1233 15435 1279 15474
rect 1233 15401 1239 15435
rect 1273 15401 1279 15435
rect 1233 15362 1279 15401
rect 1233 15328 1239 15362
rect 1273 15328 1279 15362
rect 1233 15289 1279 15328
rect 1233 15255 1239 15289
rect 1273 15255 1279 15289
rect 1233 15216 1279 15255
rect 1233 15182 1239 15216
rect 1273 15182 1279 15216
rect 1233 15143 1279 15182
rect 1233 15109 1239 15143
rect 1273 15109 1279 15143
tri 1043 15072 1046 15075 sw
tri 1230 15072 1233 15075 se
rect 1233 15072 1279 15109
rect 1469 15508 1515 15520
rect 1469 15474 1475 15508
rect 1509 15474 1515 15508
rect 1469 15435 1515 15474
rect 1469 15401 1475 15435
rect 1509 15401 1515 15435
rect 1469 15362 1515 15401
rect 1469 15328 1475 15362
rect 1509 15328 1515 15362
rect 1469 15289 1515 15328
rect 1469 15255 1475 15289
rect 1509 15255 1515 15289
rect 1469 15216 1515 15255
rect 1469 15182 1475 15216
rect 1509 15182 1515 15216
rect 1469 15143 1515 15182
rect 1469 15109 1475 15143
rect 1509 15109 1515 15143
tri 1279 15072 1282 15075 sw
tri 1466 15072 1469 15075 se
rect 1469 15072 1515 15109
rect 1705 15508 1751 15520
rect 1705 15474 1711 15508
rect 1745 15474 1751 15508
rect 1705 15435 1751 15474
rect 1705 15401 1711 15435
rect 1745 15401 1751 15435
rect 1705 15362 1751 15401
rect 1705 15328 1711 15362
rect 1745 15328 1751 15362
rect 1705 15289 1751 15328
rect 1705 15255 1711 15289
rect 1745 15255 1751 15289
rect 1705 15216 1751 15255
rect 1705 15182 1711 15216
rect 1745 15182 1751 15216
rect 1705 15143 1751 15182
rect 1705 15109 1711 15143
rect 1745 15109 1751 15143
tri 1515 15072 1518 15075 sw
tri 1702 15072 1705 15075 se
rect 1705 15072 1751 15109
rect 1941 15508 1987 15520
rect 1941 15474 1947 15508
rect 1981 15474 1987 15508
rect 1941 15435 1987 15474
rect 1941 15401 1947 15435
rect 1981 15401 1987 15435
rect 1941 15362 1987 15401
rect 1941 15328 1947 15362
rect 1981 15328 1987 15362
rect 1941 15289 1987 15328
rect 1941 15255 1947 15289
rect 1981 15255 1987 15289
rect 1941 15216 1987 15255
rect 1941 15182 1947 15216
rect 1981 15182 1987 15216
rect 1941 15143 1987 15182
rect 1941 15109 1947 15143
rect 1981 15109 1987 15143
tri 1751 15072 1754 15075 sw
tri 1938 15072 1941 15075 se
rect 1941 15072 1987 15109
rect 2177 15508 2223 15520
rect 2177 15474 2183 15508
rect 2217 15474 2223 15508
rect 2177 15435 2223 15474
rect 2177 15401 2183 15435
rect 2217 15401 2223 15435
rect 2177 15362 2223 15401
rect 2177 15328 2183 15362
rect 2217 15328 2223 15362
rect 2177 15289 2223 15328
rect 2177 15255 2183 15289
rect 2217 15255 2223 15289
rect 2177 15216 2223 15255
rect 2177 15182 2183 15216
rect 2217 15182 2223 15216
rect 2177 15143 2223 15182
rect 2177 15109 2183 15143
rect 2217 15109 2223 15143
tri 1987 15072 1990 15075 sw
tri 2174 15072 2177 15075 se
rect 2177 15072 2223 15109
rect 2413 15508 2459 15520
rect 2413 15474 2419 15508
rect 2453 15474 2459 15508
rect 2413 15435 2459 15474
rect 2413 15401 2419 15435
rect 2453 15401 2459 15435
rect 2413 15362 2459 15401
rect 2413 15328 2419 15362
rect 2453 15328 2459 15362
rect 2413 15289 2459 15328
rect 2413 15255 2419 15289
rect 2453 15255 2459 15289
rect 2413 15216 2459 15255
rect 2413 15182 2419 15216
rect 2453 15182 2459 15216
rect 2413 15143 2459 15182
rect 2413 15109 2419 15143
rect 2453 15109 2459 15143
tri 2223 15072 2226 15075 sw
tri 2410 15072 2413 15075 se
rect 2413 15072 2459 15109
rect 2649 15508 2695 15520
rect 2649 15474 2655 15508
rect 2689 15474 2695 15508
rect 2649 15435 2695 15474
rect 2649 15401 2655 15435
rect 2689 15401 2695 15435
rect 2649 15362 2695 15401
rect 2649 15328 2655 15362
rect 2689 15328 2695 15362
rect 2649 15289 2695 15328
rect 2649 15255 2655 15289
rect 2689 15255 2695 15289
rect 2649 15216 2695 15255
rect 2649 15182 2655 15216
rect 2689 15182 2695 15216
rect 2649 15143 2695 15182
rect 2649 15109 2655 15143
rect 2689 15109 2695 15143
tri 2459 15072 2462 15075 sw
tri 2646 15072 2649 15075 se
rect 2649 15072 2695 15109
rect 2885 15508 3076 15528
rect 2885 15474 2891 15508
rect 2925 15490 3076 15508
rect 2925 15474 3036 15490
rect 2885 15456 3036 15474
rect 3070 15456 3076 15490
rect 2885 15435 3076 15456
rect 2885 15401 2891 15435
rect 2925 15418 3076 15435
rect 2925 15401 3036 15418
rect 2885 15384 3036 15401
rect 3070 15384 3076 15418
rect 2885 15362 3076 15384
rect 2885 15328 2891 15362
rect 2925 15346 3076 15362
rect 2925 15328 3036 15346
rect 2885 15312 3036 15328
rect 3070 15312 3076 15346
rect 2885 15289 3076 15312
rect 2885 15255 2891 15289
rect 2925 15274 3076 15289
rect 2925 15255 3036 15274
rect 2885 15240 3036 15255
rect 3070 15240 3076 15274
rect 2885 15216 3076 15240
rect 2885 15182 2891 15216
rect 2925 15202 3076 15216
rect 2925 15182 3036 15202
rect 2885 15168 3036 15182
rect 3070 15168 3076 15202
rect 2885 15143 3076 15168
rect 2885 15109 2891 15143
rect 2925 15130 3076 15143
rect 2925 15109 3036 15130
rect 2885 15096 3036 15109
rect 3070 15096 3076 15130
tri 2695 15072 2698 15075 sw
tri 2882 15072 2885 15075 se
rect 2885 15072 3076 15096
rect 380 15070 574 15072
tri 574 15070 576 15072 sw
tri 756 15070 758 15072 se
rect 758 15070 810 15072
tri 810 15070 812 15072 sw
tri 992 15070 994 15072 se
rect 994 15070 1046 15072
tri 1046 15070 1048 15072 sw
tri 1228 15070 1230 15072 se
rect 1230 15070 1282 15072
tri 1282 15070 1284 15072 sw
tri 1464 15070 1466 15072 se
rect 1466 15070 1518 15072
tri 1518 15070 1520 15072 sw
tri 1700 15070 1702 15072 se
rect 1702 15070 1754 15072
tri 1754 15070 1756 15072 sw
tri 1936 15070 1938 15072 se
rect 1938 15070 1990 15072
tri 1990 15070 1992 15072 sw
tri 2172 15070 2174 15072 se
rect 2174 15070 2226 15072
tri 2226 15070 2228 15072 sw
tri 2408 15070 2410 15072 se
rect 2410 15070 2462 15072
tri 2462 15070 2464 15072 sw
tri 2644 15070 2646 15072 se
rect 2646 15070 2698 15072
tri 2698 15070 2700 15072 sw
tri 2880 15070 2882 15072 se
rect 2882 15070 3076 15072
rect 380 15039 531 15070
rect 380 15005 386 15039
rect 420 15036 531 15039
rect 565 15041 576 15070
tri 576 15041 605 15070 sw
tri 727 15041 756 15070 se
rect 756 15041 767 15070
rect 565 15036 767 15041
rect 801 15041 812 15070
tri 812 15041 841 15070 sw
tri 963 15041 992 15070 se
rect 992 15041 1003 15070
rect 801 15036 1003 15041
rect 1037 15041 1048 15070
tri 1048 15041 1077 15070 sw
tri 1199 15041 1228 15070 se
rect 1228 15041 1239 15070
rect 1037 15036 1239 15041
rect 1273 15041 1284 15070
tri 1284 15041 1313 15070 sw
tri 1435 15041 1464 15070 se
rect 1464 15041 1475 15070
rect 1273 15036 1475 15041
rect 1509 15041 1520 15070
tri 1520 15041 1549 15070 sw
tri 1671 15041 1700 15070 se
rect 1700 15041 1711 15070
rect 1509 15036 1711 15041
rect 1745 15041 1756 15070
tri 1756 15041 1785 15070 sw
tri 1907 15041 1936 15070 se
rect 1936 15041 1947 15070
rect 1745 15036 1947 15041
rect 1981 15041 1992 15070
tri 1992 15041 2021 15070 sw
tri 2143 15041 2172 15070 se
rect 2172 15041 2183 15070
rect 1981 15036 2183 15041
rect 2217 15041 2228 15070
tri 2228 15041 2257 15070 sw
tri 2379 15041 2408 15070 se
rect 2408 15041 2419 15070
rect 2217 15036 2419 15041
rect 2453 15041 2464 15070
tri 2464 15041 2493 15070 sw
tri 2615 15041 2644 15070 se
rect 2644 15041 2655 15070
rect 2453 15036 2655 15041
rect 2689 15041 2700 15070
tri 2700 15041 2729 15070 sw
tri 2851 15041 2880 15070 se
rect 2880 15041 2891 15070
rect 2689 15036 2891 15041
rect 2925 15058 3076 15070
rect 2925 15036 3036 15058
rect 420 15024 3036 15036
rect 3070 15024 3076 15058
rect 420 15009 3076 15024
rect 420 15005 697 15009
rect 380 14997 697 15005
rect 380 14967 531 14997
rect 380 14933 386 14967
rect 420 14963 531 14967
rect 565 14963 697 14997
rect 420 14957 697 14963
rect 749 14957 765 15009
rect 817 14957 833 15009
rect 885 14957 901 15009
rect 953 14957 969 15009
rect 1021 14997 1037 15009
rect 1021 14957 1037 14963
rect 1089 14957 1105 15009
rect 1157 14957 1173 15009
rect 1225 14997 1241 15009
rect 1293 14997 2097 15009
rect 1225 14963 1239 14997
rect 1293 14963 1475 14997
rect 1509 14963 1711 14997
rect 1745 14963 1947 14997
rect 1981 14963 2097 14997
rect 1225 14957 1241 14963
rect 1293 14957 2097 14963
rect 2149 14957 2165 15009
rect 2217 14957 2233 15009
rect 2285 14957 2301 15009
rect 2353 14957 2369 15009
rect 2421 14997 2437 15009
rect 2421 14957 2437 14963
rect 2489 14957 2505 15009
rect 2557 14957 2573 15009
rect 2625 14957 2641 15009
rect 2693 14997 3076 15009
rect 2693 14963 2891 14997
rect 2925 14986 3076 14997
rect 2925 14963 3036 14986
rect 2693 14957 3036 14963
rect 420 14952 3036 14957
rect 3070 14952 3076 14986
rect 420 14945 3076 14952
rect 420 14933 697 14945
rect 380 14924 697 14933
rect 380 14895 531 14924
rect 380 14861 386 14895
rect 420 14890 531 14895
rect 565 14893 697 14924
rect 749 14893 765 14945
rect 817 14893 833 14945
rect 885 14893 901 14945
rect 953 14893 969 14945
rect 1021 14924 1037 14945
rect 1089 14893 1105 14945
rect 1157 14893 1173 14945
rect 1225 14924 1241 14945
rect 1293 14924 2097 14945
rect 1225 14893 1239 14924
rect 1293 14893 1475 14924
rect 565 14890 767 14893
rect 801 14890 1003 14893
rect 1037 14890 1239 14893
rect 1273 14890 1475 14893
rect 1509 14890 1711 14924
rect 1745 14890 1947 14924
rect 1981 14893 2097 14924
rect 2149 14893 2165 14945
rect 2217 14893 2233 14945
rect 2285 14893 2301 14945
rect 2353 14893 2369 14945
rect 2421 14924 2437 14945
rect 2489 14893 2505 14945
rect 2557 14893 2573 14945
rect 2625 14893 2641 14945
rect 2693 14924 3076 14945
rect 2693 14893 2891 14924
rect 1981 14890 2183 14893
rect 2217 14890 2419 14893
rect 2453 14890 2655 14893
rect 2689 14890 2891 14893
rect 2925 14914 3076 14924
rect 2925 14890 3036 14914
rect 420 14881 3036 14890
rect 420 14861 697 14881
rect 380 14851 697 14861
rect 380 14823 531 14851
rect 380 14789 386 14823
rect 420 14817 531 14823
rect 565 14829 697 14851
rect 749 14829 765 14881
rect 817 14829 833 14881
rect 885 14829 901 14881
rect 953 14829 969 14881
rect 1021 14851 1037 14881
rect 1089 14829 1105 14881
rect 1157 14829 1173 14881
rect 1225 14851 1241 14881
rect 1293 14851 2097 14881
rect 1225 14829 1239 14851
rect 1293 14829 1475 14851
rect 565 14817 767 14829
rect 801 14817 1003 14829
rect 1037 14817 1239 14829
rect 1273 14817 1475 14829
rect 1509 14817 1711 14851
rect 1745 14817 1947 14851
rect 1981 14829 2097 14851
rect 2149 14829 2165 14881
rect 2217 14829 2233 14881
rect 2285 14829 2301 14881
rect 2353 14829 2369 14881
rect 2421 14851 2437 14881
rect 2489 14829 2505 14881
rect 2557 14829 2573 14881
rect 2625 14829 2641 14881
rect 2693 14880 3036 14881
rect 3070 14880 3076 14914
rect 2693 14851 3076 14880
rect 2693 14829 2891 14851
rect 1981 14817 2183 14829
rect 2217 14817 2419 14829
rect 2453 14817 2655 14829
rect 2689 14817 2891 14829
rect 2925 14842 3076 14851
rect 2925 14817 3036 14842
rect 420 14789 697 14817
rect 380 14778 697 14789
rect 380 14751 531 14778
rect 380 14717 386 14751
rect 420 14744 531 14751
rect 565 14765 697 14778
rect 749 14765 765 14817
rect 817 14765 833 14817
rect 885 14765 901 14817
rect 953 14765 969 14817
rect 1021 14778 1037 14817
rect 1089 14765 1105 14817
rect 1157 14765 1173 14817
rect 1225 14778 1241 14817
rect 1293 14778 2097 14817
rect 1225 14765 1239 14778
rect 1293 14765 1475 14778
rect 565 14753 767 14765
rect 801 14753 1003 14765
rect 1037 14753 1239 14765
rect 1273 14753 1475 14765
rect 565 14744 697 14753
rect 420 14717 697 14744
rect 380 14705 697 14717
rect 380 14679 531 14705
rect 380 14645 386 14679
rect 420 14671 531 14679
rect 565 14701 697 14705
rect 749 14701 765 14753
rect 817 14701 833 14753
rect 885 14701 901 14753
rect 953 14701 969 14753
rect 1021 14705 1037 14744
rect 1089 14701 1105 14753
rect 1157 14701 1173 14753
rect 1225 14744 1239 14753
rect 1293 14744 1475 14753
rect 1509 14744 1711 14778
rect 1745 14744 1947 14778
rect 1981 14765 2097 14778
rect 2149 14765 2165 14817
rect 2217 14765 2233 14817
rect 2285 14765 2301 14817
rect 2353 14765 2369 14817
rect 2421 14778 2437 14817
rect 2489 14765 2505 14817
rect 2557 14765 2573 14817
rect 2625 14765 2641 14817
rect 2693 14808 3036 14817
rect 3070 14808 3076 14842
rect 2693 14778 3076 14808
rect 2693 14765 2891 14778
rect 1981 14753 2183 14765
rect 2217 14753 2419 14765
rect 2453 14753 2655 14765
rect 2689 14753 2891 14765
rect 1981 14744 2097 14753
rect 1225 14705 1241 14744
rect 1293 14705 2097 14744
rect 1225 14701 1239 14705
rect 1293 14701 1475 14705
rect 565 14689 767 14701
rect 801 14689 1003 14701
rect 1037 14689 1239 14701
rect 1273 14689 1475 14701
rect 565 14671 697 14689
rect 420 14645 697 14671
rect 380 14637 697 14645
rect 749 14637 765 14689
rect 817 14637 833 14689
rect 885 14637 901 14689
rect 953 14637 969 14689
rect 1021 14637 1037 14671
rect 1089 14637 1105 14689
rect 1157 14637 1173 14689
rect 1225 14671 1239 14689
rect 1293 14671 1475 14689
rect 1509 14671 1711 14705
rect 1745 14671 1947 14705
rect 1981 14701 2097 14705
rect 2149 14701 2165 14753
rect 2217 14701 2233 14753
rect 2285 14701 2301 14753
rect 2353 14701 2369 14753
rect 2421 14705 2437 14744
rect 2489 14701 2505 14753
rect 2557 14701 2573 14753
rect 2625 14701 2641 14753
rect 2693 14744 2891 14753
rect 2925 14770 3076 14778
rect 2925 14744 3036 14770
rect 2693 14736 3036 14744
rect 3070 14736 3076 14770
rect 2693 14705 3076 14736
rect 2693 14701 2891 14705
rect 1981 14689 2183 14701
rect 2217 14689 2419 14701
rect 2453 14689 2655 14701
rect 2689 14689 2891 14701
rect 1981 14671 2097 14689
rect 1225 14637 1241 14671
rect 1293 14637 2097 14671
rect 2149 14637 2165 14689
rect 2217 14637 2233 14689
rect 2285 14637 2301 14689
rect 2353 14637 2369 14689
rect 2421 14637 2437 14671
rect 2489 14637 2505 14689
rect 2557 14637 2573 14689
rect 2625 14637 2641 14689
rect 2693 14671 2891 14689
rect 2925 14698 3076 14705
rect 2925 14671 3036 14698
rect 2693 14664 3036 14671
rect 3070 14664 3076 14698
rect 2693 14637 3076 14664
rect 380 14632 3076 14637
rect 380 14607 531 14632
rect 380 14573 386 14607
rect 420 14598 531 14607
rect 565 14625 767 14632
rect 801 14625 1003 14632
rect 1037 14625 1239 14632
rect 1273 14625 1475 14632
rect 565 14598 697 14625
rect 420 14573 697 14598
rect 749 14573 765 14625
rect 817 14573 833 14625
rect 885 14573 901 14625
rect 953 14573 969 14625
rect 1021 14573 1037 14598
rect 1089 14573 1105 14625
rect 1157 14573 1173 14625
rect 1225 14598 1239 14625
rect 1293 14598 1475 14625
rect 1509 14598 1711 14632
rect 1745 14598 1947 14632
rect 1981 14625 2183 14632
rect 2217 14625 2419 14632
rect 2453 14625 2655 14632
rect 2689 14625 2891 14632
rect 1981 14598 2097 14625
rect 1225 14573 1241 14598
rect 1293 14573 2097 14598
rect 2149 14573 2165 14625
rect 2217 14573 2233 14625
rect 2285 14573 2301 14625
rect 2353 14573 2369 14625
rect 2421 14573 2437 14598
rect 2489 14573 2505 14625
rect 2557 14573 2573 14625
rect 2625 14573 2641 14625
rect 2693 14598 2891 14625
rect 2925 14626 3076 14632
rect 2925 14598 3036 14626
rect 2693 14592 3036 14598
rect 3070 14592 3076 14626
rect 2693 14573 3076 14592
rect 380 14561 3076 14573
rect 380 14558 697 14561
rect 380 14535 531 14558
rect 380 14501 386 14535
rect 420 14524 531 14535
rect 565 14524 697 14558
rect 420 14509 697 14524
rect 749 14509 765 14561
rect 817 14509 833 14561
rect 885 14509 901 14561
rect 953 14509 969 14561
rect 1021 14558 1037 14561
rect 1021 14509 1037 14524
rect 1089 14509 1105 14561
rect 1157 14509 1173 14561
rect 1225 14558 1241 14561
rect 1293 14558 2097 14561
rect 1225 14524 1239 14558
rect 1293 14524 1475 14558
rect 1509 14524 1711 14558
rect 1745 14524 1947 14558
rect 1981 14524 2097 14558
rect 1225 14509 1241 14524
rect 1293 14509 2097 14524
rect 2149 14509 2165 14561
rect 2217 14509 2233 14561
rect 2285 14509 2301 14561
rect 2353 14509 2369 14561
rect 2421 14558 2437 14561
rect 2421 14509 2437 14524
rect 2489 14509 2505 14561
rect 2557 14509 2573 14561
rect 2625 14509 2641 14561
rect 2693 14558 3076 14561
rect 2693 14524 2891 14558
rect 2925 14554 3076 14558
rect 2925 14524 3036 14554
rect 2693 14520 3036 14524
rect 3070 14520 3076 14554
rect 2693 14509 3076 14520
rect 420 14501 3076 14509
rect 380 14497 3076 14501
rect 380 14484 697 14497
rect 380 14463 531 14484
rect 380 14429 386 14463
rect 420 14450 531 14463
rect 565 14450 697 14484
rect 420 14445 697 14450
rect 749 14445 765 14497
rect 817 14445 833 14497
rect 885 14445 901 14497
rect 953 14445 969 14497
rect 1021 14484 1037 14497
rect 1021 14445 1037 14450
rect 1089 14445 1105 14497
rect 1157 14445 1173 14497
rect 1225 14484 1241 14497
rect 1293 14484 2097 14497
rect 1225 14450 1239 14484
rect 1293 14450 1475 14484
rect 1509 14450 1711 14484
rect 1745 14450 1947 14484
rect 1981 14450 2097 14484
rect 1225 14445 1241 14450
rect 1293 14445 2097 14450
rect 2149 14445 2165 14497
rect 2217 14445 2233 14497
rect 2285 14445 2301 14497
rect 2353 14445 2369 14497
rect 2421 14484 2437 14497
rect 2421 14445 2437 14450
rect 2489 14445 2505 14497
rect 2557 14445 2573 14497
rect 2625 14445 2641 14497
rect 2693 14484 3076 14497
rect 2693 14450 2891 14484
rect 2925 14482 3076 14484
rect 2925 14450 3036 14482
rect 2693 14448 3036 14450
rect 3070 14448 3076 14482
rect 2693 14445 3076 14448
rect 420 14433 3076 14445
rect 420 14429 697 14433
rect 380 14410 697 14429
rect 380 14391 531 14410
rect 380 14357 386 14391
rect 420 14376 531 14391
rect 565 14381 697 14410
rect 749 14381 765 14433
rect 817 14381 833 14433
rect 885 14381 901 14433
rect 953 14381 969 14433
rect 1021 14410 1037 14433
rect 1089 14381 1105 14433
rect 1157 14381 1173 14433
rect 1225 14410 1241 14433
rect 1293 14410 2097 14433
rect 1225 14381 1239 14410
rect 1293 14381 1475 14410
rect 565 14376 767 14381
rect 801 14376 1003 14381
rect 1037 14376 1239 14381
rect 1273 14376 1475 14381
rect 1509 14376 1711 14410
rect 1745 14376 1947 14410
rect 1981 14381 2097 14410
rect 2149 14381 2165 14433
rect 2217 14381 2233 14433
rect 2285 14381 2301 14433
rect 2353 14381 2369 14433
rect 2421 14410 2437 14433
rect 2489 14381 2505 14433
rect 2557 14381 2573 14433
rect 2625 14381 2641 14433
rect 2693 14410 3076 14433
rect 2693 14381 2891 14410
rect 1981 14376 2183 14381
rect 2217 14376 2419 14381
rect 2453 14376 2655 14381
rect 2689 14376 2891 14381
rect 2925 14376 3036 14410
rect 3070 14376 3076 14410
rect 420 14369 3076 14376
rect 420 14357 697 14369
rect 380 14336 697 14357
rect 380 14319 531 14336
rect 380 14285 386 14319
rect 420 14302 531 14319
rect 565 14317 697 14336
rect 749 14317 765 14369
rect 817 14317 833 14369
rect 885 14317 901 14369
rect 953 14317 969 14369
rect 1021 14336 1037 14369
rect 1089 14317 1105 14369
rect 1157 14317 1173 14369
rect 1225 14336 1241 14369
rect 1293 14336 2097 14369
rect 1225 14317 1239 14336
rect 1293 14317 1475 14336
rect 565 14305 767 14317
rect 801 14305 1003 14317
rect 1037 14305 1239 14317
rect 1273 14305 1475 14317
rect 565 14302 697 14305
rect 420 14285 697 14302
rect 380 14262 697 14285
rect 380 14247 531 14262
rect 380 14213 386 14247
rect 420 14228 531 14247
rect 565 14253 697 14262
rect 749 14253 765 14305
rect 817 14253 833 14305
rect 885 14253 901 14305
rect 953 14253 969 14305
rect 1021 14262 1037 14302
rect 1089 14253 1105 14305
rect 1157 14253 1173 14305
rect 1225 14302 1239 14305
rect 1293 14302 1475 14305
rect 1509 14302 1711 14336
rect 1745 14302 1947 14336
rect 1981 14317 2097 14336
rect 2149 14317 2165 14369
rect 2217 14317 2233 14369
rect 2285 14317 2301 14369
rect 2353 14317 2369 14369
rect 2421 14336 2437 14369
rect 2489 14317 2505 14369
rect 2557 14317 2573 14369
rect 2625 14317 2641 14369
rect 2693 14338 3076 14369
rect 2693 14336 3036 14338
rect 2693 14317 2891 14336
rect 1981 14305 2183 14317
rect 2217 14305 2419 14317
rect 2453 14305 2655 14317
rect 2689 14305 2891 14317
rect 1981 14302 2097 14305
rect 1225 14262 1241 14302
rect 1293 14262 2097 14302
rect 1225 14253 1239 14262
rect 1293 14253 1475 14262
rect 565 14241 767 14253
rect 801 14241 1003 14253
rect 1037 14241 1239 14253
rect 1273 14241 1475 14253
rect 565 14228 697 14241
rect 420 14213 697 14228
rect 380 14189 697 14213
rect 749 14189 765 14241
rect 817 14189 833 14241
rect 885 14189 901 14241
rect 953 14189 969 14241
rect 1021 14189 1037 14228
rect 1089 14189 1105 14241
rect 1157 14189 1173 14241
rect 1225 14228 1239 14241
rect 1293 14228 1475 14241
rect 1509 14228 1711 14262
rect 1745 14228 1947 14262
rect 1981 14253 2097 14262
rect 2149 14253 2165 14305
rect 2217 14253 2233 14305
rect 2285 14253 2301 14305
rect 2353 14253 2369 14305
rect 2421 14262 2437 14302
rect 2489 14253 2505 14305
rect 2557 14253 2573 14305
rect 2625 14253 2641 14305
rect 2693 14302 2891 14305
rect 2925 14304 3036 14336
rect 3070 14304 3076 14338
rect 2925 14302 3076 14304
rect 2693 14266 3076 14302
rect 2693 14262 3036 14266
rect 2693 14253 2891 14262
rect 1981 14241 2183 14253
rect 2217 14241 2419 14253
rect 2453 14241 2655 14253
rect 2689 14241 2891 14253
rect 1981 14228 2097 14241
rect 1225 14189 1241 14228
rect 1293 14189 2097 14228
rect 2149 14189 2165 14241
rect 2217 14189 2233 14241
rect 2285 14189 2301 14241
rect 2353 14189 2369 14241
rect 2421 14189 2437 14228
rect 2489 14189 2505 14241
rect 2557 14189 2573 14241
rect 2625 14189 2641 14241
rect 2693 14228 2891 14241
rect 2925 14232 3036 14262
rect 3070 14232 3076 14266
rect 2925 14228 3076 14232
rect 2693 14194 3076 14228
rect 2693 14189 3036 14194
rect 380 14188 3036 14189
rect 380 14175 531 14188
rect 380 14141 386 14175
rect 420 14154 531 14175
rect 565 14177 767 14188
rect 801 14177 1003 14188
rect 1037 14177 1239 14188
rect 1273 14177 1475 14188
rect 565 14154 697 14177
rect 420 14141 697 14154
rect 380 14125 697 14141
rect 749 14125 765 14177
rect 817 14125 833 14177
rect 885 14125 901 14177
rect 953 14125 969 14177
rect 1021 14125 1037 14154
rect 1089 14125 1105 14177
rect 1157 14125 1173 14177
rect 1225 14154 1239 14177
rect 1293 14154 1475 14177
rect 1509 14154 1711 14188
rect 1745 14154 1947 14188
rect 1981 14177 2183 14188
rect 2217 14177 2419 14188
rect 2453 14177 2655 14188
rect 2689 14177 2891 14188
rect 1981 14154 2097 14177
rect 1225 14125 1241 14154
rect 1293 14125 2097 14154
rect 2149 14125 2165 14177
rect 2217 14125 2233 14177
rect 2285 14125 2301 14177
rect 2353 14125 2369 14177
rect 2421 14125 2437 14154
rect 2489 14125 2505 14177
rect 2557 14125 2573 14177
rect 2625 14125 2641 14177
rect 2693 14154 2891 14177
rect 2925 14160 3036 14188
rect 3070 14160 3076 14194
rect 2925 14154 3076 14160
rect 2693 14125 3076 14154
rect 380 14122 3076 14125
rect 380 14114 3036 14122
rect 380 14103 531 14114
rect 380 14069 386 14103
rect 420 14080 531 14103
rect 565 14113 767 14114
rect 801 14113 1003 14114
rect 1037 14113 1239 14114
rect 1273 14113 1475 14114
rect 565 14080 697 14113
rect 420 14069 697 14080
rect 380 14061 697 14069
rect 749 14061 765 14113
rect 817 14061 833 14113
rect 885 14061 901 14113
rect 953 14061 969 14113
rect 1021 14061 1037 14080
rect 1089 14061 1105 14113
rect 1157 14061 1173 14113
rect 1225 14080 1239 14113
rect 1293 14080 1475 14113
rect 1509 14080 1711 14114
rect 1745 14080 1947 14114
rect 1981 14113 2183 14114
rect 2217 14113 2419 14114
rect 2453 14113 2655 14114
rect 2689 14113 2891 14114
rect 1981 14080 2097 14113
rect 1225 14061 1241 14080
rect 1293 14061 2097 14080
rect 2149 14061 2165 14113
rect 2217 14061 2233 14113
rect 2285 14061 2301 14113
rect 2353 14061 2369 14113
rect 2421 14061 2437 14080
rect 2489 14061 2505 14113
rect 2557 14061 2573 14113
rect 2625 14061 2641 14113
rect 2693 14080 2891 14113
rect 2925 14088 3036 14114
rect 3070 14088 3076 14122
rect 2925 14080 3076 14088
rect 2693 14061 3076 14080
rect 380 14050 3076 14061
rect 380 14041 3036 14050
rect 380 14040 604 14041
tri 604 14040 605 14041 nw
tri 727 14040 728 14041 ne
rect 728 14040 840 14041
tri 840 14040 841 14041 nw
tri 963 14040 964 14041 ne
rect 964 14040 1076 14041
tri 1076 14040 1077 14041 nw
tri 1199 14040 1200 14041 ne
rect 1200 14040 1312 14041
tri 1312 14040 1313 14041 nw
tri 1435 14040 1436 14041 ne
rect 1436 14040 1548 14041
tri 1548 14040 1549 14041 nw
tri 1671 14040 1672 14041 ne
rect 1672 14040 1784 14041
tri 1784 14040 1785 14041 nw
tri 1907 14040 1908 14041 ne
rect 1908 14040 2020 14041
tri 2020 14040 2021 14041 nw
tri 2143 14040 2144 14041 ne
rect 2144 14040 2256 14041
tri 2256 14040 2257 14041 nw
tri 2379 14040 2380 14041 ne
rect 2380 14040 2492 14041
tri 2492 14040 2493 14041 nw
tri 2615 14040 2616 14041 ne
rect 2616 14040 2728 14041
tri 2728 14040 2729 14041 nw
tri 2851 14040 2852 14041 ne
rect 2852 14040 3036 14041
rect 380 14031 531 14040
rect 380 13997 386 14031
rect 420 14006 531 14031
rect 565 14006 571 14040
tri 571 14007 604 14040 nw
tri 728 14007 761 14040 ne
rect 420 13997 571 14006
rect 380 13966 571 13997
rect 380 13959 531 13966
rect 380 13925 386 13959
rect 420 13932 531 13959
rect 565 13932 571 13966
rect 420 13925 571 13932
rect 380 13892 571 13925
rect 380 13887 531 13892
rect 380 13853 386 13887
rect 420 13858 531 13887
rect 565 13858 571 13892
rect 420 13853 571 13858
rect 380 13818 571 13853
rect 380 13815 531 13818
rect 380 13781 386 13815
rect 420 13784 531 13815
rect 565 13784 571 13818
rect 420 13781 571 13784
rect 380 13744 571 13781
rect 380 13743 531 13744
rect 380 13709 386 13743
rect 420 13710 531 13743
rect 565 13710 571 13744
rect 420 13709 571 13710
rect 380 13671 571 13709
rect 380 13637 386 13671
rect 420 13670 571 13671
rect 420 13637 531 13670
rect 380 13636 531 13637
rect 565 13636 571 13670
rect 380 13599 571 13636
rect 380 13565 386 13599
rect 420 13596 571 13599
rect 420 13565 531 13596
rect 380 13562 531 13565
rect 565 13562 571 13596
rect 380 13527 571 13562
rect 761 14006 767 14040
rect 801 14006 807 14040
tri 807 14007 840 14040 nw
tri 964 14007 997 14040 ne
rect 761 13966 807 14006
rect 761 13932 767 13966
rect 801 13932 807 13966
rect 761 13892 807 13932
rect 761 13858 767 13892
rect 801 13858 807 13892
rect 761 13818 807 13858
rect 761 13784 767 13818
rect 801 13784 807 13818
rect 761 13744 807 13784
rect 761 13710 767 13744
rect 801 13710 807 13744
rect 761 13670 807 13710
rect 761 13636 767 13670
rect 801 13636 807 13670
rect 761 13596 807 13636
rect 761 13562 767 13596
rect 801 13562 807 13596
rect 761 13550 807 13562
rect 997 14006 1003 14040
rect 1037 14006 1043 14040
tri 1043 14007 1076 14040 nw
tri 1200 14007 1233 14040 ne
rect 997 13966 1043 14006
rect 997 13932 1003 13966
rect 1037 13932 1043 13966
rect 997 13892 1043 13932
rect 997 13858 1003 13892
rect 1037 13858 1043 13892
rect 997 13818 1043 13858
rect 997 13784 1003 13818
rect 1037 13784 1043 13818
rect 997 13744 1043 13784
rect 997 13710 1003 13744
rect 1037 13710 1043 13744
rect 997 13670 1043 13710
rect 997 13636 1003 13670
rect 1037 13636 1043 13670
rect 997 13596 1043 13636
rect 997 13562 1003 13596
rect 1037 13562 1043 13596
rect 997 13550 1043 13562
rect 1233 14006 1239 14040
rect 1273 14006 1279 14040
tri 1279 14007 1312 14040 nw
tri 1436 14007 1469 14040 ne
rect 1233 13966 1279 14006
rect 1233 13932 1239 13966
rect 1273 13932 1279 13966
rect 1233 13892 1279 13932
rect 1233 13858 1239 13892
rect 1273 13858 1279 13892
rect 1233 13818 1279 13858
rect 1233 13784 1239 13818
rect 1273 13784 1279 13818
rect 1233 13744 1279 13784
rect 1233 13710 1239 13744
rect 1273 13710 1279 13744
rect 1233 13670 1279 13710
rect 1233 13636 1239 13670
rect 1273 13636 1279 13670
rect 1233 13596 1279 13636
rect 1233 13562 1239 13596
rect 1273 13562 1279 13596
rect 1233 13550 1279 13562
rect 1469 14006 1475 14040
rect 1509 14006 1515 14040
tri 1515 14007 1548 14040 nw
tri 1672 14007 1705 14040 ne
rect 1469 13966 1515 14006
rect 1469 13932 1475 13966
rect 1509 13932 1515 13966
rect 1469 13892 1515 13932
rect 1469 13858 1475 13892
rect 1509 13858 1515 13892
rect 1469 13818 1515 13858
rect 1469 13784 1475 13818
rect 1509 13784 1515 13818
rect 1469 13744 1515 13784
rect 1469 13710 1475 13744
rect 1509 13710 1515 13744
rect 1469 13670 1515 13710
rect 1469 13636 1475 13670
rect 1509 13636 1515 13670
rect 1469 13596 1515 13636
rect 1469 13562 1475 13596
rect 1509 13562 1515 13596
rect 1469 13550 1515 13562
rect 1705 14006 1711 14040
rect 1745 14006 1751 14040
tri 1751 14007 1784 14040 nw
tri 1908 14007 1941 14040 ne
rect 1705 13966 1751 14006
rect 1705 13932 1711 13966
rect 1745 13932 1751 13966
rect 1705 13892 1751 13932
rect 1705 13858 1711 13892
rect 1745 13858 1751 13892
rect 1705 13818 1751 13858
rect 1705 13784 1711 13818
rect 1745 13784 1751 13818
rect 1705 13744 1751 13784
rect 1705 13710 1711 13744
rect 1745 13710 1751 13744
rect 1705 13670 1751 13710
rect 1705 13636 1711 13670
rect 1745 13636 1751 13670
rect 1705 13596 1751 13636
rect 1705 13562 1711 13596
rect 1745 13562 1751 13596
rect 1705 13550 1751 13562
rect 1941 14006 1947 14040
rect 1981 14006 1987 14040
tri 1987 14007 2020 14040 nw
tri 2144 14007 2177 14040 ne
rect 1941 13966 1987 14006
rect 1941 13932 1947 13966
rect 1981 13932 1987 13966
rect 1941 13892 1987 13932
rect 1941 13858 1947 13892
rect 1981 13858 1987 13892
rect 1941 13818 1987 13858
rect 1941 13784 1947 13818
rect 1981 13784 1987 13818
rect 1941 13744 1987 13784
rect 1941 13710 1947 13744
rect 1981 13710 1987 13744
rect 1941 13670 1987 13710
rect 1941 13636 1947 13670
rect 1981 13636 1987 13670
rect 1941 13596 1987 13636
rect 1941 13562 1947 13596
rect 1981 13562 1987 13596
rect 1941 13550 1987 13562
rect 2177 14006 2183 14040
rect 2217 14006 2223 14040
tri 2223 14007 2256 14040 nw
tri 2380 14007 2413 14040 ne
rect 2177 13966 2223 14006
rect 2177 13932 2183 13966
rect 2217 13932 2223 13966
rect 2177 13892 2223 13932
rect 2177 13858 2183 13892
rect 2217 13858 2223 13892
rect 2177 13818 2223 13858
rect 2177 13784 2183 13818
rect 2217 13784 2223 13818
rect 2177 13744 2223 13784
rect 2177 13710 2183 13744
rect 2217 13710 2223 13744
rect 2177 13670 2223 13710
rect 2177 13636 2183 13670
rect 2217 13636 2223 13670
rect 2177 13596 2223 13636
rect 2177 13562 2183 13596
rect 2217 13562 2223 13596
rect 2177 13550 2223 13562
rect 2413 14006 2419 14040
rect 2453 14006 2459 14040
tri 2459 14007 2492 14040 nw
tri 2616 14007 2649 14040 ne
rect 2413 13966 2459 14006
rect 2413 13932 2419 13966
rect 2453 13932 2459 13966
rect 2413 13892 2459 13932
rect 2413 13858 2419 13892
rect 2453 13858 2459 13892
rect 2413 13818 2459 13858
rect 2413 13784 2419 13818
rect 2453 13784 2459 13818
rect 2413 13744 2459 13784
rect 2413 13710 2419 13744
rect 2453 13710 2459 13744
rect 2413 13670 2459 13710
rect 2413 13636 2419 13670
rect 2453 13636 2459 13670
rect 2413 13596 2459 13636
rect 2413 13562 2419 13596
rect 2453 13562 2459 13596
rect 2413 13550 2459 13562
rect 2649 14006 2655 14040
rect 2689 14006 2695 14040
tri 2695 14007 2728 14040 nw
tri 2852 14007 2885 14040 ne
rect 2649 13966 2695 14006
rect 2649 13932 2655 13966
rect 2689 13932 2695 13966
rect 2649 13892 2695 13932
rect 2649 13858 2655 13892
rect 2689 13858 2695 13892
rect 2649 13818 2695 13858
rect 2649 13784 2655 13818
rect 2689 13784 2695 13818
rect 2649 13744 2695 13784
rect 2649 13710 2655 13744
rect 2689 13710 2695 13744
rect 2649 13670 2695 13710
rect 2649 13636 2655 13670
rect 2689 13636 2695 13670
rect 2649 13596 2695 13636
rect 2649 13562 2655 13596
rect 2689 13562 2695 13596
rect 2649 13550 2695 13562
rect 2885 14006 2891 14040
rect 2925 14016 3036 14040
rect 3070 14016 3076 14050
rect 2925 14006 3076 14016
rect 2885 13978 3076 14006
rect 2885 13966 3036 13978
rect 2885 13932 2891 13966
rect 2925 13944 3036 13966
rect 3070 13944 3076 13978
rect 2925 13932 3076 13944
rect 2885 13906 3076 13932
rect 2885 13892 3036 13906
rect 2885 13858 2891 13892
rect 2925 13872 3036 13892
rect 3070 13872 3076 13906
rect 2925 13858 3076 13872
rect 2885 13834 3076 13858
rect 2885 13818 3036 13834
rect 2885 13784 2891 13818
rect 2925 13800 3036 13818
rect 3070 13800 3076 13834
rect 2925 13784 3076 13800
rect 2885 13762 3076 13784
rect 2885 13744 3036 13762
rect 2885 13710 2891 13744
rect 2925 13728 3036 13744
rect 3070 13728 3076 13762
rect 2925 13710 3076 13728
rect 2885 13690 3076 13710
rect 2885 13670 3036 13690
rect 2885 13636 2891 13670
rect 2925 13656 3036 13670
rect 3070 13656 3076 13690
rect 2925 13636 3076 13656
rect 2885 13618 3076 13636
rect 2885 13596 3036 13618
rect 2885 13562 2891 13596
rect 2925 13584 3036 13596
rect 3070 13584 3076 13618
rect 2925 13562 3076 13584
rect 380 13493 386 13527
rect 420 13493 571 13527
rect 2885 13546 3076 13562
rect 2885 13512 3036 13546
rect 3070 13512 3076 13546
rect 380 13455 571 13493
rect 380 13421 386 13455
rect 420 13421 571 13455
rect 613 13494 1501 13503
rect 1553 13494 1569 13503
rect 1621 13494 1636 13503
rect 1688 13494 1703 13503
rect 1755 13494 1770 13503
rect 1822 13494 1837 13503
rect 1889 13494 2830 13503
rect 613 13460 625 13494
rect 659 13460 700 13494
rect 734 13460 775 13494
rect 809 13460 850 13494
rect 884 13460 925 13494
rect 959 13460 1000 13494
rect 1034 13460 1075 13494
rect 1109 13460 1150 13494
rect 1184 13460 1225 13494
rect 1259 13460 1300 13494
rect 1334 13460 1375 13494
rect 1409 13460 1450 13494
rect 1484 13460 1501 13494
rect 1559 13460 1569 13494
rect 1634 13460 1636 13494
rect 1889 13460 1896 13494
rect 1930 13460 1970 13494
rect 2004 13460 2044 13494
rect 2078 13460 2118 13494
rect 2152 13460 2192 13494
rect 2226 13460 2266 13494
rect 2300 13460 2340 13494
rect 2374 13460 2414 13494
rect 2448 13460 2488 13494
rect 2522 13460 2562 13494
rect 2596 13460 2636 13494
rect 2670 13460 2710 13494
rect 2744 13460 2784 13494
rect 2818 13460 2830 13494
rect 613 13451 1501 13460
rect 1553 13451 1569 13460
rect 1621 13451 1636 13460
rect 1688 13451 1703 13460
rect 1755 13451 1770 13460
rect 1822 13451 1837 13460
rect 1889 13451 2830 13460
rect 2885 13474 3076 13512
rect 380 13392 571 13421
rect 2885 13440 3036 13474
rect 3070 13440 3076 13474
rect 380 13383 531 13392
rect 380 13349 386 13383
rect 420 13358 531 13383
rect 565 13358 571 13392
rect 420 13349 571 13358
rect 380 13319 571 13349
rect 380 13311 531 13319
rect 380 13277 386 13311
rect 420 13285 531 13311
rect 565 13285 571 13319
rect 420 13277 571 13285
rect 380 13246 571 13277
rect 380 13239 531 13246
rect 380 13205 386 13239
rect 420 13212 531 13239
rect 565 13212 571 13246
rect 420 13205 571 13212
rect 380 13173 571 13205
rect 380 13167 531 13173
rect 380 13133 386 13167
rect 420 13139 531 13167
rect 565 13139 571 13173
rect 420 13133 571 13139
rect 380 13100 571 13133
rect 380 13095 531 13100
rect 380 13061 386 13095
rect 420 13066 531 13095
rect 565 13066 571 13100
rect 420 13061 571 13066
rect 380 13027 571 13061
rect 380 13023 531 13027
rect 380 12989 386 13023
rect 420 12993 531 13023
rect 565 12993 571 13027
rect 420 12989 571 12993
rect 380 12954 571 12989
rect 761 13392 807 13404
rect 761 13358 767 13392
rect 801 13358 807 13392
rect 761 13319 807 13358
rect 761 13285 767 13319
rect 801 13285 807 13319
rect 761 13246 807 13285
rect 761 13212 767 13246
rect 801 13212 807 13246
rect 761 13173 807 13212
rect 761 13139 767 13173
rect 801 13139 807 13173
rect 761 13100 807 13139
rect 761 13066 767 13100
rect 801 13066 807 13100
rect 761 13027 807 13066
rect 761 12993 767 13027
rect 801 12993 807 13027
tri 571 12954 581 12964 sw
tri 751 12954 761 12964 se
rect 761 12954 807 12993
rect 997 13392 1043 13404
rect 997 13358 1003 13392
rect 1037 13358 1043 13392
rect 997 13319 1043 13358
rect 997 13285 1003 13319
rect 1037 13285 1043 13319
rect 997 13246 1043 13285
rect 997 13212 1003 13246
rect 1037 13212 1043 13246
rect 997 13173 1043 13212
rect 997 13139 1003 13173
rect 1037 13139 1043 13173
rect 997 13100 1043 13139
rect 997 13066 1003 13100
rect 1037 13066 1043 13100
rect 997 13027 1043 13066
rect 997 12993 1003 13027
rect 1037 12993 1043 13027
tri 807 12954 817 12964 sw
tri 987 12954 997 12964 se
rect 997 12954 1043 12993
rect 1233 13392 1279 13404
rect 1233 13358 1239 13392
rect 1273 13358 1279 13392
rect 1233 13319 1279 13358
rect 1233 13285 1239 13319
rect 1273 13285 1279 13319
rect 1233 13246 1279 13285
rect 1233 13212 1239 13246
rect 1273 13212 1279 13246
rect 1233 13173 1279 13212
rect 1233 13139 1239 13173
rect 1273 13139 1279 13173
rect 1233 13100 1279 13139
rect 1233 13066 1239 13100
rect 1273 13066 1279 13100
rect 1233 13027 1279 13066
rect 1233 12993 1239 13027
rect 1273 12993 1279 13027
tri 1043 12954 1053 12964 sw
tri 1223 12954 1233 12964 se
rect 1233 12954 1279 12993
rect 1469 13392 1515 13404
rect 1469 13358 1475 13392
rect 1509 13358 1515 13392
rect 1469 13319 1515 13358
rect 1469 13285 1475 13319
rect 1509 13285 1515 13319
rect 1469 13246 1515 13285
rect 1469 13212 1475 13246
rect 1509 13212 1515 13246
rect 1469 13173 1515 13212
rect 1469 13139 1475 13173
rect 1509 13139 1515 13173
rect 1469 13100 1515 13139
rect 1469 13066 1475 13100
rect 1509 13066 1515 13100
rect 1469 13027 1515 13066
rect 1469 12993 1475 13027
rect 1509 12993 1515 13027
tri 1279 12954 1289 12964 sw
tri 1459 12954 1469 12964 se
rect 1469 12954 1515 12993
rect 1705 13392 1751 13404
rect 1705 13358 1711 13392
rect 1745 13358 1751 13392
rect 1705 13319 1751 13358
rect 1705 13285 1711 13319
rect 1745 13285 1751 13319
rect 1705 13246 1751 13285
rect 1705 13212 1711 13246
rect 1745 13212 1751 13246
rect 1705 13173 1751 13212
rect 1705 13139 1711 13173
rect 1745 13139 1751 13173
rect 1705 13100 1751 13139
rect 1705 13066 1711 13100
rect 1745 13066 1751 13100
rect 1705 13027 1751 13066
rect 1705 12993 1711 13027
rect 1745 12993 1751 13027
tri 1515 12954 1525 12964 sw
tri 1695 12954 1705 12964 se
rect 1705 12954 1751 12993
rect 1941 13392 1987 13404
rect 1941 13358 1947 13392
rect 1981 13358 1987 13392
rect 1941 13319 1987 13358
rect 1941 13285 1947 13319
rect 1981 13285 1987 13319
rect 1941 13246 1987 13285
rect 1941 13212 1947 13246
rect 1981 13212 1987 13246
rect 1941 13173 1987 13212
rect 1941 13139 1947 13173
rect 1981 13139 1987 13173
rect 1941 13100 1987 13139
rect 1941 13066 1947 13100
rect 1981 13066 1987 13100
rect 1941 13027 1987 13066
rect 1941 12993 1947 13027
rect 1981 12993 1987 13027
tri 1751 12954 1761 12964 sw
tri 1931 12954 1941 12964 se
rect 1941 12954 1987 12993
rect 2177 13392 2223 13404
rect 2177 13358 2183 13392
rect 2217 13358 2223 13392
rect 2177 13319 2223 13358
rect 2177 13285 2183 13319
rect 2217 13285 2223 13319
rect 2177 13246 2223 13285
rect 2177 13212 2183 13246
rect 2217 13212 2223 13246
rect 2177 13173 2223 13212
rect 2177 13139 2183 13173
rect 2217 13139 2223 13173
rect 2177 13100 2223 13139
rect 2177 13066 2183 13100
rect 2217 13066 2223 13100
rect 2177 13027 2223 13066
rect 2177 12993 2183 13027
rect 2217 12993 2223 13027
tri 1987 12954 1997 12964 sw
tri 2167 12954 2177 12964 se
rect 2177 12954 2223 12993
rect 2413 13392 2459 13404
rect 2413 13358 2419 13392
rect 2453 13358 2459 13392
rect 2413 13319 2459 13358
rect 2413 13285 2419 13319
rect 2453 13285 2459 13319
rect 2413 13246 2459 13285
rect 2413 13212 2419 13246
rect 2453 13212 2459 13246
rect 2413 13173 2459 13212
rect 2413 13139 2419 13173
rect 2453 13139 2459 13173
rect 2413 13100 2459 13139
rect 2413 13066 2419 13100
rect 2453 13066 2459 13100
rect 2413 13027 2459 13066
rect 2413 12993 2419 13027
rect 2453 12993 2459 13027
tri 2223 12954 2233 12964 sw
tri 2403 12954 2413 12964 se
rect 2413 12954 2459 12993
rect 2649 13392 2695 13404
rect 2649 13358 2655 13392
rect 2689 13358 2695 13392
rect 2649 13319 2695 13358
rect 2649 13285 2655 13319
rect 2689 13285 2695 13319
rect 2649 13246 2695 13285
rect 2649 13212 2655 13246
rect 2689 13212 2695 13246
rect 2649 13173 2695 13212
rect 2649 13139 2655 13173
rect 2689 13139 2695 13173
rect 2649 13100 2695 13139
rect 2649 13066 2655 13100
rect 2689 13066 2695 13100
rect 2649 13027 2695 13066
rect 2649 12993 2655 13027
rect 2689 12993 2695 13027
tri 2459 12954 2469 12964 sw
tri 2639 12954 2649 12964 se
rect 2649 12954 2695 12993
rect 2885 13402 3076 13440
rect 2885 13392 3036 13402
rect 2885 13358 2891 13392
rect 2925 13368 3036 13392
rect 3070 13368 3076 13402
rect 2925 13358 3076 13368
rect 2885 13330 3076 13358
rect 2885 13319 3036 13330
rect 2885 13285 2891 13319
rect 2925 13296 3036 13319
rect 3070 13296 3076 13330
rect 2925 13285 3076 13296
rect 2885 13258 3076 13285
rect 2885 13246 3036 13258
rect 2885 13212 2891 13246
rect 2925 13224 3036 13246
rect 3070 13224 3076 13258
rect 2925 13212 3076 13224
rect 2885 13186 3076 13212
rect 2885 13173 3036 13186
rect 2885 13139 2891 13173
rect 2925 13152 3036 13173
rect 3070 13152 3076 13186
rect 2925 13139 3076 13152
rect 2885 13114 3076 13139
rect 2885 13100 3036 13114
rect 2885 13066 2891 13100
rect 2925 13080 3036 13100
rect 3070 13080 3076 13114
rect 2925 13066 3076 13080
rect 2885 13042 3076 13066
rect 2885 13027 3036 13042
rect 2885 12993 2891 13027
rect 2925 13008 3036 13027
rect 3070 13008 3076 13042
rect 2925 12993 3076 13008
rect 2885 12970 3076 12993
tri 2695 12954 2705 12964 sw
tri 2875 12954 2885 12964 se
rect 2885 12954 3036 12970
rect 380 12951 531 12954
rect 380 12917 386 12951
rect 420 12920 531 12951
rect 565 12930 581 12954
tri 581 12930 605 12954 sw
tri 727 12930 751 12954 se
rect 751 12930 767 12954
rect 565 12920 767 12930
rect 801 12930 817 12954
tri 817 12930 841 12954 sw
tri 963 12930 987 12954 se
rect 987 12930 1003 12954
rect 801 12920 1003 12930
rect 1037 12930 1053 12954
tri 1053 12930 1077 12954 sw
tri 1199 12930 1223 12954 se
rect 1223 12930 1239 12954
rect 1037 12920 1239 12930
rect 1273 12930 1289 12954
tri 1289 12930 1313 12954 sw
tri 1435 12930 1459 12954 se
rect 1459 12930 1475 12954
rect 1273 12920 1475 12930
rect 1509 12930 1525 12954
tri 1525 12930 1549 12954 sw
tri 1671 12930 1695 12954 se
rect 1695 12930 1711 12954
rect 1509 12920 1711 12930
rect 1745 12930 1761 12954
tri 1761 12930 1785 12954 sw
tri 1907 12930 1931 12954 se
rect 1931 12930 1947 12954
rect 1745 12920 1947 12930
rect 1981 12930 1997 12954
tri 1997 12930 2021 12954 sw
tri 2143 12930 2167 12954 se
rect 2167 12930 2183 12954
rect 1981 12920 2183 12930
rect 2217 12930 2233 12954
tri 2233 12930 2257 12954 sw
tri 2379 12930 2403 12954 se
rect 2403 12930 2419 12954
rect 2217 12920 2419 12930
rect 2453 12930 2469 12954
tri 2469 12930 2493 12954 sw
tri 2615 12930 2639 12954 se
rect 2639 12930 2655 12954
rect 2453 12920 2655 12930
rect 2689 12930 2705 12954
tri 2705 12930 2729 12954 sw
tri 2851 12930 2875 12954 se
rect 2875 12930 2891 12954
rect 2689 12920 2891 12930
rect 2925 12936 3036 12954
rect 3070 12936 3076 12970
rect 2925 12920 3076 12936
rect 420 12917 3076 12920
rect 380 12907 3076 12917
rect 380 12881 697 12907
rect 380 12879 531 12881
rect 380 12845 386 12879
rect 420 12847 531 12879
rect 565 12855 697 12881
rect 749 12855 765 12907
rect 817 12855 833 12907
rect 885 12855 901 12907
rect 953 12855 969 12907
rect 1021 12881 1037 12907
rect 1089 12855 1105 12907
rect 1157 12855 1173 12907
rect 1225 12881 1241 12907
rect 1293 12881 2097 12907
rect 1225 12855 1239 12881
rect 1293 12855 1475 12881
rect 565 12847 767 12855
rect 801 12847 1003 12855
rect 1037 12847 1239 12855
rect 1273 12847 1475 12855
rect 1509 12847 1711 12881
rect 1745 12847 1947 12881
rect 1981 12855 2097 12881
rect 2149 12855 2165 12907
rect 2217 12855 2233 12907
rect 2285 12855 2301 12907
rect 2353 12855 2369 12907
rect 2421 12881 2437 12907
rect 2489 12855 2505 12907
rect 2557 12855 2573 12907
rect 2625 12855 2641 12907
rect 2693 12898 3076 12907
rect 2693 12881 3036 12898
rect 2693 12855 2891 12881
rect 1981 12847 2183 12855
rect 2217 12847 2419 12855
rect 2453 12847 2655 12855
rect 2689 12847 2891 12855
rect 2925 12864 3036 12881
rect 3070 12864 3076 12898
rect 2925 12847 3076 12864
rect 420 12845 3076 12847
rect 380 12843 3076 12845
rect 380 12808 697 12843
rect 380 12807 531 12808
rect 380 12773 386 12807
rect 420 12774 531 12807
rect 565 12791 697 12808
rect 749 12791 765 12843
rect 817 12791 833 12843
rect 885 12791 901 12843
rect 953 12791 969 12843
rect 1021 12808 1037 12843
rect 1089 12791 1105 12843
rect 1157 12791 1173 12843
rect 1225 12808 1241 12843
rect 1293 12808 2097 12843
rect 1225 12791 1239 12808
rect 1293 12791 1475 12808
rect 565 12779 767 12791
rect 801 12779 1003 12791
rect 1037 12779 1239 12791
rect 1273 12779 1475 12791
rect 565 12774 697 12779
rect 420 12773 697 12774
rect 380 12735 697 12773
rect 380 12701 386 12735
rect 420 12701 531 12735
rect 565 12727 697 12735
rect 749 12727 765 12779
rect 817 12727 833 12779
rect 885 12727 901 12779
rect 953 12727 969 12779
rect 1021 12735 1037 12774
rect 1089 12727 1105 12779
rect 1157 12727 1173 12779
rect 1225 12774 1239 12779
rect 1293 12774 1475 12779
rect 1509 12774 1711 12808
rect 1745 12774 1947 12808
rect 1981 12791 2097 12808
rect 2149 12791 2165 12843
rect 2217 12791 2233 12843
rect 2285 12791 2301 12843
rect 2353 12791 2369 12843
rect 2421 12808 2437 12843
rect 2489 12791 2505 12843
rect 2557 12791 2573 12843
rect 2625 12791 2641 12843
rect 2693 12826 3076 12843
rect 2693 12808 3036 12826
rect 2693 12791 2891 12808
rect 1981 12779 2183 12791
rect 2217 12779 2419 12791
rect 2453 12779 2655 12791
rect 2689 12779 2891 12791
rect 1981 12774 2097 12779
rect 1225 12735 1241 12774
rect 1293 12735 2097 12774
rect 1225 12727 1239 12735
rect 1293 12727 1475 12735
rect 565 12715 767 12727
rect 801 12715 1003 12727
rect 1037 12715 1239 12727
rect 1273 12715 1475 12727
rect 565 12701 697 12715
rect 380 12663 697 12701
rect 749 12663 765 12715
rect 817 12663 833 12715
rect 885 12663 901 12715
rect 953 12663 969 12715
rect 1021 12663 1037 12701
rect 1089 12663 1105 12715
rect 1157 12663 1173 12715
rect 1225 12701 1239 12715
rect 1293 12701 1475 12715
rect 1509 12701 1711 12735
rect 1745 12701 1947 12735
rect 1981 12727 2097 12735
rect 2149 12727 2165 12779
rect 2217 12727 2233 12779
rect 2285 12727 2301 12779
rect 2353 12727 2369 12779
rect 2421 12735 2437 12774
rect 2489 12727 2505 12779
rect 2557 12727 2573 12779
rect 2625 12727 2641 12779
rect 2693 12774 2891 12779
rect 2925 12792 3036 12808
rect 3070 12792 3076 12826
rect 2925 12774 3076 12792
rect 2693 12754 3076 12774
rect 2693 12735 3036 12754
rect 2693 12727 2891 12735
rect 1981 12715 2183 12727
rect 2217 12715 2419 12727
rect 2453 12715 2655 12727
rect 2689 12715 2891 12727
rect 1981 12701 2097 12715
rect 1225 12663 1241 12701
rect 1293 12663 2097 12701
rect 2149 12663 2165 12715
rect 2217 12663 2233 12715
rect 2285 12663 2301 12715
rect 2353 12663 2369 12715
rect 2421 12663 2437 12701
rect 2489 12663 2505 12715
rect 2557 12663 2573 12715
rect 2625 12663 2641 12715
rect 2693 12701 2891 12715
rect 2925 12720 3036 12735
rect 3070 12720 3076 12754
rect 2925 12701 3076 12720
rect 2693 12682 3076 12701
rect 2693 12663 3036 12682
rect 380 12629 386 12663
rect 420 12662 3036 12663
rect 420 12629 531 12662
rect 380 12628 531 12629
rect 565 12651 767 12662
rect 801 12651 1003 12662
rect 1037 12651 1239 12662
rect 1273 12651 1475 12662
rect 565 12628 697 12651
rect 380 12599 697 12628
rect 749 12599 765 12651
rect 817 12599 833 12651
rect 885 12599 901 12651
rect 953 12599 969 12651
rect 1021 12599 1037 12628
rect 1089 12599 1105 12651
rect 1157 12599 1173 12651
rect 1225 12628 1239 12651
rect 1293 12628 1475 12651
rect 1509 12628 1711 12662
rect 1745 12628 1947 12662
rect 1981 12651 2183 12662
rect 2217 12651 2419 12662
rect 2453 12651 2655 12662
rect 2689 12651 2891 12662
rect 1981 12628 2097 12651
rect 1225 12599 1241 12628
rect 1293 12599 2097 12628
rect 2149 12599 2165 12651
rect 2217 12599 2233 12651
rect 2285 12599 2301 12651
rect 2353 12599 2369 12651
rect 2421 12599 2437 12628
rect 2489 12599 2505 12651
rect 2557 12599 2573 12651
rect 2625 12599 2641 12651
rect 2693 12628 2891 12651
rect 2925 12648 3036 12662
rect 3070 12648 3076 12682
rect 2925 12628 3076 12648
rect 2693 12610 3076 12628
rect 2693 12599 3036 12610
rect 380 12591 3036 12599
rect 380 12557 386 12591
rect 420 12589 3036 12591
rect 420 12557 531 12589
rect 380 12555 531 12557
rect 565 12587 767 12589
rect 801 12587 1003 12589
rect 1037 12587 1239 12589
rect 1273 12587 1475 12589
rect 565 12555 697 12587
rect 380 12535 697 12555
rect 749 12535 765 12587
rect 817 12535 833 12587
rect 885 12535 901 12587
rect 953 12535 969 12587
rect 1021 12535 1037 12555
rect 1089 12535 1105 12587
rect 1157 12535 1173 12587
rect 1225 12555 1239 12587
rect 1293 12555 1475 12587
rect 1509 12555 1711 12589
rect 1745 12555 1947 12589
rect 1981 12587 2183 12589
rect 2217 12587 2419 12589
rect 2453 12587 2655 12589
rect 2689 12587 2891 12589
rect 1981 12555 2097 12587
rect 1225 12535 1241 12555
rect 1293 12535 2097 12555
rect 2149 12535 2165 12587
rect 2217 12535 2233 12587
rect 2285 12535 2301 12587
rect 2353 12535 2369 12587
rect 2421 12535 2437 12555
rect 2489 12535 2505 12587
rect 2557 12535 2573 12587
rect 2625 12535 2641 12587
rect 2693 12555 2891 12587
rect 2925 12576 3036 12589
rect 3070 12576 3076 12610
rect 2925 12555 3076 12576
rect 2693 12538 3076 12555
rect 2693 12535 3036 12538
rect 380 12523 3036 12535
rect 380 12519 697 12523
rect 380 12485 386 12519
rect 420 12516 697 12519
rect 420 12485 531 12516
rect 380 12482 531 12485
rect 565 12482 697 12516
rect 380 12471 697 12482
rect 749 12471 765 12523
rect 817 12471 833 12523
rect 885 12471 901 12523
rect 953 12471 969 12523
rect 1021 12516 1037 12523
rect 1021 12471 1037 12482
rect 1089 12471 1105 12523
rect 1157 12471 1173 12523
rect 1225 12516 1241 12523
rect 1293 12516 2097 12523
rect 1225 12482 1239 12516
rect 1293 12482 1475 12516
rect 1509 12482 1711 12516
rect 1745 12482 1947 12516
rect 1981 12482 2097 12516
rect 1225 12471 1241 12482
rect 1293 12471 2097 12482
rect 2149 12471 2165 12523
rect 2217 12471 2233 12523
rect 2285 12471 2301 12523
rect 2353 12471 2369 12523
rect 2421 12516 2437 12523
rect 2421 12471 2437 12482
rect 2489 12471 2505 12523
rect 2557 12471 2573 12523
rect 2625 12471 2641 12523
rect 2693 12516 3036 12523
rect 2693 12482 2891 12516
rect 2925 12504 3036 12516
rect 3070 12504 3076 12538
rect 2925 12482 3076 12504
rect 2693 12471 3076 12482
rect 380 12466 3076 12471
rect 380 12459 3036 12466
rect 380 12447 697 12459
rect 380 12413 386 12447
rect 420 12442 697 12447
rect 420 12413 531 12442
rect 380 12408 531 12413
rect 565 12408 697 12442
rect 380 12407 697 12408
rect 749 12407 765 12459
rect 817 12407 833 12459
rect 885 12407 901 12459
rect 953 12407 969 12459
rect 1021 12442 1037 12459
rect 1021 12407 1037 12408
rect 1089 12407 1105 12459
rect 1157 12407 1173 12459
rect 1225 12442 1241 12459
rect 1293 12442 2097 12459
rect 1225 12408 1239 12442
rect 1293 12408 1475 12442
rect 1509 12408 1711 12442
rect 1745 12408 1947 12442
rect 1981 12408 2097 12442
rect 1225 12407 1241 12408
rect 1293 12407 2097 12408
rect 2149 12407 2165 12459
rect 2217 12407 2233 12459
rect 2285 12407 2301 12459
rect 2353 12407 2369 12459
rect 2421 12442 2437 12459
rect 2421 12407 2437 12408
rect 2489 12407 2505 12459
rect 2557 12407 2573 12459
rect 2625 12407 2641 12459
rect 2693 12442 3036 12459
rect 2693 12408 2891 12442
rect 2925 12432 3036 12442
rect 3070 12432 3076 12466
rect 2925 12408 3076 12432
rect 2693 12407 3076 12408
rect 380 12395 3076 12407
rect 380 12375 697 12395
rect 380 12341 386 12375
rect 420 12368 697 12375
rect 420 12341 531 12368
rect 380 12334 531 12341
rect 565 12343 697 12368
rect 749 12343 765 12395
rect 817 12343 833 12395
rect 885 12343 901 12395
rect 953 12343 969 12395
rect 1021 12368 1037 12395
rect 1089 12343 1105 12395
rect 1157 12343 1173 12395
rect 1225 12368 1241 12395
rect 1293 12368 2097 12395
rect 1225 12343 1239 12368
rect 1293 12343 1475 12368
rect 565 12334 767 12343
rect 801 12334 1003 12343
rect 1037 12334 1239 12343
rect 1273 12334 1475 12343
rect 1509 12334 1711 12368
rect 1745 12334 1947 12368
rect 1981 12343 2097 12368
rect 2149 12343 2165 12395
rect 2217 12343 2233 12395
rect 2285 12343 2301 12395
rect 2353 12343 2369 12395
rect 2421 12368 2437 12395
rect 2489 12343 2505 12395
rect 2557 12343 2573 12395
rect 2625 12343 2641 12395
rect 2693 12394 3076 12395
rect 2693 12368 3036 12394
rect 2693 12343 2891 12368
rect 1981 12334 2183 12343
rect 2217 12334 2419 12343
rect 2453 12334 2655 12343
rect 2689 12334 2891 12343
rect 2925 12360 3036 12368
rect 3070 12360 3076 12394
rect 2925 12334 3076 12360
rect 380 12331 3076 12334
rect 380 12303 697 12331
rect 380 12269 386 12303
rect 420 12294 697 12303
rect 420 12269 531 12294
rect 380 12260 531 12269
rect 565 12279 697 12294
rect 749 12279 765 12331
rect 817 12279 833 12331
rect 885 12279 901 12331
rect 953 12279 969 12331
rect 1021 12294 1037 12331
rect 1089 12279 1105 12331
rect 1157 12279 1173 12331
rect 1225 12294 1241 12331
rect 1293 12294 2097 12331
rect 1225 12279 1239 12294
rect 1293 12279 1475 12294
rect 565 12267 767 12279
rect 801 12267 1003 12279
rect 1037 12267 1239 12279
rect 1273 12267 1475 12279
rect 565 12260 697 12267
rect 380 12231 697 12260
rect 380 12197 386 12231
rect 420 12220 697 12231
rect 420 12197 531 12220
rect 380 12186 531 12197
rect 565 12215 697 12220
rect 749 12215 765 12267
rect 817 12215 833 12267
rect 885 12215 901 12267
rect 953 12215 969 12267
rect 1021 12220 1037 12260
rect 1089 12215 1105 12267
rect 1157 12215 1173 12267
rect 1225 12260 1239 12267
rect 1293 12260 1475 12267
rect 1509 12260 1711 12294
rect 1745 12260 1947 12294
rect 1981 12279 2097 12294
rect 2149 12279 2165 12331
rect 2217 12279 2233 12331
rect 2285 12279 2301 12331
rect 2353 12279 2369 12331
rect 2421 12294 2437 12331
rect 2489 12279 2505 12331
rect 2557 12279 2573 12331
rect 2625 12279 2641 12331
rect 2693 12322 3076 12331
rect 2693 12294 3036 12322
rect 2693 12279 2891 12294
rect 1981 12267 2183 12279
rect 2217 12267 2419 12279
rect 2453 12267 2655 12279
rect 2689 12267 2891 12279
rect 1981 12260 2097 12267
rect 1225 12220 1241 12260
rect 1293 12220 2097 12260
rect 1225 12215 1239 12220
rect 1293 12215 1475 12220
rect 565 12203 767 12215
rect 801 12203 1003 12215
rect 1037 12203 1239 12215
rect 1273 12203 1475 12215
rect 565 12186 697 12203
rect 380 12159 697 12186
rect 380 12125 386 12159
rect 420 12151 697 12159
rect 749 12151 765 12203
rect 817 12151 833 12203
rect 885 12151 901 12203
rect 953 12151 969 12203
rect 1021 12151 1037 12186
rect 1089 12151 1105 12203
rect 1157 12151 1173 12203
rect 1225 12186 1239 12203
rect 1293 12186 1475 12203
rect 1509 12186 1711 12220
rect 1745 12186 1947 12220
rect 1981 12215 2097 12220
rect 2149 12215 2165 12267
rect 2217 12215 2233 12267
rect 2285 12215 2301 12267
rect 2353 12215 2369 12267
rect 2421 12220 2437 12260
rect 2489 12215 2505 12267
rect 2557 12215 2573 12267
rect 2625 12215 2641 12267
rect 2693 12260 2891 12267
rect 2925 12288 3036 12294
rect 3070 12288 3076 12322
rect 2925 12260 3076 12288
rect 2693 12250 3076 12260
rect 2693 12220 3036 12250
rect 2693 12215 2891 12220
rect 1981 12203 2183 12215
rect 2217 12203 2419 12215
rect 2453 12203 2655 12215
rect 2689 12203 2891 12215
rect 1981 12186 2097 12203
rect 1225 12151 1241 12186
rect 1293 12151 2097 12186
rect 2149 12151 2165 12203
rect 2217 12151 2233 12203
rect 2285 12151 2301 12203
rect 2353 12151 2369 12203
rect 2421 12151 2437 12186
rect 2489 12151 2505 12203
rect 2557 12151 2573 12203
rect 2625 12151 2641 12203
rect 2693 12186 2891 12203
rect 2925 12216 3036 12220
rect 3070 12216 3076 12250
rect 2925 12186 3076 12216
rect 2693 12178 3076 12186
rect 2693 12151 3036 12178
rect 420 12146 3036 12151
rect 420 12125 531 12146
rect 380 12112 531 12125
rect 565 12139 767 12146
rect 801 12139 1003 12146
rect 1037 12139 1239 12146
rect 1273 12139 1475 12146
rect 565 12112 697 12139
rect 380 12087 697 12112
rect 749 12087 765 12139
rect 817 12087 833 12139
rect 885 12087 901 12139
rect 953 12087 969 12139
rect 1021 12087 1037 12112
rect 1089 12087 1105 12139
rect 1157 12087 1173 12139
rect 1225 12112 1239 12139
rect 1293 12112 1475 12139
rect 1509 12112 1711 12146
rect 1745 12112 1947 12146
rect 1981 12139 2183 12146
rect 2217 12139 2419 12146
rect 2453 12139 2655 12146
rect 2689 12139 2891 12146
rect 1981 12112 2097 12139
rect 1225 12087 1241 12112
rect 1293 12087 2097 12112
rect 2149 12087 2165 12139
rect 2217 12087 2233 12139
rect 2285 12087 2301 12139
rect 2353 12087 2369 12139
rect 2421 12087 2437 12112
rect 2489 12087 2505 12139
rect 2557 12087 2573 12139
rect 2625 12087 2641 12139
rect 2693 12112 2891 12139
rect 2925 12144 3036 12146
rect 3070 12144 3076 12178
rect 2925 12112 3076 12144
rect 2693 12106 3076 12112
rect 2693 12087 3036 12106
rect 380 12053 386 12087
rect 420 12075 3036 12087
rect 420 12072 697 12075
rect 420 12053 531 12072
rect 380 12038 531 12053
rect 565 12038 697 12072
rect 380 12023 697 12038
rect 749 12023 765 12075
rect 817 12023 833 12075
rect 885 12023 901 12075
rect 953 12023 969 12075
rect 1021 12072 1037 12075
rect 1021 12023 1037 12038
rect 1089 12023 1105 12075
rect 1157 12023 1173 12075
rect 1225 12072 1241 12075
rect 1293 12072 2097 12075
rect 1225 12038 1239 12072
rect 1293 12038 1475 12072
rect 1509 12038 1711 12072
rect 1745 12038 1947 12072
rect 1981 12038 2097 12072
rect 1225 12023 1241 12038
rect 1293 12023 2097 12038
rect 2149 12023 2165 12075
rect 2217 12023 2233 12075
rect 2285 12023 2301 12075
rect 2353 12023 2369 12075
rect 2421 12072 2437 12075
rect 2421 12023 2437 12038
rect 2489 12023 2505 12075
rect 2557 12023 2573 12075
rect 2625 12023 2641 12075
rect 2693 12072 3036 12075
rect 3070 12072 3076 12106
rect 2693 12038 2891 12072
rect 2925 12038 3076 12072
rect 2693 12034 3076 12038
rect 2693 12023 3036 12034
rect 380 12015 3036 12023
rect 380 11981 386 12015
rect 420 12011 3036 12015
rect 420 11998 697 12011
rect 420 11981 531 11998
rect 380 11964 531 11981
rect 565 11964 697 11998
rect 380 11959 697 11964
rect 749 11959 765 12011
rect 817 11959 833 12011
rect 885 11959 901 12011
rect 953 11959 969 12011
rect 1021 11998 1037 12011
rect 1021 11959 1037 11964
rect 1089 11959 1105 12011
rect 1157 11959 1173 12011
rect 1225 11998 1241 12011
rect 1293 11998 2097 12011
rect 1225 11964 1239 11998
rect 1293 11964 1475 11998
rect 1509 11964 1711 11998
rect 1745 11964 1947 11998
rect 1981 11964 2097 11998
rect 1225 11959 1241 11964
rect 1293 11959 2097 11964
rect 2149 11959 2165 12011
rect 2217 11959 2233 12011
rect 2285 11959 2301 12011
rect 2353 11959 2369 12011
rect 2421 11998 2437 12011
rect 2421 11959 2437 11964
rect 2489 11959 2505 12011
rect 2557 11959 2573 12011
rect 2625 11959 2641 12011
rect 2693 12000 3036 12011
rect 3070 12000 3076 12034
rect 2693 11998 3076 12000
rect 2693 11964 2891 11998
rect 2925 11964 3076 11998
rect 2693 11962 3076 11964
rect 2693 11959 3036 11962
rect 380 11943 3036 11959
rect 380 11909 386 11943
rect 420 11930 3036 11943
rect 420 11928 603 11930
tri 603 11928 605 11930 nw
tri 727 11928 729 11930 ne
rect 729 11928 839 11930
tri 839 11928 841 11930 nw
tri 963 11928 965 11930 ne
rect 965 11928 1075 11930
tri 1075 11928 1077 11930 nw
tri 1199 11928 1201 11930 ne
rect 1201 11928 1311 11930
tri 1311 11928 1313 11930 nw
tri 1435 11928 1437 11930 ne
rect 1437 11928 1547 11930
tri 1547 11928 1549 11930 nw
tri 1671 11928 1673 11930 ne
rect 1673 11928 1783 11930
tri 1783 11928 1785 11930 nw
tri 1907 11928 1909 11930 ne
rect 1909 11928 2019 11930
tri 2019 11928 2021 11930 nw
tri 2143 11928 2145 11930 ne
rect 2145 11928 2255 11930
tri 2255 11928 2257 11930 nw
tri 2379 11928 2381 11930 ne
rect 2381 11928 2491 11930
tri 2491 11928 2493 11930 nw
tri 2615 11928 2617 11930 ne
rect 2617 11928 2727 11930
tri 2727 11928 2729 11930 nw
tri 2851 11928 2853 11930 ne
rect 2853 11928 3036 11930
rect 3070 11928 3076 11962
rect 420 11924 599 11928
tri 599 11924 603 11928 nw
tri 729 11924 733 11928 ne
rect 733 11924 835 11928
tri 835 11924 839 11928 nw
tri 965 11924 969 11928 ne
rect 969 11924 1071 11928
tri 1071 11924 1075 11928 nw
tri 1201 11924 1205 11928 ne
rect 1205 11924 1307 11928
tri 1307 11924 1311 11928 nw
tri 1437 11924 1441 11928 ne
rect 1441 11924 1543 11928
tri 1543 11924 1547 11928 nw
tri 1673 11924 1677 11928 ne
rect 1677 11924 1779 11928
tri 1779 11924 1783 11928 nw
tri 1909 11924 1913 11928 ne
rect 1913 11924 2015 11928
tri 2015 11924 2019 11928 nw
tri 2145 11924 2149 11928 ne
rect 2149 11924 2251 11928
tri 2251 11924 2255 11928 nw
tri 2381 11924 2385 11928 ne
rect 2385 11924 2487 11928
tri 2487 11924 2491 11928 nw
tri 2617 11924 2621 11928 ne
rect 2621 11924 2723 11928
tri 2723 11924 2727 11928 nw
tri 2853 11924 2857 11928 ne
rect 2857 11924 3076 11928
rect 420 11909 531 11924
rect 380 11890 531 11909
rect 565 11890 571 11924
tri 571 11896 599 11924 nw
tri 733 11896 761 11924 ne
rect 380 11871 571 11890
rect 380 11837 386 11871
rect 420 11850 571 11871
rect 420 11837 531 11850
rect 380 11816 531 11837
rect 565 11816 571 11850
rect 380 11799 571 11816
rect 380 11765 386 11799
rect 420 11776 571 11799
rect 420 11765 531 11776
rect 380 11742 531 11765
rect 565 11742 571 11776
rect 380 11727 571 11742
rect 380 11693 386 11727
rect 420 11702 571 11727
rect 420 11693 531 11702
rect 380 11668 531 11693
rect 565 11668 571 11702
rect 380 11655 571 11668
rect 380 11621 386 11655
rect 420 11628 571 11655
rect 420 11621 531 11628
rect 380 11594 531 11621
rect 565 11594 571 11628
rect 380 11583 571 11594
rect 380 11549 386 11583
rect 420 11554 571 11583
rect 420 11549 531 11554
rect 380 11520 531 11549
rect 565 11520 571 11554
rect 380 11511 571 11520
rect 380 11477 386 11511
rect 420 11480 571 11511
rect 420 11477 531 11480
rect 380 11446 531 11477
rect 565 11446 571 11480
rect 380 11439 571 11446
rect 380 11405 386 11439
rect 420 11405 571 11439
rect 761 11890 767 11924
rect 801 11890 807 11924
tri 807 11896 835 11924 nw
tri 969 11896 997 11924 ne
rect 761 11850 807 11890
rect 761 11816 767 11850
rect 801 11816 807 11850
rect 761 11776 807 11816
rect 761 11742 767 11776
rect 801 11742 807 11776
rect 761 11702 807 11742
rect 761 11668 767 11702
rect 801 11668 807 11702
rect 761 11628 807 11668
rect 761 11594 767 11628
rect 801 11594 807 11628
rect 761 11554 807 11594
rect 761 11520 767 11554
rect 801 11520 807 11554
rect 761 11480 807 11520
rect 761 11446 767 11480
rect 801 11446 807 11480
rect 761 11434 807 11446
rect 997 11890 1003 11924
rect 1037 11890 1043 11924
tri 1043 11896 1071 11924 nw
tri 1205 11896 1233 11924 ne
rect 997 11850 1043 11890
rect 997 11816 1003 11850
rect 1037 11816 1043 11850
rect 997 11776 1043 11816
rect 997 11742 1003 11776
rect 1037 11742 1043 11776
rect 997 11702 1043 11742
rect 997 11668 1003 11702
rect 1037 11668 1043 11702
rect 997 11628 1043 11668
rect 997 11594 1003 11628
rect 1037 11594 1043 11628
rect 997 11554 1043 11594
rect 997 11520 1003 11554
rect 1037 11520 1043 11554
rect 997 11480 1043 11520
rect 997 11446 1003 11480
rect 1037 11446 1043 11480
rect 997 11434 1043 11446
rect 1233 11890 1239 11924
rect 1273 11890 1279 11924
tri 1279 11896 1307 11924 nw
tri 1441 11896 1469 11924 ne
rect 1233 11850 1279 11890
rect 1233 11816 1239 11850
rect 1273 11816 1279 11850
rect 1233 11776 1279 11816
rect 1233 11742 1239 11776
rect 1273 11742 1279 11776
rect 1233 11702 1279 11742
rect 1233 11668 1239 11702
rect 1273 11668 1279 11702
rect 1233 11628 1279 11668
rect 1233 11594 1239 11628
rect 1273 11594 1279 11628
rect 1233 11554 1279 11594
rect 1233 11520 1239 11554
rect 1273 11520 1279 11554
rect 1233 11480 1279 11520
rect 1233 11446 1239 11480
rect 1273 11446 1279 11480
rect 1233 11434 1279 11446
rect 1469 11890 1475 11924
rect 1509 11890 1515 11924
tri 1515 11896 1543 11924 nw
tri 1677 11896 1705 11924 ne
rect 1469 11850 1515 11890
rect 1469 11816 1475 11850
rect 1509 11816 1515 11850
rect 1469 11776 1515 11816
rect 1469 11742 1475 11776
rect 1509 11742 1515 11776
rect 1469 11702 1515 11742
rect 1469 11668 1475 11702
rect 1509 11668 1515 11702
rect 1469 11628 1515 11668
rect 1469 11594 1475 11628
rect 1509 11594 1515 11628
rect 1469 11554 1515 11594
rect 1469 11520 1475 11554
rect 1509 11520 1515 11554
rect 1469 11480 1515 11520
rect 1469 11446 1475 11480
rect 1509 11446 1515 11480
rect 1469 11434 1515 11446
rect 1705 11890 1711 11924
rect 1745 11890 1751 11924
tri 1751 11896 1779 11924 nw
tri 1913 11896 1941 11924 ne
rect 1705 11850 1751 11890
rect 1705 11816 1711 11850
rect 1745 11816 1751 11850
rect 1705 11776 1751 11816
rect 1705 11742 1711 11776
rect 1745 11742 1751 11776
rect 1705 11702 1751 11742
rect 1705 11668 1711 11702
rect 1745 11668 1751 11702
rect 1705 11628 1751 11668
rect 1705 11594 1711 11628
rect 1745 11594 1751 11628
rect 1705 11554 1751 11594
rect 1705 11520 1711 11554
rect 1745 11520 1751 11554
rect 1705 11480 1751 11520
rect 1705 11446 1711 11480
rect 1745 11446 1751 11480
rect 1705 11434 1751 11446
rect 1941 11890 1947 11924
rect 1981 11890 1987 11924
tri 1987 11896 2015 11924 nw
tri 2149 11896 2177 11924 ne
rect 1941 11850 1987 11890
rect 1941 11816 1947 11850
rect 1981 11816 1987 11850
rect 1941 11776 1987 11816
rect 1941 11742 1947 11776
rect 1981 11742 1987 11776
rect 1941 11702 1987 11742
rect 1941 11668 1947 11702
rect 1981 11668 1987 11702
rect 1941 11628 1987 11668
rect 1941 11594 1947 11628
rect 1981 11594 1987 11628
rect 1941 11554 1987 11594
rect 1941 11520 1947 11554
rect 1981 11520 1987 11554
rect 1941 11480 1987 11520
rect 1941 11446 1947 11480
rect 1981 11446 1987 11480
rect 1941 11434 1987 11446
rect 2177 11890 2183 11924
rect 2217 11890 2223 11924
tri 2223 11896 2251 11924 nw
tri 2385 11896 2413 11924 ne
rect 2177 11850 2223 11890
rect 2177 11816 2183 11850
rect 2217 11816 2223 11850
rect 2177 11776 2223 11816
rect 2177 11742 2183 11776
rect 2217 11742 2223 11776
rect 2177 11702 2223 11742
rect 2177 11668 2183 11702
rect 2217 11668 2223 11702
rect 2177 11628 2223 11668
rect 2177 11594 2183 11628
rect 2217 11594 2223 11628
rect 2177 11554 2223 11594
rect 2177 11520 2183 11554
rect 2217 11520 2223 11554
rect 2177 11480 2223 11520
rect 2177 11446 2183 11480
rect 2217 11446 2223 11480
rect 2177 11434 2223 11446
rect 2413 11890 2419 11924
rect 2453 11890 2459 11924
tri 2459 11896 2487 11924 nw
tri 2621 11896 2649 11924 ne
rect 2413 11850 2459 11890
rect 2413 11816 2419 11850
rect 2453 11816 2459 11850
rect 2413 11776 2459 11816
rect 2413 11742 2419 11776
rect 2453 11742 2459 11776
rect 2413 11702 2459 11742
rect 2413 11668 2419 11702
rect 2453 11668 2459 11702
rect 2413 11628 2459 11668
rect 2413 11594 2419 11628
rect 2453 11594 2459 11628
rect 2413 11554 2459 11594
rect 2413 11520 2419 11554
rect 2453 11520 2459 11554
rect 2413 11480 2459 11520
rect 2413 11446 2419 11480
rect 2453 11446 2459 11480
rect 2413 11434 2459 11446
rect 2649 11890 2655 11924
rect 2689 11890 2695 11924
tri 2695 11896 2723 11924 nw
tri 2857 11896 2885 11924 ne
rect 2649 11850 2695 11890
rect 2649 11816 2655 11850
rect 2689 11816 2695 11850
rect 2649 11776 2695 11816
rect 2649 11742 2655 11776
rect 2689 11742 2695 11776
rect 2649 11702 2695 11742
rect 2649 11668 2655 11702
rect 2689 11668 2695 11702
rect 2649 11628 2695 11668
rect 2649 11594 2655 11628
rect 2689 11594 2695 11628
rect 2649 11554 2695 11594
rect 2649 11520 2655 11554
rect 2689 11520 2695 11554
rect 2649 11480 2695 11520
rect 2649 11446 2655 11480
rect 2689 11446 2695 11480
rect 2649 11434 2695 11446
rect 2885 11890 2891 11924
rect 2925 11890 3076 11924
rect 2885 11856 3036 11890
rect 3070 11856 3076 11890
rect 2885 11850 3076 11856
rect 2885 11816 2891 11850
rect 2925 11818 3076 11850
rect 2925 11816 3036 11818
rect 2885 11784 3036 11816
rect 3070 11784 3076 11818
rect 2885 11776 3076 11784
rect 2885 11742 2891 11776
rect 2925 11746 3076 11776
rect 2925 11742 3036 11746
rect 2885 11712 3036 11742
rect 3070 11712 3076 11746
rect 2885 11702 3076 11712
rect 2885 11668 2891 11702
rect 2925 11674 3076 11702
rect 2925 11668 3036 11674
rect 2885 11640 3036 11668
rect 3070 11640 3076 11674
rect 2885 11628 3076 11640
rect 2885 11594 2891 11628
rect 2925 11602 3076 11628
rect 2925 11594 3036 11602
rect 2885 11568 3036 11594
rect 3070 11568 3076 11602
rect 2885 11554 3076 11568
rect 2885 11520 2891 11554
rect 2925 11530 3076 11554
rect 2925 11520 3036 11530
rect 2885 11496 3036 11520
rect 3070 11496 3076 11530
rect 2885 11480 3076 11496
rect 2885 11446 2891 11480
rect 2925 11458 3076 11480
rect 2925 11446 3036 11458
rect 380 11367 571 11405
rect 2885 11424 3036 11446
rect 3070 11424 3076 11458
rect 2885 11386 3076 11424
rect 380 11333 386 11367
rect 420 11333 571 11367
rect 380 11295 571 11333
rect 613 11364 1501 11373
rect 1553 11364 1569 11373
rect 1621 11364 1636 11373
rect 1688 11364 1703 11373
rect 1755 11364 1770 11373
rect 1822 11364 1837 11373
rect 1889 11364 2830 11373
rect 613 11330 625 11364
rect 659 11330 700 11364
rect 734 11330 775 11364
rect 809 11330 850 11364
rect 884 11330 925 11364
rect 959 11330 1000 11364
rect 1034 11330 1075 11364
rect 1109 11330 1150 11364
rect 1184 11330 1225 11364
rect 1259 11330 1300 11364
rect 1334 11330 1375 11364
rect 1409 11330 1450 11364
rect 1484 11330 1501 11364
rect 1559 11330 1569 11364
rect 1634 11330 1636 11364
rect 1889 11330 1896 11364
rect 1930 11330 1970 11364
rect 2004 11330 2044 11364
rect 2078 11330 2118 11364
rect 2152 11330 2192 11364
rect 2226 11330 2266 11364
rect 2300 11330 2340 11364
rect 2374 11330 2414 11364
rect 2448 11330 2488 11364
rect 2522 11330 2562 11364
rect 2596 11330 2636 11364
rect 2670 11330 2710 11364
rect 2744 11330 2784 11364
rect 2818 11330 2830 11364
rect 613 11321 1501 11330
rect 1553 11321 1569 11330
rect 1621 11321 1636 11330
rect 1688 11321 1703 11330
rect 1755 11321 1770 11330
rect 1822 11321 1837 11330
rect 1889 11321 2830 11330
rect 2885 11352 3036 11386
rect 3070 11352 3076 11386
rect 380 11261 386 11295
rect 420 11261 571 11295
rect 380 11248 571 11261
rect 2885 11314 3076 11352
rect 2885 11280 3036 11314
rect 3070 11280 3076 11314
rect 380 11223 531 11248
rect 380 11189 386 11223
rect 420 11214 531 11223
rect 565 11214 571 11248
rect 420 11189 571 11214
rect 380 11175 571 11189
rect 380 11151 531 11175
rect 380 11117 386 11151
rect 420 11141 531 11151
rect 565 11141 571 11175
rect 420 11117 571 11141
rect 380 11102 571 11117
rect 380 11079 531 11102
rect 380 11045 386 11079
rect 420 11068 531 11079
rect 565 11068 571 11102
rect 420 11045 571 11068
rect 380 11029 571 11045
rect 380 11007 531 11029
rect 380 10973 386 11007
rect 420 10995 531 11007
rect 565 10995 571 11029
rect 420 10973 571 10995
rect 380 10956 571 10973
rect 380 10935 531 10956
rect 380 10901 386 10935
rect 420 10922 531 10935
rect 565 10922 571 10956
rect 420 10901 571 10922
rect 380 10883 571 10901
rect 380 10863 531 10883
rect 380 10829 386 10863
rect 420 10849 531 10863
rect 565 10849 571 10883
rect 761 11248 807 11260
rect 761 11214 767 11248
rect 801 11214 807 11248
rect 761 11175 807 11214
rect 761 11141 767 11175
rect 801 11141 807 11175
rect 761 11102 807 11141
rect 761 11068 767 11102
rect 801 11068 807 11102
rect 761 11029 807 11068
rect 761 10995 767 11029
rect 801 10995 807 11029
rect 761 10956 807 10995
rect 761 10922 767 10956
rect 801 10922 807 10956
rect 761 10883 807 10922
tri 571 10849 591 10869 sw
tri 741 10849 761 10869 se
rect 761 10849 767 10883
rect 801 10849 807 10883
rect 997 11248 1043 11260
rect 997 11214 1003 11248
rect 1037 11214 1043 11248
rect 997 11175 1043 11214
rect 997 11141 1003 11175
rect 1037 11141 1043 11175
rect 997 11102 1043 11141
rect 997 11068 1003 11102
rect 1037 11068 1043 11102
rect 997 11029 1043 11068
rect 997 10995 1003 11029
rect 1037 10995 1043 11029
rect 997 10956 1043 10995
rect 997 10922 1003 10956
rect 1037 10922 1043 10956
rect 997 10883 1043 10922
tri 807 10849 827 10869 sw
tri 977 10849 997 10869 se
rect 997 10849 1003 10883
rect 1037 10849 1043 10883
rect 1233 11248 1279 11260
rect 1233 11214 1239 11248
rect 1273 11214 1279 11248
rect 1233 11175 1279 11214
rect 1233 11141 1239 11175
rect 1273 11141 1279 11175
rect 1233 11102 1279 11141
rect 1233 11068 1239 11102
rect 1273 11068 1279 11102
rect 1233 11029 1279 11068
rect 1233 10995 1239 11029
rect 1273 10995 1279 11029
rect 1233 10956 1279 10995
rect 1233 10922 1239 10956
rect 1273 10922 1279 10956
rect 1233 10883 1279 10922
tri 1043 10849 1063 10869 sw
tri 1213 10849 1233 10869 se
rect 1233 10849 1239 10883
rect 1273 10849 1279 10883
rect 1469 11248 1515 11260
rect 1469 11214 1475 11248
rect 1509 11214 1515 11248
rect 1469 11175 1515 11214
rect 1469 11141 1475 11175
rect 1509 11141 1515 11175
rect 1469 11102 1515 11141
rect 1469 11068 1475 11102
rect 1509 11068 1515 11102
rect 1469 11029 1515 11068
rect 1469 10995 1475 11029
rect 1509 10995 1515 11029
rect 1469 10956 1515 10995
rect 1469 10922 1475 10956
rect 1509 10922 1515 10956
rect 1469 10883 1515 10922
tri 1279 10849 1299 10869 sw
tri 1449 10849 1469 10869 se
rect 1469 10849 1475 10883
rect 1509 10849 1515 10883
rect 1705 11248 1751 11260
rect 1705 11214 1711 11248
rect 1745 11214 1751 11248
rect 1705 11175 1751 11214
rect 1705 11141 1711 11175
rect 1745 11141 1751 11175
rect 1705 11102 1751 11141
rect 1705 11068 1711 11102
rect 1745 11068 1751 11102
rect 1705 11029 1751 11068
rect 1705 10995 1711 11029
rect 1745 10995 1751 11029
rect 1705 10956 1751 10995
rect 1705 10922 1711 10956
rect 1745 10922 1751 10956
rect 1705 10883 1751 10922
tri 1515 10849 1535 10869 sw
tri 1685 10849 1705 10869 se
rect 1705 10849 1711 10883
rect 1745 10849 1751 10883
rect 1941 11248 1987 11260
rect 1941 11214 1947 11248
rect 1981 11214 1987 11248
rect 1941 11175 1987 11214
rect 1941 11141 1947 11175
rect 1981 11141 1987 11175
rect 1941 11102 1987 11141
rect 1941 11068 1947 11102
rect 1981 11068 1987 11102
rect 1941 11029 1987 11068
rect 1941 10995 1947 11029
rect 1981 10995 1987 11029
rect 1941 10956 1987 10995
rect 1941 10922 1947 10956
rect 1981 10922 1987 10956
rect 1941 10883 1987 10922
tri 1751 10849 1771 10869 sw
tri 1921 10849 1941 10869 se
rect 1941 10849 1947 10883
rect 1981 10849 1987 10883
rect 2177 11248 2223 11260
rect 2177 11214 2183 11248
rect 2217 11214 2223 11248
rect 2177 11175 2223 11214
rect 2177 11141 2183 11175
rect 2217 11141 2223 11175
rect 2177 11102 2223 11141
rect 2177 11068 2183 11102
rect 2217 11068 2223 11102
rect 2177 11029 2223 11068
rect 2177 10995 2183 11029
rect 2217 10995 2223 11029
rect 2177 10956 2223 10995
rect 2177 10922 2183 10956
rect 2217 10922 2223 10956
rect 2177 10883 2223 10922
tri 1987 10849 2007 10869 sw
tri 2157 10849 2177 10869 se
rect 2177 10849 2183 10883
rect 2217 10849 2223 10883
rect 2413 11248 2459 11260
rect 2413 11214 2419 11248
rect 2453 11214 2459 11248
rect 2413 11175 2459 11214
rect 2413 11141 2419 11175
rect 2453 11141 2459 11175
rect 2413 11102 2459 11141
rect 2413 11068 2419 11102
rect 2453 11068 2459 11102
rect 2413 11029 2459 11068
rect 2413 10995 2419 11029
rect 2453 10995 2459 11029
rect 2413 10956 2459 10995
rect 2413 10922 2419 10956
rect 2453 10922 2459 10956
rect 2413 10883 2459 10922
tri 2223 10849 2243 10869 sw
tri 2393 10849 2413 10869 se
rect 2413 10849 2419 10883
rect 2453 10849 2459 10883
rect 2649 11248 2695 11260
rect 2649 11214 2655 11248
rect 2689 11214 2695 11248
rect 2649 11175 2695 11214
rect 2649 11141 2655 11175
rect 2689 11141 2695 11175
rect 2649 11102 2695 11141
rect 2649 11068 2655 11102
rect 2689 11068 2695 11102
rect 2649 11029 2695 11068
rect 2649 10995 2655 11029
rect 2689 10995 2695 11029
rect 2649 10956 2695 10995
rect 2649 10922 2655 10956
rect 2689 10922 2695 10956
rect 2649 10883 2695 10922
tri 2459 10849 2479 10869 sw
tri 2629 10849 2649 10869 se
rect 2649 10849 2655 10883
rect 2689 10849 2695 10883
rect 2885 11248 3076 11280
rect 2885 11214 2891 11248
rect 2925 11242 3076 11248
rect 2925 11214 3036 11242
rect 2885 11208 3036 11214
rect 3070 11208 3076 11242
rect 2885 11175 3076 11208
rect 2885 11141 2891 11175
rect 2925 11170 3076 11175
rect 2925 11141 3036 11170
rect 2885 11136 3036 11141
rect 3070 11136 3076 11170
rect 2885 11102 3076 11136
rect 2885 11068 2891 11102
rect 2925 11098 3076 11102
rect 2925 11068 3036 11098
rect 2885 11064 3036 11068
rect 3070 11064 3076 11098
rect 2885 11029 3076 11064
rect 2885 10995 2891 11029
rect 2925 11026 3076 11029
rect 2925 10995 3036 11026
rect 2885 10992 3036 10995
rect 3070 10992 3076 11026
rect 2885 10956 3076 10992
rect 2885 10922 2891 10956
rect 2925 10954 3076 10956
rect 2925 10922 3036 10954
rect 2885 10920 3036 10922
rect 3070 10920 3076 10954
rect 2885 10883 3076 10920
tri 2695 10849 2715 10869 sw
tri 2865 10849 2885 10869 se
rect 2885 10849 2891 10883
rect 2925 10882 3076 10883
rect 2925 10849 3036 10882
rect 420 10848 591 10849
tri 591 10848 592 10849 sw
tri 740 10848 741 10849 se
rect 741 10848 827 10849
tri 827 10848 828 10849 sw
tri 976 10848 977 10849 se
rect 977 10848 1063 10849
tri 1063 10848 1064 10849 sw
tri 1212 10848 1213 10849 se
rect 1213 10848 1299 10849
tri 1299 10848 1300 10849 sw
tri 1448 10848 1449 10849 se
rect 1449 10848 1535 10849
tri 1535 10848 1536 10849 sw
tri 1684 10848 1685 10849 se
rect 1685 10848 1771 10849
tri 1771 10848 1772 10849 sw
tri 1920 10848 1921 10849 se
rect 1921 10848 2007 10849
tri 2007 10848 2008 10849 sw
tri 2156 10848 2157 10849 se
rect 2157 10848 2243 10849
tri 2243 10848 2244 10849 sw
tri 2392 10848 2393 10849 se
rect 2393 10848 2479 10849
tri 2479 10848 2480 10849 sw
tri 2628 10848 2629 10849 se
rect 2629 10848 2715 10849
tri 2715 10848 2716 10849 sw
tri 2864 10848 2865 10849 se
rect 2865 10848 3036 10849
rect 3070 10848 3076 10882
rect 420 10835 592 10848
tri 592 10835 605 10848 sw
tri 727 10835 740 10848 se
rect 740 10835 828 10848
tri 828 10835 841 10848 sw
tri 963 10835 976 10848 se
rect 976 10835 1064 10848
tri 1064 10835 1077 10848 sw
tri 1199 10835 1212 10848 se
rect 1212 10835 1300 10848
tri 1300 10835 1313 10848 sw
tri 1435 10835 1448 10848 se
rect 1448 10835 1536 10848
tri 1536 10835 1549 10848 sw
tri 1671 10835 1684 10848 se
rect 1684 10835 1772 10848
tri 1772 10835 1785 10848 sw
tri 1907 10835 1920 10848 se
rect 1920 10835 2008 10848
tri 2008 10835 2021 10848 sw
tri 2143 10835 2156 10848 se
rect 2156 10835 2244 10848
tri 2244 10835 2257 10848 sw
tri 2379 10835 2392 10848 se
rect 2392 10835 2480 10848
tri 2480 10835 2493 10848 sw
tri 2615 10835 2628 10848 se
rect 2628 10835 2716 10848
tri 2716 10835 2729 10848 sw
tri 2851 10835 2864 10848 se
rect 2864 10835 3076 10848
rect 420 10829 3076 10835
rect 380 10813 3076 10829
rect 380 10810 697 10813
rect 380 10791 531 10810
rect 380 10757 386 10791
rect 420 10776 531 10791
rect 565 10776 697 10810
rect 420 10761 697 10776
rect 749 10761 765 10813
rect 817 10761 833 10813
rect 885 10761 901 10813
rect 953 10761 969 10813
rect 1021 10810 1037 10813
rect 1021 10761 1037 10776
rect 1089 10761 1105 10813
rect 1157 10761 1173 10813
rect 1225 10810 1241 10813
rect 1293 10810 2097 10813
rect 1225 10776 1239 10810
rect 1293 10776 1475 10810
rect 1509 10776 1711 10810
rect 1745 10776 1947 10810
rect 1981 10776 2097 10810
rect 1225 10761 1241 10776
rect 1293 10761 2097 10776
rect 2149 10761 2165 10813
rect 2217 10761 2233 10813
rect 2285 10761 2301 10813
rect 2353 10761 2369 10813
rect 2421 10810 2437 10813
rect 2421 10761 2437 10776
rect 2489 10761 2505 10813
rect 2557 10761 2573 10813
rect 2625 10761 2641 10813
rect 2693 10810 3076 10813
rect 2693 10776 2891 10810
rect 2925 10776 3036 10810
rect 3070 10776 3076 10810
rect 2693 10761 3076 10776
rect 420 10757 3076 10761
rect 380 10749 3076 10757
rect 380 10737 697 10749
rect 380 10719 531 10737
rect 380 10685 386 10719
rect 420 10703 531 10719
rect 565 10703 697 10737
rect 420 10697 697 10703
rect 749 10697 765 10749
rect 817 10697 833 10749
rect 885 10697 901 10749
rect 953 10697 969 10749
rect 1021 10737 1037 10749
rect 1021 10697 1037 10703
rect 1089 10697 1105 10749
rect 1157 10697 1173 10749
rect 1225 10737 1241 10749
rect 1293 10737 2097 10749
rect 1225 10703 1239 10737
rect 1293 10703 1475 10737
rect 1509 10703 1711 10737
rect 1745 10703 1947 10737
rect 1981 10703 2097 10737
rect 1225 10697 1241 10703
rect 1293 10697 2097 10703
rect 2149 10697 2165 10749
rect 2217 10697 2233 10749
rect 2285 10697 2301 10749
rect 2353 10697 2369 10749
rect 2421 10737 2437 10749
rect 2421 10697 2437 10703
rect 2489 10697 2505 10749
rect 2557 10697 2573 10749
rect 2625 10697 2641 10749
rect 2693 10738 3076 10749
rect 2693 10737 3036 10738
rect 2693 10703 2891 10737
rect 2925 10704 3036 10737
rect 3070 10704 3076 10738
rect 2925 10703 3076 10704
rect 2693 10697 3076 10703
rect 420 10685 3076 10697
rect 380 10664 697 10685
rect 380 10647 531 10664
rect 380 10613 386 10647
rect 420 10630 531 10647
rect 565 10633 697 10664
rect 749 10633 765 10685
rect 817 10633 833 10685
rect 885 10633 901 10685
rect 953 10633 969 10685
rect 1021 10664 1037 10685
rect 1089 10633 1105 10685
rect 1157 10633 1173 10685
rect 1225 10664 1241 10685
rect 1293 10664 2097 10685
rect 1225 10633 1239 10664
rect 1293 10633 1475 10664
rect 565 10630 767 10633
rect 801 10630 1003 10633
rect 1037 10630 1239 10633
rect 1273 10630 1475 10633
rect 1509 10630 1711 10664
rect 1745 10630 1947 10664
rect 1981 10633 2097 10664
rect 2149 10633 2165 10685
rect 2217 10633 2233 10685
rect 2285 10633 2301 10685
rect 2353 10633 2369 10685
rect 2421 10664 2437 10685
rect 2489 10633 2505 10685
rect 2557 10633 2573 10685
rect 2625 10633 2641 10685
rect 2693 10666 3076 10685
rect 2693 10664 3036 10666
rect 2693 10633 2891 10664
rect 1981 10630 2183 10633
rect 2217 10630 2419 10633
rect 2453 10630 2655 10633
rect 2689 10630 2891 10633
rect 2925 10632 3036 10664
rect 3070 10632 3076 10666
rect 2925 10630 3076 10632
rect 420 10621 3076 10630
rect 420 10613 697 10621
rect 380 10591 697 10613
rect 380 10575 531 10591
rect 380 10541 386 10575
rect 420 10557 531 10575
rect 565 10569 697 10591
rect 749 10569 765 10621
rect 817 10569 833 10621
rect 885 10569 901 10621
rect 953 10569 969 10621
rect 1021 10591 1037 10621
rect 1089 10569 1105 10621
rect 1157 10569 1173 10621
rect 1225 10591 1241 10621
rect 1293 10591 2097 10621
rect 1225 10569 1239 10591
rect 1293 10569 1475 10591
rect 565 10557 767 10569
rect 801 10557 1003 10569
rect 1037 10557 1239 10569
rect 1273 10557 1475 10569
rect 1509 10557 1711 10591
rect 1745 10557 1947 10591
rect 1981 10569 2097 10591
rect 2149 10569 2165 10621
rect 2217 10569 2233 10621
rect 2285 10569 2301 10621
rect 2353 10569 2369 10621
rect 2421 10591 2437 10621
rect 2489 10569 2505 10621
rect 2557 10569 2573 10621
rect 2625 10569 2641 10621
rect 2693 10594 3076 10621
rect 2693 10591 3036 10594
rect 2693 10569 2891 10591
rect 1981 10557 2183 10569
rect 2217 10557 2419 10569
rect 2453 10557 2655 10569
rect 2689 10557 2891 10569
rect 2925 10560 3036 10591
rect 3070 10560 3076 10594
rect 2925 10557 3076 10560
rect 420 10541 697 10557
rect 380 10518 697 10541
rect 380 10503 531 10518
rect 380 10469 386 10503
rect 420 10484 531 10503
rect 565 10505 697 10518
rect 749 10505 765 10557
rect 817 10505 833 10557
rect 885 10505 901 10557
rect 953 10505 969 10557
rect 1021 10518 1037 10557
rect 1089 10505 1105 10557
rect 1157 10505 1173 10557
rect 1225 10518 1241 10557
rect 1293 10518 2097 10557
rect 1225 10505 1239 10518
rect 1293 10505 1475 10518
rect 565 10493 767 10505
rect 801 10493 1003 10505
rect 1037 10493 1239 10505
rect 1273 10493 1475 10505
rect 565 10484 697 10493
rect 420 10469 697 10484
rect 380 10445 697 10469
rect 380 10431 531 10445
rect 380 10397 386 10431
rect 420 10411 531 10431
rect 565 10441 697 10445
rect 749 10441 765 10493
rect 817 10441 833 10493
rect 885 10441 901 10493
rect 953 10441 969 10493
rect 1021 10445 1037 10484
rect 1089 10441 1105 10493
rect 1157 10441 1173 10493
rect 1225 10484 1239 10493
rect 1293 10484 1475 10493
rect 1509 10484 1711 10518
rect 1745 10484 1947 10518
rect 1981 10505 2097 10518
rect 2149 10505 2165 10557
rect 2217 10505 2233 10557
rect 2285 10505 2301 10557
rect 2353 10505 2369 10557
rect 2421 10518 2437 10557
rect 2489 10505 2505 10557
rect 2557 10505 2573 10557
rect 2625 10505 2641 10557
rect 2693 10522 3076 10557
rect 2693 10518 3036 10522
rect 2693 10505 2891 10518
rect 1981 10493 2183 10505
rect 2217 10493 2419 10505
rect 2453 10493 2655 10505
rect 2689 10493 2891 10505
rect 1981 10484 2097 10493
rect 1225 10445 1241 10484
rect 1293 10445 2097 10484
rect 1225 10441 1239 10445
rect 1293 10441 1475 10445
rect 565 10429 767 10441
rect 801 10429 1003 10441
rect 1037 10429 1239 10441
rect 1273 10429 1475 10441
rect 565 10411 697 10429
rect 420 10397 697 10411
rect 380 10377 697 10397
rect 749 10377 765 10429
rect 817 10377 833 10429
rect 885 10377 901 10429
rect 953 10377 969 10429
rect 1021 10377 1037 10411
rect 1089 10377 1105 10429
rect 1157 10377 1173 10429
rect 1225 10411 1239 10429
rect 1293 10411 1475 10429
rect 1509 10411 1711 10445
rect 1745 10411 1947 10445
rect 1981 10441 2097 10445
rect 2149 10441 2165 10493
rect 2217 10441 2233 10493
rect 2285 10441 2301 10493
rect 2353 10441 2369 10493
rect 2421 10445 2437 10484
rect 2489 10441 2505 10493
rect 2557 10441 2573 10493
rect 2625 10441 2641 10493
rect 2693 10484 2891 10493
rect 2925 10488 3036 10518
rect 3070 10488 3076 10522
rect 2925 10484 3076 10488
rect 2693 10450 3076 10484
rect 2693 10445 3036 10450
rect 2693 10441 2891 10445
rect 1981 10429 2183 10441
rect 2217 10429 2419 10441
rect 2453 10429 2655 10441
rect 2689 10429 2891 10441
rect 1981 10411 2097 10429
rect 1225 10377 1241 10411
rect 1293 10377 2097 10411
rect 2149 10377 2165 10429
rect 2217 10377 2233 10429
rect 2285 10377 2301 10429
rect 2353 10377 2369 10429
rect 2421 10377 2437 10411
rect 2489 10377 2505 10429
rect 2557 10377 2573 10429
rect 2625 10377 2641 10429
rect 2693 10411 2891 10429
rect 2925 10416 3036 10445
rect 3070 10416 3076 10450
rect 2925 10411 3076 10416
rect 2693 10378 3076 10411
rect 2693 10377 3036 10378
rect 380 10372 3036 10377
rect 380 10359 531 10372
rect 380 10325 386 10359
rect 420 10338 531 10359
rect 565 10365 767 10372
rect 801 10365 1003 10372
rect 1037 10365 1239 10372
rect 1273 10365 1475 10372
rect 565 10338 697 10365
rect 420 10325 697 10338
rect 380 10313 697 10325
rect 749 10313 765 10365
rect 817 10313 833 10365
rect 885 10313 901 10365
rect 953 10313 969 10365
rect 1021 10313 1037 10338
rect 1089 10313 1105 10365
rect 1157 10313 1173 10365
rect 1225 10338 1239 10365
rect 1293 10338 1475 10365
rect 1509 10338 1711 10372
rect 1745 10338 1947 10372
rect 1981 10365 2183 10372
rect 2217 10365 2419 10372
rect 2453 10365 2655 10372
rect 2689 10365 2891 10372
rect 1981 10338 2097 10365
rect 1225 10313 1241 10338
rect 1293 10313 2097 10338
rect 2149 10313 2165 10365
rect 2217 10313 2233 10365
rect 2285 10313 2301 10365
rect 2353 10313 2369 10365
rect 2421 10313 2437 10338
rect 2489 10313 2505 10365
rect 2557 10313 2573 10365
rect 2625 10313 2641 10365
rect 2693 10338 2891 10365
rect 2925 10344 3036 10372
rect 3070 10344 3076 10378
rect 2925 10338 3076 10344
rect 2693 10313 3076 10338
rect 380 10306 3076 10313
rect 380 10301 3036 10306
rect 380 10298 697 10301
rect 380 10287 531 10298
rect 380 10253 386 10287
rect 420 10264 531 10287
rect 565 10264 697 10298
rect 420 10253 697 10264
rect 380 10249 697 10253
rect 749 10249 765 10301
rect 817 10249 833 10301
rect 885 10249 901 10301
rect 953 10249 969 10301
rect 1021 10298 1037 10301
rect 1021 10249 1037 10264
rect 1089 10249 1105 10301
rect 1157 10249 1173 10301
rect 1225 10298 1241 10301
rect 1293 10298 2097 10301
rect 1225 10264 1239 10298
rect 1293 10264 1475 10298
rect 1509 10264 1711 10298
rect 1745 10264 1947 10298
rect 1981 10264 2097 10298
rect 1225 10249 1241 10264
rect 1293 10249 2097 10264
rect 2149 10249 2165 10301
rect 2217 10249 2233 10301
rect 2285 10249 2301 10301
rect 2353 10249 2369 10301
rect 2421 10298 2437 10301
rect 2421 10249 2437 10264
rect 2489 10249 2505 10301
rect 2557 10249 2573 10301
rect 2625 10249 2641 10301
rect 2693 10298 3036 10301
rect 2693 10264 2891 10298
rect 2925 10272 3036 10298
rect 3070 10272 3076 10306
rect 2925 10264 3076 10272
rect 2693 10249 3076 10264
rect 380 10237 3076 10249
rect 380 10224 697 10237
rect 380 10215 531 10224
rect 380 10181 386 10215
rect 420 10190 531 10215
rect 565 10190 697 10224
rect 420 10185 697 10190
rect 749 10185 765 10237
rect 817 10185 833 10237
rect 885 10185 901 10237
rect 953 10185 969 10237
rect 1021 10224 1037 10237
rect 1021 10185 1037 10190
rect 1089 10185 1105 10237
rect 1157 10185 1173 10237
rect 1225 10224 1241 10237
rect 1293 10224 2097 10237
rect 1225 10190 1239 10224
rect 1293 10190 1475 10224
rect 1509 10190 1711 10224
rect 1745 10190 1947 10224
rect 1981 10190 2097 10224
rect 1225 10185 1241 10190
rect 1293 10185 2097 10190
rect 2149 10185 2165 10237
rect 2217 10185 2233 10237
rect 2285 10185 2301 10237
rect 2353 10185 2369 10237
rect 2421 10224 2437 10237
rect 2421 10185 2437 10190
rect 2489 10185 2505 10237
rect 2557 10185 2573 10237
rect 2625 10185 2641 10237
rect 2693 10234 3076 10237
rect 2693 10224 3036 10234
rect 2693 10190 2891 10224
rect 2925 10200 3036 10224
rect 3070 10200 3076 10234
rect 2925 10190 3076 10200
rect 2693 10185 3076 10190
rect 420 10181 3076 10185
rect 380 10173 3076 10181
rect 380 10150 697 10173
rect 380 10143 531 10150
rect 380 10109 386 10143
rect 420 10116 531 10143
rect 565 10121 697 10150
rect 749 10121 765 10173
rect 817 10121 833 10173
rect 885 10121 901 10173
rect 953 10121 969 10173
rect 1021 10150 1037 10173
rect 1089 10121 1105 10173
rect 1157 10121 1173 10173
rect 1225 10150 1241 10173
rect 1293 10150 2097 10173
rect 1225 10121 1239 10150
rect 1293 10121 1475 10150
rect 565 10116 767 10121
rect 801 10116 1003 10121
rect 1037 10116 1239 10121
rect 1273 10116 1475 10121
rect 1509 10116 1711 10150
rect 1745 10116 1947 10150
rect 1981 10121 2097 10150
rect 2149 10121 2165 10173
rect 2217 10121 2233 10173
rect 2285 10121 2301 10173
rect 2353 10121 2369 10173
rect 2421 10150 2437 10173
rect 2489 10121 2505 10173
rect 2557 10121 2573 10173
rect 2625 10121 2641 10173
rect 2693 10162 3076 10173
rect 2693 10150 3036 10162
rect 2693 10121 2891 10150
rect 1981 10116 2183 10121
rect 2217 10116 2419 10121
rect 2453 10116 2655 10121
rect 2689 10116 2891 10121
rect 2925 10128 3036 10150
rect 3070 10128 3076 10162
rect 2925 10116 3076 10128
rect 420 10109 3076 10116
rect 380 10076 697 10109
rect 380 10071 531 10076
rect 380 10037 386 10071
rect 420 10042 531 10071
rect 565 10057 697 10076
rect 749 10057 765 10109
rect 817 10057 833 10109
rect 885 10057 901 10109
rect 953 10057 969 10109
rect 1021 10076 1037 10109
rect 1089 10057 1105 10109
rect 1157 10057 1173 10109
rect 1225 10076 1241 10109
rect 1293 10076 2097 10109
rect 1225 10057 1239 10076
rect 1293 10057 1475 10076
rect 565 10045 767 10057
rect 801 10045 1003 10057
rect 1037 10045 1239 10057
rect 1273 10045 1475 10057
rect 565 10042 697 10045
rect 420 10037 697 10042
rect 380 10002 697 10037
rect 380 9999 531 10002
rect 380 9965 386 9999
rect 420 9968 531 9999
rect 565 9993 697 10002
rect 749 9993 765 10045
rect 817 9993 833 10045
rect 885 9993 901 10045
rect 953 9993 969 10045
rect 1021 10002 1037 10042
rect 1089 9993 1105 10045
rect 1157 9993 1173 10045
rect 1225 10042 1239 10045
rect 1293 10042 1475 10045
rect 1509 10042 1711 10076
rect 1745 10042 1947 10076
rect 1981 10057 2097 10076
rect 2149 10057 2165 10109
rect 2217 10057 2233 10109
rect 2285 10057 2301 10109
rect 2353 10057 2369 10109
rect 2421 10076 2437 10109
rect 2489 10057 2505 10109
rect 2557 10057 2573 10109
rect 2625 10057 2641 10109
rect 2693 10090 3076 10109
rect 2693 10076 3036 10090
rect 2693 10057 2891 10076
rect 1981 10045 2183 10057
rect 2217 10045 2419 10057
rect 2453 10045 2655 10057
rect 2689 10045 2891 10057
rect 1981 10042 2097 10045
rect 1225 10002 1241 10042
rect 1293 10002 2097 10042
rect 1225 9993 1239 10002
rect 1293 9993 1475 10002
rect 565 9981 767 9993
rect 801 9981 1003 9993
rect 1037 9981 1239 9993
rect 1273 9981 1475 9993
rect 565 9968 697 9981
rect 420 9965 697 9968
rect 380 9929 697 9965
rect 749 9929 765 9981
rect 817 9929 833 9981
rect 885 9929 901 9981
rect 953 9929 969 9981
rect 1021 9929 1037 9968
rect 1089 9929 1105 9981
rect 1157 9929 1173 9981
rect 1225 9968 1239 9981
rect 1293 9968 1475 9981
rect 1509 9968 1711 10002
rect 1745 9968 1947 10002
rect 1981 9993 2097 10002
rect 2149 9993 2165 10045
rect 2217 9993 2233 10045
rect 2285 9993 2301 10045
rect 2353 9993 2369 10045
rect 2421 10002 2437 10042
rect 2489 9993 2505 10045
rect 2557 9993 2573 10045
rect 2625 9993 2641 10045
rect 2693 10042 2891 10045
rect 2925 10056 3036 10076
rect 3070 10056 3076 10090
rect 2925 10042 3076 10056
rect 2693 10018 3076 10042
rect 2693 10002 3036 10018
rect 2693 9993 2891 10002
rect 1981 9981 2183 9993
rect 2217 9981 2419 9993
rect 2453 9981 2655 9993
rect 2689 9981 2891 9993
rect 1981 9968 2097 9981
rect 1225 9929 1241 9968
rect 1293 9929 2097 9968
rect 2149 9929 2165 9981
rect 2217 9929 2233 9981
rect 2285 9929 2301 9981
rect 2353 9929 2369 9981
rect 2421 9929 2437 9968
rect 2489 9929 2505 9981
rect 2557 9929 2573 9981
rect 2625 9929 2641 9981
rect 2693 9968 2891 9981
rect 2925 9984 3036 10002
rect 3070 9984 3076 10018
rect 2925 9968 3076 9984
rect 2693 9946 3076 9968
rect 2693 9929 3036 9946
rect 380 9928 3036 9929
rect 380 9927 531 9928
rect 380 9893 386 9927
rect 420 9894 531 9927
rect 565 9917 767 9928
rect 801 9917 1003 9928
rect 1037 9917 1239 9928
rect 1273 9917 1475 9928
rect 565 9894 697 9917
rect 420 9893 697 9894
rect 380 9865 697 9893
rect 749 9865 765 9917
rect 817 9865 833 9917
rect 885 9865 901 9917
rect 953 9865 969 9917
rect 1021 9865 1037 9894
rect 1089 9865 1105 9917
rect 1157 9865 1173 9917
rect 1225 9894 1239 9917
rect 1293 9894 1475 9917
rect 1509 9894 1711 9928
rect 1745 9894 1947 9928
rect 1981 9917 2183 9928
rect 2217 9917 2419 9928
rect 2453 9917 2655 9928
rect 2689 9917 2891 9928
rect 1981 9894 2097 9917
rect 1225 9865 1241 9894
rect 1293 9865 2097 9894
rect 2149 9865 2165 9917
rect 2217 9865 2233 9917
rect 2285 9865 2301 9917
rect 2353 9865 2369 9917
rect 2421 9865 2437 9894
rect 2489 9865 2505 9917
rect 2557 9865 2573 9917
rect 2625 9865 2641 9917
rect 2693 9894 2891 9917
rect 2925 9912 3036 9928
rect 3070 9912 3076 9946
rect 2925 9894 3076 9912
rect 2693 9874 3076 9894
rect 2693 9865 3036 9874
rect 380 9855 3036 9865
rect 380 9821 386 9855
rect 420 9854 3036 9855
rect 420 9821 531 9854
rect 380 9820 531 9821
rect 565 9835 767 9854
rect 565 9820 590 9835
tri 590 9820 605 9835 nw
tri 727 9820 742 9835 ne
rect 742 9820 767 9835
rect 801 9835 1003 9854
rect 801 9820 826 9835
tri 826 9820 841 9835 nw
tri 963 9820 978 9835 ne
rect 978 9820 1003 9835
rect 1037 9835 1239 9854
rect 1037 9820 1062 9835
tri 1062 9820 1077 9835 nw
tri 1199 9820 1214 9835 ne
rect 1214 9820 1239 9835
rect 1273 9835 1475 9854
rect 1273 9820 1298 9835
tri 1298 9820 1313 9835 nw
tri 1435 9820 1450 9835 ne
rect 1450 9820 1475 9835
rect 1509 9835 1711 9854
rect 1509 9820 1534 9835
tri 1534 9820 1549 9835 nw
tri 1671 9820 1686 9835 ne
rect 1686 9820 1711 9835
rect 1745 9835 1947 9854
rect 1745 9820 1770 9835
tri 1770 9820 1785 9835 nw
tri 1907 9820 1922 9835 ne
rect 1922 9820 1947 9835
rect 1981 9835 2183 9854
rect 1981 9820 2006 9835
tri 2006 9820 2021 9835 nw
tri 2143 9820 2158 9835 ne
rect 2158 9820 2183 9835
rect 2217 9835 2419 9854
rect 2217 9820 2242 9835
tri 2242 9820 2257 9835 nw
tri 2379 9820 2394 9835 ne
rect 2394 9820 2419 9835
rect 2453 9835 2655 9854
rect 2453 9820 2478 9835
tri 2478 9820 2493 9835 nw
tri 2615 9820 2630 9835 ne
rect 2630 9820 2655 9835
rect 2689 9835 2891 9854
rect 2689 9820 2714 9835
tri 2714 9820 2729 9835 nw
tri 2851 9820 2866 9835 ne
rect 2866 9820 2891 9835
rect 2925 9840 3036 9854
rect 3070 9840 3076 9874
rect 2925 9820 3076 9840
rect 380 9816 586 9820
tri 586 9816 590 9820 nw
tri 742 9816 746 9820 ne
rect 746 9816 822 9820
tri 822 9816 826 9820 nw
tri 978 9816 982 9820 ne
rect 982 9816 1058 9820
tri 1058 9816 1062 9820 nw
tri 1214 9816 1218 9820 ne
rect 1218 9816 1294 9820
tri 1294 9816 1298 9820 nw
tri 1450 9816 1454 9820 ne
rect 1454 9816 1530 9820
tri 1530 9816 1534 9820 nw
tri 1686 9816 1690 9820 ne
rect 1690 9816 1766 9820
tri 1766 9816 1770 9820 nw
tri 1922 9816 1926 9820 ne
rect 1926 9816 2002 9820
tri 2002 9816 2006 9820 nw
tri 2158 9816 2162 9820 ne
rect 2162 9816 2238 9820
tri 2238 9816 2242 9820 nw
tri 2394 9816 2398 9820 ne
rect 2398 9816 2474 9820
tri 2474 9816 2478 9820 nw
tri 2630 9816 2634 9820 ne
rect 2634 9816 2710 9820
tri 2710 9816 2714 9820 nw
tri 2866 9816 2870 9820 ne
rect 2870 9816 3076 9820
rect 380 9802 572 9816
tri 572 9802 586 9816 nw
tri 746 9802 760 9816 ne
rect 760 9802 808 9816
tri 808 9802 822 9816 nw
tri 982 9802 996 9816 ne
rect 996 9802 1044 9816
tri 1044 9802 1058 9816 nw
tri 1218 9802 1232 9816 ne
rect 1232 9802 1280 9816
tri 1280 9802 1294 9816 nw
tri 1454 9802 1468 9816 ne
rect 1468 9802 1516 9816
tri 1516 9802 1530 9816 nw
tri 1690 9802 1704 9816 ne
rect 1704 9802 1752 9816
tri 1752 9802 1766 9816 nw
tri 1926 9802 1940 9816 ne
rect 1940 9802 1988 9816
tri 1988 9802 2002 9816 nw
tri 2162 9802 2176 9816 ne
rect 2176 9802 2224 9816
tri 2224 9802 2238 9816 nw
tri 2398 9802 2412 9816 ne
rect 2412 9802 2460 9816
tri 2460 9802 2474 9816 nw
tri 2634 9802 2648 9816 ne
rect 2648 9802 2696 9816
tri 2696 9802 2710 9816 nw
tri 2870 9802 2884 9816 ne
rect 2884 9802 3076 9816
rect 380 9783 571 9802
tri 571 9801 572 9802 nw
tri 760 9801 761 9802 ne
rect 380 9749 386 9783
rect 420 9780 571 9783
rect 420 9749 531 9780
rect 380 9746 531 9749
rect 565 9746 571 9780
rect 380 9711 571 9746
rect 380 9677 386 9711
rect 420 9706 571 9711
rect 420 9677 531 9706
rect 380 9672 531 9677
rect 565 9672 571 9706
rect 380 9639 571 9672
rect 380 9605 386 9639
rect 420 9632 571 9639
rect 420 9605 531 9632
rect 380 9598 531 9605
rect 565 9598 571 9632
rect 380 9567 571 9598
rect 380 9533 386 9567
rect 420 9558 571 9567
rect 420 9533 531 9558
rect 380 9524 531 9533
rect 565 9524 571 9558
rect 380 9495 571 9524
rect 380 9461 386 9495
rect 420 9484 571 9495
rect 420 9461 531 9484
rect 380 9450 531 9461
rect 565 9450 571 9484
rect 380 9423 571 9450
rect 380 9389 386 9423
rect 420 9410 571 9423
rect 420 9389 531 9410
rect 380 9376 531 9389
rect 565 9376 571 9410
rect 380 9351 571 9376
rect 380 9317 386 9351
rect 420 9336 571 9351
rect 420 9317 531 9336
rect 380 9302 531 9317
rect 565 9302 571 9336
rect 380 9279 571 9302
rect 761 9780 807 9802
tri 807 9801 808 9802 nw
tri 996 9801 997 9802 ne
rect 761 9746 767 9780
rect 801 9746 807 9780
rect 761 9706 807 9746
rect 761 9672 767 9706
rect 801 9672 807 9706
rect 761 9632 807 9672
rect 761 9598 767 9632
rect 801 9598 807 9632
rect 761 9558 807 9598
rect 761 9524 767 9558
rect 801 9524 807 9558
rect 761 9484 807 9524
rect 761 9450 767 9484
rect 801 9450 807 9484
rect 761 9410 807 9450
rect 761 9376 767 9410
rect 801 9376 807 9410
rect 761 9336 807 9376
rect 761 9302 767 9336
rect 801 9302 807 9336
rect 761 9290 807 9302
rect 997 9780 1043 9802
tri 1043 9801 1044 9802 nw
tri 1232 9801 1233 9802 ne
rect 997 9746 1003 9780
rect 1037 9746 1043 9780
rect 997 9706 1043 9746
rect 997 9672 1003 9706
rect 1037 9672 1043 9706
rect 997 9632 1043 9672
rect 997 9598 1003 9632
rect 1037 9598 1043 9632
rect 997 9558 1043 9598
rect 997 9524 1003 9558
rect 1037 9524 1043 9558
rect 997 9484 1043 9524
rect 997 9450 1003 9484
rect 1037 9450 1043 9484
rect 997 9410 1043 9450
rect 997 9376 1003 9410
rect 1037 9376 1043 9410
rect 997 9336 1043 9376
rect 997 9302 1003 9336
rect 1037 9302 1043 9336
rect 997 9290 1043 9302
rect 1233 9780 1279 9802
tri 1279 9801 1280 9802 nw
tri 1468 9801 1469 9802 ne
rect 1233 9746 1239 9780
rect 1273 9746 1279 9780
rect 1233 9706 1279 9746
rect 1233 9672 1239 9706
rect 1273 9672 1279 9706
rect 1233 9632 1279 9672
rect 1233 9598 1239 9632
rect 1273 9598 1279 9632
rect 1233 9558 1279 9598
rect 1233 9524 1239 9558
rect 1273 9524 1279 9558
rect 1233 9484 1279 9524
rect 1233 9450 1239 9484
rect 1273 9450 1279 9484
rect 1233 9410 1279 9450
rect 1233 9376 1239 9410
rect 1273 9376 1279 9410
rect 1233 9336 1279 9376
rect 1233 9302 1239 9336
rect 1273 9302 1279 9336
rect 1233 9290 1279 9302
rect 1469 9780 1515 9802
tri 1515 9801 1516 9802 nw
tri 1704 9801 1705 9802 ne
rect 1469 9746 1475 9780
rect 1509 9746 1515 9780
rect 1469 9706 1515 9746
rect 1469 9672 1475 9706
rect 1509 9672 1515 9706
rect 1469 9632 1515 9672
rect 1469 9598 1475 9632
rect 1509 9598 1515 9632
rect 1469 9558 1515 9598
rect 1469 9524 1475 9558
rect 1509 9524 1515 9558
rect 1469 9484 1515 9524
rect 1469 9450 1475 9484
rect 1509 9450 1515 9484
rect 1469 9410 1515 9450
rect 1469 9376 1475 9410
rect 1509 9376 1515 9410
rect 1469 9336 1515 9376
rect 1469 9302 1475 9336
rect 1509 9302 1515 9336
rect 1469 9290 1515 9302
rect 1705 9780 1751 9802
tri 1751 9801 1752 9802 nw
tri 1940 9801 1941 9802 ne
rect 1705 9746 1711 9780
rect 1745 9746 1751 9780
rect 1705 9706 1751 9746
rect 1705 9672 1711 9706
rect 1745 9672 1751 9706
rect 1705 9632 1751 9672
rect 1705 9598 1711 9632
rect 1745 9598 1751 9632
rect 1705 9558 1751 9598
rect 1705 9524 1711 9558
rect 1745 9524 1751 9558
rect 1705 9484 1751 9524
rect 1705 9450 1711 9484
rect 1745 9450 1751 9484
rect 1705 9410 1751 9450
rect 1705 9376 1711 9410
rect 1745 9376 1751 9410
rect 1705 9336 1751 9376
rect 1705 9302 1711 9336
rect 1745 9302 1751 9336
rect 1705 9290 1751 9302
rect 1941 9780 1987 9802
tri 1987 9801 1988 9802 nw
tri 2176 9801 2177 9802 ne
rect 1941 9746 1947 9780
rect 1981 9746 1987 9780
rect 1941 9706 1987 9746
rect 1941 9672 1947 9706
rect 1981 9672 1987 9706
rect 1941 9632 1987 9672
rect 1941 9598 1947 9632
rect 1981 9598 1987 9632
rect 1941 9558 1987 9598
rect 1941 9524 1947 9558
rect 1981 9524 1987 9558
rect 1941 9484 1987 9524
rect 1941 9450 1947 9484
rect 1981 9450 1987 9484
rect 1941 9410 1987 9450
rect 1941 9376 1947 9410
rect 1981 9376 1987 9410
rect 1941 9336 1987 9376
rect 1941 9302 1947 9336
rect 1981 9302 1987 9336
rect 1941 9290 1987 9302
rect 2177 9780 2223 9802
tri 2223 9801 2224 9802 nw
tri 2412 9801 2413 9802 ne
rect 2177 9746 2183 9780
rect 2217 9746 2223 9780
rect 2177 9706 2223 9746
rect 2177 9672 2183 9706
rect 2217 9672 2223 9706
rect 2177 9632 2223 9672
rect 2177 9598 2183 9632
rect 2217 9598 2223 9632
rect 2177 9558 2223 9598
rect 2177 9524 2183 9558
rect 2217 9524 2223 9558
rect 2177 9484 2223 9524
rect 2177 9450 2183 9484
rect 2217 9450 2223 9484
rect 2177 9410 2223 9450
rect 2177 9376 2183 9410
rect 2217 9376 2223 9410
rect 2177 9336 2223 9376
rect 2177 9302 2183 9336
rect 2217 9302 2223 9336
rect 2177 9290 2223 9302
rect 2413 9780 2459 9802
tri 2459 9801 2460 9802 nw
tri 2648 9801 2649 9802 ne
rect 2413 9746 2419 9780
rect 2453 9746 2459 9780
rect 2413 9706 2459 9746
rect 2413 9672 2419 9706
rect 2453 9672 2459 9706
rect 2413 9632 2459 9672
rect 2413 9598 2419 9632
rect 2453 9598 2459 9632
rect 2413 9558 2459 9598
rect 2413 9524 2419 9558
rect 2453 9524 2459 9558
rect 2413 9484 2459 9524
rect 2413 9450 2419 9484
rect 2453 9450 2459 9484
rect 2413 9410 2459 9450
rect 2413 9376 2419 9410
rect 2453 9376 2459 9410
rect 2413 9336 2459 9376
rect 2413 9302 2419 9336
rect 2453 9302 2459 9336
rect 2413 9290 2459 9302
rect 2649 9780 2695 9802
tri 2695 9801 2696 9802 nw
tri 2884 9801 2885 9802 ne
rect 2649 9746 2655 9780
rect 2689 9746 2695 9780
rect 2649 9706 2695 9746
rect 2649 9672 2655 9706
rect 2689 9672 2695 9706
rect 2649 9632 2695 9672
rect 2649 9598 2655 9632
rect 2689 9598 2695 9632
rect 2649 9558 2695 9598
rect 2649 9524 2655 9558
rect 2689 9524 2695 9558
rect 2649 9484 2695 9524
rect 2649 9450 2655 9484
rect 2689 9450 2695 9484
rect 2649 9410 2695 9450
rect 2649 9376 2655 9410
rect 2689 9376 2695 9410
rect 2649 9336 2695 9376
rect 2649 9302 2655 9336
rect 2689 9302 2695 9336
rect 2649 9290 2695 9302
rect 2885 9780 3036 9802
rect 2885 9746 2891 9780
rect 2925 9768 3036 9780
rect 3070 9768 3076 9802
rect 2925 9746 3076 9768
rect 2885 9730 3076 9746
rect 2885 9706 3036 9730
rect 2885 9672 2891 9706
rect 2925 9696 3036 9706
rect 3070 9696 3076 9730
rect 2925 9672 3076 9696
rect 2885 9658 3076 9672
rect 2885 9632 3036 9658
rect 2885 9598 2891 9632
rect 2925 9624 3036 9632
rect 3070 9624 3076 9658
rect 2925 9598 3076 9624
rect 2885 9586 3076 9598
rect 2885 9558 3036 9586
rect 2885 9524 2891 9558
rect 2925 9552 3036 9558
rect 3070 9552 3076 9586
rect 2925 9524 3076 9552
rect 2885 9514 3076 9524
rect 2885 9484 3036 9514
rect 2885 9450 2891 9484
rect 2925 9480 3036 9484
rect 3070 9480 3076 9514
rect 2925 9450 3076 9480
rect 2885 9442 3076 9450
rect 2885 9410 3036 9442
rect 2885 9376 2891 9410
rect 2925 9408 3036 9410
rect 3070 9408 3076 9442
rect 2925 9376 3076 9408
rect 2885 9370 3076 9376
rect 2885 9336 3036 9370
rect 3070 9336 3076 9370
rect 2885 9302 2891 9336
rect 2925 9302 3076 9336
rect 2885 9298 3076 9302
rect 380 9245 386 9279
rect 420 9245 571 9279
rect 380 9207 571 9245
rect 2885 9264 3036 9298
rect 3070 9264 3076 9298
rect 380 9173 386 9207
rect 420 9173 571 9207
rect 613 9234 1501 9243
rect 1553 9234 1569 9243
rect 1621 9234 1636 9243
rect 1688 9234 1703 9243
rect 1755 9234 1770 9243
rect 1822 9234 1837 9243
rect 1889 9234 2830 9243
rect 613 9200 625 9234
rect 659 9200 700 9234
rect 734 9200 775 9234
rect 809 9200 850 9234
rect 884 9200 925 9234
rect 959 9200 1000 9234
rect 1034 9200 1075 9234
rect 1109 9200 1150 9234
rect 1184 9200 1225 9234
rect 1259 9200 1300 9234
rect 1334 9200 1375 9234
rect 1409 9200 1450 9234
rect 1484 9200 1501 9234
rect 1559 9200 1569 9234
rect 1634 9200 1636 9234
rect 1889 9200 1896 9234
rect 1930 9200 1970 9234
rect 2004 9200 2044 9234
rect 2078 9200 2118 9234
rect 2152 9200 2192 9234
rect 2226 9200 2266 9234
rect 2300 9200 2340 9234
rect 2374 9200 2414 9234
rect 2448 9200 2488 9234
rect 2522 9200 2562 9234
rect 2596 9200 2636 9234
rect 2670 9200 2710 9234
rect 2744 9200 2784 9234
rect 2818 9200 2830 9234
rect 613 9191 1501 9200
rect 1553 9191 1569 9200
rect 1621 9191 1636 9200
rect 1688 9191 1703 9200
rect 1755 9191 1770 9200
rect 1822 9191 1837 9200
rect 1889 9191 2830 9200
rect 2885 9226 3076 9264
rect 2885 9192 3036 9226
rect 3070 9192 3076 9226
rect 380 9135 571 9173
rect 2885 9154 3076 9192
rect 380 9101 386 9135
rect 420 9132 571 9135
rect 420 9101 531 9132
rect 380 9098 531 9101
rect 565 9098 571 9132
rect 380 9063 571 9098
rect 380 9029 386 9063
rect 420 9059 571 9063
rect 420 9029 531 9059
rect 380 9025 531 9029
rect 565 9025 571 9059
rect 380 8991 571 9025
rect 380 8957 386 8991
rect 420 8986 571 8991
rect 420 8957 531 8986
rect 380 8952 531 8957
rect 565 8952 571 8986
rect 380 8919 571 8952
rect 380 8885 386 8919
rect 420 8913 571 8919
rect 420 8885 531 8913
rect 380 8879 531 8885
rect 565 8879 571 8913
rect 380 8847 571 8879
rect 380 8813 386 8847
rect 420 8840 571 8847
rect 420 8813 531 8840
rect 380 8806 531 8813
rect 565 8806 571 8840
rect 380 8775 571 8806
rect 380 8741 386 8775
rect 420 8767 571 8775
rect 420 8741 531 8767
rect 380 8733 531 8741
rect 565 8733 571 8767
rect 380 8703 571 8733
rect 380 8669 386 8703
rect 420 8694 571 8703
rect 420 8669 531 8694
rect 380 8660 531 8669
rect 565 8660 571 8694
rect 761 9132 807 9144
rect 761 9098 767 9132
rect 801 9098 807 9132
rect 761 9059 807 9098
rect 761 9025 767 9059
rect 801 9025 807 9059
rect 761 8986 807 9025
rect 761 8952 767 8986
rect 801 8952 807 8986
rect 761 8913 807 8952
rect 761 8879 767 8913
rect 801 8879 807 8913
rect 761 8840 807 8879
rect 761 8806 767 8840
rect 801 8806 807 8840
rect 761 8767 807 8806
rect 761 8733 767 8767
rect 801 8733 807 8767
rect 761 8694 807 8733
tri 571 8660 583 8672 sw
tri 749 8660 761 8672 se
rect 761 8660 767 8694
rect 801 8660 807 8694
rect 997 9132 1043 9144
rect 997 9098 1003 9132
rect 1037 9098 1043 9132
rect 997 9059 1043 9098
rect 997 9025 1003 9059
rect 1037 9025 1043 9059
rect 997 8986 1043 9025
rect 997 8952 1003 8986
rect 1037 8952 1043 8986
rect 997 8913 1043 8952
rect 997 8879 1003 8913
rect 1037 8879 1043 8913
rect 997 8840 1043 8879
rect 997 8806 1003 8840
rect 1037 8806 1043 8840
rect 997 8767 1043 8806
rect 997 8733 1003 8767
rect 1037 8733 1043 8767
rect 997 8694 1043 8733
tri 807 8660 819 8672 sw
tri 985 8660 997 8672 se
rect 997 8660 1003 8694
rect 1037 8660 1043 8694
rect 1233 9132 1279 9144
rect 1233 9098 1239 9132
rect 1273 9098 1279 9132
rect 1233 9059 1279 9098
rect 1233 9025 1239 9059
rect 1273 9025 1279 9059
rect 1233 8986 1279 9025
rect 1233 8952 1239 8986
rect 1273 8952 1279 8986
rect 1233 8913 1279 8952
rect 1233 8879 1239 8913
rect 1273 8879 1279 8913
rect 1233 8840 1279 8879
rect 1233 8806 1239 8840
rect 1273 8806 1279 8840
rect 1233 8767 1279 8806
rect 1233 8733 1239 8767
rect 1273 8733 1279 8767
rect 1233 8694 1279 8733
tri 1043 8660 1055 8672 sw
tri 1221 8660 1233 8672 se
rect 1233 8660 1239 8694
rect 1273 8660 1279 8694
rect 1469 9132 1515 9144
rect 1469 9098 1475 9132
rect 1509 9098 1515 9132
rect 1469 9059 1515 9098
rect 1469 9025 1475 9059
rect 1509 9025 1515 9059
rect 1469 8986 1515 9025
rect 1469 8952 1475 8986
rect 1509 8952 1515 8986
rect 1469 8913 1515 8952
rect 1469 8879 1475 8913
rect 1509 8879 1515 8913
rect 1469 8840 1515 8879
rect 1469 8806 1475 8840
rect 1509 8806 1515 8840
rect 1469 8767 1515 8806
rect 1469 8733 1475 8767
rect 1509 8733 1515 8767
rect 1469 8694 1515 8733
tri 1279 8660 1291 8672 sw
tri 1457 8660 1469 8672 se
rect 1469 8660 1475 8694
rect 1509 8660 1515 8694
rect 1705 9132 1751 9144
rect 1705 9098 1711 9132
rect 1745 9098 1751 9132
rect 1705 9059 1751 9098
rect 1705 9025 1711 9059
rect 1745 9025 1751 9059
rect 1705 8986 1751 9025
rect 1705 8952 1711 8986
rect 1745 8952 1751 8986
rect 1705 8913 1751 8952
rect 1705 8879 1711 8913
rect 1745 8879 1751 8913
rect 1705 8840 1751 8879
rect 1705 8806 1711 8840
rect 1745 8806 1751 8840
rect 1705 8767 1751 8806
rect 1705 8733 1711 8767
rect 1745 8733 1751 8767
rect 1705 8694 1751 8733
tri 1515 8660 1527 8672 sw
tri 1693 8660 1705 8672 se
rect 1705 8660 1711 8694
rect 1745 8660 1751 8694
rect 1941 9132 1987 9144
rect 1941 9098 1947 9132
rect 1981 9098 1987 9132
rect 1941 9059 1987 9098
rect 1941 9025 1947 9059
rect 1981 9025 1987 9059
rect 1941 8986 1987 9025
rect 1941 8952 1947 8986
rect 1981 8952 1987 8986
rect 1941 8913 1987 8952
rect 1941 8879 1947 8913
rect 1981 8879 1987 8913
rect 1941 8840 1987 8879
rect 1941 8806 1947 8840
rect 1981 8806 1987 8840
rect 1941 8767 1987 8806
rect 1941 8733 1947 8767
rect 1981 8733 1987 8767
rect 1941 8694 1987 8733
tri 1751 8660 1763 8672 sw
tri 1929 8660 1941 8672 se
rect 1941 8660 1947 8694
rect 1981 8660 1987 8694
rect 2177 9132 2223 9144
rect 2177 9098 2183 9132
rect 2217 9098 2223 9132
rect 2177 9059 2223 9098
rect 2177 9025 2183 9059
rect 2217 9025 2223 9059
rect 2177 8986 2223 9025
rect 2177 8952 2183 8986
rect 2217 8952 2223 8986
rect 2177 8913 2223 8952
rect 2177 8879 2183 8913
rect 2217 8879 2223 8913
rect 2177 8840 2223 8879
rect 2177 8806 2183 8840
rect 2217 8806 2223 8840
rect 2177 8767 2223 8806
rect 2177 8733 2183 8767
rect 2217 8733 2223 8767
rect 2177 8694 2223 8733
tri 1987 8660 1999 8672 sw
tri 2165 8660 2177 8672 se
rect 2177 8660 2183 8694
rect 2217 8660 2223 8694
rect 2413 9132 2459 9144
rect 2413 9098 2419 9132
rect 2453 9098 2459 9132
rect 2413 9059 2459 9098
rect 2413 9025 2419 9059
rect 2453 9025 2459 9059
rect 2413 8986 2459 9025
rect 2413 8952 2419 8986
rect 2453 8952 2459 8986
rect 2413 8913 2459 8952
rect 2413 8879 2419 8913
rect 2453 8879 2459 8913
rect 2413 8840 2459 8879
rect 2413 8806 2419 8840
rect 2453 8806 2459 8840
rect 2413 8767 2459 8806
rect 2413 8733 2419 8767
rect 2453 8733 2459 8767
rect 2413 8694 2459 8733
tri 2223 8660 2235 8672 sw
tri 2401 8660 2413 8672 se
rect 2413 8660 2419 8694
rect 2453 8660 2459 8694
rect 2649 9132 2695 9144
rect 2649 9098 2655 9132
rect 2689 9098 2695 9132
rect 2649 9059 2695 9098
rect 2649 9025 2655 9059
rect 2689 9025 2695 9059
rect 2649 8986 2695 9025
rect 2649 8952 2655 8986
rect 2689 8952 2695 8986
rect 2649 8913 2695 8952
rect 2649 8879 2655 8913
rect 2689 8879 2695 8913
rect 2649 8840 2695 8879
rect 2649 8806 2655 8840
rect 2689 8806 2695 8840
rect 2649 8767 2695 8806
rect 2649 8733 2655 8767
rect 2689 8733 2695 8767
rect 2649 8694 2695 8733
tri 2459 8660 2471 8672 sw
tri 2637 8660 2649 8672 se
rect 2649 8660 2655 8694
rect 2689 8660 2695 8694
rect 2885 9132 3036 9154
rect 2885 9098 2891 9132
rect 2925 9120 3036 9132
rect 3070 9120 3076 9154
rect 2925 9098 3076 9120
rect 2885 9082 3076 9098
rect 2885 9059 3036 9082
rect 2885 9025 2891 9059
rect 2925 9048 3036 9059
rect 3070 9048 3076 9082
rect 2925 9025 3076 9048
rect 2885 9010 3076 9025
rect 2885 8986 3036 9010
rect 2885 8952 2891 8986
rect 2925 8976 3036 8986
rect 3070 8976 3076 9010
rect 2925 8952 3076 8976
rect 2885 8938 3076 8952
rect 2885 8913 3036 8938
rect 2885 8879 2891 8913
rect 2925 8904 3036 8913
rect 3070 8904 3076 8938
rect 2925 8879 3076 8904
rect 2885 8866 3076 8879
rect 2885 8840 3036 8866
rect 2885 8806 2891 8840
rect 2925 8832 3036 8840
rect 3070 8832 3076 8866
rect 2925 8806 3076 8832
rect 2885 8794 3076 8806
rect 2885 8767 3036 8794
rect 2885 8733 2891 8767
rect 2925 8760 3036 8767
rect 3070 8760 3076 8794
rect 2925 8733 3076 8760
rect 2885 8722 3076 8733
rect 2885 8694 3036 8722
tri 2695 8660 2707 8672 sw
tri 2873 8660 2885 8672 se
rect 2885 8660 2891 8694
rect 2925 8688 3036 8694
rect 3070 8688 3076 8722
rect 2925 8660 3076 8688
rect 380 8650 583 8660
tri 583 8650 593 8660 sw
tri 739 8650 749 8660 se
rect 749 8650 819 8660
tri 819 8650 829 8660 sw
tri 975 8650 985 8660 se
rect 985 8650 1055 8660
tri 1055 8650 1065 8660 sw
tri 1211 8650 1221 8660 se
rect 1221 8650 1291 8660
tri 1291 8650 1301 8660 sw
tri 1447 8650 1457 8660 se
rect 1457 8650 1527 8660
tri 1527 8650 1537 8660 sw
tri 1683 8650 1693 8660 se
rect 1693 8650 1763 8660
tri 1763 8650 1773 8660 sw
tri 1919 8650 1929 8660 se
rect 1929 8650 1999 8660
tri 1999 8650 2009 8660 sw
tri 2155 8650 2165 8660 se
rect 2165 8650 2235 8660
tri 2235 8650 2245 8660 sw
tri 2391 8650 2401 8660 se
rect 2401 8650 2471 8660
tri 2471 8650 2481 8660 sw
tri 2627 8650 2637 8660 se
rect 2637 8650 2707 8660
tri 2707 8650 2717 8660 sw
tri 2863 8650 2873 8660 se
rect 2873 8650 3076 8660
rect 380 8638 593 8650
tri 593 8638 605 8650 sw
tri 727 8638 739 8650 se
rect 739 8638 829 8650
tri 829 8638 841 8650 sw
tri 963 8638 975 8650 se
rect 975 8638 1065 8650
tri 1065 8638 1077 8650 sw
tri 1199 8638 1211 8650 se
rect 1211 8638 1301 8650
tri 1301 8638 1313 8650 sw
tri 1435 8638 1447 8650 se
rect 1447 8638 1537 8650
tri 1537 8638 1549 8650 sw
tri 1671 8638 1683 8650 se
rect 1683 8638 1773 8650
tri 1773 8638 1785 8650 sw
tri 1907 8638 1919 8650 se
rect 1919 8638 2009 8650
tri 2009 8638 2021 8650 sw
tri 2143 8638 2155 8650 se
rect 2155 8638 2245 8650
tri 2245 8638 2257 8650 sw
tri 2379 8638 2391 8650 se
rect 2391 8638 2481 8650
tri 2481 8638 2493 8650 sw
tri 2615 8638 2627 8650 se
rect 2627 8638 2717 8650
tri 2717 8638 2729 8650 sw
tri 2851 8638 2863 8650 se
rect 2863 8638 3036 8650
rect 380 8631 3036 8638
rect 380 8597 386 8631
rect 420 8621 3036 8631
rect 420 8597 531 8621
rect 380 8587 531 8597
rect 565 8611 767 8621
rect 801 8611 1003 8621
rect 1037 8611 1239 8621
rect 1273 8611 1475 8621
rect 565 8587 697 8611
rect 380 8559 697 8587
rect 749 8559 765 8611
rect 817 8559 833 8611
rect 885 8559 901 8611
rect 953 8559 969 8611
rect 1021 8559 1037 8587
rect 1089 8559 1105 8611
rect 1157 8559 1173 8611
rect 1225 8587 1239 8611
rect 1293 8587 1475 8611
rect 1509 8587 1711 8621
rect 1745 8587 1947 8621
rect 1981 8611 2183 8621
rect 2217 8611 2419 8621
rect 2453 8611 2655 8621
rect 2689 8611 2891 8621
rect 1981 8587 2097 8611
rect 1225 8559 1241 8587
rect 1293 8559 2097 8587
rect 2149 8559 2165 8611
rect 2217 8559 2233 8611
rect 2285 8559 2301 8611
rect 2353 8559 2369 8611
rect 2421 8559 2437 8587
rect 2489 8559 2505 8611
rect 2557 8559 2573 8611
rect 2625 8559 2641 8611
rect 2693 8587 2891 8611
rect 2925 8616 3036 8621
rect 3070 8616 3076 8650
rect 2925 8587 3076 8616
rect 2693 8578 3076 8587
rect 2693 8559 3036 8578
rect 380 8525 386 8559
rect 420 8548 3036 8559
rect 420 8525 531 8548
rect 380 8514 531 8525
rect 565 8547 767 8548
rect 801 8547 1003 8548
rect 1037 8547 1239 8548
rect 1273 8547 1475 8548
rect 565 8514 697 8547
rect 380 8495 697 8514
rect 749 8495 765 8547
rect 817 8495 833 8547
rect 885 8495 901 8547
rect 953 8495 969 8547
rect 1021 8495 1037 8514
rect 1089 8495 1105 8547
rect 1157 8495 1173 8547
rect 1225 8514 1239 8547
rect 1293 8514 1475 8547
rect 1509 8514 1711 8548
rect 1745 8514 1947 8548
rect 1981 8547 2183 8548
rect 2217 8547 2419 8548
rect 2453 8547 2655 8548
rect 2689 8547 2891 8548
rect 1981 8514 2097 8547
rect 1225 8495 1241 8514
rect 1293 8495 2097 8514
rect 2149 8495 2165 8547
rect 2217 8495 2233 8547
rect 2285 8495 2301 8547
rect 2353 8495 2369 8547
rect 2421 8495 2437 8514
rect 2489 8495 2505 8547
rect 2557 8495 2573 8547
rect 2625 8495 2641 8547
rect 2693 8514 2891 8547
rect 2925 8544 3036 8548
rect 3070 8544 3076 8578
rect 2925 8514 3076 8544
rect 2693 8506 3076 8514
rect 2693 8495 3036 8506
rect 380 8487 3036 8495
rect 380 8453 386 8487
rect 420 8483 3036 8487
rect 420 8475 697 8483
rect 420 8453 531 8475
rect 380 8441 531 8453
rect 565 8441 697 8475
rect 380 8431 697 8441
rect 749 8431 765 8483
rect 817 8431 833 8483
rect 885 8431 901 8483
rect 953 8431 969 8483
rect 1021 8475 1037 8483
rect 1021 8431 1037 8441
rect 1089 8431 1105 8483
rect 1157 8431 1173 8483
rect 1225 8475 1241 8483
rect 1293 8475 2097 8483
rect 1225 8441 1239 8475
rect 1293 8441 1475 8475
rect 1509 8441 1711 8475
rect 1745 8441 1947 8475
rect 1981 8441 2097 8475
rect 1225 8431 1241 8441
rect 1293 8431 2097 8441
rect 2149 8431 2165 8483
rect 2217 8431 2233 8483
rect 2285 8431 2301 8483
rect 2353 8431 2369 8483
rect 2421 8475 2437 8483
rect 2421 8431 2437 8441
rect 2489 8431 2505 8483
rect 2557 8431 2573 8483
rect 2625 8431 2641 8483
rect 2693 8475 3036 8483
rect 2693 8441 2891 8475
rect 2925 8472 3036 8475
rect 3070 8472 3076 8506
rect 2925 8441 3076 8472
rect 2693 8434 3076 8441
rect 2693 8431 3036 8434
rect 380 8419 3036 8431
rect 380 8415 697 8419
rect 380 8381 386 8415
rect 420 8402 697 8415
rect 420 8381 531 8402
rect 380 8368 531 8381
rect 565 8368 697 8402
rect 380 8367 697 8368
rect 749 8367 765 8419
rect 817 8367 833 8419
rect 885 8367 901 8419
rect 953 8367 969 8419
rect 1021 8402 1037 8419
rect 1021 8367 1037 8368
rect 1089 8367 1105 8419
rect 1157 8367 1173 8419
rect 1225 8402 1241 8419
rect 1293 8402 2097 8419
rect 1225 8368 1239 8402
rect 1293 8368 1475 8402
rect 1509 8368 1711 8402
rect 1745 8368 1947 8402
rect 1981 8368 2097 8402
rect 1225 8367 1241 8368
rect 1293 8367 2097 8368
rect 2149 8367 2165 8419
rect 2217 8367 2233 8419
rect 2285 8367 2301 8419
rect 2353 8367 2369 8419
rect 2421 8402 2437 8419
rect 2421 8367 2437 8368
rect 2489 8367 2505 8419
rect 2557 8367 2573 8419
rect 2625 8367 2641 8419
rect 2693 8402 3036 8419
rect 2693 8368 2891 8402
rect 2925 8400 3036 8402
rect 3070 8400 3076 8434
rect 2925 8368 3076 8400
rect 2693 8367 3076 8368
rect 380 8362 3076 8367
rect 380 8355 3036 8362
rect 380 8343 697 8355
rect 380 8309 386 8343
rect 420 8329 697 8343
rect 420 8309 531 8329
rect 380 8295 531 8309
rect 565 8303 697 8329
rect 749 8303 765 8355
rect 817 8303 833 8355
rect 885 8303 901 8355
rect 953 8303 969 8355
rect 1021 8329 1037 8355
rect 1089 8303 1105 8355
rect 1157 8303 1173 8355
rect 1225 8329 1241 8355
rect 1293 8329 2097 8355
rect 1225 8303 1239 8329
rect 1293 8303 1475 8329
rect 565 8295 767 8303
rect 801 8295 1003 8303
rect 1037 8295 1239 8303
rect 1273 8295 1475 8303
rect 1509 8295 1711 8329
rect 1745 8295 1947 8329
rect 1981 8303 2097 8329
rect 2149 8303 2165 8355
rect 2217 8303 2233 8355
rect 2285 8303 2301 8355
rect 2353 8303 2369 8355
rect 2421 8329 2437 8355
rect 2489 8303 2505 8355
rect 2557 8303 2573 8355
rect 2625 8303 2641 8355
rect 2693 8329 3036 8355
rect 2693 8303 2891 8329
rect 1981 8295 2183 8303
rect 2217 8295 2419 8303
rect 2453 8295 2655 8303
rect 2689 8295 2891 8303
rect 2925 8328 3036 8329
rect 3070 8328 3076 8362
rect 2925 8295 3076 8328
rect 380 8291 3076 8295
rect 380 8271 697 8291
rect 380 8237 386 8271
rect 420 8256 697 8271
rect 420 8237 531 8256
rect 380 8222 531 8237
rect 565 8239 697 8256
rect 749 8239 765 8291
rect 817 8239 833 8291
rect 885 8239 901 8291
rect 953 8239 969 8291
rect 1021 8256 1037 8291
rect 1089 8239 1105 8291
rect 1157 8239 1173 8291
rect 1225 8256 1241 8291
rect 1293 8256 2097 8291
rect 1225 8239 1239 8256
rect 1293 8239 1475 8256
rect 565 8227 767 8239
rect 801 8227 1003 8239
rect 1037 8227 1239 8239
rect 1273 8227 1475 8239
rect 565 8222 697 8227
rect 380 8199 697 8222
rect 380 8165 386 8199
rect 420 8182 697 8199
rect 420 8165 531 8182
rect 380 8148 531 8165
rect 565 8175 697 8182
rect 749 8175 765 8227
rect 817 8175 833 8227
rect 885 8175 901 8227
rect 953 8175 969 8227
rect 1021 8182 1037 8222
rect 1089 8175 1105 8227
rect 1157 8175 1173 8227
rect 1225 8222 1239 8227
rect 1293 8222 1475 8227
rect 1509 8222 1711 8256
rect 1745 8222 1947 8256
rect 1981 8239 2097 8256
rect 2149 8239 2165 8291
rect 2217 8239 2233 8291
rect 2285 8239 2301 8291
rect 2353 8239 2369 8291
rect 2421 8256 2437 8291
rect 2489 8239 2505 8291
rect 2557 8239 2573 8291
rect 2625 8239 2641 8291
rect 2693 8290 3076 8291
rect 2693 8256 3036 8290
rect 3070 8256 3076 8290
rect 2693 8239 2891 8256
rect 1981 8227 2183 8239
rect 2217 8227 2419 8239
rect 2453 8227 2655 8239
rect 2689 8227 2891 8239
rect 1981 8222 2097 8227
rect 1225 8182 1241 8222
rect 1293 8182 2097 8222
rect 1225 8175 1239 8182
rect 1293 8175 1475 8182
rect 565 8163 767 8175
rect 801 8163 1003 8175
rect 1037 8163 1239 8175
rect 1273 8163 1475 8175
rect 565 8148 697 8163
rect 380 8127 697 8148
rect 380 8093 386 8127
rect 420 8111 697 8127
rect 749 8111 765 8163
rect 817 8111 833 8163
rect 885 8111 901 8163
rect 953 8111 969 8163
rect 1021 8111 1037 8148
rect 1089 8111 1105 8163
rect 1157 8111 1173 8163
rect 1225 8148 1239 8163
rect 1293 8148 1475 8163
rect 1509 8148 1711 8182
rect 1745 8148 1947 8182
rect 1981 8175 2097 8182
rect 2149 8175 2165 8227
rect 2217 8175 2233 8227
rect 2285 8175 2301 8227
rect 2353 8175 2369 8227
rect 2421 8182 2437 8222
rect 2489 8175 2505 8227
rect 2557 8175 2573 8227
rect 2625 8175 2641 8227
rect 2693 8222 2891 8227
rect 2925 8222 3076 8256
rect 2693 8218 3076 8222
rect 2693 8184 3036 8218
rect 3070 8184 3076 8218
rect 2693 8182 3076 8184
rect 2693 8175 2891 8182
rect 1981 8163 2183 8175
rect 2217 8163 2419 8175
rect 2453 8163 2655 8175
rect 2689 8163 2891 8175
rect 1981 8148 2097 8163
rect 1225 8111 1241 8148
rect 1293 8111 2097 8148
rect 2149 8111 2165 8163
rect 2217 8111 2233 8163
rect 2285 8111 2301 8163
rect 2353 8111 2369 8163
rect 2421 8111 2437 8148
rect 2489 8111 2505 8163
rect 2557 8111 2573 8163
rect 2625 8111 2641 8163
rect 2693 8148 2891 8163
rect 2925 8148 3076 8182
rect 2693 8146 3076 8148
rect 2693 8112 3036 8146
rect 3070 8112 3076 8146
rect 2693 8111 3076 8112
rect 420 8108 3076 8111
rect 420 8093 531 8108
rect 380 8074 531 8093
rect 565 8099 767 8108
rect 801 8099 1003 8108
rect 1037 8099 1239 8108
rect 1273 8099 1475 8108
rect 565 8074 697 8099
rect 380 8055 697 8074
rect 380 8021 386 8055
rect 420 8047 697 8055
rect 749 8047 765 8099
rect 817 8047 833 8099
rect 885 8047 901 8099
rect 953 8047 969 8099
rect 1021 8047 1037 8074
rect 1089 8047 1105 8099
rect 1157 8047 1173 8099
rect 1225 8074 1239 8099
rect 1293 8074 1475 8099
rect 1509 8074 1711 8108
rect 1745 8074 1947 8108
rect 1981 8099 2183 8108
rect 2217 8099 2419 8108
rect 2453 8099 2655 8108
rect 2689 8099 2891 8108
rect 1981 8074 2097 8099
rect 1225 8047 1241 8074
rect 1293 8047 2097 8074
rect 2149 8047 2165 8099
rect 2217 8047 2233 8099
rect 2285 8047 2301 8099
rect 2353 8047 2369 8099
rect 2421 8047 2437 8074
rect 2489 8047 2505 8099
rect 2557 8047 2573 8099
rect 2625 8047 2641 8099
rect 2693 8074 2891 8099
rect 2925 8074 3076 8108
rect 2693 8047 3036 8074
rect 420 8040 3036 8047
rect 3070 8040 3076 8074
rect 420 8035 3076 8040
rect 420 8034 697 8035
rect 420 8021 531 8034
rect 380 8000 531 8021
rect 565 8000 697 8034
rect 380 7983 697 8000
rect 749 7983 765 8035
rect 817 7983 833 8035
rect 885 7983 901 8035
rect 953 7983 969 8035
rect 1021 8034 1037 8035
rect 1021 7983 1037 8000
rect 1089 7983 1105 8035
rect 1157 7983 1173 8035
rect 1225 8034 1241 8035
rect 1293 8034 2097 8035
rect 1225 8000 1239 8034
rect 1293 8000 1475 8034
rect 1509 8000 1711 8034
rect 1745 8000 1947 8034
rect 1981 8000 2097 8034
rect 1225 7983 1241 8000
rect 1293 7983 2097 8000
rect 2149 7983 2165 8035
rect 2217 7983 2233 8035
rect 2285 7983 2301 8035
rect 2353 7983 2369 8035
rect 2421 8034 2437 8035
rect 2421 7983 2437 8000
rect 2489 7983 2505 8035
rect 2557 7983 2573 8035
rect 2625 7983 2641 8035
rect 2693 8034 3076 8035
rect 2693 8000 2891 8034
rect 2925 8002 3076 8034
rect 2925 8000 3036 8002
rect 2693 7983 3036 8000
rect 380 7949 386 7983
rect 420 7971 3036 7983
rect 420 7960 697 7971
rect 420 7949 531 7960
rect 380 7926 531 7949
rect 565 7926 697 7960
rect 380 7919 697 7926
rect 749 7919 765 7971
rect 817 7919 833 7971
rect 885 7919 901 7971
rect 953 7919 969 7971
rect 1021 7960 1037 7971
rect 1021 7919 1037 7926
rect 1089 7919 1105 7971
rect 1157 7919 1173 7971
rect 1225 7960 1241 7971
rect 1293 7960 2097 7971
rect 1225 7926 1239 7960
rect 1293 7926 1475 7960
rect 1509 7926 1711 7960
rect 1745 7926 1947 7960
rect 1981 7926 2097 7960
rect 1225 7919 1241 7926
rect 1293 7919 2097 7926
rect 2149 7919 2165 7971
rect 2217 7919 2233 7971
rect 2285 7919 2301 7971
rect 2353 7919 2369 7971
rect 2421 7960 2437 7971
rect 2421 7919 2437 7926
rect 2489 7919 2505 7971
rect 2557 7919 2573 7971
rect 2625 7919 2641 7971
rect 2693 7968 3036 7971
rect 3070 7968 3076 8002
rect 2693 7960 3076 7968
rect 2693 7926 2891 7960
rect 2925 7930 3076 7960
rect 2925 7926 3036 7930
rect 2693 7919 3036 7926
rect 380 7911 3036 7919
rect 380 7877 386 7911
rect 420 7907 3036 7911
rect 420 7886 697 7907
rect 420 7877 531 7886
rect 380 7852 531 7877
rect 565 7855 697 7886
rect 749 7855 765 7907
rect 817 7855 833 7907
rect 885 7855 901 7907
rect 953 7855 969 7907
rect 1021 7886 1037 7907
rect 1089 7855 1105 7907
rect 1157 7855 1173 7907
rect 1225 7886 1241 7907
rect 1293 7886 2097 7907
rect 1225 7855 1239 7886
rect 1293 7855 1475 7886
rect 565 7852 767 7855
rect 801 7852 1003 7855
rect 1037 7852 1239 7855
rect 1273 7852 1475 7855
rect 1509 7852 1711 7886
rect 1745 7852 1947 7886
rect 1981 7855 2097 7886
rect 2149 7855 2165 7907
rect 2217 7855 2233 7907
rect 2285 7855 2301 7907
rect 2353 7855 2369 7907
rect 2421 7886 2437 7907
rect 2489 7855 2505 7907
rect 2557 7855 2573 7907
rect 2625 7855 2641 7907
rect 2693 7896 3036 7907
rect 3070 7896 3076 7930
rect 2693 7886 3076 7896
rect 2693 7855 2891 7886
rect 1981 7852 2183 7855
rect 2217 7852 2419 7855
rect 2453 7852 2655 7855
rect 2689 7852 2891 7855
rect 2925 7858 3076 7886
rect 2925 7852 3036 7858
rect 380 7843 3036 7852
rect 380 7839 697 7843
rect 380 7805 386 7839
rect 420 7812 697 7839
rect 420 7805 531 7812
rect 380 7778 531 7805
rect 565 7791 697 7812
rect 749 7791 765 7843
rect 817 7791 833 7843
rect 885 7791 901 7843
rect 953 7791 969 7843
rect 1021 7812 1037 7843
rect 1089 7791 1105 7843
rect 1157 7791 1173 7843
rect 1225 7812 1241 7843
rect 1293 7812 2097 7843
rect 1225 7791 1239 7812
rect 1293 7791 1475 7812
rect 565 7779 767 7791
rect 801 7779 1003 7791
rect 1037 7779 1239 7791
rect 1273 7779 1475 7791
rect 565 7778 697 7779
rect 380 7767 697 7778
rect 380 7733 386 7767
rect 420 7738 697 7767
rect 420 7733 531 7738
rect 380 7704 531 7733
rect 565 7727 697 7738
rect 749 7727 765 7779
rect 817 7727 833 7779
rect 885 7727 901 7779
rect 953 7727 969 7779
rect 1021 7738 1037 7778
rect 1089 7727 1105 7779
rect 1157 7727 1173 7779
rect 1225 7778 1239 7779
rect 1293 7778 1475 7779
rect 1509 7778 1711 7812
rect 1745 7778 1947 7812
rect 1981 7791 2097 7812
rect 2149 7791 2165 7843
rect 2217 7791 2233 7843
rect 2285 7791 2301 7843
rect 2353 7791 2369 7843
rect 2421 7812 2437 7843
rect 2489 7791 2505 7843
rect 2557 7791 2573 7843
rect 2625 7791 2641 7843
rect 2693 7824 3036 7843
rect 3070 7824 3076 7858
rect 2693 7812 3076 7824
rect 2693 7791 2891 7812
rect 1981 7779 2183 7791
rect 2217 7779 2419 7791
rect 2453 7779 2655 7791
rect 2689 7779 2891 7791
rect 1981 7778 2097 7779
rect 1225 7738 1241 7778
rect 1293 7738 2097 7778
rect 1225 7727 1239 7738
rect 1293 7727 1475 7738
rect 565 7715 767 7727
rect 801 7715 1003 7727
rect 1037 7715 1239 7727
rect 1273 7715 1475 7727
rect 565 7704 697 7715
rect 380 7695 697 7704
rect 380 7661 386 7695
rect 420 7664 697 7695
rect 420 7661 531 7664
rect 380 7630 531 7661
rect 565 7663 697 7664
rect 749 7663 765 7715
rect 817 7663 833 7715
rect 885 7663 901 7715
rect 953 7663 969 7715
rect 1021 7664 1037 7704
rect 1089 7663 1105 7715
rect 1157 7663 1173 7715
rect 1225 7704 1239 7715
rect 1293 7704 1475 7715
rect 1509 7704 1711 7738
rect 1745 7704 1947 7738
rect 1981 7727 2097 7738
rect 2149 7727 2165 7779
rect 2217 7727 2233 7779
rect 2285 7727 2301 7779
rect 2353 7727 2369 7779
rect 2421 7738 2437 7778
rect 2489 7727 2505 7779
rect 2557 7727 2573 7779
rect 2625 7727 2641 7779
rect 2693 7778 2891 7779
rect 2925 7786 3076 7812
rect 2925 7778 3036 7786
rect 2693 7752 3036 7778
rect 3070 7752 3076 7786
rect 2693 7738 3076 7752
rect 2693 7727 2891 7738
rect 1981 7715 2183 7727
rect 2217 7715 2419 7727
rect 2453 7715 2655 7727
rect 2689 7715 2891 7727
rect 1981 7704 2097 7715
rect 1225 7664 1241 7704
rect 1293 7664 2097 7704
rect 1225 7663 1239 7664
rect 1293 7663 1475 7664
rect 565 7638 767 7663
rect 565 7630 597 7638
tri 597 7630 605 7638 nw
tri 727 7630 735 7638 ne
rect 735 7630 767 7638
rect 801 7638 1003 7663
rect 801 7630 833 7638
tri 833 7630 841 7638 nw
tri 963 7630 971 7638 ne
rect 971 7630 1003 7638
rect 1037 7638 1239 7663
rect 1037 7630 1069 7638
tri 1069 7630 1077 7638 nw
tri 1199 7630 1207 7638 ne
rect 1207 7630 1239 7638
rect 1273 7638 1475 7663
rect 1273 7630 1305 7638
tri 1305 7630 1313 7638 nw
tri 1435 7630 1443 7638 ne
rect 1443 7630 1475 7638
rect 1509 7638 1711 7664
rect 1509 7630 1541 7638
tri 1541 7630 1549 7638 nw
tri 1671 7630 1679 7638 ne
rect 1679 7630 1711 7638
rect 1745 7638 1947 7664
rect 1745 7630 1777 7638
tri 1777 7630 1785 7638 nw
tri 1907 7630 1915 7638 ne
rect 1915 7630 1947 7638
rect 1981 7663 2097 7664
rect 2149 7663 2165 7715
rect 2217 7663 2233 7715
rect 2285 7663 2301 7715
rect 2353 7663 2369 7715
rect 2421 7664 2437 7704
rect 2489 7663 2505 7715
rect 2557 7663 2573 7715
rect 2625 7663 2641 7715
rect 2693 7704 2891 7715
rect 2925 7714 3076 7738
rect 2925 7704 3036 7714
rect 2693 7680 3036 7704
rect 3070 7680 3076 7714
rect 2693 7664 3076 7680
rect 2693 7663 2891 7664
rect 1981 7638 2183 7663
rect 1981 7630 2013 7638
tri 2013 7630 2021 7638 nw
tri 2143 7630 2151 7638 ne
rect 2151 7630 2183 7638
rect 2217 7638 2419 7663
rect 2217 7630 2249 7638
tri 2249 7630 2257 7638 nw
tri 2379 7630 2387 7638 ne
rect 2387 7630 2419 7638
rect 2453 7638 2655 7663
rect 2453 7630 2485 7638
tri 2485 7630 2493 7638 nw
tri 2615 7630 2623 7638 ne
rect 2623 7630 2655 7638
rect 2689 7638 2891 7663
rect 2689 7630 2721 7638
tri 2721 7630 2729 7638 nw
tri 2851 7630 2859 7638 ne
rect 2859 7630 2891 7638
rect 2925 7642 3076 7664
rect 2925 7630 3036 7642
rect 380 7623 575 7630
rect 380 7589 386 7623
rect 420 7608 575 7623
tri 575 7608 597 7630 nw
tri 735 7608 757 7630 ne
rect 757 7608 811 7630
tri 811 7608 833 7630 nw
tri 971 7608 993 7630 ne
rect 993 7608 1047 7630
tri 1047 7608 1069 7630 nw
tri 1207 7608 1229 7630 ne
rect 1229 7608 1283 7630
tri 1283 7608 1305 7630 nw
tri 1443 7608 1465 7630 ne
rect 1465 7608 1519 7630
tri 1519 7608 1541 7630 nw
tri 1679 7608 1701 7630 ne
rect 1701 7608 1755 7630
tri 1755 7608 1777 7630 nw
tri 1915 7608 1937 7630 ne
rect 1937 7608 1991 7630
tri 1991 7608 2013 7630 nw
tri 2151 7608 2173 7630 ne
rect 2173 7608 2227 7630
tri 2227 7608 2249 7630 nw
tri 2387 7608 2409 7630 ne
rect 2409 7608 2463 7630
tri 2463 7608 2485 7630 nw
tri 2623 7608 2645 7630 ne
rect 2645 7608 2699 7630
tri 2699 7608 2721 7630 nw
tri 2859 7608 2881 7630 ne
rect 2881 7608 3036 7630
rect 3070 7608 3076 7642
rect 420 7590 571 7608
tri 571 7604 575 7608 nw
tri 757 7604 761 7608 ne
rect 420 7589 531 7590
rect 380 7556 531 7589
rect 565 7556 571 7590
rect 380 7551 571 7556
rect 380 7517 386 7551
rect 420 7517 571 7551
rect 380 7516 571 7517
rect 380 7482 531 7516
rect 565 7482 571 7516
rect 380 7479 571 7482
rect 380 7445 386 7479
rect 420 7445 571 7479
rect 380 7442 571 7445
rect 380 7408 531 7442
rect 565 7408 571 7442
rect 380 7407 571 7408
rect 380 7373 386 7407
rect 420 7373 571 7407
rect 380 7368 571 7373
rect 380 7335 531 7368
rect 380 7301 386 7335
rect 420 7334 531 7335
rect 565 7334 571 7368
rect 420 7301 571 7334
rect 380 7294 571 7301
rect 380 7263 531 7294
rect 380 7229 386 7263
rect 420 7260 531 7263
rect 565 7260 571 7294
rect 420 7229 571 7260
rect 380 7220 571 7229
rect 380 7191 531 7220
rect 380 7157 386 7191
rect 420 7186 531 7191
rect 565 7186 571 7220
rect 420 7157 571 7186
rect 761 7590 807 7608
tri 807 7604 811 7608 nw
tri 993 7604 997 7608 ne
rect 761 7556 767 7590
rect 801 7556 807 7590
rect 761 7516 807 7556
rect 761 7482 767 7516
rect 801 7482 807 7516
rect 761 7442 807 7482
rect 761 7408 767 7442
rect 801 7408 807 7442
rect 761 7368 807 7408
rect 761 7334 767 7368
rect 801 7334 807 7368
rect 761 7294 807 7334
rect 761 7260 767 7294
rect 801 7260 807 7294
rect 761 7220 807 7260
rect 761 7186 767 7220
rect 801 7186 807 7220
rect 761 7174 807 7186
rect 997 7590 1043 7608
tri 1043 7604 1047 7608 nw
tri 1229 7604 1233 7608 ne
rect 997 7556 1003 7590
rect 1037 7556 1043 7590
rect 997 7516 1043 7556
rect 997 7482 1003 7516
rect 1037 7482 1043 7516
rect 997 7442 1043 7482
rect 997 7408 1003 7442
rect 1037 7408 1043 7442
rect 997 7368 1043 7408
rect 997 7334 1003 7368
rect 1037 7334 1043 7368
rect 997 7294 1043 7334
rect 997 7260 1003 7294
rect 1037 7260 1043 7294
rect 997 7220 1043 7260
rect 997 7186 1003 7220
rect 1037 7186 1043 7220
rect 997 7174 1043 7186
rect 1233 7590 1279 7608
tri 1279 7604 1283 7608 nw
tri 1465 7604 1469 7608 ne
rect 1233 7556 1239 7590
rect 1273 7556 1279 7590
rect 1233 7516 1279 7556
rect 1233 7482 1239 7516
rect 1273 7482 1279 7516
rect 1233 7442 1279 7482
rect 1233 7408 1239 7442
rect 1273 7408 1279 7442
rect 1233 7368 1279 7408
rect 1233 7334 1239 7368
rect 1273 7334 1279 7368
rect 1233 7294 1279 7334
rect 1233 7260 1239 7294
rect 1273 7260 1279 7294
rect 1233 7220 1279 7260
rect 1233 7186 1239 7220
rect 1273 7186 1279 7220
rect 1233 7174 1279 7186
rect 1469 7590 1515 7608
tri 1515 7604 1519 7608 nw
tri 1701 7604 1705 7608 ne
rect 1469 7556 1475 7590
rect 1509 7556 1515 7590
rect 1469 7516 1515 7556
rect 1469 7482 1475 7516
rect 1509 7482 1515 7516
rect 1469 7442 1515 7482
rect 1469 7408 1475 7442
rect 1509 7408 1515 7442
rect 1469 7368 1515 7408
rect 1469 7334 1475 7368
rect 1509 7334 1515 7368
rect 1469 7294 1515 7334
rect 1469 7260 1475 7294
rect 1509 7260 1515 7294
rect 1469 7220 1515 7260
rect 1469 7186 1475 7220
rect 1509 7186 1515 7220
rect 1469 7174 1515 7186
rect 1705 7590 1751 7608
tri 1751 7604 1755 7608 nw
tri 1937 7604 1941 7608 ne
rect 1705 7556 1711 7590
rect 1745 7556 1751 7590
rect 1705 7516 1751 7556
rect 1705 7482 1711 7516
rect 1745 7482 1751 7516
rect 1705 7442 1751 7482
rect 1705 7408 1711 7442
rect 1745 7408 1751 7442
rect 1705 7368 1751 7408
rect 1705 7334 1711 7368
rect 1745 7334 1751 7368
rect 1705 7294 1751 7334
rect 1705 7260 1711 7294
rect 1745 7260 1751 7294
rect 1705 7220 1751 7260
rect 1705 7186 1711 7220
rect 1745 7186 1751 7220
rect 1705 7174 1751 7186
rect 1941 7590 1987 7608
tri 1987 7604 1991 7608 nw
tri 2173 7604 2177 7608 ne
rect 1941 7556 1947 7590
rect 1981 7556 1987 7590
rect 1941 7516 1987 7556
rect 1941 7482 1947 7516
rect 1981 7482 1987 7516
rect 1941 7442 1987 7482
rect 1941 7408 1947 7442
rect 1981 7408 1987 7442
rect 1941 7368 1987 7408
rect 1941 7334 1947 7368
rect 1981 7334 1987 7368
rect 1941 7294 1987 7334
rect 1941 7260 1947 7294
rect 1981 7260 1987 7294
rect 1941 7220 1987 7260
rect 1941 7186 1947 7220
rect 1981 7186 1987 7220
rect 1941 7174 1987 7186
rect 2177 7590 2223 7608
tri 2223 7604 2227 7608 nw
tri 2409 7604 2413 7608 ne
rect 2177 7556 2183 7590
rect 2217 7556 2223 7590
rect 2177 7516 2223 7556
rect 2177 7482 2183 7516
rect 2217 7482 2223 7516
rect 2177 7442 2223 7482
rect 2177 7408 2183 7442
rect 2217 7408 2223 7442
rect 2177 7368 2223 7408
rect 2177 7334 2183 7368
rect 2217 7334 2223 7368
rect 2177 7294 2223 7334
rect 2177 7260 2183 7294
rect 2217 7260 2223 7294
rect 2177 7220 2223 7260
rect 2177 7186 2183 7220
rect 2217 7186 2223 7220
rect 2177 7174 2223 7186
rect 2413 7590 2459 7608
tri 2459 7604 2463 7608 nw
tri 2645 7604 2649 7608 ne
rect 2413 7556 2419 7590
rect 2453 7556 2459 7590
rect 2413 7516 2459 7556
rect 2413 7482 2419 7516
rect 2453 7482 2459 7516
rect 2413 7442 2459 7482
rect 2413 7408 2419 7442
rect 2453 7408 2459 7442
rect 2413 7368 2459 7408
rect 2413 7334 2419 7368
rect 2453 7334 2459 7368
rect 2413 7294 2459 7334
rect 2413 7260 2419 7294
rect 2453 7260 2459 7294
rect 2413 7220 2459 7260
rect 2413 7186 2419 7220
rect 2453 7186 2459 7220
rect 2413 7174 2459 7186
rect 2649 7590 2695 7608
tri 2695 7604 2699 7608 nw
tri 2881 7604 2885 7608 ne
rect 2649 7556 2655 7590
rect 2689 7556 2695 7590
rect 2649 7516 2695 7556
rect 2649 7482 2655 7516
rect 2689 7482 2695 7516
rect 2649 7442 2695 7482
rect 2649 7408 2655 7442
rect 2689 7408 2695 7442
rect 2649 7368 2695 7408
rect 2649 7334 2655 7368
rect 2689 7334 2695 7368
rect 2649 7294 2695 7334
rect 2649 7260 2655 7294
rect 2689 7260 2695 7294
rect 2649 7220 2695 7260
rect 2649 7186 2655 7220
rect 2689 7186 2695 7220
rect 2649 7174 2695 7186
rect 2885 7590 3076 7608
rect 2885 7556 2891 7590
rect 2925 7570 3076 7590
rect 2925 7556 3036 7570
rect 2885 7536 3036 7556
rect 3070 7536 3076 7570
rect 2885 7516 3076 7536
rect 2885 7482 2891 7516
rect 2925 7498 3076 7516
rect 2925 7482 3036 7498
rect 2885 7464 3036 7482
rect 3070 7464 3076 7498
rect 2885 7442 3076 7464
rect 2885 7408 2891 7442
rect 2925 7426 3076 7442
rect 2925 7408 3036 7426
rect 2885 7392 3036 7408
rect 3070 7392 3076 7426
rect 2885 7368 3076 7392
rect 2885 7334 2891 7368
rect 2925 7354 3076 7368
rect 2925 7334 3036 7354
rect 2885 7320 3036 7334
rect 3070 7320 3076 7354
rect 2885 7294 3076 7320
rect 2885 7260 2891 7294
rect 2925 7282 3076 7294
rect 2925 7260 3036 7282
rect 2885 7248 3036 7260
rect 3070 7248 3076 7282
rect 2885 7220 3076 7248
rect 2885 7186 2891 7220
rect 2925 7210 3076 7220
rect 2925 7186 3036 7210
rect 2885 7176 3036 7186
rect 3070 7176 3076 7210
rect 380 7119 571 7157
rect 380 7085 386 7119
rect 420 7085 571 7119
rect 2885 7138 3076 7176
rect 380 7047 571 7085
rect 613 7104 1501 7113
rect 1553 7104 1569 7113
rect 1621 7104 1636 7113
rect 1688 7104 1703 7113
rect 1755 7104 1770 7113
rect 1822 7104 1837 7113
rect 1889 7104 2830 7113
rect 613 7070 625 7104
rect 659 7070 700 7104
rect 734 7070 775 7104
rect 809 7070 850 7104
rect 884 7070 925 7104
rect 959 7070 1000 7104
rect 1034 7070 1075 7104
rect 1109 7070 1150 7104
rect 1184 7070 1225 7104
rect 1259 7070 1300 7104
rect 1334 7070 1375 7104
rect 1409 7070 1450 7104
rect 1484 7070 1501 7104
rect 1559 7070 1569 7104
rect 1634 7070 1636 7104
rect 1889 7070 1896 7104
rect 1930 7070 1970 7104
rect 2004 7070 2044 7104
rect 2078 7070 2118 7104
rect 2152 7070 2192 7104
rect 2226 7070 2266 7104
rect 2300 7070 2340 7104
rect 2374 7070 2414 7104
rect 2448 7070 2488 7104
rect 2522 7070 2562 7104
rect 2596 7070 2636 7104
rect 2670 7070 2710 7104
rect 2744 7070 2784 7104
rect 2818 7070 2830 7104
rect 613 7061 1501 7070
rect 1553 7061 1569 7070
rect 1621 7061 1636 7070
rect 1688 7061 1703 7070
rect 1755 7061 1770 7070
rect 1822 7061 1837 7070
rect 1889 7061 2830 7070
rect 2885 7104 3036 7138
rect 3070 7104 3076 7138
rect 2885 7066 3076 7104
rect 380 7013 386 7047
rect 420 7013 571 7047
rect 380 6988 571 7013
rect 2885 7032 3036 7066
rect 3070 7032 3076 7066
rect 380 6975 531 6988
rect 380 6941 386 6975
rect 420 6954 531 6975
rect 565 6954 571 6988
rect 420 6941 571 6954
rect 380 6915 571 6941
rect 380 6903 531 6915
rect 380 6869 386 6903
rect 420 6881 531 6903
rect 565 6881 571 6915
rect 420 6869 571 6881
rect 380 6842 571 6869
rect 380 6831 531 6842
rect 380 6797 386 6831
rect 420 6808 531 6831
rect 565 6808 571 6842
rect 420 6797 571 6808
rect 380 6769 571 6797
rect 380 6759 531 6769
rect 380 6725 386 6759
rect 420 6735 531 6759
rect 565 6735 571 6769
rect 420 6725 571 6735
rect 380 6696 571 6725
rect 380 6687 531 6696
rect 380 6653 386 6687
rect 420 6662 531 6687
rect 565 6662 571 6696
rect 420 6653 571 6662
rect 380 6623 571 6653
rect 380 6615 531 6623
rect 380 6581 386 6615
rect 420 6589 531 6615
rect 565 6589 571 6623
rect 420 6581 571 6589
rect 380 6550 571 6581
rect 761 6988 807 7000
rect 761 6954 767 6988
rect 801 6954 807 6988
rect 761 6915 807 6954
rect 761 6881 767 6915
rect 801 6881 807 6915
rect 761 6842 807 6881
rect 761 6808 767 6842
rect 801 6808 807 6842
rect 761 6769 807 6808
rect 761 6735 767 6769
rect 801 6735 807 6769
rect 761 6696 807 6735
rect 761 6662 767 6696
rect 801 6662 807 6696
rect 761 6623 807 6662
rect 761 6589 767 6623
rect 801 6589 807 6623
tri 571 6550 582 6561 sw
tri 750 6550 761 6561 se
rect 761 6550 807 6589
rect 997 6988 1043 7000
rect 997 6954 1003 6988
rect 1037 6954 1043 6988
rect 997 6915 1043 6954
rect 997 6881 1003 6915
rect 1037 6881 1043 6915
rect 997 6842 1043 6881
rect 997 6808 1003 6842
rect 1037 6808 1043 6842
rect 997 6769 1043 6808
rect 997 6735 1003 6769
rect 1037 6735 1043 6769
rect 997 6696 1043 6735
rect 997 6662 1003 6696
rect 1037 6662 1043 6696
rect 997 6623 1043 6662
rect 997 6589 1003 6623
rect 1037 6589 1043 6623
tri 807 6550 818 6561 sw
tri 986 6550 997 6561 se
rect 997 6550 1043 6589
rect 1233 6988 1279 7000
rect 1233 6954 1239 6988
rect 1273 6954 1279 6988
rect 1233 6915 1279 6954
rect 1233 6881 1239 6915
rect 1273 6881 1279 6915
rect 1233 6842 1279 6881
rect 1233 6808 1239 6842
rect 1273 6808 1279 6842
rect 1233 6769 1279 6808
rect 1233 6735 1239 6769
rect 1273 6735 1279 6769
rect 1233 6696 1279 6735
rect 1233 6662 1239 6696
rect 1273 6662 1279 6696
rect 1233 6623 1279 6662
rect 1233 6589 1239 6623
rect 1273 6589 1279 6623
tri 1043 6550 1054 6561 sw
tri 1222 6550 1233 6561 se
rect 1233 6550 1279 6589
rect 1469 6988 1515 7000
rect 1469 6954 1475 6988
rect 1509 6954 1515 6988
rect 1469 6915 1515 6954
rect 1469 6881 1475 6915
rect 1509 6881 1515 6915
rect 1469 6842 1515 6881
rect 1469 6808 1475 6842
rect 1509 6808 1515 6842
rect 1469 6769 1515 6808
rect 1469 6735 1475 6769
rect 1509 6735 1515 6769
rect 1469 6696 1515 6735
rect 1469 6662 1475 6696
rect 1509 6662 1515 6696
rect 1469 6623 1515 6662
rect 1469 6589 1475 6623
rect 1509 6589 1515 6623
tri 1279 6550 1290 6561 sw
tri 1458 6550 1469 6561 se
rect 1469 6550 1515 6589
rect 1705 6988 1751 7000
rect 1705 6954 1711 6988
rect 1745 6954 1751 6988
rect 1705 6915 1751 6954
rect 1705 6881 1711 6915
rect 1745 6881 1751 6915
rect 1705 6842 1751 6881
rect 1705 6808 1711 6842
rect 1745 6808 1751 6842
rect 1705 6769 1751 6808
rect 1705 6735 1711 6769
rect 1745 6735 1751 6769
rect 1705 6696 1751 6735
rect 1705 6662 1711 6696
rect 1745 6662 1751 6696
rect 1705 6623 1751 6662
rect 1705 6589 1711 6623
rect 1745 6589 1751 6623
tri 1515 6550 1526 6561 sw
tri 1694 6550 1705 6561 se
rect 1705 6550 1751 6589
rect 1941 6988 1987 7000
rect 1941 6954 1947 6988
rect 1981 6954 1987 6988
rect 1941 6915 1987 6954
rect 1941 6881 1947 6915
rect 1981 6881 1987 6915
rect 1941 6842 1987 6881
rect 1941 6808 1947 6842
rect 1981 6808 1987 6842
rect 1941 6769 1987 6808
rect 1941 6735 1947 6769
rect 1981 6735 1987 6769
rect 1941 6696 1987 6735
rect 1941 6662 1947 6696
rect 1981 6662 1987 6696
rect 1941 6623 1987 6662
rect 1941 6589 1947 6623
rect 1981 6589 1987 6623
tri 1751 6550 1762 6561 sw
tri 1930 6550 1941 6561 se
rect 1941 6550 1987 6589
rect 2177 6988 2223 7000
rect 2177 6954 2183 6988
rect 2217 6954 2223 6988
rect 2177 6915 2223 6954
rect 2177 6881 2183 6915
rect 2217 6881 2223 6915
rect 2177 6842 2223 6881
rect 2177 6808 2183 6842
rect 2217 6808 2223 6842
rect 2177 6769 2223 6808
rect 2177 6735 2183 6769
rect 2217 6735 2223 6769
rect 2177 6696 2223 6735
rect 2177 6662 2183 6696
rect 2217 6662 2223 6696
rect 2177 6623 2223 6662
rect 2177 6589 2183 6623
rect 2217 6589 2223 6623
tri 1987 6550 1998 6561 sw
tri 2166 6550 2177 6561 se
rect 2177 6550 2223 6589
rect 2413 6988 2459 7000
rect 2413 6954 2419 6988
rect 2453 6954 2459 6988
rect 2413 6915 2459 6954
rect 2413 6881 2419 6915
rect 2453 6881 2459 6915
rect 2413 6842 2459 6881
rect 2413 6808 2419 6842
rect 2453 6808 2459 6842
rect 2413 6769 2459 6808
rect 2413 6735 2419 6769
rect 2453 6735 2459 6769
rect 2413 6696 2459 6735
rect 2413 6662 2419 6696
rect 2453 6662 2459 6696
rect 2413 6623 2459 6662
rect 2413 6589 2419 6623
rect 2453 6589 2459 6623
tri 2223 6550 2234 6561 sw
tri 2402 6550 2413 6561 se
rect 2413 6550 2459 6589
rect 2649 6988 2695 7000
rect 2649 6954 2655 6988
rect 2689 6954 2695 6988
rect 2649 6915 2695 6954
rect 2649 6881 2655 6915
rect 2689 6881 2695 6915
rect 2649 6842 2695 6881
rect 2649 6808 2655 6842
rect 2689 6808 2695 6842
rect 2649 6769 2695 6808
rect 2649 6735 2655 6769
rect 2689 6735 2695 6769
rect 2649 6696 2695 6735
rect 2649 6662 2655 6696
rect 2689 6662 2695 6696
rect 2649 6623 2695 6662
rect 2649 6589 2655 6623
rect 2689 6589 2695 6623
tri 2459 6550 2470 6561 sw
tri 2638 6550 2649 6561 se
rect 2649 6550 2695 6589
rect 2885 6994 3076 7032
rect 2885 6988 3036 6994
rect 2885 6954 2891 6988
rect 2925 6960 3036 6988
rect 3070 6960 3076 6994
rect 2925 6954 3076 6960
rect 2885 6922 3076 6954
rect 2885 6915 3036 6922
rect 2885 6881 2891 6915
rect 2925 6888 3036 6915
rect 3070 6888 3076 6922
rect 2925 6881 3076 6888
rect 2885 6850 3076 6881
rect 2885 6842 3036 6850
rect 2885 6808 2891 6842
rect 2925 6816 3036 6842
rect 3070 6816 3076 6850
rect 2925 6808 3076 6816
rect 2885 6778 3076 6808
rect 2885 6769 3036 6778
rect 2885 6735 2891 6769
rect 2925 6744 3036 6769
rect 3070 6744 3076 6778
rect 2925 6735 3076 6744
rect 2885 6706 3076 6735
rect 2885 6696 3036 6706
rect 2885 6662 2891 6696
rect 2925 6672 3036 6696
rect 3070 6672 3076 6706
rect 2925 6662 3076 6672
rect 2885 6634 3076 6662
rect 2885 6623 3036 6634
rect 2885 6589 2891 6623
rect 2925 6600 3036 6623
rect 3070 6600 3076 6634
rect 2925 6589 3076 6600
rect 2885 6562 3076 6589
tri 2695 6550 2706 6561 sw
tri 2874 6550 2885 6561 se
rect 2885 6550 3036 6562
rect 380 6543 531 6550
rect 380 6509 386 6543
rect 420 6516 531 6543
rect 565 6527 582 6550
tri 582 6527 605 6550 sw
tri 727 6527 750 6550 se
rect 750 6527 767 6550
rect 565 6516 767 6527
rect 801 6527 818 6550
tri 818 6527 841 6550 sw
tri 963 6527 986 6550 se
rect 986 6527 1003 6550
rect 801 6516 1003 6527
rect 1037 6527 1054 6550
tri 1054 6527 1077 6550 sw
tri 1199 6527 1222 6550 se
rect 1222 6527 1239 6550
rect 1037 6516 1239 6527
rect 1273 6527 1290 6550
tri 1290 6527 1313 6550 sw
tri 1435 6527 1458 6550 se
rect 1458 6527 1475 6550
rect 1273 6516 1475 6527
rect 1509 6527 1526 6550
tri 1526 6527 1549 6550 sw
tri 1671 6527 1694 6550 se
rect 1694 6527 1711 6550
rect 1509 6516 1711 6527
rect 1745 6527 1762 6550
tri 1762 6527 1785 6550 sw
tri 1907 6527 1930 6550 se
rect 1930 6527 1947 6550
rect 1745 6516 1947 6527
rect 1981 6527 1998 6550
tri 1998 6527 2021 6550 sw
tri 2143 6527 2166 6550 se
rect 2166 6527 2183 6550
rect 1981 6516 2183 6527
rect 2217 6527 2234 6550
tri 2234 6527 2257 6550 sw
tri 2379 6527 2402 6550 se
rect 2402 6527 2419 6550
rect 2217 6516 2419 6527
rect 2453 6527 2470 6550
tri 2470 6527 2493 6550 sw
tri 2615 6527 2638 6550 se
rect 2638 6527 2655 6550
rect 2453 6516 2655 6527
rect 2689 6527 2706 6550
tri 2706 6527 2729 6550 sw
tri 2851 6527 2874 6550 se
rect 2874 6527 2891 6550
rect 2689 6516 2891 6527
rect 2925 6528 3036 6550
rect 3070 6528 3076 6562
rect 2925 6516 3076 6528
rect 420 6509 3076 6516
rect 380 6501 3076 6509
rect 380 6477 697 6501
rect 380 6471 531 6477
rect 380 6437 386 6471
rect 420 6443 531 6471
rect 565 6449 697 6477
rect 749 6449 765 6501
rect 817 6449 833 6501
rect 885 6449 901 6501
rect 953 6449 969 6501
rect 1021 6477 1037 6501
rect 1089 6449 1105 6501
rect 1157 6449 1173 6501
rect 1225 6477 1241 6501
rect 1293 6477 2097 6501
rect 1225 6449 1239 6477
rect 1293 6449 1475 6477
rect 565 6443 767 6449
rect 801 6443 1003 6449
rect 1037 6443 1239 6449
rect 1273 6443 1475 6449
rect 1509 6443 1711 6477
rect 1745 6443 1947 6477
rect 1981 6449 2097 6477
rect 2149 6449 2165 6501
rect 2217 6449 2233 6501
rect 2285 6449 2301 6501
rect 2353 6449 2369 6501
rect 2421 6477 2437 6501
rect 2489 6449 2505 6501
rect 2557 6449 2573 6501
rect 2625 6449 2641 6501
rect 2693 6490 3076 6501
rect 2693 6477 3036 6490
rect 2693 6449 2891 6477
rect 1981 6443 2183 6449
rect 2217 6443 2419 6449
rect 2453 6443 2655 6449
rect 2689 6443 2891 6449
rect 2925 6456 3036 6477
rect 3070 6456 3076 6490
rect 2925 6443 3076 6456
rect 420 6437 3076 6443
rect 380 6404 697 6437
rect 380 6399 531 6404
rect 380 6365 386 6399
rect 420 6370 531 6399
rect 565 6385 697 6404
rect 749 6385 765 6437
rect 817 6385 833 6437
rect 885 6385 901 6437
rect 953 6385 969 6437
rect 1021 6404 1037 6437
rect 1089 6385 1105 6437
rect 1157 6385 1173 6437
rect 1225 6404 1241 6437
rect 1293 6404 2097 6437
rect 1225 6385 1239 6404
rect 1293 6385 1475 6404
rect 565 6373 767 6385
rect 801 6373 1003 6385
rect 1037 6373 1239 6385
rect 1273 6373 1475 6385
rect 565 6370 697 6373
rect 420 6365 697 6370
rect 380 6331 697 6365
rect 380 6327 531 6331
rect 380 6293 386 6327
rect 420 6297 531 6327
rect 565 6321 697 6331
rect 749 6321 765 6373
rect 817 6321 833 6373
rect 885 6321 901 6373
rect 953 6321 969 6373
rect 1021 6331 1037 6370
rect 1089 6321 1105 6373
rect 1157 6321 1173 6373
rect 1225 6370 1239 6373
rect 1293 6370 1475 6373
rect 1509 6370 1711 6404
rect 1745 6370 1947 6404
rect 1981 6385 2097 6404
rect 2149 6385 2165 6437
rect 2217 6385 2233 6437
rect 2285 6385 2301 6437
rect 2353 6385 2369 6437
rect 2421 6404 2437 6437
rect 2489 6385 2505 6437
rect 2557 6385 2573 6437
rect 2625 6385 2641 6437
rect 2693 6418 3076 6437
rect 2693 6404 3036 6418
rect 2693 6385 2891 6404
rect 1981 6373 2183 6385
rect 2217 6373 2419 6385
rect 2453 6373 2655 6385
rect 2689 6373 2891 6385
rect 1981 6370 2097 6373
rect 1225 6331 1241 6370
rect 1293 6331 2097 6370
rect 1225 6321 1239 6331
rect 1293 6321 1475 6331
rect 565 6309 767 6321
rect 801 6309 1003 6321
rect 1037 6309 1239 6321
rect 1273 6309 1475 6321
rect 565 6297 697 6309
rect 420 6293 697 6297
rect 380 6258 697 6293
rect 380 6255 531 6258
rect 380 6221 386 6255
rect 420 6224 531 6255
rect 565 6257 697 6258
rect 749 6257 765 6309
rect 817 6257 833 6309
rect 885 6257 901 6309
rect 953 6257 969 6309
rect 1021 6258 1037 6297
rect 1089 6257 1105 6309
rect 1157 6257 1173 6309
rect 1225 6297 1239 6309
rect 1293 6297 1475 6309
rect 1509 6297 1711 6331
rect 1745 6297 1947 6331
rect 1981 6321 2097 6331
rect 2149 6321 2165 6373
rect 2217 6321 2233 6373
rect 2285 6321 2301 6373
rect 2353 6321 2369 6373
rect 2421 6331 2437 6370
rect 2489 6321 2505 6373
rect 2557 6321 2573 6373
rect 2625 6321 2641 6373
rect 2693 6370 2891 6373
rect 2925 6384 3036 6404
rect 3070 6384 3076 6418
rect 2925 6370 3076 6384
rect 2693 6346 3076 6370
rect 2693 6331 3036 6346
rect 2693 6321 2891 6331
rect 1981 6309 2183 6321
rect 2217 6309 2419 6321
rect 2453 6309 2655 6321
rect 2689 6309 2891 6321
rect 1981 6297 2097 6309
rect 1225 6258 1241 6297
rect 1293 6258 2097 6297
rect 1225 6257 1239 6258
rect 1293 6257 1475 6258
rect 565 6245 767 6257
rect 801 6245 1003 6257
rect 1037 6245 1239 6257
rect 1273 6245 1475 6257
rect 565 6224 697 6245
rect 420 6221 697 6224
rect 380 6193 697 6221
rect 749 6193 765 6245
rect 817 6193 833 6245
rect 885 6193 901 6245
rect 953 6193 969 6245
rect 1021 6193 1037 6224
rect 1089 6193 1105 6245
rect 1157 6193 1173 6245
rect 1225 6224 1239 6245
rect 1293 6224 1475 6245
rect 1509 6224 1711 6258
rect 1745 6224 1947 6258
rect 1981 6257 2097 6258
rect 2149 6257 2165 6309
rect 2217 6257 2233 6309
rect 2285 6257 2301 6309
rect 2353 6257 2369 6309
rect 2421 6258 2437 6297
rect 2489 6257 2505 6309
rect 2557 6257 2573 6309
rect 2625 6257 2641 6309
rect 2693 6297 2891 6309
rect 2925 6312 3036 6331
rect 3070 6312 3076 6346
rect 2925 6297 3076 6312
rect 2693 6274 3076 6297
rect 2693 6258 3036 6274
rect 2693 6257 2891 6258
rect 1981 6245 2183 6257
rect 2217 6245 2419 6257
rect 2453 6245 2655 6257
rect 2689 6245 2891 6257
rect 1981 6224 2097 6245
rect 1225 6193 1241 6224
rect 1293 6193 2097 6224
rect 2149 6193 2165 6245
rect 2217 6193 2233 6245
rect 2285 6193 2301 6245
rect 2353 6193 2369 6245
rect 2421 6193 2437 6224
rect 2489 6193 2505 6245
rect 2557 6193 2573 6245
rect 2625 6193 2641 6245
rect 2693 6224 2891 6245
rect 2925 6240 3036 6258
rect 3070 6240 3076 6274
rect 2925 6224 3076 6240
rect 2693 6202 3076 6224
rect 2693 6193 3036 6202
rect 380 6185 3036 6193
rect 380 6183 531 6185
rect 380 6149 386 6183
rect 420 6151 531 6183
rect 565 6181 767 6185
rect 801 6181 1003 6185
rect 1037 6181 1239 6185
rect 1273 6181 1475 6185
rect 565 6151 697 6181
rect 420 6149 697 6151
rect 380 6129 697 6149
rect 749 6129 765 6181
rect 817 6129 833 6181
rect 885 6129 901 6181
rect 953 6129 969 6181
rect 1021 6129 1037 6151
rect 1089 6129 1105 6181
rect 1157 6129 1173 6181
rect 1225 6151 1239 6181
rect 1293 6151 1475 6181
rect 1509 6151 1711 6185
rect 1745 6151 1947 6185
rect 1981 6181 2183 6185
rect 2217 6181 2419 6185
rect 2453 6181 2655 6185
rect 2689 6181 2891 6185
rect 1981 6151 2097 6181
rect 1225 6129 1241 6151
rect 1293 6129 2097 6151
rect 2149 6129 2165 6181
rect 2217 6129 2233 6181
rect 2285 6129 2301 6181
rect 2353 6129 2369 6181
rect 2421 6129 2437 6151
rect 2489 6129 2505 6181
rect 2557 6129 2573 6181
rect 2625 6129 2641 6181
rect 2693 6151 2891 6181
rect 2925 6168 3036 6185
rect 3070 6168 3076 6202
rect 2925 6151 3076 6168
rect 2693 6130 3076 6151
rect 2693 6129 3036 6130
rect 380 6117 3036 6129
rect 380 6112 697 6117
rect 380 6111 531 6112
rect 380 6077 386 6111
rect 420 6078 531 6111
rect 565 6078 697 6112
rect 420 6077 697 6078
rect 380 6065 697 6077
rect 749 6065 765 6117
rect 817 6065 833 6117
rect 885 6065 901 6117
rect 953 6065 969 6117
rect 1021 6112 1037 6117
rect 1021 6065 1037 6078
rect 1089 6065 1105 6117
rect 1157 6065 1173 6117
rect 1225 6112 1241 6117
rect 1293 6112 2097 6117
rect 1225 6078 1239 6112
rect 1293 6078 1475 6112
rect 1509 6078 1711 6112
rect 1745 6078 1947 6112
rect 1981 6078 2097 6112
rect 1225 6065 1241 6078
rect 1293 6065 2097 6078
rect 2149 6065 2165 6117
rect 2217 6065 2233 6117
rect 2285 6065 2301 6117
rect 2353 6065 2369 6117
rect 2421 6112 2437 6117
rect 2421 6065 2437 6078
rect 2489 6065 2505 6117
rect 2557 6065 2573 6117
rect 2625 6065 2641 6117
rect 2693 6112 3036 6117
rect 2693 6078 2891 6112
rect 2925 6096 3036 6112
rect 3070 6096 3076 6130
rect 2925 6078 3076 6096
rect 2693 6065 3076 6078
rect 380 6058 3076 6065
rect 380 6053 3036 6058
rect 380 6039 697 6053
rect 380 6005 386 6039
rect 420 6038 697 6039
rect 420 6005 531 6038
rect 380 6004 531 6005
rect 565 6004 697 6038
rect 380 6001 697 6004
rect 749 6001 765 6053
rect 817 6001 833 6053
rect 885 6001 901 6053
rect 953 6001 969 6053
rect 1021 6038 1037 6053
rect 1021 6001 1037 6004
rect 1089 6001 1105 6053
rect 1157 6001 1173 6053
rect 1225 6038 1241 6053
rect 1293 6038 2097 6053
rect 1225 6004 1239 6038
rect 1293 6004 1475 6038
rect 1509 6004 1711 6038
rect 1745 6004 1947 6038
rect 1981 6004 2097 6038
rect 1225 6001 1241 6004
rect 1293 6001 2097 6004
rect 2149 6001 2165 6053
rect 2217 6001 2233 6053
rect 2285 6001 2301 6053
rect 2353 6001 2369 6053
rect 2421 6038 2437 6053
rect 2421 6001 2437 6004
rect 2489 6001 2505 6053
rect 2557 6001 2573 6053
rect 2625 6001 2641 6053
rect 2693 6038 3036 6053
rect 2693 6004 2891 6038
rect 2925 6024 3036 6038
rect 3070 6024 3076 6058
rect 2925 6004 3076 6024
rect 2693 6001 3076 6004
rect 380 5989 3076 6001
rect 380 5967 697 5989
rect 380 5933 386 5967
rect 420 5964 697 5967
rect 420 5933 531 5964
rect 380 5930 531 5933
rect 565 5937 697 5964
rect 749 5937 765 5989
rect 817 5937 833 5989
rect 885 5937 901 5989
rect 953 5937 969 5989
rect 1021 5964 1037 5989
rect 1089 5937 1105 5989
rect 1157 5937 1173 5989
rect 1225 5964 1241 5989
rect 1293 5964 2097 5989
rect 1225 5937 1239 5964
rect 1293 5937 1475 5964
rect 565 5930 767 5937
rect 801 5930 1003 5937
rect 1037 5930 1239 5937
rect 1273 5930 1475 5937
rect 1509 5930 1711 5964
rect 1745 5930 1947 5964
rect 1981 5937 2097 5964
rect 2149 5937 2165 5989
rect 2217 5937 2233 5989
rect 2285 5937 2301 5989
rect 2353 5937 2369 5989
rect 2421 5964 2437 5989
rect 2489 5937 2505 5989
rect 2557 5937 2573 5989
rect 2625 5937 2641 5989
rect 2693 5986 3076 5989
rect 2693 5964 3036 5986
rect 2693 5937 2891 5964
rect 1981 5930 2183 5937
rect 2217 5930 2419 5937
rect 2453 5930 2655 5937
rect 2689 5930 2891 5937
rect 2925 5952 3036 5964
rect 3070 5952 3076 5986
rect 2925 5930 3076 5952
rect 380 5925 3076 5930
rect 380 5895 697 5925
rect 380 5861 386 5895
rect 420 5890 697 5895
rect 420 5861 531 5890
rect 380 5856 531 5861
rect 565 5873 697 5890
rect 749 5873 765 5925
rect 817 5873 833 5925
rect 885 5873 901 5925
rect 953 5873 969 5925
rect 1021 5890 1037 5925
rect 1089 5873 1105 5925
rect 1157 5873 1173 5925
rect 1225 5890 1241 5925
rect 1293 5890 2097 5925
rect 1225 5873 1239 5890
rect 1293 5873 1475 5890
rect 565 5861 767 5873
rect 801 5861 1003 5873
rect 1037 5861 1239 5873
rect 1273 5861 1475 5873
rect 565 5856 697 5861
rect 380 5823 697 5856
rect 380 5789 386 5823
rect 420 5816 697 5823
rect 420 5789 531 5816
rect 380 5782 531 5789
rect 565 5809 697 5816
rect 749 5809 765 5861
rect 817 5809 833 5861
rect 885 5809 901 5861
rect 953 5809 969 5861
rect 1021 5816 1037 5856
rect 1089 5809 1105 5861
rect 1157 5809 1173 5861
rect 1225 5856 1239 5861
rect 1293 5856 1475 5861
rect 1509 5856 1711 5890
rect 1745 5856 1947 5890
rect 1981 5873 2097 5890
rect 2149 5873 2165 5925
rect 2217 5873 2233 5925
rect 2285 5873 2301 5925
rect 2353 5873 2369 5925
rect 2421 5890 2437 5925
rect 2489 5873 2505 5925
rect 2557 5873 2573 5925
rect 2625 5873 2641 5925
rect 2693 5914 3076 5925
rect 2693 5890 3036 5914
rect 2693 5873 2891 5890
rect 1981 5861 2183 5873
rect 2217 5861 2419 5873
rect 2453 5861 2655 5873
rect 2689 5861 2891 5873
rect 1981 5856 2097 5861
rect 1225 5816 1241 5856
rect 1293 5816 2097 5856
rect 1225 5809 1239 5816
rect 1293 5809 1475 5816
rect 565 5797 767 5809
rect 801 5797 1003 5809
rect 1037 5797 1239 5809
rect 1273 5797 1475 5809
rect 565 5782 697 5797
rect 380 5751 697 5782
rect 380 5717 386 5751
rect 420 5745 697 5751
rect 749 5745 765 5797
rect 817 5745 833 5797
rect 885 5745 901 5797
rect 953 5745 969 5797
rect 1021 5745 1037 5782
rect 1089 5745 1105 5797
rect 1157 5745 1173 5797
rect 1225 5782 1239 5797
rect 1293 5782 1475 5797
rect 1509 5782 1711 5816
rect 1745 5782 1947 5816
rect 1981 5809 2097 5816
rect 2149 5809 2165 5861
rect 2217 5809 2233 5861
rect 2285 5809 2301 5861
rect 2353 5809 2369 5861
rect 2421 5816 2437 5856
rect 2489 5809 2505 5861
rect 2557 5809 2573 5861
rect 2625 5809 2641 5861
rect 2693 5856 2891 5861
rect 2925 5880 3036 5890
rect 3070 5880 3076 5914
rect 2925 5856 3076 5880
rect 2693 5842 3076 5856
rect 2693 5816 3036 5842
rect 2693 5809 2891 5816
rect 1981 5797 2183 5809
rect 2217 5797 2419 5809
rect 2453 5797 2655 5809
rect 2689 5797 2891 5809
rect 1981 5782 2097 5797
rect 1225 5745 1241 5782
rect 1293 5745 2097 5782
rect 2149 5745 2165 5797
rect 2217 5745 2233 5797
rect 2285 5745 2301 5797
rect 2353 5745 2369 5797
rect 2421 5745 2437 5782
rect 2489 5745 2505 5797
rect 2557 5745 2573 5797
rect 2625 5745 2641 5797
rect 2693 5782 2891 5797
rect 2925 5808 3036 5816
rect 3070 5808 3076 5842
rect 2925 5782 3076 5808
rect 2693 5770 3076 5782
rect 2693 5745 3036 5770
rect 420 5742 3036 5745
rect 420 5717 531 5742
rect 380 5708 531 5717
rect 565 5733 767 5742
rect 801 5733 1003 5742
rect 1037 5733 1239 5742
rect 1273 5733 1475 5742
rect 565 5708 697 5733
rect 380 5681 697 5708
rect 749 5681 765 5733
rect 817 5681 833 5733
rect 885 5681 901 5733
rect 953 5681 969 5733
rect 1021 5681 1037 5708
rect 1089 5681 1105 5733
rect 1157 5681 1173 5733
rect 1225 5708 1239 5733
rect 1293 5708 1475 5733
rect 1509 5708 1711 5742
rect 1745 5708 1947 5742
rect 1981 5733 2183 5742
rect 2217 5733 2419 5742
rect 2453 5733 2655 5742
rect 2689 5733 2891 5742
rect 1981 5708 2097 5733
rect 1225 5681 1241 5708
rect 1293 5681 2097 5708
rect 2149 5681 2165 5733
rect 2217 5681 2233 5733
rect 2285 5681 2301 5733
rect 2353 5681 2369 5733
rect 2421 5681 2437 5708
rect 2489 5681 2505 5733
rect 2557 5681 2573 5733
rect 2625 5681 2641 5733
rect 2693 5708 2891 5733
rect 2925 5736 3036 5742
rect 3070 5736 3076 5770
rect 2925 5708 3076 5736
rect 2693 5698 3076 5708
rect 2693 5681 3036 5698
rect 380 5679 3036 5681
rect 380 5645 386 5679
rect 420 5669 3036 5679
rect 420 5668 697 5669
rect 420 5645 531 5668
rect 380 5634 531 5645
rect 565 5634 697 5668
rect 380 5617 697 5634
rect 749 5617 765 5669
rect 817 5617 833 5669
rect 885 5617 901 5669
rect 953 5617 969 5669
rect 1021 5668 1037 5669
rect 1021 5617 1037 5634
rect 1089 5617 1105 5669
rect 1157 5617 1173 5669
rect 1225 5668 1241 5669
rect 1293 5668 2097 5669
rect 1225 5634 1239 5668
rect 1293 5634 1475 5668
rect 1509 5634 1711 5668
rect 1745 5634 1947 5668
rect 1981 5634 2097 5668
rect 1225 5617 1241 5634
rect 1293 5617 2097 5634
rect 2149 5617 2165 5669
rect 2217 5617 2233 5669
rect 2285 5617 2301 5669
rect 2353 5617 2369 5669
rect 2421 5668 2437 5669
rect 2421 5617 2437 5634
rect 2489 5617 2505 5669
rect 2557 5617 2573 5669
rect 2625 5617 2641 5669
rect 2693 5668 3036 5669
rect 2693 5634 2891 5668
rect 2925 5664 3036 5668
rect 3070 5664 3076 5698
rect 2925 5634 3076 5664
rect 2693 5626 3076 5634
rect 2693 5617 3036 5626
rect 380 5607 3036 5617
rect 380 5573 386 5607
rect 420 5605 3036 5607
rect 420 5594 697 5605
rect 420 5573 531 5594
rect 380 5560 531 5573
rect 565 5560 697 5594
rect 380 5553 697 5560
rect 749 5553 765 5605
rect 817 5553 833 5605
rect 885 5553 901 5605
rect 953 5553 969 5605
rect 1021 5594 1037 5605
rect 1021 5553 1037 5560
rect 1089 5553 1105 5605
rect 1157 5553 1173 5605
rect 1225 5594 1241 5605
rect 1293 5594 2097 5605
rect 1225 5560 1239 5594
rect 1293 5560 1475 5594
rect 1509 5560 1711 5594
rect 1745 5560 1947 5594
rect 1981 5560 2097 5594
rect 1225 5553 1241 5560
rect 1293 5553 2097 5560
rect 2149 5553 2165 5605
rect 2217 5553 2233 5605
rect 2285 5553 2301 5605
rect 2353 5553 2369 5605
rect 2421 5594 2437 5605
rect 2421 5553 2437 5560
rect 2489 5553 2505 5605
rect 2557 5553 2573 5605
rect 2625 5553 2641 5605
rect 2693 5594 3036 5605
rect 2693 5560 2891 5594
rect 2925 5592 3036 5594
rect 3070 5592 3076 5626
rect 2925 5560 3076 5592
rect 2693 5554 3076 5560
rect 2693 5553 3036 5554
rect 380 5535 3036 5553
rect 380 5501 386 5535
rect 420 5527 3036 5535
rect 420 5520 598 5527
tri 598 5520 605 5527 nw
tri 727 5520 734 5527 ne
rect 734 5520 834 5527
tri 834 5520 841 5527 nw
tri 963 5520 970 5527 ne
rect 970 5520 1070 5527
tri 1070 5520 1077 5527 nw
tri 1199 5520 1206 5527 ne
rect 1206 5520 1306 5527
tri 1306 5520 1313 5527 nw
tri 1435 5520 1442 5527 ne
rect 1442 5520 1542 5527
tri 1542 5520 1549 5527 nw
tri 1671 5520 1678 5527 ne
rect 1678 5520 1778 5527
tri 1778 5520 1785 5527 nw
tri 1907 5520 1914 5527 ne
rect 1914 5520 2014 5527
tri 2014 5520 2021 5527 nw
tri 2143 5520 2150 5527 ne
rect 2150 5520 2250 5527
tri 2250 5520 2257 5527 nw
tri 2379 5520 2386 5527 ne
rect 2386 5520 2486 5527
tri 2486 5520 2493 5527 nw
tri 2615 5520 2622 5527 ne
rect 2622 5520 2722 5527
tri 2722 5520 2729 5527 nw
tri 2851 5520 2858 5527 ne
rect 2858 5520 3036 5527
rect 3070 5520 3076 5554
rect 420 5501 531 5520
rect 380 5486 531 5501
rect 565 5486 571 5520
tri 571 5493 598 5520 nw
tri 734 5493 761 5520 ne
rect 380 5463 571 5486
rect 380 5429 386 5463
rect 420 5446 571 5463
rect 420 5429 531 5446
rect 380 5412 531 5429
rect 565 5412 571 5446
rect 380 5391 571 5412
rect 380 5357 386 5391
rect 420 5372 571 5391
rect 420 5357 531 5372
rect 380 5338 531 5357
rect 565 5338 571 5372
rect 380 5319 571 5338
rect 380 5285 386 5319
rect 420 5298 571 5319
rect 420 5285 531 5298
rect 380 5264 531 5285
rect 565 5264 571 5298
rect 380 5247 571 5264
rect 380 5213 386 5247
rect 420 5224 571 5247
rect 420 5213 531 5224
rect 380 5190 531 5213
rect 565 5190 571 5224
rect 380 5175 571 5190
rect 380 5141 386 5175
rect 420 5150 571 5175
rect 420 5141 531 5150
rect 380 5116 531 5141
rect 565 5116 571 5150
rect 380 5103 571 5116
rect 380 5069 386 5103
rect 420 5076 571 5103
rect 420 5069 531 5076
rect 380 5042 531 5069
rect 565 5042 571 5076
rect 380 5031 571 5042
rect 380 4997 386 5031
rect 420 4997 571 5031
rect 761 5486 767 5520
rect 801 5486 807 5520
tri 807 5493 834 5520 nw
tri 970 5493 997 5520 ne
rect 761 5446 807 5486
rect 761 5412 767 5446
rect 801 5412 807 5446
rect 761 5372 807 5412
rect 761 5338 767 5372
rect 801 5338 807 5372
rect 761 5298 807 5338
rect 761 5264 767 5298
rect 801 5264 807 5298
rect 761 5224 807 5264
rect 761 5190 767 5224
rect 801 5190 807 5224
rect 761 5150 807 5190
rect 761 5116 767 5150
rect 801 5116 807 5150
rect 761 5076 807 5116
rect 761 5042 767 5076
rect 801 5042 807 5076
rect 761 5030 807 5042
rect 997 5486 1003 5520
rect 1037 5486 1043 5520
tri 1043 5493 1070 5520 nw
tri 1206 5493 1233 5520 ne
rect 997 5446 1043 5486
rect 997 5412 1003 5446
rect 1037 5412 1043 5446
rect 997 5372 1043 5412
rect 997 5338 1003 5372
rect 1037 5338 1043 5372
rect 997 5298 1043 5338
rect 997 5264 1003 5298
rect 1037 5264 1043 5298
rect 997 5224 1043 5264
rect 997 5190 1003 5224
rect 1037 5190 1043 5224
rect 997 5150 1043 5190
rect 997 5116 1003 5150
rect 1037 5116 1043 5150
rect 997 5076 1043 5116
rect 997 5042 1003 5076
rect 1037 5042 1043 5076
rect 997 5030 1043 5042
rect 1233 5486 1239 5520
rect 1273 5486 1279 5520
tri 1279 5493 1306 5520 nw
tri 1442 5493 1469 5520 ne
rect 1233 5446 1279 5486
rect 1233 5412 1239 5446
rect 1273 5412 1279 5446
rect 1233 5372 1279 5412
rect 1233 5338 1239 5372
rect 1273 5338 1279 5372
rect 1233 5298 1279 5338
rect 1233 5264 1239 5298
rect 1273 5264 1279 5298
rect 1233 5224 1279 5264
rect 1233 5190 1239 5224
rect 1273 5190 1279 5224
rect 1233 5150 1279 5190
rect 1233 5116 1239 5150
rect 1273 5116 1279 5150
rect 1233 5076 1279 5116
rect 1233 5042 1239 5076
rect 1273 5042 1279 5076
rect 1233 5030 1279 5042
rect 1469 5486 1475 5520
rect 1509 5486 1515 5520
tri 1515 5493 1542 5520 nw
tri 1678 5493 1705 5520 ne
rect 1469 5446 1515 5486
rect 1469 5412 1475 5446
rect 1509 5412 1515 5446
rect 1469 5372 1515 5412
rect 1469 5338 1475 5372
rect 1509 5338 1515 5372
rect 1469 5298 1515 5338
rect 1469 5264 1475 5298
rect 1509 5264 1515 5298
rect 1469 5224 1515 5264
rect 1469 5190 1475 5224
rect 1509 5190 1515 5224
rect 1469 5150 1515 5190
rect 1469 5116 1475 5150
rect 1509 5116 1515 5150
rect 1469 5076 1515 5116
rect 1469 5042 1475 5076
rect 1509 5042 1515 5076
rect 1469 5030 1515 5042
rect 1705 5486 1711 5520
rect 1745 5486 1751 5520
tri 1751 5493 1778 5520 nw
tri 1914 5493 1941 5520 ne
rect 1705 5446 1751 5486
rect 1705 5412 1711 5446
rect 1745 5412 1751 5446
rect 1705 5372 1751 5412
rect 1705 5338 1711 5372
rect 1745 5338 1751 5372
rect 1705 5298 1751 5338
rect 1705 5264 1711 5298
rect 1745 5264 1751 5298
rect 1705 5224 1751 5264
rect 1705 5190 1711 5224
rect 1745 5190 1751 5224
rect 1705 5150 1751 5190
rect 1705 5116 1711 5150
rect 1745 5116 1751 5150
rect 1705 5076 1751 5116
rect 1705 5042 1711 5076
rect 1745 5042 1751 5076
rect 1705 5030 1751 5042
rect 1941 5486 1947 5520
rect 1981 5486 1987 5520
tri 1987 5493 2014 5520 nw
tri 2150 5493 2177 5520 ne
rect 1941 5446 1987 5486
rect 1941 5412 1947 5446
rect 1981 5412 1987 5446
rect 1941 5372 1987 5412
rect 1941 5338 1947 5372
rect 1981 5338 1987 5372
rect 1941 5298 1987 5338
rect 1941 5264 1947 5298
rect 1981 5264 1987 5298
rect 1941 5224 1987 5264
rect 1941 5190 1947 5224
rect 1981 5190 1987 5224
rect 1941 5150 1987 5190
rect 1941 5116 1947 5150
rect 1981 5116 1987 5150
rect 1941 5076 1987 5116
rect 1941 5042 1947 5076
rect 1981 5042 1987 5076
rect 1941 5030 1987 5042
rect 2177 5486 2183 5520
rect 2217 5486 2223 5520
tri 2223 5493 2250 5520 nw
tri 2386 5493 2413 5520 ne
rect 2177 5446 2223 5486
rect 2177 5412 2183 5446
rect 2217 5412 2223 5446
rect 2177 5372 2223 5412
rect 2177 5338 2183 5372
rect 2217 5338 2223 5372
rect 2177 5298 2223 5338
rect 2177 5264 2183 5298
rect 2217 5264 2223 5298
rect 2177 5224 2223 5264
rect 2177 5190 2183 5224
rect 2217 5190 2223 5224
rect 2177 5150 2223 5190
rect 2177 5116 2183 5150
rect 2217 5116 2223 5150
rect 2177 5076 2223 5116
rect 2177 5042 2183 5076
rect 2217 5042 2223 5076
rect 2177 5030 2223 5042
rect 2413 5486 2419 5520
rect 2453 5486 2459 5520
tri 2459 5493 2486 5520 nw
tri 2622 5493 2649 5520 ne
rect 2413 5446 2459 5486
rect 2413 5412 2419 5446
rect 2453 5412 2459 5446
rect 2413 5372 2459 5412
rect 2413 5338 2419 5372
rect 2453 5338 2459 5372
rect 2413 5298 2459 5338
rect 2413 5264 2419 5298
rect 2453 5264 2459 5298
rect 2413 5224 2459 5264
rect 2413 5190 2419 5224
rect 2453 5190 2459 5224
rect 2413 5150 2459 5190
rect 2413 5116 2419 5150
rect 2453 5116 2459 5150
rect 2413 5076 2459 5116
rect 2413 5042 2419 5076
rect 2453 5042 2459 5076
rect 2413 5030 2459 5042
rect 2649 5486 2655 5520
rect 2689 5486 2695 5520
tri 2695 5493 2722 5520 nw
tri 2858 5493 2885 5520 ne
rect 2649 5446 2695 5486
rect 2649 5412 2655 5446
rect 2689 5412 2695 5446
rect 2649 5372 2695 5412
rect 2649 5338 2655 5372
rect 2689 5338 2695 5372
rect 2649 5298 2695 5338
rect 2649 5264 2655 5298
rect 2689 5264 2695 5298
rect 2649 5224 2695 5264
rect 2649 5190 2655 5224
rect 2689 5190 2695 5224
rect 2649 5150 2695 5190
rect 2649 5116 2655 5150
rect 2689 5116 2695 5150
rect 2649 5076 2695 5116
rect 2649 5042 2655 5076
rect 2689 5042 2695 5076
rect 2649 5030 2695 5042
rect 2885 5486 2891 5520
rect 2925 5486 3076 5520
rect 2885 5482 3076 5486
rect 2885 5448 3036 5482
rect 3070 5448 3076 5482
rect 2885 5446 3076 5448
rect 2885 5412 2891 5446
rect 2925 5412 3076 5446
rect 2885 5410 3076 5412
rect 2885 5376 3036 5410
rect 3070 5376 3076 5410
rect 2885 5372 3076 5376
rect 2885 5338 2891 5372
rect 2925 5338 3076 5372
rect 2885 5304 3036 5338
rect 3070 5304 3076 5338
rect 2885 5298 3076 5304
rect 2885 5264 2891 5298
rect 2925 5266 3076 5298
rect 2925 5264 3036 5266
rect 2885 5232 3036 5264
rect 3070 5232 3076 5266
rect 2885 5224 3076 5232
rect 2885 5190 2891 5224
rect 2925 5194 3076 5224
rect 2925 5190 3036 5194
rect 2885 5160 3036 5190
rect 3070 5160 3076 5194
rect 2885 5150 3076 5160
rect 2885 5116 2891 5150
rect 2925 5122 3076 5150
rect 2925 5116 3036 5122
rect 2885 5088 3036 5116
rect 3070 5088 3076 5122
rect 2885 5076 3076 5088
rect 2885 5042 2891 5076
rect 2925 5050 3076 5076
rect 2925 5042 3036 5050
rect 380 4959 571 4997
rect 2885 5016 3036 5042
rect 3070 5016 3076 5050
rect 380 4925 386 4959
rect 420 4925 571 4959
rect 613 4974 1501 4983
rect 1553 4974 1569 4983
rect 1621 4974 1636 4983
rect 1688 4974 1703 4983
rect 1755 4974 1770 4983
rect 1822 4974 1837 4983
rect 1889 4974 2830 4983
rect 613 4940 625 4974
rect 659 4940 700 4974
rect 734 4940 775 4974
rect 809 4940 850 4974
rect 884 4940 925 4974
rect 959 4940 1000 4974
rect 1034 4940 1075 4974
rect 1109 4940 1150 4974
rect 1184 4940 1225 4974
rect 1259 4940 1300 4974
rect 1334 4940 1375 4974
rect 1409 4940 1450 4974
rect 1484 4940 1501 4974
rect 1559 4940 1569 4974
rect 1634 4940 1636 4974
rect 1889 4940 1896 4974
rect 1930 4940 1970 4974
rect 2004 4940 2044 4974
rect 2078 4940 2118 4974
rect 2152 4940 2192 4974
rect 2226 4940 2266 4974
rect 2300 4940 2340 4974
rect 2374 4940 2414 4974
rect 2448 4940 2488 4974
rect 2522 4940 2562 4974
rect 2596 4940 2636 4974
rect 2670 4940 2710 4974
rect 2744 4940 2784 4974
rect 2818 4940 2830 4974
rect 613 4931 1501 4940
rect 1553 4931 1569 4940
rect 1621 4931 1636 4940
rect 1688 4931 1703 4940
rect 1755 4931 1770 4940
rect 1822 4931 1837 4940
rect 1889 4931 2830 4940
rect 2885 4978 3076 5016
rect 2885 4944 3036 4978
rect 3070 4944 3076 4978
rect 380 4887 571 4925
rect 380 4853 386 4887
rect 420 4872 571 4887
rect 2885 4906 3076 4944
rect 420 4853 531 4872
rect 380 4838 531 4853
rect 565 4838 571 4872
rect 380 4815 571 4838
rect 380 4781 386 4815
rect 420 4799 571 4815
rect 420 4781 531 4799
rect 380 4765 531 4781
rect 565 4765 571 4799
rect 380 4743 571 4765
rect 380 4709 386 4743
rect 420 4726 571 4743
rect 420 4709 531 4726
rect 380 4692 531 4709
rect 565 4692 571 4726
rect 380 4671 571 4692
rect 380 4637 386 4671
rect 420 4653 571 4671
rect 420 4637 531 4653
rect 380 4619 531 4637
rect 565 4619 571 4653
rect 380 4599 571 4619
rect 380 4565 386 4599
rect 420 4580 571 4599
rect 420 4565 531 4580
rect 380 4546 531 4565
rect 565 4546 571 4580
rect 380 4527 571 4546
rect 380 4493 386 4527
rect 420 4507 571 4527
rect 420 4493 531 4507
rect 380 4473 531 4493
rect 565 4473 571 4507
rect 761 4872 807 4884
rect 761 4838 767 4872
rect 801 4838 807 4872
rect 761 4799 807 4838
rect 761 4765 767 4799
rect 801 4765 807 4799
rect 761 4726 807 4765
rect 761 4692 767 4726
rect 801 4692 807 4726
rect 761 4653 807 4692
rect 761 4619 767 4653
rect 801 4619 807 4653
rect 761 4580 807 4619
rect 761 4546 767 4580
rect 801 4546 807 4580
rect 761 4507 807 4546
tri 571 4473 591 4493 sw
tri 741 4473 761 4493 se
rect 761 4473 767 4507
rect 801 4473 807 4507
rect 997 4872 1043 4884
rect 997 4838 1003 4872
rect 1037 4838 1043 4872
rect 997 4799 1043 4838
rect 997 4765 1003 4799
rect 1037 4765 1043 4799
rect 997 4726 1043 4765
rect 997 4692 1003 4726
rect 1037 4692 1043 4726
rect 997 4653 1043 4692
rect 997 4619 1003 4653
rect 1037 4619 1043 4653
rect 997 4580 1043 4619
rect 997 4546 1003 4580
rect 1037 4546 1043 4580
rect 997 4507 1043 4546
tri 807 4473 827 4493 sw
tri 977 4473 997 4493 se
rect 997 4473 1003 4507
rect 1037 4473 1043 4507
rect 1233 4872 1279 4884
rect 1233 4838 1239 4872
rect 1273 4838 1279 4872
rect 1233 4799 1279 4838
rect 1233 4765 1239 4799
rect 1273 4765 1279 4799
rect 1233 4726 1279 4765
rect 1233 4692 1239 4726
rect 1273 4692 1279 4726
rect 1233 4653 1279 4692
rect 1233 4619 1239 4653
rect 1273 4619 1279 4653
rect 1233 4580 1279 4619
rect 1233 4546 1239 4580
rect 1273 4546 1279 4580
rect 1233 4507 1279 4546
tri 1043 4473 1063 4493 sw
tri 1213 4473 1233 4493 se
rect 1233 4473 1239 4507
rect 1273 4473 1279 4507
rect 1469 4872 1515 4884
rect 1469 4838 1475 4872
rect 1509 4838 1515 4872
rect 1469 4799 1515 4838
rect 1469 4765 1475 4799
rect 1509 4765 1515 4799
rect 1469 4726 1515 4765
rect 1469 4692 1475 4726
rect 1509 4692 1515 4726
rect 1469 4653 1515 4692
rect 1469 4619 1475 4653
rect 1509 4619 1515 4653
rect 1469 4580 1515 4619
rect 1469 4546 1475 4580
rect 1509 4546 1515 4580
rect 1469 4507 1515 4546
tri 1279 4473 1299 4493 sw
tri 1449 4473 1469 4493 se
rect 1469 4473 1475 4507
rect 1509 4473 1515 4507
rect 1705 4872 1751 4884
rect 1705 4838 1711 4872
rect 1745 4838 1751 4872
rect 1705 4799 1751 4838
rect 1705 4765 1711 4799
rect 1745 4765 1751 4799
rect 1705 4726 1751 4765
rect 1705 4692 1711 4726
rect 1745 4692 1751 4726
rect 1705 4653 1751 4692
rect 1705 4619 1711 4653
rect 1745 4619 1751 4653
rect 1705 4580 1751 4619
rect 1705 4546 1711 4580
rect 1745 4546 1751 4580
rect 1705 4507 1751 4546
tri 1515 4473 1535 4493 sw
tri 1685 4473 1705 4493 se
rect 1705 4473 1711 4507
rect 1745 4473 1751 4507
rect 1941 4872 1987 4884
rect 1941 4838 1947 4872
rect 1981 4838 1987 4872
rect 1941 4799 1987 4838
rect 1941 4765 1947 4799
rect 1981 4765 1987 4799
rect 1941 4726 1987 4765
rect 1941 4692 1947 4726
rect 1981 4692 1987 4726
rect 1941 4653 1987 4692
rect 1941 4619 1947 4653
rect 1981 4619 1987 4653
rect 1941 4580 1987 4619
rect 1941 4546 1947 4580
rect 1981 4546 1987 4580
rect 1941 4507 1987 4546
tri 1751 4473 1771 4493 sw
tri 1921 4473 1941 4493 se
rect 1941 4473 1947 4507
rect 1981 4473 1987 4507
rect 2177 4872 2223 4884
rect 2177 4838 2183 4872
rect 2217 4838 2223 4872
rect 2177 4799 2223 4838
rect 2177 4765 2183 4799
rect 2217 4765 2223 4799
rect 2177 4726 2223 4765
rect 2177 4692 2183 4726
rect 2217 4692 2223 4726
rect 2177 4653 2223 4692
rect 2177 4619 2183 4653
rect 2217 4619 2223 4653
rect 2177 4580 2223 4619
rect 2177 4546 2183 4580
rect 2217 4546 2223 4580
rect 2177 4507 2223 4546
tri 1987 4473 2007 4493 sw
tri 2157 4473 2177 4493 se
rect 2177 4473 2183 4507
rect 2217 4473 2223 4507
rect 2413 4872 2459 4884
rect 2413 4838 2419 4872
rect 2453 4838 2459 4872
rect 2413 4799 2459 4838
rect 2413 4765 2419 4799
rect 2453 4765 2459 4799
rect 2413 4726 2459 4765
rect 2413 4692 2419 4726
rect 2453 4692 2459 4726
rect 2413 4653 2459 4692
rect 2413 4619 2419 4653
rect 2453 4619 2459 4653
rect 2413 4580 2459 4619
rect 2413 4546 2419 4580
rect 2453 4546 2459 4580
rect 2413 4507 2459 4546
tri 2223 4473 2243 4493 sw
tri 2393 4473 2413 4493 se
rect 2413 4473 2419 4507
rect 2453 4473 2459 4507
rect 2649 4872 2695 4884
rect 2649 4838 2655 4872
rect 2689 4838 2695 4872
rect 2649 4799 2695 4838
rect 2649 4765 2655 4799
rect 2689 4765 2695 4799
rect 2649 4726 2695 4765
rect 2649 4692 2655 4726
rect 2689 4692 2695 4726
rect 2649 4653 2695 4692
rect 2649 4619 2655 4653
rect 2689 4619 2695 4653
rect 2649 4580 2695 4619
rect 2649 4546 2655 4580
rect 2689 4546 2695 4580
rect 2649 4507 2695 4546
tri 2459 4473 2479 4493 sw
tri 2629 4473 2649 4493 se
rect 2649 4473 2655 4507
rect 2689 4473 2695 4507
rect 2885 4872 3036 4906
rect 3070 4872 3076 4906
rect 2885 4838 2891 4872
rect 2925 4838 3076 4872
rect 2885 4834 3076 4838
rect 2885 4800 3036 4834
rect 3070 4800 3076 4834
rect 2885 4799 3076 4800
rect 2885 4765 2891 4799
rect 2925 4765 3076 4799
rect 2885 4762 3076 4765
rect 2885 4728 3036 4762
rect 3070 4728 3076 4762
rect 2885 4726 3076 4728
rect 2885 4692 2891 4726
rect 2925 4692 3076 4726
rect 2885 4690 3076 4692
rect 2885 4656 3036 4690
rect 3070 4656 3076 4690
rect 2885 4653 3076 4656
rect 2885 4619 2891 4653
rect 2925 4619 3076 4653
rect 2885 4618 3076 4619
rect 2885 4584 3036 4618
rect 3070 4584 3076 4618
rect 2885 4580 3076 4584
rect 2885 4546 2891 4580
rect 2925 4546 3076 4580
rect 2885 4512 3036 4546
rect 3070 4512 3076 4546
rect 2885 4507 3076 4512
tri 2695 4473 2715 4493 sw
tri 2865 4473 2885 4493 se
rect 2885 4473 2891 4507
rect 2925 4474 3076 4507
rect 2925 4473 3036 4474
rect 380 4459 591 4473
tri 591 4459 605 4473 sw
tri 727 4459 741 4473 se
rect 741 4459 827 4473
tri 827 4459 841 4473 sw
tri 963 4459 977 4473 se
rect 977 4459 1063 4473
tri 1063 4459 1077 4473 sw
tri 1199 4459 1213 4473 se
rect 1213 4459 1299 4473
tri 1299 4459 1313 4473 sw
tri 1435 4459 1449 4473 se
rect 1449 4459 1535 4473
tri 1535 4459 1549 4473 sw
tri 1671 4459 1685 4473 se
rect 1685 4459 1771 4473
tri 1771 4459 1785 4473 sw
tri 1907 4459 1921 4473 se
rect 1921 4459 2007 4473
tri 2007 4459 2021 4473 sw
tri 2143 4459 2157 4473 se
rect 2157 4459 2243 4473
tri 2243 4459 2257 4473 sw
tri 2379 4459 2393 4473 se
rect 2393 4459 2479 4473
tri 2479 4459 2493 4473 sw
tri 2615 4459 2629 4473 se
rect 2629 4459 2715 4473
tri 2715 4459 2729 4473 sw
tri 2851 4459 2865 4473 se
rect 2865 4459 3036 4473
rect 380 4455 3036 4459
rect 380 4421 386 4455
rect 420 4440 3036 4455
rect 3070 4440 3076 4474
rect 420 4437 3076 4440
rect 420 4434 697 4437
rect 420 4421 531 4434
rect 380 4400 531 4421
rect 565 4400 697 4434
rect 380 4385 697 4400
rect 749 4385 765 4437
rect 817 4385 833 4437
rect 885 4385 901 4437
rect 953 4385 969 4437
rect 1021 4434 1037 4437
rect 1021 4385 1037 4400
rect 1089 4385 1105 4437
rect 1157 4385 1173 4437
rect 1225 4434 1241 4437
rect 1293 4434 2097 4437
rect 1225 4400 1239 4434
rect 1293 4400 1475 4434
rect 1509 4400 1711 4434
rect 1745 4400 1947 4434
rect 1981 4400 2097 4434
rect 1225 4385 1241 4400
rect 1293 4385 2097 4400
rect 2149 4385 2165 4437
rect 2217 4385 2233 4437
rect 2285 4385 2301 4437
rect 2353 4385 2369 4437
rect 2421 4434 2437 4437
rect 2421 4385 2437 4400
rect 2489 4385 2505 4437
rect 2557 4385 2573 4437
rect 2625 4385 2641 4437
rect 2693 4434 3076 4437
rect 2693 4400 2891 4434
rect 2925 4402 3076 4434
rect 2925 4400 3036 4402
rect 2693 4385 3036 4400
rect 380 4383 3036 4385
rect 380 4349 386 4383
rect 420 4373 3036 4383
rect 420 4361 697 4373
rect 420 4349 531 4361
rect 380 4327 531 4349
rect 565 4327 697 4361
rect 380 4321 697 4327
rect 749 4321 765 4373
rect 817 4321 833 4373
rect 885 4321 901 4373
rect 953 4321 969 4373
rect 1021 4361 1037 4373
rect 1021 4321 1037 4327
rect 1089 4321 1105 4373
rect 1157 4321 1173 4373
rect 1225 4361 1241 4373
rect 1293 4361 2097 4373
rect 1225 4327 1239 4361
rect 1293 4327 1475 4361
rect 1509 4327 1711 4361
rect 1745 4327 1947 4361
rect 1981 4327 2097 4361
rect 1225 4321 1241 4327
rect 1293 4321 2097 4327
rect 2149 4321 2165 4373
rect 2217 4321 2233 4373
rect 2285 4321 2301 4373
rect 2353 4321 2369 4373
rect 2421 4361 2437 4373
rect 2421 4321 2437 4327
rect 2489 4321 2505 4373
rect 2557 4321 2573 4373
rect 2625 4321 2641 4373
rect 2693 4368 3036 4373
rect 3070 4368 3076 4402
rect 2693 4361 3076 4368
rect 2693 4327 2891 4361
rect 2925 4330 3076 4361
rect 2925 4327 3036 4330
rect 2693 4321 3036 4327
rect 380 4311 3036 4321
rect 380 4277 386 4311
rect 420 4309 3036 4311
rect 420 4288 697 4309
rect 420 4277 531 4288
rect 380 4254 531 4277
rect 565 4257 697 4288
rect 749 4257 765 4309
rect 817 4257 833 4309
rect 885 4257 901 4309
rect 953 4257 969 4309
rect 1021 4288 1037 4309
rect 1089 4257 1105 4309
rect 1157 4257 1173 4309
rect 1225 4288 1241 4309
rect 1293 4288 2097 4309
rect 1225 4257 1239 4288
rect 1293 4257 1475 4288
rect 565 4254 767 4257
rect 801 4254 1003 4257
rect 1037 4254 1239 4257
rect 1273 4254 1475 4257
rect 1509 4254 1711 4288
rect 1745 4254 1947 4288
rect 1981 4257 2097 4288
rect 2149 4257 2165 4309
rect 2217 4257 2233 4309
rect 2285 4257 2301 4309
rect 2353 4257 2369 4309
rect 2421 4288 2437 4309
rect 2489 4257 2505 4309
rect 2557 4257 2573 4309
rect 2625 4257 2641 4309
rect 2693 4296 3036 4309
rect 3070 4296 3076 4330
rect 2693 4288 3076 4296
rect 2693 4257 2891 4288
rect 1981 4254 2183 4257
rect 2217 4254 2419 4257
rect 2453 4254 2655 4257
rect 2689 4254 2891 4257
rect 2925 4258 3076 4288
rect 2925 4254 3036 4258
rect 380 4245 3036 4254
rect 380 4239 697 4245
rect 380 4205 386 4239
rect 420 4215 697 4239
rect 420 4205 531 4215
rect 380 4181 531 4205
rect 565 4193 697 4215
rect 749 4193 765 4245
rect 817 4193 833 4245
rect 885 4193 901 4245
rect 953 4193 969 4245
rect 1021 4215 1037 4245
rect 1089 4193 1105 4245
rect 1157 4193 1173 4245
rect 1225 4215 1241 4245
rect 1293 4215 2097 4245
rect 1225 4193 1239 4215
rect 1293 4193 1475 4215
rect 565 4181 767 4193
rect 801 4181 1003 4193
rect 1037 4181 1239 4193
rect 1273 4181 1475 4193
rect 1509 4181 1711 4215
rect 1745 4181 1947 4215
rect 1981 4193 2097 4215
rect 2149 4193 2165 4245
rect 2217 4193 2233 4245
rect 2285 4193 2301 4245
rect 2353 4193 2369 4245
rect 2421 4215 2437 4245
rect 2489 4193 2505 4245
rect 2557 4193 2573 4245
rect 2625 4193 2641 4245
rect 2693 4224 3036 4245
rect 3070 4224 3076 4258
rect 2693 4215 3076 4224
rect 2693 4193 2891 4215
rect 1981 4181 2183 4193
rect 2217 4181 2419 4193
rect 2453 4181 2655 4193
rect 2689 4181 2891 4193
rect 2925 4186 3076 4215
rect 2925 4181 3036 4186
rect 380 4167 697 4181
rect 380 4133 386 4167
rect 420 4142 697 4167
rect 420 4133 531 4142
rect 380 4108 531 4133
rect 565 4129 697 4142
rect 749 4129 765 4181
rect 817 4129 833 4181
rect 885 4129 901 4181
rect 953 4129 969 4181
rect 1021 4142 1037 4181
rect 1089 4129 1105 4181
rect 1157 4129 1173 4181
rect 1225 4142 1241 4181
rect 1293 4142 2097 4181
rect 1225 4129 1239 4142
rect 1293 4129 1475 4142
rect 565 4117 767 4129
rect 801 4117 1003 4129
rect 1037 4117 1239 4129
rect 1273 4117 1475 4129
rect 565 4108 697 4117
rect 380 4095 697 4108
rect 380 4061 386 4095
rect 420 4069 697 4095
rect 420 4061 531 4069
rect 380 4035 531 4061
rect 565 4065 697 4069
rect 749 4065 765 4117
rect 817 4065 833 4117
rect 885 4065 901 4117
rect 953 4065 969 4117
rect 1021 4069 1037 4108
rect 1089 4065 1105 4117
rect 1157 4065 1173 4117
rect 1225 4108 1239 4117
rect 1293 4108 1475 4117
rect 1509 4108 1711 4142
rect 1745 4108 1947 4142
rect 1981 4129 2097 4142
rect 2149 4129 2165 4181
rect 2217 4129 2233 4181
rect 2285 4129 2301 4181
rect 2353 4129 2369 4181
rect 2421 4142 2437 4181
rect 2489 4129 2505 4181
rect 2557 4129 2573 4181
rect 2625 4129 2641 4181
rect 2693 4152 3036 4181
rect 3070 4152 3076 4186
rect 2693 4142 3076 4152
rect 2693 4129 2891 4142
rect 1981 4117 2183 4129
rect 2217 4117 2419 4129
rect 2453 4117 2655 4129
rect 2689 4117 2891 4129
rect 1981 4108 2097 4117
rect 1225 4069 1241 4108
rect 1293 4069 2097 4108
rect 1225 4065 1239 4069
rect 1293 4065 1475 4069
rect 565 4053 767 4065
rect 801 4053 1003 4065
rect 1037 4053 1239 4065
rect 1273 4053 1475 4065
rect 565 4035 697 4053
rect 380 4023 697 4035
rect 380 3989 386 4023
rect 420 4001 697 4023
rect 749 4001 765 4053
rect 817 4001 833 4053
rect 885 4001 901 4053
rect 953 4001 969 4053
rect 1021 4001 1037 4035
rect 1089 4001 1105 4053
rect 1157 4001 1173 4053
rect 1225 4035 1239 4053
rect 1293 4035 1475 4053
rect 1509 4035 1711 4069
rect 1745 4035 1947 4069
rect 1981 4065 2097 4069
rect 2149 4065 2165 4117
rect 2217 4065 2233 4117
rect 2285 4065 2301 4117
rect 2353 4065 2369 4117
rect 2421 4069 2437 4108
rect 2489 4065 2505 4117
rect 2557 4065 2573 4117
rect 2625 4065 2641 4117
rect 2693 4108 2891 4117
rect 2925 4114 3076 4142
rect 2925 4108 3036 4114
rect 2693 4080 3036 4108
rect 3070 4080 3076 4114
rect 2693 4069 3076 4080
rect 2693 4065 2891 4069
rect 1981 4053 2183 4065
rect 2217 4053 2419 4065
rect 2453 4053 2655 4065
rect 2689 4053 2891 4065
rect 1981 4035 2097 4053
rect 1225 4001 1241 4035
rect 1293 4001 2097 4035
rect 2149 4001 2165 4053
rect 2217 4001 2233 4053
rect 2285 4001 2301 4053
rect 2353 4001 2369 4053
rect 2421 4001 2437 4035
rect 2489 4001 2505 4053
rect 2557 4001 2573 4053
rect 2625 4001 2641 4053
rect 2693 4035 2891 4053
rect 2925 4042 3076 4069
rect 2925 4035 3036 4042
rect 2693 4008 3036 4035
rect 3070 4008 3076 4042
rect 2693 4001 3076 4008
rect 420 3996 3076 4001
rect 420 3989 531 3996
rect 380 3962 531 3989
rect 565 3989 767 3996
rect 801 3989 1003 3996
rect 1037 3989 1239 3996
rect 1273 3989 1475 3996
rect 565 3962 697 3989
rect 380 3951 697 3962
rect 380 3917 386 3951
rect 420 3937 697 3951
rect 749 3937 765 3989
rect 817 3937 833 3989
rect 885 3937 901 3989
rect 953 3937 969 3989
rect 1021 3937 1037 3962
rect 1089 3937 1105 3989
rect 1157 3937 1173 3989
rect 1225 3962 1239 3989
rect 1293 3962 1475 3989
rect 1509 3962 1711 3996
rect 1745 3962 1947 3996
rect 1981 3989 2183 3996
rect 2217 3989 2419 3996
rect 2453 3989 2655 3996
rect 2689 3989 2891 3996
rect 1981 3962 2097 3989
rect 1225 3937 1241 3962
rect 1293 3937 2097 3962
rect 2149 3937 2165 3989
rect 2217 3937 2233 3989
rect 2285 3937 2301 3989
rect 2353 3937 2369 3989
rect 2421 3937 2437 3962
rect 2489 3937 2505 3989
rect 2557 3937 2573 3989
rect 2625 3937 2641 3989
rect 2693 3962 2891 3989
rect 2925 3970 3076 3996
rect 2925 3962 3036 3970
rect 2693 3937 3036 3962
rect 420 3936 3036 3937
rect 3070 3936 3076 3970
rect 420 3925 3076 3936
rect 420 3922 697 3925
rect 420 3917 531 3922
rect 380 3888 531 3917
rect 565 3888 697 3922
rect 380 3879 697 3888
rect 380 3845 386 3879
rect 420 3873 697 3879
rect 749 3873 765 3925
rect 817 3873 833 3925
rect 885 3873 901 3925
rect 953 3873 969 3925
rect 1021 3922 1037 3925
rect 1021 3873 1037 3888
rect 1089 3873 1105 3925
rect 1157 3873 1173 3925
rect 1225 3922 1241 3925
rect 1293 3922 2097 3925
rect 1225 3888 1239 3922
rect 1293 3888 1475 3922
rect 1509 3888 1711 3922
rect 1745 3888 1947 3922
rect 1981 3888 2097 3922
rect 1225 3873 1241 3888
rect 1293 3873 2097 3888
rect 2149 3873 2165 3925
rect 2217 3873 2233 3925
rect 2285 3873 2301 3925
rect 2353 3873 2369 3925
rect 2421 3922 2437 3925
rect 2421 3873 2437 3888
rect 2489 3873 2505 3925
rect 2557 3873 2573 3925
rect 2625 3873 2641 3925
rect 2693 3922 3076 3925
rect 2693 3888 2891 3922
rect 2925 3898 3076 3922
rect 2925 3888 3036 3898
rect 2693 3873 3036 3888
rect 420 3864 3036 3873
rect 3070 3864 3076 3898
rect 420 3861 3076 3864
rect 420 3848 697 3861
rect 420 3845 531 3848
rect 380 3814 531 3845
rect 565 3814 697 3848
rect 380 3809 697 3814
rect 749 3809 765 3861
rect 817 3809 833 3861
rect 885 3809 901 3861
rect 953 3809 969 3861
rect 1021 3848 1037 3861
rect 1021 3809 1037 3814
rect 1089 3809 1105 3861
rect 1157 3809 1173 3861
rect 1225 3848 1241 3861
rect 1293 3848 2097 3861
rect 1225 3814 1239 3848
rect 1293 3814 1475 3848
rect 1509 3814 1711 3848
rect 1745 3814 1947 3848
rect 1981 3814 2097 3848
rect 1225 3809 1241 3814
rect 1293 3809 2097 3814
rect 2149 3809 2165 3861
rect 2217 3809 2233 3861
rect 2285 3809 2301 3861
rect 2353 3809 2369 3861
rect 2421 3848 2437 3861
rect 2421 3809 2437 3814
rect 2489 3809 2505 3861
rect 2557 3809 2573 3861
rect 2625 3809 2641 3861
rect 2693 3848 3076 3861
rect 2693 3814 2891 3848
rect 2925 3826 3076 3848
rect 2925 3814 3036 3826
rect 2693 3809 3036 3814
rect 380 3807 3036 3809
rect 380 3773 386 3807
rect 420 3797 3036 3807
rect 420 3774 697 3797
rect 420 3773 531 3774
rect 380 3740 531 3773
rect 565 3745 697 3774
rect 749 3745 765 3797
rect 817 3745 833 3797
rect 885 3745 901 3797
rect 953 3745 969 3797
rect 1021 3774 1037 3797
rect 1089 3745 1105 3797
rect 1157 3745 1173 3797
rect 1225 3774 1241 3797
rect 1293 3774 2097 3797
rect 1225 3745 1239 3774
rect 1293 3745 1475 3774
rect 565 3740 767 3745
rect 801 3740 1003 3745
rect 1037 3740 1239 3745
rect 1273 3740 1475 3745
rect 1509 3740 1711 3774
rect 1745 3740 1947 3774
rect 1981 3745 2097 3774
rect 2149 3745 2165 3797
rect 2217 3745 2233 3797
rect 2285 3745 2301 3797
rect 2353 3745 2369 3797
rect 2421 3774 2437 3797
rect 2489 3745 2505 3797
rect 2557 3745 2573 3797
rect 2625 3745 2641 3797
rect 2693 3792 3036 3797
rect 3070 3792 3076 3826
rect 2693 3774 3076 3792
rect 2693 3745 2891 3774
rect 1981 3740 2183 3745
rect 2217 3740 2419 3745
rect 2453 3740 2655 3745
rect 2689 3740 2891 3745
rect 2925 3754 3076 3774
rect 2925 3740 3036 3754
rect 380 3735 3036 3740
rect 380 3701 386 3735
rect 420 3733 3036 3735
rect 420 3701 697 3733
rect 380 3700 697 3701
rect 380 3666 531 3700
rect 565 3681 697 3700
rect 749 3681 765 3733
rect 817 3681 833 3733
rect 885 3681 901 3733
rect 953 3681 969 3733
rect 1021 3700 1037 3733
rect 1089 3681 1105 3733
rect 1157 3681 1173 3733
rect 1225 3700 1241 3733
rect 1293 3700 2097 3733
rect 1225 3681 1239 3700
rect 1293 3681 1475 3700
rect 565 3669 767 3681
rect 801 3669 1003 3681
rect 1037 3669 1239 3681
rect 1273 3669 1475 3681
rect 565 3666 697 3669
rect 380 3663 697 3666
rect 380 3629 386 3663
rect 420 3629 697 3663
rect 380 3626 697 3629
rect 380 3592 531 3626
rect 565 3617 697 3626
rect 749 3617 765 3669
rect 817 3617 833 3669
rect 885 3617 901 3669
rect 953 3617 969 3669
rect 1021 3626 1037 3666
rect 1089 3617 1105 3669
rect 1157 3617 1173 3669
rect 1225 3666 1239 3669
rect 1293 3666 1475 3669
rect 1509 3666 1711 3700
rect 1745 3666 1947 3700
rect 1981 3681 2097 3700
rect 2149 3681 2165 3733
rect 2217 3681 2233 3733
rect 2285 3681 2301 3733
rect 2353 3681 2369 3733
rect 2421 3700 2437 3733
rect 2489 3681 2505 3733
rect 2557 3681 2573 3733
rect 2625 3681 2641 3733
rect 2693 3720 3036 3733
rect 3070 3720 3076 3754
rect 2693 3700 3076 3720
rect 2693 3681 2891 3700
rect 1981 3669 2183 3681
rect 2217 3669 2419 3681
rect 2453 3669 2655 3681
rect 2689 3669 2891 3681
rect 1981 3666 2097 3669
rect 1225 3626 1241 3666
rect 1293 3626 2097 3666
rect 1225 3617 1239 3626
rect 1293 3617 1475 3626
rect 565 3605 767 3617
rect 801 3605 1003 3617
rect 1037 3605 1239 3617
rect 1273 3605 1475 3617
rect 565 3592 697 3605
rect 380 3591 697 3592
rect 380 3557 386 3591
rect 420 3557 697 3591
rect 380 3553 697 3557
rect 749 3553 765 3605
rect 817 3553 833 3605
rect 885 3553 901 3605
rect 953 3553 969 3605
rect 1021 3553 1037 3592
rect 1089 3553 1105 3605
rect 1157 3553 1173 3605
rect 1225 3592 1239 3605
rect 1293 3592 1475 3605
rect 1509 3592 1711 3626
rect 1745 3592 1947 3626
rect 1981 3617 2097 3626
rect 2149 3617 2165 3669
rect 2217 3617 2233 3669
rect 2285 3617 2301 3669
rect 2353 3617 2369 3669
rect 2421 3626 2437 3666
rect 2489 3617 2505 3669
rect 2557 3617 2573 3669
rect 2625 3617 2641 3669
rect 2693 3666 2891 3669
rect 2925 3682 3076 3700
rect 2925 3666 3036 3682
rect 2693 3648 3036 3666
rect 3070 3648 3076 3682
rect 2693 3626 3076 3648
rect 2693 3617 2891 3626
rect 1981 3605 2183 3617
rect 2217 3605 2419 3617
rect 2453 3605 2655 3617
rect 2689 3605 2891 3617
rect 1981 3592 2097 3605
rect 1225 3553 1241 3592
rect 1293 3553 2097 3592
rect 2149 3553 2165 3605
rect 2217 3553 2233 3605
rect 2285 3553 2301 3605
rect 2353 3553 2369 3605
rect 2421 3553 2437 3592
rect 2489 3553 2505 3605
rect 2557 3553 2573 3605
rect 2625 3553 2641 3605
rect 2693 3592 2891 3605
rect 2925 3610 3076 3626
rect 2925 3592 3036 3610
rect 2693 3576 3036 3592
rect 3070 3576 3076 3610
rect 2693 3553 3076 3576
rect 380 3552 3076 3553
rect 380 3519 531 3552
rect 380 3485 386 3519
rect 420 3518 531 3519
rect 565 3541 767 3552
rect 801 3541 1003 3552
rect 1037 3541 1239 3552
rect 1273 3541 1475 3552
rect 565 3518 697 3541
rect 420 3489 697 3518
rect 749 3489 765 3541
rect 817 3489 833 3541
rect 885 3489 901 3541
rect 953 3489 969 3541
rect 1021 3489 1037 3518
rect 1089 3489 1105 3541
rect 1157 3489 1173 3541
rect 1225 3518 1239 3541
rect 1293 3518 1475 3541
rect 1509 3518 1711 3552
rect 1745 3518 1947 3552
rect 1981 3541 2183 3552
rect 2217 3541 2419 3552
rect 2453 3541 2655 3552
rect 2689 3541 2891 3552
rect 1981 3518 2097 3541
rect 1225 3489 1241 3518
rect 1293 3489 2097 3518
rect 2149 3489 2165 3541
rect 2217 3489 2233 3541
rect 2285 3489 2301 3541
rect 2353 3489 2369 3541
rect 2421 3489 2437 3518
rect 2489 3489 2505 3541
rect 2557 3489 2573 3541
rect 2625 3489 2641 3541
rect 2693 3518 2891 3541
rect 2925 3538 3076 3552
rect 2925 3518 3036 3538
rect 2693 3504 3036 3518
rect 3070 3504 3076 3538
rect 2693 3489 3076 3504
rect 420 3485 3076 3489
rect 380 3478 3076 3485
rect 380 3447 531 3478
rect 380 3413 386 3447
rect 420 3444 531 3447
rect 565 3459 767 3478
rect 565 3444 590 3459
tri 590 3444 605 3459 nw
tri 727 3444 742 3459 ne
rect 742 3444 767 3459
rect 801 3459 1003 3478
rect 801 3444 826 3459
tri 826 3444 841 3459 nw
tri 963 3444 978 3459 ne
rect 978 3444 1003 3459
rect 1037 3459 1239 3478
rect 1037 3444 1062 3459
tri 1062 3444 1077 3459 nw
tri 1199 3444 1214 3459 ne
rect 1214 3444 1239 3459
rect 1273 3459 1475 3478
rect 1273 3444 1298 3459
tri 1298 3444 1313 3459 nw
tri 1435 3444 1450 3459 ne
rect 1450 3444 1475 3459
rect 1509 3459 1711 3478
rect 1509 3444 1534 3459
tri 1534 3444 1549 3459 nw
tri 1671 3444 1686 3459 ne
rect 1686 3444 1711 3459
rect 1745 3459 1947 3478
rect 1745 3444 1770 3459
tri 1770 3444 1785 3459 nw
tri 1907 3444 1922 3459 ne
rect 1922 3444 1947 3459
rect 1981 3459 2183 3478
rect 1981 3444 2006 3459
tri 2006 3444 2021 3459 nw
tri 2143 3444 2158 3459 ne
rect 2158 3444 2183 3459
rect 2217 3459 2419 3478
rect 2217 3444 2242 3459
tri 2242 3444 2257 3459 nw
tri 2379 3444 2394 3459 ne
rect 2394 3444 2419 3459
rect 2453 3459 2655 3478
rect 2453 3444 2478 3459
tri 2478 3444 2493 3459 nw
tri 2615 3444 2630 3459 ne
rect 2630 3444 2655 3459
rect 2689 3459 2891 3478
rect 2689 3444 2714 3459
tri 2714 3444 2729 3459 nw
tri 2851 3444 2866 3459 ne
rect 2866 3444 2891 3459
rect 2925 3466 3076 3478
rect 2925 3444 3036 3466
rect 420 3432 578 3444
tri 578 3432 590 3444 nw
tri 742 3432 754 3444 ne
rect 754 3432 814 3444
tri 814 3432 826 3444 nw
tri 978 3432 990 3444 ne
rect 990 3432 1050 3444
tri 1050 3432 1062 3444 nw
tri 1214 3432 1226 3444 ne
rect 1226 3432 1286 3444
tri 1286 3432 1298 3444 nw
tri 1450 3432 1462 3444 ne
rect 1462 3432 1522 3444
tri 1522 3432 1534 3444 nw
tri 1686 3432 1698 3444 ne
rect 1698 3432 1758 3444
tri 1758 3432 1770 3444 nw
tri 1922 3432 1934 3444 ne
rect 1934 3432 1994 3444
tri 1994 3432 2006 3444 nw
tri 2158 3432 2170 3444 ne
rect 2170 3432 2230 3444
tri 2230 3432 2242 3444 nw
tri 2394 3432 2406 3444 ne
rect 2406 3432 2466 3444
tri 2466 3432 2478 3444 nw
tri 2630 3432 2642 3444 ne
rect 2642 3432 2702 3444
tri 2702 3432 2714 3444 nw
tri 2866 3432 2878 3444 ne
rect 2878 3432 3036 3444
rect 3070 3432 3076 3466
rect 420 3413 571 3432
tri 571 3425 578 3432 nw
tri 754 3425 761 3432 ne
rect 380 3404 571 3413
rect 380 3375 531 3404
rect 380 3341 386 3375
rect 420 3370 531 3375
rect 565 3370 571 3404
rect 420 3341 571 3370
rect 380 3330 571 3341
rect 380 3303 531 3330
rect 380 3269 386 3303
rect 420 3296 531 3303
rect 565 3296 571 3330
rect 420 3269 571 3296
rect 380 3256 571 3269
rect 380 3231 531 3256
rect 380 3197 386 3231
rect 420 3222 531 3231
rect 565 3222 571 3256
rect 420 3197 571 3222
rect 380 3182 571 3197
rect 380 3159 531 3182
rect 380 3125 386 3159
rect 420 3148 531 3159
rect 565 3148 571 3182
rect 420 3125 571 3148
rect 380 3108 571 3125
rect 380 3087 531 3108
rect 380 3053 386 3087
rect 420 3074 531 3087
rect 565 3074 571 3108
rect 420 3053 571 3074
rect 380 3034 571 3053
rect 380 3015 531 3034
rect 380 2981 386 3015
rect 420 3000 531 3015
rect 565 3000 571 3034
rect 420 2981 571 3000
rect 380 2960 571 2981
rect 380 2943 531 2960
rect 380 2909 386 2943
rect 420 2926 531 2943
rect 565 2926 571 2960
rect 420 2909 571 2926
rect 761 3404 807 3432
tri 807 3425 814 3432 nw
tri 990 3425 997 3432 ne
rect 761 3370 767 3404
rect 801 3370 807 3404
rect 761 3330 807 3370
rect 761 3296 767 3330
rect 801 3296 807 3330
rect 761 3256 807 3296
rect 761 3222 767 3256
rect 801 3222 807 3256
rect 761 3182 807 3222
rect 761 3148 767 3182
rect 801 3148 807 3182
rect 761 3108 807 3148
rect 761 3074 767 3108
rect 801 3074 807 3108
rect 761 3034 807 3074
rect 761 3000 767 3034
rect 801 3000 807 3034
rect 761 2960 807 3000
rect 761 2926 767 2960
rect 801 2926 807 2960
rect 761 2914 807 2926
rect 997 3404 1043 3432
tri 1043 3425 1050 3432 nw
tri 1226 3425 1233 3432 ne
rect 997 3370 1003 3404
rect 1037 3370 1043 3404
rect 997 3330 1043 3370
rect 997 3296 1003 3330
rect 1037 3296 1043 3330
rect 997 3256 1043 3296
rect 997 3222 1003 3256
rect 1037 3222 1043 3256
rect 997 3182 1043 3222
rect 997 3148 1003 3182
rect 1037 3148 1043 3182
rect 997 3108 1043 3148
rect 997 3074 1003 3108
rect 1037 3074 1043 3108
rect 997 3034 1043 3074
rect 997 3000 1003 3034
rect 1037 3000 1043 3034
rect 997 2960 1043 3000
rect 997 2926 1003 2960
rect 1037 2926 1043 2960
rect 997 2914 1043 2926
rect 1233 3404 1279 3432
tri 1279 3425 1286 3432 nw
tri 1462 3425 1469 3432 ne
rect 1233 3370 1239 3404
rect 1273 3370 1279 3404
rect 1233 3330 1279 3370
rect 1233 3296 1239 3330
rect 1273 3296 1279 3330
rect 1233 3256 1279 3296
rect 1233 3222 1239 3256
rect 1273 3222 1279 3256
rect 1233 3182 1279 3222
rect 1233 3148 1239 3182
rect 1273 3148 1279 3182
rect 1233 3108 1279 3148
rect 1233 3074 1239 3108
rect 1273 3074 1279 3108
rect 1233 3034 1279 3074
rect 1233 3000 1239 3034
rect 1273 3000 1279 3034
rect 1233 2960 1279 3000
rect 1233 2926 1239 2960
rect 1273 2926 1279 2960
rect 1233 2914 1279 2926
rect 1469 3404 1515 3432
tri 1515 3425 1522 3432 nw
tri 1698 3425 1705 3432 ne
rect 1469 3370 1475 3404
rect 1509 3370 1515 3404
rect 1469 3330 1515 3370
rect 1469 3296 1475 3330
rect 1509 3296 1515 3330
rect 1469 3256 1515 3296
rect 1469 3222 1475 3256
rect 1509 3222 1515 3256
rect 1469 3182 1515 3222
rect 1469 3148 1475 3182
rect 1509 3148 1515 3182
rect 1469 3108 1515 3148
rect 1469 3074 1475 3108
rect 1509 3074 1515 3108
rect 1469 3034 1515 3074
rect 1469 3000 1475 3034
rect 1509 3000 1515 3034
rect 1469 2960 1515 3000
rect 1469 2926 1475 2960
rect 1509 2926 1515 2960
rect 1469 2914 1515 2926
rect 1705 3404 1751 3432
tri 1751 3425 1758 3432 nw
tri 1934 3425 1941 3432 ne
rect 1705 3370 1711 3404
rect 1745 3370 1751 3404
rect 1705 3330 1751 3370
rect 1705 3296 1711 3330
rect 1745 3296 1751 3330
rect 1705 3256 1751 3296
rect 1705 3222 1711 3256
rect 1745 3222 1751 3256
rect 1705 3182 1751 3222
rect 1705 3148 1711 3182
rect 1745 3148 1751 3182
rect 1705 3108 1751 3148
rect 1705 3074 1711 3108
rect 1745 3074 1751 3108
rect 1705 3034 1751 3074
rect 1705 3000 1711 3034
rect 1745 3000 1751 3034
rect 1705 2960 1751 3000
rect 1705 2926 1711 2960
rect 1745 2926 1751 2960
rect 1705 2914 1751 2926
rect 1941 3404 1987 3432
tri 1987 3425 1994 3432 nw
tri 2170 3425 2177 3432 ne
rect 1941 3370 1947 3404
rect 1981 3370 1987 3404
rect 1941 3330 1987 3370
rect 1941 3296 1947 3330
rect 1981 3296 1987 3330
rect 1941 3256 1987 3296
rect 1941 3222 1947 3256
rect 1981 3222 1987 3256
rect 1941 3182 1987 3222
rect 1941 3148 1947 3182
rect 1981 3148 1987 3182
rect 1941 3108 1987 3148
rect 1941 3074 1947 3108
rect 1981 3074 1987 3108
rect 1941 3034 1987 3074
rect 1941 3000 1947 3034
rect 1981 3000 1987 3034
rect 1941 2960 1987 3000
rect 1941 2926 1947 2960
rect 1981 2926 1987 2960
rect 1941 2914 1987 2926
rect 2177 3404 2223 3432
tri 2223 3425 2230 3432 nw
tri 2406 3425 2413 3432 ne
rect 2177 3370 2183 3404
rect 2217 3370 2223 3404
rect 2177 3330 2223 3370
rect 2177 3296 2183 3330
rect 2217 3296 2223 3330
rect 2177 3256 2223 3296
rect 2177 3222 2183 3256
rect 2217 3222 2223 3256
rect 2177 3182 2223 3222
rect 2177 3148 2183 3182
rect 2217 3148 2223 3182
rect 2177 3108 2223 3148
rect 2177 3074 2183 3108
rect 2217 3074 2223 3108
rect 2177 3034 2223 3074
rect 2177 3000 2183 3034
rect 2217 3000 2223 3034
rect 2177 2960 2223 3000
rect 2177 2926 2183 2960
rect 2217 2926 2223 2960
rect 2177 2914 2223 2926
rect 2413 3404 2459 3432
tri 2459 3425 2466 3432 nw
tri 2642 3425 2649 3432 ne
rect 2413 3370 2419 3404
rect 2453 3370 2459 3404
rect 2413 3330 2459 3370
rect 2413 3296 2419 3330
rect 2453 3296 2459 3330
rect 2413 3256 2459 3296
rect 2413 3222 2419 3256
rect 2453 3222 2459 3256
rect 2413 3182 2459 3222
rect 2413 3148 2419 3182
rect 2453 3148 2459 3182
rect 2413 3108 2459 3148
rect 2413 3074 2419 3108
rect 2453 3074 2459 3108
rect 2413 3034 2459 3074
rect 2413 3000 2419 3034
rect 2453 3000 2459 3034
rect 2413 2960 2459 3000
rect 2413 2926 2419 2960
rect 2453 2926 2459 2960
rect 2413 2914 2459 2926
rect 2649 3404 2695 3432
tri 2695 3425 2702 3432 nw
tri 2878 3425 2885 3432 ne
rect 2649 3370 2655 3404
rect 2689 3370 2695 3404
rect 2649 3330 2695 3370
rect 2649 3296 2655 3330
rect 2689 3296 2695 3330
rect 2649 3256 2695 3296
rect 2649 3222 2655 3256
rect 2689 3222 2695 3256
rect 2649 3182 2695 3222
rect 2649 3148 2655 3182
rect 2689 3148 2695 3182
rect 2649 3108 2695 3148
rect 2649 3074 2655 3108
rect 2689 3074 2695 3108
rect 2649 3034 2695 3074
rect 2649 3000 2655 3034
rect 2689 3000 2695 3034
rect 2649 2960 2695 3000
rect 2649 2926 2655 2960
rect 2689 2926 2695 2960
rect 2649 2914 2695 2926
rect 2885 3404 3076 3432
rect 2885 3370 2891 3404
rect 2925 3394 3076 3404
rect 2925 3370 3036 3394
rect 2885 3360 3036 3370
rect 3070 3360 3076 3394
rect 2885 3330 3076 3360
rect 2885 3296 2891 3330
rect 2925 3322 3076 3330
rect 2925 3296 3036 3322
rect 2885 3288 3036 3296
rect 3070 3288 3076 3322
rect 2885 3256 3076 3288
rect 2885 3222 2891 3256
rect 2925 3250 3076 3256
rect 2925 3222 3036 3250
rect 2885 3216 3036 3222
rect 3070 3216 3076 3250
rect 2885 3182 3076 3216
rect 2885 3148 2891 3182
rect 2925 3178 3076 3182
rect 2925 3148 3036 3178
rect 2885 3144 3036 3148
rect 3070 3144 3076 3178
rect 2885 3108 3076 3144
rect 2885 3074 2891 3108
rect 2925 3106 3076 3108
rect 2925 3074 3036 3106
rect 2885 3072 3036 3074
rect 3070 3072 3076 3106
rect 2885 3034 3076 3072
rect 2885 3000 2891 3034
rect 2925 3000 3036 3034
rect 3070 3000 3076 3034
rect 2885 2962 3076 3000
rect 2885 2960 3036 2962
rect 2885 2926 2891 2960
rect 2925 2928 3036 2960
rect 3070 2928 3076 2962
rect 2925 2926 3076 2928
rect 380 2871 571 2909
rect 380 2837 386 2871
rect 420 2837 571 2871
rect 2885 2890 3076 2926
rect 2885 2856 3036 2890
rect 3070 2856 3076 2890
rect 380 2799 571 2837
rect 613 2844 1501 2853
rect 1553 2844 1569 2853
rect 1621 2844 1636 2853
rect 1688 2844 1703 2853
rect 1755 2844 1770 2853
rect 1822 2844 1837 2853
rect 1889 2844 2830 2853
rect 613 2810 625 2844
rect 659 2810 700 2844
rect 734 2810 775 2844
rect 809 2810 850 2844
rect 884 2810 925 2844
rect 959 2810 1000 2844
rect 1034 2810 1075 2844
rect 1109 2810 1150 2844
rect 1184 2810 1225 2844
rect 1259 2810 1300 2844
rect 1334 2810 1375 2844
rect 1409 2810 1450 2844
rect 1484 2810 1501 2844
rect 1559 2810 1569 2844
rect 1634 2810 1636 2844
rect 1889 2810 1896 2844
rect 1930 2810 1970 2844
rect 2004 2810 2044 2844
rect 2078 2810 2118 2844
rect 2152 2810 2192 2844
rect 2226 2810 2266 2844
rect 2300 2810 2340 2844
rect 2374 2810 2414 2844
rect 2448 2810 2488 2844
rect 2522 2810 2562 2844
rect 2596 2810 2636 2844
rect 2670 2810 2710 2844
rect 2744 2810 2784 2844
rect 2818 2810 2830 2844
rect 613 2801 1501 2810
rect 1553 2801 1569 2810
rect 1621 2801 1636 2810
rect 1688 2801 1703 2810
rect 1755 2801 1770 2810
rect 1822 2801 1837 2810
rect 1889 2801 2830 2810
rect 2885 2818 3076 2856
rect 380 2765 386 2799
rect 420 2765 571 2799
rect 380 2727 571 2765
rect 2885 2784 3036 2818
rect 3070 2784 3076 2818
rect 2885 2746 3076 2784
rect 380 2693 386 2727
rect 420 2720 571 2727
rect 420 2693 531 2720
rect 380 2686 531 2693
rect 565 2686 571 2720
rect 380 2655 571 2686
rect 380 2621 386 2655
rect 420 2647 571 2655
rect 420 2621 531 2647
rect 380 2613 531 2621
rect 565 2613 571 2647
rect 380 2583 571 2613
rect 380 2549 386 2583
rect 420 2574 571 2583
rect 420 2549 531 2574
rect 380 2540 531 2549
rect 565 2540 571 2574
rect 380 2511 571 2540
rect 380 2477 386 2511
rect 420 2501 571 2511
rect 420 2477 531 2501
rect 380 2467 531 2477
rect 565 2467 571 2501
rect 380 2439 571 2467
rect 380 2405 386 2439
rect 420 2428 571 2439
rect 420 2405 531 2428
rect 380 2394 531 2405
rect 565 2394 571 2428
rect 380 2367 571 2394
rect 380 2333 386 2367
rect 420 2355 571 2367
rect 420 2333 531 2355
rect 380 2321 531 2333
rect 565 2321 571 2355
rect 380 2295 571 2321
rect 761 2720 807 2732
rect 761 2686 767 2720
rect 801 2686 807 2720
rect 761 2647 807 2686
rect 761 2613 767 2647
rect 801 2613 807 2647
rect 761 2574 807 2613
rect 761 2540 767 2574
rect 801 2540 807 2574
rect 761 2501 807 2540
rect 761 2467 767 2501
rect 801 2467 807 2501
rect 761 2428 807 2467
rect 761 2394 767 2428
rect 801 2394 807 2428
rect 761 2355 807 2394
rect 761 2321 767 2355
rect 801 2321 807 2355
rect 380 2261 386 2295
rect 420 2282 571 2295
tri 571 2282 590 2301 sw
tri 742 2282 761 2301 se
rect 761 2282 807 2321
rect 997 2720 1043 2732
rect 997 2686 1003 2720
rect 1037 2686 1043 2720
rect 997 2647 1043 2686
rect 997 2613 1003 2647
rect 1037 2613 1043 2647
rect 997 2574 1043 2613
rect 997 2540 1003 2574
rect 1037 2540 1043 2574
rect 997 2501 1043 2540
rect 997 2467 1003 2501
rect 1037 2467 1043 2501
rect 997 2428 1043 2467
rect 997 2394 1003 2428
rect 1037 2394 1043 2428
rect 997 2355 1043 2394
rect 997 2321 1003 2355
rect 1037 2321 1043 2355
tri 807 2282 826 2301 sw
tri 978 2282 997 2301 se
rect 997 2282 1043 2321
rect 1233 2720 1279 2732
rect 1233 2686 1239 2720
rect 1273 2686 1279 2720
rect 1233 2647 1279 2686
rect 1233 2613 1239 2647
rect 1273 2613 1279 2647
rect 1233 2574 1279 2613
rect 1233 2540 1239 2574
rect 1273 2540 1279 2574
rect 1233 2501 1279 2540
rect 1233 2467 1239 2501
rect 1273 2467 1279 2501
rect 1233 2428 1279 2467
rect 1233 2394 1239 2428
rect 1273 2394 1279 2428
rect 1233 2355 1279 2394
rect 1233 2321 1239 2355
rect 1273 2321 1279 2355
tri 1043 2282 1062 2301 sw
tri 1214 2282 1233 2301 se
rect 1233 2282 1279 2321
rect 1469 2720 1515 2732
rect 1469 2686 1475 2720
rect 1509 2686 1515 2720
rect 1469 2647 1515 2686
rect 1469 2613 1475 2647
rect 1509 2613 1515 2647
rect 1469 2574 1515 2613
rect 1469 2540 1475 2574
rect 1509 2540 1515 2574
rect 1469 2501 1515 2540
rect 1469 2467 1475 2501
rect 1509 2467 1515 2501
rect 1469 2428 1515 2467
rect 1469 2394 1475 2428
rect 1509 2394 1515 2428
rect 1469 2355 1515 2394
rect 1469 2321 1475 2355
rect 1509 2321 1515 2355
tri 1279 2282 1298 2301 sw
tri 1450 2282 1469 2301 se
rect 1469 2282 1515 2321
rect 1705 2720 1751 2732
rect 1705 2686 1711 2720
rect 1745 2686 1751 2720
rect 1705 2647 1751 2686
rect 1705 2613 1711 2647
rect 1745 2613 1751 2647
rect 1705 2574 1751 2613
rect 1705 2540 1711 2574
rect 1745 2540 1751 2574
rect 1705 2501 1751 2540
rect 1705 2467 1711 2501
rect 1745 2467 1751 2501
rect 1705 2428 1751 2467
rect 1705 2394 1711 2428
rect 1745 2394 1751 2428
rect 1705 2355 1751 2394
rect 1705 2321 1711 2355
rect 1745 2321 1751 2355
tri 1515 2282 1534 2301 sw
tri 1686 2282 1705 2301 se
rect 1705 2282 1751 2321
rect 1941 2720 1987 2732
rect 1941 2686 1947 2720
rect 1981 2686 1987 2720
rect 1941 2647 1987 2686
rect 1941 2613 1947 2647
rect 1981 2613 1987 2647
rect 1941 2574 1987 2613
rect 1941 2540 1947 2574
rect 1981 2540 1987 2574
rect 1941 2501 1987 2540
rect 1941 2467 1947 2501
rect 1981 2467 1987 2501
rect 1941 2428 1987 2467
rect 1941 2394 1947 2428
rect 1981 2394 1987 2428
rect 1941 2355 1987 2394
rect 1941 2321 1947 2355
rect 1981 2321 1987 2355
tri 1751 2282 1770 2301 sw
tri 1922 2282 1941 2301 se
rect 1941 2282 1987 2321
rect 2177 2720 2223 2732
rect 2177 2686 2183 2720
rect 2217 2686 2223 2720
rect 2177 2647 2223 2686
rect 2177 2613 2183 2647
rect 2217 2613 2223 2647
rect 2177 2574 2223 2613
rect 2177 2540 2183 2574
rect 2217 2540 2223 2574
rect 2177 2501 2223 2540
rect 2177 2467 2183 2501
rect 2217 2467 2223 2501
rect 2177 2428 2223 2467
rect 2177 2394 2183 2428
rect 2217 2394 2223 2428
rect 2177 2355 2223 2394
rect 2177 2321 2183 2355
rect 2217 2321 2223 2355
tri 1987 2282 2006 2301 sw
tri 2158 2282 2177 2301 se
rect 2177 2282 2223 2321
rect 2413 2720 2459 2732
rect 2413 2686 2419 2720
rect 2453 2686 2459 2720
rect 2413 2647 2459 2686
rect 2413 2613 2419 2647
rect 2453 2613 2459 2647
rect 2413 2574 2459 2613
rect 2413 2540 2419 2574
rect 2453 2540 2459 2574
rect 2413 2501 2459 2540
rect 2413 2467 2419 2501
rect 2453 2467 2459 2501
rect 2413 2428 2459 2467
rect 2413 2394 2419 2428
rect 2453 2394 2459 2428
rect 2413 2355 2459 2394
rect 2413 2321 2419 2355
rect 2453 2321 2459 2355
tri 2223 2282 2242 2301 sw
tri 2394 2282 2413 2301 se
rect 2413 2282 2459 2321
rect 2649 2720 2695 2732
rect 2649 2686 2655 2720
rect 2689 2686 2695 2720
rect 2649 2647 2695 2686
rect 2649 2613 2655 2647
rect 2689 2613 2695 2647
rect 2649 2574 2695 2613
rect 2649 2540 2655 2574
rect 2689 2540 2695 2574
rect 2649 2501 2695 2540
rect 2649 2467 2655 2501
rect 2689 2467 2695 2501
rect 2649 2428 2695 2467
rect 2649 2394 2655 2428
rect 2689 2394 2695 2428
rect 2649 2355 2695 2394
rect 2649 2321 2655 2355
rect 2689 2321 2695 2355
tri 2459 2282 2478 2301 sw
tri 2630 2282 2649 2301 se
rect 2649 2282 2695 2321
rect 2885 2712 3036 2746
rect 3070 2712 3076 2746
rect 2885 2678 2891 2712
rect 2925 2678 3076 2712
rect 2885 2674 3076 2678
rect 2885 2640 3036 2674
rect 3070 2640 3076 2674
rect 2885 2639 3076 2640
rect 2885 2605 2891 2639
rect 2925 2605 3076 2639
rect 2885 2602 3076 2605
rect 2885 2568 3036 2602
rect 3070 2568 3076 2602
rect 2885 2566 3076 2568
rect 2885 2532 2891 2566
rect 2925 2532 3076 2566
rect 2885 2530 3076 2532
rect 2885 2496 3036 2530
rect 3070 2496 3076 2530
rect 2885 2493 3076 2496
rect 2885 2459 2891 2493
rect 2925 2459 3076 2493
rect 2885 2458 3076 2459
rect 2885 2424 3036 2458
rect 3070 2424 3076 2458
rect 2885 2420 3076 2424
rect 2885 2386 2891 2420
rect 2925 2386 3076 2420
rect 2885 2352 3036 2386
rect 3070 2352 3076 2386
rect 2885 2347 3076 2352
rect 2885 2313 2891 2347
rect 2925 2314 3076 2347
rect 2925 2313 3036 2314
rect 420 2261 531 2282
rect 380 2248 531 2261
rect 565 2267 590 2282
tri 590 2267 605 2282 sw
tri 727 2267 742 2282 se
rect 742 2267 767 2282
rect 565 2248 767 2267
rect 801 2267 826 2282
tri 826 2267 841 2282 sw
tri 963 2267 978 2282 se
rect 978 2267 1003 2282
rect 801 2248 1003 2267
rect 1037 2267 1062 2282
tri 1062 2267 1077 2282 sw
tri 1199 2267 1214 2282 se
rect 1214 2267 1239 2282
rect 1037 2248 1239 2267
rect 1273 2267 1298 2282
tri 1298 2267 1313 2282 sw
tri 1435 2267 1450 2282 se
rect 1450 2267 1475 2282
rect 1273 2248 1475 2267
rect 1509 2267 1534 2282
tri 1534 2267 1549 2282 sw
tri 1671 2267 1686 2282 se
rect 1686 2267 1711 2282
rect 1509 2248 1711 2267
rect 1745 2267 1770 2282
tri 1770 2267 1785 2282 sw
tri 1907 2267 1922 2282 se
rect 1922 2267 1947 2282
rect 1745 2248 1947 2267
rect 1981 2267 2006 2282
tri 2006 2267 2021 2282 sw
tri 2143 2267 2158 2282 se
rect 2158 2267 2183 2282
rect 1981 2248 2183 2267
rect 2217 2267 2242 2282
tri 2242 2267 2257 2282 sw
tri 2379 2267 2394 2282 se
rect 2394 2267 2419 2282
rect 2217 2248 2419 2267
rect 2453 2267 2478 2282
tri 2478 2267 2493 2282 sw
tri 2615 2267 2630 2282 se
rect 2630 2267 2655 2282
rect 2453 2248 2655 2267
rect 2689 2280 2695 2282
tri 2695 2280 2716 2301 sw
tri 2864 2280 2885 2301 se
rect 2885 2280 3036 2313
rect 3070 2280 3076 2314
rect 2689 2276 2716 2280
tri 2716 2276 2720 2280 sw
tri 2860 2276 2864 2280 se
rect 2864 2276 3076 2280
rect 2689 2274 2720 2276
tri 2720 2274 2722 2276 sw
tri 2858 2274 2860 2276 se
rect 2860 2274 3076 2276
rect 2689 2267 2722 2274
tri 2722 2267 2729 2274 sw
tri 2851 2267 2858 2274 se
rect 2858 2267 2891 2274
rect 2689 2248 2891 2267
rect 380 2243 2891 2248
rect 380 2223 697 2243
rect 380 2189 386 2223
rect 420 2209 697 2223
rect 420 2189 531 2209
rect 380 2175 531 2189
rect 565 2191 697 2209
rect 749 2191 765 2243
rect 817 2191 833 2243
rect 885 2191 901 2243
rect 953 2191 969 2243
rect 1021 2209 1037 2243
rect 1089 2191 1105 2243
rect 1157 2191 1173 2243
rect 1225 2209 1241 2243
rect 1293 2209 2097 2243
rect 1225 2191 1239 2209
rect 1293 2191 1475 2209
rect 565 2179 767 2191
rect 801 2179 1003 2191
rect 1037 2179 1239 2191
rect 1273 2179 1475 2191
rect 565 2175 697 2179
rect 380 2151 697 2175
rect 380 2117 386 2151
rect 420 2136 697 2151
rect 420 2117 531 2136
rect 380 2102 531 2117
rect 565 2127 697 2136
rect 749 2127 765 2179
rect 817 2127 833 2179
rect 885 2127 901 2179
rect 953 2127 969 2179
rect 1021 2136 1037 2175
rect 1089 2127 1105 2179
rect 1157 2127 1173 2179
rect 1225 2175 1239 2179
rect 1293 2175 1475 2179
rect 1509 2175 1711 2209
rect 1745 2175 1947 2209
rect 1981 2191 2097 2209
rect 2149 2191 2165 2243
rect 2217 2191 2233 2243
rect 2285 2191 2301 2243
rect 2353 2191 2369 2243
rect 2421 2209 2437 2243
rect 2489 2191 2505 2243
rect 2557 2191 2573 2243
rect 2625 2191 2641 2243
rect 2693 2240 2891 2243
rect 2925 2242 3076 2274
rect 2925 2240 3036 2242
rect 2693 2208 3036 2240
rect 3070 2208 3076 2242
rect 2693 2201 3076 2208
rect 2693 2191 2891 2201
rect 1981 2179 2183 2191
rect 2217 2179 2419 2191
rect 2453 2179 2655 2191
rect 2689 2179 2891 2191
rect 1981 2175 2097 2179
rect 1225 2136 1241 2175
rect 1293 2136 2097 2175
rect 1225 2127 1239 2136
rect 1293 2127 1475 2136
rect 565 2115 767 2127
rect 801 2115 1003 2127
rect 1037 2115 1239 2127
rect 1273 2115 1475 2127
rect 565 2102 697 2115
rect 380 2079 697 2102
rect 380 2045 386 2079
rect 420 2063 697 2079
rect 749 2063 765 2115
rect 817 2063 833 2115
rect 885 2063 901 2115
rect 953 2063 969 2115
rect 1021 2063 1037 2102
rect 1089 2063 1105 2115
rect 1157 2063 1173 2115
rect 1225 2102 1239 2115
rect 1293 2102 1475 2115
rect 1509 2102 1711 2136
rect 1745 2102 1947 2136
rect 1981 2127 2097 2136
rect 2149 2127 2165 2179
rect 2217 2127 2233 2179
rect 2285 2127 2301 2179
rect 2353 2127 2369 2179
rect 2421 2136 2437 2175
rect 2489 2127 2505 2179
rect 2557 2127 2573 2179
rect 2625 2127 2641 2179
rect 2693 2167 2891 2179
rect 2925 2170 3076 2201
rect 2925 2167 3036 2170
rect 2693 2136 3036 2167
rect 3070 2136 3076 2170
rect 2693 2128 3076 2136
rect 2693 2127 2891 2128
rect 1981 2115 2183 2127
rect 2217 2115 2419 2127
rect 2453 2115 2655 2127
rect 2689 2115 2891 2127
rect 1981 2102 2097 2115
rect 1225 2063 1241 2102
rect 1293 2063 2097 2102
rect 2149 2063 2165 2115
rect 2217 2063 2233 2115
rect 2285 2063 2301 2115
rect 2353 2063 2369 2115
rect 2421 2063 2437 2102
rect 2489 2063 2505 2115
rect 2557 2063 2573 2115
rect 2625 2063 2641 2115
rect 2693 2094 2891 2115
rect 2925 2098 3076 2128
rect 2925 2094 3036 2098
rect 2693 2064 3036 2094
rect 3070 2064 3076 2098
rect 2693 2063 3076 2064
rect 420 2045 531 2063
rect 380 2029 531 2045
rect 565 2051 767 2063
rect 801 2051 1003 2063
rect 1037 2051 1239 2063
rect 1273 2051 1475 2063
rect 565 2029 697 2051
rect 380 2007 697 2029
rect 380 1973 386 2007
rect 420 1999 697 2007
rect 749 1999 765 2051
rect 817 1999 833 2051
rect 885 1999 901 2051
rect 953 1999 969 2051
rect 1021 1999 1037 2029
rect 1089 1999 1105 2051
rect 1157 1999 1173 2051
rect 1225 2029 1239 2051
rect 1293 2029 1475 2051
rect 1509 2029 1711 2063
rect 1745 2029 1947 2063
rect 1981 2051 2183 2063
rect 2217 2051 2419 2063
rect 2453 2051 2655 2063
rect 2689 2055 3076 2063
rect 2689 2051 2891 2055
rect 1981 2029 2097 2051
rect 1225 1999 1241 2029
rect 1293 1999 2097 2029
rect 2149 1999 2165 2051
rect 2217 1999 2233 2051
rect 2285 1999 2301 2051
rect 2353 1999 2369 2051
rect 2421 1999 2437 2029
rect 2489 1999 2505 2051
rect 2557 1999 2573 2051
rect 2625 1999 2641 2051
rect 2693 2021 2891 2051
rect 2925 2026 3076 2055
rect 2925 2021 3036 2026
rect 2693 1999 3036 2021
rect 420 1992 3036 1999
rect 3070 1992 3076 2026
rect 420 1990 3076 1992
rect 420 1973 531 1990
rect 380 1956 531 1973
rect 565 1987 767 1990
rect 801 1987 1003 1990
rect 1037 1987 1239 1990
rect 1273 1987 1475 1990
rect 565 1956 697 1987
rect 380 1935 697 1956
rect 749 1935 765 1987
rect 817 1935 833 1987
rect 885 1935 901 1987
rect 953 1935 969 1987
rect 1021 1935 1037 1956
rect 1089 1935 1105 1987
rect 1157 1935 1173 1987
rect 1225 1956 1239 1987
rect 1293 1956 1475 1987
rect 1509 1956 1711 1990
rect 1745 1956 1947 1990
rect 1981 1987 2183 1990
rect 2217 1987 2419 1990
rect 2453 1987 2655 1990
rect 2689 1987 3076 1990
rect 1981 1956 2097 1987
rect 1225 1935 1241 1956
rect 1293 1935 2097 1956
rect 2149 1935 2165 1987
rect 2217 1935 2233 1987
rect 2285 1935 2301 1987
rect 2353 1935 2369 1987
rect 2421 1935 2437 1956
rect 2489 1935 2505 1987
rect 2557 1935 2573 1987
rect 2625 1935 2641 1987
rect 2693 1982 3076 1987
rect 2693 1948 2891 1982
rect 2925 1953 3076 1982
rect 2925 1948 3036 1953
rect 2693 1935 3036 1948
rect 380 1901 386 1935
rect 420 1923 3036 1935
rect 420 1917 697 1923
rect 420 1901 531 1917
rect 380 1883 531 1901
rect 565 1883 697 1917
rect 380 1871 697 1883
rect 749 1871 765 1923
rect 817 1871 833 1923
rect 885 1871 901 1923
rect 953 1871 969 1923
rect 1021 1917 1037 1923
rect 1021 1871 1037 1883
rect 1089 1871 1105 1923
rect 1157 1871 1173 1923
rect 1225 1917 1241 1923
rect 1293 1917 2097 1923
rect 1225 1883 1239 1917
rect 1293 1883 1475 1917
rect 1509 1883 1711 1917
rect 1745 1883 1947 1917
rect 1981 1883 2097 1917
rect 1225 1871 1241 1883
rect 1293 1871 2097 1883
rect 2149 1871 2165 1923
rect 2217 1871 2233 1923
rect 2285 1871 2301 1923
rect 2353 1871 2369 1923
rect 2421 1917 2437 1923
rect 2421 1871 2437 1883
rect 2489 1871 2505 1923
rect 2557 1871 2573 1923
rect 2625 1871 2641 1923
rect 2693 1919 3036 1923
rect 3070 1919 3076 1953
rect 2693 1909 3076 1919
rect 2693 1875 2891 1909
rect 2925 1880 3076 1909
rect 2925 1875 3036 1880
rect 2693 1871 3036 1875
rect 380 1863 3036 1871
rect 380 1829 386 1863
rect 420 1859 3036 1863
rect 420 1844 697 1859
rect 420 1829 531 1844
rect 380 1810 531 1829
rect 565 1810 697 1844
rect 380 1807 697 1810
rect 749 1807 765 1859
rect 817 1807 833 1859
rect 885 1807 901 1859
rect 953 1807 969 1859
rect 1021 1844 1037 1859
rect 1021 1807 1037 1810
rect 1089 1807 1105 1859
rect 1157 1807 1173 1859
rect 1225 1844 1241 1859
rect 1293 1844 2097 1859
rect 1225 1810 1239 1844
rect 1293 1810 1475 1844
rect 1509 1810 1711 1844
rect 1745 1810 1947 1844
rect 1981 1810 2097 1844
rect 1225 1807 1241 1810
rect 1293 1807 2097 1810
rect 2149 1807 2165 1859
rect 2217 1807 2233 1859
rect 2285 1807 2301 1859
rect 2353 1807 2369 1859
rect 2421 1844 2437 1859
rect 2421 1807 2437 1810
rect 2489 1807 2505 1859
rect 2557 1807 2573 1859
rect 2625 1807 2641 1859
rect 2693 1846 3036 1859
rect 3070 1846 3076 1880
rect 2693 1836 3076 1846
rect 2693 1807 2891 1836
rect 380 1802 2891 1807
rect 2925 1807 3076 1836
rect 2925 1802 3036 1807
rect 380 1795 3036 1802
rect 380 1791 697 1795
rect 380 1757 386 1791
rect 420 1770 697 1791
rect 420 1757 531 1770
rect 380 1736 531 1757
rect 565 1743 697 1770
rect 749 1743 765 1795
rect 817 1743 833 1795
rect 885 1743 901 1795
rect 953 1743 969 1795
rect 1021 1770 1037 1795
rect 1089 1743 1105 1795
rect 1157 1743 1173 1795
rect 1225 1770 1241 1795
rect 1293 1770 2097 1795
rect 1225 1743 1239 1770
rect 1293 1743 1475 1770
rect 565 1736 767 1743
rect 801 1736 1003 1743
rect 1037 1736 1239 1743
rect 1273 1736 1475 1743
rect 1509 1736 1711 1770
rect 1745 1736 1947 1770
rect 1981 1743 2097 1770
rect 2149 1743 2165 1795
rect 2217 1743 2233 1795
rect 2285 1743 2301 1795
rect 2353 1743 2369 1795
rect 2421 1770 2437 1795
rect 2489 1743 2505 1795
rect 2557 1743 2573 1795
rect 2625 1743 2641 1795
rect 2693 1773 3036 1795
rect 3070 1773 3076 1807
rect 2693 1762 3076 1773
rect 2693 1743 2891 1762
rect 1981 1736 2183 1743
rect 2217 1736 2419 1743
rect 2453 1736 2655 1743
rect 2689 1736 2891 1743
rect 380 1731 2891 1736
rect 380 1719 697 1731
rect 380 1685 386 1719
rect 420 1696 697 1719
rect 420 1685 531 1696
rect 380 1662 531 1685
rect 565 1679 697 1696
rect 749 1679 765 1731
rect 817 1679 833 1731
rect 885 1679 901 1731
rect 953 1679 969 1731
rect 1021 1696 1037 1731
rect 1089 1679 1105 1731
rect 1157 1679 1173 1731
rect 1225 1696 1241 1731
rect 1293 1696 2097 1731
rect 1225 1679 1239 1696
rect 1293 1679 1475 1696
rect 565 1667 767 1679
rect 801 1667 1003 1679
rect 1037 1667 1239 1679
rect 1273 1667 1475 1679
rect 565 1662 697 1667
rect 380 1647 697 1662
rect 380 1613 386 1647
rect 420 1622 697 1647
rect 420 1613 531 1622
rect 380 1588 531 1613
rect 565 1615 697 1622
rect 749 1615 765 1667
rect 817 1615 833 1667
rect 885 1615 901 1667
rect 953 1615 969 1667
rect 1021 1622 1037 1662
rect 1089 1615 1105 1667
rect 1157 1615 1173 1667
rect 1225 1662 1239 1667
rect 1293 1662 1475 1667
rect 1509 1662 1711 1696
rect 1745 1662 1947 1696
rect 1981 1679 2097 1696
rect 2149 1679 2165 1731
rect 2217 1679 2233 1731
rect 2285 1679 2301 1731
rect 2353 1679 2369 1731
rect 2421 1696 2437 1731
rect 2489 1679 2505 1731
rect 2557 1679 2573 1731
rect 2625 1679 2641 1731
rect 2693 1728 2891 1731
rect 2925 1734 3076 1762
rect 2925 1728 3036 1734
rect 2693 1700 3036 1728
rect 3070 1700 3076 1734
rect 2693 1688 3076 1700
rect 2693 1679 2891 1688
rect 1981 1667 2183 1679
rect 2217 1667 2419 1679
rect 2453 1667 2655 1679
rect 2689 1667 2891 1679
rect 1981 1662 2097 1667
rect 1225 1622 1241 1662
rect 1293 1622 2097 1662
rect 1225 1615 1239 1622
rect 1293 1615 1475 1622
rect 565 1603 767 1615
rect 801 1603 1003 1615
rect 1037 1603 1239 1615
rect 1273 1603 1475 1615
rect 565 1588 697 1603
rect 380 1575 697 1588
rect 380 1541 386 1575
rect 420 1551 697 1575
rect 749 1551 765 1603
rect 817 1551 833 1603
rect 885 1551 901 1603
rect 953 1551 969 1603
rect 1021 1551 1037 1588
rect 1089 1551 1105 1603
rect 1157 1551 1173 1603
rect 1225 1588 1239 1603
rect 1293 1588 1475 1603
rect 1509 1588 1711 1622
rect 1745 1588 1947 1622
rect 1981 1615 2097 1622
rect 2149 1615 2165 1667
rect 2217 1615 2233 1667
rect 2285 1615 2301 1667
rect 2353 1615 2369 1667
rect 2421 1622 2437 1662
rect 2489 1615 2505 1667
rect 2557 1615 2573 1667
rect 2625 1615 2641 1667
rect 2693 1654 2891 1667
rect 2925 1661 3076 1688
rect 2925 1654 3036 1661
rect 2693 1627 3036 1654
rect 3070 1627 3076 1661
rect 2693 1615 3076 1627
rect 1981 1603 2183 1615
rect 2217 1603 2419 1615
rect 2453 1603 2655 1615
rect 2689 1614 3076 1615
rect 2689 1603 2891 1614
rect 1981 1588 2097 1603
rect 1225 1551 1241 1588
rect 1293 1551 2097 1588
rect 2149 1551 2165 1603
rect 2217 1551 2233 1603
rect 2285 1551 2301 1603
rect 2353 1551 2369 1603
rect 2421 1551 2437 1588
rect 2489 1551 2505 1603
rect 2557 1551 2573 1603
rect 2625 1551 2641 1603
rect 2693 1580 2891 1603
rect 2925 1588 3076 1614
rect 2925 1580 3036 1588
rect 2693 1554 3036 1580
rect 3070 1554 3076 1588
rect 2693 1551 3076 1554
rect 420 1548 3076 1551
rect 420 1541 531 1548
rect 380 1514 531 1541
rect 565 1539 767 1548
rect 801 1539 1003 1548
rect 1037 1539 1239 1548
rect 1273 1539 1475 1548
rect 565 1514 697 1539
rect 380 1503 697 1514
rect 380 1469 386 1503
rect 420 1487 697 1503
rect 749 1487 765 1539
rect 817 1487 833 1539
rect 885 1487 901 1539
rect 953 1487 969 1539
rect 1021 1487 1037 1514
rect 1089 1487 1105 1539
rect 1157 1487 1173 1539
rect 1225 1514 1239 1539
rect 1293 1514 1475 1539
rect 1509 1514 1711 1548
rect 1745 1514 1947 1548
rect 1981 1539 2183 1548
rect 2217 1539 2419 1548
rect 2453 1539 2655 1548
rect 2689 1540 3076 1548
rect 2689 1539 2891 1540
rect 1981 1514 2097 1539
rect 1225 1487 1241 1514
rect 1293 1487 2097 1514
rect 2149 1487 2165 1539
rect 2217 1487 2233 1539
rect 2285 1487 2301 1539
rect 2353 1487 2369 1539
rect 2421 1487 2437 1514
rect 2489 1487 2505 1539
rect 2557 1487 2573 1539
rect 2625 1487 2641 1539
rect 2693 1506 2891 1539
rect 2925 1515 3076 1540
rect 2925 1506 3036 1515
rect 2693 1487 3036 1506
rect 420 1481 3036 1487
rect 3070 1481 3076 1515
rect 420 1475 3076 1481
rect 420 1474 697 1475
rect 420 1469 531 1474
rect 380 1440 531 1469
rect 565 1440 697 1474
rect 380 1431 697 1440
rect 380 1397 386 1431
rect 420 1423 697 1431
rect 749 1423 765 1475
rect 817 1423 833 1475
rect 885 1423 901 1475
rect 953 1423 969 1475
rect 1021 1474 1037 1475
rect 1021 1423 1037 1440
rect 1089 1423 1105 1475
rect 1157 1423 1173 1475
rect 1225 1474 1241 1475
rect 1293 1474 2097 1475
rect 1225 1440 1239 1474
rect 1293 1440 1475 1474
rect 1509 1440 1711 1474
rect 1745 1440 1947 1474
rect 1981 1440 2097 1474
rect 1225 1423 1241 1440
rect 1293 1423 2097 1440
rect 2149 1423 2165 1475
rect 2217 1423 2233 1475
rect 2285 1423 2301 1475
rect 2353 1423 2369 1475
rect 2421 1474 2437 1475
rect 2421 1423 2437 1440
rect 2489 1423 2505 1475
rect 2557 1423 2573 1475
rect 2625 1423 2641 1475
rect 2693 1466 3076 1475
rect 2693 1432 2891 1466
rect 2925 1442 3076 1466
rect 2925 1432 3036 1442
rect 2693 1423 3036 1432
rect 420 1411 3036 1423
rect 420 1400 697 1411
rect 420 1397 531 1400
rect 380 1366 531 1397
rect 565 1366 697 1400
rect 380 1359 697 1366
rect 749 1359 765 1411
rect 817 1359 833 1411
rect 885 1359 901 1411
rect 953 1359 969 1411
rect 1021 1400 1037 1411
rect 1021 1359 1037 1366
rect 1089 1359 1105 1411
rect 1157 1359 1173 1411
rect 1225 1400 1241 1411
rect 1293 1400 2097 1411
rect 1225 1366 1239 1400
rect 1293 1366 1475 1400
rect 1509 1366 1711 1400
rect 1745 1366 1947 1400
rect 1981 1366 2097 1400
rect 1225 1359 1241 1366
rect 1293 1359 2097 1366
rect 2149 1359 2165 1411
rect 2217 1359 2233 1411
rect 2285 1359 2301 1411
rect 2353 1359 2369 1411
rect 2421 1400 2437 1411
rect 2421 1359 2437 1366
rect 2489 1359 2505 1411
rect 2557 1359 2573 1411
rect 2625 1359 2641 1411
rect 2693 1408 3036 1411
rect 3070 1408 3076 1442
rect 2693 1392 3076 1408
rect 2693 1359 2891 1392
rect 380 1325 386 1359
rect 420 1358 2891 1359
rect 2925 1369 3076 1392
rect 2925 1358 3036 1369
rect 420 1347 3036 1358
rect 420 1326 697 1347
rect 420 1325 531 1326
rect 380 1292 531 1325
rect 565 1295 697 1326
rect 749 1295 765 1347
rect 817 1295 833 1347
rect 885 1295 901 1347
rect 953 1295 969 1347
rect 1021 1326 1037 1347
rect 1089 1295 1105 1347
rect 1157 1295 1173 1347
rect 1225 1326 1241 1347
rect 1293 1326 2097 1347
rect 1225 1295 1239 1326
rect 1293 1295 1475 1326
rect 565 1292 767 1295
rect 801 1292 1003 1295
rect 1037 1292 1239 1295
rect 1273 1292 1475 1295
rect 1509 1292 1711 1326
rect 1745 1292 1947 1326
rect 1981 1295 2097 1326
rect 2149 1295 2165 1347
rect 2217 1295 2233 1347
rect 2285 1295 2301 1347
rect 2353 1295 2369 1347
rect 2421 1326 2437 1347
rect 2489 1295 2505 1347
rect 2557 1295 2573 1347
rect 2625 1295 2641 1347
rect 2693 1335 3036 1347
rect 3070 1335 3076 1369
rect 2693 1318 3076 1335
rect 2693 1295 2891 1318
rect 1981 1292 2183 1295
rect 2217 1292 2419 1295
rect 2453 1292 2655 1295
rect 2689 1292 2891 1295
rect 380 1287 2891 1292
rect 380 1253 386 1287
rect 420 1284 2891 1287
rect 2925 1296 3076 1318
rect 2925 1284 3036 1296
rect 420 1267 3036 1284
rect 420 1262 600 1267
tri 600 1262 605 1267 nw
tri 727 1262 732 1267 ne
rect 732 1262 836 1267
tri 836 1262 841 1267 nw
tri 963 1262 968 1267 ne
rect 968 1262 1072 1267
tri 1072 1262 1077 1267 nw
tri 1199 1262 1204 1267 ne
rect 1204 1262 1308 1267
tri 1308 1262 1313 1267 nw
tri 1435 1262 1440 1267 ne
rect 1440 1262 1544 1267
tri 1544 1262 1549 1267 nw
tri 1671 1262 1676 1267 ne
rect 1676 1262 1780 1267
tri 1780 1262 1785 1267 nw
tri 1907 1262 1912 1267 ne
rect 1912 1262 2016 1267
tri 2016 1262 2021 1267 nw
tri 2143 1262 2148 1267 ne
rect 2148 1262 2252 1267
tri 2252 1262 2257 1267 nw
tri 2379 1262 2384 1267 ne
rect 2384 1262 2488 1267
tri 2488 1262 2493 1267 nw
tri 2615 1262 2620 1267 ne
rect 2620 1262 2724 1267
tri 2724 1262 2729 1267 nw
tri 2851 1262 2856 1267 ne
rect 2856 1262 3036 1267
rect 3070 1262 3076 1296
rect 420 1254 592 1262
tri 592 1254 600 1262 nw
tri 732 1254 740 1262 ne
rect 740 1254 828 1262
tri 828 1254 836 1262 nw
tri 968 1254 976 1262 ne
rect 976 1254 1064 1262
tri 1064 1254 1072 1262 nw
tri 1204 1254 1212 1262 ne
rect 1212 1254 1300 1262
tri 1300 1254 1308 1262 nw
tri 1440 1254 1448 1262 ne
rect 1448 1254 1536 1262
tri 1536 1254 1544 1262 nw
tri 1676 1254 1684 1262 ne
rect 1684 1254 1772 1262
tri 1772 1254 1780 1262 nw
tri 1912 1254 1920 1262 ne
rect 1920 1254 2008 1262
tri 2008 1254 2016 1262 nw
tri 2148 1254 2156 1262 ne
rect 2156 1254 2244 1262
tri 2244 1254 2252 1262 nw
tri 2384 1254 2392 1262 ne
rect 2392 1254 2480 1262
tri 2480 1254 2488 1262 nw
tri 2620 1254 2628 1262 ne
rect 2628 1254 2716 1262
tri 2716 1254 2724 1262 nw
tri 2856 1254 2864 1262 ne
rect 2864 1254 3076 1262
rect 420 1253 590 1254
rect 380 1252 590 1253
tri 590 1252 592 1254 nw
tri 740 1252 742 1254 ne
rect 742 1252 826 1254
tri 826 1252 828 1254 nw
tri 976 1252 978 1254 ne
rect 978 1252 1062 1254
tri 1062 1252 1064 1254 nw
tri 1212 1252 1214 1254 ne
rect 1214 1252 1298 1254
tri 1298 1252 1300 1254 nw
tri 1448 1252 1450 1254 ne
rect 1450 1252 1534 1254
tri 1534 1252 1536 1254 nw
tri 1684 1252 1686 1254 ne
rect 1686 1252 1770 1254
tri 1770 1252 1772 1254 nw
tri 1920 1252 1922 1254 ne
rect 1922 1252 2006 1254
tri 2006 1252 2008 1254 nw
tri 2156 1252 2158 1254 ne
rect 2158 1252 2242 1254
tri 2242 1252 2244 1254 nw
tri 2392 1252 2394 1254 ne
rect 2394 1252 2478 1254
tri 2478 1252 2480 1254 nw
tri 2628 1252 2630 1254 ne
rect 2630 1252 2706 1254
rect 380 1218 531 1252
rect 565 1218 571 1252
tri 571 1233 590 1252 nw
tri 742 1233 761 1252 ne
rect 380 1215 571 1218
rect 380 1181 386 1215
rect 420 1181 571 1215
rect 380 1178 571 1181
rect 380 1144 531 1178
rect 565 1144 571 1178
rect 380 1143 571 1144
rect 380 1109 386 1143
rect 420 1109 571 1143
rect 380 1104 571 1109
rect 380 1071 531 1104
rect 380 1037 386 1071
rect 420 1070 531 1071
rect 565 1070 571 1104
rect 420 1037 571 1070
rect 380 1030 571 1037
rect 380 999 531 1030
rect 380 965 386 999
rect 420 996 531 999
rect 565 996 571 1030
rect 420 965 571 996
rect 380 956 571 965
rect 380 927 531 956
rect 380 893 386 927
rect 420 922 531 927
rect 565 922 571 956
rect 420 893 571 922
rect 380 882 571 893
rect 380 855 531 882
rect 380 821 386 855
rect 420 848 531 855
rect 565 848 571 882
rect 420 821 571 848
rect 380 808 571 821
rect 380 783 531 808
rect 380 749 386 783
rect 420 774 531 783
rect 565 774 571 808
rect 420 749 571 774
rect 761 1218 767 1252
rect 801 1218 807 1252
tri 807 1233 826 1252 nw
tri 978 1233 997 1252 ne
rect 761 1178 807 1218
rect 761 1144 767 1178
rect 801 1144 807 1178
rect 761 1104 807 1144
rect 761 1070 767 1104
rect 801 1070 807 1104
rect 761 1030 807 1070
rect 761 996 767 1030
rect 801 996 807 1030
rect 761 956 807 996
rect 761 922 767 956
rect 801 922 807 956
rect 761 882 807 922
rect 761 848 767 882
rect 801 848 807 882
rect 761 808 807 848
rect 761 774 767 808
rect 801 774 807 808
rect 761 762 807 774
rect 997 1218 1003 1252
rect 1037 1218 1043 1252
tri 1043 1233 1062 1252 nw
tri 1214 1233 1233 1252 ne
rect 997 1178 1043 1218
rect 997 1144 1003 1178
rect 1037 1144 1043 1178
rect 997 1104 1043 1144
rect 997 1070 1003 1104
rect 1037 1070 1043 1104
rect 997 1030 1043 1070
rect 997 996 1003 1030
rect 1037 996 1043 1030
rect 997 956 1043 996
rect 997 922 1003 956
rect 1037 922 1043 956
rect 997 882 1043 922
rect 997 848 1003 882
rect 1037 848 1043 882
rect 997 808 1043 848
rect 997 774 1003 808
rect 1037 774 1043 808
rect 997 762 1043 774
rect 1233 1218 1239 1252
rect 1273 1218 1279 1252
tri 1279 1233 1298 1252 nw
tri 1450 1233 1469 1252 ne
rect 1233 1178 1279 1218
rect 1233 1144 1239 1178
rect 1273 1144 1279 1178
rect 1233 1104 1279 1144
rect 1233 1070 1239 1104
rect 1273 1070 1279 1104
rect 1233 1030 1279 1070
rect 1233 996 1239 1030
rect 1273 996 1279 1030
rect 1233 956 1279 996
rect 1233 922 1239 956
rect 1273 922 1279 956
rect 1233 882 1279 922
rect 1233 848 1239 882
rect 1273 848 1279 882
rect 1233 808 1279 848
rect 1233 774 1239 808
rect 1273 774 1279 808
rect 1233 762 1279 774
rect 1469 1218 1475 1252
rect 1509 1218 1515 1252
tri 1515 1233 1534 1252 nw
tri 1686 1233 1705 1252 ne
rect 1469 1178 1515 1218
rect 1469 1144 1475 1178
rect 1509 1144 1515 1178
rect 1469 1104 1515 1144
rect 1469 1070 1475 1104
rect 1509 1070 1515 1104
rect 1469 1030 1515 1070
rect 1469 996 1475 1030
rect 1509 996 1515 1030
rect 1469 956 1515 996
rect 1469 922 1475 956
rect 1509 922 1515 956
rect 1469 882 1515 922
rect 1469 848 1475 882
rect 1509 848 1515 882
rect 1469 808 1515 848
rect 1469 774 1475 808
rect 1509 774 1515 808
rect 1469 762 1515 774
rect 1705 1218 1711 1252
rect 1745 1218 1751 1252
tri 1751 1233 1770 1252 nw
tri 1922 1233 1941 1252 ne
rect 1705 1178 1751 1218
rect 1705 1144 1711 1178
rect 1745 1144 1751 1178
rect 1705 1104 1751 1144
rect 1705 1070 1711 1104
rect 1745 1070 1751 1104
rect 1705 1030 1751 1070
rect 1705 996 1711 1030
rect 1745 996 1751 1030
rect 1705 956 1751 996
rect 1705 922 1711 956
rect 1745 922 1751 956
rect 1705 882 1751 922
rect 1705 848 1711 882
rect 1745 848 1751 882
rect 1705 808 1751 848
rect 1705 774 1711 808
rect 1745 774 1751 808
rect 1705 762 1751 774
rect 1941 1218 1947 1252
rect 1981 1218 1987 1252
tri 1987 1233 2006 1252 nw
tri 2158 1233 2177 1252 ne
rect 1941 1178 1987 1218
rect 1941 1144 1947 1178
rect 1981 1144 1987 1178
rect 1941 1104 1987 1144
rect 1941 1070 1947 1104
rect 1981 1070 1987 1104
rect 1941 1030 1987 1070
rect 1941 996 1947 1030
rect 1981 996 1987 1030
rect 1941 956 1987 996
rect 1941 922 1947 956
rect 1981 922 1987 956
rect 1941 882 1987 922
rect 1941 848 1947 882
rect 1981 848 1987 882
rect 1941 808 1987 848
rect 1941 774 1947 808
rect 1981 774 1987 808
rect 1941 762 1987 774
rect 2177 1218 2183 1252
rect 2217 1218 2223 1252
tri 2223 1233 2242 1252 nw
tri 2394 1233 2413 1252 ne
rect 2177 1178 2223 1218
rect 2177 1144 2183 1178
rect 2217 1144 2223 1178
rect 2177 1104 2223 1144
rect 2177 1070 2183 1104
rect 2217 1070 2223 1104
rect 2177 1030 2223 1070
rect 2177 996 2183 1030
rect 2217 996 2223 1030
rect 2177 956 2223 996
rect 2177 922 2183 956
rect 2217 922 2223 956
rect 2177 882 2223 922
rect 2177 848 2183 882
rect 2217 848 2223 882
rect 2177 808 2223 848
rect 2177 774 2183 808
rect 2217 774 2223 808
rect 2177 762 2223 774
rect 2413 1218 2419 1252
rect 2453 1218 2459 1252
tri 2459 1233 2478 1252 nw
tri 2630 1233 2649 1252 ne
rect 2413 1178 2459 1218
rect 2413 1144 2419 1178
rect 2453 1144 2459 1178
rect 2413 1104 2459 1144
rect 2413 1070 2419 1104
rect 2453 1070 2459 1104
rect 2413 1030 2459 1070
rect 2413 996 2419 1030
rect 2453 996 2459 1030
rect 2413 956 2459 996
rect 2413 922 2419 956
rect 2453 922 2459 956
rect 2413 882 2459 922
rect 2413 848 2419 882
rect 2453 848 2459 882
rect 2413 808 2459 848
rect 2413 774 2419 808
rect 2453 774 2459 808
rect 2413 762 2459 774
rect 2649 1218 2655 1252
rect 2689 1244 2706 1252
tri 2706 1244 2716 1254 nw
tri 2864 1244 2874 1254 ne
rect 2874 1244 3076 1254
rect 2689 1218 2695 1244
tri 2695 1233 2706 1244 nw
tri 2874 1233 2885 1244 ne
rect 2649 1178 2695 1218
rect 2649 1144 2655 1178
rect 2689 1144 2695 1178
rect 2649 1104 2695 1144
rect 2649 1070 2655 1104
rect 2689 1070 2695 1104
rect 2649 1030 2695 1070
rect 2649 996 2655 1030
rect 2689 996 2695 1030
rect 2649 956 2695 996
rect 2649 922 2655 956
rect 2689 922 2695 956
rect 2649 882 2695 922
rect 2649 848 2655 882
rect 2689 848 2695 882
rect 2649 808 2695 848
rect 2649 774 2655 808
rect 2689 774 2695 808
rect 2649 762 2695 774
rect 2885 1210 2891 1244
rect 2925 1223 3076 1244
rect 2925 1210 3036 1223
rect 2885 1189 3036 1210
rect 3070 1189 3076 1223
rect 2885 1170 3076 1189
rect 2885 1136 2891 1170
rect 2925 1150 3076 1170
rect 2925 1136 3036 1150
rect 2885 1116 3036 1136
rect 3070 1116 3076 1150
rect 2885 1096 3076 1116
rect 2885 1062 2891 1096
rect 2925 1077 3076 1096
rect 2925 1062 3036 1077
rect 2885 1043 3036 1062
rect 3070 1043 3076 1077
rect 2885 1022 3076 1043
rect 2885 988 2891 1022
rect 2925 1004 3076 1022
rect 2925 988 3036 1004
rect 2885 970 3036 988
rect 3070 970 3076 1004
rect 2885 948 3076 970
rect 2885 914 2891 948
rect 2925 931 3076 948
rect 2925 914 3036 931
rect 2885 897 3036 914
rect 3070 897 3076 931
rect 2885 874 3076 897
rect 2885 840 2891 874
rect 2925 858 3076 874
rect 2925 840 3036 858
rect 2885 824 3036 840
rect 3070 824 3076 858
rect 2885 800 3076 824
rect 2885 766 2891 800
rect 2925 785 3076 800
rect 2925 766 3036 785
rect 380 711 571 749
rect 2885 751 3036 766
rect 3070 751 3076 785
rect 380 677 386 711
rect 420 677 571 711
rect 380 639 571 677
rect 613 714 1501 723
rect 1553 714 1569 723
rect 1621 714 1636 723
rect 1688 714 1703 723
rect 1755 714 1770 723
rect 1822 714 1837 723
rect 1889 714 2830 723
rect 613 680 625 714
rect 659 680 700 714
rect 734 680 775 714
rect 809 680 850 714
rect 884 680 925 714
rect 959 680 1000 714
rect 1034 680 1075 714
rect 1109 680 1150 714
rect 1184 680 1225 714
rect 1259 680 1300 714
rect 1334 680 1375 714
rect 1409 680 1450 714
rect 1484 680 1501 714
rect 1559 680 1569 714
rect 1634 680 1636 714
rect 1889 680 1896 714
rect 1930 680 1970 714
rect 2004 680 2044 714
rect 2078 680 2118 714
rect 2152 680 2192 714
rect 2226 680 2266 714
rect 2300 680 2340 714
rect 2374 680 2414 714
rect 2448 680 2488 714
rect 2522 680 2562 714
rect 2596 680 2636 714
rect 2670 680 2710 714
rect 2744 680 2784 714
rect 2818 680 2830 714
rect 613 671 1501 680
rect 1553 671 1569 680
rect 1621 671 1636 680
rect 1688 671 1703 680
rect 1755 671 1770 680
rect 1822 671 1837 680
rect 1889 671 2830 680
rect 2885 712 3076 751
rect 2885 678 3036 712
rect 3070 678 3076 712
rect 380 605 386 639
rect 420 605 571 639
rect 2885 639 3076 678
tri 571 605 573 607 sw
tri 2883 605 2885 607 se
rect 2885 605 3036 639
rect 3070 605 3076 639
rect 380 597 573 605
tri 573 597 581 605 sw
tri 2875 597 2883 605 se
rect 2883 597 3076 605
rect 380 573 581 597
tri 581 573 605 597 sw
tri 2851 573 2875 597 se
rect 2875 573 3076 597
rect 380 567 3076 573
rect 380 533 458 567
rect 492 533 532 567
rect 566 533 606 567
rect 640 533 680 567
rect 714 533 754 567
rect 788 533 828 567
rect 862 533 902 567
rect 936 533 976 567
rect 1010 533 1050 567
rect 1084 533 1124 567
rect 1158 533 1198 567
rect 1232 533 1272 567
rect 1306 533 1346 567
rect 1380 533 1420 567
rect 1454 533 1494 567
rect 1528 533 1568 567
rect 1602 533 1642 567
rect 1676 533 1716 567
rect 1750 533 1790 567
rect 1824 533 1864 567
rect 1898 533 1938 567
rect 1972 533 2012 567
rect 2046 533 2086 567
rect 2120 533 2160 567
rect 2194 533 2233 567
rect 2267 533 2306 567
rect 2340 533 2379 567
rect 2413 533 2452 567
rect 2486 533 2525 567
rect 2559 533 2598 567
rect 2632 533 2671 567
rect 2705 533 2744 567
rect 2778 533 2817 567
rect 2851 533 2890 567
rect 2924 533 2963 567
rect 2997 533 3076 567
rect 380 527 3076 533
rect 3287 39154 3339 39192
rect 3287 39120 3296 39154
rect 3330 39120 3339 39154
rect 3287 39082 3339 39120
rect 3287 39048 3296 39082
rect 3330 39048 3339 39082
rect 3287 39010 3339 39048
rect 3287 38976 3296 39010
rect 3330 38976 3339 39010
rect 3287 38938 3339 38976
rect 3287 38904 3296 38938
rect 3330 38904 3339 38938
rect 3287 38866 3339 38904
rect 3287 38832 3296 38866
rect 3330 38832 3339 38866
rect 3287 38794 3339 38832
rect 3287 38760 3296 38794
rect 3330 38760 3339 38794
rect 3287 38722 3339 38760
rect 3287 38688 3296 38722
rect 3330 38688 3339 38722
rect 3287 38650 3339 38688
rect 3287 38616 3296 38650
rect 3330 38616 3339 38650
rect 3287 38578 3339 38616
rect 3287 38544 3296 38578
rect 3330 38544 3339 38578
rect 3287 38506 3339 38544
rect 3287 38472 3296 38506
rect 3330 38472 3339 38506
rect 3287 38434 3339 38472
rect 3287 38400 3296 38434
rect 3330 38400 3339 38434
rect 3287 38362 3339 38400
rect 3287 38328 3296 38362
rect 3330 38328 3339 38362
rect 3287 38290 3339 38328
rect 3287 38256 3296 38290
rect 3330 38256 3339 38290
rect 3287 38218 3339 38256
rect 3287 38184 3296 38218
rect 3330 38184 3339 38218
rect 3287 38146 3339 38184
rect 3287 38112 3296 38146
rect 3330 38112 3339 38146
rect 3287 38074 3339 38112
rect 3287 38040 3296 38074
rect 3330 38040 3339 38074
rect 3287 38002 3339 38040
rect 3287 37968 3296 38002
rect 3330 37968 3339 38002
rect 3287 37930 3339 37968
rect 3287 37896 3296 37930
rect 3330 37896 3339 37930
rect 3287 37858 3339 37896
rect 3287 37824 3296 37858
rect 3330 37824 3339 37858
rect 3287 37786 3339 37824
rect 3287 37752 3296 37786
rect 3330 37752 3339 37786
rect 3287 37714 3339 37752
rect 3287 37680 3296 37714
rect 3330 37680 3339 37714
rect 3287 37642 3339 37680
rect 3287 37608 3296 37642
rect 3330 37608 3339 37642
rect 3287 37570 3339 37608
rect 3287 37536 3296 37570
rect 3330 37536 3339 37570
rect 3287 37498 3339 37536
rect 3287 37464 3296 37498
rect 3330 37464 3339 37498
rect 3287 37426 3339 37464
rect 3287 37392 3296 37426
rect 3330 37392 3339 37426
rect 3287 37354 3339 37392
rect 3287 37320 3296 37354
rect 3330 37320 3339 37354
rect 3287 37282 3339 37320
rect 3287 37248 3296 37282
rect 3330 37248 3339 37282
rect 3287 37210 3339 37248
rect 3287 37176 3296 37210
rect 3330 37176 3339 37210
rect 3287 37138 3339 37176
rect 3287 37104 3296 37138
rect 3330 37104 3339 37138
rect 3287 37066 3339 37104
rect 3287 37032 3296 37066
rect 3330 37032 3339 37066
rect 3287 36994 3339 37032
rect 3287 36960 3296 36994
rect 3330 36960 3339 36994
rect 3287 36922 3339 36960
rect 3287 36888 3296 36922
rect 3330 36888 3339 36922
rect 3287 36850 3339 36888
rect 3287 36816 3296 36850
rect 3330 36816 3339 36850
rect 3287 36778 3339 36816
rect 3287 36744 3296 36778
rect 3330 36744 3339 36778
rect 3287 36706 3339 36744
rect 3287 36672 3296 36706
rect 3330 36672 3339 36706
rect 3287 36634 3339 36672
rect 3287 36600 3296 36634
rect 3330 36600 3339 36634
rect 3287 36562 3339 36600
rect 3287 36528 3296 36562
rect 3330 36528 3339 36562
rect 3287 36490 3339 36528
rect 3287 36456 3296 36490
rect 3330 36456 3339 36490
rect 3287 36418 3339 36456
rect 3287 36384 3296 36418
rect 3330 36384 3339 36418
rect 3287 36346 3339 36384
rect 3287 36312 3296 36346
rect 3330 36312 3339 36346
rect 3287 36274 3339 36312
rect 3287 36240 3296 36274
rect 3330 36240 3339 36274
rect 3287 36202 3339 36240
rect 3287 36168 3296 36202
rect 3330 36168 3339 36202
rect 3287 36130 3339 36168
rect 3287 36096 3296 36130
rect 3330 36096 3339 36130
rect 3287 36058 3339 36096
rect 3287 36024 3296 36058
rect 3330 36024 3339 36058
rect 3287 35986 3339 36024
rect 3287 35952 3296 35986
rect 3330 35952 3339 35986
rect 3287 35914 3339 35952
rect 3287 35880 3296 35914
rect 3330 35880 3339 35914
rect 3287 35842 3339 35880
rect 3287 35808 3296 35842
rect 3330 35808 3339 35842
rect 3287 35770 3339 35808
rect 3287 35736 3296 35770
rect 3330 35736 3339 35770
rect 3287 35698 3339 35736
rect 3287 35664 3296 35698
rect 3330 35664 3339 35698
rect 3287 35626 3339 35664
rect 3287 35592 3296 35626
rect 3330 35592 3339 35626
rect 3287 35554 3339 35592
rect 3287 35520 3296 35554
rect 3330 35520 3339 35554
rect 3287 35482 3339 35520
rect 3287 35448 3296 35482
rect 3330 35448 3339 35482
rect 3287 35410 3339 35448
rect 3287 35376 3296 35410
rect 3330 35376 3339 35410
rect 3287 35338 3339 35376
rect 3287 35304 3296 35338
rect 3330 35304 3339 35338
rect 3287 35266 3339 35304
rect 3287 35232 3296 35266
rect 3330 35232 3339 35266
rect 3287 35194 3339 35232
rect 3287 35160 3296 35194
rect 3330 35160 3339 35194
rect 3287 35122 3339 35160
rect 3287 35088 3296 35122
rect 3330 35088 3339 35122
rect 3287 35050 3339 35088
rect 3287 35016 3296 35050
rect 3330 35016 3339 35050
rect 3287 34978 3339 35016
rect 3287 34944 3296 34978
rect 3330 34944 3339 34978
rect 3287 34906 3339 34944
rect 3287 34872 3296 34906
rect 3330 34872 3339 34906
rect 3287 34834 3339 34872
rect 3287 34800 3296 34834
rect 3330 34800 3339 34834
rect 3287 34762 3339 34800
rect 3287 34728 3296 34762
rect 3330 34728 3339 34762
rect 3287 34690 3339 34728
rect 3287 34656 3296 34690
rect 3330 34656 3339 34690
rect 3287 34618 3339 34656
rect 3287 34584 3296 34618
rect 3330 34584 3339 34618
rect 3287 34546 3339 34584
rect 3287 34512 3296 34546
rect 3330 34512 3339 34546
rect 3287 34474 3339 34512
rect 3287 34440 3296 34474
rect 3330 34440 3339 34474
rect 3287 34402 3339 34440
rect 3287 34368 3296 34402
rect 3330 34368 3339 34402
rect 3287 34330 3339 34368
rect 3287 34296 3296 34330
rect 3330 34296 3339 34330
rect 3287 34258 3339 34296
rect 3287 34224 3296 34258
rect 3330 34224 3339 34258
rect 3287 34186 3339 34224
rect 3287 34152 3296 34186
rect 3330 34152 3339 34186
rect 3287 34114 3339 34152
rect 3287 34080 3296 34114
rect 3330 34080 3339 34114
rect 3287 34042 3339 34080
rect 3287 34008 3296 34042
rect 3330 34008 3339 34042
rect 3287 33970 3339 34008
rect 3287 33936 3296 33970
rect 3330 33936 3339 33970
rect 3287 33898 3339 33936
rect 3287 33864 3296 33898
rect 3330 33864 3339 33898
rect 3287 33826 3339 33864
rect 3287 33792 3296 33826
rect 3330 33792 3339 33826
rect 3287 33754 3339 33792
rect 3287 33720 3296 33754
rect 3330 33720 3339 33754
rect 3287 33682 3339 33720
rect 3287 33648 3296 33682
rect 3330 33648 3339 33682
rect 3287 33610 3339 33648
rect 3287 33576 3296 33610
rect 3330 33576 3339 33610
rect 3287 33538 3339 33576
rect 3287 33504 3296 33538
rect 3330 33504 3339 33538
rect 3287 33466 3339 33504
rect 3287 33432 3296 33466
rect 3330 33432 3339 33466
rect 3287 33394 3339 33432
rect 3287 33360 3296 33394
rect 3330 33360 3339 33394
rect 3287 33322 3339 33360
rect 3287 33288 3296 33322
rect 3330 33288 3339 33322
rect 3287 33250 3339 33288
rect 3287 33216 3296 33250
rect 3330 33216 3339 33250
rect 3287 33178 3339 33216
rect 3287 33144 3296 33178
rect 3330 33144 3339 33178
rect 3287 33106 3339 33144
rect 3287 33072 3296 33106
rect 3330 33072 3339 33106
rect 3287 33034 3339 33072
rect 3287 33000 3296 33034
rect 3330 33000 3339 33034
rect 3287 32962 3339 33000
rect 3287 32928 3296 32962
rect 3330 32928 3339 32962
rect 3287 32890 3339 32928
rect 3287 32856 3296 32890
rect 3330 32856 3339 32890
rect 3287 32818 3339 32856
rect 3287 32784 3296 32818
rect 3330 32784 3339 32818
rect 3287 32746 3339 32784
rect 3287 32712 3296 32746
rect 3330 32712 3339 32746
rect 3287 32674 3339 32712
rect 3287 32640 3296 32674
rect 3330 32640 3339 32674
rect 3287 32602 3339 32640
rect 3287 32568 3296 32602
rect 3330 32568 3339 32602
rect 3287 32530 3339 32568
rect 3287 32496 3296 32530
rect 3330 32496 3339 32530
rect 3287 32458 3339 32496
rect 3287 32424 3296 32458
rect 3330 32424 3339 32458
rect 3287 32386 3339 32424
rect 3287 32352 3296 32386
rect 3330 32352 3339 32386
rect 3287 32314 3339 32352
rect 3287 32280 3296 32314
rect 3330 32280 3339 32314
rect 3287 32242 3339 32280
rect 3287 32208 3296 32242
rect 3330 32208 3339 32242
rect 3287 32170 3339 32208
rect 3287 32136 3296 32170
rect 3330 32136 3339 32170
rect 3287 32098 3339 32136
rect 3287 32064 3296 32098
rect 3330 32064 3339 32098
rect 3287 32026 3339 32064
rect 3287 31992 3296 32026
rect 3330 31992 3339 32026
rect 3287 31954 3339 31992
rect 3287 31920 3296 31954
rect 3330 31920 3339 31954
rect 3287 31882 3339 31920
rect 3287 31848 3296 31882
rect 3330 31848 3339 31882
rect 3287 31810 3339 31848
rect 3287 31776 3296 31810
rect 3330 31776 3339 31810
rect 3287 31738 3339 31776
rect 3287 31704 3296 31738
rect 3330 31704 3339 31738
rect 3287 31666 3339 31704
rect 3287 31632 3296 31666
rect 3330 31632 3339 31666
rect 3287 31594 3339 31632
rect 3287 31560 3296 31594
rect 3330 31560 3339 31594
rect 3287 31522 3339 31560
rect 3287 31488 3296 31522
rect 3330 31488 3339 31522
rect 3287 31450 3339 31488
rect 3287 31416 3296 31450
rect 3330 31416 3339 31450
rect 3287 31378 3339 31416
rect 3287 31344 3296 31378
rect 3330 31344 3339 31378
rect 3287 31306 3339 31344
rect 3287 31272 3296 31306
rect 3330 31272 3339 31306
rect 3287 31234 3339 31272
rect 3287 31200 3296 31234
rect 3330 31200 3339 31234
rect 3287 31162 3339 31200
rect 3287 31128 3296 31162
rect 3330 31128 3339 31162
rect 3287 31090 3339 31128
rect 3287 31056 3296 31090
rect 3330 31056 3339 31090
rect 3287 31018 3339 31056
rect 3287 30984 3296 31018
rect 3330 30984 3339 31018
rect 3287 30946 3339 30984
rect 3287 30912 3296 30946
rect 3330 30912 3339 30946
rect 3287 30874 3339 30912
rect 3287 30840 3296 30874
rect 3330 30840 3339 30874
rect 3287 30802 3339 30840
rect 3287 30768 3296 30802
rect 3330 30768 3339 30802
rect 3287 30730 3339 30768
rect 3287 30696 3296 30730
rect 3330 30696 3339 30730
rect 3287 30658 3339 30696
rect 3287 30624 3296 30658
rect 3330 30624 3339 30658
rect 3287 30586 3339 30624
rect 3287 30552 3296 30586
rect 3330 30552 3339 30586
rect 3287 30514 3339 30552
rect 3287 30480 3296 30514
rect 3330 30480 3339 30514
rect 3287 30442 3339 30480
rect 3287 30408 3296 30442
rect 3330 30408 3339 30442
rect 3287 30370 3339 30408
rect 3287 30336 3296 30370
rect 3330 30336 3339 30370
rect 3287 30298 3339 30336
rect 3287 30264 3296 30298
rect 3330 30264 3339 30298
rect 3287 30226 3339 30264
rect 3287 30192 3296 30226
rect 3330 30192 3339 30226
rect 3287 30154 3339 30192
rect 3287 30120 3296 30154
rect 3330 30120 3339 30154
rect 3287 30082 3339 30120
rect 3287 30048 3296 30082
rect 3330 30048 3339 30082
rect 3287 30010 3339 30048
rect 3287 29976 3296 30010
rect 3330 29976 3339 30010
rect 3287 29938 3339 29976
rect 3287 29904 3296 29938
rect 3330 29904 3339 29938
rect 3287 29866 3339 29904
rect 3287 29832 3296 29866
rect 3330 29832 3339 29866
rect 3287 29794 3339 29832
rect 3287 29760 3296 29794
rect 3330 29760 3339 29794
rect 3287 29722 3339 29760
rect 3287 29688 3296 29722
rect 3330 29688 3339 29722
rect 3287 29650 3339 29688
rect 3287 29616 3296 29650
rect 3330 29616 3339 29650
rect 3287 29578 3339 29616
rect 3287 29544 3296 29578
rect 3330 29544 3339 29578
rect 3287 29506 3339 29544
rect 3287 29472 3296 29506
rect 3330 29472 3339 29506
rect 3287 29434 3339 29472
rect 3287 29400 3296 29434
rect 3330 29400 3339 29434
rect 3287 29362 3339 29400
rect 3287 29328 3296 29362
rect 3330 29328 3339 29362
rect 3287 29290 3339 29328
rect 3287 29256 3296 29290
rect 3330 29256 3339 29290
rect 3287 29218 3339 29256
rect 3287 29184 3296 29218
rect 3330 29184 3339 29218
rect 3287 29146 3339 29184
rect 3287 29112 3296 29146
rect 3330 29112 3339 29146
rect 3287 29074 3339 29112
rect 3287 29040 3296 29074
rect 3330 29040 3339 29074
rect 3287 29002 3339 29040
rect 3287 28968 3296 29002
rect 3330 28968 3339 29002
rect 3287 28930 3339 28968
rect 3287 28896 3296 28930
rect 3330 28896 3339 28930
rect 3287 28858 3339 28896
rect 3287 28824 3296 28858
rect 3330 28824 3339 28858
rect 3287 28786 3339 28824
rect 3287 28752 3296 28786
rect 3330 28752 3339 28786
rect 3287 28714 3339 28752
rect 3287 28680 3296 28714
rect 3330 28680 3339 28714
rect 3287 28642 3339 28680
rect 3287 28608 3296 28642
rect 3330 28608 3339 28642
rect 3287 28570 3339 28608
rect 3287 28536 3296 28570
rect 3330 28536 3339 28570
rect 3287 28498 3339 28536
rect 3287 28464 3296 28498
rect 3330 28464 3339 28498
rect 3287 28426 3339 28464
rect 3287 28392 3296 28426
rect 3330 28392 3339 28426
rect 3287 28354 3339 28392
rect 3287 28320 3296 28354
rect 3330 28320 3339 28354
rect 3287 28282 3339 28320
rect 3287 28248 3296 28282
rect 3330 28248 3339 28282
rect 3287 28210 3339 28248
rect 3287 28176 3296 28210
rect 3330 28176 3339 28210
rect 3287 28138 3339 28176
rect 3287 28104 3296 28138
rect 3330 28104 3339 28138
rect 3287 28066 3339 28104
rect 3287 28032 3296 28066
rect 3330 28032 3339 28066
rect 3287 27994 3339 28032
rect 3287 27960 3296 27994
rect 3330 27960 3339 27994
rect 3287 27922 3339 27960
rect 3287 27888 3296 27922
rect 3330 27888 3339 27922
rect 3287 27850 3339 27888
rect 3287 27816 3296 27850
rect 3330 27816 3339 27850
rect 3287 27778 3339 27816
rect 3287 27744 3296 27778
rect 3330 27744 3339 27778
rect 3287 27706 3339 27744
rect 3287 27672 3296 27706
rect 3330 27672 3339 27706
rect 3287 27634 3339 27672
rect 3287 27600 3296 27634
rect 3330 27600 3339 27634
rect 3287 27562 3339 27600
rect 3287 27528 3296 27562
rect 3330 27528 3339 27562
rect 3287 27490 3339 27528
rect 3287 27456 3296 27490
rect 3330 27456 3339 27490
rect 3287 27418 3339 27456
rect 3287 27384 3296 27418
rect 3330 27384 3339 27418
rect 3287 27346 3339 27384
rect 3287 27312 3296 27346
rect 3330 27312 3339 27346
rect 3287 27274 3339 27312
rect 3287 27240 3296 27274
rect 3330 27240 3339 27274
rect 3287 27202 3339 27240
rect 3287 27168 3296 27202
rect 3330 27168 3339 27202
rect 3287 27130 3339 27168
rect 3287 27096 3296 27130
rect 3330 27096 3339 27130
rect 3287 27058 3339 27096
rect 3287 27024 3296 27058
rect 3330 27024 3339 27058
rect 3287 26986 3339 27024
rect 3287 26952 3296 26986
rect 3330 26952 3339 26986
rect 3287 26914 3339 26952
rect 3287 26880 3296 26914
rect 3330 26880 3339 26914
rect 3287 26842 3339 26880
rect 3287 26808 3296 26842
rect 3330 26808 3339 26842
rect 3287 26770 3339 26808
rect 3287 26736 3296 26770
rect 3330 26736 3339 26770
rect 3287 26698 3339 26736
rect 3287 26664 3296 26698
rect 3330 26664 3339 26698
rect 3287 26626 3339 26664
rect 3287 26592 3296 26626
rect 3330 26592 3339 26626
rect 3287 26554 3339 26592
rect 3287 26520 3296 26554
rect 3330 26520 3339 26554
rect 3287 26482 3339 26520
rect 3287 26448 3296 26482
rect 3330 26448 3339 26482
rect 3287 26410 3339 26448
rect 3287 26376 3296 26410
rect 3330 26376 3339 26410
rect 3287 26338 3339 26376
rect 3287 26304 3296 26338
rect 3330 26304 3339 26338
rect 3287 26266 3339 26304
rect 3287 26232 3296 26266
rect 3330 26232 3339 26266
rect 3287 26194 3339 26232
rect 3287 26160 3296 26194
rect 3330 26160 3339 26194
rect 3287 26122 3339 26160
rect 3287 26088 3296 26122
rect 3330 26088 3339 26122
rect 3287 26050 3339 26088
rect 3287 26016 3296 26050
rect 3330 26016 3339 26050
rect 3287 25978 3339 26016
rect 3287 25944 3296 25978
rect 3330 25944 3339 25978
rect 3287 25906 3339 25944
rect 3287 25872 3296 25906
rect 3330 25872 3339 25906
rect 3287 25834 3339 25872
rect 3287 25800 3296 25834
rect 3330 25800 3339 25834
rect 3287 25762 3339 25800
rect 3287 25728 3296 25762
rect 3330 25728 3339 25762
rect 3287 25690 3339 25728
rect 3287 25656 3296 25690
rect 3330 25656 3339 25690
rect 3287 25618 3339 25656
rect 3287 25584 3296 25618
rect 3330 25584 3339 25618
rect 3287 25546 3339 25584
rect 3287 25512 3296 25546
rect 3330 25512 3339 25546
rect 3287 25474 3339 25512
rect 3287 25440 3296 25474
rect 3330 25440 3339 25474
rect 3287 25402 3339 25440
rect 3287 25368 3296 25402
rect 3330 25368 3339 25402
rect 3287 25330 3339 25368
rect 3287 25296 3296 25330
rect 3330 25296 3339 25330
rect 3287 25258 3339 25296
rect 3287 25224 3296 25258
rect 3330 25224 3339 25258
rect 3287 25186 3339 25224
rect 3287 25152 3296 25186
rect 3330 25152 3339 25186
rect 3287 25114 3339 25152
rect 3287 25080 3296 25114
rect 3330 25080 3339 25114
rect 3287 25042 3339 25080
rect 3287 25008 3296 25042
rect 3330 25008 3339 25042
rect 3287 24970 3339 25008
rect 3287 24936 3296 24970
rect 3330 24936 3339 24970
rect 3287 24898 3339 24936
rect 3287 24864 3296 24898
rect 3330 24864 3339 24898
rect 3287 24826 3339 24864
rect 3287 24792 3296 24826
rect 3330 24792 3339 24826
rect 3287 24754 3339 24792
rect 3287 24720 3296 24754
rect 3330 24720 3339 24754
rect 3287 24682 3339 24720
rect 3287 24648 3296 24682
rect 3330 24648 3339 24682
rect 3287 24610 3339 24648
rect 3287 24576 3296 24610
rect 3330 24576 3339 24610
rect 3287 24538 3339 24576
rect 3287 24504 3296 24538
rect 3330 24504 3339 24538
rect 3287 24466 3339 24504
rect 3287 24432 3296 24466
rect 3330 24432 3339 24466
rect 3287 24394 3339 24432
rect 3287 24360 3296 24394
rect 3330 24360 3339 24394
rect 3287 24322 3339 24360
rect 3287 24288 3296 24322
rect 3330 24288 3339 24322
rect 3287 24250 3339 24288
rect 3287 24216 3296 24250
rect 3330 24216 3339 24250
rect 3287 24178 3339 24216
rect 3287 24144 3296 24178
rect 3330 24144 3339 24178
rect 3287 24106 3339 24144
rect 3287 24072 3296 24106
rect 3330 24072 3339 24106
rect 3287 24034 3339 24072
rect 3287 24000 3296 24034
rect 3330 24000 3339 24034
rect 3287 23962 3339 24000
rect 3287 23928 3296 23962
rect 3330 23928 3339 23962
rect 3287 23890 3339 23928
rect 3287 23856 3296 23890
rect 3330 23856 3339 23890
rect 3287 23818 3339 23856
rect 3287 23784 3296 23818
rect 3330 23784 3339 23818
rect 3287 23746 3339 23784
rect 3287 23712 3296 23746
rect 3330 23712 3339 23746
rect 3287 23674 3339 23712
rect 3287 23640 3296 23674
rect 3330 23640 3339 23674
rect 3287 23602 3339 23640
rect 3287 23568 3296 23602
rect 3330 23568 3339 23602
rect 3287 23530 3339 23568
rect 3287 23496 3296 23530
rect 3330 23496 3339 23530
rect 3287 23458 3339 23496
rect 3287 23424 3296 23458
rect 3330 23424 3339 23458
rect 3287 23386 3339 23424
rect 3287 23352 3296 23386
rect 3330 23352 3339 23386
rect 3287 23314 3339 23352
rect 3287 23280 3296 23314
rect 3330 23280 3339 23314
rect 3287 23242 3339 23280
rect 3287 23208 3296 23242
rect 3330 23208 3339 23242
rect 3287 23170 3339 23208
rect 3287 23136 3296 23170
rect 3330 23136 3339 23170
rect 3287 23098 3339 23136
rect 3287 23064 3296 23098
rect 3330 23064 3339 23098
rect 3287 23026 3339 23064
rect 3287 22992 3296 23026
rect 3330 22992 3339 23026
rect 3287 22954 3339 22992
rect 3287 22920 3296 22954
rect 3330 22920 3339 22954
rect 3287 22882 3339 22920
rect 3287 22848 3296 22882
rect 3330 22848 3339 22882
rect 3287 22810 3339 22848
rect 3287 22776 3296 22810
rect 3330 22776 3339 22810
rect 3287 22738 3339 22776
rect 3287 22704 3296 22738
rect 3330 22704 3339 22738
rect 3287 22666 3339 22704
rect 3287 22632 3296 22666
rect 3330 22632 3339 22666
rect 3287 22594 3339 22632
rect 3287 22560 3296 22594
rect 3330 22560 3339 22594
rect 3287 22522 3339 22560
rect 3287 22488 3296 22522
rect 3330 22488 3339 22522
rect 3287 22450 3339 22488
rect 3287 22416 3296 22450
rect 3330 22416 3339 22450
rect 3287 22378 3339 22416
rect 3287 22344 3296 22378
rect 3330 22344 3339 22378
rect 3287 22306 3339 22344
rect 3287 22272 3296 22306
rect 3330 22272 3339 22306
rect 3287 22234 3339 22272
rect 3287 22200 3296 22234
rect 3330 22200 3339 22234
rect 3287 22162 3339 22200
rect 3287 22128 3296 22162
rect 3330 22128 3339 22162
rect 3287 22090 3339 22128
rect 3287 22056 3296 22090
rect 3330 22056 3339 22090
rect 3287 22018 3339 22056
rect 3287 21984 3296 22018
rect 3330 21984 3339 22018
rect 3287 21946 3339 21984
rect 3287 21912 3296 21946
rect 3330 21912 3339 21946
rect 3287 21874 3339 21912
rect 3287 21840 3296 21874
rect 3330 21840 3339 21874
rect 3287 21802 3339 21840
rect 3287 21768 3296 21802
rect 3330 21768 3339 21802
rect 3287 21730 3339 21768
rect 3287 21696 3296 21730
rect 3330 21696 3339 21730
rect 3287 21658 3339 21696
rect 3287 21624 3296 21658
rect 3330 21624 3339 21658
rect 3287 21586 3339 21624
rect 3287 21552 3296 21586
rect 3330 21552 3339 21586
rect 3287 21514 3339 21552
rect 3287 21480 3296 21514
rect 3330 21480 3339 21514
rect 3287 21442 3339 21480
rect 3287 21408 3296 21442
rect 3330 21408 3339 21442
rect 3287 21370 3339 21408
rect 3287 21336 3296 21370
rect 3330 21336 3339 21370
rect 3287 21298 3339 21336
rect 3287 21264 3296 21298
rect 3330 21264 3339 21298
rect 3287 21226 3339 21264
rect 3287 21192 3296 21226
rect 3330 21192 3339 21226
rect 3287 21154 3339 21192
rect 3287 21120 3296 21154
rect 3330 21120 3339 21154
rect 3287 21082 3339 21120
rect 3287 21048 3296 21082
rect 3330 21048 3339 21082
rect 3287 21010 3339 21048
rect 3287 20976 3296 21010
rect 3330 20976 3339 21010
rect 3287 20938 3339 20976
rect 3287 20904 3296 20938
rect 3330 20904 3339 20938
rect 3287 20866 3339 20904
rect 3287 20832 3296 20866
rect 3330 20832 3339 20866
rect 3287 20794 3339 20832
rect 3287 20760 3296 20794
rect 3330 20760 3339 20794
rect 3287 20722 3339 20760
rect 3287 20688 3296 20722
rect 3330 20688 3339 20722
rect 3287 20650 3339 20688
rect 3287 20616 3296 20650
rect 3330 20616 3339 20650
rect 3287 20578 3339 20616
rect 3287 20544 3296 20578
rect 3330 20544 3339 20578
rect 3287 20506 3339 20544
rect 3287 20472 3296 20506
rect 3330 20472 3339 20506
rect 3287 20434 3339 20472
rect 3287 20400 3296 20434
rect 3330 20400 3339 20434
rect 3287 20362 3339 20400
rect 3287 20328 3296 20362
rect 3330 20328 3339 20362
rect 3287 20290 3339 20328
rect 3287 20256 3296 20290
rect 3330 20256 3339 20290
rect 3287 20218 3339 20256
rect 3287 20184 3296 20218
rect 3330 20184 3339 20218
rect 3287 20146 3339 20184
rect 3287 20112 3296 20146
rect 3330 20112 3339 20146
rect 3287 20074 3339 20112
rect 3287 20040 3296 20074
rect 3330 20040 3339 20074
rect 3287 20002 3339 20040
rect 3287 19968 3296 20002
rect 3330 19968 3339 20002
rect 3287 19930 3339 19968
rect 3287 19896 3296 19930
rect 3330 19896 3339 19930
rect 3287 19858 3339 19896
rect 3287 19824 3296 19858
rect 3330 19824 3339 19858
rect 3287 19786 3339 19824
rect 3287 19752 3296 19786
rect 3330 19752 3339 19786
rect 3287 19714 3339 19752
rect 3287 19680 3296 19714
rect 3330 19680 3339 19714
rect 3287 19642 3339 19680
rect 3287 19608 3296 19642
rect 3330 19608 3339 19642
rect 3287 19570 3339 19608
rect 3287 19536 3296 19570
rect 3330 19536 3339 19570
rect 3287 19498 3339 19536
rect 3287 19464 3296 19498
rect 3330 19464 3339 19498
rect 3287 19426 3339 19464
rect 3287 19392 3296 19426
rect 3330 19392 3339 19426
rect 3287 19354 3339 19392
rect 3287 19320 3296 19354
rect 3330 19320 3339 19354
rect 3287 19282 3339 19320
rect 3287 19248 3296 19282
rect 3330 19248 3339 19282
rect 3287 19210 3339 19248
rect 3287 19176 3296 19210
rect 3330 19176 3339 19210
rect 3287 19138 3339 19176
rect 3287 19104 3296 19138
rect 3330 19104 3339 19138
rect 3287 19066 3339 19104
rect 3287 19032 3296 19066
rect 3330 19032 3339 19066
rect 3287 18994 3339 19032
rect 3287 18960 3296 18994
rect 3330 18960 3339 18994
rect 3287 18922 3339 18960
rect 3287 18888 3296 18922
rect 3330 18888 3339 18922
rect 3287 18850 3339 18888
rect 3287 18816 3296 18850
rect 3330 18816 3339 18850
rect 3287 18778 3339 18816
rect 3287 18744 3296 18778
rect 3330 18744 3339 18778
rect 3287 18706 3339 18744
rect 3287 18672 3296 18706
rect 3330 18672 3339 18706
rect 3287 18634 3339 18672
rect 3287 18600 3296 18634
rect 3330 18600 3339 18634
rect 3287 18562 3339 18600
rect 3287 18528 3296 18562
rect 3330 18528 3339 18562
rect 3287 18490 3339 18528
rect 3287 18456 3296 18490
rect 3330 18456 3339 18490
rect 3287 18418 3339 18456
rect 3287 18384 3296 18418
rect 3330 18384 3339 18418
rect 3287 18346 3339 18384
rect 3287 18312 3296 18346
rect 3330 18312 3339 18346
rect 3287 18274 3339 18312
rect 3287 18240 3296 18274
rect 3330 18240 3339 18274
rect 3287 18202 3339 18240
rect 3287 18168 3296 18202
rect 3330 18168 3339 18202
rect 3287 18130 3339 18168
rect 3287 18096 3296 18130
rect 3330 18096 3339 18130
rect 3287 18058 3339 18096
rect 3287 18024 3296 18058
rect 3330 18024 3339 18058
rect 3287 17986 3339 18024
rect 3287 17952 3296 17986
rect 3330 17952 3339 17986
rect 3287 17914 3339 17952
rect 3287 17880 3296 17914
rect 3330 17880 3339 17914
rect 3287 17842 3339 17880
rect 3287 17808 3296 17842
rect 3330 17808 3339 17842
rect 3287 17770 3339 17808
rect 3287 17736 3296 17770
rect 3330 17736 3339 17770
rect 3287 17698 3339 17736
rect 3287 17664 3296 17698
rect 3330 17664 3339 17698
rect 3287 17626 3339 17664
rect 3287 17592 3296 17626
rect 3330 17592 3339 17626
rect 3287 17554 3339 17592
rect 3287 17520 3296 17554
rect 3330 17520 3339 17554
rect 3287 17482 3339 17520
rect 3287 17448 3296 17482
rect 3330 17448 3339 17482
rect 3287 17410 3339 17448
rect 3287 17376 3296 17410
rect 3330 17376 3339 17410
rect 3287 17338 3339 17376
rect 3287 17304 3296 17338
rect 3330 17304 3339 17338
rect 3287 17266 3339 17304
rect 3287 17232 3296 17266
rect 3330 17232 3339 17266
rect 3287 17194 3339 17232
rect 3287 17160 3296 17194
rect 3330 17160 3339 17194
rect 3287 17122 3339 17160
rect 3287 17088 3296 17122
rect 3330 17088 3339 17122
rect 3287 17050 3339 17088
rect 3287 17016 3296 17050
rect 3330 17016 3339 17050
rect 3287 16978 3339 17016
rect 3287 16944 3296 16978
rect 3330 16944 3339 16978
rect 3287 16906 3339 16944
rect 3287 16872 3296 16906
rect 3330 16872 3339 16906
rect 3287 16834 3339 16872
rect 3287 16800 3296 16834
rect 3330 16800 3339 16834
rect 3287 16762 3339 16800
rect 3287 16728 3296 16762
rect 3330 16728 3339 16762
rect 3287 16690 3339 16728
rect 3287 16656 3296 16690
rect 3330 16656 3339 16690
rect 3287 16618 3339 16656
rect 3287 16584 3296 16618
rect 3330 16584 3339 16618
rect 3287 16546 3339 16584
rect 3287 16512 3296 16546
rect 3330 16512 3339 16546
rect 3287 16474 3339 16512
rect 3287 16440 3296 16474
rect 3330 16440 3339 16474
rect 3287 16402 3339 16440
rect 3287 16368 3296 16402
rect 3330 16368 3339 16402
rect 3287 16330 3339 16368
rect 3287 16296 3296 16330
rect 3330 16296 3339 16330
rect 3287 16258 3339 16296
rect 3287 16224 3296 16258
rect 3330 16224 3339 16258
rect 3287 16186 3339 16224
rect 3287 16152 3296 16186
rect 3330 16152 3339 16186
rect 3287 16114 3339 16152
rect 3287 16080 3296 16114
rect 3330 16080 3339 16114
rect 3287 16042 3339 16080
rect 3287 16008 3296 16042
rect 3330 16008 3339 16042
rect 3287 15970 3339 16008
rect 3287 15936 3296 15970
rect 3330 15936 3339 15970
rect 3287 15898 3339 15936
rect 3287 15864 3296 15898
rect 3330 15864 3339 15898
rect 3287 15826 3339 15864
rect 3287 15792 3296 15826
rect 3330 15792 3339 15826
rect 3287 15754 3339 15792
rect 3287 15720 3296 15754
rect 3330 15720 3339 15754
rect 3287 15682 3339 15720
rect 3287 15648 3296 15682
rect 3330 15648 3339 15682
rect 3287 15610 3339 15648
rect 3287 15576 3296 15610
rect 3330 15576 3339 15610
rect 3287 15538 3339 15576
rect 3287 15504 3296 15538
rect 3330 15504 3339 15538
rect 3287 15466 3339 15504
rect 3287 15432 3296 15466
rect 3330 15432 3339 15466
rect 3287 15394 3339 15432
rect 3287 15360 3296 15394
rect 3330 15360 3339 15394
rect 3287 15322 3339 15360
rect 3287 15288 3296 15322
rect 3330 15288 3339 15322
rect 3287 15250 3339 15288
rect 3287 15216 3296 15250
rect 3330 15216 3339 15250
rect 3287 15178 3339 15216
rect 3287 15144 3296 15178
rect 3330 15144 3339 15178
rect 3287 15106 3339 15144
rect 3287 15072 3296 15106
rect 3330 15072 3339 15106
rect 3287 15034 3339 15072
rect 3287 15000 3296 15034
rect 3330 15000 3339 15034
rect 3287 14962 3339 15000
rect 3287 14928 3296 14962
rect 3330 14928 3339 14962
rect 3287 14890 3339 14928
rect 3287 14856 3296 14890
rect 3330 14856 3339 14890
rect 3287 14818 3339 14856
rect 3287 14784 3296 14818
rect 3330 14784 3339 14818
rect 3287 14746 3339 14784
rect 3287 14712 3296 14746
rect 3330 14712 3339 14746
rect 3287 14674 3339 14712
rect 3287 14640 3296 14674
rect 3330 14640 3339 14674
rect 3287 14602 3339 14640
rect 3287 14568 3296 14602
rect 3330 14568 3339 14602
rect 3287 14530 3339 14568
rect 3287 14496 3296 14530
rect 3330 14496 3339 14530
rect 3287 14458 3339 14496
rect 3287 14424 3296 14458
rect 3330 14424 3339 14458
rect 3287 14386 3339 14424
rect 3287 14352 3296 14386
rect 3330 14352 3339 14386
rect 3287 14314 3339 14352
rect 3287 14280 3296 14314
rect 3330 14280 3339 14314
rect 3287 14242 3339 14280
rect 3287 14208 3296 14242
rect 3330 14208 3339 14242
rect 3287 14170 3339 14208
rect 3287 14136 3296 14170
rect 3330 14136 3339 14170
rect 3287 14098 3339 14136
rect 3287 14064 3296 14098
rect 3330 14064 3339 14098
rect 3287 14026 3339 14064
rect 3287 13992 3296 14026
rect 3330 13992 3339 14026
rect 3287 13954 3339 13992
rect 3287 13920 3296 13954
rect 3330 13920 3339 13954
rect 3287 13882 3339 13920
rect 3287 13848 3296 13882
rect 3330 13848 3339 13882
rect 3287 13810 3339 13848
rect 3287 13776 3296 13810
rect 3330 13776 3339 13810
rect 3287 13738 3339 13776
rect 3287 13704 3296 13738
rect 3330 13704 3339 13738
rect 3287 13701 3339 13704
rect 3287 13633 3296 13649
rect 3330 13633 3339 13649
rect 3287 13565 3296 13581
rect 3330 13565 3339 13581
rect 3287 13496 3296 13513
rect 3330 13496 3339 13513
rect 3287 13427 3296 13444
rect 3330 13427 3339 13444
rect 3287 13358 3296 13375
rect 3330 13358 3339 13375
rect 3287 13289 3296 13306
rect 3330 13289 3339 13306
rect 3287 13234 3339 13237
rect 3287 13220 3296 13234
rect 3330 13220 3339 13234
rect 3287 13162 3339 13168
rect 3287 13151 3296 13162
rect 3330 13151 3339 13162
rect 3287 13090 3339 13099
rect 3287 13082 3296 13090
rect 3330 13082 3339 13090
rect 3287 13018 3339 13030
rect 3287 13013 3296 13018
rect 3330 13013 3339 13018
rect 3287 12946 3339 12961
rect 3287 12944 3296 12946
rect 3330 12944 3339 12946
rect 3287 12875 3339 12892
rect 3287 12802 3339 12823
rect 3287 12768 3296 12802
rect 3330 12768 3339 12802
rect 3287 12730 3339 12768
rect 3287 12696 3296 12730
rect 3330 12696 3339 12730
rect 3287 12658 3339 12696
rect 3287 12624 3296 12658
rect 3330 12624 3339 12658
rect 3287 12586 3339 12624
rect 3287 12552 3296 12586
rect 3330 12552 3339 12586
rect 3287 12514 3339 12552
rect 3287 12480 3296 12514
rect 3330 12480 3339 12514
rect 3287 12442 3339 12480
rect 3287 12408 3296 12442
rect 3330 12408 3339 12442
rect 3287 12370 3339 12408
rect 3287 12336 3296 12370
rect 3330 12336 3339 12370
rect 3287 12298 3339 12336
rect 3287 12264 3296 12298
rect 3330 12264 3339 12298
rect 3287 12226 3339 12264
rect 3287 12192 3296 12226
rect 3330 12192 3339 12226
rect 3287 12154 3339 12192
rect 3287 12120 3296 12154
rect 3330 12120 3339 12154
rect 3287 12082 3339 12120
rect 3287 12048 3296 12082
rect 3330 12048 3339 12082
rect 3287 12010 3339 12048
rect 3287 11976 3296 12010
rect 3330 11976 3339 12010
rect 3287 11938 3339 11976
rect 3287 11904 3296 11938
rect 3330 11904 3339 11938
rect 3287 11866 3339 11904
rect 3287 11832 3296 11866
rect 3330 11832 3339 11866
rect 3287 11794 3339 11832
rect 3287 11760 3296 11794
rect 3330 11760 3339 11794
rect 3287 11722 3339 11760
rect 3287 11688 3296 11722
rect 3330 11688 3339 11722
rect 3287 11650 3339 11688
rect 3287 11616 3296 11650
rect 3330 11616 3339 11650
rect 3287 11578 3339 11616
rect 3287 11544 3296 11578
rect 3330 11544 3339 11578
rect 3287 11506 3339 11544
rect 3287 11472 3296 11506
rect 3330 11472 3339 11506
rect 3287 11434 3339 11472
rect 3287 11400 3296 11434
rect 3330 11400 3339 11434
rect 3287 11362 3339 11400
rect 3287 11328 3296 11362
rect 3330 11328 3339 11362
rect 3287 11290 3339 11328
rect 3287 11256 3296 11290
rect 3330 11256 3339 11290
rect 3287 11218 3339 11256
rect 3287 11184 3296 11218
rect 3330 11184 3339 11218
rect 3287 11146 3339 11184
rect 3287 11112 3296 11146
rect 3330 11112 3339 11146
rect 3287 11074 3339 11112
rect 3287 11040 3296 11074
rect 3330 11040 3339 11074
rect 3287 11002 3339 11040
rect 3287 10968 3296 11002
rect 3330 10968 3339 11002
rect 3287 10930 3339 10968
rect 3287 10896 3296 10930
rect 3330 10896 3339 10930
rect 3287 10858 3339 10896
rect 3287 10824 3296 10858
rect 3330 10824 3339 10858
rect 3287 10786 3339 10824
rect 3287 10752 3296 10786
rect 3330 10752 3339 10786
rect 3287 10714 3339 10752
rect 3287 10680 3296 10714
rect 3330 10680 3339 10714
rect 3287 10642 3339 10680
rect 3287 10608 3296 10642
rect 3330 10608 3339 10642
rect 3287 10570 3339 10608
rect 3287 10536 3296 10570
rect 3330 10536 3339 10570
rect 3287 10498 3339 10536
rect 3287 10464 3296 10498
rect 3330 10464 3339 10498
rect 3287 10426 3339 10464
rect 3287 10392 3296 10426
rect 3330 10392 3339 10426
rect 3287 10354 3339 10392
rect 3287 10320 3296 10354
rect 3330 10320 3339 10354
rect 3287 10282 3339 10320
rect 3287 10248 3296 10282
rect 3330 10248 3339 10282
rect 3287 10210 3339 10248
rect 3287 10176 3296 10210
rect 3330 10176 3339 10210
rect 3287 10138 3339 10176
rect 3287 10104 3296 10138
rect 3330 10104 3339 10138
rect 3287 10066 3339 10104
rect 3287 10032 3296 10066
rect 3330 10032 3339 10066
rect 3287 9994 3339 10032
rect 3287 9960 3296 9994
rect 3330 9960 3339 9994
rect 3287 9922 3339 9960
rect 3287 9888 3296 9922
rect 3330 9888 3339 9922
rect 3287 9850 3339 9888
rect 3287 9816 3296 9850
rect 3330 9816 3339 9850
rect 3287 9778 3339 9816
rect 3287 9744 3296 9778
rect 3330 9744 3339 9778
rect 3287 9706 3339 9744
rect 3287 9672 3296 9706
rect 3330 9672 3339 9706
rect 3287 9634 3339 9672
rect 3287 9600 3296 9634
rect 3330 9600 3339 9634
rect 3287 9562 3339 9600
rect 3287 9528 3296 9562
rect 3330 9528 3339 9562
rect 3287 9490 3339 9528
rect 3287 9456 3296 9490
rect 3330 9456 3339 9490
rect 3287 9418 3339 9456
rect 3287 9384 3296 9418
rect 3330 9384 3339 9418
rect 3287 9346 3339 9384
rect 3287 9312 3296 9346
rect 3330 9312 3339 9346
rect 3287 9274 3339 9312
rect 3287 9240 3296 9274
rect 3330 9240 3339 9274
rect 3287 9202 3339 9240
rect 3287 9168 3296 9202
rect 3330 9168 3339 9202
rect 3287 9130 3339 9168
rect 3287 9096 3296 9130
rect 3330 9096 3339 9130
rect 3287 9058 3339 9096
rect 3287 9024 3296 9058
rect 3330 9024 3339 9058
rect 3287 8986 3339 9024
rect 3287 8952 3296 8986
rect 3330 8952 3339 8986
rect 3287 8914 3339 8952
rect 3287 8880 3296 8914
rect 3330 8880 3339 8914
rect 3287 8842 3339 8880
rect 3287 8808 3296 8842
rect 3330 8808 3339 8842
rect 3287 8770 3339 8808
rect 3287 8736 3296 8770
rect 3330 8736 3339 8770
rect 3287 8698 3339 8736
rect 3287 8664 3296 8698
rect 3330 8664 3339 8698
rect 3287 8626 3339 8664
rect 3287 8592 3296 8626
rect 3330 8592 3339 8626
rect 3287 8554 3339 8592
rect 3287 8520 3296 8554
rect 3330 8520 3339 8554
rect 3287 8482 3339 8520
rect 3287 8448 3296 8482
rect 3330 8448 3339 8482
rect 3287 8410 3339 8448
rect 3287 8376 3296 8410
rect 3330 8376 3339 8410
rect 3287 8338 3339 8376
rect 3287 8304 3296 8338
rect 3330 8304 3339 8338
rect 3287 8266 3339 8304
rect 3287 8232 3296 8266
rect 3330 8232 3339 8266
rect 3287 8194 3339 8232
rect 3287 8160 3296 8194
rect 3330 8160 3339 8194
rect 3287 8122 3339 8160
rect 3287 8088 3296 8122
rect 3330 8088 3339 8122
rect 3287 8050 3339 8088
rect 3287 8016 3296 8050
rect 3330 8016 3339 8050
rect 3287 7978 3339 8016
rect 3287 7944 3296 7978
rect 3330 7944 3339 7978
rect 3287 7906 3339 7944
rect 3287 7872 3296 7906
rect 3330 7872 3339 7906
rect 3287 7834 3339 7872
rect 3287 7800 3296 7834
rect 3330 7800 3339 7834
rect 3287 7762 3339 7800
rect 3287 7728 3296 7762
rect 3330 7728 3339 7762
rect 3287 7690 3339 7728
rect 3287 7656 3296 7690
rect 3330 7656 3339 7690
rect 3287 7618 3339 7656
rect 3287 7584 3296 7618
rect 3330 7584 3339 7618
rect 3287 7546 3339 7584
rect 3287 7512 3296 7546
rect 3330 7512 3339 7546
rect 3287 7474 3339 7512
rect 3287 7440 3296 7474
rect 3330 7440 3339 7474
rect 3287 7402 3339 7440
rect 3287 7368 3296 7402
rect 3330 7368 3339 7402
rect 3287 7330 3339 7368
rect 3287 7296 3296 7330
rect 3330 7296 3339 7330
rect 3287 7258 3339 7296
rect 3287 7224 3296 7258
rect 3330 7224 3339 7258
rect 3287 7186 3339 7224
rect 3287 7152 3296 7186
rect 3330 7152 3339 7186
rect 3287 7114 3339 7152
rect 3287 7080 3296 7114
rect 3330 7080 3339 7114
rect 3287 7042 3339 7080
rect 3287 7008 3296 7042
rect 3330 7008 3339 7042
rect 3287 6970 3339 7008
rect 3287 6936 3296 6970
rect 3330 6936 3339 6970
rect 3287 6898 3339 6936
rect 3287 6864 3296 6898
rect 3330 6864 3339 6898
rect 3287 6826 3339 6864
rect 3287 6792 3296 6826
rect 3330 6792 3339 6826
rect 3287 6754 3339 6792
rect 3287 6720 3296 6754
rect 3330 6720 3339 6754
rect 3287 6682 3339 6720
rect 3287 6648 3296 6682
rect 3330 6648 3339 6682
rect 3287 6610 3339 6648
rect 3287 6576 3296 6610
rect 3330 6576 3339 6610
rect 3287 6538 3339 6576
rect 3287 6504 3296 6538
rect 3330 6504 3339 6538
rect 3287 6466 3339 6504
rect 3287 6432 3296 6466
rect 3330 6432 3339 6466
rect 3287 6394 3339 6432
rect 3287 6360 3296 6394
rect 3330 6360 3339 6394
rect 3287 6322 3339 6360
rect 3287 6288 3296 6322
rect 3330 6288 3339 6322
rect 3287 6250 3339 6288
rect 3287 6216 3296 6250
rect 3330 6216 3339 6250
rect 3287 6178 3339 6216
rect 3287 6144 3296 6178
rect 3330 6144 3339 6178
rect 3287 6106 3339 6144
rect 3287 6072 3296 6106
rect 3330 6072 3339 6106
rect 3287 6034 3339 6072
rect 3287 6000 3296 6034
rect 3330 6000 3339 6034
rect 3287 5962 3339 6000
rect 3287 5928 3296 5962
rect 3330 5928 3339 5962
rect 3287 5890 3339 5928
rect 3287 5856 3296 5890
rect 3330 5856 3339 5890
rect 3287 5818 3339 5856
rect 3287 5784 3296 5818
rect 3330 5784 3339 5818
rect 3287 5746 3339 5784
rect 3287 5712 3296 5746
rect 3330 5712 3339 5746
rect 3287 5674 3339 5712
rect 3287 5640 3296 5674
rect 3330 5640 3339 5674
rect 3287 5602 3339 5640
rect 3287 5568 3296 5602
rect 3330 5568 3339 5602
rect 3287 5530 3339 5568
rect 3287 5496 3296 5530
rect 3330 5496 3339 5530
rect 3287 5458 3339 5496
rect 3287 5424 3296 5458
rect 3330 5424 3339 5458
rect 3287 5386 3339 5424
rect 3287 5352 3296 5386
rect 3330 5352 3339 5386
rect 3287 5314 3339 5352
rect 3287 5280 3296 5314
rect 3330 5280 3339 5314
rect 3287 5242 3339 5280
rect 3287 5208 3296 5242
rect 3330 5208 3339 5242
rect 3287 5170 3339 5208
rect 3287 5136 3296 5170
rect 3330 5136 3339 5170
rect 3287 5098 3339 5136
rect 3287 5064 3296 5098
rect 3330 5064 3339 5098
rect 3287 5026 3339 5064
rect 3287 4992 3296 5026
rect 3330 4992 3339 5026
rect 3287 4954 3339 4992
rect 3287 4920 3296 4954
rect 3330 4920 3339 4954
rect 3287 4882 3339 4920
rect 3287 4848 3296 4882
rect 3330 4848 3339 4882
rect 3287 4810 3339 4848
rect 3287 4776 3296 4810
rect 3330 4776 3339 4810
rect 3287 4738 3339 4776
rect 3287 4704 3296 4738
rect 3330 4704 3339 4738
rect 3287 4666 3339 4704
rect 3287 4632 3296 4666
rect 3330 4632 3339 4666
rect 3287 4594 3339 4632
rect 3287 4560 3296 4594
rect 3330 4560 3339 4594
rect 3287 4522 3339 4560
rect 3287 4488 3296 4522
rect 3330 4488 3339 4522
rect 3287 4450 3339 4488
rect 3287 4416 3296 4450
rect 3330 4416 3339 4450
rect 3287 4378 3339 4416
rect 3287 4344 3296 4378
rect 3330 4344 3339 4378
rect 3287 4306 3339 4344
rect 3287 4272 3296 4306
rect 3330 4272 3339 4306
rect 3287 4234 3339 4272
rect 3287 4200 3296 4234
rect 3330 4200 3339 4234
rect 3287 4162 3339 4200
rect 3287 4128 3296 4162
rect 3330 4128 3339 4162
rect 3287 4090 3339 4128
rect 3287 4056 3296 4090
rect 3330 4056 3339 4090
rect 3287 4018 3339 4056
rect 3287 3984 3296 4018
rect 3330 3984 3339 4018
rect 3287 3946 3339 3984
rect 3287 3912 3296 3946
rect 3330 3912 3339 3946
rect 3287 3874 3339 3912
rect 3287 3840 3296 3874
rect 3330 3840 3339 3874
rect 3287 3802 3339 3840
rect 3287 3768 3296 3802
rect 3330 3768 3339 3802
rect 3287 3730 3339 3768
rect 3287 3696 3296 3730
rect 3330 3696 3339 3730
rect 3287 3658 3339 3696
rect 3287 3624 3296 3658
rect 3330 3624 3339 3658
rect 3287 3586 3339 3624
rect 3287 3552 3296 3586
rect 3330 3552 3339 3586
rect 3287 3514 3339 3552
rect 3287 3480 3296 3514
rect 3330 3480 3339 3514
rect 3287 3442 3339 3480
rect 3287 3408 3296 3442
rect 3330 3408 3339 3442
rect 3287 3370 3339 3408
rect 3287 3336 3296 3370
rect 3330 3336 3339 3370
rect 3287 3298 3339 3336
rect 3287 3264 3296 3298
rect 3330 3264 3339 3298
rect 3287 3225 3339 3264
rect 3287 3191 3296 3225
rect 3330 3191 3339 3225
rect 3287 3152 3339 3191
rect 3287 3118 3296 3152
rect 3330 3118 3339 3152
rect 3287 3079 3339 3118
rect 3287 3045 3296 3079
rect 3330 3045 3339 3079
rect 3287 3006 3339 3045
rect 3287 2972 3296 3006
rect 3330 2972 3339 3006
rect 3287 2933 3339 2972
rect 3287 2899 3296 2933
rect 3330 2899 3339 2933
rect 3287 2860 3339 2899
rect 3287 2826 3296 2860
rect 3330 2826 3339 2860
rect 3287 2787 3339 2826
rect 3287 2753 3296 2787
rect 3330 2753 3339 2787
rect 3287 2714 3339 2753
rect 3287 2680 3296 2714
rect 3330 2680 3339 2714
rect 3287 2641 3339 2680
rect 3287 2607 3296 2641
rect 3330 2607 3339 2641
rect 3287 2568 3339 2607
rect 3287 2534 3296 2568
rect 3330 2534 3339 2568
rect 3287 2495 3339 2534
rect 3287 2461 3296 2495
rect 3330 2461 3339 2495
rect 3287 2422 3339 2461
rect 3287 2388 3296 2422
rect 3330 2388 3339 2422
rect 3287 2349 3339 2388
rect 3287 2315 3296 2349
rect 3330 2315 3339 2349
rect 3287 2276 3339 2315
rect 3287 2242 3296 2276
rect 3330 2242 3339 2276
rect 3287 2203 3339 2242
rect 3287 2169 3296 2203
rect 3330 2169 3339 2203
rect 3287 2130 3339 2169
rect 3287 2096 3296 2130
rect 3330 2096 3339 2130
rect 3287 2057 3339 2096
rect 3287 2023 3296 2057
rect 3330 2023 3339 2057
rect 3287 1984 3339 2023
rect 3287 1950 3296 1984
rect 3330 1950 3339 1984
rect 3287 1911 3339 1950
rect 3287 1877 3296 1911
rect 3330 1877 3339 1911
rect 3287 1838 3339 1877
rect 3287 1804 3296 1838
rect 3330 1804 3339 1838
rect 3287 1765 3339 1804
rect 3287 1731 3296 1765
rect 3330 1731 3339 1765
rect 3287 1692 3339 1731
rect 3287 1658 3296 1692
rect 3330 1658 3339 1692
rect 3287 1619 3339 1658
rect 3287 1585 3296 1619
rect 3330 1585 3339 1619
rect 3287 1546 3339 1585
rect 3287 1512 3296 1546
rect 3330 1512 3339 1546
rect 3287 1473 3339 1512
rect 3287 1439 3296 1473
rect 3330 1439 3339 1473
rect 3287 1400 3339 1439
rect 3287 1366 3296 1400
rect 3330 1366 3339 1400
rect 3287 1327 3339 1366
rect 3287 1293 3296 1327
rect 3330 1293 3339 1327
rect 3287 1254 3339 1293
rect 3287 1220 3296 1254
rect 3330 1220 3339 1254
rect 3287 1181 3339 1220
rect 3287 1147 3296 1181
rect 3330 1147 3339 1181
rect 3287 1108 3339 1147
rect 3287 1074 3296 1108
rect 3330 1074 3339 1108
rect 3287 1035 3339 1074
rect 3287 1001 3296 1035
rect 3330 1001 3339 1035
rect 3287 962 3339 1001
rect 3287 928 3296 962
rect 3330 928 3339 962
rect 3287 889 3339 928
rect 3287 855 3296 889
rect 3330 855 3339 889
rect 3287 816 3339 855
rect 3287 782 3296 816
rect 3330 782 3339 816
rect 3287 743 3339 782
rect 3287 709 3296 743
rect 3330 709 3339 743
rect 3287 670 3339 709
rect 3287 636 3296 670
rect 3330 636 3339 670
rect 3287 597 3339 636
rect 3287 563 3296 597
rect 3330 563 3339 597
rect 117 486 126 520
rect 160 486 169 520
rect 117 448 169 486
rect 117 414 126 448
rect 160 414 169 448
rect 117 376 169 414
rect 117 342 126 376
rect 160 342 169 376
rect 117 304 169 342
rect 117 270 126 304
rect 160 270 169 304
rect 117 232 169 270
rect 117 198 126 232
rect 160 198 169 232
rect 3287 524 3339 563
rect 3287 490 3296 524
rect 3330 490 3339 524
rect 3287 451 3339 490
rect 3287 417 3296 451
rect 3330 417 3339 451
rect 3287 378 3339 417
rect 3287 344 3296 378
rect 3330 344 3339 378
rect 3287 305 3339 344
rect 3287 271 3296 305
rect 3330 271 3339 305
rect 3287 232 3339 271
tri 169 198 171 200 sw
tri 3285 198 3287 200 se
rect 3287 198 3296 232
rect 3330 198 3339 232
rect 117 166 171 198
tri 171 166 203 198 sw
tri 3253 166 3285 198 se
rect 3285 166 3339 198
rect 117 160 3339 166
rect 117 126 198 160
rect 232 126 271 160
rect 305 126 344 160
rect 378 126 416 160
rect 450 126 488 160
rect 522 126 560 160
rect 594 126 632 160
rect 666 126 704 160
rect 738 126 776 160
rect 810 126 848 160
rect 882 126 920 160
rect 954 126 992 160
rect 1026 126 1064 160
rect 1098 126 1136 160
rect 1170 126 1208 160
rect 1242 126 1280 160
rect 1314 126 1352 160
rect 1386 126 1424 160
rect 1458 126 1496 160
rect 1530 126 1568 160
rect 1602 126 1640 160
rect 1674 126 1712 160
rect 1746 126 1784 160
rect 1818 126 1856 160
rect 1890 126 1928 160
rect 1962 126 2000 160
rect 2034 126 2072 160
rect 2106 126 2144 160
rect 2178 126 2216 160
rect 2250 126 2288 160
rect 2322 126 2360 160
rect 2394 126 2432 160
rect 2466 126 2504 160
rect 2538 126 2576 160
rect 2610 126 2648 160
rect 2682 126 2720 160
rect 2754 126 2792 160
rect 2826 126 2864 160
rect 2898 126 2936 160
rect 2970 126 3008 160
rect 3042 126 3080 160
rect 3114 126 3152 160
rect 3186 126 3224 160
rect 3258 126 3339 160
rect 117 120 3339 126
<< via1 >>
rect 117 13696 169 13701
rect 117 13662 126 13696
rect 126 13662 160 13696
rect 160 13662 169 13696
rect 117 13649 169 13662
rect 117 13624 169 13633
rect 117 13590 126 13624
rect 126 13590 160 13624
rect 160 13590 169 13624
rect 117 13581 169 13590
rect 117 13552 169 13565
rect 117 13518 126 13552
rect 126 13518 160 13552
rect 160 13518 169 13552
rect 117 13513 169 13518
rect 117 13480 169 13496
rect 117 13446 126 13480
rect 126 13446 160 13480
rect 160 13446 169 13480
rect 117 13444 169 13446
rect 117 13408 169 13427
rect 117 13375 126 13408
rect 126 13375 160 13408
rect 160 13375 169 13408
rect 117 13336 169 13358
rect 117 13306 126 13336
rect 126 13306 160 13336
rect 160 13306 169 13336
rect 117 13264 169 13289
rect 117 13237 126 13264
rect 126 13237 160 13264
rect 160 13237 169 13264
rect 117 13192 169 13220
rect 117 13168 126 13192
rect 126 13168 160 13192
rect 160 13168 169 13192
rect 117 13120 169 13151
rect 117 13099 126 13120
rect 126 13099 160 13120
rect 160 13099 169 13120
rect 117 13048 169 13082
rect 117 13030 126 13048
rect 126 13030 160 13048
rect 160 13030 169 13048
rect 117 12976 169 13013
rect 117 12961 126 12976
rect 126 12961 160 12976
rect 160 12961 169 12976
rect 117 12942 126 12944
rect 126 12942 160 12944
rect 160 12942 169 12944
rect 117 12904 169 12942
rect 117 12892 126 12904
rect 126 12892 160 12904
rect 160 12892 169 12904
rect 117 12870 126 12875
rect 126 12870 160 12875
rect 160 12870 169 12875
rect 117 12832 169 12870
rect 117 12823 126 12832
rect 126 12823 160 12832
rect 160 12823 169 12832
rect 1501 39011 1553 39063
rect 1569 39011 1621 39063
rect 1636 39011 1688 39063
rect 1703 39011 1755 39063
rect 1770 39011 1822 39063
rect 1837 39011 1889 39063
rect 697 38371 749 38423
rect 765 38419 767 38423
rect 767 38419 801 38423
rect 801 38419 817 38423
rect 765 38380 817 38419
rect 765 38371 767 38380
rect 767 38371 801 38380
rect 801 38371 817 38380
rect 833 38371 885 38423
rect 901 38371 953 38423
rect 969 38419 1003 38423
rect 1003 38419 1021 38423
rect 969 38380 1021 38419
rect 969 38371 1003 38380
rect 1003 38371 1021 38380
rect 1037 38371 1089 38423
rect 1105 38371 1157 38423
rect 1173 38371 1225 38423
rect 1241 38419 1273 38423
rect 1273 38419 1293 38423
rect 1241 38380 1293 38419
rect 1241 38371 1273 38380
rect 1273 38371 1293 38380
rect 697 38307 749 38359
rect 765 38346 767 38359
rect 767 38346 801 38359
rect 801 38346 817 38359
rect 765 38307 817 38346
rect 833 38307 885 38359
rect 901 38307 953 38359
rect 969 38346 1003 38359
rect 1003 38346 1021 38359
rect 969 38307 1021 38346
rect 1037 38307 1089 38359
rect 1105 38307 1157 38359
rect 1173 38307 1225 38359
rect 1241 38346 1273 38359
rect 1273 38346 1293 38359
rect 2097 38371 2149 38423
rect 2165 38419 2183 38423
rect 2183 38419 2217 38423
rect 2165 38380 2217 38419
rect 2165 38371 2183 38380
rect 2183 38371 2217 38380
rect 2233 38371 2285 38423
rect 2301 38371 2353 38423
rect 2369 38419 2419 38423
rect 2419 38419 2421 38423
rect 2437 38419 2453 38423
rect 2453 38419 2489 38423
rect 2369 38380 2421 38419
rect 2437 38380 2489 38419
rect 2369 38371 2419 38380
rect 2419 38371 2421 38380
rect 2437 38371 2453 38380
rect 2453 38371 2489 38380
rect 2505 38371 2557 38423
rect 2573 38371 2625 38423
rect 2641 38419 2655 38423
rect 2655 38419 2689 38423
rect 2689 38419 2693 38423
rect 2641 38380 2693 38419
rect 2641 38371 2655 38380
rect 2655 38371 2689 38380
rect 2689 38371 2693 38380
rect 1241 38307 1293 38346
rect 2097 38307 2149 38359
rect 2165 38346 2183 38359
rect 2183 38346 2217 38359
rect 2165 38307 2217 38346
rect 2233 38307 2285 38359
rect 2301 38307 2353 38359
rect 2369 38346 2419 38359
rect 2419 38346 2421 38359
rect 2437 38346 2453 38359
rect 2453 38346 2489 38359
rect 2369 38307 2421 38346
rect 2437 38307 2489 38346
rect 2505 38307 2557 38359
rect 2573 38307 2625 38359
rect 2641 38346 2655 38359
rect 2655 38346 2689 38359
rect 2689 38346 2693 38359
rect 2641 38307 2693 38346
rect 697 38243 749 38295
rect 765 38273 767 38295
rect 767 38273 801 38295
rect 801 38273 817 38295
rect 765 38243 817 38273
rect 833 38243 885 38295
rect 901 38243 953 38295
rect 969 38273 1003 38295
rect 1003 38273 1021 38295
rect 969 38243 1021 38273
rect 1037 38243 1089 38295
rect 1105 38243 1157 38295
rect 1173 38243 1225 38295
rect 1241 38273 1273 38295
rect 1273 38273 1293 38295
rect 1241 38243 1293 38273
rect 2097 38243 2149 38295
rect 2165 38273 2183 38295
rect 2183 38273 2217 38295
rect 2165 38243 2217 38273
rect 2233 38243 2285 38295
rect 2301 38243 2353 38295
rect 2369 38273 2419 38295
rect 2419 38273 2421 38295
rect 2437 38273 2453 38295
rect 2453 38273 2489 38295
rect 2369 38243 2421 38273
rect 2437 38243 2489 38273
rect 2505 38243 2557 38295
rect 2573 38243 2625 38295
rect 2641 38273 2655 38295
rect 2655 38273 2689 38295
rect 2689 38273 2693 38295
rect 2641 38243 2693 38273
rect 697 38179 749 38231
rect 765 38200 767 38231
rect 767 38200 801 38231
rect 801 38200 817 38231
rect 765 38179 817 38200
rect 833 38179 885 38231
rect 901 38179 953 38231
rect 969 38200 1003 38231
rect 1003 38200 1021 38231
rect 969 38179 1021 38200
rect 1037 38179 1089 38231
rect 1105 38179 1157 38231
rect 1173 38179 1225 38231
rect 1241 38200 1273 38231
rect 1273 38200 1293 38231
rect 1241 38179 1293 38200
rect 2097 38179 2149 38231
rect 2165 38200 2183 38231
rect 2183 38200 2217 38231
rect 2165 38179 2217 38200
rect 2233 38179 2285 38231
rect 2301 38179 2353 38231
rect 2369 38200 2419 38231
rect 2419 38200 2421 38231
rect 2437 38200 2453 38231
rect 2453 38200 2489 38231
rect 2369 38179 2421 38200
rect 2437 38179 2489 38200
rect 2505 38179 2557 38231
rect 2573 38179 2625 38231
rect 2641 38200 2655 38231
rect 2655 38200 2689 38231
rect 2689 38200 2693 38231
rect 2641 38179 2693 38200
rect 697 38115 749 38167
rect 765 38161 817 38167
rect 765 38127 767 38161
rect 767 38127 801 38161
rect 801 38127 817 38161
rect 765 38115 817 38127
rect 833 38115 885 38167
rect 901 38115 953 38167
rect 969 38161 1021 38167
rect 969 38127 1003 38161
rect 1003 38127 1021 38161
rect 969 38115 1021 38127
rect 1037 38115 1089 38167
rect 1105 38115 1157 38167
rect 1173 38115 1225 38167
rect 1241 38161 1293 38167
rect 1241 38127 1273 38161
rect 1273 38127 1293 38161
rect 1241 38115 1293 38127
rect 2097 38115 2149 38167
rect 2165 38161 2217 38167
rect 2165 38127 2183 38161
rect 2183 38127 2217 38161
rect 2165 38115 2217 38127
rect 2233 38115 2285 38167
rect 2301 38115 2353 38167
rect 2369 38161 2421 38167
rect 2437 38161 2489 38167
rect 2369 38127 2419 38161
rect 2419 38127 2421 38161
rect 2437 38127 2453 38161
rect 2453 38127 2489 38161
rect 2369 38115 2421 38127
rect 2437 38115 2489 38127
rect 2505 38115 2557 38167
rect 2573 38115 2625 38167
rect 2641 38161 2693 38167
rect 2641 38127 2655 38161
rect 2655 38127 2689 38161
rect 2689 38127 2693 38161
rect 2641 38115 2693 38127
rect 697 38051 749 38103
rect 765 38088 817 38103
rect 765 38054 767 38088
rect 767 38054 801 38088
rect 801 38054 817 38088
rect 765 38051 817 38054
rect 833 38051 885 38103
rect 901 38051 953 38103
rect 969 38088 1021 38103
rect 969 38054 1003 38088
rect 1003 38054 1021 38088
rect 969 38051 1021 38054
rect 1037 38051 1089 38103
rect 1105 38051 1157 38103
rect 1173 38051 1225 38103
rect 1241 38088 1293 38103
rect 1241 38054 1273 38088
rect 1273 38054 1293 38088
rect 1241 38051 1293 38054
rect 2097 38051 2149 38103
rect 2165 38088 2217 38103
rect 2165 38054 2183 38088
rect 2183 38054 2217 38088
rect 2165 38051 2217 38054
rect 2233 38051 2285 38103
rect 2301 38051 2353 38103
rect 2369 38088 2421 38103
rect 2437 38088 2489 38103
rect 2369 38054 2419 38088
rect 2419 38054 2421 38088
rect 2437 38054 2453 38088
rect 2453 38054 2489 38088
rect 2369 38051 2421 38054
rect 2437 38051 2489 38054
rect 2505 38051 2557 38103
rect 2573 38051 2625 38103
rect 2641 38088 2693 38103
rect 2641 38054 2655 38088
rect 2655 38054 2689 38088
rect 2689 38054 2693 38088
rect 2641 38051 2693 38054
rect 697 37987 749 38039
rect 765 38014 817 38039
rect 765 37987 767 38014
rect 767 37987 801 38014
rect 801 37987 817 38014
rect 833 37987 885 38039
rect 901 37987 953 38039
rect 969 38014 1021 38039
rect 969 37987 1003 38014
rect 1003 37987 1021 38014
rect 1037 37987 1089 38039
rect 1105 37987 1157 38039
rect 1173 37987 1225 38039
rect 1241 38014 1293 38039
rect 1241 37987 1273 38014
rect 1273 37987 1293 38014
rect 2097 37987 2149 38039
rect 2165 38014 2217 38039
rect 2165 37987 2183 38014
rect 2183 37987 2217 38014
rect 2233 37987 2285 38039
rect 2301 37987 2353 38039
rect 2369 38014 2421 38039
rect 2437 38014 2489 38039
rect 2369 37987 2419 38014
rect 2419 37987 2421 38014
rect 2437 37987 2453 38014
rect 2453 37987 2489 38014
rect 2505 37987 2557 38039
rect 2573 37987 2625 38039
rect 2641 38014 2693 38039
rect 2641 37987 2655 38014
rect 2655 37987 2689 38014
rect 2689 37987 2693 38014
rect 697 37923 749 37975
rect 765 37940 817 37975
rect 765 37923 767 37940
rect 767 37923 801 37940
rect 801 37923 817 37940
rect 833 37923 885 37975
rect 901 37923 953 37975
rect 969 37940 1021 37975
rect 969 37923 1003 37940
rect 1003 37923 1021 37940
rect 1037 37923 1089 37975
rect 1105 37923 1157 37975
rect 1173 37923 1225 37975
rect 1241 37940 1293 37975
rect 1241 37923 1273 37940
rect 1273 37923 1293 37940
rect 697 37859 749 37911
rect 765 37906 767 37911
rect 767 37906 801 37911
rect 801 37906 817 37911
rect 765 37866 817 37906
rect 765 37859 767 37866
rect 767 37859 801 37866
rect 801 37859 817 37866
rect 833 37859 885 37911
rect 901 37859 953 37911
rect 969 37906 1003 37911
rect 1003 37906 1021 37911
rect 969 37866 1021 37906
rect 969 37859 1003 37866
rect 1003 37859 1021 37866
rect 1037 37859 1089 37911
rect 1105 37859 1157 37911
rect 1173 37859 1225 37911
rect 1241 37906 1273 37911
rect 1273 37906 1293 37911
rect 2097 37923 2149 37975
rect 2165 37940 2217 37975
rect 2165 37923 2183 37940
rect 2183 37923 2217 37940
rect 2233 37923 2285 37975
rect 2301 37923 2353 37975
rect 2369 37940 2421 37975
rect 2437 37940 2489 37975
rect 2369 37923 2419 37940
rect 2419 37923 2421 37940
rect 2437 37923 2453 37940
rect 2453 37923 2489 37940
rect 2505 37923 2557 37975
rect 2573 37923 2625 37975
rect 2641 37940 2693 37975
rect 2641 37923 2655 37940
rect 2655 37923 2689 37940
rect 2689 37923 2693 37940
rect 1241 37866 1293 37906
rect 1241 37859 1273 37866
rect 1273 37859 1293 37866
rect 697 37795 749 37847
rect 765 37832 767 37847
rect 767 37832 801 37847
rect 801 37832 817 37847
rect 765 37795 817 37832
rect 833 37795 885 37847
rect 901 37795 953 37847
rect 969 37832 1003 37847
rect 1003 37832 1021 37847
rect 969 37795 1021 37832
rect 1037 37795 1089 37847
rect 1105 37795 1157 37847
rect 1173 37795 1225 37847
rect 1241 37832 1273 37847
rect 1273 37832 1293 37847
rect 2097 37859 2149 37911
rect 2165 37906 2183 37911
rect 2183 37906 2217 37911
rect 2165 37866 2217 37906
rect 2165 37859 2183 37866
rect 2183 37859 2217 37866
rect 2233 37859 2285 37911
rect 2301 37859 2353 37911
rect 2369 37906 2419 37911
rect 2419 37906 2421 37911
rect 2437 37906 2453 37911
rect 2453 37906 2489 37911
rect 2369 37866 2421 37906
rect 2437 37866 2489 37906
rect 2369 37859 2419 37866
rect 2419 37859 2421 37866
rect 2437 37859 2453 37866
rect 2453 37859 2489 37866
rect 2505 37859 2557 37911
rect 2573 37859 2625 37911
rect 2641 37906 2655 37911
rect 2655 37906 2689 37911
rect 2689 37906 2693 37911
rect 2641 37866 2693 37906
rect 2641 37859 2655 37866
rect 2655 37859 2689 37866
rect 2689 37859 2693 37866
rect 1241 37795 1293 37832
rect 2097 37795 2149 37847
rect 2165 37832 2183 37847
rect 2183 37832 2217 37847
rect 2165 37795 2217 37832
rect 2233 37795 2285 37847
rect 2301 37795 2353 37847
rect 2369 37832 2419 37847
rect 2419 37832 2421 37847
rect 2437 37832 2453 37847
rect 2453 37832 2489 37847
rect 2369 37795 2421 37832
rect 2437 37795 2489 37832
rect 2505 37795 2557 37847
rect 2573 37795 2625 37847
rect 2641 37832 2655 37847
rect 2655 37832 2689 37847
rect 2689 37832 2693 37847
rect 2641 37795 2693 37832
rect 697 37731 749 37783
rect 765 37758 767 37783
rect 767 37758 801 37783
rect 801 37758 817 37783
rect 765 37731 817 37758
rect 833 37731 885 37783
rect 901 37731 953 37783
rect 969 37758 1003 37783
rect 1003 37758 1021 37783
rect 969 37731 1021 37758
rect 1037 37731 1089 37783
rect 1105 37731 1157 37783
rect 1173 37731 1225 37783
rect 1241 37758 1273 37783
rect 1273 37758 1293 37783
rect 1241 37731 1293 37758
rect 2097 37731 2149 37783
rect 2165 37758 2183 37783
rect 2183 37758 2217 37783
rect 2165 37731 2217 37758
rect 2233 37731 2285 37783
rect 2301 37731 2353 37783
rect 2369 37758 2419 37783
rect 2419 37758 2421 37783
rect 2437 37758 2453 37783
rect 2453 37758 2489 37783
rect 2369 37731 2421 37758
rect 2437 37731 2489 37758
rect 2505 37731 2557 37783
rect 2573 37731 2625 37783
rect 2641 37758 2655 37783
rect 2655 37758 2689 37783
rect 2689 37758 2693 37783
rect 2641 37731 2693 37758
rect 697 37667 749 37719
rect 765 37718 817 37719
rect 765 37684 767 37718
rect 767 37684 801 37718
rect 801 37684 817 37718
rect 765 37667 817 37684
rect 833 37667 885 37719
rect 901 37667 953 37719
rect 969 37718 1021 37719
rect 969 37684 1003 37718
rect 1003 37684 1021 37718
rect 969 37667 1021 37684
rect 1037 37667 1089 37719
rect 1105 37667 1157 37719
rect 1173 37667 1225 37719
rect 1241 37718 1293 37719
rect 1241 37684 1273 37718
rect 1273 37684 1293 37718
rect 1241 37667 1293 37684
rect 2097 37667 2149 37719
rect 2165 37718 2217 37719
rect 2165 37684 2183 37718
rect 2183 37684 2217 37718
rect 2165 37667 2217 37684
rect 2233 37667 2285 37719
rect 2301 37667 2353 37719
rect 2369 37718 2421 37719
rect 2437 37718 2489 37719
rect 2369 37684 2419 37718
rect 2419 37684 2421 37718
rect 2437 37684 2453 37718
rect 2453 37684 2489 37718
rect 2369 37667 2421 37684
rect 2437 37667 2489 37684
rect 2505 37667 2557 37719
rect 2573 37667 2625 37719
rect 2641 37718 2693 37719
rect 2641 37684 2655 37718
rect 2655 37684 2689 37718
rect 2689 37684 2693 37718
rect 2641 37667 2693 37684
rect 697 37603 749 37655
rect 765 37644 817 37655
rect 765 37610 767 37644
rect 767 37610 801 37644
rect 801 37610 817 37644
rect 765 37603 817 37610
rect 833 37603 885 37655
rect 901 37603 953 37655
rect 969 37644 1021 37655
rect 969 37610 1003 37644
rect 1003 37610 1021 37644
rect 969 37603 1021 37610
rect 1037 37603 1089 37655
rect 1105 37603 1157 37655
rect 1173 37603 1225 37655
rect 1241 37644 1293 37655
rect 1241 37610 1273 37644
rect 1273 37610 1293 37644
rect 1241 37603 1293 37610
rect 2097 37603 2149 37655
rect 2165 37644 2217 37655
rect 2165 37610 2183 37644
rect 2183 37610 2217 37644
rect 2165 37603 2217 37610
rect 2233 37603 2285 37655
rect 2301 37603 2353 37655
rect 2369 37644 2421 37655
rect 2437 37644 2489 37655
rect 2369 37610 2419 37644
rect 2419 37610 2421 37644
rect 2437 37610 2453 37644
rect 2453 37610 2489 37644
rect 2369 37603 2421 37610
rect 2437 37603 2489 37610
rect 2505 37603 2557 37655
rect 2573 37603 2625 37655
rect 2641 37644 2693 37655
rect 2641 37610 2655 37644
rect 2655 37610 2689 37644
rect 2689 37610 2693 37644
rect 2641 37603 2693 37610
rect 697 37539 749 37591
rect 765 37570 817 37591
rect 765 37539 767 37570
rect 767 37539 801 37570
rect 801 37539 817 37570
rect 833 37539 885 37591
rect 901 37539 953 37591
rect 969 37570 1021 37591
rect 969 37539 1003 37570
rect 1003 37539 1021 37570
rect 1037 37539 1089 37591
rect 1105 37539 1157 37591
rect 1173 37539 1225 37591
rect 1241 37570 1293 37591
rect 1241 37539 1273 37570
rect 1273 37539 1293 37570
rect 2097 37539 2149 37591
rect 2165 37570 2217 37591
rect 2165 37539 2183 37570
rect 2183 37539 2217 37570
rect 2233 37539 2285 37591
rect 2301 37539 2353 37591
rect 2369 37570 2421 37591
rect 2437 37570 2489 37591
rect 2369 37539 2419 37570
rect 2419 37539 2421 37570
rect 2437 37539 2453 37570
rect 2453 37539 2489 37570
rect 2505 37539 2557 37591
rect 2573 37539 2625 37591
rect 2641 37570 2693 37591
rect 2641 37539 2655 37570
rect 2655 37539 2689 37570
rect 2689 37539 2693 37570
rect 697 37475 749 37527
rect 765 37496 817 37527
rect 765 37475 767 37496
rect 767 37475 801 37496
rect 801 37475 817 37496
rect 833 37475 885 37527
rect 901 37475 953 37527
rect 969 37496 1021 37527
rect 969 37475 1003 37496
rect 1003 37475 1021 37496
rect 1037 37475 1089 37527
rect 1105 37475 1157 37527
rect 1173 37475 1225 37527
rect 1241 37496 1293 37527
rect 1241 37475 1273 37496
rect 1273 37475 1293 37496
rect 2097 37475 2149 37527
rect 2165 37496 2217 37527
rect 2165 37475 2183 37496
rect 2183 37475 2217 37496
rect 2233 37475 2285 37527
rect 2301 37475 2353 37527
rect 2369 37496 2421 37527
rect 2437 37496 2489 37527
rect 2369 37475 2419 37496
rect 2419 37475 2421 37496
rect 2437 37475 2453 37496
rect 2453 37475 2489 37496
rect 2505 37475 2557 37527
rect 2573 37475 2625 37527
rect 2641 37496 2693 37527
rect 2641 37475 2655 37496
rect 2655 37475 2689 37496
rect 2689 37475 2693 37496
rect 1501 36924 1553 36933
rect 1569 36924 1621 36933
rect 1636 36924 1688 36933
rect 1703 36924 1755 36933
rect 1770 36924 1822 36933
rect 1837 36924 1889 36933
rect 1501 36890 1525 36924
rect 1525 36890 1553 36924
rect 1569 36890 1600 36924
rect 1600 36890 1621 36924
rect 1636 36890 1674 36924
rect 1674 36890 1688 36924
rect 1703 36890 1708 36924
rect 1708 36890 1748 36924
rect 1748 36890 1755 36924
rect 1770 36890 1782 36924
rect 1782 36890 1822 36924
rect 1837 36890 1856 36924
rect 1856 36890 1889 36924
rect 1501 36881 1553 36890
rect 1569 36881 1621 36890
rect 1636 36881 1688 36890
rect 1703 36881 1755 36890
rect 1770 36881 1822 36890
rect 1837 36881 1889 36890
rect 697 36317 749 36369
rect 765 36350 767 36369
rect 767 36350 801 36369
rect 801 36350 817 36369
rect 765 36317 817 36350
rect 833 36317 885 36369
rect 901 36317 953 36369
rect 969 36350 1003 36369
rect 1003 36350 1021 36369
rect 969 36317 1021 36350
rect 1037 36317 1089 36369
rect 1105 36317 1157 36369
rect 1173 36317 1225 36369
rect 1241 36350 1273 36369
rect 1273 36350 1293 36369
rect 1241 36317 1293 36350
rect 2097 36317 2149 36369
rect 2165 36350 2183 36369
rect 2183 36350 2217 36369
rect 2165 36317 2217 36350
rect 2233 36317 2285 36369
rect 2301 36317 2353 36369
rect 2369 36350 2419 36369
rect 2419 36350 2421 36369
rect 2437 36350 2453 36369
rect 2453 36350 2489 36369
rect 2369 36317 2421 36350
rect 2437 36317 2489 36350
rect 2505 36317 2557 36369
rect 2573 36317 2625 36369
rect 2641 36350 2655 36369
rect 2655 36350 2689 36369
rect 2689 36350 2693 36369
rect 2641 36317 2693 36350
rect 697 36253 749 36305
rect 765 36277 767 36305
rect 767 36277 801 36305
rect 801 36277 817 36305
rect 765 36253 817 36277
rect 833 36253 885 36305
rect 901 36253 953 36305
rect 969 36277 1003 36305
rect 1003 36277 1021 36305
rect 969 36253 1021 36277
rect 1037 36253 1089 36305
rect 1105 36253 1157 36305
rect 1173 36253 1225 36305
rect 1241 36277 1273 36305
rect 1273 36277 1293 36305
rect 1241 36253 1293 36277
rect 2097 36253 2149 36305
rect 2165 36277 2183 36305
rect 2183 36277 2217 36305
rect 2165 36253 2217 36277
rect 2233 36253 2285 36305
rect 2301 36253 2353 36305
rect 2369 36277 2419 36305
rect 2419 36277 2421 36305
rect 2437 36277 2453 36305
rect 2453 36277 2489 36305
rect 2369 36253 2421 36277
rect 2437 36253 2489 36277
rect 2505 36253 2557 36305
rect 2573 36253 2625 36305
rect 2641 36277 2655 36305
rect 2655 36277 2689 36305
rect 2689 36277 2693 36305
rect 2641 36253 2693 36277
rect 697 36189 749 36241
rect 765 36238 817 36241
rect 765 36204 767 36238
rect 767 36204 801 36238
rect 801 36204 817 36238
rect 765 36189 817 36204
rect 833 36189 885 36241
rect 901 36189 953 36241
rect 969 36238 1021 36241
rect 969 36204 1003 36238
rect 1003 36204 1021 36238
rect 969 36189 1021 36204
rect 1037 36189 1089 36241
rect 1105 36189 1157 36241
rect 1173 36189 1225 36241
rect 1241 36238 1293 36241
rect 1241 36204 1273 36238
rect 1273 36204 1293 36238
rect 1241 36189 1293 36204
rect 2097 36189 2149 36241
rect 2165 36238 2217 36241
rect 2165 36204 2183 36238
rect 2183 36204 2217 36238
rect 2165 36189 2217 36204
rect 2233 36189 2285 36241
rect 2301 36189 2353 36241
rect 2369 36238 2421 36241
rect 2437 36238 2489 36241
rect 2369 36204 2419 36238
rect 2419 36204 2421 36238
rect 2437 36204 2453 36238
rect 2453 36204 2489 36238
rect 2369 36189 2421 36204
rect 2437 36189 2489 36204
rect 2505 36189 2557 36241
rect 2573 36189 2625 36241
rect 2641 36238 2693 36241
rect 2641 36204 2655 36238
rect 2655 36204 2689 36238
rect 2689 36204 2693 36238
rect 2641 36189 2693 36204
rect 697 36125 749 36177
rect 765 36165 817 36177
rect 765 36131 767 36165
rect 767 36131 801 36165
rect 801 36131 817 36165
rect 765 36125 817 36131
rect 833 36125 885 36177
rect 901 36125 953 36177
rect 969 36165 1021 36177
rect 969 36131 1003 36165
rect 1003 36131 1021 36165
rect 969 36125 1021 36131
rect 1037 36125 1089 36177
rect 1105 36125 1157 36177
rect 1173 36125 1225 36177
rect 1241 36165 1293 36177
rect 1241 36131 1273 36165
rect 1273 36131 1293 36165
rect 1241 36125 1293 36131
rect 2097 36125 2149 36177
rect 2165 36165 2217 36177
rect 2165 36131 2183 36165
rect 2183 36131 2217 36165
rect 2165 36125 2217 36131
rect 2233 36125 2285 36177
rect 2301 36125 2353 36177
rect 2369 36165 2421 36177
rect 2437 36165 2489 36177
rect 2369 36131 2419 36165
rect 2419 36131 2421 36165
rect 2437 36131 2453 36165
rect 2453 36131 2489 36165
rect 2369 36125 2421 36131
rect 2437 36125 2489 36131
rect 2505 36125 2557 36177
rect 2573 36125 2625 36177
rect 2641 36165 2693 36177
rect 2641 36131 2655 36165
rect 2655 36131 2689 36165
rect 2689 36131 2693 36165
rect 2641 36125 2693 36131
rect 697 36061 749 36113
rect 765 36092 817 36113
rect 765 36061 767 36092
rect 767 36061 801 36092
rect 801 36061 817 36092
rect 833 36061 885 36113
rect 901 36061 953 36113
rect 969 36092 1021 36113
rect 969 36061 1003 36092
rect 1003 36061 1021 36092
rect 1037 36061 1089 36113
rect 1105 36061 1157 36113
rect 1173 36061 1225 36113
rect 1241 36092 1293 36113
rect 1241 36061 1273 36092
rect 1273 36061 1293 36092
rect 2097 36061 2149 36113
rect 2165 36092 2217 36113
rect 2165 36061 2183 36092
rect 2183 36061 2217 36092
rect 2233 36061 2285 36113
rect 2301 36061 2353 36113
rect 2369 36092 2421 36113
rect 2437 36092 2489 36113
rect 2369 36061 2419 36092
rect 2419 36061 2421 36092
rect 2437 36061 2453 36092
rect 2453 36061 2489 36092
rect 2505 36061 2557 36113
rect 2573 36061 2625 36113
rect 2641 36092 2693 36113
rect 2641 36061 2655 36092
rect 2655 36061 2689 36092
rect 2689 36061 2693 36092
rect 697 35997 749 36049
rect 765 36019 817 36049
rect 765 35997 767 36019
rect 767 35997 801 36019
rect 801 35997 817 36019
rect 833 35997 885 36049
rect 901 35997 953 36049
rect 969 36019 1021 36049
rect 969 35997 1003 36019
rect 1003 35997 1021 36019
rect 1037 35997 1089 36049
rect 1105 35997 1157 36049
rect 1173 35997 1225 36049
rect 1241 36019 1293 36049
rect 1241 35997 1273 36019
rect 1273 35997 1293 36019
rect 2097 35997 2149 36049
rect 2165 36019 2217 36049
rect 2165 35997 2183 36019
rect 2183 35997 2217 36019
rect 2233 35997 2285 36049
rect 2301 35997 2353 36049
rect 2369 36019 2421 36049
rect 2437 36019 2489 36049
rect 2369 35997 2419 36019
rect 2419 35997 2421 36019
rect 2437 35997 2453 36019
rect 2453 35997 2489 36019
rect 2505 35997 2557 36049
rect 2573 35997 2625 36049
rect 2641 36019 2693 36049
rect 2641 35997 2655 36019
rect 2655 35997 2689 36019
rect 2689 35997 2693 36019
rect 697 35933 749 35985
rect 765 35946 817 35985
rect 765 35933 767 35946
rect 767 35933 801 35946
rect 801 35933 817 35946
rect 833 35933 885 35985
rect 901 35933 953 35985
rect 969 35946 1021 35985
rect 969 35933 1003 35946
rect 1003 35933 1021 35946
rect 1037 35933 1089 35985
rect 1105 35933 1157 35985
rect 1173 35933 1225 35985
rect 1241 35946 1293 35985
rect 1241 35933 1273 35946
rect 1273 35933 1293 35946
rect 697 35869 749 35921
rect 765 35912 767 35921
rect 767 35912 801 35921
rect 801 35912 817 35921
rect 765 35872 817 35912
rect 765 35869 767 35872
rect 767 35869 801 35872
rect 801 35869 817 35872
rect 833 35869 885 35921
rect 901 35869 953 35921
rect 969 35912 1003 35921
rect 1003 35912 1021 35921
rect 969 35872 1021 35912
rect 969 35869 1003 35872
rect 1003 35869 1021 35872
rect 1037 35869 1089 35921
rect 1105 35869 1157 35921
rect 1173 35869 1225 35921
rect 1241 35912 1273 35921
rect 1273 35912 1293 35921
rect 2097 35933 2149 35985
rect 2165 35946 2217 35985
rect 2165 35933 2183 35946
rect 2183 35933 2217 35946
rect 2233 35933 2285 35985
rect 2301 35933 2353 35985
rect 2369 35946 2421 35985
rect 2437 35946 2489 35985
rect 2369 35933 2419 35946
rect 2419 35933 2421 35946
rect 2437 35933 2453 35946
rect 2453 35933 2489 35946
rect 2505 35933 2557 35985
rect 2573 35933 2625 35985
rect 2641 35946 2693 35985
rect 2641 35933 2655 35946
rect 2655 35933 2689 35946
rect 2689 35933 2693 35946
rect 1241 35872 1293 35912
rect 1241 35869 1273 35872
rect 1273 35869 1293 35872
rect 697 35805 749 35857
rect 765 35838 767 35857
rect 767 35838 801 35857
rect 801 35838 817 35857
rect 765 35805 817 35838
rect 833 35805 885 35857
rect 901 35805 953 35857
rect 969 35838 1003 35857
rect 1003 35838 1021 35857
rect 969 35805 1021 35838
rect 1037 35805 1089 35857
rect 1105 35805 1157 35857
rect 1173 35805 1225 35857
rect 1241 35838 1273 35857
rect 1273 35838 1293 35857
rect 2097 35869 2149 35921
rect 2165 35912 2183 35921
rect 2183 35912 2217 35921
rect 2165 35872 2217 35912
rect 2165 35869 2183 35872
rect 2183 35869 2217 35872
rect 2233 35869 2285 35921
rect 2301 35869 2353 35921
rect 2369 35912 2419 35921
rect 2419 35912 2421 35921
rect 2437 35912 2453 35921
rect 2453 35912 2489 35921
rect 2369 35872 2421 35912
rect 2437 35872 2489 35912
rect 2369 35869 2419 35872
rect 2419 35869 2421 35872
rect 2437 35869 2453 35872
rect 2453 35869 2489 35872
rect 2505 35869 2557 35921
rect 2573 35869 2625 35921
rect 2641 35912 2655 35921
rect 2655 35912 2689 35921
rect 2689 35912 2693 35921
rect 2641 35872 2693 35912
rect 2641 35869 2655 35872
rect 2655 35869 2689 35872
rect 2689 35869 2693 35872
rect 1241 35805 1293 35838
rect 2097 35805 2149 35857
rect 2165 35838 2183 35857
rect 2183 35838 2217 35857
rect 2165 35805 2217 35838
rect 2233 35805 2285 35857
rect 2301 35805 2353 35857
rect 2369 35838 2419 35857
rect 2419 35838 2421 35857
rect 2437 35838 2453 35857
rect 2453 35838 2489 35857
rect 2369 35805 2421 35838
rect 2437 35805 2489 35838
rect 2505 35805 2557 35857
rect 2573 35805 2625 35857
rect 2641 35838 2655 35857
rect 2655 35838 2689 35857
rect 2689 35838 2693 35857
rect 2641 35805 2693 35838
rect 697 35741 749 35793
rect 765 35764 767 35793
rect 767 35764 801 35793
rect 801 35764 817 35793
rect 765 35741 817 35764
rect 833 35741 885 35793
rect 901 35741 953 35793
rect 969 35764 1003 35793
rect 1003 35764 1021 35793
rect 969 35741 1021 35764
rect 1037 35741 1089 35793
rect 1105 35741 1157 35793
rect 1173 35741 1225 35793
rect 1241 35764 1273 35793
rect 1273 35764 1293 35793
rect 1241 35741 1293 35764
rect 2097 35741 2149 35793
rect 2165 35764 2183 35793
rect 2183 35764 2217 35793
rect 2165 35741 2217 35764
rect 2233 35741 2285 35793
rect 2301 35741 2353 35793
rect 2369 35764 2419 35793
rect 2419 35764 2421 35793
rect 2437 35764 2453 35793
rect 2453 35764 2489 35793
rect 2369 35741 2421 35764
rect 2437 35741 2489 35764
rect 2505 35741 2557 35793
rect 2573 35741 2625 35793
rect 2641 35764 2655 35793
rect 2655 35764 2689 35793
rect 2689 35764 2693 35793
rect 2641 35741 2693 35764
rect 697 35677 749 35729
rect 765 35724 817 35729
rect 765 35690 767 35724
rect 767 35690 801 35724
rect 801 35690 817 35724
rect 765 35677 817 35690
rect 833 35677 885 35729
rect 901 35677 953 35729
rect 969 35724 1021 35729
rect 969 35690 1003 35724
rect 1003 35690 1021 35724
rect 969 35677 1021 35690
rect 1037 35677 1089 35729
rect 1105 35677 1157 35729
rect 1173 35677 1225 35729
rect 1241 35724 1293 35729
rect 1241 35690 1273 35724
rect 1273 35690 1293 35724
rect 1241 35677 1293 35690
rect 2097 35677 2149 35729
rect 2165 35724 2217 35729
rect 2165 35690 2183 35724
rect 2183 35690 2217 35724
rect 2165 35677 2217 35690
rect 2233 35677 2285 35729
rect 2301 35677 2353 35729
rect 2369 35724 2421 35729
rect 2437 35724 2489 35729
rect 2369 35690 2419 35724
rect 2419 35690 2421 35724
rect 2437 35690 2453 35724
rect 2453 35690 2489 35724
rect 2369 35677 2421 35690
rect 2437 35677 2489 35690
rect 2505 35677 2557 35729
rect 2573 35677 2625 35729
rect 2641 35724 2693 35729
rect 2641 35690 2655 35724
rect 2655 35690 2689 35724
rect 2689 35690 2693 35724
rect 2641 35677 2693 35690
rect 697 35613 749 35665
rect 765 35650 817 35665
rect 765 35616 767 35650
rect 767 35616 801 35650
rect 801 35616 817 35650
rect 765 35613 817 35616
rect 833 35613 885 35665
rect 901 35613 953 35665
rect 969 35650 1021 35665
rect 969 35616 1003 35650
rect 1003 35616 1021 35650
rect 969 35613 1021 35616
rect 1037 35613 1089 35665
rect 1105 35613 1157 35665
rect 1173 35613 1225 35665
rect 1241 35650 1293 35665
rect 1241 35616 1273 35650
rect 1273 35616 1293 35650
rect 1241 35613 1293 35616
rect 2097 35613 2149 35665
rect 2165 35650 2217 35665
rect 2165 35616 2183 35650
rect 2183 35616 2217 35650
rect 2165 35613 2217 35616
rect 2233 35613 2285 35665
rect 2301 35613 2353 35665
rect 2369 35650 2421 35665
rect 2437 35650 2489 35665
rect 2369 35616 2419 35650
rect 2419 35616 2421 35650
rect 2437 35616 2453 35650
rect 2453 35616 2489 35650
rect 2369 35613 2421 35616
rect 2437 35613 2489 35616
rect 2505 35613 2557 35665
rect 2573 35613 2625 35665
rect 2641 35650 2693 35665
rect 2641 35616 2655 35650
rect 2655 35616 2689 35650
rect 2689 35616 2693 35650
rect 2641 35613 2693 35616
rect 697 35549 749 35601
rect 765 35576 817 35601
rect 765 35549 767 35576
rect 767 35549 801 35576
rect 801 35549 817 35576
rect 833 35549 885 35601
rect 901 35549 953 35601
rect 969 35576 1021 35601
rect 969 35549 1003 35576
rect 1003 35549 1021 35576
rect 1037 35549 1089 35601
rect 1105 35549 1157 35601
rect 1173 35549 1225 35601
rect 1241 35576 1293 35601
rect 1241 35549 1273 35576
rect 1273 35549 1293 35576
rect 2097 35549 2149 35601
rect 2165 35576 2217 35601
rect 2165 35549 2183 35576
rect 2183 35549 2217 35576
rect 2233 35549 2285 35601
rect 2301 35549 2353 35601
rect 2369 35576 2421 35601
rect 2437 35576 2489 35601
rect 2369 35549 2419 35576
rect 2419 35549 2421 35576
rect 2437 35549 2453 35576
rect 2453 35549 2489 35576
rect 2505 35549 2557 35601
rect 2573 35549 2625 35601
rect 2641 35576 2693 35601
rect 2641 35549 2655 35576
rect 2655 35549 2689 35576
rect 2689 35549 2693 35576
rect 697 35485 749 35537
rect 765 35502 817 35537
rect 765 35485 767 35502
rect 767 35485 801 35502
rect 801 35485 817 35502
rect 833 35485 885 35537
rect 901 35485 953 35537
rect 969 35502 1021 35537
rect 969 35485 1003 35502
rect 1003 35485 1021 35502
rect 1037 35485 1089 35537
rect 1105 35485 1157 35537
rect 1173 35485 1225 35537
rect 1241 35502 1293 35537
rect 1241 35485 1273 35502
rect 1273 35485 1293 35502
rect 697 35421 749 35473
rect 765 35468 767 35473
rect 767 35468 801 35473
rect 801 35468 817 35473
rect 765 35428 817 35468
rect 765 35421 767 35428
rect 767 35421 801 35428
rect 801 35421 817 35428
rect 833 35421 885 35473
rect 901 35421 953 35473
rect 969 35468 1003 35473
rect 1003 35468 1021 35473
rect 969 35428 1021 35468
rect 969 35421 1003 35428
rect 1003 35421 1021 35428
rect 1037 35421 1089 35473
rect 1105 35421 1157 35473
rect 1173 35421 1225 35473
rect 1241 35468 1273 35473
rect 1273 35468 1293 35473
rect 2097 35485 2149 35537
rect 2165 35502 2217 35537
rect 2165 35485 2183 35502
rect 2183 35485 2217 35502
rect 2233 35485 2285 35537
rect 2301 35485 2353 35537
rect 2369 35502 2421 35537
rect 2437 35502 2489 35537
rect 2369 35485 2419 35502
rect 2419 35485 2421 35502
rect 2437 35485 2453 35502
rect 2453 35485 2489 35502
rect 2505 35485 2557 35537
rect 2573 35485 2625 35537
rect 2641 35502 2693 35537
rect 2641 35485 2655 35502
rect 2655 35485 2689 35502
rect 2689 35485 2693 35502
rect 1241 35428 1293 35468
rect 1241 35421 1273 35428
rect 1273 35421 1293 35428
rect 2097 35421 2149 35473
rect 2165 35468 2183 35473
rect 2183 35468 2217 35473
rect 2165 35428 2217 35468
rect 2165 35421 2183 35428
rect 2183 35421 2217 35428
rect 2233 35421 2285 35473
rect 2301 35421 2353 35473
rect 2369 35468 2419 35473
rect 2419 35468 2421 35473
rect 2437 35468 2453 35473
rect 2453 35468 2489 35473
rect 2369 35428 2421 35468
rect 2437 35428 2489 35468
rect 2369 35421 2419 35428
rect 2419 35421 2421 35428
rect 2437 35421 2453 35428
rect 2453 35421 2489 35428
rect 2505 35421 2557 35473
rect 2573 35421 2625 35473
rect 2641 35468 2655 35473
rect 2655 35468 2689 35473
rect 2689 35468 2693 35473
rect 2641 35428 2693 35468
rect 2641 35421 2655 35428
rect 2655 35421 2689 35428
rect 2689 35421 2693 35428
rect 1501 34794 1553 34803
rect 1569 34794 1621 34803
rect 1636 34794 1688 34803
rect 1703 34794 1755 34803
rect 1770 34794 1822 34803
rect 1837 34794 1889 34803
rect 1501 34760 1525 34794
rect 1525 34760 1553 34794
rect 1569 34760 1600 34794
rect 1600 34760 1621 34794
rect 1636 34760 1674 34794
rect 1674 34760 1688 34794
rect 1703 34760 1708 34794
rect 1708 34760 1748 34794
rect 1748 34760 1755 34794
rect 1770 34760 1782 34794
rect 1782 34760 1822 34794
rect 1837 34760 1856 34794
rect 1856 34760 1889 34794
rect 1501 34751 1553 34760
rect 1569 34751 1621 34760
rect 1636 34751 1688 34760
rect 1703 34751 1755 34760
rect 1770 34751 1822 34760
rect 1837 34751 1889 34760
rect 697 34098 749 34150
rect 765 34147 767 34150
rect 767 34147 801 34150
rect 801 34147 817 34150
rect 765 34108 817 34147
rect 765 34098 767 34108
rect 767 34098 801 34108
rect 801 34098 817 34108
rect 833 34098 885 34150
rect 901 34098 953 34150
rect 969 34147 1003 34150
rect 1003 34147 1021 34150
rect 969 34108 1021 34147
rect 969 34098 1003 34108
rect 1003 34098 1021 34108
rect 1037 34098 1089 34150
rect 1105 34098 1157 34150
rect 1173 34098 1225 34150
rect 1241 34147 1273 34150
rect 1273 34147 1293 34150
rect 1241 34108 1293 34147
rect 1241 34098 1273 34108
rect 1273 34098 1293 34108
rect 697 34034 749 34086
rect 765 34074 767 34086
rect 767 34074 801 34086
rect 801 34074 817 34086
rect 765 34035 817 34074
rect 765 34034 767 34035
rect 767 34034 801 34035
rect 801 34034 817 34035
rect 833 34034 885 34086
rect 901 34034 953 34086
rect 969 34074 1003 34086
rect 1003 34074 1021 34086
rect 969 34035 1021 34074
rect 969 34034 1003 34035
rect 1003 34034 1021 34035
rect 1037 34034 1089 34086
rect 1105 34034 1157 34086
rect 1173 34034 1225 34086
rect 1241 34074 1273 34086
rect 1273 34074 1293 34086
rect 2097 34098 2149 34150
rect 2165 34147 2183 34150
rect 2183 34147 2217 34150
rect 2165 34108 2217 34147
rect 2165 34098 2183 34108
rect 2183 34098 2217 34108
rect 2233 34098 2285 34150
rect 2301 34098 2353 34150
rect 2369 34147 2419 34150
rect 2419 34147 2421 34150
rect 2437 34147 2453 34150
rect 2453 34147 2489 34150
rect 2369 34108 2421 34147
rect 2437 34108 2489 34147
rect 2369 34098 2419 34108
rect 2419 34098 2421 34108
rect 2437 34098 2453 34108
rect 2453 34098 2489 34108
rect 2505 34098 2557 34150
rect 2573 34098 2625 34150
rect 2641 34147 2655 34150
rect 2655 34147 2689 34150
rect 2689 34147 2693 34150
rect 2641 34108 2693 34147
rect 2641 34098 2655 34108
rect 2655 34098 2689 34108
rect 2689 34098 2693 34108
rect 1241 34035 1293 34074
rect 1241 34034 1273 34035
rect 1273 34034 1293 34035
rect 697 33970 749 34022
rect 765 34001 767 34022
rect 767 34001 801 34022
rect 801 34001 817 34022
rect 765 33970 817 34001
rect 833 33970 885 34022
rect 901 33970 953 34022
rect 969 34001 1003 34022
rect 1003 34001 1021 34022
rect 969 33970 1021 34001
rect 1037 33970 1089 34022
rect 1105 33970 1157 34022
rect 1173 33970 1225 34022
rect 1241 34001 1273 34022
rect 1273 34001 1293 34022
rect 2097 34034 2149 34086
rect 2165 34074 2183 34086
rect 2183 34074 2217 34086
rect 2165 34035 2217 34074
rect 2165 34034 2183 34035
rect 2183 34034 2217 34035
rect 2233 34034 2285 34086
rect 2301 34034 2353 34086
rect 2369 34074 2419 34086
rect 2419 34074 2421 34086
rect 2437 34074 2453 34086
rect 2453 34074 2489 34086
rect 2369 34035 2421 34074
rect 2437 34035 2489 34074
rect 2369 34034 2419 34035
rect 2419 34034 2421 34035
rect 2437 34034 2453 34035
rect 2453 34034 2489 34035
rect 2505 34034 2557 34086
rect 2573 34034 2625 34086
rect 2641 34074 2655 34086
rect 2655 34074 2689 34086
rect 2689 34074 2693 34086
rect 2641 34035 2693 34074
rect 2641 34034 2655 34035
rect 2655 34034 2689 34035
rect 2689 34034 2693 34035
rect 1241 33970 1293 34001
rect 2097 33970 2149 34022
rect 2165 34001 2183 34022
rect 2183 34001 2217 34022
rect 2165 33970 2217 34001
rect 2233 33970 2285 34022
rect 2301 33970 2353 34022
rect 2369 34001 2419 34022
rect 2419 34001 2421 34022
rect 2437 34001 2453 34022
rect 2453 34001 2489 34022
rect 2369 33970 2421 34001
rect 2437 33970 2489 34001
rect 2505 33970 2557 34022
rect 2573 33970 2625 34022
rect 2641 34001 2655 34022
rect 2655 34001 2689 34022
rect 2689 34001 2693 34022
rect 2641 33970 2693 34001
rect 697 33906 749 33958
rect 765 33928 767 33958
rect 767 33928 801 33958
rect 801 33928 817 33958
rect 765 33906 817 33928
rect 833 33906 885 33958
rect 901 33906 953 33958
rect 969 33928 1003 33958
rect 1003 33928 1021 33958
rect 969 33906 1021 33928
rect 1037 33906 1089 33958
rect 1105 33906 1157 33958
rect 1173 33906 1225 33958
rect 1241 33928 1273 33958
rect 1273 33928 1293 33958
rect 1241 33906 1293 33928
rect 2097 33906 2149 33958
rect 2165 33928 2183 33958
rect 2183 33928 2217 33958
rect 2165 33906 2217 33928
rect 2233 33906 2285 33958
rect 2301 33906 2353 33958
rect 2369 33928 2419 33958
rect 2419 33928 2421 33958
rect 2437 33928 2453 33958
rect 2453 33928 2489 33958
rect 2369 33906 2421 33928
rect 2437 33906 2489 33928
rect 2505 33906 2557 33958
rect 2573 33906 2625 33958
rect 2641 33928 2655 33958
rect 2655 33928 2689 33958
rect 2689 33928 2693 33958
rect 2641 33906 2693 33928
rect 697 33842 749 33894
rect 765 33889 817 33894
rect 765 33855 767 33889
rect 767 33855 801 33889
rect 801 33855 817 33889
rect 765 33842 817 33855
rect 833 33842 885 33894
rect 901 33842 953 33894
rect 969 33889 1021 33894
rect 969 33855 1003 33889
rect 1003 33855 1021 33889
rect 969 33842 1021 33855
rect 1037 33842 1089 33894
rect 1105 33842 1157 33894
rect 1173 33842 1225 33894
rect 1241 33889 1293 33894
rect 1241 33855 1273 33889
rect 1273 33855 1293 33889
rect 1241 33842 1293 33855
rect 2097 33842 2149 33894
rect 2165 33889 2217 33894
rect 2165 33855 2183 33889
rect 2183 33855 2217 33889
rect 2165 33842 2217 33855
rect 2233 33842 2285 33894
rect 2301 33842 2353 33894
rect 2369 33889 2421 33894
rect 2437 33889 2489 33894
rect 2369 33855 2419 33889
rect 2419 33855 2421 33889
rect 2437 33855 2453 33889
rect 2453 33855 2489 33889
rect 2369 33842 2421 33855
rect 2437 33842 2489 33855
rect 2505 33842 2557 33894
rect 2573 33842 2625 33894
rect 2641 33889 2693 33894
rect 2641 33855 2655 33889
rect 2655 33855 2689 33889
rect 2689 33855 2693 33889
rect 2641 33842 2693 33855
rect 697 33778 749 33830
rect 765 33816 817 33830
rect 765 33782 767 33816
rect 767 33782 801 33816
rect 801 33782 817 33816
rect 765 33778 817 33782
rect 833 33778 885 33830
rect 901 33778 953 33830
rect 969 33816 1021 33830
rect 969 33782 1003 33816
rect 1003 33782 1021 33816
rect 969 33778 1021 33782
rect 1037 33778 1089 33830
rect 1105 33778 1157 33830
rect 1173 33778 1225 33830
rect 1241 33816 1293 33830
rect 1241 33782 1273 33816
rect 1273 33782 1293 33816
rect 1241 33778 1293 33782
rect 2097 33778 2149 33830
rect 2165 33816 2217 33830
rect 2165 33782 2183 33816
rect 2183 33782 2217 33816
rect 2165 33778 2217 33782
rect 2233 33778 2285 33830
rect 2301 33778 2353 33830
rect 2369 33816 2421 33830
rect 2437 33816 2489 33830
rect 2369 33782 2419 33816
rect 2419 33782 2421 33816
rect 2437 33782 2453 33816
rect 2453 33782 2489 33816
rect 2369 33778 2421 33782
rect 2437 33778 2489 33782
rect 2505 33778 2557 33830
rect 2573 33778 2625 33830
rect 2641 33816 2693 33830
rect 2641 33782 2655 33816
rect 2655 33782 2689 33816
rect 2689 33782 2693 33816
rect 2641 33778 2693 33782
rect 697 33714 749 33766
rect 765 33742 817 33766
rect 765 33714 767 33742
rect 767 33714 801 33742
rect 801 33714 817 33742
rect 833 33714 885 33766
rect 901 33714 953 33766
rect 969 33742 1021 33766
rect 969 33714 1003 33742
rect 1003 33714 1021 33742
rect 1037 33714 1089 33766
rect 1105 33714 1157 33766
rect 1173 33714 1225 33766
rect 1241 33742 1293 33766
rect 1241 33714 1273 33742
rect 1273 33714 1293 33742
rect 2097 33714 2149 33766
rect 2165 33742 2217 33766
rect 2165 33714 2183 33742
rect 2183 33714 2217 33742
rect 2233 33714 2285 33766
rect 2301 33714 2353 33766
rect 2369 33742 2421 33766
rect 2437 33742 2489 33766
rect 2369 33714 2419 33742
rect 2419 33714 2421 33742
rect 2437 33714 2453 33742
rect 2453 33714 2489 33742
rect 2505 33714 2557 33766
rect 2573 33714 2625 33766
rect 2641 33742 2693 33766
rect 2641 33714 2655 33742
rect 2655 33714 2689 33742
rect 2689 33714 2693 33742
rect 697 33650 749 33702
rect 765 33668 817 33702
rect 765 33650 767 33668
rect 767 33650 801 33668
rect 801 33650 817 33668
rect 833 33650 885 33702
rect 901 33650 953 33702
rect 969 33668 1021 33702
rect 969 33650 1003 33668
rect 1003 33650 1021 33668
rect 1037 33650 1089 33702
rect 1105 33650 1157 33702
rect 1173 33650 1225 33702
rect 1241 33668 1293 33702
rect 1241 33650 1273 33668
rect 1273 33650 1293 33668
rect 697 33586 749 33638
rect 765 33634 767 33638
rect 767 33634 801 33638
rect 801 33634 817 33638
rect 765 33594 817 33634
rect 765 33586 767 33594
rect 767 33586 801 33594
rect 801 33586 817 33594
rect 833 33586 885 33638
rect 901 33586 953 33638
rect 969 33634 1003 33638
rect 1003 33634 1021 33638
rect 969 33594 1021 33634
rect 969 33586 1003 33594
rect 1003 33586 1021 33594
rect 1037 33586 1089 33638
rect 1105 33586 1157 33638
rect 1173 33586 1225 33638
rect 1241 33634 1273 33638
rect 1273 33634 1293 33638
rect 2097 33650 2149 33702
rect 2165 33668 2217 33702
rect 2165 33650 2183 33668
rect 2183 33650 2217 33668
rect 2233 33650 2285 33702
rect 2301 33650 2353 33702
rect 2369 33668 2421 33702
rect 2437 33668 2489 33702
rect 2369 33650 2419 33668
rect 2419 33650 2421 33668
rect 2437 33650 2453 33668
rect 2453 33650 2489 33668
rect 2505 33650 2557 33702
rect 2573 33650 2625 33702
rect 2641 33668 2693 33702
rect 2641 33650 2655 33668
rect 2655 33650 2689 33668
rect 2689 33650 2693 33668
rect 1241 33594 1293 33634
rect 1241 33586 1273 33594
rect 1273 33586 1293 33594
rect 697 33522 749 33574
rect 765 33560 767 33574
rect 767 33560 801 33574
rect 801 33560 817 33574
rect 765 33522 817 33560
rect 833 33522 885 33574
rect 901 33522 953 33574
rect 969 33560 1003 33574
rect 1003 33560 1021 33574
rect 969 33522 1021 33560
rect 1037 33522 1089 33574
rect 1105 33522 1157 33574
rect 1173 33522 1225 33574
rect 1241 33560 1273 33574
rect 1273 33560 1293 33574
rect 2097 33586 2149 33638
rect 2165 33634 2183 33638
rect 2183 33634 2217 33638
rect 2165 33594 2217 33634
rect 2165 33586 2183 33594
rect 2183 33586 2217 33594
rect 2233 33586 2285 33638
rect 2301 33586 2353 33638
rect 2369 33634 2419 33638
rect 2419 33634 2421 33638
rect 2437 33634 2453 33638
rect 2453 33634 2489 33638
rect 2369 33594 2421 33634
rect 2437 33594 2489 33634
rect 2369 33586 2419 33594
rect 2419 33586 2421 33594
rect 2437 33586 2453 33594
rect 2453 33586 2489 33594
rect 2505 33586 2557 33638
rect 2573 33586 2625 33638
rect 2641 33634 2655 33638
rect 2655 33634 2689 33638
rect 2689 33634 2693 33638
rect 2641 33594 2693 33634
rect 2641 33586 2655 33594
rect 2655 33586 2689 33594
rect 2689 33586 2693 33594
rect 1241 33522 1293 33560
rect 2097 33522 2149 33574
rect 2165 33560 2183 33574
rect 2183 33560 2217 33574
rect 2165 33522 2217 33560
rect 2233 33522 2285 33574
rect 2301 33522 2353 33574
rect 2369 33560 2419 33574
rect 2419 33560 2421 33574
rect 2437 33560 2453 33574
rect 2453 33560 2489 33574
rect 2369 33522 2421 33560
rect 2437 33522 2489 33560
rect 2505 33522 2557 33574
rect 2573 33522 2625 33574
rect 2641 33560 2655 33574
rect 2655 33560 2689 33574
rect 2689 33560 2693 33574
rect 2641 33522 2693 33560
rect 697 33458 749 33510
rect 765 33486 767 33510
rect 767 33486 801 33510
rect 801 33486 817 33510
rect 765 33458 817 33486
rect 833 33458 885 33510
rect 901 33458 953 33510
rect 969 33486 1003 33510
rect 1003 33486 1021 33510
rect 969 33458 1021 33486
rect 1037 33458 1089 33510
rect 1105 33458 1157 33510
rect 1173 33458 1225 33510
rect 1241 33486 1273 33510
rect 1273 33486 1293 33510
rect 1241 33458 1293 33486
rect 2097 33458 2149 33510
rect 2165 33486 2183 33510
rect 2183 33486 2217 33510
rect 2165 33458 2217 33486
rect 2233 33458 2285 33510
rect 2301 33458 2353 33510
rect 2369 33486 2419 33510
rect 2419 33486 2421 33510
rect 2437 33486 2453 33510
rect 2453 33486 2489 33510
rect 2369 33458 2421 33486
rect 2437 33458 2489 33486
rect 2505 33458 2557 33510
rect 2573 33458 2625 33510
rect 2641 33486 2655 33510
rect 2655 33486 2689 33510
rect 2689 33486 2693 33510
rect 2641 33458 2693 33486
rect 697 33394 749 33446
rect 765 33412 767 33446
rect 767 33412 801 33446
rect 801 33412 817 33446
rect 765 33394 817 33412
rect 833 33394 885 33446
rect 901 33394 953 33446
rect 969 33412 1003 33446
rect 1003 33412 1021 33446
rect 969 33394 1021 33412
rect 1037 33394 1089 33446
rect 1105 33394 1157 33446
rect 1173 33394 1225 33446
rect 1241 33412 1273 33446
rect 1273 33412 1293 33446
rect 1241 33394 1293 33412
rect 2097 33394 2149 33446
rect 2165 33412 2183 33446
rect 2183 33412 2217 33446
rect 2165 33394 2217 33412
rect 2233 33394 2285 33446
rect 2301 33394 2353 33446
rect 2369 33412 2419 33446
rect 2419 33412 2421 33446
rect 2437 33412 2453 33446
rect 2453 33412 2489 33446
rect 2369 33394 2421 33412
rect 2437 33394 2489 33412
rect 2505 33394 2557 33446
rect 2573 33394 2625 33446
rect 2641 33412 2655 33446
rect 2655 33412 2689 33446
rect 2689 33412 2693 33446
rect 2641 33394 2693 33412
rect 697 33330 749 33382
rect 765 33372 817 33382
rect 765 33338 767 33372
rect 767 33338 801 33372
rect 801 33338 817 33372
rect 765 33330 817 33338
rect 833 33330 885 33382
rect 901 33330 953 33382
rect 969 33372 1021 33382
rect 969 33338 1003 33372
rect 1003 33338 1021 33372
rect 969 33330 1021 33338
rect 1037 33330 1089 33382
rect 1105 33330 1157 33382
rect 1173 33330 1225 33382
rect 1241 33372 1293 33382
rect 1241 33338 1273 33372
rect 1273 33338 1293 33372
rect 1241 33330 1293 33338
rect 2097 33330 2149 33382
rect 2165 33372 2217 33382
rect 2165 33338 2183 33372
rect 2183 33338 2217 33372
rect 2165 33330 2217 33338
rect 2233 33330 2285 33382
rect 2301 33330 2353 33382
rect 2369 33372 2421 33382
rect 2437 33372 2489 33382
rect 2369 33338 2419 33372
rect 2419 33338 2421 33372
rect 2437 33338 2453 33372
rect 2453 33338 2489 33372
rect 2369 33330 2421 33338
rect 2437 33330 2489 33338
rect 2505 33330 2557 33382
rect 2573 33330 2625 33382
rect 2641 33372 2693 33382
rect 2641 33338 2655 33372
rect 2655 33338 2689 33372
rect 2689 33338 2693 33372
rect 2641 33330 2693 33338
rect 697 33266 749 33318
rect 765 33298 817 33318
rect 765 33266 767 33298
rect 767 33266 801 33298
rect 801 33266 817 33298
rect 833 33266 885 33318
rect 901 33266 953 33318
rect 969 33298 1021 33318
rect 969 33266 1003 33298
rect 1003 33266 1021 33298
rect 1037 33266 1089 33318
rect 1105 33266 1157 33318
rect 1173 33266 1225 33318
rect 1241 33298 1293 33318
rect 1241 33266 1273 33298
rect 1273 33266 1293 33298
rect 2097 33266 2149 33318
rect 2165 33298 2217 33318
rect 2165 33266 2183 33298
rect 2183 33266 2217 33298
rect 2233 33266 2285 33318
rect 2301 33266 2353 33318
rect 2369 33298 2421 33318
rect 2437 33298 2489 33318
rect 2369 33266 2419 33298
rect 2419 33266 2421 33298
rect 2437 33266 2453 33298
rect 2453 33266 2489 33298
rect 2505 33266 2557 33318
rect 2573 33266 2625 33318
rect 2641 33298 2693 33318
rect 2641 33266 2655 33298
rect 2655 33266 2689 33298
rect 2689 33266 2693 33298
rect 697 33202 749 33254
rect 765 33224 817 33254
rect 765 33202 767 33224
rect 767 33202 801 33224
rect 801 33202 817 33224
rect 833 33202 885 33254
rect 901 33202 953 33254
rect 969 33224 1021 33254
rect 969 33202 1003 33224
rect 1003 33202 1021 33224
rect 1037 33202 1089 33254
rect 1105 33202 1157 33254
rect 1173 33202 1225 33254
rect 1241 33224 1293 33254
rect 1241 33202 1273 33224
rect 1273 33202 1293 33224
rect 2097 33202 2149 33254
rect 2165 33224 2217 33254
rect 2165 33202 2183 33224
rect 2183 33202 2217 33224
rect 2233 33202 2285 33254
rect 2301 33202 2353 33254
rect 2369 33224 2421 33254
rect 2437 33224 2489 33254
rect 2369 33202 2419 33224
rect 2419 33202 2421 33224
rect 2437 33202 2453 33224
rect 2453 33202 2489 33224
rect 2505 33202 2557 33254
rect 2573 33202 2625 33254
rect 2641 33224 2693 33254
rect 2641 33202 2655 33224
rect 2655 33202 2689 33224
rect 2689 33202 2693 33224
rect 1501 32664 1553 32673
rect 1569 32664 1621 32673
rect 1636 32664 1688 32673
rect 1703 32664 1755 32673
rect 1770 32664 1822 32673
rect 1837 32664 1889 32673
rect 1501 32630 1525 32664
rect 1525 32630 1553 32664
rect 1569 32630 1600 32664
rect 1600 32630 1621 32664
rect 1636 32630 1674 32664
rect 1674 32630 1688 32664
rect 1703 32630 1708 32664
rect 1708 32630 1748 32664
rect 1748 32630 1755 32664
rect 1770 32630 1782 32664
rect 1782 32630 1822 32664
rect 1837 32630 1856 32664
rect 1856 32630 1889 32664
rect 1501 32621 1553 32630
rect 1569 32621 1621 32630
rect 1636 32621 1688 32630
rect 1703 32621 1755 32630
rect 1770 32621 1822 32630
rect 1837 32621 1889 32630
rect 697 31969 749 32021
rect 765 32003 767 32021
rect 767 32003 801 32021
rect 801 32003 817 32021
rect 765 31969 817 32003
rect 833 31969 885 32021
rect 901 31969 953 32021
rect 969 32003 1003 32021
rect 1003 32003 1021 32021
rect 969 31969 1021 32003
rect 1037 31969 1089 32021
rect 1105 31969 1157 32021
rect 1173 31969 1225 32021
rect 1241 32003 1273 32021
rect 1273 32003 1293 32021
rect 1241 31969 1293 32003
rect 2097 31969 2149 32021
rect 2165 32003 2183 32021
rect 2183 32003 2217 32021
rect 2165 31969 2217 32003
rect 2233 31969 2285 32021
rect 2301 31969 2353 32021
rect 2369 32003 2419 32021
rect 2419 32003 2421 32021
rect 2437 32003 2453 32021
rect 2453 32003 2489 32021
rect 2369 31969 2421 32003
rect 2437 31969 2489 32003
rect 2505 31969 2557 32021
rect 2573 31969 2625 32021
rect 2641 32003 2655 32021
rect 2655 32003 2689 32021
rect 2689 32003 2693 32021
rect 2641 31969 2693 32003
rect 697 31905 749 31957
rect 765 31930 767 31957
rect 767 31930 801 31957
rect 801 31930 817 31957
rect 765 31905 817 31930
rect 833 31905 885 31957
rect 901 31905 953 31957
rect 969 31930 1003 31957
rect 1003 31930 1021 31957
rect 969 31905 1021 31930
rect 1037 31905 1089 31957
rect 1105 31905 1157 31957
rect 1173 31905 1225 31957
rect 1241 31930 1273 31957
rect 1273 31930 1293 31957
rect 1241 31905 1293 31930
rect 2097 31905 2149 31957
rect 2165 31930 2183 31957
rect 2183 31930 2217 31957
rect 2165 31905 2217 31930
rect 2233 31905 2285 31957
rect 2301 31905 2353 31957
rect 2369 31930 2419 31957
rect 2419 31930 2421 31957
rect 2437 31930 2453 31957
rect 2453 31930 2489 31957
rect 2369 31905 2421 31930
rect 2437 31905 2489 31930
rect 2505 31905 2557 31957
rect 2573 31905 2625 31957
rect 2641 31930 2655 31957
rect 2655 31930 2689 31957
rect 2689 31930 2693 31957
rect 2641 31905 2693 31930
rect 697 31841 749 31893
rect 765 31891 817 31893
rect 765 31857 767 31891
rect 767 31857 801 31891
rect 801 31857 817 31891
rect 765 31841 817 31857
rect 833 31841 885 31893
rect 901 31841 953 31893
rect 969 31891 1021 31893
rect 969 31857 1003 31891
rect 1003 31857 1021 31891
rect 969 31841 1021 31857
rect 1037 31841 1089 31893
rect 1105 31841 1157 31893
rect 1173 31841 1225 31893
rect 1241 31891 1293 31893
rect 1241 31857 1273 31891
rect 1273 31857 1293 31891
rect 1241 31841 1293 31857
rect 2097 31841 2149 31893
rect 2165 31891 2217 31893
rect 2165 31857 2183 31891
rect 2183 31857 2217 31891
rect 2165 31841 2217 31857
rect 2233 31841 2285 31893
rect 2301 31841 2353 31893
rect 2369 31891 2421 31893
rect 2437 31891 2489 31893
rect 2369 31857 2419 31891
rect 2419 31857 2421 31891
rect 2437 31857 2453 31891
rect 2453 31857 2489 31891
rect 2369 31841 2421 31857
rect 2437 31841 2489 31857
rect 2505 31841 2557 31893
rect 2573 31841 2625 31893
rect 2641 31891 2693 31893
rect 2641 31857 2655 31891
rect 2655 31857 2689 31891
rect 2689 31857 2693 31891
rect 2641 31841 2693 31857
rect 697 31777 749 31829
rect 765 31818 817 31829
rect 765 31784 767 31818
rect 767 31784 801 31818
rect 801 31784 817 31818
rect 765 31777 817 31784
rect 833 31777 885 31829
rect 901 31777 953 31829
rect 969 31818 1021 31829
rect 969 31784 1003 31818
rect 1003 31784 1021 31818
rect 969 31777 1021 31784
rect 1037 31777 1089 31829
rect 1105 31777 1157 31829
rect 1173 31777 1225 31829
rect 1241 31818 1293 31829
rect 1241 31784 1273 31818
rect 1273 31784 1293 31818
rect 1241 31777 1293 31784
rect 2097 31777 2149 31829
rect 2165 31818 2217 31829
rect 2165 31784 2183 31818
rect 2183 31784 2217 31818
rect 2165 31777 2217 31784
rect 2233 31777 2285 31829
rect 2301 31777 2353 31829
rect 2369 31818 2421 31829
rect 2437 31818 2489 31829
rect 2369 31784 2419 31818
rect 2419 31784 2421 31818
rect 2437 31784 2453 31818
rect 2453 31784 2489 31818
rect 2369 31777 2421 31784
rect 2437 31777 2489 31784
rect 2505 31777 2557 31829
rect 2573 31777 2625 31829
rect 2641 31818 2693 31829
rect 2641 31784 2655 31818
rect 2655 31784 2689 31818
rect 2689 31784 2693 31818
rect 2641 31777 2693 31784
rect 697 31713 749 31765
rect 765 31745 817 31765
rect 765 31713 767 31745
rect 767 31713 801 31745
rect 801 31713 817 31745
rect 833 31713 885 31765
rect 901 31713 953 31765
rect 969 31745 1021 31765
rect 969 31713 1003 31745
rect 1003 31713 1021 31745
rect 1037 31713 1089 31765
rect 1105 31713 1157 31765
rect 1173 31713 1225 31765
rect 1241 31745 1293 31765
rect 1241 31713 1273 31745
rect 1273 31713 1293 31745
rect 2097 31713 2149 31765
rect 2165 31745 2217 31765
rect 2165 31713 2183 31745
rect 2183 31713 2217 31745
rect 2233 31713 2285 31765
rect 2301 31713 2353 31765
rect 2369 31745 2421 31765
rect 2437 31745 2489 31765
rect 2369 31713 2419 31745
rect 2419 31713 2421 31745
rect 2437 31713 2453 31745
rect 2453 31713 2489 31745
rect 2505 31713 2557 31765
rect 2573 31713 2625 31765
rect 2641 31745 2693 31765
rect 2641 31713 2655 31745
rect 2655 31713 2689 31745
rect 2689 31713 2693 31745
rect 697 31649 749 31701
rect 765 31672 817 31701
rect 765 31649 767 31672
rect 767 31649 801 31672
rect 801 31649 817 31672
rect 833 31649 885 31701
rect 901 31649 953 31701
rect 969 31672 1021 31701
rect 969 31649 1003 31672
rect 1003 31649 1021 31672
rect 1037 31649 1089 31701
rect 1105 31649 1157 31701
rect 1173 31649 1225 31701
rect 1241 31672 1293 31701
rect 1241 31649 1273 31672
rect 1273 31649 1293 31672
rect 2097 31649 2149 31701
rect 2165 31672 2217 31701
rect 2165 31649 2183 31672
rect 2183 31649 2217 31672
rect 2233 31649 2285 31701
rect 2301 31649 2353 31701
rect 2369 31672 2421 31701
rect 2437 31672 2489 31701
rect 2369 31649 2419 31672
rect 2419 31649 2421 31672
rect 2437 31649 2453 31672
rect 2453 31649 2489 31672
rect 2505 31649 2557 31701
rect 2573 31649 2625 31701
rect 2641 31672 2693 31701
rect 2641 31649 2655 31672
rect 2655 31649 2689 31672
rect 2689 31649 2693 31672
rect 697 31585 749 31637
rect 765 31598 817 31637
rect 765 31585 767 31598
rect 767 31585 801 31598
rect 801 31585 817 31598
rect 833 31585 885 31637
rect 901 31585 953 31637
rect 969 31598 1021 31637
rect 969 31585 1003 31598
rect 1003 31585 1021 31598
rect 1037 31585 1089 31637
rect 1105 31585 1157 31637
rect 1173 31585 1225 31637
rect 1241 31598 1293 31637
rect 1241 31585 1273 31598
rect 1273 31585 1293 31598
rect 697 31521 749 31573
rect 765 31564 767 31573
rect 767 31564 801 31573
rect 801 31564 817 31573
rect 765 31524 817 31564
rect 765 31521 767 31524
rect 767 31521 801 31524
rect 801 31521 817 31524
rect 833 31521 885 31573
rect 901 31521 953 31573
rect 969 31564 1003 31573
rect 1003 31564 1021 31573
rect 969 31524 1021 31564
rect 969 31521 1003 31524
rect 1003 31521 1021 31524
rect 1037 31521 1089 31573
rect 1105 31521 1157 31573
rect 1173 31521 1225 31573
rect 1241 31564 1273 31573
rect 1273 31564 1293 31573
rect 2097 31585 2149 31637
rect 2165 31598 2217 31637
rect 2165 31585 2183 31598
rect 2183 31585 2217 31598
rect 2233 31585 2285 31637
rect 2301 31585 2353 31637
rect 2369 31598 2421 31637
rect 2437 31598 2489 31637
rect 2369 31585 2419 31598
rect 2419 31585 2421 31598
rect 2437 31585 2453 31598
rect 2453 31585 2489 31598
rect 2505 31585 2557 31637
rect 2573 31585 2625 31637
rect 2641 31598 2693 31637
rect 2641 31585 2655 31598
rect 2655 31585 2689 31598
rect 2689 31585 2693 31598
rect 1241 31524 1293 31564
rect 1241 31521 1273 31524
rect 1273 31521 1293 31524
rect 697 31457 749 31509
rect 765 31490 767 31509
rect 767 31490 801 31509
rect 801 31490 817 31509
rect 765 31457 817 31490
rect 833 31457 885 31509
rect 901 31457 953 31509
rect 969 31490 1003 31509
rect 1003 31490 1021 31509
rect 969 31457 1021 31490
rect 1037 31457 1089 31509
rect 1105 31457 1157 31509
rect 1173 31457 1225 31509
rect 1241 31490 1273 31509
rect 1273 31490 1293 31509
rect 2097 31521 2149 31573
rect 2165 31564 2183 31573
rect 2183 31564 2217 31573
rect 2165 31524 2217 31564
rect 2165 31521 2183 31524
rect 2183 31521 2217 31524
rect 2233 31521 2285 31573
rect 2301 31521 2353 31573
rect 2369 31564 2419 31573
rect 2419 31564 2421 31573
rect 2437 31564 2453 31573
rect 2453 31564 2489 31573
rect 2369 31524 2421 31564
rect 2437 31524 2489 31564
rect 2369 31521 2419 31524
rect 2419 31521 2421 31524
rect 2437 31521 2453 31524
rect 2453 31521 2489 31524
rect 2505 31521 2557 31573
rect 2573 31521 2625 31573
rect 2641 31564 2655 31573
rect 2655 31564 2689 31573
rect 2689 31564 2693 31573
rect 2641 31524 2693 31564
rect 2641 31521 2655 31524
rect 2655 31521 2689 31524
rect 2689 31521 2693 31524
rect 1241 31457 1293 31490
rect 2097 31457 2149 31509
rect 2165 31490 2183 31509
rect 2183 31490 2217 31509
rect 2165 31457 2217 31490
rect 2233 31457 2285 31509
rect 2301 31457 2353 31509
rect 2369 31490 2419 31509
rect 2419 31490 2421 31509
rect 2437 31490 2453 31509
rect 2453 31490 2489 31509
rect 2369 31457 2421 31490
rect 2437 31457 2489 31490
rect 2505 31457 2557 31509
rect 2573 31457 2625 31509
rect 2641 31490 2655 31509
rect 2655 31490 2689 31509
rect 2689 31490 2693 31509
rect 2641 31457 2693 31490
rect 697 31393 749 31445
rect 765 31416 767 31445
rect 767 31416 801 31445
rect 801 31416 817 31445
rect 765 31393 817 31416
rect 833 31393 885 31445
rect 901 31393 953 31445
rect 969 31416 1003 31445
rect 1003 31416 1021 31445
rect 969 31393 1021 31416
rect 1037 31393 1089 31445
rect 1105 31393 1157 31445
rect 1173 31393 1225 31445
rect 1241 31416 1273 31445
rect 1273 31416 1293 31445
rect 1241 31393 1293 31416
rect 2097 31393 2149 31445
rect 2165 31416 2183 31445
rect 2183 31416 2217 31445
rect 2165 31393 2217 31416
rect 2233 31393 2285 31445
rect 2301 31393 2353 31445
rect 2369 31416 2419 31445
rect 2419 31416 2421 31445
rect 2437 31416 2453 31445
rect 2453 31416 2489 31445
rect 2369 31393 2421 31416
rect 2437 31393 2489 31416
rect 2505 31393 2557 31445
rect 2573 31393 2625 31445
rect 2641 31416 2655 31445
rect 2655 31416 2689 31445
rect 2689 31416 2693 31445
rect 2641 31393 2693 31416
rect 697 31329 749 31381
rect 765 31376 817 31381
rect 765 31342 767 31376
rect 767 31342 801 31376
rect 801 31342 817 31376
rect 765 31329 817 31342
rect 833 31329 885 31381
rect 901 31329 953 31381
rect 969 31376 1021 31381
rect 969 31342 1003 31376
rect 1003 31342 1021 31376
rect 969 31329 1021 31342
rect 1037 31329 1089 31381
rect 1105 31329 1157 31381
rect 1173 31329 1225 31381
rect 1241 31376 1293 31381
rect 1241 31342 1273 31376
rect 1273 31342 1293 31376
rect 1241 31329 1293 31342
rect 2097 31329 2149 31381
rect 2165 31376 2217 31381
rect 2165 31342 2183 31376
rect 2183 31342 2217 31376
rect 2165 31329 2217 31342
rect 2233 31329 2285 31381
rect 2301 31329 2353 31381
rect 2369 31376 2421 31381
rect 2437 31376 2489 31381
rect 2369 31342 2419 31376
rect 2419 31342 2421 31376
rect 2437 31342 2453 31376
rect 2453 31342 2489 31376
rect 2369 31329 2421 31342
rect 2437 31329 2489 31342
rect 2505 31329 2557 31381
rect 2573 31329 2625 31381
rect 2641 31376 2693 31381
rect 2641 31342 2655 31376
rect 2655 31342 2689 31376
rect 2689 31342 2693 31376
rect 2641 31329 2693 31342
rect 697 31265 749 31317
rect 765 31302 817 31317
rect 765 31268 767 31302
rect 767 31268 801 31302
rect 801 31268 817 31302
rect 765 31265 817 31268
rect 833 31265 885 31317
rect 901 31265 953 31317
rect 969 31302 1021 31317
rect 969 31268 1003 31302
rect 1003 31268 1021 31302
rect 969 31265 1021 31268
rect 1037 31265 1089 31317
rect 1105 31265 1157 31317
rect 1173 31265 1225 31317
rect 1241 31302 1293 31317
rect 1241 31268 1273 31302
rect 1273 31268 1293 31302
rect 1241 31265 1293 31268
rect 2097 31265 2149 31317
rect 2165 31302 2217 31317
rect 2165 31268 2183 31302
rect 2183 31268 2217 31302
rect 2165 31265 2217 31268
rect 2233 31265 2285 31317
rect 2301 31265 2353 31317
rect 2369 31302 2421 31317
rect 2437 31302 2489 31317
rect 2369 31268 2419 31302
rect 2419 31268 2421 31302
rect 2437 31268 2453 31302
rect 2453 31268 2489 31302
rect 2369 31265 2421 31268
rect 2437 31265 2489 31268
rect 2505 31265 2557 31317
rect 2573 31265 2625 31317
rect 2641 31302 2693 31317
rect 2641 31268 2655 31302
rect 2655 31268 2689 31302
rect 2689 31268 2693 31302
rect 2641 31265 2693 31268
rect 697 31201 749 31253
rect 765 31228 817 31253
rect 765 31201 767 31228
rect 767 31201 801 31228
rect 801 31201 817 31228
rect 833 31201 885 31253
rect 901 31201 953 31253
rect 969 31228 1021 31253
rect 969 31201 1003 31228
rect 1003 31201 1021 31228
rect 1037 31201 1089 31253
rect 1105 31201 1157 31253
rect 1173 31201 1225 31253
rect 1241 31228 1293 31253
rect 1241 31201 1273 31228
rect 1273 31201 1293 31228
rect 2097 31201 2149 31253
rect 2165 31228 2217 31253
rect 2165 31201 2183 31228
rect 2183 31201 2217 31228
rect 2233 31201 2285 31253
rect 2301 31201 2353 31253
rect 2369 31228 2421 31253
rect 2437 31228 2489 31253
rect 2369 31201 2419 31228
rect 2419 31201 2421 31228
rect 2437 31201 2453 31228
rect 2453 31201 2489 31228
rect 2505 31201 2557 31253
rect 2573 31201 2625 31253
rect 2641 31228 2693 31253
rect 2641 31201 2655 31228
rect 2655 31201 2689 31228
rect 2689 31201 2693 31228
rect 697 31137 749 31189
rect 765 31154 817 31189
rect 765 31137 767 31154
rect 767 31137 801 31154
rect 801 31137 817 31154
rect 833 31137 885 31189
rect 901 31137 953 31189
rect 969 31154 1021 31189
rect 969 31137 1003 31154
rect 1003 31137 1021 31154
rect 1037 31137 1089 31189
rect 1105 31137 1157 31189
rect 1173 31137 1225 31189
rect 1241 31154 1293 31189
rect 1241 31137 1273 31154
rect 1273 31137 1293 31154
rect 697 31073 749 31125
rect 765 31120 767 31125
rect 767 31120 801 31125
rect 801 31120 817 31125
rect 765 31080 817 31120
rect 765 31073 767 31080
rect 767 31073 801 31080
rect 801 31073 817 31080
rect 833 31073 885 31125
rect 901 31073 953 31125
rect 969 31120 1003 31125
rect 1003 31120 1021 31125
rect 969 31080 1021 31120
rect 969 31073 1003 31080
rect 1003 31073 1021 31080
rect 1037 31073 1089 31125
rect 1105 31073 1157 31125
rect 1173 31073 1225 31125
rect 1241 31120 1273 31125
rect 1273 31120 1293 31125
rect 2097 31137 2149 31189
rect 2165 31154 2217 31189
rect 2165 31137 2183 31154
rect 2183 31137 2217 31154
rect 2233 31137 2285 31189
rect 2301 31137 2353 31189
rect 2369 31154 2421 31189
rect 2437 31154 2489 31189
rect 2369 31137 2419 31154
rect 2419 31137 2421 31154
rect 2437 31137 2453 31154
rect 2453 31137 2489 31154
rect 2505 31137 2557 31189
rect 2573 31137 2625 31189
rect 2641 31154 2693 31189
rect 2641 31137 2655 31154
rect 2655 31137 2689 31154
rect 2689 31137 2693 31154
rect 1241 31080 1293 31120
rect 1241 31073 1273 31080
rect 1273 31073 1293 31080
rect 2097 31073 2149 31125
rect 2165 31120 2183 31125
rect 2183 31120 2217 31125
rect 2165 31080 2217 31120
rect 2165 31073 2183 31080
rect 2183 31073 2217 31080
rect 2233 31073 2285 31125
rect 2301 31073 2353 31125
rect 2369 31120 2419 31125
rect 2419 31120 2421 31125
rect 2437 31120 2453 31125
rect 2453 31120 2489 31125
rect 2369 31080 2421 31120
rect 2437 31080 2489 31120
rect 2369 31073 2419 31080
rect 2419 31073 2421 31080
rect 2437 31073 2453 31080
rect 2453 31073 2489 31080
rect 2505 31073 2557 31125
rect 2573 31073 2625 31125
rect 2641 31120 2655 31125
rect 2655 31120 2689 31125
rect 2689 31120 2693 31125
rect 2641 31080 2693 31120
rect 2641 31073 2655 31080
rect 2655 31073 2689 31080
rect 2689 31073 2693 31080
rect 1501 30534 1553 30543
rect 1569 30534 1621 30543
rect 1636 30534 1688 30543
rect 1703 30534 1755 30543
rect 1770 30534 1822 30543
rect 1837 30534 1889 30543
rect 1501 30500 1525 30534
rect 1525 30500 1553 30534
rect 1569 30500 1600 30534
rect 1600 30500 1621 30534
rect 1636 30500 1674 30534
rect 1674 30500 1688 30534
rect 1703 30500 1708 30534
rect 1708 30500 1748 30534
rect 1748 30500 1755 30534
rect 1770 30500 1782 30534
rect 1782 30500 1822 30534
rect 1837 30500 1856 30534
rect 1856 30500 1889 30534
rect 1501 30491 1553 30500
rect 1569 30491 1621 30500
rect 1636 30491 1688 30500
rect 1703 30491 1755 30500
rect 1770 30491 1822 30500
rect 1837 30491 1889 30500
rect 697 29820 749 29872
rect 765 29848 817 29872
rect 765 29820 767 29848
rect 767 29820 801 29848
rect 801 29820 817 29848
rect 833 29820 885 29872
rect 901 29820 953 29872
rect 969 29848 1021 29872
rect 969 29820 1003 29848
rect 1003 29820 1021 29848
rect 1037 29820 1089 29872
rect 1105 29820 1157 29872
rect 1173 29820 1225 29872
rect 1241 29848 1293 29872
rect 1241 29820 1273 29848
rect 1273 29820 1293 29848
rect 2097 29820 2149 29872
rect 2165 29848 2217 29872
rect 2165 29820 2183 29848
rect 2183 29820 2217 29848
rect 2233 29820 2285 29872
rect 2301 29820 2353 29872
rect 2369 29848 2421 29872
rect 2437 29848 2489 29872
rect 2369 29820 2419 29848
rect 2419 29820 2421 29848
rect 2437 29820 2453 29848
rect 2453 29820 2489 29848
rect 2505 29820 2557 29872
rect 2573 29820 2625 29872
rect 2641 29848 2693 29872
rect 2641 29820 2655 29848
rect 2655 29820 2689 29848
rect 2689 29820 2693 29848
rect 697 29756 749 29808
rect 765 29775 817 29808
rect 765 29756 767 29775
rect 767 29756 801 29775
rect 801 29756 817 29775
rect 833 29756 885 29808
rect 901 29756 953 29808
rect 969 29775 1021 29808
rect 969 29756 1003 29775
rect 1003 29756 1021 29775
rect 1037 29756 1089 29808
rect 1105 29756 1157 29808
rect 1173 29756 1225 29808
rect 1241 29775 1293 29808
rect 1241 29756 1273 29775
rect 1273 29756 1293 29775
rect 697 29692 749 29744
rect 765 29741 767 29744
rect 767 29741 801 29744
rect 801 29741 817 29744
rect 765 29702 817 29741
rect 765 29692 767 29702
rect 767 29692 801 29702
rect 801 29692 817 29702
rect 833 29692 885 29744
rect 901 29692 953 29744
rect 969 29741 1003 29744
rect 1003 29741 1021 29744
rect 969 29702 1021 29741
rect 969 29692 1003 29702
rect 1003 29692 1021 29702
rect 1037 29692 1089 29744
rect 1105 29692 1157 29744
rect 1173 29692 1225 29744
rect 1241 29741 1273 29744
rect 1273 29741 1293 29744
rect 2097 29756 2149 29808
rect 2165 29775 2217 29808
rect 2165 29756 2183 29775
rect 2183 29756 2217 29775
rect 2233 29756 2285 29808
rect 2301 29756 2353 29808
rect 2369 29775 2421 29808
rect 2437 29775 2489 29808
rect 2369 29756 2419 29775
rect 2419 29756 2421 29775
rect 2437 29756 2453 29775
rect 2453 29756 2489 29775
rect 2505 29756 2557 29808
rect 2573 29756 2625 29808
rect 2641 29775 2693 29808
rect 2641 29756 2655 29775
rect 2655 29756 2689 29775
rect 2689 29756 2693 29775
rect 1241 29702 1293 29741
rect 1241 29692 1273 29702
rect 1273 29692 1293 29702
rect 697 29628 749 29680
rect 765 29668 767 29680
rect 767 29668 801 29680
rect 801 29668 817 29680
rect 765 29629 817 29668
rect 765 29628 767 29629
rect 767 29628 801 29629
rect 801 29628 817 29629
rect 833 29628 885 29680
rect 901 29628 953 29680
rect 969 29668 1003 29680
rect 1003 29668 1021 29680
rect 969 29629 1021 29668
rect 969 29628 1003 29629
rect 1003 29628 1021 29629
rect 1037 29628 1089 29680
rect 1105 29628 1157 29680
rect 1173 29628 1225 29680
rect 1241 29668 1273 29680
rect 1273 29668 1293 29680
rect 2097 29692 2149 29744
rect 2165 29741 2183 29744
rect 2183 29741 2217 29744
rect 2165 29702 2217 29741
rect 2165 29692 2183 29702
rect 2183 29692 2217 29702
rect 2233 29692 2285 29744
rect 2301 29692 2353 29744
rect 2369 29741 2419 29744
rect 2419 29741 2421 29744
rect 2437 29741 2453 29744
rect 2453 29741 2489 29744
rect 2369 29702 2421 29741
rect 2437 29702 2489 29741
rect 2369 29692 2419 29702
rect 2419 29692 2421 29702
rect 2437 29692 2453 29702
rect 2453 29692 2489 29702
rect 2505 29692 2557 29744
rect 2573 29692 2625 29744
rect 2641 29741 2655 29744
rect 2655 29741 2689 29744
rect 2689 29741 2693 29744
rect 2641 29702 2693 29741
rect 2641 29692 2655 29702
rect 2655 29692 2689 29702
rect 2689 29692 2693 29702
rect 1241 29629 1293 29668
rect 1241 29628 1273 29629
rect 1273 29628 1293 29629
rect 697 29564 749 29616
rect 765 29595 767 29616
rect 767 29595 801 29616
rect 801 29595 817 29616
rect 765 29564 817 29595
rect 833 29564 885 29616
rect 901 29564 953 29616
rect 969 29595 1003 29616
rect 1003 29595 1021 29616
rect 969 29564 1021 29595
rect 1037 29564 1089 29616
rect 1105 29564 1157 29616
rect 1173 29564 1225 29616
rect 1241 29595 1273 29616
rect 1273 29595 1293 29616
rect 2097 29628 2149 29680
rect 2165 29668 2183 29680
rect 2183 29668 2217 29680
rect 2165 29629 2217 29668
rect 2165 29628 2183 29629
rect 2183 29628 2217 29629
rect 2233 29628 2285 29680
rect 2301 29628 2353 29680
rect 2369 29668 2419 29680
rect 2419 29668 2421 29680
rect 2437 29668 2453 29680
rect 2453 29668 2489 29680
rect 2369 29629 2421 29668
rect 2437 29629 2489 29668
rect 2369 29628 2419 29629
rect 2419 29628 2421 29629
rect 2437 29628 2453 29629
rect 2453 29628 2489 29629
rect 2505 29628 2557 29680
rect 2573 29628 2625 29680
rect 2641 29668 2655 29680
rect 2655 29668 2689 29680
rect 2689 29668 2693 29680
rect 2641 29629 2693 29668
rect 2641 29628 2655 29629
rect 2655 29628 2689 29629
rect 2689 29628 2693 29629
rect 1241 29564 1293 29595
rect 2097 29564 2149 29616
rect 2165 29595 2183 29616
rect 2183 29595 2217 29616
rect 2165 29564 2217 29595
rect 2233 29564 2285 29616
rect 2301 29564 2353 29616
rect 2369 29595 2419 29616
rect 2419 29595 2421 29616
rect 2437 29595 2453 29616
rect 2453 29595 2489 29616
rect 2369 29564 2421 29595
rect 2437 29564 2489 29595
rect 2505 29564 2557 29616
rect 2573 29564 2625 29616
rect 2641 29595 2655 29616
rect 2655 29595 2689 29616
rect 2689 29595 2693 29616
rect 2641 29564 2693 29595
rect 697 29500 749 29552
rect 765 29522 767 29552
rect 767 29522 801 29552
rect 801 29522 817 29552
rect 765 29500 817 29522
rect 833 29500 885 29552
rect 901 29500 953 29552
rect 969 29522 1003 29552
rect 1003 29522 1021 29552
rect 969 29500 1021 29522
rect 1037 29500 1089 29552
rect 1105 29500 1157 29552
rect 1173 29500 1225 29552
rect 1241 29522 1273 29552
rect 1273 29522 1293 29552
rect 1241 29500 1293 29522
rect 2097 29500 2149 29552
rect 2165 29522 2183 29552
rect 2183 29522 2217 29552
rect 2165 29500 2217 29522
rect 2233 29500 2285 29552
rect 2301 29500 2353 29552
rect 2369 29522 2419 29552
rect 2419 29522 2421 29552
rect 2437 29522 2453 29552
rect 2453 29522 2489 29552
rect 2369 29500 2421 29522
rect 2437 29500 2489 29522
rect 2505 29500 2557 29552
rect 2573 29500 2625 29552
rect 2641 29522 2655 29552
rect 2655 29522 2689 29552
rect 2689 29522 2693 29552
rect 2641 29500 2693 29522
rect 697 29436 749 29488
rect 765 29482 817 29488
rect 765 29448 767 29482
rect 767 29448 801 29482
rect 801 29448 817 29482
rect 765 29436 817 29448
rect 833 29436 885 29488
rect 901 29436 953 29488
rect 969 29482 1021 29488
rect 969 29448 1003 29482
rect 1003 29448 1021 29482
rect 969 29436 1021 29448
rect 1037 29436 1089 29488
rect 1105 29436 1157 29488
rect 1173 29436 1225 29488
rect 1241 29482 1293 29488
rect 1241 29448 1273 29482
rect 1273 29448 1293 29482
rect 1241 29436 1293 29448
rect 2097 29436 2149 29488
rect 2165 29482 2217 29488
rect 2165 29448 2183 29482
rect 2183 29448 2217 29482
rect 2165 29436 2217 29448
rect 2233 29436 2285 29488
rect 2301 29436 2353 29488
rect 2369 29482 2421 29488
rect 2437 29482 2489 29488
rect 2369 29448 2419 29482
rect 2419 29448 2421 29482
rect 2437 29448 2453 29482
rect 2453 29448 2489 29482
rect 2369 29436 2421 29448
rect 2437 29436 2489 29448
rect 2505 29436 2557 29488
rect 2573 29436 2625 29488
rect 2641 29482 2693 29488
rect 2641 29448 2655 29482
rect 2655 29448 2689 29482
rect 2689 29448 2693 29482
rect 2641 29436 2693 29448
rect 697 29372 749 29424
rect 765 29408 817 29424
rect 765 29374 767 29408
rect 767 29374 801 29408
rect 801 29374 817 29408
rect 765 29372 817 29374
rect 833 29372 885 29424
rect 901 29372 953 29424
rect 969 29408 1021 29424
rect 969 29374 1003 29408
rect 1003 29374 1021 29408
rect 969 29372 1021 29374
rect 1037 29372 1089 29424
rect 1105 29372 1157 29424
rect 1173 29372 1225 29424
rect 1241 29408 1293 29424
rect 1241 29374 1273 29408
rect 1273 29374 1293 29408
rect 1241 29372 1293 29374
rect 2097 29372 2149 29424
rect 2165 29408 2217 29424
rect 2165 29374 2183 29408
rect 2183 29374 2217 29408
rect 2165 29372 2217 29374
rect 2233 29372 2285 29424
rect 2301 29372 2353 29424
rect 2369 29408 2421 29424
rect 2437 29408 2489 29424
rect 2369 29374 2419 29408
rect 2419 29374 2421 29408
rect 2437 29374 2453 29408
rect 2453 29374 2489 29408
rect 2369 29372 2421 29374
rect 2437 29372 2489 29374
rect 2505 29372 2557 29424
rect 2573 29372 2625 29424
rect 2641 29408 2693 29424
rect 2641 29374 2655 29408
rect 2655 29374 2689 29408
rect 2689 29374 2693 29408
rect 2641 29372 2693 29374
rect 697 29308 749 29360
rect 765 29334 817 29360
rect 765 29308 767 29334
rect 767 29308 801 29334
rect 801 29308 817 29334
rect 833 29308 885 29360
rect 901 29308 953 29360
rect 969 29334 1021 29360
rect 969 29308 1003 29334
rect 1003 29308 1021 29334
rect 1037 29308 1089 29360
rect 1105 29308 1157 29360
rect 1173 29308 1225 29360
rect 1241 29334 1293 29360
rect 1241 29308 1273 29334
rect 1273 29308 1293 29334
rect 2097 29308 2149 29360
rect 2165 29334 2217 29360
rect 2165 29308 2183 29334
rect 2183 29308 2217 29334
rect 2233 29308 2285 29360
rect 2301 29308 2353 29360
rect 2369 29334 2421 29360
rect 2437 29334 2489 29360
rect 2369 29308 2419 29334
rect 2419 29308 2421 29334
rect 2437 29308 2453 29334
rect 2453 29308 2489 29334
rect 2505 29308 2557 29360
rect 2573 29308 2625 29360
rect 2641 29334 2693 29360
rect 2641 29308 2655 29334
rect 2655 29308 2689 29334
rect 2689 29308 2693 29334
rect 697 29244 749 29296
rect 765 29260 817 29296
rect 765 29244 767 29260
rect 767 29244 801 29260
rect 801 29244 817 29260
rect 833 29244 885 29296
rect 901 29244 953 29296
rect 969 29260 1021 29296
rect 969 29244 1003 29260
rect 1003 29244 1021 29260
rect 1037 29244 1089 29296
rect 1105 29244 1157 29296
rect 1173 29244 1225 29296
rect 1241 29260 1293 29296
rect 1241 29244 1273 29260
rect 1273 29244 1293 29260
rect 697 29180 749 29232
rect 765 29226 767 29232
rect 767 29226 801 29232
rect 801 29226 817 29232
rect 765 29186 817 29226
rect 765 29180 767 29186
rect 767 29180 801 29186
rect 801 29180 817 29186
rect 833 29180 885 29232
rect 901 29180 953 29232
rect 969 29226 1003 29232
rect 1003 29226 1021 29232
rect 969 29186 1021 29226
rect 969 29180 1003 29186
rect 1003 29180 1021 29186
rect 1037 29180 1089 29232
rect 1105 29180 1157 29232
rect 1173 29180 1225 29232
rect 1241 29226 1273 29232
rect 1273 29226 1293 29232
rect 2097 29244 2149 29296
rect 2165 29260 2217 29296
rect 2165 29244 2183 29260
rect 2183 29244 2217 29260
rect 2233 29244 2285 29296
rect 2301 29244 2353 29296
rect 2369 29260 2421 29296
rect 2437 29260 2489 29296
rect 2369 29244 2419 29260
rect 2419 29244 2421 29260
rect 2437 29244 2453 29260
rect 2453 29244 2489 29260
rect 2505 29244 2557 29296
rect 2573 29244 2625 29296
rect 2641 29260 2693 29296
rect 2641 29244 2655 29260
rect 2655 29244 2689 29260
rect 2689 29244 2693 29260
rect 1241 29186 1293 29226
rect 1241 29180 1273 29186
rect 1273 29180 1293 29186
rect 697 29116 749 29168
rect 765 29152 767 29168
rect 767 29152 801 29168
rect 801 29152 817 29168
rect 765 29116 817 29152
rect 833 29116 885 29168
rect 901 29116 953 29168
rect 969 29152 1003 29168
rect 1003 29152 1021 29168
rect 969 29116 1021 29152
rect 1037 29116 1089 29168
rect 1105 29116 1157 29168
rect 1173 29116 1225 29168
rect 1241 29152 1273 29168
rect 1273 29152 1293 29168
rect 2097 29180 2149 29232
rect 2165 29226 2183 29232
rect 2183 29226 2217 29232
rect 2165 29186 2217 29226
rect 2165 29180 2183 29186
rect 2183 29180 2217 29186
rect 2233 29180 2285 29232
rect 2301 29180 2353 29232
rect 2369 29226 2419 29232
rect 2419 29226 2421 29232
rect 2437 29226 2453 29232
rect 2453 29226 2489 29232
rect 2369 29186 2421 29226
rect 2437 29186 2489 29226
rect 2369 29180 2419 29186
rect 2419 29180 2421 29186
rect 2437 29180 2453 29186
rect 2453 29180 2489 29186
rect 2505 29180 2557 29232
rect 2573 29180 2625 29232
rect 2641 29226 2655 29232
rect 2655 29226 2689 29232
rect 2689 29226 2693 29232
rect 2641 29186 2693 29226
rect 2641 29180 2655 29186
rect 2655 29180 2689 29186
rect 2689 29180 2693 29186
rect 1241 29116 1293 29152
rect 2097 29116 2149 29168
rect 2165 29152 2183 29168
rect 2183 29152 2217 29168
rect 2165 29116 2217 29152
rect 2233 29116 2285 29168
rect 2301 29116 2353 29168
rect 2369 29152 2419 29168
rect 2419 29152 2421 29168
rect 2437 29152 2453 29168
rect 2453 29152 2489 29168
rect 2369 29116 2421 29152
rect 2437 29116 2489 29152
rect 2505 29116 2557 29168
rect 2573 29116 2625 29168
rect 2641 29152 2655 29168
rect 2655 29152 2689 29168
rect 2689 29152 2693 29168
rect 2641 29116 2693 29152
rect 697 29052 749 29104
rect 765 29078 767 29104
rect 767 29078 801 29104
rect 801 29078 817 29104
rect 765 29052 817 29078
rect 833 29052 885 29104
rect 901 29052 953 29104
rect 969 29078 1003 29104
rect 1003 29078 1021 29104
rect 969 29052 1021 29078
rect 1037 29052 1089 29104
rect 1105 29052 1157 29104
rect 1173 29052 1225 29104
rect 1241 29078 1273 29104
rect 1273 29078 1293 29104
rect 1241 29052 1293 29078
rect 2097 29052 2149 29104
rect 2165 29078 2183 29104
rect 2183 29078 2217 29104
rect 2165 29052 2217 29078
rect 2233 29052 2285 29104
rect 2301 29052 2353 29104
rect 2369 29078 2419 29104
rect 2419 29078 2421 29104
rect 2437 29078 2453 29104
rect 2453 29078 2489 29104
rect 2369 29052 2421 29078
rect 2437 29052 2489 29078
rect 2505 29052 2557 29104
rect 2573 29052 2625 29104
rect 2641 29078 2655 29104
rect 2655 29078 2689 29104
rect 2689 29078 2693 29104
rect 2641 29052 2693 29078
rect 697 28988 749 29040
rect 765 29038 817 29040
rect 765 29004 767 29038
rect 767 29004 801 29038
rect 801 29004 817 29038
rect 765 28988 817 29004
rect 833 28988 885 29040
rect 901 28988 953 29040
rect 969 29038 1021 29040
rect 969 29004 1003 29038
rect 1003 29004 1021 29038
rect 969 28988 1021 29004
rect 1037 28988 1089 29040
rect 1105 28988 1157 29040
rect 1173 28988 1225 29040
rect 1241 29038 1293 29040
rect 1241 29004 1273 29038
rect 1273 29004 1293 29038
rect 1241 28988 1293 29004
rect 2097 28988 2149 29040
rect 2165 29038 2217 29040
rect 2165 29004 2183 29038
rect 2183 29004 2217 29038
rect 2165 28988 2217 29004
rect 2233 28988 2285 29040
rect 2301 28988 2353 29040
rect 2369 29038 2421 29040
rect 2437 29038 2489 29040
rect 2369 29004 2419 29038
rect 2419 29004 2421 29038
rect 2437 29004 2453 29038
rect 2453 29004 2489 29038
rect 2369 28988 2421 29004
rect 2437 28988 2489 29004
rect 2505 28988 2557 29040
rect 2573 28988 2625 29040
rect 2641 29038 2693 29040
rect 2641 29004 2655 29038
rect 2655 29004 2689 29038
rect 2689 29004 2693 29038
rect 2641 28988 2693 29004
rect 697 28924 749 28976
rect 765 28964 817 28976
rect 765 28930 767 28964
rect 767 28930 801 28964
rect 801 28930 817 28964
rect 765 28924 817 28930
rect 833 28924 885 28976
rect 901 28924 953 28976
rect 969 28964 1021 28976
rect 969 28930 1003 28964
rect 1003 28930 1021 28964
rect 969 28924 1021 28930
rect 1037 28924 1089 28976
rect 1105 28924 1157 28976
rect 1173 28924 1225 28976
rect 1241 28964 1293 28976
rect 1241 28930 1273 28964
rect 1273 28930 1293 28964
rect 1241 28924 1293 28930
rect 2097 28924 2149 28976
rect 2165 28964 2217 28976
rect 2165 28930 2183 28964
rect 2183 28930 2217 28964
rect 2165 28924 2217 28930
rect 2233 28924 2285 28976
rect 2301 28924 2353 28976
rect 2369 28964 2421 28976
rect 2437 28964 2489 28976
rect 2369 28930 2419 28964
rect 2419 28930 2421 28964
rect 2437 28930 2453 28964
rect 2453 28930 2489 28964
rect 2369 28924 2421 28930
rect 2437 28924 2489 28930
rect 2505 28924 2557 28976
rect 2573 28924 2625 28976
rect 2641 28964 2693 28976
rect 2641 28930 2655 28964
rect 2655 28930 2689 28964
rect 2689 28930 2693 28964
rect 2641 28924 2693 28930
rect 1501 28404 1553 28413
rect 1569 28404 1621 28413
rect 1636 28404 1688 28413
rect 1703 28404 1755 28413
rect 1770 28404 1822 28413
rect 1837 28404 1889 28413
rect 1501 28370 1525 28404
rect 1525 28370 1553 28404
rect 1569 28370 1600 28404
rect 1600 28370 1621 28404
rect 1636 28370 1674 28404
rect 1674 28370 1688 28404
rect 1703 28370 1708 28404
rect 1708 28370 1748 28404
rect 1748 28370 1755 28404
rect 1770 28370 1782 28404
rect 1782 28370 1822 28404
rect 1837 28370 1856 28404
rect 1856 28370 1889 28404
rect 1501 28361 1553 28370
rect 1569 28361 1621 28370
rect 1636 28361 1688 28370
rect 1703 28361 1755 28370
rect 1770 28361 1822 28370
rect 1837 28361 1889 28370
rect 697 27813 749 27865
rect 765 27850 817 27865
rect 765 27816 767 27850
rect 767 27816 801 27850
rect 801 27816 817 27850
rect 765 27813 817 27816
rect 833 27813 885 27865
rect 901 27813 953 27865
rect 969 27850 1021 27865
rect 969 27816 1003 27850
rect 1003 27816 1021 27850
rect 969 27813 1021 27816
rect 1037 27813 1089 27865
rect 1105 27813 1157 27865
rect 1173 27813 1225 27865
rect 1241 27850 1293 27865
rect 1241 27816 1273 27850
rect 1273 27816 1293 27850
rect 1241 27813 1293 27816
rect 2097 27813 2149 27865
rect 2165 27850 2217 27865
rect 2165 27816 2183 27850
rect 2183 27816 2217 27850
rect 2165 27813 2217 27816
rect 2233 27813 2285 27865
rect 2301 27813 2353 27865
rect 2369 27850 2421 27865
rect 2437 27850 2489 27865
rect 2369 27816 2419 27850
rect 2419 27816 2421 27850
rect 2437 27816 2453 27850
rect 2453 27816 2489 27850
rect 2369 27813 2421 27816
rect 2437 27813 2489 27816
rect 2505 27813 2557 27865
rect 2573 27813 2625 27865
rect 2641 27850 2693 27865
rect 2641 27816 2655 27850
rect 2655 27816 2689 27850
rect 2689 27816 2693 27850
rect 2641 27813 2693 27816
rect 697 27749 749 27801
rect 765 27777 817 27801
rect 765 27749 767 27777
rect 767 27749 801 27777
rect 801 27749 817 27777
rect 833 27749 885 27801
rect 901 27749 953 27801
rect 969 27777 1021 27801
rect 969 27749 1003 27777
rect 1003 27749 1021 27777
rect 1037 27749 1089 27801
rect 1105 27749 1157 27801
rect 1173 27749 1225 27801
rect 1241 27777 1293 27801
rect 1241 27749 1273 27777
rect 1273 27749 1293 27777
rect 2097 27749 2149 27801
rect 2165 27777 2217 27801
rect 2165 27749 2183 27777
rect 2183 27749 2217 27777
rect 2233 27749 2285 27801
rect 2301 27749 2353 27801
rect 2369 27777 2421 27801
rect 2437 27777 2489 27801
rect 2369 27749 2419 27777
rect 2419 27749 2421 27777
rect 2437 27749 2453 27777
rect 2453 27749 2489 27777
rect 2505 27749 2557 27801
rect 2573 27749 2625 27801
rect 2641 27777 2693 27801
rect 2641 27749 2655 27777
rect 2655 27749 2689 27777
rect 2689 27749 2693 27777
rect 697 27685 749 27737
rect 765 27704 817 27737
rect 765 27685 767 27704
rect 767 27685 801 27704
rect 801 27685 817 27704
rect 833 27685 885 27737
rect 901 27685 953 27737
rect 969 27704 1021 27737
rect 969 27685 1003 27704
rect 1003 27685 1021 27704
rect 1037 27685 1089 27737
rect 1105 27685 1157 27737
rect 1173 27685 1225 27737
rect 1241 27704 1293 27737
rect 1241 27685 1273 27704
rect 1273 27685 1293 27704
rect 697 27621 749 27673
rect 765 27670 767 27673
rect 767 27670 801 27673
rect 801 27670 817 27673
rect 765 27631 817 27670
rect 765 27621 767 27631
rect 767 27621 801 27631
rect 801 27621 817 27631
rect 833 27621 885 27673
rect 901 27621 953 27673
rect 969 27670 1003 27673
rect 1003 27670 1021 27673
rect 969 27631 1021 27670
rect 969 27621 1003 27631
rect 1003 27621 1021 27631
rect 1037 27621 1089 27673
rect 1105 27621 1157 27673
rect 1173 27621 1225 27673
rect 1241 27670 1273 27673
rect 1273 27670 1293 27673
rect 2097 27685 2149 27737
rect 2165 27704 2217 27737
rect 2165 27685 2183 27704
rect 2183 27685 2217 27704
rect 2233 27685 2285 27737
rect 2301 27685 2353 27737
rect 2369 27704 2421 27737
rect 2437 27704 2489 27737
rect 2369 27685 2419 27704
rect 2419 27685 2421 27704
rect 2437 27685 2453 27704
rect 2453 27685 2489 27704
rect 2505 27685 2557 27737
rect 2573 27685 2625 27737
rect 2641 27704 2693 27737
rect 2641 27685 2655 27704
rect 2655 27685 2689 27704
rect 2689 27685 2693 27704
rect 1241 27631 1293 27670
rect 1241 27621 1273 27631
rect 1273 27621 1293 27631
rect 697 27557 749 27609
rect 765 27597 767 27609
rect 767 27597 801 27609
rect 801 27597 817 27609
rect 765 27558 817 27597
rect 765 27557 767 27558
rect 767 27557 801 27558
rect 801 27557 817 27558
rect 833 27557 885 27609
rect 901 27557 953 27609
rect 969 27597 1003 27609
rect 1003 27597 1021 27609
rect 969 27558 1021 27597
rect 969 27557 1003 27558
rect 1003 27557 1021 27558
rect 1037 27557 1089 27609
rect 1105 27557 1157 27609
rect 1173 27557 1225 27609
rect 1241 27597 1273 27609
rect 1273 27597 1293 27609
rect 2097 27621 2149 27673
rect 2165 27670 2183 27673
rect 2183 27670 2217 27673
rect 2165 27631 2217 27670
rect 2165 27621 2183 27631
rect 2183 27621 2217 27631
rect 2233 27621 2285 27673
rect 2301 27621 2353 27673
rect 2369 27670 2419 27673
rect 2419 27670 2421 27673
rect 2437 27670 2453 27673
rect 2453 27670 2489 27673
rect 2369 27631 2421 27670
rect 2437 27631 2489 27670
rect 2369 27621 2419 27631
rect 2419 27621 2421 27631
rect 2437 27621 2453 27631
rect 2453 27621 2489 27631
rect 2505 27621 2557 27673
rect 2573 27621 2625 27673
rect 2641 27670 2655 27673
rect 2655 27670 2689 27673
rect 2689 27670 2693 27673
rect 2641 27631 2693 27670
rect 2641 27621 2655 27631
rect 2655 27621 2689 27631
rect 2689 27621 2693 27631
rect 1241 27558 1293 27597
rect 1241 27557 1273 27558
rect 1273 27557 1293 27558
rect 697 27493 749 27545
rect 765 27524 767 27545
rect 767 27524 801 27545
rect 801 27524 817 27545
rect 765 27493 817 27524
rect 833 27493 885 27545
rect 901 27493 953 27545
rect 969 27524 1003 27545
rect 1003 27524 1021 27545
rect 969 27493 1021 27524
rect 1037 27493 1089 27545
rect 1105 27493 1157 27545
rect 1173 27493 1225 27545
rect 1241 27524 1273 27545
rect 1273 27524 1293 27545
rect 2097 27557 2149 27609
rect 2165 27597 2183 27609
rect 2183 27597 2217 27609
rect 2165 27558 2217 27597
rect 2165 27557 2183 27558
rect 2183 27557 2217 27558
rect 2233 27557 2285 27609
rect 2301 27557 2353 27609
rect 2369 27597 2419 27609
rect 2419 27597 2421 27609
rect 2437 27597 2453 27609
rect 2453 27597 2489 27609
rect 2369 27558 2421 27597
rect 2437 27558 2489 27597
rect 2369 27557 2419 27558
rect 2419 27557 2421 27558
rect 2437 27557 2453 27558
rect 2453 27557 2489 27558
rect 2505 27557 2557 27609
rect 2573 27557 2625 27609
rect 2641 27597 2655 27609
rect 2655 27597 2689 27609
rect 2689 27597 2693 27609
rect 2641 27558 2693 27597
rect 2641 27557 2655 27558
rect 2655 27557 2689 27558
rect 2689 27557 2693 27558
rect 1241 27493 1293 27524
rect 2097 27493 2149 27545
rect 2165 27524 2183 27545
rect 2183 27524 2217 27545
rect 2165 27493 2217 27524
rect 2233 27493 2285 27545
rect 2301 27493 2353 27545
rect 2369 27524 2419 27545
rect 2419 27524 2421 27545
rect 2437 27524 2453 27545
rect 2453 27524 2489 27545
rect 2369 27493 2421 27524
rect 2437 27493 2489 27524
rect 2505 27493 2557 27545
rect 2573 27493 2625 27545
rect 2641 27524 2655 27545
rect 2655 27524 2689 27545
rect 2689 27524 2693 27545
rect 2641 27493 2693 27524
rect 697 27429 749 27481
rect 765 27451 767 27481
rect 767 27451 801 27481
rect 801 27451 817 27481
rect 765 27429 817 27451
rect 833 27429 885 27481
rect 901 27429 953 27481
rect 969 27451 1003 27481
rect 1003 27451 1021 27481
rect 969 27429 1021 27451
rect 1037 27429 1089 27481
rect 1105 27429 1157 27481
rect 1173 27429 1225 27481
rect 1241 27451 1273 27481
rect 1273 27451 1293 27481
rect 1241 27429 1293 27451
rect 2097 27429 2149 27481
rect 2165 27451 2183 27481
rect 2183 27451 2217 27481
rect 2165 27429 2217 27451
rect 2233 27429 2285 27481
rect 2301 27429 2353 27481
rect 2369 27451 2419 27481
rect 2419 27451 2421 27481
rect 2437 27451 2453 27481
rect 2453 27451 2489 27481
rect 2369 27429 2421 27451
rect 2437 27429 2489 27451
rect 2505 27429 2557 27481
rect 2573 27429 2625 27481
rect 2641 27451 2655 27481
rect 2655 27451 2689 27481
rect 2689 27451 2693 27481
rect 2641 27429 2693 27451
rect 697 27365 749 27417
rect 765 27412 817 27417
rect 765 27378 767 27412
rect 767 27378 801 27412
rect 801 27378 817 27412
rect 765 27365 817 27378
rect 833 27365 885 27417
rect 901 27365 953 27417
rect 969 27412 1021 27417
rect 969 27378 1003 27412
rect 1003 27378 1021 27412
rect 969 27365 1021 27378
rect 1037 27365 1089 27417
rect 1105 27365 1157 27417
rect 1173 27365 1225 27417
rect 1241 27412 1293 27417
rect 1241 27378 1273 27412
rect 1273 27378 1293 27412
rect 1241 27365 1293 27378
rect 2097 27365 2149 27417
rect 2165 27412 2217 27417
rect 2165 27378 2183 27412
rect 2183 27378 2217 27412
rect 2165 27365 2217 27378
rect 2233 27365 2285 27417
rect 2301 27365 2353 27417
rect 2369 27412 2421 27417
rect 2437 27412 2489 27417
rect 2369 27378 2419 27412
rect 2419 27378 2421 27412
rect 2437 27378 2453 27412
rect 2453 27378 2489 27412
rect 2369 27365 2421 27378
rect 2437 27365 2489 27378
rect 2505 27365 2557 27417
rect 2573 27365 2625 27417
rect 2641 27412 2693 27417
rect 2641 27378 2655 27412
rect 2655 27378 2689 27412
rect 2689 27378 2693 27412
rect 2641 27365 2693 27378
rect 697 27301 749 27353
rect 765 27338 817 27353
rect 765 27304 767 27338
rect 767 27304 801 27338
rect 801 27304 817 27338
rect 765 27301 817 27304
rect 833 27301 885 27353
rect 901 27301 953 27353
rect 969 27338 1021 27353
rect 969 27304 1003 27338
rect 1003 27304 1021 27338
rect 969 27301 1021 27304
rect 1037 27301 1089 27353
rect 1105 27301 1157 27353
rect 1173 27301 1225 27353
rect 1241 27338 1293 27353
rect 1241 27304 1273 27338
rect 1273 27304 1293 27338
rect 1241 27301 1293 27304
rect 2097 27301 2149 27353
rect 2165 27338 2217 27353
rect 2165 27304 2183 27338
rect 2183 27304 2217 27338
rect 2165 27301 2217 27304
rect 2233 27301 2285 27353
rect 2301 27301 2353 27353
rect 2369 27338 2421 27353
rect 2437 27338 2489 27353
rect 2369 27304 2419 27338
rect 2419 27304 2421 27338
rect 2437 27304 2453 27338
rect 2453 27304 2489 27338
rect 2369 27301 2421 27304
rect 2437 27301 2489 27304
rect 2505 27301 2557 27353
rect 2573 27301 2625 27353
rect 2641 27338 2693 27353
rect 2641 27304 2655 27338
rect 2655 27304 2689 27338
rect 2689 27304 2693 27338
rect 2641 27301 2693 27304
rect 697 27237 749 27289
rect 765 27264 817 27289
rect 765 27237 767 27264
rect 767 27237 801 27264
rect 801 27237 817 27264
rect 833 27237 885 27289
rect 901 27237 953 27289
rect 969 27264 1021 27289
rect 969 27237 1003 27264
rect 1003 27237 1021 27264
rect 1037 27237 1089 27289
rect 1105 27237 1157 27289
rect 1173 27237 1225 27289
rect 1241 27264 1293 27289
rect 1241 27237 1273 27264
rect 1273 27237 1293 27264
rect 2097 27237 2149 27289
rect 2165 27264 2217 27289
rect 2165 27237 2183 27264
rect 2183 27237 2217 27264
rect 2233 27237 2285 27289
rect 2301 27237 2353 27289
rect 2369 27264 2421 27289
rect 2437 27264 2489 27289
rect 2369 27237 2419 27264
rect 2419 27237 2421 27264
rect 2437 27237 2453 27264
rect 2453 27237 2489 27264
rect 2505 27237 2557 27289
rect 2573 27237 2625 27289
rect 2641 27264 2693 27289
rect 2641 27237 2655 27264
rect 2655 27237 2689 27264
rect 2689 27237 2693 27264
rect 697 27173 749 27225
rect 765 27190 817 27225
rect 765 27173 767 27190
rect 767 27173 801 27190
rect 801 27173 817 27190
rect 833 27173 885 27225
rect 901 27173 953 27225
rect 969 27190 1021 27225
rect 969 27173 1003 27190
rect 1003 27173 1021 27190
rect 1037 27173 1089 27225
rect 1105 27173 1157 27225
rect 1173 27173 1225 27225
rect 1241 27190 1293 27225
rect 1241 27173 1273 27190
rect 1273 27173 1293 27190
rect 697 27109 749 27161
rect 765 27156 767 27161
rect 767 27156 801 27161
rect 801 27156 817 27161
rect 765 27116 817 27156
rect 765 27109 767 27116
rect 767 27109 801 27116
rect 801 27109 817 27116
rect 833 27109 885 27161
rect 901 27109 953 27161
rect 969 27156 1003 27161
rect 1003 27156 1021 27161
rect 969 27116 1021 27156
rect 969 27109 1003 27116
rect 1003 27109 1021 27116
rect 1037 27109 1089 27161
rect 1105 27109 1157 27161
rect 1173 27109 1225 27161
rect 1241 27156 1273 27161
rect 1273 27156 1293 27161
rect 2097 27173 2149 27225
rect 2165 27190 2217 27225
rect 2165 27173 2183 27190
rect 2183 27173 2217 27190
rect 2233 27173 2285 27225
rect 2301 27173 2353 27225
rect 2369 27190 2421 27225
rect 2437 27190 2489 27225
rect 2369 27173 2419 27190
rect 2419 27173 2421 27190
rect 2437 27173 2453 27190
rect 2453 27173 2489 27190
rect 2505 27173 2557 27225
rect 2573 27173 2625 27225
rect 2641 27190 2693 27225
rect 2641 27173 2655 27190
rect 2655 27173 2689 27190
rect 2689 27173 2693 27190
rect 1241 27116 1293 27156
rect 1241 27109 1273 27116
rect 1273 27109 1293 27116
rect 697 27045 749 27097
rect 765 27082 767 27097
rect 767 27082 801 27097
rect 801 27082 817 27097
rect 765 27045 817 27082
rect 833 27045 885 27097
rect 901 27045 953 27097
rect 969 27082 1003 27097
rect 1003 27082 1021 27097
rect 969 27045 1021 27082
rect 1037 27045 1089 27097
rect 1105 27045 1157 27097
rect 1173 27045 1225 27097
rect 1241 27082 1273 27097
rect 1273 27082 1293 27097
rect 2097 27109 2149 27161
rect 2165 27156 2183 27161
rect 2183 27156 2217 27161
rect 2165 27116 2217 27156
rect 2165 27109 2183 27116
rect 2183 27109 2217 27116
rect 2233 27109 2285 27161
rect 2301 27109 2353 27161
rect 2369 27156 2419 27161
rect 2419 27156 2421 27161
rect 2437 27156 2453 27161
rect 2453 27156 2489 27161
rect 2369 27116 2421 27156
rect 2437 27116 2489 27156
rect 2369 27109 2419 27116
rect 2419 27109 2421 27116
rect 2437 27109 2453 27116
rect 2453 27109 2489 27116
rect 2505 27109 2557 27161
rect 2573 27109 2625 27161
rect 2641 27156 2655 27161
rect 2655 27156 2689 27161
rect 2689 27156 2693 27161
rect 2641 27116 2693 27156
rect 2641 27109 2655 27116
rect 2655 27109 2689 27116
rect 2689 27109 2693 27116
rect 1241 27045 1293 27082
rect 2097 27045 2149 27097
rect 2165 27082 2183 27097
rect 2183 27082 2217 27097
rect 2165 27045 2217 27082
rect 2233 27045 2285 27097
rect 2301 27045 2353 27097
rect 2369 27082 2419 27097
rect 2419 27082 2421 27097
rect 2437 27082 2453 27097
rect 2453 27082 2489 27097
rect 2369 27045 2421 27082
rect 2437 27045 2489 27082
rect 2505 27045 2557 27097
rect 2573 27045 2625 27097
rect 2641 27082 2655 27097
rect 2655 27082 2689 27097
rect 2689 27082 2693 27097
rect 2641 27045 2693 27082
rect 697 26981 749 27033
rect 765 27008 767 27033
rect 767 27008 801 27033
rect 801 27008 817 27033
rect 765 26981 817 27008
rect 833 26981 885 27033
rect 901 26981 953 27033
rect 969 27008 1003 27033
rect 1003 27008 1021 27033
rect 969 26981 1021 27008
rect 1037 26981 1089 27033
rect 1105 26981 1157 27033
rect 1173 26981 1225 27033
rect 1241 27008 1273 27033
rect 1273 27008 1293 27033
rect 1241 26981 1293 27008
rect 2097 26981 2149 27033
rect 2165 27008 2183 27033
rect 2183 27008 2217 27033
rect 2165 26981 2217 27008
rect 2233 26981 2285 27033
rect 2301 26981 2353 27033
rect 2369 27008 2419 27033
rect 2419 27008 2421 27033
rect 2437 27008 2453 27033
rect 2453 27008 2489 27033
rect 2369 26981 2421 27008
rect 2437 26981 2489 27008
rect 2505 26981 2557 27033
rect 2573 26981 2625 27033
rect 2641 27008 2655 27033
rect 2655 27008 2689 27033
rect 2689 27008 2693 27033
rect 2641 26981 2693 27008
rect 697 26917 749 26969
rect 765 26968 817 26969
rect 765 26934 767 26968
rect 767 26934 801 26968
rect 801 26934 817 26968
rect 765 26917 817 26934
rect 833 26917 885 26969
rect 901 26917 953 26969
rect 969 26968 1021 26969
rect 969 26934 1003 26968
rect 1003 26934 1021 26968
rect 969 26917 1021 26934
rect 1037 26917 1089 26969
rect 1105 26917 1157 26969
rect 1173 26917 1225 26969
rect 1241 26968 1293 26969
rect 1241 26934 1273 26968
rect 1273 26934 1293 26968
rect 1241 26917 1293 26934
rect 2097 26917 2149 26969
rect 2165 26968 2217 26969
rect 2165 26934 2183 26968
rect 2183 26934 2217 26968
rect 2165 26917 2217 26934
rect 2233 26917 2285 26969
rect 2301 26917 2353 26969
rect 2369 26968 2421 26969
rect 2437 26968 2489 26969
rect 2369 26934 2419 26968
rect 2419 26934 2421 26968
rect 2437 26934 2453 26968
rect 2453 26934 2489 26968
rect 2369 26917 2421 26934
rect 2437 26917 2489 26934
rect 2505 26917 2557 26969
rect 2573 26917 2625 26969
rect 2641 26968 2693 26969
rect 2641 26934 2655 26968
rect 2655 26934 2689 26968
rect 2689 26934 2693 26968
rect 2641 26917 2693 26934
rect 1501 26274 1553 26283
rect 1569 26274 1621 26283
rect 1636 26274 1688 26283
rect 1703 26274 1755 26283
rect 1770 26274 1822 26283
rect 1837 26274 1889 26283
rect 1501 26240 1525 26274
rect 1525 26240 1553 26274
rect 1569 26240 1600 26274
rect 1600 26240 1621 26274
rect 1636 26240 1674 26274
rect 1674 26240 1688 26274
rect 1703 26240 1708 26274
rect 1708 26240 1748 26274
rect 1748 26240 1755 26274
rect 1770 26240 1782 26274
rect 1782 26240 1822 26274
rect 1837 26240 1856 26274
rect 1856 26240 1889 26274
rect 1501 26231 1553 26240
rect 1569 26231 1621 26240
rect 1636 26231 1688 26240
rect 1703 26231 1755 26240
rect 1770 26231 1822 26240
rect 1837 26231 1889 26240
rect 697 25627 749 25679
rect 765 25661 817 25679
rect 765 25627 767 25661
rect 767 25627 801 25661
rect 801 25627 817 25661
rect 833 25627 885 25679
rect 901 25627 953 25679
rect 969 25661 1021 25679
rect 969 25627 1003 25661
rect 1003 25627 1021 25661
rect 1037 25627 1089 25679
rect 1105 25627 1157 25679
rect 1173 25627 1225 25679
rect 1241 25661 1293 25679
rect 1241 25627 1273 25661
rect 1273 25627 1293 25661
rect 2097 25627 2149 25679
rect 2165 25661 2217 25679
rect 2165 25627 2183 25661
rect 2183 25627 2217 25661
rect 2233 25627 2285 25679
rect 2301 25627 2353 25679
rect 2369 25661 2421 25679
rect 2437 25661 2489 25679
rect 2369 25627 2419 25661
rect 2419 25627 2421 25661
rect 2437 25627 2453 25661
rect 2453 25627 2489 25661
rect 2505 25627 2557 25679
rect 2573 25627 2625 25679
rect 2641 25661 2693 25679
rect 2641 25627 2655 25661
rect 2655 25627 2689 25661
rect 2689 25627 2693 25661
rect 697 25563 749 25615
rect 765 25588 817 25615
rect 765 25563 767 25588
rect 767 25563 801 25588
rect 801 25563 817 25588
rect 833 25563 885 25615
rect 901 25563 953 25615
rect 969 25588 1021 25615
rect 969 25563 1003 25588
rect 1003 25563 1021 25588
rect 1037 25563 1089 25615
rect 1105 25563 1157 25615
rect 1173 25563 1225 25615
rect 1241 25588 1293 25615
rect 1241 25563 1273 25588
rect 1273 25563 1293 25588
rect 2097 25563 2149 25615
rect 2165 25588 2217 25615
rect 2165 25563 2183 25588
rect 2183 25563 2217 25588
rect 2233 25563 2285 25615
rect 2301 25563 2353 25615
rect 2369 25588 2421 25615
rect 2437 25588 2489 25615
rect 2369 25563 2419 25588
rect 2419 25563 2421 25588
rect 2437 25563 2453 25588
rect 2453 25563 2489 25588
rect 2505 25563 2557 25615
rect 2573 25563 2625 25615
rect 2641 25588 2693 25615
rect 2641 25563 2655 25588
rect 2655 25563 2689 25588
rect 2689 25563 2693 25588
rect 697 25499 749 25551
rect 765 25515 817 25551
rect 765 25499 767 25515
rect 767 25499 801 25515
rect 801 25499 817 25515
rect 833 25499 885 25551
rect 901 25499 953 25551
rect 969 25515 1021 25551
rect 969 25499 1003 25515
rect 1003 25499 1021 25515
rect 1037 25499 1089 25551
rect 1105 25499 1157 25551
rect 1173 25499 1225 25551
rect 1241 25515 1293 25551
rect 1241 25499 1273 25515
rect 1273 25499 1293 25515
rect 697 25435 749 25487
rect 765 25481 767 25487
rect 767 25481 801 25487
rect 801 25481 817 25487
rect 765 25442 817 25481
rect 765 25435 767 25442
rect 767 25435 801 25442
rect 801 25435 817 25442
rect 833 25435 885 25487
rect 901 25435 953 25487
rect 969 25481 1003 25487
rect 1003 25481 1021 25487
rect 969 25442 1021 25481
rect 969 25435 1003 25442
rect 1003 25435 1021 25442
rect 1037 25435 1089 25487
rect 1105 25435 1157 25487
rect 1173 25435 1225 25487
rect 1241 25481 1273 25487
rect 1273 25481 1293 25487
rect 2097 25499 2149 25551
rect 2165 25515 2217 25551
rect 2165 25499 2183 25515
rect 2183 25499 2217 25515
rect 2233 25499 2285 25551
rect 2301 25499 2353 25551
rect 2369 25515 2421 25551
rect 2437 25515 2489 25551
rect 2369 25499 2419 25515
rect 2419 25499 2421 25515
rect 2437 25499 2453 25515
rect 2453 25499 2489 25515
rect 2505 25499 2557 25551
rect 2573 25499 2625 25551
rect 2641 25515 2693 25551
rect 2641 25499 2655 25515
rect 2655 25499 2689 25515
rect 2689 25499 2693 25515
rect 1241 25442 1293 25481
rect 1241 25435 1273 25442
rect 1273 25435 1293 25442
rect 697 25371 749 25423
rect 765 25408 767 25423
rect 767 25408 801 25423
rect 801 25408 817 25423
rect 765 25371 817 25408
rect 833 25371 885 25423
rect 901 25371 953 25423
rect 969 25408 1003 25423
rect 1003 25408 1021 25423
rect 969 25371 1021 25408
rect 1037 25371 1089 25423
rect 1105 25371 1157 25423
rect 1173 25371 1225 25423
rect 1241 25408 1273 25423
rect 1273 25408 1293 25423
rect 2097 25435 2149 25487
rect 2165 25481 2183 25487
rect 2183 25481 2217 25487
rect 2165 25442 2217 25481
rect 2165 25435 2183 25442
rect 2183 25435 2217 25442
rect 2233 25435 2285 25487
rect 2301 25435 2353 25487
rect 2369 25481 2419 25487
rect 2419 25481 2421 25487
rect 2437 25481 2453 25487
rect 2453 25481 2489 25487
rect 2369 25442 2421 25481
rect 2437 25442 2489 25481
rect 2369 25435 2419 25442
rect 2419 25435 2421 25442
rect 2437 25435 2453 25442
rect 2453 25435 2489 25442
rect 2505 25435 2557 25487
rect 2573 25435 2625 25487
rect 2641 25481 2655 25487
rect 2655 25481 2689 25487
rect 2689 25481 2693 25487
rect 2641 25442 2693 25481
rect 2641 25435 2655 25442
rect 2655 25435 2689 25442
rect 2689 25435 2693 25442
rect 1241 25371 1293 25408
rect 2097 25371 2149 25423
rect 2165 25408 2183 25423
rect 2183 25408 2217 25423
rect 2165 25371 2217 25408
rect 2233 25371 2285 25423
rect 2301 25371 2353 25423
rect 2369 25408 2419 25423
rect 2419 25408 2421 25423
rect 2437 25408 2453 25423
rect 2453 25408 2489 25423
rect 2369 25371 2421 25408
rect 2437 25371 2489 25408
rect 2505 25371 2557 25423
rect 2573 25371 2625 25423
rect 2641 25408 2655 25423
rect 2655 25408 2689 25423
rect 2689 25408 2693 25423
rect 2641 25371 2693 25408
rect 697 25307 749 25359
rect 765 25335 767 25359
rect 767 25335 801 25359
rect 801 25335 817 25359
rect 765 25307 817 25335
rect 833 25307 885 25359
rect 901 25307 953 25359
rect 969 25335 1003 25359
rect 1003 25335 1021 25359
rect 969 25307 1021 25335
rect 1037 25307 1089 25359
rect 1105 25307 1157 25359
rect 1173 25307 1225 25359
rect 1241 25335 1273 25359
rect 1273 25335 1293 25359
rect 1241 25307 1293 25335
rect 2097 25307 2149 25359
rect 2165 25335 2183 25359
rect 2183 25335 2217 25359
rect 2165 25307 2217 25335
rect 2233 25307 2285 25359
rect 2301 25307 2353 25359
rect 2369 25335 2419 25359
rect 2419 25335 2421 25359
rect 2437 25335 2453 25359
rect 2453 25335 2489 25359
rect 2369 25307 2421 25335
rect 2437 25307 2489 25335
rect 2505 25307 2557 25359
rect 2573 25307 2625 25359
rect 2641 25335 2655 25359
rect 2655 25335 2689 25359
rect 2689 25335 2693 25359
rect 2641 25307 2693 25335
rect 697 25243 749 25295
rect 765 25262 767 25295
rect 767 25262 801 25295
rect 801 25262 817 25295
rect 765 25243 817 25262
rect 833 25243 885 25295
rect 901 25243 953 25295
rect 969 25262 1003 25295
rect 1003 25262 1021 25295
rect 969 25243 1021 25262
rect 1037 25243 1089 25295
rect 1105 25243 1157 25295
rect 1173 25243 1225 25295
rect 1241 25262 1273 25295
rect 1273 25262 1293 25295
rect 1241 25243 1293 25262
rect 2097 25243 2149 25295
rect 2165 25262 2183 25295
rect 2183 25262 2217 25295
rect 2165 25243 2217 25262
rect 2233 25243 2285 25295
rect 2301 25243 2353 25295
rect 2369 25262 2419 25295
rect 2419 25262 2421 25295
rect 2437 25262 2453 25295
rect 2453 25262 2489 25295
rect 2369 25243 2421 25262
rect 2437 25243 2489 25262
rect 2505 25243 2557 25295
rect 2573 25243 2625 25295
rect 2641 25262 2655 25295
rect 2655 25262 2689 25295
rect 2689 25262 2693 25295
rect 2641 25243 2693 25262
rect 697 25179 749 25231
rect 765 25222 817 25231
rect 765 25188 767 25222
rect 767 25188 801 25222
rect 801 25188 817 25222
rect 765 25179 817 25188
rect 833 25179 885 25231
rect 901 25179 953 25231
rect 969 25222 1021 25231
rect 969 25188 1003 25222
rect 1003 25188 1021 25222
rect 969 25179 1021 25188
rect 1037 25179 1089 25231
rect 1105 25179 1157 25231
rect 1173 25179 1225 25231
rect 1241 25222 1293 25231
rect 1241 25188 1273 25222
rect 1273 25188 1293 25222
rect 1241 25179 1293 25188
rect 2097 25179 2149 25231
rect 2165 25222 2217 25231
rect 2165 25188 2183 25222
rect 2183 25188 2217 25222
rect 2165 25179 2217 25188
rect 2233 25179 2285 25231
rect 2301 25179 2353 25231
rect 2369 25222 2421 25231
rect 2437 25222 2489 25231
rect 2369 25188 2419 25222
rect 2419 25188 2421 25222
rect 2437 25188 2453 25222
rect 2453 25188 2489 25222
rect 2369 25179 2421 25188
rect 2437 25179 2489 25188
rect 2505 25179 2557 25231
rect 2573 25179 2625 25231
rect 2641 25222 2693 25231
rect 2641 25188 2655 25222
rect 2655 25188 2689 25222
rect 2689 25188 2693 25222
rect 2641 25179 2693 25188
rect 697 25115 749 25167
rect 765 25148 817 25167
rect 765 25115 767 25148
rect 767 25115 801 25148
rect 801 25115 817 25148
rect 833 25115 885 25167
rect 901 25115 953 25167
rect 969 25148 1021 25167
rect 969 25115 1003 25148
rect 1003 25115 1021 25148
rect 1037 25115 1089 25167
rect 1105 25115 1157 25167
rect 1173 25115 1225 25167
rect 1241 25148 1293 25167
rect 1241 25115 1273 25148
rect 1273 25115 1293 25148
rect 2097 25115 2149 25167
rect 2165 25148 2217 25167
rect 2165 25115 2183 25148
rect 2183 25115 2217 25148
rect 2233 25115 2285 25167
rect 2301 25115 2353 25167
rect 2369 25148 2421 25167
rect 2437 25148 2489 25167
rect 2369 25115 2419 25148
rect 2419 25115 2421 25148
rect 2437 25115 2453 25148
rect 2453 25115 2489 25148
rect 2505 25115 2557 25167
rect 2573 25115 2625 25167
rect 2641 25148 2693 25167
rect 2641 25115 2655 25148
rect 2655 25115 2689 25148
rect 2689 25115 2693 25148
rect 697 25051 749 25103
rect 765 25074 817 25103
rect 765 25051 767 25074
rect 767 25051 801 25074
rect 801 25051 817 25074
rect 833 25051 885 25103
rect 901 25051 953 25103
rect 969 25074 1021 25103
rect 969 25051 1003 25074
rect 1003 25051 1021 25074
rect 1037 25051 1089 25103
rect 1105 25051 1157 25103
rect 1173 25051 1225 25103
rect 1241 25074 1293 25103
rect 1241 25051 1273 25074
rect 1273 25051 1293 25074
rect 2097 25051 2149 25103
rect 2165 25074 2217 25103
rect 2165 25051 2183 25074
rect 2183 25051 2217 25074
rect 2233 25051 2285 25103
rect 2301 25051 2353 25103
rect 2369 25074 2421 25103
rect 2437 25074 2489 25103
rect 2369 25051 2419 25074
rect 2419 25051 2421 25074
rect 2437 25051 2453 25074
rect 2453 25051 2489 25074
rect 2505 25051 2557 25103
rect 2573 25051 2625 25103
rect 2641 25074 2693 25103
rect 2641 25051 2655 25074
rect 2655 25051 2689 25074
rect 2689 25051 2693 25074
rect 697 24987 749 25039
rect 765 25000 817 25039
rect 765 24987 767 25000
rect 767 24987 801 25000
rect 801 24987 817 25000
rect 833 24987 885 25039
rect 901 24987 953 25039
rect 969 25000 1021 25039
rect 969 24987 1003 25000
rect 1003 24987 1021 25000
rect 1037 24987 1089 25039
rect 1105 24987 1157 25039
rect 1173 24987 1225 25039
rect 1241 25000 1293 25039
rect 1241 24987 1273 25000
rect 1273 24987 1293 25000
rect 697 24923 749 24975
rect 765 24966 767 24975
rect 767 24966 801 24975
rect 801 24966 817 24975
rect 765 24926 817 24966
rect 765 24923 767 24926
rect 767 24923 801 24926
rect 801 24923 817 24926
rect 833 24923 885 24975
rect 901 24923 953 24975
rect 969 24966 1003 24975
rect 1003 24966 1021 24975
rect 969 24926 1021 24966
rect 969 24923 1003 24926
rect 1003 24923 1021 24926
rect 1037 24923 1089 24975
rect 1105 24923 1157 24975
rect 1173 24923 1225 24975
rect 1241 24966 1273 24975
rect 1273 24966 1293 24975
rect 2097 24987 2149 25039
rect 2165 25000 2217 25039
rect 2165 24987 2183 25000
rect 2183 24987 2217 25000
rect 2233 24987 2285 25039
rect 2301 24987 2353 25039
rect 2369 25000 2421 25039
rect 2437 25000 2489 25039
rect 2369 24987 2419 25000
rect 2419 24987 2421 25000
rect 2437 24987 2453 25000
rect 2453 24987 2489 25000
rect 2505 24987 2557 25039
rect 2573 24987 2625 25039
rect 2641 25000 2693 25039
rect 2641 24987 2655 25000
rect 2655 24987 2689 25000
rect 2689 24987 2693 25000
rect 1241 24926 1293 24966
rect 1241 24923 1273 24926
rect 1273 24923 1293 24926
rect 697 24859 749 24911
rect 765 24892 767 24911
rect 767 24892 801 24911
rect 801 24892 817 24911
rect 765 24859 817 24892
rect 833 24859 885 24911
rect 901 24859 953 24911
rect 969 24892 1003 24911
rect 1003 24892 1021 24911
rect 969 24859 1021 24892
rect 1037 24859 1089 24911
rect 1105 24859 1157 24911
rect 1173 24859 1225 24911
rect 1241 24892 1273 24911
rect 1273 24892 1293 24911
rect 2097 24923 2149 24975
rect 2165 24966 2183 24975
rect 2183 24966 2217 24975
rect 2165 24926 2217 24966
rect 2165 24923 2183 24926
rect 2183 24923 2217 24926
rect 2233 24923 2285 24975
rect 2301 24923 2353 24975
rect 2369 24966 2419 24975
rect 2419 24966 2421 24975
rect 2437 24966 2453 24975
rect 2453 24966 2489 24975
rect 2369 24926 2421 24966
rect 2437 24926 2489 24966
rect 2369 24923 2419 24926
rect 2419 24923 2421 24926
rect 2437 24923 2453 24926
rect 2453 24923 2489 24926
rect 2505 24923 2557 24975
rect 2573 24923 2625 24975
rect 2641 24966 2655 24975
rect 2655 24966 2689 24975
rect 2689 24966 2693 24975
rect 2641 24926 2693 24966
rect 2641 24923 2655 24926
rect 2655 24923 2689 24926
rect 2689 24923 2693 24926
rect 1241 24859 1293 24892
rect 2097 24859 2149 24911
rect 2165 24892 2183 24911
rect 2183 24892 2217 24911
rect 2165 24859 2217 24892
rect 2233 24859 2285 24911
rect 2301 24859 2353 24911
rect 2369 24892 2419 24911
rect 2419 24892 2421 24911
rect 2437 24892 2453 24911
rect 2453 24892 2489 24911
rect 2369 24859 2421 24892
rect 2437 24859 2489 24892
rect 2505 24859 2557 24911
rect 2573 24859 2625 24911
rect 2641 24892 2655 24911
rect 2655 24892 2689 24911
rect 2689 24892 2693 24911
rect 2641 24859 2693 24892
rect 697 24795 749 24847
rect 765 24818 767 24847
rect 767 24818 801 24847
rect 801 24818 817 24847
rect 765 24795 817 24818
rect 833 24795 885 24847
rect 901 24795 953 24847
rect 969 24818 1003 24847
rect 1003 24818 1021 24847
rect 969 24795 1021 24818
rect 1037 24795 1089 24847
rect 1105 24795 1157 24847
rect 1173 24795 1225 24847
rect 1241 24818 1273 24847
rect 1273 24818 1293 24847
rect 1241 24795 1293 24818
rect 2097 24795 2149 24847
rect 2165 24818 2183 24847
rect 2183 24818 2217 24847
rect 2165 24795 2217 24818
rect 2233 24795 2285 24847
rect 2301 24795 2353 24847
rect 2369 24818 2419 24847
rect 2419 24818 2421 24847
rect 2437 24818 2453 24847
rect 2453 24818 2489 24847
rect 2369 24795 2421 24818
rect 2437 24795 2489 24818
rect 2505 24795 2557 24847
rect 2573 24795 2625 24847
rect 2641 24818 2655 24847
rect 2655 24818 2689 24847
rect 2689 24818 2693 24847
rect 2641 24795 2693 24818
rect 697 24731 749 24783
rect 765 24778 817 24783
rect 765 24744 767 24778
rect 767 24744 801 24778
rect 801 24744 817 24778
rect 765 24731 817 24744
rect 833 24731 885 24783
rect 901 24731 953 24783
rect 969 24778 1021 24783
rect 969 24744 1003 24778
rect 1003 24744 1021 24778
rect 969 24731 1021 24744
rect 1037 24731 1089 24783
rect 1105 24731 1157 24783
rect 1173 24731 1225 24783
rect 1241 24778 1293 24783
rect 1241 24744 1273 24778
rect 1273 24744 1293 24778
rect 1241 24731 1293 24744
rect 2097 24731 2149 24783
rect 2165 24778 2217 24783
rect 2165 24744 2183 24778
rect 2183 24744 2217 24778
rect 2165 24731 2217 24744
rect 2233 24731 2285 24783
rect 2301 24731 2353 24783
rect 2369 24778 2421 24783
rect 2437 24778 2489 24783
rect 2369 24744 2419 24778
rect 2419 24744 2421 24778
rect 2437 24744 2453 24778
rect 2453 24744 2489 24778
rect 2369 24731 2421 24744
rect 2437 24731 2489 24744
rect 2505 24731 2557 24783
rect 2573 24731 2625 24783
rect 2641 24778 2693 24783
rect 2641 24744 2655 24778
rect 2655 24744 2689 24778
rect 2689 24744 2693 24778
rect 2641 24731 2693 24744
rect 1501 24144 1553 24153
rect 1569 24144 1621 24153
rect 1636 24144 1688 24153
rect 1703 24144 1755 24153
rect 1770 24144 1822 24153
rect 1837 24144 1889 24153
rect 1501 24110 1525 24144
rect 1525 24110 1553 24144
rect 1569 24110 1600 24144
rect 1600 24110 1621 24144
rect 1636 24110 1674 24144
rect 1674 24110 1688 24144
rect 1703 24110 1708 24144
rect 1708 24110 1748 24144
rect 1748 24110 1755 24144
rect 1770 24110 1782 24144
rect 1782 24110 1822 24144
rect 1837 24110 1856 24144
rect 1856 24110 1889 24144
rect 1501 24101 1553 24110
rect 1569 24101 1621 24110
rect 1636 24101 1688 24110
rect 1703 24101 1755 24110
rect 1770 24101 1822 24110
rect 1837 24101 1889 24110
rect 697 23479 749 23531
rect 765 23517 817 23531
rect 765 23483 767 23517
rect 767 23483 801 23517
rect 801 23483 817 23517
rect 765 23479 817 23483
rect 833 23479 885 23531
rect 901 23479 953 23531
rect 969 23517 1021 23531
rect 969 23483 1003 23517
rect 1003 23483 1021 23517
rect 969 23479 1021 23483
rect 1037 23479 1089 23531
rect 1105 23479 1157 23531
rect 1173 23479 1225 23531
rect 1241 23517 1293 23531
rect 1241 23483 1273 23517
rect 1273 23483 1293 23517
rect 1241 23479 1293 23483
rect 2097 23479 2149 23531
rect 2165 23517 2217 23531
rect 2165 23483 2183 23517
rect 2183 23483 2217 23517
rect 2165 23479 2217 23483
rect 2233 23479 2285 23531
rect 2301 23479 2353 23531
rect 2369 23517 2421 23531
rect 2437 23517 2489 23531
rect 2369 23483 2419 23517
rect 2419 23483 2421 23517
rect 2437 23483 2453 23517
rect 2453 23483 2489 23517
rect 2369 23479 2421 23483
rect 2437 23479 2489 23483
rect 2505 23479 2557 23531
rect 2573 23479 2625 23531
rect 2641 23517 2693 23531
rect 2641 23483 2655 23517
rect 2655 23483 2689 23517
rect 2689 23483 2693 23517
rect 2641 23479 2693 23483
rect 697 23415 749 23467
rect 765 23444 817 23467
rect 765 23415 767 23444
rect 767 23415 801 23444
rect 801 23415 817 23444
rect 833 23415 885 23467
rect 901 23415 953 23467
rect 969 23444 1021 23467
rect 969 23415 1003 23444
rect 1003 23415 1021 23444
rect 1037 23415 1089 23467
rect 1105 23415 1157 23467
rect 1173 23415 1225 23467
rect 1241 23444 1293 23467
rect 1241 23415 1273 23444
rect 1273 23415 1293 23444
rect 2097 23415 2149 23467
rect 2165 23444 2217 23467
rect 2165 23415 2183 23444
rect 2183 23415 2217 23444
rect 2233 23415 2285 23467
rect 2301 23415 2353 23467
rect 2369 23444 2421 23467
rect 2437 23444 2489 23467
rect 2369 23415 2419 23444
rect 2419 23415 2421 23444
rect 2437 23415 2453 23444
rect 2453 23415 2489 23444
rect 2505 23415 2557 23467
rect 2573 23415 2625 23467
rect 2641 23444 2693 23467
rect 2641 23415 2655 23444
rect 2655 23415 2689 23444
rect 2689 23415 2693 23444
rect 697 23351 749 23403
rect 765 23371 817 23403
rect 765 23351 767 23371
rect 767 23351 801 23371
rect 801 23351 817 23371
rect 833 23351 885 23403
rect 901 23351 953 23403
rect 969 23371 1021 23403
rect 969 23351 1003 23371
rect 1003 23351 1021 23371
rect 1037 23351 1089 23403
rect 1105 23351 1157 23403
rect 1173 23351 1225 23403
rect 1241 23371 1293 23403
rect 1241 23351 1273 23371
rect 1273 23351 1293 23371
rect 697 23287 749 23339
rect 765 23337 767 23339
rect 767 23337 801 23339
rect 801 23337 817 23339
rect 765 23298 817 23337
rect 765 23287 767 23298
rect 767 23287 801 23298
rect 801 23287 817 23298
rect 833 23287 885 23339
rect 901 23287 953 23339
rect 969 23337 1003 23339
rect 1003 23337 1021 23339
rect 969 23298 1021 23337
rect 969 23287 1003 23298
rect 1003 23287 1021 23298
rect 1037 23287 1089 23339
rect 1105 23287 1157 23339
rect 1173 23287 1225 23339
rect 1241 23337 1273 23339
rect 1273 23337 1293 23339
rect 2097 23351 2149 23403
rect 2165 23371 2217 23403
rect 2165 23351 2183 23371
rect 2183 23351 2217 23371
rect 2233 23351 2285 23403
rect 2301 23351 2353 23403
rect 2369 23371 2421 23403
rect 2437 23371 2489 23403
rect 2369 23351 2419 23371
rect 2419 23351 2421 23371
rect 2437 23351 2453 23371
rect 2453 23351 2489 23371
rect 2505 23351 2557 23403
rect 2573 23351 2625 23403
rect 2641 23371 2693 23403
rect 2641 23351 2655 23371
rect 2655 23351 2689 23371
rect 2689 23351 2693 23371
rect 1241 23298 1293 23337
rect 1241 23287 1273 23298
rect 1273 23287 1293 23298
rect 697 23223 749 23275
rect 765 23264 767 23275
rect 767 23264 801 23275
rect 801 23264 817 23275
rect 765 23225 817 23264
rect 765 23223 767 23225
rect 767 23223 801 23225
rect 801 23223 817 23225
rect 833 23223 885 23275
rect 901 23223 953 23275
rect 969 23264 1003 23275
rect 1003 23264 1021 23275
rect 969 23225 1021 23264
rect 969 23223 1003 23225
rect 1003 23223 1021 23225
rect 1037 23223 1089 23275
rect 1105 23223 1157 23275
rect 1173 23223 1225 23275
rect 1241 23264 1273 23275
rect 1273 23264 1293 23275
rect 2097 23287 2149 23339
rect 2165 23337 2183 23339
rect 2183 23337 2217 23339
rect 2165 23298 2217 23337
rect 2165 23287 2183 23298
rect 2183 23287 2217 23298
rect 2233 23287 2285 23339
rect 2301 23287 2353 23339
rect 2369 23337 2419 23339
rect 2419 23337 2421 23339
rect 2437 23337 2453 23339
rect 2453 23337 2489 23339
rect 2369 23298 2421 23337
rect 2437 23298 2489 23337
rect 2369 23287 2419 23298
rect 2419 23287 2421 23298
rect 2437 23287 2453 23298
rect 2453 23287 2489 23298
rect 2505 23287 2557 23339
rect 2573 23287 2625 23339
rect 2641 23337 2655 23339
rect 2655 23337 2689 23339
rect 2689 23337 2693 23339
rect 2641 23298 2693 23337
rect 2641 23287 2655 23298
rect 2655 23287 2689 23298
rect 2689 23287 2693 23298
rect 1241 23225 1293 23264
rect 1241 23223 1273 23225
rect 1273 23223 1293 23225
rect 697 23159 749 23211
rect 765 23191 767 23211
rect 767 23191 801 23211
rect 801 23191 817 23211
rect 765 23159 817 23191
rect 833 23159 885 23211
rect 901 23159 953 23211
rect 969 23191 1003 23211
rect 1003 23191 1021 23211
rect 969 23159 1021 23191
rect 1037 23159 1089 23211
rect 1105 23159 1157 23211
rect 1173 23159 1225 23211
rect 1241 23191 1273 23211
rect 1273 23191 1293 23211
rect 2097 23223 2149 23275
rect 2165 23264 2183 23275
rect 2183 23264 2217 23275
rect 2165 23225 2217 23264
rect 2165 23223 2183 23225
rect 2183 23223 2217 23225
rect 2233 23223 2285 23275
rect 2301 23223 2353 23275
rect 2369 23264 2419 23275
rect 2419 23264 2421 23275
rect 2437 23264 2453 23275
rect 2453 23264 2489 23275
rect 2369 23225 2421 23264
rect 2437 23225 2489 23264
rect 2369 23223 2419 23225
rect 2419 23223 2421 23225
rect 2437 23223 2453 23225
rect 2453 23223 2489 23225
rect 2505 23223 2557 23275
rect 2573 23223 2625 23275
rect 2641 23264 2655 23275
rect 2655 23264 2689 23275
rect 2689 23264 2693 23275
rect 2641 23225 2693 23264
rect 2641 23223 2655 23225
rect 2655 23223 2689 23225
rect 2689 23223 2693 23225
rect 1241 23159 1293 23191
rect 2097 23159 2149 23211
rect 2165 23191 2183 23211
rect 2183 23191 2217 23211
rect 2165 23159 2217 23191
rect 2233 23159 2285 23211
rect 2301 23159 2353 23211
rect 2369 23191 2419 23211
rect 2419 23191 2421 23211
rect 2437 23191 2453 23211
rect 2453 23191 2489 23211
rect 2369 23159 2421 23191
rect 2437 23159 2489 23191
rect 2505 23159 2557 23211
rect 2573 23159 2625 23211
rect 2641 23191 2655 23211
rect 2655 23191 2689 23211
rect 2689 23191 2693 23211
rect 2641 23159 2693 23191
rect 697 23095 749 23147
rect 765 23118 767 23147
rect 767 23118 801 23147
rect 801 23118 817 23147
rect 765 23095 817 23118
rect 833 23095 885 23147
rect 901 23095 953 23147
rect 969 23118 1003 23147
rect 1003 23118 1021 23147
rect 969 23095 1021 23118
rect 1037 23095 1089 23147
rect 1105 23095 1157 23147
rect 1173 23095 1225 23147
rect 1241 23118 1273 23147
rect 1273 23118 1293 23147
rect 1241 23095 1293 23118
rect 2097 23095 2149 23147
rect 2165 23118 2183 23147
rect 2183 23118 2217 23147
rect 2165 23095 2217 23118
rect 2233 23095 2285 23147
rect 2301 23095 2353 23147
rect 2369 23118 2419 23147
rect 2419 23118 2421 23147
rect 2437 23118 2453 23147
rect 2453 23118 2489 23147
rect 2369 23095 2421 23118
rect 2437 23095 2489 23118
rect 2505 23095 2557 23147
rect 2573 23095 2625 23147
rect 2641 23118 2655 23147
rect 2655 23118 2689 23147
rect 2689 23118 2693 23147
rect 2641 23095 2693 23118
rect 697 23031 749 23083
rect 765 23078 817 23083
rect 765 23044 767 23078
rect 767 23044 801 23078
rect 801 23044 817 23078
rect 765 23031 817 23044
rect 833 23031 885 23083
rect 901 23031 953 23083
rect 969 23078 1021 23083
rect 969 23044 1003 23078
rect 1003 23044 1021 23078
rect 969 23031 1021 23044
rect 1037 23031 1089 23083
rect 1105 23031 1157 23083
rect 1173 23031 1225 23083
rect 1241 23078 1293 23083
rect 1241 23044 1273 23078
rect 1273 23044 1293 23078
rect 1241 23031 1293 23044
rect 2097 23031 2149 23083
rect 2165 23078 2217 23083
rect 2165 23044 2183 23078
rect 2183 23044 2217 23078
rect 2165 23031 2217 23044
rect 2233 23031 2285 23083
rect 2301 23031 2353 23083
rect 2369 23078 2421 23083
rect 2437 23078 2489 23083
rect 2369 23044 2419 23078
rect 2419 23044 2421 23078
rect 2437 23044 2453 23078
rect 2453 23044 2489 23078
rect 2369 23031 2421 23044
rect 2437 23031 2489 23044
rect 2505 23031 2557 23083
rect 2573 23031 2625 23083
rect 2641 23078 2693 23083
rect 2641 23044 2655 23078
rect 2655 23044 2689 23078
rect 2689 23044 2693 23078
rect 2641 23031 2693 23044
rect 697 22967 749 23019
rect 765 23004 817 23019
rect 765 22970 767 23004
rect 767 22970 801 23004
rect 801 22970 817 23004
rect 765 22967 817 22970
rect 833 22967 885 23019
rect 901 22967 953 23019
rect 969 23004 1021 23019
rect 969 22970 1003 23004
rect 1003 22970 1021 23004
rect 969 22967 1021 22970
rect 1037 22967 1089 23019
rect 1105 22967 1157 23019
rect 1173 22967 1225 23019
rect 1241 23004 1293 23019
rect 1241 22970 1273 23004
rect 1273 22970 1293 23004
rect 1241 22967 1293 22970
rect 2097 22967 2149 23019
rect 2165 23004 2217 23019
rect 2165 22970 2183 23004
rect 2183 22970 2217 23004
rect 2165 22967 2217 22970
rect 2233 22967 2285 23019
rect 2301 22967 2353 23019
rect 2369 23004 2421 23019
rect 2437 23004 2489 23019
rect 2369 22970 2419 23004
rect 2419 22970 2421 23004
rect 2437 22970 2453 23004
rect 2453 22970 2489 23004
rect 2369 22967 2421 22970
rect 2437 22967 2489 22970
rect 2505 22967 2557 23019
rect 2573 22967 2625 23019
rect 2641 23004 2693 23019
rect 2641 22970 2655 23004
rect 2655 22970 2689 23004
rect 2689 22970 2693 23004
rect 2641 22967 2693 22970
rect 697 22903 749 22955
rect 765 22930 817 22955
rect 765 22903 767 22930
rect 767 22903 801 22930
rect 801 22903 817 22930
rect 833 22903 885 22955
rect 901 22903 953 22955
rect 969 22930 1021 22955
rect 969 22903 1003 22930
rect 1003 22903 1021 22930
rect 1037 22903 1089 22955
rect 1105 22903 1157 22955
rect 1173 22903 1225 22955
rect 1241 22930 1293 22955
rect 1241 22903 1273 22930
rect 1273 22903 1293 22930
rect 2097 22903 2149 22955
rect 2165 22930 2217 22955
rect 2165 22903 2183 22930
rect 2183 22903 2217 22930
rect 2233 22903 2285 22955
rect 2301 22903 2353 22955
rect 2369 22930 2421 22955
rect 2437 22930 2489 22955
rect 2369 22903 2419 22930
rect 2419 22903 2421 22930
rect 2437 22903 2453 22930
rect 2453 22903 2489 22930
rect 2505 22903 2557 22955
rect 2573 22903 2625 22955
rect 2641 22930 2693 22955
rect 2641 22903 2655 22930
rect 2655 22903 2689 22930
rect 2689 22903 2693 22930
rect 697 22839 749 22891
rect 765 22856 817 22891
rect 765 22839 767 22856
rect 767 22839 801 22856
rect 801 22839 817 22856
rect 833 22839 885 22891
rect 901 22839 953 22891
rect 969 22856 1021 22891
rect 969 22839 1003 22856
rect 1003 22839 1021 22856
rect 1037 22839 1089 22891
rect 1105 22839 1157 22891
rect 1173 22839 1225 22891
rect 1241 22856 1293 22891
rect 1241 22839 1273 22856
rect 1273 22839 1293 22856
rect 697 22775 749 22827
rect 765 22822 767 22827
rect 767 22822 801 22827
rect 801 22822 817 22827
rect 765 22782 817 22822
rect 765 22775 767 22782
rect 767 22775 801 22782
rect 801 22775 817 22782
rect 833 22775 885 22827
rect 901 22775 953 22827
rect 969 22822 1003 22827
rect 1003 22822 1021 22827
rect 969 22782 1021 22822
rect 969 22775 1003 22782
rect 1003 22775 1021 22782
rect 1037 22775 1089 22827
rect 1105 22775 1157 22827
rect 1173 22775 1225 22827
rect 1241 22822 1273 22827
rect 1273 22822 1293 22827
rect 2097 22839 2149 22891
rect 2165 22856 2217 22891
rect 2165 22839 2183 22856
rect 2183 22839 2217 22856
rect 2233 22839 2285 22891
rect 2301 22839 2353 22891
rect 2369 22856 2421 22891
rect 2437 22856 2489 22891
rect 2369 22839 2419 22856
rect 2419 22839 2421 22856
rect 2437 22839 2453 22856
rect 2453 22839 2489 22856
rect 2505 22839 2557 22891
rect 2573 22839 2625 22891
rect 2641 22856 2693 22891
rect 2641 22839 2655 22856
rect 2655 22839 2689 22856
rect 2689 22839 2693 22856
rect 1241 22782 1293 22822
rect 1241 22775 1273 22782
rect 1273 22775 1293 22782
rect 697 22711 749 22763
rect 765 22748 767 22763
rect 767 22748 801 22763
rect 801 22748 817 22763
rect 765 22711 817 22748
rect 833 22711 885 22763
rect 901 22711 953 22763
rect 969 22748 1003 22763
rect 1003 22748 1021 22763
rect 969 22711 1021 22748
rect 1037 22711 1089 22763
rect 1105 22711 1157 22763
rect 1173 22711 1225 22763
rect 1241 22748 1273 22763
rect 1273 22748 1293 22763
rect 2097 22775 2149 22827
rect 2165 22822 2183 22827
rect 2183 22822 2217 22827
rect 2165 22782 2217 22822
rect 2165 22775 2183 22782
rect 2183 22775 2217 22782
rect 2233 22775 2285 22827
rect 2301 22775 2353 22827
rect 2369 22822 2419 22827
rect 2419 22822 2421 22827
rect 2437 22822 2453 22827
rect 2453 22822 2489 22827
rect 2369 22782 2421 22822
rect 2437 22782 2489 22822
rect 2369 22775 2419 22782
rect 2419 22775 2421 22782
rect 2437 22775 2453 22782
rect 2453 22775 2489 22782
rect 2505 22775 2557 22827
rect 2573 22775 2625 22827
rect 2641 22822 2655 22827
rect 2655 22822 2689 22827
rect 2689 22822 2693 22827
rect 2641 22782 2693 22822
rect 2641 22775 2655 22782
rect 2655 22775 2689 22782
rect 2689 22775 2693 22782
rect 1241 22711 1293 22748
rect 2097 22711 2149 22763
rect 2165 22748 2183 22763
rect 2183 22748 2217 22763
rect 2165 22711 2217 22748
rect 2233 22711 2285 22763
rect 2301 22711 2353 22763
rect 2369 22748 2419 22763
rect 2419 22748 2421 22763
rect 2437 22748 2453 22763
rect 2453 22748 2489 22763
rect 2369 22711 2421 22748
rect 2437 22711 2489 22748
rect 2505 22711 2557 22763
rect 2573 22711 2625 22763
rect 2641 22748 2655 22763
rect 2655 22748 2689 22763
rect 2689 22748 2693 22763
rect 2641 22711 2693 22748
rect 697 22647 749 22699
rect 765 22674 767 22699
rect 767 22674 801 22699
rect 801 22674 817 22699
rect 765 22647 817 22674
rect 833 22647 885 22699
rect 901 22647 953 22699
rect 969 22674 1003 22699
rect 1003 22674 1021 22699
rect 969 22647 1021 22674
rect 1037 22647 1089 22699
rect 1105 22647 1157 22699
rect 1173 22647 1225 22699
rect 1241 22674 1273 22699
rect 1273 22674 1293 22699
rect 1241 22647 1293 22674
rect 2097 22647 2149 22699
rect 2165 22674 2183 22699
rect 2183 22674 2217 22699
rect 2165 22647 2217 22674
rect 2233 22647 2285 22699
rect 2301 22647 2353 22699
rect 2369 22674 2419 22699
rect 2419 22674 2421 22699
rect 2437 22674 2453 22699
rect 2453 22674 2489 22699
rect 2369 22647 2421 22674
rect 2437 22647 2489 22674
rect 2505 22647 2557 22699
rect 2573 22647 2625 22699
rect 2641 22674 2655 22699
rect 2655 22674 2689 22699
rect 2689 22674 2693 22699
rect 2641 22647 2693 22674
rect 697 22583 749 22635
rect 765 22634 817 22635
rect 765 22600 767 22634
rect 767 22600 801 22634
rect 801 22600 817 22634
rect 765 22583 817 22600
rect 833 22583 885 22635
rect 901 22583 953 22635
rect 969 22634 1021 22635
rect 969 22600 1003 22634
rect 1003 22600 1021 22634
rect 969 22583 1021 22600
rect 1037 22583 1089 22635
rect 1105 22583 1157 22635
rect 1173 22583 1225 22635
rect 1241 22634 1293 22635
rect 1241 22600 1273 22634
rect 1273 22600 1293 22634
rect 1241 22583 1293 22600
rect 2097 22583 2149 22635
rect 2165 22634 2217 22635
rect 2165 22600 2183 22634
rect 2183 22600 2217 22634
rect 2165 22583 2217 22600
rect 2233 22583 2285 22635
rect 2301 22583 2353 22635
rect 2369 22634 2421 22635
rect 2437 22634 2489 22635
rect 2369 22600 2419 22634
rect 2419 22600 2421 22634
rect 2437 22600 2453 22634
rect 2453 22600 2489 22634
rect 2369 22583 2421 22600
rect 2437 22583 2489 22600
rect 2505 22583 2557 22635
rect 2573 22583 2625 22635
rect 2641 22634 2693 22635
rect 2641 22600 2655 22634
rect 2655 22600 2689 22634
rect 2689 22600 2693 22634
rect 2641 22583 2693 22600
rect 1501 22014 1553 22023
rect 1569 22014 1621 22023
rect 1636 22014 1688 22023
rect 1703 22014 1755 22023
rect 1770 22014 1822 22023
rect 1837 22014 1889 22023
rect 1501 21980 1525 22014
rect 1525 21980 1553 22014
rect 1569 21980 1600 22014
rect 1600 21980 1621 22014
rect 1636 21980 1674 22014
rect 1674 21980 1688 22014
rect 1703 21980 1708 22014
rect 1708 21980 1748 22014
rect 1748 21980 1755 22014
rect 1770 21980 1782 22014
rect 1782 21980 1822 22014
rect 1837 21980 1856 22014
rect 1856 21980 1889 22014
rect 1501 21971 1553 21980
rect 1569 21971 1621 21980
rect 1636 21971 1688 21980
rect 1703 21971 1755 21980
rect 1770 21971 1822 21980
rect 1837 21971 1889 21980
rect 697 21309 749 21361
rect 765 21328 817 21361
rect 765 21309 767 21328
rect 767 21309 801 21328
rect 801 21309 817 21328
rect 833 21309 885 21361
rect 901 21309 953 21361
rect 969 21328 1021 21361
rect 969 21309 1003 21328
rect 1003 21309 1021 21328
rect 1037 21309 1089 21361
rect 1105 21309 1157 21361
rect 1173 21309 1225 21361
rect 1241 21328 1293 21361
rect 1241 21309 1273 21328
rect 1273 21309 1293 21328
rect 697 21245 749 21297
rect 765 21294 767 21297
rect 767 21294 801 21297
rect 801 21294 817 21297
rect 765 21255 817 21294
rect 765 21245 767 21255
rect 767 21245 801 21255
rect 801 21245 817 21255
rect 833 21245 885 21297
rect 901 21245 953 21297
rect 969 21294 1003 21297
rect 1003 21294 1021 21297
rect 969 21255 1021 21294
rect 969 21245 1003 21255
rect 1003 21245 1021 21255
rect 1037 21245 1089 21297
rect 1105 21245 1157 21297
rect 1173 21245 1225 21297
rect 1241 21294 1273 21297
rect 1273 21294 1293 21297
rect 2097 21309 2149 21361
rect 2165 21328 2217 21361
rect 2165 21309 2183 21328
rect 2183 21309 2217 21328
rect 2233 21309 2285 21361
rect 2301 21309 2353 21361
rect 2369 21328 2421 21361
rect 2437 21328 2489 21361
rect 2369 21309 2419 21328
rect 2419 21309 2421 21328
rect 2437 21309 2453 21328
rect 2453 21309 2489 21328
rect 2505 21309 2557 21361
rect 2573 21309 2625 21361
rect 2641 21328 2693 21361
rect 2641 21309 2655 21328
rect 2655 21309 2689 21328
rect 2689 21309 2693 21328
rect 1241 21255 1293 21294
rect 1241 21245 1273 21255
rect 1273 21245 1293 21255
rect 697 21181 749 21233
rect 765 21221 767 21233
rect 767 21221 801 21233
rect 801 21221 817 21233
rect 765 21182 817 21221
rect 765 21181 767 21182
rect 767 21181 801 21182
rect 801 21181 817 21182
rect 833 21181 885 21233
rect 901 21181 953 21233
rect 969 21221 1003 21233
rect 1003 21221 1021 21233
rect 969 21182 1021 21221
rect 969 21181 1003 21182
rect 1003 21181 1021 21182
rect 1037 21181 1089 21233
rect 1105 21181 1157 21233
rect 1173 21181 1225 21233
rect 1241 21221 1273 21233
rect 1273 21221 1293 21233
rect 2097 21245 2149 21297
rect 2165 21294 2183 21297
rect 2183 21294 2217 21297
rect 2165 21255 2217 21294
rect 2165 21245 2183 21255
rect 2183 21245 2217 21255
rect 2233 21245 2285 21297
rect 2301 21245 2353 21297
rect 2369 21294 2419 21297
rect 2419 21294 2421 21297
rect 2437 21294 2453 21297
rect 2453 21294 2489 21297
rect 2369 21255 2421 21294
rect 2437 21255 2489 21294
rect 2369 21245 2419 21255
rect 2419 21245 2421 21255
rect 2437 21245 2453 21255
rect 2453 21245 2489 21255
rect 2505 21245 2557 21297
rect 2573 21245 2625 21297
rect 2641 21294 2655 21297
rect 2655 21294 2689 21297
rect 2689 21294 2693 21297
rect 2641 21255 2693 21294
rect 2641 21245 2655 21255
rect 2655 21245 2689 21255
rect 2689 21245 2693 21255
rect 1241 21182 1293 21221
rect 1241 21181 1273 21182
rect 1273 21181 1293 21182
rect 697 21117 749 21169
rect 765 21148 767 21169
rect 767 21148 801 21169
rect 801 21148 817 21169
rect 765 21117 817 21148
rect 833 21117 885 21169
rect 901 21117 953 21169
rect 969 21148 1003 21169
rect 1003 21148 1021 21169
rect 969 21117 1021 21148
rect 1037 21117 1089 21169
rect 1105 21117 1157 21169
rect 1173 21117 1225 21169
rect 1241 21148 1273 21169
rect 1273 21148 1293 21169
rect 2097 21181 2149 21233
rect 2165 21221 2183 21233
rect 2183 21221 2217 21233
rect 2165 21182 2217 21221
rect 2165 21181 2183 21182
rect 2183 21181 2217 21182
rect 2233 21181 2285 21233
rect 2301 21181 2353 21233
rect 2369 21221 2419 21233
rect 2419 21221 2421 21233
rect 2437 21221 2453 21233
rect 2453 21221 2489 21233
rect 2369 21182 2421 21221
rect 2437 21182 2489 21221
rect 2369 21181 2419 21182
rect 2419 21181 2421 21182
rect 2437 21181 2453 21182
rect 2453 21181 2489 21182
rect 2505 21181 2557 21233
rect 2573 21181 2625 21233
rect 2641 21221 2655 21233
rect 2655 21221 2689 21233
rect 2689 21221 2693 21233
rect 2641 21182 2693 21221
rect 2641 21181 2655 21182
rect 2655 21181 2689 21182
rect 2689 21181 2693 21182
rect 1241 21117 1293 21148
rect 2097 21117 2149 21169
rect 2165 21148 2183 21169
rect 2183 21148 2217 21169
rect 2165 21117 2217 21148
rect 2233 21117 2285 21169
rect 2301 21117 2353 21169
rect 2369 21148 2419 21169
rect 2419 21148 2421 21169
rect 2437 21148 2453 21169
rect 2453 21148 2489 21169
rect 2369 21117 2421 21148
rect 2437 21117 2489 21148
rect 2505 21117 2557 21169
rect 2573 21117 2625 21169
rect 2641 21148 2655 21169
rect 2655 21148 2689 21169
rect 2689 21148 2693 21169
rect 2641 21117 2693 21148
rect 697 21053 749 21105
rect 765 21075 767 21105
rect 767 21075 801 21105
rect 801 21075 817 21105
rect 765 21053 817 21075
rect 833 21053 885 21105
rect 901 21053 953 21105
rect 969 21075 1003 21105
rect 1003 21075 1021 21105
rect 969 21053 1021 21075
rect 1037 21053 1089 21105
rect 1105 21053 1157 21105
rect 1173 21053 1225 21105
rect 1241 21075 1273 21105
rect 1273 21075 1293 21105
rect 1241 21053 1293 21075
rect 2097 21053 2149 21105
rect 2165 21075 2183 21105
rect 2183 21075 2217 21105
rect 2165 21053 2217 21075
rect 2233 21053 2285 21105
rect 2301 21053 2353 21105
rect 2369 21075 2419 21105
rect 2419 21075 2421 21105
rect 2437 21075 2453 21105
rect 2453 21075 2489 21105
rect 2369 21053 2421 21075
rect 2437 21053 2489 21075
rect 2505 21053 2557 21105
rect 2573 21053 2625 21105
rect 2641 21075 2655 21105
rect 2655 21075 2689 21105
rect 2689 21075 2693 21105
rect 2641 21053 2693 21075
rect 697 20989 749 21041
rect 765 21036 817 21041
rect 765 21002 767 21036
rect 767 21002 801 21036
rect 801 21002 817 21036
rect 765 20989 817 21002
rect 833 20989 885 21041
rect 901 20989 953 21041
rect 969 21036 1021 21041
rect 969 21002 1003 21036
rect 1003 21002 1021 21036
rect 969 20989 1021 21002
rect 1037 20989 1089 21041
rect 1105 20989 1157 21041
rect 1173 20989 1225 21041
rect 1241 21036 1293 21041
rect 1241 21002 1273 21036
rect 1273 21002 1293 21036
rect 1241 20989 1293 21002
rect 2097 20989 2149 21041
rect 2165 21036 2217 21041
rect 2165 21002 2183 21036
rect 2183 21002 2217 21036
rect 2165 20989 2217 21002
rect 2233 20989 2285 21041
rect 2301 20989 2353 21041
rect 2369 21036 2421 21041
rect 2437 21036 2489 21041
rect 2369 21002 2419 21036
rect 2419 21002 2421 21036
rect 2437 21002 2453 21036
rect 2453 21002 2489 21036
rect 2369 20989 2421 21002
rect 2437 20989 2489 21002
rect 2505 20989 2557 21041
rect 2573 20989 2625 21041
rect 2641 21036 2693 21041
rect 2641 21002 2655 21036
rect 2655 21002 2689 21036
rect 2689 21002 2693 21036
rect 2641 20989 2693 21002
rect 697 20925 749 20977
rect 765 20962 817 20977
rect 765 20928 767 20962
rect 767 20928 801 20962
rect 801 20928 817 20962
rect 765 20925 817 20928
rect 833 20925 885 20977
rect 901 20925 953 20977
rect 969 20962 1021 20977
rect 969 20928 1003 20962
rect 1003 20928 1021 20962
rect 969 20925 1021 20928
rect 1037 20925 1089 20977
rect 1105 20925 1157 20977
rect 1173 20925 1225 20977
rect 1241 20962 1293 20977
rect 1241 20928 1273 20962
rect 1273 20928 1293 20962
rect 1241 20925 1293 20928
rect 2097 20925 2149 20977
rect 2165 20962 2217 20977
rect 2165 20928 2183 20962
rect 2183 20928 2217 20962
rect 2165 20925 2217 20928
rect 2233 20925 2285 20977
rect 2301 20925 2353 20977
rect 2369 20962 2421 20977
rect 2437 20962 2489 20977
rect 2369 20928 2419 20962
rect 2419 20928 2421 20962
rect 2437 20928 2453 20962
rect 2453 20928 2489 20962
rect 2369 20925 2421 20928
rect 2437 20925 2489 20928
rect 2505 20925 2557 20977
rect 2573 20925 2625 20977
rect 2641 20962 2693 20977
rect 2641 20928 2655 20962
rect 2655 20928 2689 20962
rect 2689 20928 2693 20962
rect 2641 20925 2693 20928
rect 697 20861 749 20913
rect 765 20888 817 20913
rect 765 20861 767 20888
rect 767 20861 801 20888
rect 801 20861 817 20888
rect 833 20861 885 20913
rect 901 20861 953 20913
rect 969 20888 1021 20913
rect 969 20861 1003 20888
rect 1003 20861 1021 20888
rect 1037 20861 1089 20913
rect 1105 20861 1157 20913
rect 1173 20861 1225 20913
rect 1241 20888 1293 20913
rect 1241 20861 1273 20888
rect 1273 20861 1293 20888
rect 2097 20861 2149 20913
rect 2165 20888 2217 20913
rect 2165 20861 2183 20888
rect 2183 20861 2217 20888
rect 2233 20861 2285 20913
rect 2301 20861 2353 20913
rect 2369 20888 2421 20913
rect 2437 20888 2489 20913
rect 2369 20861 2419 20888
rect 2419 20861 2421 20888
rect 2437 20861 2453 20888
rect 2453 20861 2489 20888
rect 2505 20861 2557 20913
rect 2573 20861 2625 20913
rect 2641 20888 2693 20913
rect 2641 20861 2655 20888
rect 2655 20861 2689 20888
rect 2689 20861 2693 20888
rect 697 20797 749 20849
rect 765 20814 817 20849
rect 765 20797 767 20814
rect 767 20797 801 20814
rect 801 20797 817 20814
rect 833 20797 885 20849
rect 901 20797 953 20849
rect 969 20814 1021 20849
rect 969 20797 1003 20814
rect 1003 20797 1021 20814
rect 1037 20797 1089 20849
rect 1105 20797 1157 20849
rect 1173 20797 1225 20849
rect 1241 20814 1293 20849
rect 1241 20797 1273 20814
rect 1273 20797 1293 20814
rect 697 20733 749 20785
rect 765 20780 767 20785
rect 767 20780 801 20785
rect 801 20780 817 20785
rect 765 20740 817 20780
rect 765 20733 767 20740
rect 767 20733 801 20740
rect 801 20733 817 20740
rect 833 20733 885 20785
rect 901 20733 953 20785
rect 969 20780 1003 20785
rect 1003 20780 1021 20785
rect 969 20740 1021 20780
rect 969 20733 1003 20740
rect 1003 20733 1021 20740
rect 1037 20733 1089 20785
rect 1105 20733 1157 20785
rect 1173 20733 1225 20785
rect 1241 20780 1273 20785
rect 1273 20780 1293 20785
rect 2097 20797 2149 20849
rect 2165 20814 2217 20849
rect 2165 20797 2183 20814
rect 2183 20797 2217 20814
rect 2233 20797 2285 20849
rect 2301 20797 2353 20849
rect 2369 20814 2421 20849
rect 2437 20814 2489 20849
rect 2369 20797 2419 20814
rect 2419 20797 2421 20814
rect 2437 20797 2453 20814
rect 2453 20797 2489 20814
rect 2505 20797 2557 20849
rect 2573 20797 2625 20849
rect 2641 20814 2693 20849
rect 2641 20797 2655 20814
rect 2655 20797 2689 20814
rect 2689 20797 2693 20814
rect 1241 20740 1293 20780
rect 1241 20733 1273 20740
rect 1273 20733 1293 20740
rect 697 20669 749 20721
rect 765 20706 767 20721
rect 767 20706 801 20721
rect 801 20706 817 20721
rect 765 20669 817 20706
rect 833 20669 885 20721
rect 901 20669 953 20721
rect 969 20706 1003 20721
rect 1003 20706 1021 20721
rect 969 20669 1021 20706
rect 1037 20669 1089 20721
rect 1105 20669 1157 20721
rect 1173 20669 1225 20721
rect 1241 20706 1273 20721
rect 1273 20706 1293 20721
rect 2097 20733 2149 20785
rect 2165 20780 2183 20785
rect 2183 20780 2217 20785
rect 2165 20740 2217 20780
rect 2165 20733 2183 20740
rect 2183 20733 2217 20740
rect 2233 20733 2285 20785
rect 2301 20733 2353 20785
rect 2369 20780 2419 20785
rect 2419 20780 2421 20785
rect 2437 20780 2453 20785
rect 2453 20780 2489 20785
rect 2369 20740 2421 20780
rect 2437 20740 2489 20780
rect 2369 20733 2419 20740
rect 2419 20733 2421 20740
rect 2437 20733 2453 20740
rect 2453 20733 2489 20740
rect 2505 20733 2557 20785
rect 2573 20733 2625 20785
rect 2641 20780 2655 20785
rect 2655 20780 2689 20785
rect 2689 20780 2693 20785
rect 2641 20740 2693 20780
rect 2641 20733 2655 20740
rect 2655 20733 2689 20740
rect 2689 20733 2693 20740
rect 1241 20669 1293 20706
rect 2097 20669 2149 20721
rect 2165 20706 2183 20721
rect 2183 20706 2217 20721
rect 2165 20669 2217 20706
rect 2233 20669 2285 20721
rect 2301 20669 2353 20721
rect 2369 20706 2419 20721
rect 2419 20706 2421 20721
rect 2437 20706 2453 20721
rect 2453 20706 2489 20721
rect 2369 20669 2421 20706
rect 2437 20669 2489 20706
rect 2505 20669 2557 20721
rect 2573 20669 2625 20721
rect 2641 20706 2655 20721
rect 2655 20706 2689 20721
rect 2689 20706 2693 20721
rect 2641 20669 2693 20706
rect 697 20605 749 20657
rect 765 20632 767 20657
rect 767 20632 801 20657
rect 801 20632 817 20657
rect 765 20605 817 20632
rect 833 20605 885 20657
rect 901 20605 953 20657
rect 969 20632 1003 20657
rect 1003 20632 1021 20657
rect 969 20605 1021 20632
rect 1037 20605 1089 20657
rect 1105 20605 1157 20657
rect 1173 20605 1225 20657
rect 1241 20632 1273 20657
rect 1273 20632 1293 20657
rect 1241 20605 1293 20632
rect 2097 20605 2149 20657
rect 2165 20632 2183 20657
rect 2183 20632 2217 20657
rect 2165 20605 2217 20632
rect 2233 20605 2285 20657
rect 2301 20605 2353 20657
rect 2369 20632 2419 20657
rect 2419 20632 2421 20657
rect 2437 20632 2453 20657
rect 2453 20632 2489 20657
rect 2369 20605 2421 20632
rect 2437 20605 2489 20632
rect 2505 20605 2557 20657
rect 2573 20605 2625 20657
rect 2641 20632 2655 20657
rect 2655 20632 2689 20657
rect 2689 20632 2693 20657
rect 2641 20605 2693 20632
rect 697 20541 749 20593
rect 765 20592 817 20593
rect 765 20558 767 20592
rect 767 20558 801 20592
rect 801 20558 817 20592
rect 765 20541 817 20558
rect 833 20541 885 20593
rect 901 20541 953 20593
rect 969 20592 1021 20593
rect 969 20558 1003 20592
rect 1003 20558 1021 20592
rect 969 20541 1021 20558
rect 1037 20541 1089 20593
rect 1105 20541 1157 20593
rect 1173 20541 1225 20593
rect 1241 20592 1293 20593
rect 1241 20558 1273 20592
rect 1273 20558 1293 20592
rect 1241 20541 1293 20558
rect 2097 20541 2149 20593
rect 2165 20592 2217 20593
rect 2165 20558 2183 20592
rect 2183 20558 2217 20592
rect 2165 20541 2217 20558
rect 2233 20541 2285 20593
rect 2301 20541 2353 20593
rect 2369 20592 2421 20593
rect 2437 20592 2489 20593
rect 2369 20558 2419 20592
rect 2419 20558 2421 20592
rect 2437 20558 2453 20592
rect 2453 20558 2489 20592
rect 2369 20541 2421 20558
rect 2437 20541 2489 20558
rect 2505 20541 2557 20593
rect 2573 20541 2625 20593
rect 2641 20592 2693 20593
rect 2641 20558 2655 20592
rect 2655 20558 2689 20592
rect 2689 20558 2693 20592
rect 2641 20541 2693 20558
rect 697 20477 749 20529
rect 765 20518 817 20529
rect 765 20484 767 20518
rect 767 20484 801 20518
rect 801 20484 817 20518
rect 765 20477 817 20484
rect 833 20477 885 20529
rect 901 20477 953 20529
rect 969 20518 1021 20529
rect 969 20484 1003 20518
rect 1003 20484 1021 20518
rect 969 20477 1021 20484
rect 1037 20477 1089 20529
rect 1105 20477 1157 20529
rect 1173 20477 1225 20529
rect 1241 20518 1293 20529
rect 1241 20484 1273 20518
rect 1273 20484 1293 20518
rect 1241 20477 1293 20484
rect 2097 20477 2149 20529
rect 2165 20518 2217 20529
rect 2165 20484 2183 20518
rect 2183 20484 2217 20518
rect 2165 20477 2217 20484
rect 2233 20477 2285 20529
rect 2301 20477 2353 20529
rect 2369 20518 2421 20529
rect 2437 20518 2489 20529
rect 2369 20484 2419 20518
rect 2419 20484 2421 20518
rect 2437 20484 2453 20518
rect 2453 20484 2489 20518
rect 2369 20477 2421 20484
rect 2437 20477 2489 20484
rect 2505 20477 2557 20529
rect 2573 20477 2625 20529
rect 2641 20518 2693 20529
rect 2641 20484 2655 20518
rect 2655 20484 2689 20518
rect 2689 20484 2693 20518
rect 2641 20477 2693 20484
rect 697 20413 749 20465
rect 765 20444 817 20465
rect 765 20413 767 20444
rect 767 20413 801 20444
rect 801 20413 817 20444
rect 833 20413 885 20465
rect 901 20413 953 20465
rect 969 20444 1021 20465
rect 969 20413 1003 20444
rect 1003 20413 1021 20444
rect 1037 20413 1089 20465
rect 1105 20413 1157 20465
rect 1173 20413 1225 20465
rect 1241 20444 1293 20465
rect 1241 20413 1273 20444
rect 1273 20413 1293 20444
rect 2097 20413 2149 20465
rect 2165 20444 2217 20465
rect 2165 20413 2183 20444
rect 2183 20413 2217 20444
rect 2233 20413 2285 20465
rect 2301 20413 2353 20465
rect 2369 20444 2421 20465
rect 2437 20444 2489 20465
rect 2369 20413 2419 20444
rect 2419 20413 2421 20444
rect 2437 20413 2453 20444
rect 2453 20413 2489 20444
rect 2505 20413 2557 20465
rect 2573 20413 2625 20465
rect 2641 20444 2693 20465
rect 2641 20413 2655 20444
rect 2655 20413 2689 20444
rect 2689 20413 2693 20444
rect 1501 19884 1553 19893
rect 1569 19884 1621 19893
rect 1636 19884 1688 19893
rect 1703 19884 1755 19893
rect 1770 19884 1822 19893
rect 1837 19884 1889 19893
rect 1501 19850 1525 19884
rect 1525 19850 1553 19884
rect 1569 19850 1600 19884
rect 1600 19850 1621 19884
rect 1636 19850 1674 19884
rect 1674 19850 1688 19884
rect 1703 19850 1708 19884
rect 1708 19850 1748 19884
rect 1748 19850 1755 19884
rect 1770 19850 1782 19884
rect 1782 19850 1822 19884
rect 1837 19850 1856 19884
rect 1856 19850 1889 19884
rect 1501 19841 1553 19850
rect 1569 19841 1621 19850
rect 1636 19841 1688 19850
rect 1703 19841 1755 19850
rect 1770 19841 1822 19850
rect 1837 19841 1889 19850
rect 697 19205 749 19257
rect 765 19223 767 19257
rect 767 19223 801 19257
rect 801 19223 817 19257
rect 765 19205 817 19223
rect 833 19205 885 19257
rect 901 19205 953 19257
rect 969 19223 1003 19257
rect 1003 19223 1021 19257
rect 969 19205 1021 19223
rect 1037 19205 1089 19257
rect 1105 19205 1157 19257
rect 1173 19205 1225 19257
rect 1241 19223 1273 19257
rect 1273 19223 1293 19257
rect 1241 19205 1293 19223
rect 2097 19205 2149 19257
rect 2165 19223 2183 19257
rect 2183 19223 2217 19257
rect 2165 19205 2217 19223
rect 2233 19205 2285 19257
rect 2301 19205 2353 19257
rect 2369 19223 2419 19257
rect 2419 19223 2421 19257
rect 2437 19223 2453 19257
rect 2453 19223 2489 19257
rect 2369 19205 2421 19223
rect 2437 19205 2489 19223
rect 2505 19205 2557 19257
rect 2573 19205 2625 19257
rect 2641 19223 2655 19257
rect 2655 19223 2689 19257
rect 2689 19223 2693 19257
rect 2641 19205 2693 19223
rect 697 19141 749 19193
rect 765 19184 817 19193
rect 765 19150 767 19184
rect 767 19150 801 19184
rect 801 19150 817 19184
rect 765 19141 817 19150
rect 833 19141 885 19193
rect 901 19141 953 19193
rect 969 19184 1021 19193
rect 969 19150 1003 19184
rect 1003 19150 1021 19184
rect 969 19141 1021 19150
rect 1037 19141 1089 19193
rect 1105 19141 1157 19193
rect 1173 19141 1225 19193
rect 1241 19184 1293 19193
rect 1241 19150 1273 19184
rect 1273 19150 1293 19184
rect 1241 19141 1293 19150
rect 2097 19141 2149 19193
rect 2165 19184 2217 19193
rect 2165 19150 2183 19184
rect 2183 19150 2217 19184
rect 2165 19141 2217 19150
rect 2233 19141 2285 19193
rect 2301 19141 2353 19193
rect 2369 19184 2421 19193
rect 2437 19184 2489 19193
rect 2369 19150 2419 19184
rect 2419 19150 2421 19184
rect 2437 19150 2453 19184
rect 2453 19150 2489 19184
rect 2369 19141 2421 19150
rect 2437 19141 2489 19150
rect 2505 19141 2557 19193
rect 2573 19141 2625 19193
rect 2641 19184 2693 19193
rect 2641 19150 2655 19184
rect 2655 19150 2689 19184
rect 2689 19150 2693 19184
rect 2641 19141 2693 19150
rect 697 19077 749 19129
rect 765 19111 817 19129
rect 765 19077 767 19111
rect 767 19077 801 19111
rect 801 19077 817 19111
rect 833 19077 885 19129
rect 901 19077 953 19129
rect 969 19111 1021 19129
rect 969 19077 1003 19111
rect 1003 19077 1021 19111
rect 1037 19077 1089 19129
rect 1105 19077 1157 19129
rect 1173 19077 1225 19129
rect 1241 19111 1293 19129
rect 1241 19077 1273 19111
rect 1273 19077 1293 19111
rect 2097 19077 2149 19129
rect 2165 19111 2217 19129
rect 2165 19077 2183 19111
rect 2183 19077 2217 19111
rect 2233 19077 2285 19129
rect 2301 19077 2353 19129
rect 2369 19111 2421 19129
rect 2437 19111 2489 19129
rect 2369 19077 2419 19111
rect 2419 19077 2421 19111
rect 2437 19077 2453 19111
rect 2453 19077 2489 19111
rect 2505 19077 2557 19129
rect 2573 19077 2625 19129
rect 2641 19111 2693 19129
rect 2641 19077 2655 19111
rect 2655 19077 2689 19111
rect 2689 19077 2693 19111
rect 697 19013 749 19065
rect 765 19038 817 19065
rect 765 19013 767 19038
rect 767 19013 801 19038
rect 801 19013 817 19038
rect 833 19013 885 19065
rect 901 19013 953 19065
rect 969 19038 1021 19065
rect 969 19013 1003 19038
rect 1003 19013 1021 19038
rect 1037 19013 1089 19065
rect 1105 19013 1157 19065
rect 1173 19013 1225 19065
rect 1241 19038 1293 19065
rect 1241 19013 1273 19038
rect 1273 19013 1293 19038
rect 2097 19013 2149 19065
rect 2165 19038 2217 19065
rect 2165 19013 2183 19038
rect 2183 19013 2217 19038
rect 2233 19013 2285 19065
rect 2301 19013 2353 19065
rect 2369 19038 2421 19065
rect 2437 19038 2489 19065
rect 2369 19013 2419 19038
rect 2419 19013 2421 19038
rect 2437 19013 2453 19038
rect 2453 19013 2489 19038
rect 2505 19013 2557 19065
rect 2573 19013 2625 19065
rect 2641 19038 2693 19065
rect 2641 19013 2655 19038
rect 2655 19013 2689 19038
rect 2689 19013 2693 19038
rect 697 18949 749 19001
rect 765 18965 817 19001
rect 765 18949 767 18965
rect 767 18949 801 18965
rect 801 18949 817 18965
rect 833 18949 885 19001
rect 901 18949 953 19001
rect 969 18965 1021 19001
rect 969 18949 1003 18965
rect 1003 18949 1021 18965
rect 1037 18949 1089 19001
rect 1105 18949 1157 19001
rect 1173 18949 1225 19001
rect 1241 18965 1293 19001
rect 1241 18949 1273 18965
rect 1273 18949 1293 18965
rect 697 18885 749 18937
rect 765 18931 767 18937
rect 767 18931 801 18937
rect 801 18931 817 18937
rect 765 18892 817 18931
rect 765 18885 767 18892
rect 767 18885 801 18892
rect 801 18885 817 18892
rect 833 18885 885 18937
rect 901 18885 953 18937
rect 969 18931 1003 18937
rect 1003 18931 1021 18937
rect 969 18892 1021 18931
rect 969 18885 1003 18892
rect 1003 18885 1021 18892
rect 1037 18885 1089 18937
rect 1105 18885 1157 18937
rect 1173 18885 1225 18937
rect 1241 18931 1273 18937
rect 1273 18931 1293 18937
rect 2097 18949 2149 19001
rect 2165 18965 2217 19001
rect 2165 18949 2183 18965
rect 2183 18949 2217 18965
rect 2233 18949 2285 19001
rect 2301 18949 2353 19001
rect 2369 18965 2421 19001
rect 2437 18965 2489 19001
rect 2369 18949 2419 18965
rect 2419 18949 2421 18965
rect 2437 18949 2453 18965
rect 2453 18949 2489 18965
rect 2505 18949 2557 19001
rect 2573 18949 2625 19001
rect 2641 18965 2693 19001
rect 2641 18949 2655 18965
rect 2655 18949 2689 18965
rect 2689 18949 2693 18965
rect 1241 18892 1293 18931
rect 1241 18885 1273 18892
rect 1273 18885 1293 18892
rect 697 18821 749 18873
rect 765 18858 767 18873
rect 767 18858 801 18873
rect 801 18858 817 18873
rect 765 18821 817 18858
rect 833 18821 885 18873
rect 901 18821 953 18873
rect 969 18858 1003 18873
rect 1003 18858 1021 18873
rect 969 18821 1021 18858
rect 1037 18821 1089 18873
rect 1105 18821 1157 18873
rect 1173 18821 1225 18873
rect 1241 18858 1273 18873
rect 1273 18858 1293 18873
rect 2097 18885 2149 18937
rect 2165 18931 2183 18937
rect 2183 18931 2217 18937
rect 2165 18892 2217 18931
rect 2165 18885 2183 18892
rect 2183 18885 2217 18892
rect 2233 18885 2285 18937
rect 2301 18885 2353 18937
rect 2369 18931 2419 18937
rect 2419 18931 2421 18937
rect 2437 18931 2453 18937
rect 2453 18931 2489 18937
rect 2369 18892 2421 18931
rect 2437 18892 2489 18931
rect 2369 18885 2419 18892
rect 2419 18885 2421 18892
rect 2437 18885 2453 18892
rect 2453 18885 2489 18892
rect 2505 18885 2557 18937
rect 2573 18885 2625 18937
rect 2641 18931 2655 18937
rect 2655 18931 2689 18937
rect 2689 18931 2693 18937
rect 2641 18892 2693 18931
rect 2641 18885 2655 18892
rect 2655 18885 2689 18892
rect 2689 18885 2693 18892
rect 1241 18821 1293 18858
rect 2097 18821 2149 18873
rect 2165 18858 2183 18873
rect 2183 18858 2217 18873
rect 2165 18821 2217 18858
rect 2233 18821 2285 18873
rect 2301 18821 2353 18873
rect 2369 18858 2419 18873
rect 2419 18858 2421 18873
rect 2437 18858 2453 18873
rect 2453 18858 2489 18873
rect 2369 18821 2421 18858
rect 2437 18821 2489 18858
rect 2505 18821 2557 18873
rect 2573 18821 2625 18873
rect 2641 18858 2655 18873
rect 2655 18858 2689 18873
rect 2689 18858 2693 18873
rect 2641 18821 2693 18858
rect 697 18757 749 18809
rect 765 18784 767 18809
rect 767 18784 801 18809
rect 801 18784 817 18809
rect 765 18757 817 18784
rect 833 18757 885 18809
rect 901 18757 953 18809
rect 969 18784 1003 18809
rect 1003 18784 1021 18809
rect 969 18757 1021 18784
rect 1037 18757 1089 18809
rect 1105 18757 1157 18809
rect 1173 18757 1225 18809
rect 1241 18784 1273 18809
rect 1273 18784 1293 18809
rect 1241 18757 1293 18784
rect 2097 18757 2149 18809
rect 2165 18784 2183 18809
rect 2183 18784 2217 18809
rect 2165 18757 2217 18784
rect 2233 18757 2285 18809
rect 2301 18757 2353 18809
rect 2369 18784 2419 18809
rect 2419 18784 2421 18809
rect 2437 18784 2453 18809
rect 2453 18784 2489 18809
rect 2369 18757 2421 18784
rect 2437 18757 2489 18784
rect 2505 18757 2557 18809
rect 2573 18757 2625 18809
rect 2641 18784 2655 18809
rect 2655 18784 2689 18809
rect 2689 18784 2693 18809
rect 2641 18757 2693 18784
rect 697 18693 749 18745
rect 765 18744 817 18745
rect 765 18710 767 18744
rect 767 18710 801 18744
rect 801 18710 817 18744
rect 765 18693 817 18710
rect 833 18693 885 18745
rect 901 18693 953 18745
rect 969 18744 1021 18745
rect 969 18710 1003 18744
rect 1003 18710 1021 18744
rect 969 18693 1021 18710
rect 1037 18693 1089 18745
rect 1105 18693 1157 18745
rect 1173 18693 1225 18745
rect 1241 18744 1293 18745
rect 1241 18710 1273 18744
rect 1273 18710 1293 18744
rect 1241 18693 1293 18710
rect 2097 18693 2149 18745
rect 2165 18744 2217 18745
rect 2165 18710 2183 18744
rect 2183 18710 2217 18744
rect 2165 18693 2217 18710
rect 2233 18693 2285 18745
rect 2301 18693 2353 18745
rect 2369 18744 2421 18745
rect 2437 18744 2489 18745
rect 2369 18710 2419 18744
rect 2419 18710 2421 18744
rect 2437 18710 2453 18744
rect 2453 18710 2489 18744
rect 2369 18693 2421 18710
rect 2437 18693 2489 18710
rect 2505 18693 2557 18745
rect 2573 18693 2625 18745
rect 2641 18744 2693 18745
rect 2641 18710 2655 18744
rect 2655 18710 2689 18744
rect 2689 18710 2693 18744
rect 2641 18693 2693 18710
rect 697 18629 749 18681
rect 765 18670 817 18681
rect 765 18636 767 18670
rect 767 18636 801 18670
rect 801 18636 817 18670
rect 765 18629 817 18636
rect 833 18629 885 18681
rect 901 18629 953 18681
rect 969 18670 1021 18681
rect 969 18636 1003 18670
rect 1003 18636 1021 18670
rect 969 18629 1021 18636
rect 1037 18629 1089 18681
rect 1105 18629 1157 18681
rect 1173 18629 1225 18681
rect 1241 18670 1293 18681
rect 1241 18636 1273 18670
rect 1273 18636 1293 18670
rect 1241 18629 1293 18636
rect 2097 18629 2149 18681
rect 2165 18670 2217 18681
rect 2165 18636 2183 18670
rect 2183 18636 2217 18670
rect 2165 18629 2217 18636
rect 2233 18629 2285 18681
rect 2301 18629 2353 18681
rect 2369 18670 2421 18681
rect 2437 18670 2489 18681
rect 2369 18636 2419 18670
rect 2419 18636 2421 18670
rect 2437 18636 2453 18670
rect 2453 18636 2489 18670
rect 2369 18629 2421 18636
rect 2437 18629 2489 18636
rect 2505 18629 2557 18681
rect 2573 18629 2625 18681
rect 2641 18670 2693 18681
rect 2641 18636 2655 18670
rect 2655 18636 2689 18670
rect 2689 18636 2693 18670
rect 2641 18629 2693 18636
rect 697 18565 749 18617
rect 765 18596 817 18617
rect 765 18565 767 18596
rect 767 18565 801 18596
rect 801 18565 817 18596
rect 833 18565 885 18617
rect 901 18565 953 18617
rect 969 18596 1021 18617
rect 969 18565 1003 18596
rect 1003 18565 1021 18596
rect 1037 18565 1089 18617
rect 1105 18565 1157 18617
rect 1173 18565 1225 18617
rect 1241 18596 1293 18617
rect 1241 18565 1273 18596
rect 1273 18565 1293 18596
rect 2097 18565 2149 18617
rect 2165 18596 2217 18617
rect 2165 18565 2183 18596
rect 2183 18565 2217 18596
rect 2233 18565 2285 18617
rect 2301 18565 2353 18617
rect 2369 18596 2421 18617
rect 2437 18596 2489 18617
rect 2369 18565 2419 18596
rect 2419 18565 2421 18596
rect 2437 18565 2453 18596
rect 2453 18565 2489 18596
rect 2505 18565 2557 18617
rect 2573 18565 2625 18617
rect 2641 18596 2693 18617
rect 2641 18565 2655 18596
rect 2655 18565 2689 18596
rect 2689 18565 2693 18596
rect 697 18501 749 18553
rect 765 18522 817 18553
rect 765 18501 767 18522
rect 767 18501 801 18522
rect 801 18501 817 18522
rect 833 18501 885 18553
rect 901 18501 953 18553
rect 969 18522 1021 18553
rect 969 18501 1003 18522
rect 1003 18501 1021 18522
rect 1037 18501 1089 18553
rect 1105 18501 1157 18553
rect 1173 18501 1225 18553
rect 1241 18522 1293 18553
rect 1241 18501 1273 18522
rect 1273 18501 1293 18522
rect 697 18437 749 18489
rect 765 18488 767 18489
rect 767 18488 801 18489
rect 801 18488 817 18489
rect 765 18448 817 18488
rect 765 18437 767 18448
rect 767 18437 801 18448
rect 801 18437 817 18448
rect 833 18437 885 18489
rect 901 18437 953 18489
rect 969 18488 1003 18489
rect 1003 18488 1021 18489
rect 969 18448 1021 18488
rect 969 18437 1003 18448
rect 1003 18437 1021 18448
rect 1037 18437 1089 18489
rect 1105 18437 1157 18489
rect 1173 18437 1225 18489
rect 1241 18488 1273 18489
rect 1273 18488 1293 18489
rect 2097 18501 2149 18553
rect 2165 18522 2217 18553
rect 2165 18501 2183 18522
rect 2183 18501 2217 18522
rect 2233 18501 2285 18553
rect 2301 18501 2353 18553
rect 2369 18522 2421 18553
rect 2437 18522 2489 18553
rect 2369 18501 2419 18522
rect 2419 18501 2421 18522
rect 2437 18501 2453 18522
rect 2453 18501 2489 18522
rect 2505 18501 2557 18553
rect 2573 18501 2625 18553
rect 2641 18522 2693 18553
rect 2641 18501 2655 18522
rect 2655 18501 2689 18522
rect 2689 18501 2693 18522
rect 1241 18448 1293 18488
rect 1241 18437 1273 18448
rect 1273 18437 1293 18448
rect 697 18373 749 18425
rect 765 18414 767 18425
rect 767 18414 801 18425
rect 801 18414 817 18425
rect 765 18374 817 18414
rect 765 18373 767 18374
rect 767 18373 801 18374
rect 801 18373 817 18374
rect 833 18373 885 18425
rect 901 18373 953 18425
rect 969 18414 1003 18425
rect 1003 18414 1021 18425
rect 969 18374 1021 18414
rect 969 18373 1003 18374
rect 1003 18373 1021 18374
rect 1037 18373 1089 18425
rect 1105 18373 1157 18425
rect 1173 18373 1225 18425
rect 1241 18414 1273 18425
rect 1273 18414 1293 18425
rect 2097 18437 2149 18489
rect 2165 18488 2183 18489
rect 2183 18488 2217 18489
rect 2165 18448 2217 18488
rect 2165 18437 2183 18448
rect 2183 18437 2217 18448
rect 2233 18437 2285 18489
rect 2301 18437 2353 18489
rect 2369 18488 2419 18489
rect 2419 18488 2421 18489
rect 2437 18488 2453 18489
rect 2453 18488 2489 18489
rect 2369 18448 2421 18488
rect 2437 18448 2489 18488
rect 2369 18437 2419 18448
rect 2419 18437 2421 18448
rect 2437 18437 2453 18448
rect 2453 18437 2489 18448
rect 2505 18437 2557 18489
rect 2573 18437 2625 18489
rect 2641 18488 2655 18489
rect 2655 18488 2689 18489
rect 2689 18488 2693 18489
rect 2641 18448 2693 18488
rect 2641 18437 2655 18448
rect 2655 18437 2689 18448
rect 2689 18437 2693 18448
rect 1241 18374 1293 18414
rect 1241 18373 1273 18374
rect 1273 18373 1293 18374
rect 697 18309 749 18361
rect 765 18340 767 18361
rect 767 18340 801 18361
rect 801 18340 817 18361
rect 765 18309 817 18340
rect 833 18309 885 18361
rect 901 18309 953 18361
rect 969 18340 1003 18361
rect 1003 18340 1021 18361
rect 969 18309 1021 18340
rect 1037 18309 1089 18361
rect 1105 18309 1157 18361
rect 1173 18309 1225 18361
rect 1241 18340 1273 18361
rect 1273 18340 1293 18361
rect 2097 18373 2149 18425
rect 2165 18414 2183 18425
rect 2183 18414 2217 18425
rect 2165 18374 2217 18414
rect 2165 18373 2183 18374
rect 2183 18373 2217 18374
rect 2233 18373 2285 18425
rect 2301 18373 2353 18425
rect 2369 18414 2419 18425
rect 2419 18414 2421 18425
rect 2437 18414 2453 18425
rect 2453 18414 2489 18425
rect 2369 18374 2421 18414
rect 2437 18374 2489 18414
rect 2369 18373 2419 18374
rect 2419 18373 2421 18374
rect 2437 18373 2453 18374
rect 2453 18373 2489 18374
rect 2505 18373 2557 18425
rect 2573 18373 2625 18425
rect 2641 18414 2655 18425
rect 2655 18414 2689 18425
rect 2689 18414 2693 18425
rect 2641 18374 2693 18414
rect 2641 18373 2655 18374
rect 2655 18373 2689 18374
rect 2689 18373 2693 18374
rect 1241 18309 1293 18340
rect 2097 18309 2149 18361
rect 2165 18340 2183 18361
rect 2183 18340 2217 18361
rect 2165 18309 2217 18340
rect 2233 18309 2285 18361
rect 2301 18309 2353 18361
rect 2369 18340 2419 18361
rect 2419 18340 2421 18361
rect 2437 18340 2453 18361
rect 2453 18340 2489 18361
rect 2369 18309 2421 18340
rect 2437 18309 2489 18340
rect 2505 18309 2557 18361
rect 2573 18309 2625 18361
rect 2641 18340 2655 18361
rect 2655 18340 2689 18361
rect 2689 18340 2693 18361
rect 2641 18309 2693 18340
rect 1501 17754 1553 17763
rect 1569 17754 1621 17763
rect 1636 17754 1688 17763
rect 1703 17754 1755 17763
rect 1770 17754 1822 17763
rect 1837 17754 1889 17763
rect 1501 17720 1525 17754
rect 1525 17720 1553 17754
rect 1569 17720 1600 17754
rect 1600 17720 1621 17754
rect 1636 17720 1674 17754
rect 1674 17720 1688 17754
rect 1703 17720 1708 17754
rect 1708 17720 1748 17754
rect 1748 17720 1755 17754
rect 1770 17720 1782 17754
rect 1782 17720 1822 17754
rect 1837 17720 1856 17754
rect 1856 17720 1889 17754
rect 1501 17711 1553 17720
rect 1569 17711 1621 17720
rect 1636 17711 1688 17720
rect 1703 17711 1755 17720
rect 1770 17711 1822 17720
rect 1837 17711 1889 17720
rect 697 17094 749 17146
rect 765 17141 817 17146
rect 765 17107 767 17141
rect 767 17107 801 17141
rect 801 17107 817 17141
rect 765 17094 817 17107
rect 833 17094 885 17146
rect 901 17094 953 17146
rect 969 17141 1021 17146
rect 969 17107 1003 17141
rect 1003 17107 1021 17141
rect 969 17094 1021 17107
rect 1037 17094 1089 17146
rect 1105 17094 1157 17146
rect 1173 17094 1225 17146
rect 1241 17141 1293 17146
rect 1241 17107 1273 17141
rect 1273 17107 1293 17141
rect 1241 17094 1293 17107
rect 2097 17094 2149 17146
rect 2165 17141 2217 17146
rect 2165 17107 2183 17141
rect 2183 17107 2217 17141
rect 2165 17094 2217 17107
rect 2233 17094 2285 17146
rect 2301 17094 2353 17146
rect 2369 17141 2421 17146
rect 2437 17141 2489 17146
rect 2369 17107 2419 17141
rect 2419 17107 2421 17141
rect 2437 17107 2453 17141
rect 2453 17107 2489 17141
rect 2369 17094 2421 17107
rect 2437 17094 2489 17107
rect 2505 17094 2557 17146
rect 2573 17094 2625 17146
rect 2641 17141 2693 17146
rect 2641 17107 2655 17141
rect 2655 17107 2689 17141
rect 2689 17107 2693 17141
rect 2641 17094 2693 17107
rect 697 17030 749 17082
rect 765 17068 817 17082
rect 765 17034 767 17068
rect 767 17034 801 17068
rect 801 17034 817 17068
rect 765 17030 817 17034
rect 833 17030 885 17082
rect 901 17030 953 17082
rect 969 17068 1021 17082
rect 969 17034 1003 17068
rect 1003 17034 1021 17068
rect 969 17030 1021 17034
rect 1037 17030 1089 17082
rect 1105 17030 1157 17082
rect 1173 17030 1225 17082
rect 1241 17068 1293 17082
rect 1241 17034 1273 17068
rect 1273 17034 1293 17068
rect 1241 17030 1293 17034
rect 2097 17030 2149 17082
rect 2165 17068 2217 17082
rect 2165 17034 2183 17068
rect 2183 17034 2217 17068
rect 2165 17030 2217 17034
rect 2233 17030 2285 17082
rect 2301 17030 2353 17082
rect 2369 17068 2421 17082
rect 2437 17068 2489 17082
rect 2369 17034 2419 17068
rect 2419 17034 2421 17068
rect 2437 17034 2453 17068
rect 2453 17034 2489 17068
rect 2369 17030 2421 17034
rect 2437 17030 2489 17034
rect 2505 17030 2557 17082
rect 2573 17030 2625 17082
rect 2641 17068 2693 17082
rect 2641 17034 2655 17068
rect 2655 17034 2689 17068
rect 2689 17034 2693 17068
rect 2641 17030 2693 17034
rect 697 16966 749 17018
rect 765 16995 817 17018
rect 765 16966 767 16995
rect 767 16966 801 16995
rect 801 16966 817 16995
rect 833 16966 885 17018
rect 901 16966 953 17018
rect 969 16995 1021 17018
rect 969 16966 1003 16995
rect 1003 16966 1021 16995
rect 1037 16966 1089 17018
rect 1105 16966 1157 17018
rect 1173 16966 1225 17018
rect 1241 16995 1293 17018
rect 1241 16966 1273 16995
rect 1273 16966 1293 16995
rect 2097 16966 2149 17018
rect 2165 16995 2217 17018
rect 2165 16966 2183 16995
rect 2183 16966 2217 16995
rect 2233 16966 2285 17018
rect 2301 16966 2353 17018
rect 2369 16995 2421 17018
rect 2437 16995 2489 17018
rect 2369 16966 2419 16995
rect 2419 16966 2421 16995
rect 2437 16966 2453 16995
rect 2453 16966 2489 16995
rect 2505 16966 2557 17018
rect 2573 16966 2625 17018
rect 2641 16995 2693 17018
rect 2641 16966 2655 16995
rect 2655 16966 2689 16995
rect 2689 16966 2693 16995
rect 697 16902 749 16954
rect 765 16922 817 16954
rect 765 16902 767 16922
rect 767 16902 801 16922
rect 801 16902 817 16922
rect 833 16902 885 16954
rect 901 16902 953 16954
rect 969 16922 1021 16954
rect 969 16902 1003 16922
rect 1003 16902 1021 16922
rect 1037 16902 1089 16954
rect 1105 16902 1157 16954
rect 1173 16902 1225 16954
rect 1241 16922 1293 16954
rect 1241 16902 1273 16922
rect 1273 16902 1293 16922
rect 697 16838 749 16890
rect 765 16888 767 16890
rect 767 16888 801 16890
rect 801 16888 817 16890
rect 765 16849 817 16888
rect 765 16838 767 16849
rect 767 16838 801 16849
rect 801 16838 817 16849
rect 833 16838 885 16890
rect 901 16838 953 16890
rect 969 16888 1003 16890
rect 1003 16888 1021 16890
rect 969 16849 1021 16888
rect 969 16838 1003 16849
rect 1003 16838 1021 16849
rect 1037 16838 1089 16890
rect 1105 16838 1157 16890
rect 1173 16838 1225 16890
rect 1241 16888 1273 16890
rect 1273 16888 1293 16890
rect 2097 16902 2149 16954
rect 2165 16922 2217 16954
rect 2165 16902 2183 16922
rect 2183 16902 2217 16922
rect 2233 16902 2285 16954
rect 2301 16902 2353 16954
rect 2369 16922 2421 16954
rect 2437 16922 2489 16954
rect 2369 16902 2419 16922
rect 2419 16902 2421 16922
rect 2437 16902 2453 16922
rect 2453 16902 2489 16922
rect 2505 16902 2557 16954
rect 2573 16902 2625 16954
rect 2641 16922 2693 16954
rect 2641 16902 2655 16922
rect 2655 16902 2689 16922
rect 2689 16902 2693 16922
rect 1241 16849 1293 16888
rect 1241 16838 1273 16849
rect 1273 16838 1293 16849
rect 697 16774 749 16826
rect 765 16815 767 16826
rect 767 16815 801 16826
rect 801 16815 817 16826
rect 765 16776 817 16815
rect 765 16774 767 16776
rect 767 16774 801 16776
rect 801 16774 817 16776
rect 833 16774 885 16826
rect 901 16774 953 16826
rect 969 16815 1003 16826
rect 1003 16815 1021 16826
rect 969 16776 1021 16815
rect 969 16774 1003 16776
rect 1003 16774 1021 16776
rect 1037 16774 1089 16826
rect 1105 16774 1157 16826
rect 1173 16774 1225 16826
rect 1241 16815 1273 16826
rect 1273 16815 1293 16826
rect 2097 16838 2149 16890
rect 2165 16888 2183 16890
rect 2183 16888 2217 16890
rect 2165 16849 2217 16888
rect 2165 16838 2183 16849
rect 2183 16838 2217 16849
rect 2233 16838 2285 16890
rect 2301 16838 2353 16890
rect 2369 16888 2419 16890
rect 2419 16888 2421 16890
rect 2437 16888 2453 16890
rect 2453 16888 2489 16890
rect 2369 16849 2421 16888
rect 2437 16849 2489 16888
rect 2369 16838 2419 16849
rect 2419 16838 2421 16849
rect 2437 16838 2453 16849
rect 2453 16838 2489 16849
rect 2505 16838 2557 16890
rect 2573 16838 2625 16890
rect 2641 16888 2655 16890
rect 2655 16888 2689 16890
rect 2689 16888 2693 16890
rect 2641 16849 2693 16888
rect 2641 16838 2655 16849
rect 2655 16838 2689 16849
rect 2689 16838 2693 16849
rect 1241 16776 1293 16815
rect 1241 16774 1273 16776
rect 1273 16774 1293 16776
rect 697 16710 749 16762
rect 765 16742 767 16762
rect 767 16742 801 16762
rect 801 16742 817 16762
rect 765 16710 817 16742
rect 833 16710 885 16762
rect 901 16710 953 16762
rect 969 16742 1003 16762
rect 1003 16742 1021 16762
rect 969 16710 1021 16742
rect 1037 16710 1089 16762
rect 1105 16710 1157 16762
rect 1173 16710 1225 16762
rect 1241 16742 1273 16762
rect 1273 16742 1293 16762
rect 2097 16774 2149 16826
rect 2165 16815 2183 16826
rect 2183 16815 2217 16826
rect 2165 16776 2217 16815
rect 2165 16774 2183 16776
rect 2183 16774 2217 16776
rect 2233 16774 2285 16826
rect 2301 16774 2353 16826
rect 2369 16815 2419 16826
rect 2419 16815 2421 16826
rect 2437 16815 2453 16826
rect 2453 16815 2489 16826
rect 2369 16776 2421 16815
rect 2437 16776 2489 16815
rect 2369 16774 2419 16776
rect 2419 16774 2421 16776
rect 2437 16774 2453 16776
rect 2453 16774 2489 16776
rect 2505 16774 2557 16826
rect 2573 16774 2625 16826
rect 2641 16815 2655 16826
rect 2655 16815 2689 16826
rect 2689 16815 2693 16826
rect 2641 16776 2693 16815
rect 2641 16774 2655 16776
rect 2655 16774 2689 16776
rect 2689 16774 2693 16776
rect 1241 16710 1293 16742
rect 2097 16710 2149 16762
rect 2165 16742 2183 16762
rect 2183 16742 2217 16762
rect 2165 16710 2217 16742
rect 2233 16710 2285 16762
rect 2301 16710 2353 16762
rect 2369 16742 2419 16762
rect 2419 16742 2421 16762
rect 2437 16742 2453 16762
rect 2453 16742 2489 16762
rect 2369 16710 2421 16742
rect 2437 16710 2489 16742
rect 2505 16710 2557 16762
rect 2573 16710 2625 16762
rect 2641 16742 2655 16762
rect 2655 16742 2689 16762
rect 2689 16742 2693 16762
rect 2641 16710 2693 16742
rect 697 16646 749 16698
rect 765 16668 767 16698
rect 767 16668 801 16698
rect 801 16668 817 16698
rect 765 16646 817 16668
rect 833 16646 885 16698
rect 901 16646 953 16698
rect 969 16668 1003 16698
rect 1003 16668 1021 16698
rect 969 16646 1021 16668
rect 1037 16646 1089 16698
rect 1105 16646 1157 16698
rect 1173 16646 1225 16698
rect 1241 16668 1273 16698
rect 1273 16668 1293 16698
rect 1241 16646 1293 16668
rect 2097 16646 2149 16698
rect 2165 16668 2183 16698
rect 2183 16668 2217 16698
rect 2165 16646 2217 16668
rect 2233 16646 2285 16698
rect 2301 16646 2353 16698
rect 2369 16668 2419 16698
rect 2419 16668 2421 16698
rect 2437 16668 2453 16698
rect 2453 16668 2489 16698
rect 2369 16646 2421 16668
rect 2437 16646 2489 16668
rect 2505 16646 2557 16698
rect 2573 16646 2625 16698
rect 2641 16668 2655 16698
rect 2655 16668 2689 16698
rect 2689 16668 2693 16698
rect 2641 16646 2693 16668
rect 697 16582 749 16634
rect 765 16628 817 16634
rect 765 16594 767 16628
rect 767 16594 801 16628
rect 801 16594 817 16628
rect 765 16582 817 16594
rect 833 16582 885 16634
rect 901 16582 953 16634
rect 969 16628 1021 16634
rect 969 16594 1003 16628
rect 1003 16594 1021 16628
rect 969 16582 1021 16594
rect 1037 16582 1089 16634
rect 1105 16582 1157 16634
rect 1173 16582 1225 16634
rect 1241 16628 1293 16634
rect 1241 16594 1273 16628
rect 1273 16594 1293 16628
rect 1241 16582 1293 16594
rect 2097 16582 2149 16634
rect 2165 16628 2217 16634
rect 2165 16594 2183 16628
rect 2183 16594 2217 16628
rect 2165 16582 2217 16594
rect 2233 16582 2285 16634
rect 2301 16582 2353 16634
rect 2369 16628 2421 16634
rect 2437 16628 2489 16634
rect 2369 16594 2419 16628
rect 2419 16594 2421 16628
rect 2437 16594 2453 16628
rect 2453 16594 2489 16628
rect 2369 16582 2421 16594
rect 2437 16582 2489 16594
rect 2505 16582 2557 16634
rect 2573 16582 2625 16634
rect 2641 16628 2693 16634
rect 2641 16594 2655 16628
rect 2655 16594 2689 16628
rect 2689 16594 2693 16628
rect 2641 16582 2693 16594
rect 697 16518 749 16570
rect 765 16554 817 16570
rect 765 16520 767 16554
rect 767 16520 801 16554
rect 801 16520 817 16554
rect 765 16518 817 16520
rect 833 16518 885 16570
rect 901 16518 953 16570
rect 969 16554 1021 16570
rect 969 16520 1003 16554
rect 1003 16520 1021 16554
rect 969 16518 1021 16520
rect 1037 16518 1089 16570
rect 1105 16518 1157 16570
rect 1173 16518 1225 16570
rect 1241 16554 1293 16570
rect 1241 16520 1273 16554
rect 1273 16520 1293 16554
rect 1241 16518 1293 16520
rect 2097 16518 2149 16570
rect 2165 16554 2217 16570
rect 2165 16520 2183 16554
rect 2183 16520 2217 16554
rect 2165 16518 2217 16520
rect 2233 16518 2285 16570
rect 2301 16518 2353 16570
rect 2369 16554 2421 16570
rect 2437 16554 2489 16570
rect 2369 16520 2419 16554
rect 2419 16520 2421 16554
rect 2437 16520 2453 16554
rect 2453 16520 2489 16554
rect 2369 16518 2421 16520
rect 2437 16518 2489 16520
rect 2505 16518 2557 16570
rect 2573 16518 2625 16570
rect 2641 16554 2693 16570
rect 2641 16520 2655 16554
rect 2655 16520 2689 16554
rect 2689 16520 2693 16554
rect 2641 16518 2693 16520
rect 697 16454 749 16506
rect 765 16480 817 16506
rect 765 16454 767 16480
rect 767 16454 801 16480
rect 801 16454 817 16480
rect 833 16454 885 16506
rect 901 16454 953 16506
rect 969 16480 1021 16506
rect 969 16454 1003 16480
rect 1003 16454 1021 16480
rect 1037 16454 1089 16506
rect 1105 16454 1157 16506
rect 1173 16454 1225 16506
rect 1241 16480 1293 16506
rect 1241 16454 1273 16480
rect 1273 16454 1293 16480
rect 2097 16454 2149 16506
rect 2165 16480 2217 16506
rect 2165 16454 2183 16480
rect 2183 16454 2217 16480
rect 2233 16454 2285 16506
rect 2301 16454 2353 16506
rect 2369 16480 2421 16506
rect 2437 16480 2489 16506
rect 2369 16454 2419 16480
rect 2419 16454 2421 16480
rect 2437 16454 2453 16480
rect 2453 16454 2489 16480
rect 2505 16454 2557 16506
rect 2573 16454 2625 16506
rect 2641 16480 2693 16506
rect 2641 16454 2655 16480
rect 2655 16454 2689 16480
rect 2689 16454 2693 16480
rect 697 16390 749 16442
rect 765 16406 817 16442
rect 765 16390 767 16406
rect 767 16390 801 16406
rect 801 16390 817 16406
rect 833 16390 885 16442
rect 901 16390 953 16442
rect 969 16406 1021 16442
rect 969 16390 1003 16406
rect 1003 16390 1021 16406
rect 1037 16390 1089 16442
rect 1105 16390 1157 16442
rect 1173 16390 1225 16442
rect 1241 16406 1293 16442
rect 1241 16390 1273 16406
rect 1273 16390 1293 16406
rect 697 16326 749 16378
rect 765 16372 767 16378
rect 767 16372 801 16378
rect 801 16372 817 16378
rect 765 16332 817 16372
rect 765 16326 767 16332
rect 767 16326 801 16332
rect 801 16326 817 16332
rect 833 16326 885 16378
rect 901 16326 953 16378
rect 969 16372 1003 16378
rect 1003 16372 1021 16378
rect 969 16332 1021 16372
rect 969 16326 1003 16332
rect 1003 16326 1021 16332
rect 1037 16326 1089 16378
rect 1105 16326 1157 16378
rect 1173 16326 1225 16378
rect 1241 16372 1273 16378
rect 1273 16372 1293 16378
rect 2097 16390 2149 16442
rect 2165 16406 2217 16442
rect 2165 16390 2183 16406
rect 2183 16390 2217 16406
rect 2233 16390 2285 16442
rect 2301 16390 2353 16442
rect 2369 16406 2421 16442
rect 2437 16406 2489 16442
rect 2369 16390 2419 16406
rect 2419 16390 2421 16406
rect 2437 16390 2453 16406
rect 2453 16390 2489 16406
rect 2505 16390 2557 16442
rect 2573 16390 2625 16442
rect 2641 16406 2693 16442
rect 2641 16390 2655 16406
rect 2655 16390 2689 16406
rect 2689 16390 2693 16406
rect 1241 16332 1293 16372
rect 1241 16326 1273 16332
rect 1273 16326 1293 16332
rect 697 16262 749 16314
rect 765 16298 767 16314
rect 767 16298 801 16314
rect 801 16298 817 16314
rect 765 16262 817 16298
rect 833 16262 885 16314
rect 901 16262 953 16314
rect 969 16298 1003 16314
rect 1003 16298 1021 16314
rect 969 16262 1021 16298
rect 1037 16262 1089 16314
rect 1105 16262 1157 16314
rect 1173 16262 1225 16314
rect 1241 16298 1273 16314
rect 1273 16298 1293 16314
rect 2097 16326 2149 16378
rect 2165 16372 2183 16378
rect 2183 16372 2217 16378
rect 2165 16332 2217 16372
rect 2165 16326 2183 16332
rect 2183 16326 2217 16332
rect 2233 16326 2285 16378
rect 2301 16326 2353 16378
rect 2369 16372 2419 16378
rect 2419 16372 2421 16378
rect 2437 16372 2453 16378
rect 2453 16372 2489 16378
rect 2369 16332 2421 16372
rect 2437 16332 2489 16372
rect 2369 16326 2419 16332
rect 2419 16326 2421 16332
rect 2437 16326 2453 16332
rect 2453 16326 2489 16332
rect 2505 16326 2557 16378
rect 2573 16326 2625 16378
rect 2641 16372 2655 16378
rect 2655 16372 2689 16378
rect 2689 16372 2693 16378
rect 2641 16332 2693 16372
rect 2641 16326 2655 16332
rect 2655 16326 2689 16332
rect 2689 16326 2693 16332
rect 1241 16262 1293 16298
rect 2097 16262 2149 16314
rect 2165 16298 2183 16314
rect 2183 16298 2217 16314
rect 2165 16262 2217 16298
rect 2233 16262 2285 16314
rect 2301 16262 2353 16314
rect 2369 16298 2419 16314
rect 2419 16298 2421 16314
rect 2437 16298 2453 16314
rect 2453 16298 2489 16314
rect 2369 16262 2421 16298
rect 2437 16262 2489 16298
rect 2505 16262 2557 16314
rect 2573 16262 2625 16314
rect 2641 16298 2655 16314
rect 2655 16298 2689 16314
rect 2689 16298 2693 16314
rect 2641 16262 2693 16298
rect 697 16198 749 16250
rect 765 16224 767 16250
rect 767 16224 801 16250
rect 801 16224 817 16250
rect 765 16198 817 16224
rect 833 16198 885 16250
rect 901 16198 953 16250
rect 969 16224 1003 16250
rect 1003 16224 1021 16250
rect 969 16198 1021 16224
rect 1037 16198 1089 16250
rect 1105 16198 1157 16250
rect 1173 16198 1225 16250
rect 1241 16224 1273 16250
rect 1273 16224 1293 16250
rect 1241 16198 1293 16224
rect 2097 16198 2149 16250
rect 2165 16224 2183 16250
rect 2183 16224 2217 16250
rect 2165 16198 2217 16224
rect 2233 16198 2285 16250
rect 2301 16198 2353 16250
rect 2369 16224 2419 16250
rect 2419 16224 2421 16250
rect 2437 16224 2453 16250
rect 2453 16224 2489 16250
rect 2369 16198 2421 16224
rect 2437 16198 2489 16224
rect 2505 16198 2557 16250
rect 2573 16198 2625 16250
rect 2641 16224 2655 16250
rect 2655 16224 2689 16250
rect 2689 16224 2693 16250
rect 2641 16198 2693 16224
rect 1501 15624 1553 15633
rect 1569 15624 1621 15633
rect 1636 15624 1688 15633
rect 1703 15624 1755 15633
rect 1770 15624 1822 15633
rect 1837 15624 1889 15633
rect 1501 15590 1525 15624
rect 1525 15590 1553 15624
rect 1569 15590 1600 15624
rect 1600 15590 1621 15624
rect 1636 15590 1674 15624
rect 1674 15590 1688 15624
rect 1703 15590 1708 15624
rect 1708 15590 1748 15624
rect 1748 15590 1755 15624
rect 1770 15590 1782 15624
rect 1782 15590 1822 15624
rect 1837 15590 1856 15624
rect 1856 15590 1889 15624
rect 1501 15581 1553 15590
rect 1569 15581 1621 15590
rect 1636 15581 1688 15590
rect 1703 15581 1755 15590
rect 1770 15581 1822 15590
rect 1837 15581 1889 15590
rect 697 14957 749 15009
rect 765 14997 817 15009
rect 765 14963 767 14997
rect 767 14963 801 14997
rect 801 14963 817 14997
rect 765 14957 817 14963
rect 833 14957 885 15009
rect 901 14957 953 15009
rect 969 14997 1021 15009
rect 969 14963 1003 14997
rect 1003 14963 1021 14997
rect 969 14957 1021 14963
rect 1037 14957 1089 15009
rect 1105 14957 1157 15009
rect 1173 14957 1225 15009
rect 1241 14997 1293 15009
rect 1241 14963 1273 14997
rect 1273 14963 1293 14997
rect 1241 14957 1293 14963
rect 2097 14957 2149 15009
rect 2165 14997 2217 15009
rect 2165 14963 2183 14997
rect 2183 14963 2217 14997
rect 2165 14957 2217 14963
rect 2233 14957 2285 15009
rect 2301 14957 2353 15009
rect 2369 14997 2421 15009
rect 2437 14997 2489 15009
rect 2369 14963 2419 14997
rect 2419 14963 2421 14997
rect 2437 14963 2453 14997
rect 2453 14963 2489 14997
rect 2369 14957 2421 14963
rect 2437 14957 2489 14963
rect 2505 14957 2557 15009
rect 2573 14957 2625 15009
rect 2641 14997 2693 15009
rect 2641 14963 2655 14997
rect 2655 14963 2689 14997
rect 2689 14963 2693 14997
rect 2641 14957 2693 14963
rect 697 14893 749 14945
rect 765 14924 817 14945
rect 765 14893 767 14924
rect 767 14893 801 14924
rect 801 14893 817 14924
rect 833 14893 885 14945
rect 901 14893 953 14945
rect 969 14924 1021 14945
rect 969 14893 1003 14924
rect 1003 14893 1021 14924
rect 1037 14893 1089 14945
rect 1105 14893 1157 14945
rect 1173 14893 1225 14945
rect 1241 14924 1293 14945
rect 1241 14893 1273 14924
rect 1273 14893 1293 14924
rect 2097 14893 2149 14945
rect 2165 14924 2217 14945
rect 2165 14893 2183 14924
rect 2183 14893 2217 14924
rect 2233 14893 2285 14945
rect 2301 14893 2353 14945
rect 2369 14924 2421 14945
rect 2437 14924 2489 14945
rect 2369 14893 2419 14924
rect 2419 14893 2421 14924
rect 2437 14893 2453 14924
rect 2453 14893 2489 14924
rect 2505 14893 2557 14945
rect 2573 14893 2625 14945
rect 2641 14924 2693 14945
rect 2641 14893 2655 14924
rect 2655 14893 2689 14924
rect 2689 14893 2693 14924
rect 697 14829 749 14881
rect 765 14851 817 14881
rect 765 14829 767 14851
rect 767 14829 801 14851
rect 801 14829 817 14851
rect 833 14829 885 14881
rect 901 14829 953 14881
rect 969 14851 1021 14881
rect 969 14829 1003 14851
rect 1003 14829 1021 14851
rect 1037 14829 1089 14881
rect 1105 14829 1157 14881
rect 1173 14829 1225 14881
rect 1241 14851 1293 14881
rect 1241 14829 1273 14851
rect 1273 14829 1293 14851
rect 2097 14829 2149 14881
rect 2165 14851 2217 14881
rect 2165 14829 2183 14851
rect 2183 14829 2217 14851
rect 2233 14829 2285 14881
rect 2301 14829 2353 14881
rect 2369 14851 2421 14881
rect 2437 14851 2489 14881
rect 2369 14829 2419 14851
rect 2419 14829 2421 14851
rect 2437 14829 2453 14851
rect 2453 14829 2489 14851
rect 2505 14829 2557 14881
rect 2573 14829 2625 14881
rect 2641 14851 2693 14881
rect 2641 14829 2655 14851
rect 2655 14829 2689 14851
rect 2689 14829 2693 14851
rect 697 14765 749 14817
rect 765 14778 817 14817
rect 765 14765 767 14778
rect 767 14765 801 14778
rect 801 14765 817 14778
rect 833 14765 885 14817
rect 901 14765 953 14817
rect 969 14778 1021 14817
rect 969 14765 1003 14778
rect 1003 14765 1021 14778
rect 1037 14765 1089 14817
rect 1105 14765 1157 14817
rect 1173 14765 1225 14817
rect 1241 14778 1293 14817
rect 1241 14765 1273 14778
rect 1273 14765 1293 14778
rect 697 14701 749 14753
rect 765 14744 767 14753
rect 767 14744 801 14753
rect 801 14744 817 14753
rect 765 14705 817 14744
rect 765 14701 767 14705
rect 767 14701 801 14705
rect 801 14701 817 14705
rect 833 14701 885 14753
rect 901 14701 953 14753
rect 969 14744 1003 14753
rect 1003 14744 1021 14753
rect 969 14705 1021 14744
rect 969 14701 1003 14705
rect 1003 14701 1021 14705
rect 1037 14701 1089 14753
rect 1105 14701 1157 14753
rect 1173 14701 1225 14753
rect 1241 14744 1273 14753
rect 1273 14744 1293 14753
rect 2097 14765 2149 14817
rect 2165 14778 2217 14817
rect 2165 14765 2183 14778
rect 2183 14765 2217 14778
rect 2233 14765 2285 14817
rect 2301 14765 2353 14817
rect 2369 14778 2421 14817
rect 2437 14778 2489 14817
rect 2369 14765 2419 14778
rect 2419 14765 2421 14778
rect 2437 14765 2453 14778
rect 2453 14765 2489 14778
rect 2505 14765 2557 14817
rect 2573 14765 2625 14817
rect 2641 14778 2693 14817
rect 2641 14765 2655 14778
rect 2655 14765 2689 14778
rect 2689 14765 2693 14778
rect 1241 14705 1293 14744
rect 1241 14701 1273 14705
rect 1273 14701 1293 14705
rect 697 14637 749 14689
rect 765 14671 767 14689
rect 767 14671 801 14689
rect 801 14671 817 14689
rect 765 14637 817 14671
rect 833 14637 885 14689
rect 901 14637 953 14689
rect 969 14671 1003 14689
rect 1003 14671 1021 14689
rect 969 14637 1021 14671
rect 1037 14637 1089 14689
rect 1105 14637 1157 14689
rect 1173 14637 1225 14689
rect 1241 14671 1273 14689
rect 1273 14671 1293 14689
rect 2097 14701 2149 14753
rect 2165 14744 2183 14753
rect 2183 14744 2217 14753
rect 2165 14705 2217 14744
rect 2165 14701 2183 14705
rect 2183 14701 2217 14705
rect 2233 14701 2285 14753
rect 2301 14701 2353 14753
rect 2369 14744 2419 14753
rect 2419 14744 2421 14753
rect 2437 14744 2453 14753
rect 2453 14744 2489 14753
rect 2369 14705 2421 14744
rect 2437 14705 2489 14744
rect 2369 14701 2419 14705
rect 2419 14701 2421 14705
rect 2437 14701 2453 14705
rect 2453 14701 2489 14705
rect 2505 14701 2557 14753
rect 2573 14701 2625 14753
rect 2641 14744 2655 14753
rect 2655 14744 2689 14753
rect 2689 14744 2693 14753
rect 2641 14705 2693 14744
rect 2641 14701 2655 14705
rect 2655 14701 2689 14705
rect 2689 14701 2693 14705
rect 1241 14637 1293 14671
rect 2097 14637 2149 14689
rect 2165 14671 2183 14689
rect 2183 14671 2217 14689
rect 2165 14637 2217 14671
rect 2233 14637 2285 14689
rect 2301 14637 2353 14689
rect 2369 14671 2419 14689
rect 2419 14671 2421 14689
rect 2437 14671 2453 14689
rect 2453 14671 2489 14689
rect 2369 14637 2421 14671
rect 2437 14637 2489 14671
rect 2505 14637 2557 14689
rect 2573 14637 2625 14689
rect 2641 14671 2655 14689
rect 2655 14671 2689 14689
rect 2689 14671 2693 14689
rect 2641 14637 2693 14671
rect 697 14573 749 14625
rect 765 14598 767 14625
rect 767 14598 801 14625
rect 801 14598 817 14625
rect 765 14573 817 14598
rect 833 14573 885 14625
rect 901 14573 953 14625
rect 969 14598 1003 14625
rect 1003 14598 1021 14625
rect 969 14573 1021 14598
rect 1037 14573 1089 14625
rect 1105 14573 1157 14625
rect 1173 14573 1225 14625
rect 1241 14598 1273 14625
rect 1273 14598 1293 14625
rect 1241 14573 1293 14598
rect 2097 14573 2149 14625
rect 2165 14598 2183 14625
rect 2183 14598 2217 14625
rect 2165 14573 2217 14598
rect 2233 14573 2285 14625
rect 2301 14573 2353 14625
rect 2369 14598 2419 14625
rect 2419 14598 2421 14625
rect 2437 14598 2453 14625
rect 2453 14598 2489 14625
rect 2369 14573 2421 14598
rect 2437 14573 2489 14598
rect 2505 14573 2557 14625
rect 2573 14573 2625 14625
rect 2641 14598 2655 14625
rect 2655 14598 2689 14625
rect 2689 14598 2693 14625
rect 2641 14573 2693 14598
rect 697 14509 749 14561
rect 765 14558 817 14561
rect 765 14524 767 14558
rect 767 14524 801 14558
rect 801 14524 817 14558
rect 765 14509 817 14524
rect 833 14509 885 14561
rect 901 14509 953 14561
rect 969 14558 1021 14561
rect 969 14524 1003 14558
rect 1003 14524 1021 14558
rect 969 14509 1021 14524
rect 1037 14509 1089 14561
rect 1105 14509 1157 14561
rect 1173 14509 1225 14561
rect 1241 14558 1293 14561
rect 1241 14524 1273 14558
rect 1273 14524 1293 14558
rect 1241 14509 1293 14524
rect 2097 14509 2149 14561
rect 2165 14558 2217 14561
rect 2165 14524 2183 14558
rect 2183 14524 2217 14558
rect 2165 14509 2217 14524
rect 2233 14509 2285 14561
rect 2301 14509 2353 14561
rect 2369 14558 2421 14561
rect 2437 14558 2489 14561
rect 2369 14524 2419 14558
rect 2419 14524 2421 14558
rect 2437 14524 2453 14558
rect 2453 14524 2489 14558
rect 2369 14509 2421 14524
rect 2437 14509 2489 14524
rect 2505 14509 2557 14561
rect 2573 14509 2625 14561
rect 2641 14558 2693 14561
rect 2641 14524 2655 14558
rect 2655 14524 2689 14558
rect 2689 14524 2693 14558
rect 2641 14509 2693 14524
rect 697 14445 749 14497
rect 765 14484 817 14497
rect 765 14450 767 14484
rect 767 14450 801 14484
rect 801 14450 817 14484
rect 765 14445 817 14450
rect 833 14445 885 14497
rect 901 14445 953 14497
rect 969 14484 1021 14497
rect 969 14450 1003 14484
rect 1003 14450 1021 14484
rect 969 14445 1021 14450
rect 1037 14445 1089 14497
rect 1105 14445 1157 14497
rect 1173 14445 1225 14497
rect 1241 14484 1293 14497
rect 1241 14450 1273 14484
rect 1273 14450 1293 14484
rect 1241 14445 1293 14450
rect 2097 14445 2149 14497
rect 2165 14484 2217 14497
rect 2165 14450 2183 14484
rect 2183 14450 2217 14484
rect 2165 14445 2217 14450
rect 2233 14445 2285 14497
rect 2301 14445 2353 14497
rect 2369 14484 2421 14497
rect 2437 14484 2489 14497
rect 2369 14450 2419 14484
rect 2419 14450 2421 14484
rect 2437 14450 2453 14484
rect 2453 14450 2489 14484
rect 2369 14445 2421 14450
rect 2437 14445 2489 14450
rect 2505 14445 2557 14497
rect 2573 14445 2625 14497
rect 2641 14484 2693 14497
rect 2641 14450 2655 14484
rect 2655 14450 2689 14484
rect 2689 14450 2693 14484
rect 2641 14445 2693 14450
rect 697 14381 749 14433
rect 765 14410 817 14433
rect 765 14381 767 14410
rect 767 14381 801 14410
rect 801 14381 817 14410
rect 833 14381 885 14433
rect 901 14381 953 14433
rect 969 14410 1021 14433
rect 969 14381 1003 14410
rect 1003 14381 1021 14410
rect 1037 14381 1089 14433
rect 1105 14381 1157 14433
rect 1173 14381 1225 14433
rect 1241 14410 1293 14433
rect 1241 14381 1273 14410
rect 1273 14381 1293 14410
rect 2097 14381 2149 14433
rect 2165 14410 2217 14433
rect 2165 14381 2183 14410
rect 2183 14381 2217 14410
rect 2233 14381 2285 14433
rect 2301 14381 2353 14433
rect 2369 14410 2421 14433
rect 2437 14410 2489 14433
rect 2369 14381 2419 14410
rect 2419 14381 2421 14410
rect 2437 14381 2453 14410
rect 2453 14381 2489 14410
rect 2505 14381 2557 14433
rect 2573 14381 2625 14433
rect 2641 14410 2693 14433
rect 2641 14381 2655 14410
rect 2655 14381 2689 14410
rect 2689 14381 2693 14410
rect 697 14317 749 14369
rect 765 14336 817 14369
rect 765 14317 767 14336
rect 767 14317 801 14336
rect 801 14317 817 14336
rect 833 14317 885 14369
rect 901 14317 953 14369
rect 969 14336 1021 14369
rect 969 14317 1003 14336
rect 1003 14317 1021 14336
rect 1037 14317 1089 14369
rect 1105 14317 1157 14369
rect 1173 14317 1225 14369
rect 1241 14336 1293 14369
rect 1241 14317 1273 14336
rect 1273 14317 1293 14336
rect 697 14253 749 14305
rect 765 14302 767 14305
rect 767 14302 801 14305
rect 801 14302 817 14305
rect 765 14262 817 14302
rect 765 14253 767 14262
rect 767 14253 801 14262
rect 801 14253 817 14262
rect 833 14253 885 14305
rect 901 14253 953 14305
rect 969 14302 1003 14305
rect 1003 14302 1021 14305
rect 969 14262 1021 14302
rect 969 14253 1003 14262
rect 1003 14253 1021 14262
rect 1037 14253 1089 14305
rect 1105 14253 1157 14305
rect 1173 14253 1225 14305
rect 1241 14302 1273 14305
rect 1273 14302 1293 14305
rect 2097 14317 2149 14369
rect 2165 14336 2217 14369
rect 2165 14317 2183 14336
rect 2183 14317 2217 14336
rect 2233 14317 2285 14369
rect 2301 14317 2353 14369
rect 2369 14336 2421 14369
rect 2437 14336 2489 14369
rect 2369 14317 2419 14336
rect 2419 14317 2421 14336
rect 2437 14317 2453 14336
rect 2453 14317 2489 14336
rect 2505 14317 2557 14369
rect 2573 14317 2625 14369
rect 2641 14336 2693 14369
rect 2641 14317 2655 14336
rect 2655 14317 2689 14336
rect 2689 14317 2693 14336
rect 1241 14262 1293 14302
rect 1241 14253 1273 14262
rect 1273 14253 1293 14262
rect 697 14189 749 14241
rect 765 14228 767 14241
rect 767 14228 801 14241
rect 801 14228 817 14241
rect 765 14189 817 14228
rect 833 14189 885 14241
rect 901 14189 953 14241
rect 969 14228 1003 14241
rect 1003 14228 1021 14241
rect 969 14189 1021 14228
rect 1037 14189 1089 14241
rect 1105 14189 1157 14241
rect 1173 14189 1225 14241
rect 1241 14228 1273 14241
rect 1273 14228 1293 14241
rect 2097 14253 2149 14305
rect 2165 14302 2183 14305
rect 2183 14302 2217 14305
rect 2165 14262 2217 14302
rect 2165 14253 2183 14262
rect 2183 14253 2217 14262
rect 2233 14253 2285 14305
rect 2301 14253 2353 14305
rect 2369 14302 2419 14305
rect 2419 14302 2421 14305
rect 2437 14302 2453 14305
rect 2453 14302 2489 14305
rect 2369 14262 2421 14302
rect 2437 14262 2489 14302
rect 2369 14253 2419 14262
rect 2419 14253 2421 14262
rect 2437 14253 2453 14262
rect 2453 14253 2489 14262
rect 2505 14253 2557 14305
rect 2573 14253 2625 14305
rect 2641 14302 2655 14305
rect 2655 14302 2689 14305
rect 2689 14302 2693 14305
rect 2641 14262 2693 14302
rect 2641 14253 2655 14262
rect 2655 14253 2689 14262
rect 2689 14253 2693 14262
rect 1241 14189 1293 14228
rect 2097 14189 2149 14241
rect 2165 14228 2183 14241
rect 2183 14228 2217 14241
rect 2165 14189 2217 14228
rect 2233 14189 2285 14241
rect 2301 14189 2353 14241
rect 2369 14228 2419 14241
rect 2419 14228 2421 14241
rect 2437 14228 2453 14241
rect 2453 14228 2489 14241
rect 2369 14189 2421 14228
rect 2437 14189 2489 14228
rect 2505 14189 2557 14241
rect 2573 14189 2625 14241
rect 2641 14228 2655 14241
rect 2655 14228 2689 14241
rect 2689 14228 2693 14241
rect 2641 14189 2693 14228
rect 697 14125 749 14177
rect 765 14154 767 14177
rect 767 14154 801 14177
rect 801 14154 817 14177
rect 765 14125 817 14154
rect 833 14125 885 14177
rect 901 14125 953 14177
rect 969 14154 1003 14177
rect 1003 14154 1021 14177
rect 969 14125 1021 14154
rect 1037 14125 1089 14177
rect 1105 14125 1157 14177
rect 1173 14125 1225 14177
rect 1241 14154 1273 14177
rect 1273 14154 1293 14177
rect 1241 14125 1293 14154
rect 2097 14125 2149 14177
rect 2165 14154 2183 14177
rect 2183 14154 2217 14177
rect 2165 14125 2217 14154
rect 2233 14125 2285 14177
rect 2301 14125 2353 14177
rect 2369 14154 2419 14177
rect 2419 14154 2421 14177
rect 2437 14154 2453 14177
rect 2453 14154 2489 14177
rect 2369 14125 2421 14154
rect 2437 14125 2489 14154
rect 2505 14125 2557 14177
rect 2573 14125 2625 14177
rect 2641 14154 2655 14177
rect 2655 14154 2689 14177
rect 2689 14154 2693 14177
rect 2641 14125 2693 14154
rect 697 14061 749 14113
rect 765 14080 767 14113
rect 767 14080 801 14113
rect 801 14080 817 14113
rect 765 14061 817 14080
rect 833 14061 885 14113
rect 901 14061 953 14113
rect 969 14080 1003 14113
rect 1003 14080 1021 14113
rect 969 14061 1021 14080
rect 1037 14061 1089 14113
rect 1105 14061 1157 14113
rect 1173 14061 1225 14113
rect 1241 14080 1273 14113
rect 1273 14080 1293 14113
rect 1241 14061 1293 14080
rect 2097 14061 2149 14113
rect 2165 14080 2183 14113
rect 2183 14080 2217 14113
rect 2165 14061 2217 14080
rect 2233 14061 2285 14113
rect 2301 14061 2353 14113
rect 2369 14080 2419 14113
rect 2419 14080 2421 14113
rect 2437 14080 2453 14113
rect 2453 14080 2489 14113
rect 2369 14061 2421 14080
rect 2437 14061 2489 14080
rect 2505 14061 2557 14113
rect 2573 14061 2625 14113
rect 2641 14080 2655 14113
rect 2655 14080 2689 14113
rect 2689 14080 2693 14113
rect 2641 14061 2693 14080
rect 1501 13494 1553 13503
rect 1569 13494 1621 13503
rect 1636 13494 1688 13503
rect 1703 13494 1755 13503
rect 1770 13494 1822 13503
rect 1837 13494 1889 13503
rect 1501 13460 1525 13494
rect 1525 13460 1553 13494
rect 1569 13460 1600 13494
rect 1600 13460 1621 13494
rect 1636 13460 1674 13494
rect 1674 13460 1688 13494
rect 1703 13460 1708 13494
rect 1708 13460 1748 13494
rect 1748 13460 1755 13494
rect 1770 13460 1782 13494
rect 1782 13460 1822 13494
rect 1837 13460 1856 13494
rect 1856 13460 1889 13494
rect 1501 13451 1553 13460
rect 1569 13451 1621 13460
rect 1636 13451 1688 13460
rect 1703 13451 1755 13460
rect 1770 13451 1822 13460
rect 1837 13451 1889 13460
rect 697 12855 749 12907
rect 765 12881 817 12907
rect 765 12855 767 12881
rect 767 12855 801 12881
rect 801 12855 817 12881
rect 833 12855 885 12907
rect 901 12855 953 12907
rect 969 12881 1021 12907
rect 969 12855 1003 12881
rect 1003 12855 1021 12881
rect 1037 12855 1089 12907
rect 1105 12855 1157 12907
rect 1173 12855 1225 12907
rect 1241 12881 1293 12907
rect 1241 12855 1273 12881
rect 1273 12855 1293 12881
rect 2097 12855 2149 12907
rect 2165 12881 2217 12907
rect 2165 12855 2183 12881
rect 2183 12855 2217 12881
rect 2233 12855 2285 12907
rect 2301 12855 2353 12907
rect 2369 12881 2421 12907
rect 2437 12881 2489 12907
rect 2369 12855 2419 12881
rect 2419 12855 2421 12881
rect 2437 12855 2453 12881
rect 2453 12855 2489 12881
rect 2505 12855 2557 12907
rect 2573 12855 2625 12907
rect 2641 12881 2693 12907
rect 2641 12855 2655 12881
rect 2655 12855 2689 12881
rect 2689 12855 2693 12881
rect 697 12791 749 12843
rect 765 12808 817 12843
rect 765 12791 767 12808
rect 767 12791 801 12808
rect 801 12791 817 12808
rect 833 12791 885 12843
rect 901 12791 953 12843
rect 969 12808 1021 12843
rect 969 12791 1003 12808
rect 1003 12791 1021 12808
rect 1037 12791 1089 12843
rect 1105 12791 1157 12843
rect 1173 12791 1225 12843
rect 1241 12808 1293 12843
rect 1241 12791 1273 12808
rect 1273 12791 1293 12808
rect 697 12727 749 12779
rect 765 12774 767 12779
rect 767 12774 801 12779
rect 801 12774 817 12779
rect 765 12735 817 12774
rect 765 12727 767 12735
rect 767 12727 801 12735
rect 801 12727 817 12735
rect 833 12727 885 12779
rect 901 12727 953 12779
rect 969 12774 1003 12779
rect 1003 12774 1021 12779
rect 969 12735 1021 12774
rect 969 12727 1003 12735
rect 1003 12727 1021 12735
rect 1037 12727 1089 12779
rect 1105 12727 1157 12779
rect 1173 12727 1225 12779
rect 1241 12774 1273 12779
rect 1273 12774 1293 12779
rect 2097 12791 2149 12843
rect 2165 12808 2217 12843
rect 2165 12791 2183 12808
rect 2183 12791 2217 12808
rect 2233 12791 2285 12843
rect 2301 12791 2353 12843
rect 2369 12808 2421 12843
rect 2437 12808 2489 12843
rect 2369 12791 2419 12808
rect 2419 12791 2421 12808
rect 2437 12791 2453 12808
rect 2453 12791 2489 12808
rect 2505 12791 2557 12843
rect 2573 12791 2625 12843
rect 2641 12808 2693 12843
rect 2641 12791 2655 12808
rect 2655 12791 2689 12808
rect 2689 12791 2693 12808
rect 1241 12735 1293 12774
rect 1241 12727 1273 12735
rect 1273 12727 1293 12735
rect 697 12663 749 12715
rect 765 12701 767 12715
rect 767 12701 801 12715
rect 801 12701 817 12715
rect 765 12663 817 12701
rect 833 12663 885 12715
rect 901 12663 953 12715
rect 969 12701 1003 12715
rect 1003 12701 1021 12715
rect 969 12663 1021 12701
rect 1037 12663 1089 12715
rect 1105 12663 1157 12715
rect 1173 12663 1225 12715
rect 1241 12701 1273 12715
rect 1273 12701 1293 12715
rect 2097 12727 2149 12779
rect 2165 12774 2183 12779
rect 2183 12774 2217 12779
rect 2165 12735 2217 12774
rect 2165 12727 2183 12735
rect 2183 12727 2217 12735
rect 2233 12727 2285 12779
rect 2301 12727 2353 12779
rect 2369 12774 2419 12779
rect 2419 12774 2421 12779
rect 2437 12774 2453 12779
rect 2453 12774 2489 12779
rect 2369 12735 2421 12774
rect 2437 12735 2489 12774
rect 2369 12727 2419 12735
rect 2419 12727 2421 12735
rect 2437 12727 2453 12735
rect 2453 12727 2489 12735
rect 2505 12727 2557 12779
rect 2573 12727 2625 12779
rect 2641 12774 2655 12779
rect 2655 12774 2689 12779
rect 2689 12774 2693 12779
rect 2641 12735 2693 12774
rect 2641 12727 2655 12735
rect 2655 12727 2689 12735
rect 2689 12727 2693 12735
rect 1241 12663 1293 12701
rect 2097 12663 2149 12715
rect 2165 12701 2183 12715
rect 2183 12701 2217 12715
rect 2165 12663 2217 12701
rect 2233 12663 2285 12715
rect 2301 12663 2353 12715
rect 2369 12701 2419 12715
rect 2419 12701 2421 12715
rect 2437 12701 2453 12715
rect 2453 12701 2489 12715
rect 2369 12663 2421 12701
rect 2437 12663 2489 12701
rect 2505 12663 2557 12715
rect 2573 12663 2625 12715
rect 2641 12701 2655 12715
rect 2655 12701 2689 12715
rect 2689 12701 2693 12715
rect 2641 12663 2693 12701
rect 697 12599 749 12651
rect 765 12628 767 12651
rect 767 12628 801 12651
rect 801 12628 817 12651
rect 765 12599 817 12628
rect 833 12599 885 12651
rect 901 12599 953 12651
rect 969 12628 1003 12651
rect 1003 12628 1021 12651
rect 969 12599 1021 12628
rect 1037 12599 1089 12651
rect 1105 12599 1157 12651
rect 1173 12599 1225 12651
rect 1241 12628 1273 12651
rect 1273 12628 1293 12651
rect 1241 12599 1293 12628
rect 2097 12599 2149 12651
rect 2165 12628 2183 12651
rect 2183 12628 2217 12651
rect 2165 12599 2217 12628
rect 2233 12599 2285 12651
rect 2301 12599 2353 12651
rect 2369 12628 2419 12651
rect 2419 12628 2421 12651
rect 2437 12628 2453 12651
rect 2453 12628 2489 12651
rect 2369 12599 2421 12628
rect 2437 12599 2489 12628
rect 2505 12599 2557 12651
rect 2573 12599 2625 12651
rect 2641 12628 2655 12651
rect 2655 12628 2689 12651
rect 2689 12628 2693 12651
rect 2641 12599 2693 12628
rect 697 12535 749 12587
rect 765 12555 767 12587
rect 767 12555 801 12587
rect 801 12555 817 12587
rect 765 12535 817 12555
rect 833 12535 885 12587
rect 901 12535 953 12587
rect 969 12555 1003 12587
rect 1003 12555 1021 12587
rect 969 12535 1021 12555
rect 1037 12535 1089 12587
rect 1105 12535 1157 12587
rect 1173 12535 1225 12587
rect 1241 12555 1273 12587
rect 1273 12555 1293 12587
rect 1241 12535 1293 12555
rect 2097 12535 2149 12587
rect 2165 12555 2183 12587
rect 2183 12555 2217 12587
rect 2165 12535 2217 12555
rect 2233 12535 2285 12587
rect 2301 12535 2353 12587
rect 2369 12555 2419 12587
rect 2419 12555 2421 12587
rect 2437 12555 2453 12587
rect 2453 12555 2489 12587
rect 2369 12535 2421 12555
rect 2437 12535 2489 12555
rect 2505 12535 2557 12587
rect 2573 12535 2625 12587
rect 2641 12555 2655 12587
rect 2655 12555 2689 12587
rect 2689 12555 2693 12587
rect 2641 12535 2693 12555
rect 697 12471 749 12523
rect 765 12516 817 12523
rect 765 12482 767 12516
rect 767 12482 801 12516
rect 801 12482 817 12516
rect 765 12471 817 12482
rect 833 12471 885 12523
rect 901 12471 953 12523
rect 969 12516 1021 12523
rect 969 12482 1003 12516
rect 1003 12482 1021 12516
rect 969 12471 1021 12482
rect 1037 12471 1089 12523
rect 1105 12471 1157 12523
rect 1173 12471 1225 12523
rect 1241 12516 1293 12523
rect 1241 12482 1273 12516
rect 1273 12482 1293 12516
rect 1241 12471 1293 12482
rect 2097 12471 2149 12523
rect 2165 12516 2217 12523
rect 2165 12482 2183 12516
rect 2183 12482 2217 12516
rect 2165 12471 2217 12482
rect 2233 12471 2285 12523
rect 2301 12471 2353 12523
rect 2369 12516 2421 12523
rect 2437 12516 2489 12523
rect 2369 12482 2419 12516
rect 2419 12482 2421 12516
rect 2437 12482 2453 12516
rect 2453 12482 2489 12516
rect 2369 12471 2421 12482
rect 2437 12471 2489 12482
rect 2505 12471 2557 12523
rect 2573 12471 2625 12523
rect 2641 12516 2693 12523
rect 2641 12482 2655 12516
rect 2655 12482 2689 12516
rect 2689 12482 2693 12516
rect 2641 12471 2693 12482
rect 697 12407 749 12459
rect 765 12442 817 12459
rect 765 12408 767 12442
rect 767 12408 801 12442
rect 801 12408 817 12442
rect 765 12407 817 12408
rect 833 12407 885 12459
rect 901 12407 953 12459
rect 969 12442 1021 12459
rect 969 12408 1003 12442
rect 1003 12408 1021 12442
rect 969 12407 1021 12408
rect 1037 12407 1089 12459
rect 1105 12407 1157 12459
rect 1173 12407 1225 12459
rect 1241 12442 1293 12459
rect 1241 12408 1273 12442
rect 1273 12408 1293 12442
rect 1241 12407 1293 12408
rect 2097 12407 2149 12459
rect 2165 12442 2217 12459
rect 2165 12408 2183 12442
rect 2183 12408 2217 12442
rect 2165 12407 2217 12408
rect 2233 12407 2285 12459
rect 2301 12407 2353 12459
rect 2369 12442 2421 12459
rect 2437 12442 2489 12459
rect 2369 12408 2419 12442
rect 2419 12408 2421 12442
rect 2437 12408 2453 12442
rect 2453 12408 2489 12442
rect 2369 12407 2421 12408
rect 2437 12407 2489 12408
rect 2505 12407 2557 12459
rect 2573 12407 2625 12459
rect 2641 12442 2693 12459
rect 2641 12408 2655 12442
rect 2655 12408 2689 12442
rect 2689 12408 2693 12442
rect 2641 12407 2693 12408
rect 697 12343 749 12395
rect 765 12368 817 12395
rect 765 12343 767 12368
rect 767 12343 801 12368
rect 801 12343 817 12368
rect 833 12343 885 12395
rect 901 12343 953 12395
rect 969 12368 1021 12395
rect 969 12343 1003 12368
rect 1003 12343 1021 12368
rect 1037 12343 1089 12395
rect 1105 12343 1157 12395
rect 1173 12343 1225 12395
rect 1241 12368 1293 12395
rect 1241 12343 1273 12368
rect 1273 12343 1293 12368
rect 2097 12343 2149 12395
rect 2165 12368 2217 12395
rect 2165 12343 2183 12368
rect 2183 12343 2217 12368
rect 2233 12343 2285 12395
rect 2301 12343 2353 12395
rect 2369 12368 2421 12395
rect 2437 12368 2489 12395
rect 2369 12343 2419 12368
rect 2419 12343 2421 12368
rect 2437 12343 2453 12368
rect 2453 12343 2489 12368
rect 2505 12343 2557 12395
rect 2573 12343 2625 12395
rect 2641 12368 2693 12395
rect 2641 12343 2655 12368
rect 2655 12343 2689 12368
rect 2689 12343 2693 12368
rect 697 12279 749 12331
rect 765 12294 817 12331
rect 765 12279 767 12294
rect 767 12279 801 12294
rect 801 12279 817 12294
rect 833 12279 885 12331
rect 901 12279 953 12331
rect 969 12294 1021 12331
rect 969 12279 1003 12294
rect 1003 12279 1021 12294
rect 1037 12279 1089 12331
rect 1105 12279 1157 12331
rect 1173 12279 1225 12331
rect 1241 12294 1293 12331
rect 1241 12279 1273 12294
rect 1273 12279 1293 12294
rect 697 12215 749 12267
rect 765 12260 767 12267
rect 767 12260 801 12267
rect 801 12260 817 12267
rect 765 12220 817 12260
rect 765 12215 767 12220
rect 767 12215 801 12220
rect 801 12215 817 12220
rect 833 12215 885 12267
rect 901 12215 953 12267
rect 969 12260 1003 12267
rect 1003 12260 1021 12267
rect 969 12220 1021 12260
rect 969 12215 1003 12220
rect 1003 12215 1021 12220
rect 1037 12215 1089 12267
rect 1105 12215 1157 12267
rect 1173 12215 1225 12267
rect 1241 12260 1273 12267
rect 1273 12260 1293 12267
rect 2097 12279 2149 12331
rect 2165 12294 2217 12331
rect 2165 12279 2183 12294
rect 2183 12279 2217 12294
rect 2233 12279 2285 12331
rect 2301 12279 2353 12331
rect 2369 12294 2421 12331
rect 2437 12294 2489 12331
rect 2369 12279 2419 12294
rect 2419 12279 2421 12294
rect 2437 12279 2453 12294
rect 2453 12279 2489 12294
rect 2505 12279 2557 12331
rect 2573 12279 2625 12331
rect 2641 12294 2693 12331
rect 2641 12279 2655 12294
rect 2655 12279 2689 12294
rect 2689 12279 2693 12294
rect 1241 12220 1293 12260
rect 1241 12215 1273 12220
rect 1273 12215 1293 12220
rect 697 12151 749 12203
rect 765 12186 767 12203
rect 767 12186 801 12203
rect 801 12186 817 12203
rect 765 12151 817 12186
rect 833 12151 885 12203
rect 901 12151 953 12203
rect 969 12186 1003 12203
rect 1003 12186 1021 12203
rect 969 12151 1021 12186
rect 1037 12151 1089 12203
rect 1105 12151 1157 12203
rect 1173 12151 1225 12203
rect 1241 12186 1273 12203
rect 1273 12186 1293 12203
rect 2097 12215 2149 12267
rect 2165 12260 2183 12267
rect 2183 12260 2217 12267
rect 2165 12220 2217 12260
rect 2165 12215 2183 12220
rect 2183 12215 2217 12220
rect 2233 12215 2285 12267
rect 2301 12215 2353 12267
rect 2369 12260 2419 12267
rect 2419 12260 2421 12267
rect 2437 12260 2453 12267
rect 2453 12260 2489 12267
rect 2369 12220 2421 12260
rect 2437 12220 2489 12260
rect 2369 12215 2419 12220
rect 2419 12215 2421 12220
rect 2437 12215 2453 12220
rect 2453 12215 2489 12220
rect 2505 12215 2557 12267
rect 2573 12215 2625 12267
rect 2641 12260 2655 12267
rect 2655 12260 2689 12267
rect 2689 12260 2693 12267
rect 2641 12220 2693 12260
rect 2641 12215 2655 12220
rect 2655 12215 2689 12220
rect 2689 12215 2693 12220
rect 1241 12151 1293 12186
rect 2097 12151 2149 12203
rect 2165 12186 2183 12203
rect 2183 12186 2217 12203
rect 2165 12151 2217 12186
rect 2233 12151 2285 12203
rect 2301 12151 2353 12203
rect 2369 12186 2419 12203
rect 2419 12186 2421 12203
rect 2437 12186 2453 12203
rect 2453 12186 2489 12203
rect 2369 12151 2421 12186
rect 2437 12151 2489 12186
rect 2505 12151 2557 12203
rect 2573 12151 2625 12203
rect 2641 12186 2655 12203
rect 2655 12186 2689 12203
rect 2689 12186 2693 12203
rect 2641 12151 2693 12186
rect 697 12087 749 12139
rect 765 12112 767 12139
rect 767 12112 801 12139
rect 801 12112 817 12139
rect 765 12087 817 12112
rect 833 12087 885 12139
rect 901 12087 953 12139
rect 969 12112 1003 12139
rect 1003 12112 1021 12139
rect 969 12087 1021 12112
rect 1037 12087 1089 12139
rect 1105 12087 1157 12139
rect 1173 12087 1225 12139
rect 1241 12112 1273 12139
rect 1273 12112 1293 12139
rect 1241 12087 1293 12112
rect 2097 12087 2149 12139
rect 2165 12112 2183 12139
rect 2183 12112 2217 12139
rect 2165 12087 2217 12112
rect 2233 12087 2285 12139
rect 2301 12087 2353 12139
rect 2369 12112 2419 12139
rect 2419 12112 2421 12139
rect 2437 12112 2453 12139
rect 2453 12112 2489 12139
rect 2369 12087 2421 12112
rect 2437 12087 2489 12112
rect 2505 12087 2557 12139
rect 2573 12087 2625 12139
rect 2641 12112 2655 12139
rect 2655 12112 2689 12139
rect 2689 12112 2693 12139
rect 2641 12087 2693 12112
rect 697 12023 749 12075
rect 765 12072 817 12075
rect 765 12038 767 12072
rect 767 12038 801 12072
rect 801 12038 817 12072
rect 765 12023 817 12038
rect 833 12023 885 12075
rect 901 12023 953 12075
rect 969 12072 1021 12075
rect 969 12038 1003 12072
rect 1003 12038 1021 12072
rect 969 12023 1021 12038
rect 1037 12023 1089 12075
rect 1105 12023 1157 12075
rect 1173 12023 1225 12075
rect 1241 12072 1293 12075
rect 1241 12038 1273 12072
rect 1273 12038 1293 12072
rect 1241 12023 1293 12038
rect 2097 12023 2149 12075
rect 2165 12072 2217 12075
rect 2165 12038 2183 12072
rect 2183 12038 2217 12072
rect 2165 12023 2217 12038
rect 2233 12023 2285 12075
rect 2301 12023 2353 12075
rect 2369 12072 2421 12075
rect 2437 12072 2489 12075
rect 2369 12038 2419 12072
rect 2419 12038 2421 12072
rect 2437 12038 2453 12072
rect 2453 12038 2489 12072
rect 2369 12023 2421 12038
rect 2437 12023 2489 12038
rect 2505 12023 2557 12075
rect 2573 12023 2625 12075
rect 2641 12072 2693 12075
rect 2641 12038 2655 12072
rect 2655 12038 2689 12072
rect 2689 12038 2693 12072
rect 2641 12023 2693 12038
rect 697 11959 749 12011
rect 765 11998 817 12011
rect 765 11964 767 11998
rect 767 11964 801 11998
rect 801 11964 817 11998
rect 765 11959 817 11964
rect 833 11959 885 12011
rect 901 11959 953 12011
rect 969 11998 1021 12011
rect 969 11964 1003 11998
rect 1003 11964 1021 11998
rect 969 11959 1021 11964
rect 1037 11959 1089 12011
rect 1105 11959 1157 12011
rect 1173 11959 1225 12011
rect 1241 11998 1293 12011
rect 1241 11964 1273 11998
rect 1273 11964 1293 11998
rect 1241 11959 1293 11964
rect 2097 11959 2149 12011
rect 2165 11998 2217 12011
rect 2165 11964 2183 11998
rect 2183 11964 2217 11998
rect 2165 11959 2217 11964
rect 2233 11959 2285 12011
rect 2301 11959 2353 12011
rect 2369 11998 2421 12011
rect 2437 11998 2489 12011
rect 2369 11964 2419 11998
rect 2419 11964 2421 11998
rect 2437 11964 2453 11998
rect 2453 11964 2489 11998
rect 2369 11959 2421 11964
rect 2437 11959 2489 11964
rect 2505 11959 2557 12011
rect 2573 11959 2625 12011
rect 2641 11998 2693 12011
rect 2641 11964 2655 11998
rect 2655 11964 2689 11998
rect 2689 11964 2693 11998
rect 2641 11959 2693 11964
rect 1501 11364 1553 11373
rect 1569 11364 1621 11373
rect 1636 11364 1688 11373
rect 1703 11364 1755 11373
rect 1770 11364 1822 11373
rect 1837 11364 1889 11373
rect 1501 11330 1525 11364
rect 1525 11330 1553 11364
rect 1569 11330 1600 11364
rect 1600 11330 1621 11364
rect 1636 11330 1674 11364
rect 1674 11330 1688 11364
rect 1703 11330 1708 11364
rect 1708 11330 1748 11364
rect 1748 11330 1755 11364
rect 1770 11330 1782 11364
rect 1782 11330 1822 11364
rect 1837 11330 1856 11364
rect 1856 11330 1889 11364
rect 1501 11321 1553 11330
rect 1569 11321 1621 11330
rect 1636 11321 1688 11330
rect 1703 11321 1755 11330
rect 1770 11321 1822 11330
rect 1837 11321 1889 11330
rect 697 10761 749 10813
rect 765 10810 817 10813
rect 765 10776 767 10810
rect 767 10776 801 10810
rect 801 10776 817 10810
rect 765 10761 817 10776
rect 833 10761 885 10813
rect 901 10761 953 10813
rect 969 10810 1021 10813
rect 969 10776 1003 10810
rect 1003 10776 1021 10810
rect 969 10761 1021 10776
rect 1037 10761 1089 10813
rect 1105 10761 1157 10813
rect 1173 10761 1225 10813
rect 1241 10810 1293 10813
rect 1241 10776 1273 10810
rect 1273 10776 1293 10810
rect 1241 10761 1293 10776
rect 2097 10761 2149 10813
rect 2165 10810 2217 10813
rect 2165 10776 2183 10810
rect 2183 10776 2217 10810
rect 2165 10761 2217 10776
rect 2233 10761 2285 10813
rect 2301 10761 2353 10813
rect 2369 10810 2421 10813
rect 2437 10810 2489 10813
rect 2369 10776 2419 10810
rect 2419 10776 2421 10810
rect 2437 10776 2453 10810
rect 2453 10776 2489 10810
rect 2369 10761 2421 10776
rect 2437 10761 2489 10776
rect 2505 10761 2557 10813
rect 2573 10761 2625 10813
rect 2641 10810 2693 10813
rect 2641 10776 2655 10810
rect 2655 10776 2689 10810
rect 2689 10776 2693 10810
rect 2641 10761 2693 10776
rect 697 10697 749 10749
rect 765 10737 817 10749
rect 765 10703 767 10737
rect 767 10703 801 10737
rect 801 10703 817 10737
rect 765 10697 817 10703
rect 833 10697 885 10749
rect 901 10697 953 10749
rect 969 10737 1021 10749
rect 969 10703 1003 10737
rect 1003 10703 1021 10737
rect 969 10697 1021 10703
rect 1037 10697 1089 10749
rect 1105 10697 1157 10749
rect 1173 10697 1225 10749
rect 1241 10737 1293 10749
rect 1241 10703 1273 10737
rect 1273 10703 1293 10737
rect 1241 10697 1293 10703
rect 2097 10697 2149 10749
rect 2165 10737 2217 10749
rect 2165 10703 2183 10737
rect 2183 10703 2217 10737
rect 2165 10697 2217 10703
rect 2233 10697 2285 10749
rect 2301 10697 2353 10749
rect 2369 10737 2421 10749
rect 2437 10737 2489 10749
rect 2369 10703 2419 10737
rect 2419 10703 2421 10737
rect 2437 10703 2453 10737
rect 2453 10703 2489 10737
rect 2369 10697 2421 10703
rect 2437 10697 2489 10703
rect 2505 10697 2557 10749
rect 2573 10697 2625 10749
rect 2641 10737 2693 10749
rect 2641 10703 2655 10737
rect 2655 10703 2689 10737
rect 2689 10703 2693 10737
rect 2641 10697 2693 10703
rect 697 10633 749 10685
rect 765 10664 817 10685
rect 765 10633 767 10664
rect 767 10633 801 10664
rect 801 10633 817 10664
rect 833 10633 885 10685
rect 901 10633 953 10685
rect 969 10664 1021 10685
rect 969 10633 1003 10664
rect 1003 10633 1021 10664
rect 1037 10633 1089 10685
rect 1105 10633 1157 10685
rect 1173 10633 1225 10685
rect 1241 10664 1293 10685
rect 1241 10633 1273 10664
rect 1273 10633 1293 10664
rect 2097 10633 2149 10685
rect 2165 10664 2217 10685
rect 2165 10633 2183 10664
rect 2183 10633 2217 10664
rect 2233 10633 2285 10685
rect 2301 10633 2353 10685
rect 2369 10664 2421 10685
rect 2437 10664 2489 10685
rect 2369 10633 2419 10664
rect 2419 10633 2421 10664
rect 2437 10633 2453 10664
rect 2453 10633 2489 10664
rect 2505 10633 2557 10685
rect 2573 10633 2625 10685
rect 2641 10664 2693 10685
rect 2641 10633 2655 10664
rect 2655 10633 2689 10664
rect 2689 10633 2693 10664
rect 697 10569 749 10621
rect 765 10591 817 10621
rect 765 10569 767 10591
rect 767 10569 801 10591
rect 801 10569 817 10591
rect 833 10569 885 10621
rect 901 10569 953 10621
rect 969 10591 1021 10621
rect 969 10569 1003 10591
rect 1003 10569 1021 10591
rect 1037 10569 1089 10621
rect 1105 10569 1157 10621
rect 1173 10569 1225 10621
rect 1241 10591 1293 10621
rect 1241 10569 1273 10591
rect 1273 10569 1293 10591
rect 2097 10569 2149 10621
rect 2165 10591 2217 10621
rect 2165 10569 2183 10591
rect 2183 10569 2217 10591
rect 2233 10569 2285 10621
rect 2301 10569 2353 10621
rect 2369 10591 2421 10621
rect 2437 10591 2489 10621
rect 2369 10569 2419 10591
rect 2419 10569 2421 10591
rect 2437 10569 2453 10591
rect 2453 10569 2489 10591
rect 2505 10569 2557 10621
rect 2573 10569 2625 10621
rect 2641 10591 2693 10621
rect 2641 10569 2655 10591
rect 2655 10569 2689 10591
rect 2689 10569 2693 10591
rect 697 10505 749 10557
rect 765 10518 817 10557
rect 765 10505 767 10518
rect 767 10505 801 10518
rect 801 10505 817 10518
rect 833 10505 885 10557
rect 901 10505 953 10557
rect 969 10518 1021 10557
rect 969 10505 1003 10518
rect 1003 10505 1021 10518
rect 1037 10505 1089 10557
rect 1105 10505 1157 10557
rect 1173 10505 1225 10557
rect 1241 10518 1293 10557
rect 1241 10505 1273 10518
rect 1273 10505 1293 10518
rect 697 10441 749 10493
rect 765 10484 767 10493
rect 767 10484 801 10493
rect 801 10484 817 10493
rect 765 10445 817 10484
rect 765 10441 767 10445
rect 767 10441 801 10445
rect 801 10441 817 10445
rect 833 10441 885 10493
rect 901 10441 953 10493
rect 969 10484 1003 10493
rect 1003 10484 1021 10493
rect 969 10445 1021 10484
rect 969 10441 1003 10445
rect 1003 10441 1021 10445
rect 1037 10441 1089 10493
rect 1105 10441 1157 10493
rect 1173 10441 1225 10493
rect 1241 10484 1273 10493
rect 1273 10484 1293 10493
rect 2097 10505 2149 10557
rect 2165 10518 2217 10557
rect 2165 10505 2183 10518
rect 2183 10505 2217 10518
rect 2233 10505 2285 10557
rect 2301 10505 2353 10557
rect 2369 10518 2421 10557
rect 2437 10518 2489 10557
rect 2369 10505 2419 10518
rect 2419 10505 2421 10518
rect 2437 10505 2453 10518
rect 2453 10505 2489 10518
rect 2505 10505 2557 10557
rect 2573 10505 2625 10557
rect 2641 10518 2693 10557
rect 2641 10505 2655 10518
rect 2655 10505 2689 10518
rect 2689 10505 2693 10518
rect 1241 10445 1293 10484
rect 1241 10441 1273 10445
rect 1273 10441 1293 10445
rect 697 10377 749 10429
rect 765 10411 767 10429
rect 767 10411 801 10429
rect 801 10411 817 10429
rect 765 10377 817 10411
rect 833 10377 885 10429
rect 901 10377 953 10429
rect 969 10411 1003 10429
rect 1003 10411 1021 10429
rect 969 10377 1021 10411
rect 1037 10377 1089 10429
rect 1105 10377 1157 10429
rect 1173 10377 1225 10429
rect 1241 10411 1273 10429
rect 1273 10411 1293 10429
rect 2097 10441 2149 10493
rect 2165 10484 2183 10493
rect 2183 10484 2217 10493
rect 2165 10445 2217 10484
rect 2165 10441 2183 10445
rect 2183 10441 2217 10445
rect 2233 10441 2285 10493
rect 2301 10441 2353 10493
rect 2369 10484 2419 10493
rect 2419 10484 2421 10493
rect 2437 10484 2453 10493
rect 2453 10484 2489 10493
rect 2369 10445 2421 10484
rect 2437 10445 2489 10484
rect 2369 10441 2419 10445
rect 2419 10441 2421 10445
rect 2437 10441 2453 10445
rect 2453 10441 2489 10445
rect 2505 10441 2557 10493
rect 2573 10441 2625 10493
rect 2641 10484 2655 10493
rect 2655 10484 2689 10493
rect 2689 10484 2693 10493
rect 2641 10445 2693 10484
rect 2641 10441 2655 10445
rect 2655 10441 2689 10445
rect 2689 10441 2693 10445
rect 1241 10377 1293 10411
rect 2097 10377 2149 10429
rect 2165 10411 2183 10429
rect 2183 10411 2217 10429
rect 2165 10377 2217 10411
rect 2233 10377 2285 10429
rect 2301 10377 2353 10429
rect 2369 10411 2419 10429
rect 2419 10411 2421 10429
rect 2437 10411 2453 10429
rect 2453 10411 2489 10429
rect 2369 10377 2421 10411
rect 2437 10377 2489 10411
rect 2505 10377 2557 10429
rect 2573 10377 2625 10429
rect 2641 10411 2655 10429
rect 2655 10411 2689 10429
rect 2689 10411 2693 10429
rect 2641 10377 2693 10411
rect 697 10313 749 10365
rect 765 10338 767 10365
rect 767 10338 801 10365
rect 801 10338 817 10365
rect 765 10313 817 10338
rect 833 10313 885 10365
rect 901 10313 953 10365
rect 969 10338 1003 10365
rect 1003 10338 1021 10365
rect 969 10313 1021 10338
rect 1037 10313 1089 10365
rect 1105 10313 1157 10365
rect 1173 10313 1225 10365
rect 1241 10338 1273 10365
rect 1273 10338 1293 10365
rect 1241 10313 1293 10338
rect 2097 10313 2149 10365
rect 2165 10338 2183 10365
rect 2183 10338 2217 10365
rect 2165 10313 2217 10338
rect 2233 10313 2285 10365
rect 2301 10313 2353 10365
rect 2369 10338 2419 10365
rect 2419 10338 2421 10365
rect 2437 10338 2453 10365
rect 2453 10338 2489 10365
rect 2369 10313 2421 10338
rect 2437 10313 2489 10338
rect 2505 10313 2557 10365
rect 2573 10313 2625 10365
rect 2641 10338 2655 10365
rect 2655 10338 2689 10365
rect 2689 10338 2693 10365
rect 2641 10313 2693 10338
rect 697 10249 749 10301
rect 765 10298 817 10301
rect 765 10264 767 10298
rect 767 10264 801 10298
rect 801 10264 817 10298
rect 765 10249 817 10264
rect 833 10249 885 10301
rect 901 10249 953 10301
rect 969 10298 1021 10301
rect 969 10264 1003 10298
rect 1003 10264 1021 10298
rect 969 10249 1021 10264
rect 1037 10249 1089 10301
rect 1105 10249 1157 10301
rect 1173 10249 1225 10301
rect 1241 10298 1293 10301
rect 1241 10264 1273 10298
rect 1273 10264 1293 10298
rect 1241 10249 1293 10264
rect 2097 10249 2149 10301
rect 2165 10298 2217 10301
rect 2165 10264 2183 10298
rect 2183 10264 2217 10298
rect 2165 10249 2217 10264
rect 2233 10249 2285 10301
rect 2301 10249 2353 10301
rect 2369 10298 2421 10301
rect 2437 10298 2489 10301
rect 2369 10264 2419 10298
rect 2419 10264 2421 10298
rect 2437 10264 2453 10298
rect 2453 10264 2489 10298
rect 2369 10249 2421 10264
rect 2437 10249 2489 10264
rect 2505 10249 2557 10301
rect 2573 10249 2625 10301
rect 2641 10298 2693 10301
rect 2641 10264 2655 10298
rect 2655 10264 2689 10298
rect 2689 10264 2693 10298
rect 2641 10249 2693 10264
rect 697 10185 749 10237
rect 765 10224 817 10237
rect 765 10190 767 10224
rect 767 10190 801 10224
rect 801 10190 817 10224
rect 765 10185 817 10190
rect 833 10185 885 10237
rect 901 10185 953 10237
rect 969 10224 1021 10237
rect 969 10190 1003 10224
rect 1003 10190 1021 10224
rect 969 10185 1021 10190
rect 1037 10185 1089 10237
rect 1105 10185 1157 10237
rect 1173 10185 1225 10237
rect 1241 10224 1293 10237
rect 1241 10190 1273 10224
rect 1273 10190 1293 10224
rect 1241 10185 1293 10190
rect 2097 10185 2149 10237
rect 2165 10224 2217 10237
rect 2165 10190 2183 10224
rect 2183 10190 2217 10224
rect 2165 10185 2217 10190
rect 2233 10185 2285 10237
rect 2301 10185 2353 10237
rect 2369 10224 2421 10237
rect 2437 10224 2489 10237
rect 2369 10190 2419 10224
rect 2419 10190 2421 10224
rect 2437 10190 2453 10224
rect 2453 10190 2489 10224
rect 2369 10185 2421 10190
rect 2437 10185 2489 10190
rect 2505 10185 2557 10237
rect 2573 10185 2625 10237
rect 2641 10224 2693 10237
rect 2641 10190 2655 10224
rect 2655 10190 2689 10224
rect 2689 10190 2693 10224
rect 2641 10185 2693 10190
rect 697 10121 749 10173
rect 765 10150 817 10173
rect 765 10121 767 10150
rect 767 10121 801 10150
rect 801 10121 817 10150
rect 833 10121 885 10173
rect 901 10121 953 10173
rect 969 10150 1021 10173
rect 969 10121 1003 10150
rect 1003 10121 1021 10150
rect 1037 10121 1089 10173
rect 1105 10121 1157 10173
rect 1173 10121 1225 10173
rect 1241 10150 1293 10173
rect 1241 10121 1273 10150
rect 1273 10121 1293 10150
rect 2097 10121 2149 10173
rect 2165 10150 2217 10173
rect 2165 10121 2183 10150
rect 2183 10121 2217 10150
rect 2233 10121 2285 10173
rect 2301 10121 2353 10173
rect 2369 10150 2421 10173
rect 2437 10150 2489 10173
rect 2369 10121 2419 10150
rect 2419 10121 2421 10150
rect 2437 10121 2453 10150
rect 2453 10121 2489 10150
rect 2505 10121 2557 10173
rect 2573 10121 2625 10173
rect 2641 10150 2693 10173
rect 2641 10121 2655 10150
rect 2655 10121 2689 10150
rect 2689 10121 2693 10150
rect 697 10057 749 10109
rect 765 10076 817 10109
rect 765 10057 767 10076
rect 767 10057 801 10076
rect 801 10057 817 10076
rect 833 10057 885 10109
rect 901 10057 953 10109
rect 969 10076 1021 10109
rect 969 10057 1003 10076
rect 1003 10057 1021 10076
rect 1037 10057 1089 10109
rect 1105 10057 1157 10109
rect 1173 10057 1225 10109
rect 1241 10076 1293 10109
rect 1241 10057 1273 10076
rect 1273 10057 1293 10076
rect 697 9993 749 10045
rect 765 10042 767 10045
rect 767 10042 801 10045
rect 801 10042 817 10045
rect 765 10002 817 10042
rect 765 9993 767 10002
rect 767 9993 801 10002
rect 801 9993 817 10002
rect 833 9993 885 10045
rect 901 9993 953 10045
rect 969 10042 1003 10045
rect 1003 10042 1021 10045
rect 969 10002 1021 10042
rect 969 9993 1003 10002
rect 1003 9993 1021 10002
rect 1037 9993 1089 10045
rect 1105 9993 1157 10045
rect 1173 9993 1225 10045
rect 1241 10042 1273 10045
rect 1273 10042 1293 10045
rect 2097 10057 2149 10109
rect 2165 10076 2217 10109
rect 2165 10057 2183 10076
rect 2183 10057 2217 10076
rect 2233 10057 2285 10109
rect 2301 10057 2353 10109
rect 2369 10076 2421 10109
rect 2437 10076 2489 10109
rect 2369 10057 2419 10076
rect 2419 10057 2421 10076
rect 2437 10057 2453 10076
rect 2453 10057 2489 10076
rect 2505 10057 2557 10109
rect 2573 10057 2625 10109
rect 2641 10076 2693 10109
rect 2641 10057 2655 10076
rect 2655 10057 2689 10076
rect 2689 10057 2693 10076
rect 1241 10002 1293 10042
rect 1241 9993 1273 10002
rect 1273 9993 1293 10002
rect 697 9929 749 9981
rect 765 9968 767 9981
rect 767 9968 801 9981
rect 801 9968 817 9981
rect 765 9929 817 9968
rect 833 9929 885 9981
rect 901 9929 953 9981
rect 969 9968 1003 9981
rect 1003 9968 1021 9981
rect 969 9929 1021 9968
rect 1037 9929 1089 9981
rect 1105 9929 1157 9981
rect 1173 9929 1225 9981
rect 1241 9968 1273 9981
rect 1273 9968 1293 9981
rect 2097 9993 2149 10045
rect 2165 10042 2183 10045
rect 2183 10042 2217 10045
rect 2165 10002 2217 10042
rect 2165 9993 2183 10002
rect 2183 9993 2217 10002
rect 2233 9993 2285 10045
rect 2301 9993 2353 10045
rect 2369 10042 2419 10045
rect 2419 10042 2421 10045
rect 2437 10042 2453 10045
rect 2453 10042 2489 10045
rect 2369 10002 2421 10042
rect 2437 10002 2489 10042
rect 2369 9993 2419 10002
rect 2419 9993 2421 10002
rect 2437 9993 2453 10002
rect 2453 9993 2489 10002
rect 2505 9993 2557 10045
rect 2573 9993 2625 10045
rect 2641 10042 2655 10045
rect 2655 10042 2689 10045
rect 2689 10042 2693 10045
rect 2641 10002 2693 10042
rect 2641 9993 2655 10002
rect 2655 9993 2689 10002
rect 2689 9993 2693 10002
rect 1241 9929 1293 9968
rect 2097 9929 2149 9981
rect 2165 9968 2183 9981
rect 2183 9968 2217 9981
rect 2165 9929 2217 9968
rect 2233 9929 2285 9981
rect 2301 9929 2353 9981
rect 2369 9968 2419 9981
rect 2419 9968 2421 9981
rect 2437 9968 2453 9981
rect 2453 9968 2489 9981
rect 2369 9929 2421 9968
rect 2437 9929 2489 9968
rect 2505 9929 2557 9981
rect 2573 9929 2625 9981
rect 2641 9968 2655 9981
rect 2655 9968 2689 9981
rect 2689 9968 2693 9981
rect 2641 9929 2693 9968
rect 697 9865 749 9917
rect 765 9894 767 9917
rect 767 9894 801 9917
rect 801 9894 817 9917
rect 765 9865 817 9894
rect 833 9865 885 9917
rect 901 9865 953 9917
rect 969 9894 1003 9917
rect 1003 9894 1021 9917
rect 969 9865 1021 9894
rect 1037 9865 1089 9917
rect 1105 9865 1157 9917
rect 1173 9865 1225 9917
rect 1241 9894 1273 9917
rect 1273 9894 1293 9917
rect 1241 9865 1293 9894
rect 2097 9865 2149 9917
rect 2165 9894 2183 9917
rect 2183 9894 2217 9917
rect 2165 9865 2217 9894
rect 2233 9865 2285 9917
rect 2301 9865 2353 9917
rect 2369 9894 2419 9917
rect 2419 9894 2421 9917
rect 2437 9894 2453 9917
rect 2453 9894 2489 9917
rect 2369 9865 2421 9894
rect 2437 9865 2489 9894
rect 2505 9865 2557 9917
rect 2573 9865 2625 9917
rect 2641 9894 2655 9917
rect 2655 9894 2689 9917
rect 2689 9894 2693 9917
rect 2641 9865 2693 9894
rect 1501 9234 1553 9243
rect 1569 9234 1621 9243
rect 1636 9234 1688 9243
rect 1703 9234 1755 9243
rect 1770 9234 1822 9243
rect 1837 9234 1889 9243
rect 1501 9200 1525 9234
rect 1525 9200 1553 9234
rect 1569 9200 1600 9234
rect 1600 9200 1621 9234
rect 1636 9200 1674 9234
rect 1674 9200 1688 9234
rect 1703 9200 1708 9234
rect 1708 9200 1748 9234
rect 1748 9200 1755 9234
rect 1770 9200 1782 9234
rect 1782 9200 1822 9234
rect 1837 9200 1856 9234
rect 1856 9200 1889 9234
rect 1501 9191 1553 9200
rect 1569 9191 1621 9200
rect 1636 9191 1688 9200
rect 1703 9191 1755 9200
rect 1770 9191 1822 9200
rect 1837 9191 1889 9200
rect 697 8559 749 8611
rect 765 8587 767 8611
rect 767 8587 801 8611
rect 801 8587 817 8611
rect 765 8559 817 8587
rect 833 8559 885 8611
rect 901 8559 953 8611
rect 969 8587 1003 8611
rect 1003 8587 1021 8611
rect 969 8559 1021 8587
rect 1037 8559 1089 8611
rect 1105 8559 1157 8611
rect 1173 8559 1225 8611
rect 1241 8587 1273 8611
rect 1273 8587 1293 8611
rect 1241 8559 1293 8587
rect 2097 8559 2149 8611
rect 2165 8587 2183 8611
rect 2183 8587 2217 8611
rect 2165 8559 2217 8587
rect 2233 8559 2285 8611
rect 2301 8559 2353 8611
rect 2369 8587 2419 8611
rect 2419 8587 2421 8611
rect 2437 8587 2453 8611
rect 2453 8587 2489 8611
rect 2369 8559 2421 8587
rect 2437 8559 2489 8587
rect 2505 8559 2557 8611
rect 2573 8559 2625 8611
rect 2641 8587 2655 8611
rect 2655 8587 2689 8611
rect 2689 8587 2693 8611
rect 2641 8559 2693 8587
rect 697 8495 749 8547
rect 765 8514 767 8547
rect 767 8514 801 8547
rect 801 8514 817 8547
rect 765 8495 817 8514
rect 833 8495 885 8547
rect 901 8495 953 8547
rect 969 8514 1003 8547
rect 1003 8514 1021 8547
rect 969 8495 1021 8514
rect 1037 8495 1089 8547
rect 1105 8495 1157 8547
rect 1173 8495 1225 8547
rect 1241 8514 1273 8547
rect 1273 8514 1293 8547
rect 1241 8495 1293 8514
rect 2097 8495 2149 8547
rect 2165 8514 2183 8547
rect 2183 8514 2217 8547
rect 2165 8495 2217 8514
rect 2233 8495 2285 8547
rect 2301 8495 2353 8547
rect 2369 8514 2419 8547
rect 2419 8514 2421 8547
rect 2437 8514 2453 8547
rect 2453 8514 2489 8547
rect 2369 8495 2421 8514
rect 2437 8495 2489 8514
rect 2505 8495 2557 8547
rect 2573 8495 2625 8547
rect 2641 8514 2655 8547
rect 2655 8514 2689 8547
rect 2689 8514 2693 8547
rect 2641 8495 2693 8514
rect 697 8431 749 8483
rect 765 8475 817 8483
rect 765 8441 767 8475
rect 767 8441 801 8475
rect 801 8441 817 8475
rect 765 8431 817 8441
rect 833 8431 885 8483
rect 901 8431 953 8483
rect 969 8475 1021 8483
rect 969 8441 1003 8475
rect 1003 8441 1021 8475
rect 969 8431 1021 8441
rect 1037 8431 1089 8483
rect 1105 8431 1157 8483
rect 1173 8431 1225 8483
rect 1241 8475 1293 8483
rect 1241 8441 1273 8475
rect 1273 8441 1293 8475
rect 1241 8431 1293 8441
rect 2097 8431 2149 8483
rect 2165 8475 2217 8483
rect 2165 8441 2183 8475
rect 2183 8441 2217 8475
rect 2165 8431 2217 8441
rect 2233 8431 2285 8483
rect 2301 8431 2353 8483
rect 2369 8475 2421 8483
rect 2437 8475 2489 8483
rect 2369 8441 2419 8475
rect 2419 8441 2421 8475
rect 2437 8441 2453 8475
rect 2453 8441 2489 8475
rect 2369 8431 2421 8441
rect 2437 8431 2489 8441
rect 2505 8431 2557 8483
rect 2573 8431 2625 8483
rect 2641 8475 2693 8483
rect 2641 8441 2655 8475
rect 2655 8441 2689 8475
rect 2689 8441 2693 8475
rect 2641 8431 2693 8441
rect 697 8367 749 8419
rect 765 8402 817 8419
rect 765 8368 767 8402
rect 767 8368 801 8402
rect 801 8368 817 8402
rect 765 8367 817 8368
rect 833 8367 885 8419
rect 901 8367 953 8419
rect 969 8402 1021 8419
rect 969 8368 1003 8402
rect 1003 8368 1021 8402
rect 969 8367 1021 8368
rect 1037 8367 1089 8419
rect 1105 8367 1157 8419
rect 1173 8367 1225 8419
rect 1241 8402 1293 8419
rect 1241 8368 1273 8402
rect 1273 8368 1293 8402
rect 1241 8367 1293 8368
rect 2097 8367 2149 8419
rect 2165 8402 2217 8419
rect 2165 8368 2183 8402
rect 2183 8368 2217 8402
rect 2165 8367 2217 8368
rect 2233 8367 2285 8419
rect 2301 8367 2353 8419
rect 2369 8402 2421 8419
rect 2437 8402 2489 8419
rect 2369 8368 2419 8402
rect 2419 8368 2421 8402
rect 2437 8368 2453 8402
rect 2453 8368 2489 8402
rect 2369 8367 2421 8368
rect 2437 8367 2489 8368
rect 2505 8367 2557 8419
rect 2573 8367 2625 8419
rect 2641 8402 2693 8419
rect 2641 8368 2655 8402
rect 2655 8368 2689 8402
rect 2689 8368 2693 8402
rect 2641 8367 2693 8368
rect 697 8303 749 8355
rect 765 8329 817 8355
rect 765 8303 767 8329
rect 767 8303 801 8329
rect 801 8303 817 8329
rect 833 8303 885 8355
rect 901 8303 953 8355
rect 969 8329 1021 8355
rect 969 8303 1003 8329
rect 1003 8303 1021 8329
rect 1037 8303 1089 8355
rect 1105 8303 1157 8355
rect 1173 8303 1225 8355
rect 1241 8329 1293 8355
rect 1241 8303 1273 8329
rect 1273 8303 1293 8329
rect 2097 8303 2149 8355
rect 2165 8329 2217 8355
rect 2165 8303 2183 8329
rect 2183 8303 2217 8329
rect 2233 8303 2285 8355
rect 2301 8303 2353 8355
rect 2369 8329 2421 8355
rect 2437 8329 2489 8355
rect 2369 8303 2419 8329
rect 2419 8303 2421 8329
rect 2437 8303 2453 8329
rect 2453 8303 2489 8329
rect 2505 8303 2557 8355
rect 2573 8303 2625 8355
rect 2641 8329 2693 8355
rect 2641 8303 2655 8329
rect 2655 8303 2689 8329
rect 2689 8303 2693 8329
rect 697 8239 749 8291
rect 765 8256 817 8291
rect 765 8239 767 8256
rect 767 8239 801 8256
rect 801 8239 817 8256
rect 833 8239 885 8291
rect 901 8239 953 8291
rect 969 8256 1021 8291
rect 969 8239 1003 8256
rect 1003 8239 1021 8256
rect 1037 8239 1089 8291
rect 1105 8239 1157 8291
rect 1173 8239 1225 8291
rect 1241 8256 1293 8291
rect 1241 8239 1273 8256
rect 1273 8239 1293 8256
rect 697 8175 749 8227
rect 765 8222 767 8227
rect 767 8222 801 8227
rect 801 8222 817 8227
rect 765 8182 817 8222
rect 765 8175 767 8182
rect 767 8175 801 8182
rect 801 8175 817 8182
rect 833 8175 885 8227
rect 901 8175 953 8227
rect 969 8222 1003 8227
rect 1003 8222 1021 8227
rect 969 8182 1021 8222
rect 969 8175 1003 8182
rect 1003 8175 1021 8182
rect 1037 8175 1089 8227
rect 1105 8175 1157 8227
rect 1173 8175 1225 8227
rect 1241 8222 1273 8227
rect 1273 8222 1293 8227
rect 2097 8239 2149 8291
rect 2165 8256 2217 8291
rect 2165 8239 2183 8256
rect 2183 8239 2217 8256
rect 2233 8239 2285 8291
rect 2301 8239 2353 8291
rect 2369 8256 2421 8291
rect 2437 8256 2489 8291
rect 2369 8239 2419 8256
rect 2419 8239 2421 8256
rect 2437 8239 2453 8256
rect 2453 8239 2489 8256
rect 2505 8239 2557 8291
rect 2573 8239 2625 8291
rect 2641 8256 2693 8291
rect 2641 8239 2655 8256
rect 2655 8239 2689 8256
rect 2689 8239 2693 8256
rect 1241 8182 1293 8222
rect 1241 8175 1273 8182
rect 1273 8175 1293 8182
rect 697 8111 749 8163
rect 765 8148 767 8163
rect 767 8148 801 8163
rect 801 8148 817 8163
rect 765 8111 817 8148
rect 833 8111 885 8163
rect 901 8111 953 8163
rect 969 8148 1003 8163
rect 1003 8148 1021 8163
rect 969 8111 1021 8148
rect 1037 8111 1089 8163
rect 1105 8111 1157 8163
rect 1173 8111 1225 8163
rect 1241 8148 1273 8163
rect 1273 8148 1293 8163
rect 2097 8175 2149 8227
rect 2165 8222 2183 8227
rect 2183 8222 2217 8227
rect 2165 8182 2217 8222
rect 2165 8175 2183 8182
rect 2183 8175 2217 8182
rect 2233 8175 2285 8227
rect 2301 8175 2353 8227
rect 2369 8222 2419 8227
rect 2419 8222 2421 8227
rect 2437 8222 2453 8227
rect 2453 8222 2489 8227
rect 2369 8182 2421 8222
rect 2437 8182 2489 8222
rect 2369 8175 2419 8182
rect 2419 8175 2421 8182
rect 2437 8175 2453 8182
rect 2453 8175 2489 8182
rect 2505 8175 2557 8227
rect 2573 8175 2625 8227
rect 2641 8222 2655 8227
rect 2655 8222 2689 8227
rect 2689 8222 2693 8227
rect 2641 8182 2693 8222
rect 2641 8175 2655 8182
rect 2655 8175 2689 8182
rect 2689 8175 2693 8182
rect 1241 8111 1293 8148
rect 2097 8111 2149 8163
rect 2165 8148 2183 8163
rect 2183 8148 2217 8163
rect 2165 8111 2217 8148
rect 2233 8111 2285 8163
rect 2301 8111 2353 8163
rect 2369 8148 2419 8163
rect 2419 8148 2421 8163
rect 2437 8148 2453 8163
rect 2453 8148 2489 8163
rect 2369 8111 2421 8148
rect 2437 8111 2489 8148
rect 2505 8111 2557 8163
rect 2573 8111 2625 8163
rect 2641 8148 2655 8163
rect 2655 8148 2689 8163
rect 2689 8148 2693 8163
rect 2641 8111 2693 8148
rect 697 8047 749 8099
rect 765 8074 767 8099
rect 767 8074 801 8099
rect 801 8074 817 8099
rect 765 8047 817 8074
rect 833 8047 885 8099
rect 901 8047 953 8099
rect 969 8074 1003 8099
rect 1003 8074 1021 8099
rect 969 8047 1021 8074
rect 1037 8047 1089 8099
rect 1105 8047 1157 8099
rect 1173 8047 1225 8099
rect 1241 8074 1273 8099
rect 1273 8074 1293 8099
rect 1241 8047 1293 8074
rect 2097 8047 2149 8099
rect 2165 8074 2183 8099
rect 2183 8074 2217 8099
rect 2165 8047 2217 8074
rect 2233 8047 2285 8099
rect 2301 8047 2353 8099
rect 2369 8074 2419 8099
rect 2419 8074 2421 8099
rect 2437 8074 2453 8099
rect 2453 8074 2489 8099
rect 2369 8047 2421 8074
rect 2437 8047 2489 8074
rect 2505 8047 2557 8099
rect 2573 8047 2625 8099
rect 2641 8074 2655 8099
rect 2655 8074 2689 8099
rect 2689 8074 2693 8099
rect 2641 8047 2693 8074
rect 697 7983 749 8035
rect 765 8034 817 8035
rect 765 8000 767 8034
rect 767 8000 801 8034
rect 801 8000 817 8034
rect 765 7983 817 8000
rect 833 7983 885 8035
rect 901 7983 953 8035
rect 969 8034 1021 8035
rect 969 8000 1003 8034
rect 1003 8000 1021 8034
rect 969 7983 1021 8000
rect 1037 7983 1089 8035
rect 1105 7983 1157 8035
rect 1173 7983 1225 8035
rect 1241 8034 1293 8035
rect 1241 8000 1273 8034
rect 1273 8000 1293 8034
rect 1241 7983 1293 8000
rect 2097 7983 2149 8035
rect 2165 8034 2217 8035
rect 2165 8000 2183 8034
rect 2183 8000 2217 8034
rect 2165 7983 2217 8000
rect 2233 7983 2285 8035
rect 2301 7983 2353 8035
rect 2369 8034 2421 8035
rect 2437 8034 2489 8035
rect 2369 8000 2419 8034
rect 2419 8000 2421 8034
rect 2437 8000 2453 8034
rect 2453 8000 2489 8034
rect 2369 7983 2421 8000
rect 2437 7983 2489 8000
rect 2505 7983 2557 8035
rect 2573 7983 2625 8035
rect 2641 8034 2693 8035
rect 2641 8000 2655 8034
rect 2655 8000 2689 8034
rect 2689 8000 2693 8034
rect 2641 7983 2693 8000
rect 697 7919 749 7971
rect 765 7960 817 7971
rect 765 7926 767 7960
rect 767 7926 801 7960
rect 801 7926 817 7960
rect 765 7919 817 7926
rect 833 7919 885 7971
rect 901 7919 953 7971
rect 969 7960 1021 7971
rect 969 7926 1003 7960
rect 1003 7926 1021 7960
rect 969 7919 1021 7926
rect 1037 7919 1089 7971
rect 1105 7919 1157 7971
rect 1173 7919 1225 7971
rect 1241 7960 1293 7971
rect 1241 7926 1273 7960
rect 1273 7926 1293 7960
rect 1241 7919 1293 7926
rect 2097 7919 2149 7971
rect 2165 7960 2217 7971
rect 2165 7926 2183 7960
rect 2183 7926 2217 7960
rect 2165 7919 2217 7926
rect 2233 7919 2285 7971
rect 2301 7919 2353 7971
rect 2369 7960 2421 7971
rect 2437 7960 2489 7971
rect 2369 7926 2419 7960
rect 2419 7926 2421 7960
rect 2437 7926 2453 7960
rect 2453 7926 2489 7960
rect 2369 7919 2421 7926
rect 2437 7919 2489 7926
rect 2505 7919 2557 7971
rect 2573 7919 2625 7971
rect 2641 7960 2693 7971
rect 2641 7926 2655 7960
rect 2655 7926 2689 7960
rect 2689 7926 2693 7960
rect 2641 7919 2693 7926
rect 697 7855 749 7907
rect 765 7886 817 7907
rect 765 7855 767 7886
rect 767 7855 801 7886
rect 801 7855 817 7886
rect 833 7855 885 7907
rect 901 7855 953 7907
rect 969 7886 1021 7907
rect 969 7855 1003 7886
rect 1003 7855 1021 7886
rect 1037 7855 1089 7907
rect 1105 7855 1157 7907
rect 1173 7855 1225 7907
rect 1241 7886 1293 7907
rect 1241 7855 1273 7886
rect 1273 7855 1293 7886
rect 2097 7855 2149 7907
rect 2165 7886 2217 7907
rect 2165 7855 2183 7886
rect 2183 7855 2217 7886
rect 2233 7855 2285 7907
rect 2301 7855 2353 7907
rect 2369 7886 2421 7907
rect 2437 7886 2489 7907
rect 2369 7855 2419 7886
rect 2419 7855 2421 7886
rect 2437 7855 2453 7886
rect 2453 7855 2489 7886
rect 2505 7855 2557 7907
rect 2573 7855 2625 7907
rect 2641 7886 2693 7907
rect 2641 7855 2655 7886
rect 2655 7855 2689 7886
rect 2689 7855 2693 7886
rect 697 7791 749 7843
rect 765 7812 817 7843
rect 765 7791 767 7812
rect 767 7791 801 7812
rect 801 7791 817 7812
rect 833 7791 885 7843
rect 901 7791 953 7843
rect 969 7812 1021 7843
rect 969 7791 1003 7812
rect 1003 7791 1021 7812
rect 1037 7791 1089 7843
rect 1105 7791 1157 7843
rect 1173 7791 1225 7843
rect 1241 7812 1293 7843
rect 1241 7791 1273 7812
rect 1273 7791 1293 7812
rect 697 7727 749 7779
rect 765 7778 767 7779
rect 767 7778 801 7779
rect 801 7778 817 7779
rect 765 7738 817 7778
rect 765 7727 767 7738
rect 767 7727 801 7738
rect 801 7727 817 7738
rect 833 7727 885 7779
rect 901 7727 953 7779
rect 969 7778 1003 7779
rect 1003 7778 1021 7779
rect 969 7738 1021 7778
rect 969 7727 1003 7738
rect 1003 7727 1021 7738
rect 1037 7727 1089 7779
rect 1105 7727 1157 7779
rect 1173 7727 1225 7779
rect 1241 7778 1273 7779
rect 1273 7778 1293 7779
rect 2097 7791 2149 7843
rect 2165 7812 2217 7843
rect 2165 7791 2183 7812
rect 2183 7791 2217 7812
rect 2233 7791 2285 7843
rect 2301 7791 2353 7843
rect 2369 7812 2421 7843
rect 2437 7812 2489 7843
rect 2369 7791 2419 7812
rect 2419 7791 2421 7812
rect 2437 7791 2453 7812
rect 2453 7791 2489 7812
rect 2505 7791 2557 7843
rect 2573 7791 2625 7843
rect 2641 7812 2693 7843
rect 2641 7791 2655 7812
rect 2655 7791 2689 7812
rect 2689 7791 2693 7812
rect 1241 7738 1293 7778
rect 1241 7727 1273 7738
rect 1273 7727 1293 7738
rect 697 7663 749 7715
rect 765 7704 767 7715
rect 767 7704 801 7715
rect 801 7704 817 7715
rect 765 7664 817 7704
rect 765 7663 767 7664
rect 767 7663 801 7664
rect 801 7663 817 7664
rect 833 7663 885 7715
rect 901 7663 953 7715
rect 969 7704 1003 7715
rect 1003 7704 1021 7715
rect 969 7664 1021 7704
rect 969 7663 1003 7664
rect 1003 7663 1021 7664
rect 1037 7663 1089 7715
rect 1105 7663 1157 7715
rect 1173 7663 1225 7715
rect 1241 7704 1273 7715
rect 1273 7704 1293 7715
rect 2097 7727 2149 7779
rect 2165 7778 2183 7779
rect 2183 7778 2217 7779
rect 2165 7738 2217 7778
rect 2165 7727 2183 7738
rect 2183 7727 2217 7738
rect 2233 7727 2285 7779
rect 2301 7727 2353 7779
rect 2369 7778 2419 7779
rect 2419 7778 2421 7779
rect 2437 7778 2453 7779
rect 2453 7778 2489 7779
rect 2369 7738 2421 7778
rect 2437 7738 2489 7778
rect 2369 7727 2419 7738
rect 2419 7727 2421 7738
rect 2437 7727 2453 7738
rect 2453 7727 2489 7738
rect 2505 7727 2557 7779
rect 2573 7727 2625 7779
rect 2641 7778 2655 7779
rect 2655 7778 2689 7779
rect 2689 7778 2693 7779
rect 2641 7738 2693 7778
rect 2641 7727 2655 7738
rect 2655 7727 2689 7738
rect 2689 7727 2693 7738
rect 1241 7664 1293 7704
rect 1241 7663 1273 7664
rect 1273 7663 1293 7664
rect 2097 7663 2149 7715
rect 2165 7704 2183 7715
rect 2183 7704 2217 7715
rect 2165 7664 2217 7704
rect 2165 7663 2183 7664
rect 2183 7663 2217 7664
rect 2233 7663 2285 7715
rect 2301 7663 2353 7715
rect 2369 7704 2419 7715
rect 2419 7704 2421 7715
rect 2437 7704 2453 7715
rect 2453 7704 2489 7715
rect 2369 7664 2421 7704
rect 2437 7664 2489 7704
rect 2369 7663 2419 7664
rect 2419 7663 2421 7664
rect 2437 7663 2453 7664
rect 2453 7663 2489 7664
rect 2505 7663 2557 7715
rect 2573 7663 2625 7715
rect 2641 7704 2655 7715
rect 2655 7704 2689 7715
rect 2689 7704 2693 7715
rect 2641 7664 2693 7704
rect 2641 7663 2655 7664
rect 2655 7663 2689 7664
rect 2689 7663 2693 7664
rect 1501 7104 1553 7113
rect 1569 7104 1621 7113
rect 1636 7104 1688 7113
rect 1703 7104 1755 7113
rect 1770 7104 1822 7113
rect 1837 7104 1889 7113
rect 1501 7070 1525 7104
rect 1525 7070 1553 7104
rect 1569 7070 1600 7104
rect 1600 7070 1621 7104
rect 1636 7070 1674 7104
rect 1674 7070 1688 7104
rect 1703 7070 1708 7104
rect 1708 7070 1748 7104
rect 1748 7070 1755 7104
rect 1770 7070 1782 7104
rect 1782 7070 1822 7104
rect 1837 7070 1856 7104
rect 1856 7070 1889 7104
rect 1501 7061 1553 7070
rect 1569 7061 1621 7070
rect 1636 7061 1688 7070
rect 1703 7061 1755 7070
rect 1770 7061 1822 7070
rect 1837 7061 1889 7070
rect 697 6449 749 6501
rect 765 6477 817 6501
rect 765 6449 767 6477
rect 767 6449 801 6477
rect 801 6449 817 6477
rect 833 6449 885 6501
rect 901 6449 953 6501
rect 969 6477 1021 6501
rect 969 6449 1003 6477
rect 1003 6449 1021 6477
rect 1037 6449 1089 6501
rect 1105 6449 1157 6501
rect 1173 6449 1225 6501
rect 1241 6477 1293 6501
rect 1241 6449 1273 6477
rect 1273 6449 1293 6477
rect 2097 6449 2149 6501
rect 2165 6477 2217 6501
rect 2165 6449 2183 6477
rect 2183 6449 2217 6477
rect 2233 6449 2285 6501
rect 2301 6449 2353 6501
rect 2369 6477 2421 6501
rect 2437 6477 2489 6501
rect 2369 6449 2419 6477
rect 2419 6449 2421 6477
rect 2437 6449 2453 6477
rect 2453 6449 2489 6477
rect 2505 6449 2557 6501
rect 2573 6449 2625 6501
rect 2641 6477 2693 6501
rect 2641 6449 2655 6477
rect 2655 6449 2689 6477
rect 2689 6449 2693 6477
rect 697 6385 749 6437
rect 765 6404 817 6437
rect 765 6385 767 6404
rect 767 6385 801 6404
rect 801 6385 817 6404
rect 833 6385 885 6437
rect 901 6385 953 6437
rect 969 6404 1021 6437
rect 969 6385 1003 6404
rect 1003 6385 1021 6404
rect 1037 6385 1089 6437
rect 1105 6385 1157 6437
rect 1173 6385 1225 6437
rect 1241 6404 1293 6437
rect 1241 6385 1273 6404
rect 1273 6385 1293 6404
rect 697 6321 749 6373
rect 765 6370 767 6373
rect 767 6370 801 6373
rect 801 6370 817 6373
rect 765 6331 817 6370
rect 765 6321 767 6331
rect 767 6321 801 6331
rect 801 6321 817 6331
rect 833 6321 885 6373
rect 901 6321 953 6373
rect 969 6370 1003 6373
rect 1003 6370 1021 6373
rect 969 6331 1021 6370
rect 969 6321 1003 6331
rect 1003 6321 1021 6331
rect 1037 6321 1089 6373
rect 1105 6321 1157 6373
rect 1173 6321 1225 6373
rect 1241 6370 1273 6373
rect 1273 6370 1293 6373
rect 2097 6385 2149 6437
rect 2165 6404 2217 6437
rect 2165 6385 2183 6404
rect 2183 6385 2217 6404
rect 2233 6385 2285 6437
rect 2301 6385 2353 6437
rect 2369 6404 2421 6437
rect 2437 6404 2489 6437
rect 2369 6385 2419 6404
rect 2419 6385 2421 6404
rect 2437 6385 2453 6404
rect 2453 6385 2489 6404
rect 2505 6385 2557 6437
rect 2573 6385 2625 6437
rect 2641 6404 2693 6437
rect 2641 6385 2655 6404
rect 2655 6385 2689 6404
rect 2689 6385 2693 6404
rect 1241 6331 1293 6370
rect 1241 6321 1273 6331
rect 1273 6321 1293 6331
rect 697 6257 749 6309
rect 765 6297 767 6309
rect 767 6297 801 6309
rect 801 6297 817 6309
rect 765 6258 817 6297
rect 765 6257 767 6258
rect 767 6257 801 6258
rect 801 6257 817 6258
rect 833 6257 885 6309
rect 901 6257 953 6309
rect 969 6297 1003 6309
rect 1003 6297 1021 6309
rect 969 6258 1021 6297
rect 969 6257 1003 6258
rect 1003 6257 1021 6258
rect 1037 6257 1089 6309
rect 1105 6257 1157 6309
rect 1173 6257 1225 6309
rect 1241 6297 1273 6309
rect 1273 6297 1293 6309
rect 2097 6321 2149 6373
rect 2165 6370 2183 6373
rect 2183 6370 2217 6373
rect 2165 6331 2217 6370
rect 2165 6321 2183 6331
rect 2183 6321 2217 6331
rect 2233 6321 2285 6373
rect 2301 6321 2353 6373
rect 2369 6370 2419 6373
rect 2419 6370 2421 6373
rect 2437 6370 2453 6373
rect 2453 6370 2489 6373
rect 2369 6331 2421 6370
rect 2437 6331 2489 6370
rect 2369 6321 2419 6331
rect 2419 6321 2421 6331
rect 2437 6321 2453 6331
rect 2453 6321 2489 6331
rect 2505 6321 2557 6373
rect 2573 6321 2625 6373
rect 2641 6370 2655 6373
rect 2655 6370 2689 6373
rect 2689 6370 2693 6373
rect 2641 6331 2693 6370
rect 2641 6321 2655 6331
rect 2655 6321 2689 6331
rect 2689 6321 2693 6331
rect 1241 6258 1293 6297
rect 1241 6257 1273 6258
rect 1273 6257 1293 6258
rect 697 6193 749 6245
rect 765 6224 767 6245
rect 767 6224 801 6245
rect 801 6224 817 6245
rect 765 6193 817 6224
rect 833 6193 885 6245
rect 901 6193 953 6245
rect 969 6224 1003 6245
rect 1003 6224 1021 6245
rect 969 6193 1021 6224
rect 1037 6193 1089 6245
rect 1105 6193 1157 6245
rect 1173 6193 1225 6245
rect 1241 6224 1273 6245
rect 1273 6224 1293 6245
rect 2097 6257 2149 6309
rect 2165 6297 2183 6309
rect 2183 6297 2217 6309
rect 2165 6258 2217 6297
rect 2165 6257 2183 6258
rect 2183 6257 2217 6258
rect 2233 6257 2285 6309
rect 2301 6257 2353 6309
rect 2369 6297 2419 6309
rect 2419 6297 2421 6309
rect 2437 6297 2453 6309
rect 2453 6297 2489 6309
rect 2369 6258 2421 6297
rect 2437 6258 2489 6297
rect 2369 6257 2419 6258
rect 2419 6257 2421 6258
rect 2437 6257 2453 6258
rect 2453 6257 2489 6258
rect 2505 6257 2557 6309
rect 2573 6257 2625 6309
rect 2641 6297 2655 6309
rect 2655 6297 2689 6309
rect 2689 6297 2693 6309
rect 2641 6258 2693 6297
rect 2641 6257 2655 6258
rect 2655 6257 2689 6258
rect 2689 6257 2693 6258
rect 1241 6193 1293 6224
rect 2097 6193 2149 6245
rect 2165 6224 2183 6245
rect 2183 6224 2217 6245
rect 2165 6193 2217 6224
rect 2233 6193 2285 6245
rect 2301 6193 2353 6245
rect 2369 6224 2419 6245
rect 2419 6224 2421 6245
rect 2437 6224 2453 6245
rect 2453 6224 2489 6245
rect 2369 6193 2421 6224
rect 2437 6193 2489 6224
rect 2505 6193 2557 6245
rect 2573 6193 2625 6245
rect 2641 6224 2655 6245
rect 2655 6224 2689 6245
rect 2689 6224 2693 6245
rect 2641 6193 2693 6224
rect 697 6129 749 6181
rect 765 6151 767 6181
rect 767 6151 801 6181
rect 801 6151 817 6181
rect 765 6129 817 6151
rect 833 6129 885 6181
rect 901 6129 953 6181
rect 969 6151 1003 6181
rect 1003 6151 1021 6181
rect 969 6129 1021 6151
rect 1037 6129 1089 6181
rect 1105 6129 1157 6181
rect 1173 6129 1225 6181
rect 1241 6151 1273 6181
rect 1273 6151 1293 6181
rect 1241 6129 1293 6151
rect 2097 6129 2149 6181
rect 2165 6151 2183 6181
rect 2183 6151 2217 6181
rect 2165 6129 2217 6151
rect 2233 6129 2285 6181
rect 2301 6129 2353 6181
rect 2369 6151 2419 6181
rect 2419 6151 2421 6181
rect 2437 6151 2453 6181
rect 2453 6151 2489 6181
rect 2369 6129 2421 6151
rect 2437 6129 2489 6151
rect 2505 6129 2557 6181
rect 2573 6129 2625 6181
rect 2641 6151 2655 6181
rect 2655 6151 2689 6181
rect 2689 6151 2693 6181
rect 2641 6129 2693 6151
rect 697 6065 749 6117
rect 765 6112 817 6117
rect 765 6078 767 6112
rect 767 6078 801 6112
rect 801 6078 817 6112
rect 765 6065 817 6078
rect 833 6065 885 6117
rect 901 6065 953 6117
rect 969 6112 1021 6117
rect 969 6078 1003 6112
rect 1003 6078 1021 6112
rect 969 6065 1021 6078
rect 1037 6065 1089 6117
rect 1105 6065 1157 6117
rect 1173 6065 1225 6117
rect 1241 6112 1293 6117
rect 1241 6078 1273 6112
rect 1273 6078 1293 6112
rect 1241 6065 1293 6078
rect 2097 6065 2149 6117
rect 2165 6112 2217 6117
rect 2165 6078 2183 6112
rect 2183 6078 2217 6112
rect 2165 6065 2217 6078
rect 2233 6065 2285 6117
rect 2301 6065 2353 6117
rect 2369 6112 2421 6117
rect 2437 6112 2489 6117
rect 2369 6078 2419 6112
rect 2419 6078 2421 6112
rect 2437 6078 2453 6112
rect 2453 6078 2489 6112
rect 2369 6065 2421 6078
rect 2437 6065 2489 6078
rect 2505 6065 2557 6117
rect 2573 6065 2625 6117
rect 2641 6112 2693 6117
rect 2641 6078 2655 6112
rect 2655 6078 2689 6112
rect 2689 6078 2693 6112
rect 2641 6065 2693 6078
rect 697 6001 749 6053
rect 765 6038 817 6053
rect 765 6004 767 6038
rect 767 6004 801 6038
rect 801 6004 817 6038
rect 765 6001 817 6004
rect 833 6001 885 6053
rect 901 6001 953 6053
rect 969 6038 1021 6053
rect 969 6004 1003 6038
rect 1003 6004 1021 6038
rect 969 6001 1021 6004
rect 1037 6001 1089 6053
rect 1105 6001 1157 6053
rect 1173 6001 1225 6053
rect 1241 6038 1293 6053
rect 1241 6004 1273 6038
rect 1273 6004 1293 6038
rect 1241 6001 1293 6004
rect 2097 6001 2149 6053
rect 2165 6038 2217 6053
rect 2165 6004 2183 6038
rect 2183 6004 2217 6038
rect 2165 6001 2217 6004
rect 2233 6001 2285 6053
rect 2301 6001 2353 6053
rect 2369 6038 2421 6053
rect 2437 6038 2489 6053
rect 2369 6004 2419 6038
rect 2419 6004 2421 6038
rect 2437 6004 2453 6038
rect 2453 6004 2489 6038
rect 2369 6001 2421 6004
rect 2437 6001 2489 6004
rect 2505 6001 2557 6053
rect 2573 6001 2625 6053
rect 2641 6038 2693 6053
rect 2641 6004 2655 6038
rect 2655 6004 2689 6038
rect 2689 6004 2693 6038
rect 2641 6001 2693 6004
rect 697 5937 749 5989
rect 765 5964 817 5989
rect 765 5937 767 5964
rect 767 5937 801 5964
rect 801 5937 817 5964
rect 833 5937 885 5989
rect 901 5937 953 5989
rect 969 5964 1021 5989
rect 969 5937 1003 5964
rect 1003 5937 1021 5964
rect 1037 5937 1089 5989
rect 1105 5937 1157 5989
rect 1173 5937 1225 5989
rect 1241 5964 1293 5989
rect 1241 5937 1273 5964
rect 1273 5937 1293 5964
rect 2097 5937 2149 5989
rect 2165 5964 2217 5989
rect 2165 5937 2183 5964
rect 2183 5937 2217 5964
rect 2233 5937 2285 5989
rect 2301 5937 2353 5989
rect 2369 5964 2421 5989
rect 2437 5964 2489 5989
rect 2369 5937 2419 5964
rect 2419 5937 2421 5964
rect 2437 5937 2453 5964
rect 2453 5937 2489 5964
rect 2505 5937 2557 5989
rect 2573 5937 2625 5989
rect 2641 5964 2693 5989
rect 2641 5937 2655 5964
rect 2655 5937 2689 5964
rect 2689 5937 2693 5964
rect 697 5873 749 5925
rect 765 5890 817 5925
rect 765 5873 767 5890
rect 767 5873 801 5890
rect 801 5873 817 5890
rect 833 5873 885 5925
rect 901 5873 953 5925
rect 969 5890 1021 5925
rect 969 5873 1003 5890
rect 1003 5873 1021 5890
rect 1037 5873 1089 5925
rect 1105 5873 1157 5925
rect 1173 5873 1225 5925
rect 1241 5890 1293 5925
rect 1241 5873 1273 5890
rect 1273 5873 1293 5890
rect 697 5809 749 5861
rect 765 5856 767 5861
rect 767 5856 801 5861
rect 801 5856 817 5861
rect 765 5816 817 5856
rect 765 5809 767 5816
rect 767 5809 801 5816
rect 801 5809 817 5816
rect 833 5809 885 5861
rect 901 5809 953 5861
rect 969 5856 1003 5861
rect 1003 5856 1021 5861
rect 969 5816 1021 5856
rect 969 5809 1003 5816
rect 1003 5809 1021 5816
rect 1037 5809 1089 5861
rect 1105 5809 1157 5861
rect 1173 5809 1225 5861
rect 1241 5856 1273 5861
rect 1273 5856 1293 5861
rect 2097 5873 2149 5925
rect 2165 5890 2217 5925
rect 2165 5873 2183 5890
rect 2183 5873 2217 5890
rect 2233 5873 2285 5925
rect 2301 5873 2353 5925
rect 2369 5890 2421 5925
rect 2437 5890 2489 5925
rect 2369 5873 2419 5890
rect 2419 5873 2421 5890
rect 2437 5873 2453 5890
rect 2453 5873 2489 5890
rect 2505 5873 2557 5925
rect 2573 5873 2625 5925
rect 2641 5890 2693 5925
rect 2641 5873 2655 5890
rect 2655 5873 2689 5890
rect 2689 5873 2693 5890
rect 1241 5816 1293 5856
rect 1241 5809 1273 5816
rect 1273 5809 1293 5816
rect 697 5745 749 5797
rect 765 5782 767 5797
rect 767 5782 801 5797
rect 801 5782 817 5797
rect 765 5745 817 5782
rect 833 5745 885 5797
rect 901 5745 953 5797
rect 969 5782 1003 5797
rect 1003 5782 1021 5797
rect 969 5745 1021 5782
rect 1037 5745 1089 5797
rect 1105 5745 1157 5797
rect 1173 5745 1225 5797
rect 1241 5782 1273 5797
rect 1273 5782 1293 5797
rect 2097 5809 2149 5861
rect 2165 5856 2183 5861
rect 2183 5856 2217 5861
rect 2165 5816 2217 5856
rect 2165 5809 2183 5816
rect 2183 5809 2217 5816
rect 2233 5809 2285 5861
rect 2301 5809 2353 5861
rect 2369 5856 2419 5861
rect 2419 5856 2421 5861
rect 2437 5856 2453 5861
rect 2453 5856 2489 5861
rect 2369 5816 2421 5856
rect 2437 5816 2489 5856
rect 2369 5809 2419 5816
rect 2419 5809 2421 5816
rect 2437 5809 2453 5816
rect 2453 5809 2489 5816
rect 2505 5809 2557 5861
rect 2573 5809 2625 5861
rect 2641 5856 2655 5861
rect 2655 5856 2689 5861
rect 2689 5856 2693 5861
rect 2641 5816 2693 5856
rect 2641 5809 2655 5816
rect 2655 5809 2689 5816
rect 2689 5809 2693 5816
rect 1241 5745 1293 5782
rect 2097 5745 2149 5797
rect 2165 5782 2183 5797
rect 2183 5782 2217 5797
rect 2165 5745 2217 5782
rect 2233 5745 2285 5797
rect 2301 5745 2353 5797
rect 2369 5782 2419 5797
rect 2419 5782 2421 5797
rect 2437 5782 2453 5797
rect 2453 5782 2489 5797
rect 2369 5745 2421 5782
rect 2437 5745 2489 5782
rect 2505 5745 2557 5797
rect 2573 5745 2625 5797
rect 2641 5782 2655 5797
rect 2655 5782 2689 5797
rect 2689 5782 2693 5797
rect 2641 5745 2693 5782
rect 697 5681 749 5733
rect 765 5708 767 5733
rect 767 5708 801 5733
rect 801 5708 817 5733
rect 765 5681 817 5708
rect 833 5681 885 5733
rect 901 5681 953 5733
rect 969 5708 1003 5733
rect 1003 5708 1021 5733
rect 969 5681 1021 5708
rect 1037 5681 1089 5733
rect 1105 5681 1157 5733
rect 1173 5681 1225 5733
rect 1241 5708 1273 5733
rect 1273 5708 1293 5733
rect 1241 5681 1293 5708
rect 2097 5681 2149 5733
rect 2165 5708 2183 5733
rect 2183 5708 2217 5733
rect 2165 5681 2217 5708
rect 2233 5681 2285 5733
rect 2301 5681 2353 5733
rect 2369 5708 2419 5733
rect 2419 5708 2421 5733
rect 2437 5708 2453 5733
rect 2453 5708 2489 5733
rect 2369 5681 2421 5708
rect 2437 5681 2489 5708
rect 2505 5681 2557 5733
rect 2573 5681 2625 5733
rect 2641 5708 2655 5733
rect 2655 5708 2689 5733
rect 2689 5708 2693 5733
rect 2641 5681 2693 5708
rect 697 5617 749 5669
rect 765 5668 817 5669
rect 765 5634 767 5668
rect 767 5634 801 5668
rect 801 5634 817 5668
rect 765 5617 817 5634
rect 833 5617 885 5669
rect 901 5617 953 5669
rect 969 5668 1021 5669
rect 969 5634 1003 5668
rect 1003 5634 1021 5668
rect 969 5617 1021 5634
rect 1037 5617 1089 5669
rect 1105 5617 1157 5669
rect 1173 5617 1225 5669
rect 1241 5668 1293 5669
rect 1241 5634 1273 5668
rect 1273 5634 1293 5668
rect 1241 5617 1293 5634
rect 2097 5617 2149 5669
rect 2165 5668 2217 5669
rect 2165 5634 2183 5668
rect 2183 5634 2217 5668
rect 2165 5617 2217 5634
rect 2233 5617 2285 5669
rect 2301 5617 2353 5669
rect 2369 5668 2421 5669
rect 2437 5668 2489 5669
rect 2369 5634 2419 5668
rect 2419 5634 2421 5668
rect 2437 5634 2453 5668
rect 2453 5634 2489 5668
rect 2369 5617 2421 5634
rect 2437 5617 2489 5634
rect 2505 5617 2557 5669
rect 2573 5617 2625 5669
rect 2641 5668 2693 5669
rect 2641 5634 2655 5668
rect 2655 5634 2689 5668
rect 2689 5634 2693 5668
rect 2641 5617 2693 5634
rect 697 5553 749 5605
rect 765 5594 817 5605
rect 765 5560 767 5594
rect 767 5560 801 5594
rect 801 5560 817 5594
rect 765 5553 817 5560
rect 833 5553 885 5605
rect 901 5553 953 5605
rect 969 5594 1021 5605
rect 969 5560 1003 5594
rect 1003 5560 1021 5594
rect 969 5553 1021 5560
rect 1037 5553 1089 5605
rect 1105 5553 1157 5605
rect 1173 5553 1225 5605
rect 1241 5594 1293 5605
rect 1241 5560 1273 5594
rect 1273 5560 1293 5594
rect 1241 5553 1293 5560
rect 2097 5553 2149 5605
rect 2165 5594 2217 5605
rect 2165 5560 2183 5594
rect 2183 5560 2217 5594
rect 2165 5553 2217 5560
rect 2233 5553 2285 5605
rect 2301 5553 2353 5605
rect 2369 5594 2421 5605
rect 2437 5594 2489 5605
rect 2369 5560 2419 5594
rect 2419 5560 2421 5594
rect 2437 5560 2453 5594
rect 2453 5560 2489 5594
rect 2369 5553 2421 5560
rect 2437 5553 2489 5560
rect 2505 5553 2557 5605
rect 2573 5553 2625 5605
rect 2641 5594 2693 5605
rect 2641 5560 2655 5594
rect 2655 5560 2689 5594
rect 2689 5560 2693 5594
rect 2641 5553 2693 5560
rect 1501 4974 1553 4983
rect 1569 4974 1621 4983
rect 1636 4974 1688 4983
rect 1703 4974 1755 4983
rect 1770 4974 1822 4983
rect 1837 4974 1889 4983
rect 1501 4940 1525 4974
rect 1525 4940 1553 4974
rect 1569 4940 1600 4974
rect 1600 4940 1621 4974
rect 1636 4940 1674 4974
rect 1674 4940 1688 4974
rect 1703 4940 1708 4974
rect 1708 4940 1748 4974
rect 1748 4940 1755 4974
rect 1770 4940 1782 4974
rect 1782 4940 1822 4974
rect 1837 4940 1856 4974
rect 1856 4940 1889 4974
rect 1501 4931 1553 4940
rect 1569 4931 1621 4940
rect 1636 4931 1688 4940
rect 1703 4931 1755 4940
rect 1770 4931 1822 4940
rect 1837 4931 1889 4940
rect 697 4385 749 4437
rect 765 4434 817 4437
rect 765 4400 767 4434
rect 767 4400 801 4434
rect 801 4400 817 4434
rect 765 4385 817 4400
rect 833 4385 885 4437
rect 901 4385 953 4437
rect 969 4434 1021 4437
rect 969 4400 1003 4434
rect 1003 4400 1021 4434
rect 969 4385 1021 4400
rect 1037 4385 1089 4437
rect 1105 4385 1157 4437
rect 1173 4385 1225 4437
rect 1241 4434 1293 4437
rect 1241 4400 1273 4434
rect 1273 4400 1293 4434
rect 1241 4385 1293 4400
rect 2097 4385 2149 4437
rect 2165 4434 2217 4437
rect 2165 4400 2183 4434
rect 2183 4400 2217 4434
rect 2165 4385 2217 4400
rect 2233 4385 2285 4437
rect 2301 4385 2353 4437
rect 2369 4434 2421 4437
rect 2437 4434 2489 4437
rect 2369 4400 2419 4434
rect 2419 4400 2421 4434
rect 2437 4400 2453 4434
rect 2453 4400 2489 4434
rect 2369 4385 2421 4400
rect 2437 4385 2489 4400
rect 2505 4385 2557 4437
rect 2573 4385 2625 4437
rect 2641 4434 2693 4437
rect 2641 4400 2655 4434
rect 2655 4400 2689 4434
rect 2689 4400 2693 4434
rect 2641 4385 2693 4400
rect 697 4321 749 4373
rect 765 4361 817 4373
rect 765 4327 767 4361
rect 767 4327 801 4361
rect 801 4327 817 4361
rect 765 4321 817 4327
rect 833 4321 885 4373
rect 901 4321 953 4373
rect 969 4361 1021 4373
rect 969 4327 1003 4361
rect 1003 4327 1021 4361
rect 969 4321 1021 4327
rect 1037 4321 1089 4373
rect 1105 4321 1157 4373
rect 1173 4321 1225 4373
rect 1241 4361 1293 4373
rect 1241 4327 1273 4361
rect 1273 4327 1293 4361
rect 1241 4321 1293 4327
rect 2097 4321 2149 4373
rect 2165 4361 2217 4373
rect 2165 4327 2183 4361
rect 2183 4327 2217 4361
rect 2165 4321 2217 4327
rect 2233 4321 2285 4373
rect 2301 4321 2353 4373
rect 2369 4361 2421 4373
rect 2437 4361 2489 4373
rect 2369 4327 2419 4361
rect 2419 4327 2421 4361
rect 2437 4327 2453 4361
rect 2453 4327 2489 4361
rect 2369 4321 2421 4327
rect 2437 4321 2489 4327
rect 2505 4321 2557 4373
rect 2573 4321 2625 4373
rect 2641 4361 2693 4373
rect 2641 4327 2655 4361
rect 2655 4327 2689 4361
rect 2689 4327 2693 4361
rect 2641 4321 2693 4327
rect 697 4257 749 4309
rect 765 4288 817 4309
rect 765 4257 767 4288
rect 767 4257 801 4288
rect 801 4257 817 4288
rect 833 4257 885 4309
rect 901 4257 953 4309
rect 969 4288 1021 4309
rect 969 4257 1003 4288
rect 1003 4257 1021 4288
rect 1037 4257 1089 4309
rect 1105 4257 1157 4309
rect 1173 4257 1225 4309
rect 1241 4288 1293 4309
rect 1241 4257 1273 4288
rect 1273 4257 1293 4288
rect 2097 4257 2149 4309
rect 2165 4288 2217 4309
rect 2165 4257 2183 4288
rect 2183 4257 2217 4288
rect 2233 4257 2285 4309
rect 2301 4257 2353 4309
rect 2369 4288 2421 4309
rect 2437 4288 2489 4309
rect 2369 4257 2419 4288
rect 2419 4257 2421 4288
rect 2437 4257 2453 4288
rect 2453 4257 2489 4288
rect 2505 4257 2557 4309
rect 2573 4257 2625 4309
rect 2641 4288 2693 4309
rect 2641 4257 2655 4288
rect 2655 4257 2689 4288
rect 2689 4257 2693 4288
rect 697 4193 749 4245
rect 765 4215 817 4245
rect 765 4193 767 4215
rect 767 4193 801 4215
rect 801 4193 817 4215
rect 833 4193 885 4245
rect 901 4193 953 4245
rect 969 4215 1021 4245
rect 969 4193 1003 4215
rect 1003 4193 1021 4215
rect 1037 4193 1089 4245
rect 1105 4193 1157 4245
rect 1173 4193 1225 4245
rect 1241 4215 1293 4245
rect 1241 4193 1273 4215
rect 1273 4193 1293 4215
rect 2097 4193 2149 4245
rect 2165 4215 2217 4245
rect 2165 4193 2183 4215
rect 2183 4193 2217 4215
rect 2233 4193 2285 4245
rect 2301 4193 2353 4245
rect 2369 4215 2421 4245
rect 2437 4215 2489 4245
rect 2369 4193 2419 4215
rect 2419 4193 2421 4215
rect 2437 4193 2453 4215
rect 2453 4193 2489 4215
rect 2505 4193 2557 4245
rect 2573 4193 2625 4245
rect 2641 4215 2693 4245
rect 2641 4193 2655 4215
rect 2655 4193 2689 4215
rect 2689 4193 2693 4215
rect 697 4129 749 4181
rect 765 4142 817 4181
rect 765 4129 767 4142
rect 767 4129 801 4142
rect 801 4129 817 4142
rect 833 4129 885 4181
rect 901 4129 953 4181
rect 969 4142 1021 4181
rect 969 4129 1003 4142
rect 1003 4129 1021 4142
rect 1037 4129 1089 4181
rect 1105 4129 1157 4181
rect 1173 4129 1225 4181
rect 1241 4142 1293 4181
rect 1241 4129 1273 4142
rect 1273 4129 1293 4142
rect 697 4065 749 4117
rect 765 4108 767 4117
rect 767 4108 801 4117
rect 801 4108 817 4117
rect 765 4069 817 4108
rect 765 4065 767 4069
rect 767 4065 801 4069
rect 801 4065 817 4069
rect 833 4065 885 4117
rect 901 4065 953 4117
rect 969 4108 1003 4117
rect 1003 4108 1021 4117
rect 969 4069 1021 4108
rect 969 4065 1003 4069
rect 1003 4065 1021 4069
rect 1037 4065 1089 4117
rect 1105 4065 1157 4117
rect 1173 4065 1225 4117
rect 1241 4108 1273 4117
rect 1273 4108 1293 4117
rect 2097 4129 2149 4181
rect 2165 4142 2217 4181
rect 2165 4129 2183 4142
rect 2183 4129 2217 4142
rect 2233 4129 2285 4181
rect 2301 4129 2353 4181
rect 2369 4142 2421 4181
rect 2437 4142 2489 4181
rect 2369 4129 2419 4142
rect 2419 4129 2421 4142
rect 2437 4129 2453 4142
rect 2453 4129 2489 4142
rect 2505 4129 2557 4181
rect 2573 4129 2625 4181
rect 2641 4142 2693 4181
rect 2641 4129 2655 4142
rect 2655 4129 2689 4142
rect 2689 4129 2693 4142
rect 1241 4069 1293 4108
rect 1241 4065 1273 4069
rect 1273 4065 1293 4069
rect 697 4001 749 4053
rect 765 4035 767 4053
rect 767 4035 801 4053
rect 801 4035 817 4053
rect 765 4001 817 4035
rect 833 4001 885 4053
rect 901 4001 953 4053
rect 969 4035 1003 4053
rect 1003 4035 1021 4053
rect 969 4001 1021 4035
rect 1037 4001 1089 4053
rect 1105 4001 1157 4053
rect 1173 4001 1225 4053
rect 1241 4035 1273 4053
rect 1273 4035 1293 4053
rect 2097 4065 2149 4117
rect 2165 4108 2183 4117
rect 2183 4108 2217 4117
rect 2165 4069 2217 4108
rect 2165 4065 2183 4069
rect 2183 4065 2217 4069
rect 2233 4065 2285 4117
rect 2301 4065 2353 4117
rect 2369 4108 2419 4117
rect 2419 4108 2421 4117
rect 2437 4108 2453 4117
rect 2453 4108 2489 4117
rect 2369 4069 2421 4108
rect 2437 4069 2489 4108
rect 2369 4065 2419 4069
rect 2419 4065 2421 4069
rect 2437 4065 2453 4069
rect 2453 4065 2489 4069
rect 2505 4065 2557 4117
rect 2573 4065 2625 4117
rect 2641 4108 2655 4117
rect 2655 4108 2689 4117
rect 2689 4108 2693 4117
rect 2641 4069 2693 4108
rect 2641 4065 2655 4069
rect 2655 4065 2689 4069
rect 2689 4065 2693 4069
rect 1241 4001 1293 4035
rect 2097 4001 2149 4053
rect 2165 4035 2183 4053
rect 2183 4035 2217 4053
rect 2165 4001 2217 4035
rect 2233 4001 2285 4053
rect 2301 4001 2353 4053
rect 2369 4035 2419 4053
rect 2419 4035 2421 4053
rect 2437 4035 2453 4053
rect 2453 4035 2489 4053
rect 2369 4001 2421 4035
rect 2437 4001 2489 4035
rect 2505 4001 2557 4053
rect 2573 4001 2625 4053
rect 2641 4035 2655 4053
rect 2655 4035 2689 4053
rect 2689 4035 2693 4053
rect 2641 4001 2693 4035
rect 697 3937 749 3989
rect 765 3962 767 3989
rect 767 3962 801 3989
rect 801 3962 817 3989
rect 765 3937 817 3962
rect 833 3937 885 3989
rect 901 3937 953 3989
rect 969 3962 1003 3989
rect 1003 3962 1021 3989
rect 969 3937 1021 3962
rect 1037 3937 1089 3989
rect 1105 3937 1157 3989
rect 1173 3937 1225 3989
rect 1241 3962 1273 3989
rect 1273 3962 1293 3989
rect 1241 3937 1293 3962
rect 2097 3937 2149 3989
rect 2165 3962 2183 3989
rect 2183 3962 2217 3989
rect 2165 3937 2217 3962
rect 2233 3937 2285 3989
rect 2301 3937 2353 3989
rect 2369 3962 2419 3989
rect 2419 3962 2421 3989
rect 2437 3962 2453 3989
rect 2453 3962 2489 3989
rect 2369 3937 2421 3962
rect 2437 3937 2489 3962
rect 2505 3937 2557 3989
rect 2573 3937 2625 3989
rect 2641 3962 2655 3989
rect 2655 3962 2689 3989
rect 2689 3962 2693 3989
rect 2641 3937 2693 3962
rect 697 3873 749 3925
rect 765 3922 817 3925
rect 765 3888 767 3922
rect 767 3888 801 3922
rect 801 3888 817 3922
rect 765 3873 817 3888
rect 833 3873 885 3925
rect 901 3873 953 3925
rect 969 3922 1021 3925
rect 969 3888 1003 3922
rect 1003 3888 1021 3922
rect 969 3873 1021 3888
rect 1037 3873 1089 3925
rect 1105 3873 1157 3925
rect 1173 3873 1225 3925
rect 1241 3922 1293 3925
rect 1241 3888 1273 3922
rect 1273 3888 1293 3922
rect 1241 3873 1293 3888
rect 2097 3873 2149 3925
rect 2165 3922 2217 3925
rect 2165 3888 2183 3922
rect 2183 3888 2217 3922
rect 2165 3873 2217 3888
rect 2233 3873 2285 3925
rect 2301 3873 2353 3925
rect 2369 3922 2421 3925
rect 2437 3922 2489 3925
rect 2369 3888 2419 3922
rect 2419 3888 2421 3922
rect 2437 3888 2453 3922
rect 2453 3888 2489 3922
rect 2369 3873 2421 3888
rect 2437 3873 2489 3888
rect 2505 3873 2557 3925
rect 2573 3873 2625 3925
rect 2641 3922 2693 3925
rect 2641 3888 2655 3922
rect 2655 3888 2689 3922
rect 2689 3888 2693 3922
rect 2641 3873 2693 3888
rect 697 3809 749 3861
rect 765 3848 817 3861
rect 765 3814 767 3848
rect 767 3814 801 3848
rect 801 3814 817 3848
rect 765 3809 817 3814
rect 833 3809 885 3861
rect 901 3809 953 3861
rect 969 3848 1021 3861
rect 969 3814 1003 3848
rect 1003 3814 1021 3848
rect 969 3809 1021 3814
rect 1037 3809 1089 3861
rect 1105 3809 1157 3861
rect 1173 3809 1225 3861
rect 1241 3848 1293 3861
rect 1241 3814 1273 3848
rect 1273 3814 1293 3848
rect 1241 3809 1293 3814
rect 2097 3809 2149 3861
rect 2165 3848 2217 3861
rect 2165 3814 2183 3848
rect 2183 3814 2217 3848
rect 2165 3809 2217 3814
rect 2233 3809 2285 3861
rect 2301 3809 2353 3861
rect 2369 3848 2421 3861
rect 2437 3848 2489 3861
rect 2369 3814 2419 3848
rect 2419 3814 2421 3848
rect 2437 3814 2453 3848
rect 2453 3814 2489 3848
rect 2369 3809 2421 3814
rect 2437 3809 2489 3814
rect 2505 3809 2557 3861
rect 2573 3809 2625 3861
rect 2641 3848 2693 3861
rect 2641 3814 2655 3848
rect 2655 3814 2689 3848
rect 2689 3814 2693 3848
rect 2641 3809 2693 3814
rect 697 3745 749 3797
rect 765 3774 817 3797
rect 765 3745 767 3774
rect 767 3745 801 3774
rect 801 3745 817 3774
rect 833 3745 885 3797
rect 901 3745 953 3797
rect 969 3774 1021 3797
rect 969 3745 1003 3774
rect 1003 3745 1021 3774
rect 1037 3745 1089 3797
rect 1105 3745 1157 3797
rect 1173 3745 1225 3797
rect 1241 3774 1293 3797
rect 1241 3745 1273 3774
rect 1273 3745 1293 3774
rect 2097 3745 2149 3797
rect 2165 3774 2217 3797
rect 2165 3745 2183 3774
rect 2183 3745 2217 3774
rect 2233 3745 2285 3797
rect 2301 3745 2353 3797
rect 2369 3774 2421 3797
rect 2437 3774 2489 3797
rect 2369 3745 2419 3774
rect 2419 3745 2421 3774
rect 2437 3745 2453 3774
rect 2453 3745 2489 3774
rect 2505 3745 2557 3797
rect 2573 3745 2625 3797
rect 2641 3774 2693 3797
rect 2641 3745 2655 3774
rect 2655 3745 2689 3774
rect 2689 3745 2693 3774
rect 697 3681 749 3733
rect 765 3700 817 3733
rect 765 3681 767 3700
rect 767 3681 801 3700
rect 801 3681 817 3700
rect 833 3681 885 3733
rect 901 3681 953 3733
rect 969 3700 1021 3733
rect 969 3681 1003 3700
rect 1003 3681 1021 3700
rect 1037 3681 1089 3733
rect 1105 3681 1157 3733
rect 1173 3681 1225 3733
rect 1241 3700 1293 3733
rect 1241 3681 1273 3700
rect 1273 3681 1293 3700
rect 697 3617 749 3669
rect 765 3666 767 3669
rect 767 3666 801 3669
rect 801 3666 817 3669
rect 765 3626 817 3666
rect 765 3617 767 3626
rect 767 3617 801 3626
rect 801 3617 817 3626
rect 833 3617 885 3669
rect 901 3617 953 3669
rect 969 3666 1003 3669
rect 1003 3666 1021 3669
rect 969 3626 1021 3666
rect 969 3617 1003 3626
rect 1003 3617 1021 3626
rect 1037 3617 1089 3669
rect 1105 3617 1157 3669
rect 1173 3617 1225 3669
rect 1241 3666 1273 3669
rect 1273 3666 1293 3669
rect 2097 3681 2149 3733
rect 2165 3700 2217 3733
rect 2165 3681 2183 3700
rect 2183 3681 2217 3700
rect 2233 3681 2285 3733
rect 2301 3681 2353 3733
rect 2369 3700 2421 3733
rect 2437 3700 2489 3733
rect 2369 3681 2419 3700
rect 2419 3681 2421 3700
rect 2437 3681 2453 3700
rect 2453 3681 2489 3700
rect 2505 3681 2557 3733
rect 2573 3681 2625 3733
rect 2641 3700 2693 3733
rect 2641 3681 2655 3700
rect 2655 3681 2689 3700
rect 2689 3681 2693 3700
rect 1241 3626 1293 3666
rect 1241 3617 1273 3626
rect 1273 3617 1293 3626
rect 697 3553 749 3605
rect 765 3592 767 3605
rect 767 3592 801 3605
rect 801 3592 817 3605
rect 765 3553 817 3592
rect 833 3553 885 3605
rect 901 3553 953 3605
rect 969 3592 1003 3605
rect 1003 3592 1021 3605
rect 969 3553 1021 3592
rect 1037 3553 1089 3605
rect 1105 3553 1157 3605
rect 1173 3553 1225 3605
rect 1241 3592 1273 3605
rect 1273 3592 1293 3605
rect 2097 3617 2149 3669
rect 2165 3666 2183 3669
rect 2183 3666 2217 3669
rect 2165 3626 2217 3666
rect 2165 3617 2183 3626
rect 2183 3617 2217 3626
rect 2233 3617 2285 3669
rect 2301 3617 2353 3669
rect 2369 3666 2419 3669
rect 2419 3666 2421 3669
rect 2437 3666 2453 3669
rect 2453 3666 2489 3669
rect 2369 3626 2421 3666
rect 2437 3626 2489 3666
rect 2369 3617 2419 3626
rect 2419 3617 2421 3626
rect 2437 3617 2453 3626
rect 2453 3617 2489 3626
rect 2505 3617 2557 3669
rect 2573 3617 2625 3669
rect 2641 3666 2655 3669
rect 2655 3666 2689 3669
rect 2689 3666 2693 3669
rect 2641 3626 2693 3666
rect 2641 3617 2655 3626
rect 2655 3617 2689 3626
rect 2689 3617 2693 3626
rect 1241 3553 1293 3592
rect 2097 3553 2149 3605
rect 2165 3592 2183 3605
rect 2183 3592 2217 3605
rect 2165 3553 2217 3592
rect 2233 3553 2285 3605
rect 2301 3553 2353 3605
rect 2369 3592 2419 3605
rect 2419 3592 2421 3605
rect 2437 3592 2453 3605
rect 2453 3592 2489 3605
rect 2369 3553 2421 3592
rect 2437 3553 2489 3592
rect 2505 3553 2557 3605
rect 2573 3553 2625 3605
rect 2641 3592 2655 3605
rect 2655 3592 2689 3605
rect 2689 3592 2693 3605
rect 2641 3553 2693 3592
rect 697 3489 749 3541
rect 765 3518 767 3541
rect 767 3518 801 3541
rect 801 3518 817 3541
rect 765 3489 817 3518
rect 833 3489 885 3541
rect 901 3489 953 3541
rect 969 3518 1003 3541
rect 1003 3518 1021 3541
rect 969 3489 1021 3518
rect 1037 3489 1089 3541
rect 1105 3489 1157 3541
rect 1173 3489 1225 3541
rect 1241 3518 1273 3541
rect 1273 3518 1293 3541
rect 1241 3489 1293 3518
rect 2097 3489 2149 3541
rect 2165 3518 2183 3541
rect 2183 3518 2217 3541
rect 2165 3489 2217 3518
rect 2233 3489 2285 3541
rect 2301 3489 2353 3541
rect 2369 3518 2419 3541
rect 2419 3518 2421 3541
rect 2437 3518 2453 3541
rect 2453 3518 2489 3541
rect 2369 3489 2421 3518
rect 2437 3489 2489 3518
rect 2505 3489 2557 3541
rect 2573 3489 2625 3541
rect 2641 3518 2655 3541
rect 2655 3518 2689 3541
rect 2689 3518 2693 3541
rect 2641 3489 2693 3518
rect 1501 2844 1553 2853
rect 1569 2844 1621 2853
rect 1636 2844 1688 2853
rect 1703 2844 1755 2853
rect 1770 2844 1822 2853
rect 1837 2844 1889 2853
rect 1501 2810 1525 2844
rect 1525 2810 1553 2844
rect 1569 2810 1600 2844
rect 1600 2810 1621 2844
rect 1636 2810 1674 2844
rect 1674 2810 1688 2844
rect 1703 2810 1708 2844
rect 1708 2810 1748 2844
rect 1748 2810 1755 2844
rect 1770 2810 1782 2844
rect 1782 2810 1822 2844
rect 1837 2810 1856 2844
rect 1856 2810 1889 2844
rect 1501 2801 1553 2810
rect 1569 2801 1621 2810
rect 1636 2801 1688 2810
rect 1703 2801 1755 2810
rect 1770 2801 1822 2810
rect 1837 2801 1889 2810
rect 697 2191 749 2243
rect 765 2209 817 2243
rect 765 2191 767 2209
rect 767 2191 801 2209
rect 801 2191 817 2209
rect 833 2191 885 2243
rect 901 2191 953 2243
rect 969 2209 1021 2243
rect 969 2191 1003 2209
rect 1003 2191 1021 2209
rect 1037 2191 1089 2243
rect 1105 2191 1157 2243
rect 1173 2191 1225 2243
rect 1241 2209 1293 2243
rect 1241 2191 1273 2209
rect 1273 2191 1293 2209
rect 697 2127 749 2179
rect 765 2175 767 2179
rect 767 2175 801 2179
rect 801 2175 817 2179
rect 765 2136 817 2175
rect 765 2127 767 2136
rect 767 2127 801 2136
rect 801 2127 817 2136
rect 833 2127 885 2179
rect 901 2127 953 2179
rect 969 2175 1003 2179
rect 1003 2175 1021 2179
rect 969 2136 1021 2175
rect 969 2127 1003 2136
rect 1003 2127 1021 2136
rect 1037 2127 1089 2179
rect 1105 2127 1157 2179
rect 1173 2127 1225 2179
rect 1241 2175 1273 2179
rect 1273 2175 1293 2179
rect 2097 2191 2149 2243
rect 2165 2209 2217 2243
rect 2165 2191 2183 2209
rect 2183 2191 2217 2209
rect 2233 2191 2285 2243
rect 2301 2191 2353 2243
rect 2369 2209 2421 2243
rect 2437 2209 2489 2243
rect 2369 2191 2419 2209
rect 2419 2191 2421 2209
rect 2437 2191 2453 2209
rect 2453 2191 2489 2209
rect 2505 2191 2557 2243
rect 2573 2191 2625 2243
rect 2641 2209 2693 2243
rect 2641 2191 2655 2209
rect 2655 2191 2689 2209
rect 2689 2191 2693 2209
rect 1241 2136 1293 2175
rect 1241 2127 1273 2136
rect 1273 2127 1293 2136
rect 697 2063 749 2115
rect 765 2102 767 2115
rect 767 2102 801 2115
rect 801 2102 817 2115
rect 765 2063 817 2102
rect 833 2063 885 2115
rect 901 2063 953 2115
rect 969 2102 1003 2115
rect 1003 2102 1021 2115
rect 969 2063 1021 2102
rect 1037 2063 1089 2115
rect 1105 2063 1157 2115
rect 1173 2063 1225 2115
rect 1241 2102 1273 2115
rect 1273 2102 1293 2115
rect 2097 2127 2149 2179
rect 2165 2175 2183 2179
rect 2183 2175 2217 2179
rect 2165 2136 2217 2175
rect 2165 2127 2183 2136
rect 2183 2127 2217 2136
rect 2233 2127 2285 2179
rect 2301 2127 2353 2179
rect 2369 2175 2419 2179
rect 2419 2175 2421 2179
rect 2437 2175 2453 2179
rect 2453 2175 2489 2179
rect 2369 2136 2421 2175
rect 2437 2136 2489 2175
rect 2369 2127 2419 2136
rect 2419 2127 2421 2136
rect 2437 2127 2453 2136
rect 2453 2127 2489 2136
rect 2505 2127 2557 2179
rect 2573 2127 2625 2179
rect 2641 2175 2655 2179
rect 2655 2175 2689 2179
rect 2689 2175 2693 2179
rect 2641 2136 2693 2175
rect 2641 2127 2655 2136
rect 2655 2127 2689 2136
rect 2689 2127 2693 2136
rect 1241 2063 1293 2102
rect 2097 2063 2149 2115
rect 2165 2102 2183 2115
rect 2183 2102 2217 2115
rect 2165 2063 2217 2102
rect 2233 2063 2285 2115
rect 2301 2063 2353 2115
rect 2369 2102 2419 2115
rect 2419 2102 2421 2115
rect 2437 2102 2453 2115
rect 2453 2102 2489 2115
rect 2369 2063 2421 2102
rect 2437 2063 2489 2102
rect 2505 2063 2557 2115
rect 2573 2063 2625 2115
rect 2641 2102 2655 2115
rect 2655 2102 2689 2115
rect 2689 2102 2693 2115
rect 2641 2063 2693 2102
rect 697 1999 749 2051
rect 765 2029 767 2051
rect 767 2029 801 2051
rect 801 2029 817 2051
rect 765 1999 817 2029
rect 833 1999 885 2051
rect 901 1999 953 2051
rect 969 2029 1003 2051
rect 1003 2029 1021 2051
rect 969 1999 1021 2029
rect 1037 1999 1089 2051
rect 1105 1999 1157 2051
rect 1173 1999 1225 2051
rect 1241 2029 1273 2051
rect 1273 2029 1293 2051
rect 1241 1999 1293 2029
rect 2097 1999 2149 2051
rect 2165 2029 2183 2051
rect 2183 2029 2217 2051
rect 2165 1999 2217 2029
rect 2233 1999 2285 2051
rect 2301 1999 2353 2051
rect 2369 2029 2419 2051
rect 2419 2029 2421 2051
rect 2437 2029 2453 2051
rect 2453 2029 2489 2051
rect 2369 1999 2421 2029
rect 2437 1999 2489 2029
rect 2505 1999 2557 2051
rect 2573 1999 2625 2051
rect 2641 2029 2655 2051
rect 2655 2029 2689 2051
rect 2689 2029 2693 2051
rect 2641 1999 2693 2029
rect 697 1935 749 1987
rect 765 1956 767 1987
rect 767 1956 801 1987
rect 801 1956 817 1987
rect 765 1935 817 1956
rect 833 1935 885 1987
rect 901 1935 953 1987
rect 969 1956 1003 1987
rect 1003 1956 1021 1987
rect 969 1935 1021 1956
rect 1037 1935 1089 1987
rect 1105 1935 1157 1987
rect 1173 1935 1225 1987
rect 1241 1956 1273 1987
rect 1273 1956 1293 1987
rect 1241 1935 1293 1956
rect 2097 1935 2149 1987
rect 2165 1956 2183 1987
rect 2183 1956 2217 1987
rect 2165 1935 2217 1956
rect 2233 1935 2285 1987
rect 2301 1935 2353 1987
rect 2369 1956 2419 1987
rect 2419 1956 2421 1987
rect 2437 1956 2453 1987
rect 2453 1956 2489 1987
rect 2369 1935 2421 1956
rect 2437 1935 2489 1956
rect 2505 1935 2557 1987
rect 2573 1935 2625 1987
rect 2641 1956 2655 1987
rect 2655 1956 2689 1987
rect 2689 1956 2693 1987
rect 2641 1935 2693 1956
rect 697 1871 749 1923
rect 765 1917 817 1923
rect 765 1883 767 1917
rect 767 1883 801 1917
rect 801 1883 817 1917
rect 765 1871 817 1883
rect 833 1871 885 1923
rect 901 1871 953 1923
rect 969 1917 1021 1923
rect 969 1883 1003 1917
rect 1003 1883 1021 1917
rect 969 1871 1021 1883
rect 1037 1871 1089 1923
rect 1105 1871 1157 1923
rect 1173 1871 1225 1923
rect 1241 1917 1293 1923
rect 1241 1883 1273 1917
rect 1273 1883 1293 1917
rect 1241 1871 1293 1883
rect 2097 1871 2149 1923
rect 2165 1917 2217 1923
rect 2165 1883 2183 1917
rect 2183 1883 2217 1917
rect 2165 1871 2217 1883
rect 2233 1871 2285 1923
rect 2301 1871 2353 1923
rect 2369 1917 2421 1923
rect 2437 1917 2489 1923
rect 2369 1883 2419 1917
rect 2419 1883 2421 1917
rect 2437 1883 2453 1917
rect 2453 1883 2489 1917
rect 2369 1871 2421 1883
rect 2437 1871 2489 1883
rect 2505 1871 2557 1923
rect 2573 1871 2625 1923
rect 2641 1917 2693 1923
rect 2641 1883 2655 1917
rect 2655 1883 2689 1917
rect 2689 1883 2693 1917
rect 2641 1871 2693 1883
rect 697 1807 749 1859
rect 765 1844 817 1859
rect 765 1810 767 1844
rect 767 1810 801 1844
rect 801 1810 817 1844
rect 765 1807 817 1810
rect 833 1807 885 1859
rect 901 1807 953 1859
rect 969 1844 1021 1859
rect 969 1810 1003 1844
rect 1003 1810 1021 1844
rect 969 1807 1021 1810
rect 1037 1807 1089 1859
rect 1105 1807 1157 1859
rect 1173 1807 1225 1859
rect 1241 1844 1293 1859
rect 1241 1810 1273 1844
rect 1273 1810 1293 1844
rect 1241 1807 1293 1810
rect 2097 1807 2149 1859
rect 2165 1844 2217 1859
rect 2165 1810 2183 1844
rect 2183 1810 2217 1844
rect 2165 1807 2217 1810
rect 2233 1807 2285 1859
rect 2301 1807 2353 1859
rect 2369 1844 2421 1859
rect 2437 1844 2489 1859
rect 2369 1810 2419 1844
rect 2419 1810 2421 1844
rect 2437 1810 2453 1844
rect 2453 1810 2489 1844
rect 2369 1807 2421 1810
rect 2437 1807 2489 1810
rect 2505 1807 2557 1859
rect 2573 1807 2625 1859
rect 2641 1844 2693 1859
rect 2641 1810 2655 1844
rect 2655 1810 2689 1844
rect 2689 1810 2693 1844
rect 2641 1807 2693 1810
rect 697 1743 749 1795
rect 765 1770 817 1795
rect 765 1743 767 1770
rect 767 1743 801 1770
rect 801 1743 817 1770
rect 833 1743 885 1795
rect 901 1743 953 1795
rect 969 1770 1021 1795
rect 969 1743 1003 1770
rect 1003 1743 1021 1770
rect 1037 1743 1089 1795
rect 1105 1743 1157 1795
rect 1173 1743 1225 1795
rect 1241 1770 1293 1795
rect 1241 1743 1273 1770
rect 1273 1743 1293 1770
rect 2097 1743 2149 1795
rect 2165 1770 2217 1795
rect 2165 1743 2183 1770
rect 2183 1743 2217 1770
rect 2233 1743 2285 1795
rect 2301 1743 2353 1795
rect 2369 1770 2421 1795
rect 2437 1770 2489 1795
rect 2369 1743 2419 1770
rect 2419 1743 2421 1770
rect 2437 1743 2453 1770
rect 2453 1743 2489 1770
rect 2505 1743 2557 1795
rect 2573 1743 2625 1795
rect 2641 1770 2693 1795
rect 2641 1743 2655 1770
rect 2655 1743 2689 1770
rect 2689 1743 2693 1770
rect 697 1679 749 1731
rect 765 1696 817 1731
rect 765 1679 767 1696
rect 767 1679 801 1696
rect 801 1679 817 1696
rect 833 1679 885 1731
rect 901 1679 953 1731
rect 969 1696 1021 1731
rect 969 1679 1003 1696
rect 1003 1679 1021 1696
rect 1037 1679 1089 1731
rect 1105 1679 1157 1731
rect 1173 1679 1225 1731
rect 1241 1696 1293 1731
rect 1241 1679 1273 1696
rect 1273 1679 1293 1696
rect 697 1615 749 1667
rect 765 1662 767 1667
rect 767 1662 801 1667
rect 801 1662 817 1667
rect 765 1622 817 1662
rect 765 1615 767 1622
rect 767 1615 801 1622
rect 801 1615 817 1622
rect 833 1615 885 1667
rect 901 1615 953 1667
rect 969 1662 1003 1667
rect 1003 1662 1021 1667
rect 969 1622 1021 1662
rect 969 1615 1003 1622
rect 1003 1615 1021 1622
rect 1037 1615 1089 1667
rect 1105 1615 1157 1667
rect 1173 1615 1225 1667
rect 1241 1662 1273 1667
rect 1273 1662 1293 1667
rect 2097 1679 2149 1731
rect 2165 1696 2217 1731
rect 2165 1679 2183 1696
rect 2183 1679 2217 1696
rect 2233 1679 2285 1731
rect 2301 1679 2353 1731
rect 2369 1696 2421 1731
rect 2437 1696 2489 1731
rect 2369 1679 2419 1696
rect 2419 1679 2421 1696
rect 2437 1679 2453 1696
rect 2453 1679 2489 1696
rect 2505 1679 2557 1731
rect 2573 1679 2625 1731
rect 2641 1696 2693 1731
rect 2641 1679 2655 1696
rect 2655 1679 2689 1696
rect 2689 1679 2693 1696
rect 1241 1622 1293 1662
rect 1241 1615 1273 1622
rect 1273 1615 1293 1622
rect 697 1551 749 1603
rect 765 1588 767 1603
rect 767 1588 801 1603
rect 801 1588 817 1603
rect 765 1551 817 1588
rect 833 1551 885 1603
rect 901 1551 953 1603
rect 969 1588 1003 1603
rect 1003 1588 1021 1603
rect 969 1551 1021 1588
rect 1037 1551 1089 1603
rect 1105 1551 1157 1603
rect 1173 1551 1225 1603
rect 1241 1588 1273 1603
rect 1273 1588 1293 1603
rect 2097 1615 2149 1667
rect 2165 1662 2183 1667
rect 2183 1662 2217 1667
rect 2165 1622 2217 1662
rect 2165 1615 2183 1622
rect 2183 1615 2217 1622
rect 2233 1615 2285 1667
rect 2301 1615 2353 1667
rect 2369 1662 2419 1667
rect 2419 1662 2421 1667
rect 2437 1662 2453 1667
rect 2453 1662 2489 1667
rect 2369 1622 2421 1662
rect 2437 1622 2489 1662
rect 2369 1615 2419 1622
rect 2419 1615 2421 1622
rect 2437 1615 2453 1622
rect 2453 1615 2489 1622
rect 2505 1615 2557 1667
rect 2573 1615 2625 1667
rect 2641 1662 2655 1667
rect 2655 1662 2689 1667
rect 2689 1662 2693 1667
rect 2641 1622 2693 1662
rect 2641 1615 2655 1622
rect 2655 1615 2689 1622
rect 2689 1615 2693 1622
rect 1241 1551 1293 1588
rect 2097 1551 2149 1603
rect 2165 1588 2183 1603
rect 2183 1588 2217 1603
rect 2165 1551 2217 1588
rect 2233 1551 2285 1603
rect 2301 1551 2353 1603
rect 2369 1588 2419 1603
rect 2419 1588 2421 1603
rect 2437 1588 2453 1603
rect 2453 1588 2489 1603
rect 2369 1551 2421 1588
rect 2437 1551 2489 1588
rect 2505 1551 2557 1603
rect 2573 1551 2625 1603
rect 2641 1588 2655 1603
rect 2655 1588 2689 1603
rect 2689 1588 2693 1603
rect 2641 1551 2693 1588
rect 697 1487 749 1539
rect 765 1514 767 1539
rect 767 1514 801 1539
rect 801 1514 817 1539
rect 765 1487 817 1514
rect 833 1487 885 1539
rect 901 1487 953 1539
rect 969 1514 1003 1539
rect 1003 1514 1021 1539
rect 969 1487 1021 1514
rect 1037 1487 1089 1539
rect 1105 1487 1157 1539
rect 1173 1487 1225 1539
rect 1241 1514 1273 1539
rect 1273 1514 1293 1539
rect 1241 1487 1293 1514
rect 2097 1487 2149 1539
rect 2165 1514 2183 1539
rect 2183 1514 2217 1539
rect 2165 1487 2217 1514
rect 2233 1487 2285 1539
rect 2301 1487 2353 1539
rect 2369 1514 2419 1539
rect 2419 1514 2421 1539
rect 2437 1514 2453 1539
rect 2453 1514 2489 1539
rect 2369 1487 2421 1514
rect 2437 1487 2489 1514
rect 2505 1487 2557 1539
rect 2573 1487 2625 1539
rect 2641 1514 2655 1539
rect 2655 1514 2689 1539
rect 2689 1514 2693 1539
rect 2641 1487 2693 1514
rect 697 1423 749 1475
rect 765 1474 817 1475
rect 765 1440 767 1474
rect 767 1440 801 1474
rect 801 1440 817 1474
rect 765 1423 817 1440
rect 833 1423 885 1475
rect 901 1423 953 1475
rect 969 1474 1021 1475
rect 969 1440 1003 1474
rect 1003 1440 1021 1474
rect 969 1423 1021 1440
rect 1037 1423 1089 1475
rect 1105 1423 1157 1475
rect 1173 1423 1225 1475
rect 1241 1474 1293 1475
rect 1241 1440 1273 1474
rect 1273 1440 1293 1474
rect 1241 1423 1293 1440
rect 2097 1423 2149 1475
rect 2165 1474 2217 1475
rect 2165 1440 2183 1474
rect 2183 1440 2217 1474
rect 2165 1423 2217 1440
rect 2233 1423 2285 1475
rect 2301 1423 2353 1475
rect 2369 1474 2421 1475
rect 2437 1474 2489 1475
rect 2369 1440 2419 1474
rect 2419 1440 2421 1474
rect 2437 1440 2453 1474
rect 2453 1440 2489 1474
rect 2369 1423 2421 1440
rect 2437 1423 2489 1440
rect 2505 1423 2557 1475
rect 2573 1423 2625 1475
rect 2641 1474 2693 1475
rect 2641 1440 2655 1474
rect 2655 1440 2689 1474
rect 2689 1440 2693 1474
rect 2641 1423 2693 1440
rect 697 1359 749 1411
rect 765 1400 817 1411
rect 765 1366 767 1400
rect 767 1366 801 1400
rect 801 1366 817 1400
rect 765 1359 817 1366
rect 833 1359 885 1411
rect 901 1359 953 1411
rect 969 1400 1021 1411
rect 969 1366 1003 1400
rect 1003 1366 1021 1400
rect 969 1359 1021 1366
rect 1037 1359 1089 1411
rect 1105 1359 1157 1411
rect 1173 1359 1225 1411
rect 1241 1400 1293 1411
rect 1241 1366 1273 1400
rect 1273 1366 1293 1400
rect 1241 1359 1293 1366
rect 2097 1359 2149 1411
rect 2165 1400 2217 1411
rect 2165 1366 2183 1400
rect 2183 1366 2217 1400
rect 2165 1359 2217 1366
rect 2233 1359 2285 1411
rect 2301 1359 2353 1411
rect 2369 1400 2421 1411
rect 2437 1400 2489 1411
rect 2369 1366 2419 1400
rect 2419 1366 2421 1400
rect 2437 1366 2453 1400
rect 2453 1366 2489 1400
rect 2369 1359 2421 1366
rect 2437 1359 2489 1366
rect 2505 1359 2557 1411
rect 2573 1359 2625 1411
rect 2641 1400 2693 1411
rect 2641 1366 2655 1400
rect 2655 1366 2689 1400
rect 2689 1366 2693 1400
rect 2641 1359 2693 1366
rect 697 1295 749 1347
rect 765 1326 817 1347
rect 765 1295 767 1326
rect 767 1295 801 1326
rect 801 1295 817 1326
rect 833 1295 885 1347
rect 901 1295 953 1347
rect 969 1326 1021 1347
rect 969 1295 1003 1326
rect 1003 1295 1021 1326
rect 1037 1295 1089 1347
rect 1105 1295 1157 1347
rect 1173 1295 1225 1347
rect 1241 1326 1293 1347
rect 1241 1295 1273 1326
rect 1273 1295 1293 1326
rect 2097 1295 2149 1347
rect 2165 1326 2217 1347
rect 2165 1295 2183 1326
rect 2183 1295 2217 1326
rect 2233 1295 2285 1347
rect 2301 1295 2353 1347
rect 2369 1326 2421 1347
rect 2437 1326 2489 1347
rect 2369 1295 2419 1326
rect 2419 1295 2421 1326
rect 2437 1295 2453 1326
rect 2453 1295 2489 1326
rect 2505 1295 2557 1347
rect 2573 1295 2625 1347
rect 2641 1326 2693 1347
rect 2641 1295 2655 1326
rect 2655 1295 2689 1326
rect 2689 1295 2693 1326
rect 1501 714 1553 723
rect 1569 714 1621 723
rect 1636 714 1688 723
rect 1703 714 1755 723
rect 1770 714 1822 723
rect 1837 714 1889 723
rect 1501 680 1525 714
rect 1525 680 1553 714
rect 1569 680 1600 714
rect 1600 680 1621 714
rect 1636 680 1674 714
rect 1674 680 1688 714
rect 1703 680 1708 714
rect 1708 680 1748 714
rect 1748 680 1755 714
rect 1770 680 1782 714
rect 1782 680 1822 714
rect 1837 680 1856 714
rect 1856 680 1889 714
rect 1501 671 1553 680
rect 1569 671 1621 680
rect 1636 671 1688 680
rect 1703 671 1755 680
rect 1770 671 1822 680
rect 1837 671 1889 680
rect 3287 13666 3339 13701
rect 3287 13649 3296 13666
rect 3296 13649 3330 13666
rect 3330 13649 3339 13666
rect 3287 13632 3296 13633
rect 3296 13632 3330 13633
rect 3330 13632 3339 13633
rect 3287 13594 3339 13632
rect 3287 13581 3296 13594
rect 3296 13581 3330 13594
rect 3330 13581 3339 13594
rect 3287 13560 3296 13565
rect 3296 13560 3330 13565
rect 3330 13560 3339 13565
rect 3287 13522 3339 13560
rect 3287 13513 3296 13522
rect 3296 13513 3330 13522
rect 3330 13513 3339 13522
rect 3287 13488 3296 13496
rect 3296 13488 3330 13496
rect 3330 13488 3339 13496
rect 3287 13450 3339 13488
rect 3287 13444 3296 13450
rect 3296 13444 3330 13450
rect 3330 13444 3339 13450
rect 3287 13416 3296 13427
rect 3296 13416 3330 13427
rect 3330 13416 3339 13427
rect 3287 13378 3339 13416
rect 3287 13375 3296 13378
rect 3296 13375 3330 13378
rect 3330 13375 3339 13378
rect 3287 13344 3296 13358
rect 3296 13344 3330 13358
rect 3330 13344 3339 13358
rect 3287 13306 3339 13344
rect 3287 13272 3296 13289
rect 3296 13272 3330 13289
rect 3330 13272 3339 13289
rect 3287 13237 3339 13272
rect 3287 13200 3296 13220
rect 3296 13200 3330 13220
rect 3330 13200 3339 13220
rect 3287 13168 3339 13200
rect 3287 13128 3296 13151
rect 3296 13128 3330 13151
rect 3330 13128 3339 13151
rect 3287 13099 3339 13128
rect 3287 13056 3296 13082
rect 3296 13056 3330 13082
rect 3330 13056 3339 13082
rect 3287 13030 3339 13056
rect 3287 12984 3296 13013
rect 3296 12984 3330 13013
rect 3330 12984 3339 13013
rect 3287 12961 3339 12984
rect 3287 12912 3296 12944
rect 3296 12912 3330 12944
rect 3330 12912 3339 12944
rect 3287 12892 3339 12912
rect 3287 12874 3339 12875
rect 3287 12840 3296 12874
rect 3296 12840 3330 12874
rect 3330 12840 3339 12874
rect 3287 12823 3339 12840
<< metal2 >>
rect 695 39341 2695 39782
rect 695 38423 1295 39341
tri 1295 39165 1471 39341 nw
tri 1919 39165 2095 39341 ne
rect 695 38371 697 38423
rect 749 38420 765 38423
rect 817 38420 833 38423
rect 885 38420 901 38423
rect 953 38420 969 38423
rect 1021 38420 1037 38423
rect 1089 38420 1105 38423
rect 1157 38420 1173 38423
rect 1225 38420 1241 38423
rect 1293 38371 1295 38423
rect 695 38359 727 38371
rect 1263 38359 1295 38371
rect 695 38307 697 38359
rect 1293 38307 1295 38359
rect 695 38295 727 38307
rect 1263 38295 1295 38307
rect 695 38243 697 38295
rect 1293 38243 1295 38295
rect 695 38231 727 38243
rect 1263 38231 1295 38243
rect 695 38179 697 38231
rect 1293 38179 1295 38231
rect 695 38167 727 38179
rect 1263 38167 1295 38179
rect 695 38115 697 38167
rect 1293 38115 1295 38167
rect 695 38103 727 38115
rect 1263 38103 1295 38115
rect 695 38051 697 38103
rect 1293 38051 1295 38103
rect 695 38039 727 38051
rect 1263 38039 1295 38051
rect 695 37987 697 38039
rect 1293 37987 1295 38039
rect 695 37975 727 37987
rect 1263 37975 1295 37987
rect 695 37923 697 37975
rect 749 37939 765 37964
rect 817 37939 833 37964
rect 885 37939 901 37964
rect 953 37939 969 37964
rect 1021 37939 1037 37964
rect 1089 37939 1105 37964
rect 1157 37939 1173 37964
rect 1225 37939 1241 37964
rect 885 37923 887 37939
rect 953 37923 967 37939
rect 1023 37923 1037 37939
rect 1103 37923 1105 37939
rect 1293 37923 1295 37975
rect 695 37911 727 37923
rect 783 37911 807 37923
rect 863 37911 887 37923
rect 943 37911 967 37923
rect 1023 37911 1047 37923
rect 1103 37911 1127 37923
rect 1183 37911 1207 37923
rect 1263 37911 1295 37923
rect 695 37859 697 37911
rect 885 37883 887 37911
rect 953 37883 967 37911
rect 1023 37883 1037 37911
rect 1103 37883 1105 37911
rect 749 37859 765 37883
rect 817 37859 833 37883
rect 885 37859 901 37883
rect 953 37859 969 37883
rect 1021 37859 1037 37883
rect 1089 37859 1105 37883
rect 1157 37859 1173 37883
rect 1225 37859 1241 37883
rect 1293 37859 1295 37911
rect 695 37858 1295 37859
rect 695 37847 727 37858
rect 783 37847 807 37858
rect 863 37847 887 37858
rect 943 37847 967 37858
rect 1023 37847 1047 37858
rect 1103 37847 1127 37858
rect 1183 37847 1207 37858
rect 1263 37847 1295 37858
rect 695 37795 697 37847
rect 885 37802 887 37847
rect 953 37802 967 37847
rect 1023 37802 1037 37847
rect 1103 37802 1105 37847
rect 749 37795 765 37802
rect 817 37795 833 37802
rect 885 37795 901 37802
rect 953 37795 969 37802
rect 1021 37795 1037 37802
rect 1089 37795 1105 37802
rect 1157 37795 1173 37802
rect 1225 37795 1241 37802
rect 1293 37795 1295 37847
rect 695 37783 1295 37795
rect 695 37731 697 37783
rect 749 37777 765 37783
rect 817 37777 833 37783
rect 885 37777 901 37783
rect 953 37777 969 37783
rect 1021 37777 1037 37783
rect 1089 37777 1105 37783
rect 1157 37777 1173 37783
rect 1225 37777 1241 37783
rect 885 37731 887 37777
rect 953 37731 967 37777
rect 1023 37731 1037 37777
rect 1103 37731 1105 37777
rect 1293 37731 1295 37783
rect 695 37721 727 37731
rect 783 37721 807 37731
rect 863 37721 887 37731
rect 943 37721 967 37731
rect 1023 37721 1047 37731
rect 1103 37721 1127 37731
rect 1183 37721 1207 37731
rect 1263 37721 1295 37731
rect 695 37719 1295 37721
rect 695 37667 697 37719
rect 749 37696 765 37719
rect 817 37696 833 37719
rect 885 37696 901 37719
rect 953 37696 969 37719
rect 1021 37696 1037 37719
rect 1089 37696 1105 37719
rect 1157 37696 1173 37719
rect 1225 37696 1241 37719
rect 885 37667 887 37696
rect 953 37667 967 37696
rect 1023 37667 1037 37696
rect 1103 37667 1105 37696
rect 1293 37667 1295 37719
rect 695 37655 727 37667
rect 783 37655 807 37667
rect 863 37655 887 37667
rect 943 37655 967 37667
rect 1023 37655 1047 37667
rect 1103 37655 1127 37667
rect 1183 37655 1207 37667
rect 1263 37655 1295 37667
rect 695 37603 697 37655
rect 885 37640 887 37655
rect 953 37640 967 37655
rect 1023 37640 1037 37655
rect 1103 37640 1105 37655
rect 749 37615 765 37640
rect 817 37615 833 37640
rect 885 37615 901 37640
rect 953 37615 969 37640
rect 1021 37615 1037 37640
rect 1089 37615 1105 37640
rect 1157 37615 1173 37640
rect 1225 37615 1241 37640
rect 885 37603 887 37615
rect 953 37603 967 37615
rect 1023 37603 1037 37615
rect 1103 37603 1105 37615
rect 1293 37603 1295 37655
rect 695 37591 727 37603
rect 783 37591 807 37603
rect 863 37591 887 37603
rect 943 37591 967 37603
rect 1023 37591 1047 37603
rect 1103 37591 1127 37603
rect 1183 37591 1207 37603
rect 1263 37591 1295 37603
rect 695 37539 697 37591
rect 885 37559 887 37591
rect 953 37559 967 37591
rect 1023 37559 1037 37591
rect 1103 37559 1105 37591
rect 749 37539 765 37559
rect 817 37539 833 37559
rect 885 37539 901 37559
rect 953 37539 969 37559
rect 1021 37539 1037 37559
rect 1089 37539 1105 37559
rect 1157 37539 1173 37559
rect 1225 37539 1241 37559
rect 1293 37539 1295 37591
rect 695 37534 1295 37539
rect 695 37527 727 37534
rect 783 37527 807 37534
rect 863 37527 887 37534
rect 943 37527 967 37534
rect 1023 37527 1047 37534
rect 1103 37527 1127 37534
rect 1183 37527 1207 37534
rect 1263 37527 1295 37534
rect 695 37475 697 37527
rect 885 37478 887 37527
rect 953 37478 967 37527
rect 1023 37478 1037 37527
rect 1103 37478 1105 37527
rect 749 37475 765 37478
rect 817 37475 833 37478
rect 885 37475 901 37478
rect 953 37475 969 37478
rect 1021 37475 1037 37478
rect 1089 37475 1105 37478
rect 1157 37475 1173 37478
rect 1225 37475 1241 37478
rect 1293 37475 1295 37527
rect 695 36369 1295 37475
rect 695 36317 697 36369
rect 749 36366 765 36369
rect 817 36366 833 36369
rect 885 36366 901 36369
rect 953 36366 969 36369
rect 1021 36366 1037 36369
rect 1089 36366 1105 36369
rect 1157 36366 1173 36369
rect 1225 36366 1241 36369
rect 1293 36317 1295 36369
rect 695 36305 727 36317
rect 1263 36305 1295 36317
rect 695 36253 697 36305
rect 1293 36253 1295 36305
rect 695 36241 727 36253
rect 1263 36241 1295 36253
rect 695 36189 697 36241
rect 1293 36189 1295 36241
rect 695 36177 727 36189
rect 1263 36177 1295 36189
rect 695 36125 697 36177
rect 1293 36125 1295 36177
rect 695 36113 727 36125
rect 1263 36113 1295 36125
rect 695 36061 697 36113
rect 1293 36061 1295 36113
rect 695 36049 727 36061
rect 1263 36049 1295 36061
rect 695 35997 697 36049
rect 1293 35997 1295 36049
rect 695 35985 727 35997
rect 1263 35985 1295 35997
rect 695 35933 697 35985
rect 1293 35933 1295 35985
rect 695 35921 727 35933
rect 1263 35921 1295 35933
rect 695 35869 697 35921
rect 749 35885 765 35910
rect 817 35885 833 35910
rect 885 35885 901 35910
rect 953 35885 969 35910
rect 1021 35885 1037 35910
rect 1089 35885 1105 35910
rect 1157 35885 1173 35910
rect 1225 35885 1241 35910
rect 885 35869 887 35885
rect 953 35869 967 35885
rect 1023 35869 1037 35885
rect 1103 35869 1105 35885
rect 1293 35869 1295 35921
rect 695 35857 727 35869
rect 783 35857 807 35869
rect 863 35857 887 35869
rect 943 35857 967 35869
rect 1023 35857 1047 35869
rect 1103 35857 1127 35869
rect 1183 35857 1207 35869
rect 1263 35857 1295 35869
rect 695 35805 697 35857
rect 885 35829 887 35857
rect 953 35829 967 35857
rect 1023 35829 1037 35857
rect 1103 35829 1105 35857
rect 749 35805 765 35829
rect 817 35805 833 35829
rect 885 35805 901 35829
rect 953 35805 969 35829
rect 1021 35805 1037 35829
rect 1089 35805 1105 35829
rect 1157 35805 1173 35829
rect 1225 35805 1241 35829
rect 1293 35805 1295 35857
rect 695 35804 1295 35805
rect 695 35793 727 35804
rect 783 35793 807 35804
rect 863 35793 887 35804
rect 943 35793 967 35804
rect 1023 35793 1047 35804
rect 1103 35793 1127 35804
rect 1183 35793 1207 35804
rect 1263 35793 1295 35804
rect 695 35741 697 35793
rect 885 35748 887 35793
rect 953 35748 967 35793
rect 1023 35748 1037 35793
rect 1103 35748 1105 35793
rect 749 35741 765 35748
rect 817 35741 833 35748
rect 885 35741 901 35748
rect 953 35741 969 35748
rect 1021 35741 1037 35748
rect 1089 35741 1105 35748
rect 1157 35741 1173 35748
rect 1225 35741 1241 35748
rect 1293 35741 1295 35793
rect 695 35729 1295 35741
rect 695 35677 697 35729
rect 749 35723 765 35729
rect 817 35723 833 35729
rect 885 35723 901 35729
rect 953 35723 969 35729
rect 1021 35723 1037 35729
rect 1089 35723 1105 35729
rect 1157 35723 1173 35729
rect 1225 35723 1241 35729
rect 885 35677 887 35723
rect 953 35677 967 35723
rect 1023 35677 1037 35723
rect 1103 35677 1105 35723
rect 1293 35677 1295 35729
rect 695 35667 727 35677
rect 783 35667 807 35677
rect 863 35667 887 35677
rect 943 35667 967 35677
rect 1023 35667 1047 35677
rect 1103 35667 1127 35677
rect 1183 35667 1207 35677
rect 1263 35667 1295 35677
rect 695 35665 1295 35667
rect 695 35613 697 35665
rect 749 35642 765 35665
rect 817 35642 833 35665
rect 885 35642 901 35665
rect 953 35642 969 35665
rect 1021 35642 1037 35665
rect 1089 35642 1105 35665
rect 1157 35642 1173 35665
rect 1225 35642 1241 35665
rect 885 35613 887 35642
rect 953 35613 967 35642
rect 1023 35613 1037 35642
rect 1103 35613 1105 35642
rect 1293 35613 1295 35665
rect 695 35601 727 35613
rect 783 35601 807 35613
rect 863 35601 887 35613
rect 943 35601 967 35613
rect 1023 35601 1047 35613
rect 1103 35601 1127 35613
rect 1183 35601 1207 35613
rect 1263 35601 1295 35613
rect 695 35549 697 35601
rect 885 35586 887 35601
rect 953 35586 967 35601
rect 1023 35586 1037 35601
rect 1103 35586 1105 35601
rect 749 35561 765 35586
rect 817 35561 833 35586
rect 885 35561 901 35586
rect 953 35561 969 35586
rect 1021 35561 1037 35586
rect 1089 35561 1105 35586
rect 1157 35561 1173 35586
rect 1225 35561 1241 35586
rect 885 35549 887 35561
rect 953 35549 967 35561
rect 1023 35549 1037 35561
rect 1103 35549 1105 35561
rect 1293 35549 1295 35601
rect 695 35537 727 35549
rect 783 35537 807 35549
rect 863 35537 887 35549
rect 943 35537 967 35549
rect 1023 35537 1047 35549
rect 1103 35537 1127 35549
rect 1183 35537 1207 35549
rect 1263 35537 1295 35549
rect 695 35485 697 35537
rect 885 35505 887 35537
rect 953 35505 967 35537
rect 1023 35505 1037 35537
rect 1103 35505 1105 35537
rect 749 35485 765 35505
rect 817 35485 833 35505
rect 885 35485 901 35505
rect 953 35485 969 35505
rect 1021 35485 1037 35505
rect 1089 35485 1105 35505
rect 1157 35485 1173 35505
rect 1225 35485 1241 35505
rect 1293 35485 1295 35537
rect 695 35480 1295 35485
rect 695 35473 727 35480
rect 783 35473 807 35480
rect 863 35473 887 35480
rect 943 35473 967 35480
rect 1023 35473 1047 35480
rect 1103 35473 1127 35480
rect 1183 35473 1207 35480
rect 1263 35473 1295 35480
rect 695 35421 697 35473
rect 885 35424 887 35473
rect 953 35424 967 35473
rect 1023 35424 1037 35473
rect 1103 35424 1105 35473
rect 749 35421 765 35424
rect 817 35421 833 35424
rect 885 35421 901 35424
rect 953 35421 969 35424
rect 1021 35421 1037 35424
rect 1089 35421 1105 35424
rect 1157 35421 1173 35424
rect 1225 35421 1241 35424
rect 1293 35421 1295 35473
rect 695 34150 1295 35421
rect 695 34098 697 34150
rect 749 34147 765 34150
rect 817 34147 833 34150
rect 885 34147 901 34150
rect 953 34147 969 34150
rect 1021 34147 1037 34150
rect 1089 34147 1105 34150
rect 1157 34147 1173 34150
rect 1225 34147 1241 34150
rect 1293 34098 1295 34150
rect 695 34086 727 34098
rect 1263 34086 1295 34098
rect 695 34034 697 34086
rect 1293 34034 1295 34086
rect 695 34022 727 34034
rect 1263 34022 1295 34034
rect 695 33970 697 34022
rect 1293 33970 1295 34022
rect 695 33958 727 33970
rect 1263 33958 1295 33970
rect 695 33906 697 33958
rect 1293 33906 1295 33958
rect 695 33894 727 33906
rect 1263 33894 1295 33906
rect 695 33842 697 33894
rect 1293 33842 1295 33894
rect 695 33830 727 33842
rect 1263 33830 1295 33842
rect 695 33778 697 33830
rect 1293 33778 1295 33830
rect 695 33766 727 33778
rect 1263 33766 1295 33778
rect 695 33714 697 33766
rect 1293 33714 1295 33766
rect 695 33702 727 33714
rect 1263 33702 1295 33714
rect 695 33650 697 33702
rect 749 33666 765 33691
rect 817 33666 833 33691
rect 885 33666 901 33691
rect 953 33666 969 33691
rect 1021 33666 1037 33691
rect 1089 33666 1105 33691
rect 1157 33666 1173 33691
rect 1225 33666 1241 33691
rect 885 33650 887 33666
rect 953 33650 967 33666
rect 1023 33650 1037 33666
rect 1103 33650 1105 33666
rect 1293 33650 1295 33702
rect 695 33638 727 33650
rect 783 33638 807 33650
rect 863 33638 887 33650
rect 943 33638 967 33650
rect 1023 33638 1047 33650
rect 1103 33638 1127 33650
rect 1183 33638 1207 33650
rect 1263 33638 1295 33650
rect 695 33586 697 33638
rect 885 33610 887 33638
rect 953 33610 967 33638
rect 1023 33610 1037 33638
rect 1103 33610 1105 33638
rect 749 33586 765 33610
rect 817 33586 833 33610
rect 885 33586 901 33610
rect 953 33586 969 33610
rect 1021 33586 1037 33610
rect 1089 33586 1105 33610
rect 1157 33586 1173 33610
rect 1225 33586 1241 33610
rect 1293 33586 1295 33638
rect 695 33585 1295 33586
rect 695 33574 727 33585
rect 783 33574 807 33585
rect 863 33574 887 33585
rect 943 33574 967 33585
rect 1023 33574 1047 33585
rect 1103 33574 1127 33585
rect 1183 33574 1207 33585
rect 1263 33574 1295 33585
rect 695 33522 697 33574
rect 885 33529 887 33574
rect 953 33529 967 33574
rect 1023 33529 1037 33574
rect 1103 33529 1105 33574
rect 749 33522 765 33529
rect 817 33522 833 33529
rect 885 33522 901 33529
rect 953 33522 969 33529
rect 1021 33522 1037 33529
rect 1089 33522 1105 33529
rect 1157 33522 1173 33529
rect 1225 33522 1241 33529
rect 1293 33522 1295 33574
rect 695 33510 1295 33522
rect 695 33458 697 33510
rect 749 33504 765 33510
rect 817 33504 833 33510
rect 885 33504 901 33510
rect 953 33504 969 33510
rect 1021 33504 1037 33510
rect 1089 33504 1105 33510
rect 1157 33504 1173 33510
rect 1225 33504 1241 33510
rect 885 33458 887 33504
rect 953 33458 967 33504
rect 1023 33458 1037 33504
rect 1103 33458 1105 33504
rect 1293 33458 1295 33510
rect 695 33448 727 33458
rect 783 33448 807 33458
rect 863 33448 887 33458
rect 943 33448 967 33458
rect 1023 33448 1047 33458
rect 1103 33448 1127 33458
rect 1183 33448 1207 33458
rect 1263 33448 1295 33458
rect 695 33446 1295 33448
rect 695 33394 697 33446
rect 749 33423 765 33446
rect 817 33423 833 33446
rect 885 33423 901 33446
rect 953 33423 969 33446
rect 1021 33423 1037 33446
rect 1089 33423 1105 33446
rect 1157 33423 1173 33446
rect 1225 33423 1241 33446
rect 885 33394 887 33423
rect 953 33394 967 33423
rect 1023 33394 1037 33423
rect 1103 33394 1105 33423
rect 1293 33394 1295 33446
rect 695 33382 727 33394
rect 783 33382 807 33394
rect 863 33382 887 33394
rect 943 33382 967 33394
rect 1023 33382 1047 33394
rect 1103 33382 1127 33394
rect 1183 33382 1207 33394
rect 1263 33382 1295 33394
rect 695 33330 697 33382
rect 885 33367 887 33382
rect 953 33367 967 33382
rect 1023 33367 1037 33382
rect 1103 33367 1105 33382
rect 749 33342 765 33367
rect 817 33342 833 33367
rect 885 33342 901 33367
rect 953 33342 969 33367
rect 1021 33342 1037 33367
rect 1089 33342 1105 33367
rect 1157 33342 1173 33367
rect 1225 33342 1241 33367
rect 885 33330 887 33342
rect 953 33330 967 33342
rect 1023 33330 1037 33342
rect 1103 33330 1105 33342
rect 1293 33330 1295 33382
rect 695 33318 727 33330
rect 783 33318 807 33330
rect 863 33318 887 33330
rect 943 33318 967 33330
rect 1023 33318 1047 33330
rect 1103 33318 1127 33330
rect 1183 33318 1207 33330
rect 1263 33318 1295 33330
rect 695 33266 697 33318
rect 885 33286 887 33318
rect 953 33286 967 33318
rect 1023 33286 1037 33318
rect 1103 33286 1105 33318
rect 749 33266 765 33286
rect 817 33266 833 33286
rect 885 33266 901 33286
rect 953 33266 969 33286
rect 1021 33266 1037 33286
rect 1089 33266 1105 33286
rect 1157 33266 1173 33286
rect 1225 33266 1241 33286
rect 1293 33266 1295 33318
rect 695 33261 1295 33266
rect 695 33254 727 33261
rect 783 33254 807 33261
rect 863 33254 887 33261
rect 943 33254 967 33261
rect 1023 33254 1047 33261
rect 1103 33254 1127 33261
rect 1183 33254 1207 33261
rect 1263 33254 1295 33261
rect 695 33202 697 33254
rect 885 33205 887 33254
rect 953 33205 967 33254
rect 1023 33205 1037 33254
rect 1103 33205 1105 33254
rect 749 33202 765 33205
rect 817 33202 833 33205
rect 885 33202 901 33205
rect 953 33202 969 33205
rect 1021 33202 1037 33205
rect 1089 33202 1105 33205
rect 1157 33202 1173 33205
rect 1225 33202 1241 33205
rect 1293 33202 1295 33254
rect 695 32021 1295 33202
rect 695 31969 697 32021
rect 749 32018 765 32021
rect 817 32018 833 32021
rect 885 32018 901 32021
rect 953 32018 969 32021
rect 1021 32018 1037 32021
rect 1089 32018 1105 32021
rect 1157 32018 1173 32021
rect 1225 32018 1241 32021
rect 1293 31969 1295 32021
rect 695 31957 727 31969
rect 1263 31957 1295 31969
rect 695 31905 697 31957
rect 1293 31905 1295 31957
rect 695 31893 727 31905
rect 1263 31893 1295 31905
rect 695 31841 697 31893
rect 1293 31841 1295 31893
rect 695 31829 727 31841
rect 1263 31829 1295 31841
rect 695 31777 697 31829
rect 1293 31777 1295 31829
rect 695 31765 727 31777
rect 1263 31765 1295 31777
rect 695 31713 697 31765
rect 1293 31713 1295 31765
rect 695 31701 727 31713
rect 1263 31701 1295 31713
rect 695 31649 697 31701
rect 1293 31649 1295 31701
rect 695 31637 727 31649
rect 1263 31637 1295 31649
rect 695 31585 697 31637
rect 1293 31585 1295 31637
rect 695 31573 727 31585
rect 1263 31573 1295 31585
rect 695 31521 697 31573
rect 749 31537 765 31562
rect 817 31537 833 31562
rect 885 31537 901 31562
rect 953 31537 969 31562
rect 1021 31537 1037 31562
rect 1089 31537 1105 31562
rect 1157 31537 1173 31562
rect 1225 31537 1241 31562
rect 885 31521 887 31537
rect 953 31521 967 31537
rect 1023 31521 1037 31537
rect 1103 31521 1105 31537
rect 1293 31521 1295 31573
rect 695 31509 727 31521
rect 783 31509 807 31521
rect 863 31509 887 31521
rect 943 31509 967 31521
rect 1023 31509 1047 31521
rect 1103 31509 1127 31521
rect 1183 31509 1207 31521
rect 1263 31509 1295 31521
rect 695 31457 697 31509
rect 885 31481 887 31509
rect 953 31481 967 31509
rect 1023 31481 1037 31509
rect 1103 31481 1105 31509
rect 749 31457 765 31481
rect 817 31457 833 31481
rect 885 31457 901 31481
rect 953 31457 969 31481
rect 1021 31457 1037 31481
rect 1089 31457 1105 31481
rect 1157 31457 1173 31481
rect 1225 31457 1241 31481
rect 1293 31457 1295 31509
rect 695 31456 1295 31457
rect 695 31445 727 31456
rect 783 31445 807 31456
rect 863 31445 887 31456
rect 943 31445 967 31456
rect 1023 31445 1047 31456
rect 1103 31445 1127 31456
rect 1183 31445 1207 31456
rect 1263 31445 1295 31456
rect 695 31393 697 31445
rect 885 31400 887 31445
rect 953 31400 967 31445
rect 1023 31400 1037 31445
rect 1103 31400 1105 31445
rect 749 31393 765 31400
rect 817 31393 833 31400
rect 885 31393 901 31400
rect 953 31393 969 31400
rect 1021 31393 1037 31400
rect 1089 31393 1105 31400
rect 1157 31393 1173 31400
rect 1225 31393 1241 31400
rect 1293 31393 1295 31445
rect 695 31381 1295 31393
rect 695 31329 697 31381
rect 749 31375 765 31381
rect 817 31375 833 31381
rect 885 31375 901 31381
rect 953 31375 969 31381
rect 1021 31375 1037 31381
rect 1089 31375 1105 31381
rect 1157 31375 1173 31381
rect 1225 31375 1241 31381
rect 885 31329 887 31375
rect 953 31329 967 31375
rect 1023 31329 1037 31375
rect 1103 31329 1105 31375
rect 1293 31329 1295 31381
rect 695 31319 727 31329
rect 783 31319 807 31329
rect 863 31319 887 31329
rect 943 31319 967 31329
rect 1023 31319 1047 31329
rect 1103 31319 1127 31329
rect 1183 31319 1207 31329
rect 1263 31319 1295 31329
rect 695 31317 1295 31319
rect 695 31265 697 31317
rect 749 31294 765 31317
rect 817 31294 833 31317
rect 885 31294 901 31317
rect 953 31294 969 31317
rect 1021 31294 1037 31317
rect 1089 31294 1105 31317
rect 1157 31294 1173 31317
rect 1225 31294 1241 31317
rect 885 31265 887 31294
rect 953 31265 967 31294
rect 1023 31265 1037 31294
rect 1103 31265 1105 31294
rect 1293 31265 1295 31317
rect 695 31253 727 31265
rect 783 31253 807 31265
rect 863 31253 887 31265
rect 943 31253 967 31265
rect 1023 31253 1047 31265
rect 1103 31253 1127 31265
rect 1183 31253 1207 31265
rect 1263 31253 1295 31265
rect 695 31201 697 31253
rect 885 31238 887 31253
rect 953 31238 967 31253
rect 1023 31238 1037 31253
rect 1103 31238 1105 31253
rect 749 31213 765 31238
rect 817 31213 833 31238
rect 885 31213 901 31238
rect 953 31213 969 31238
rect 1021 31213 1037 31238
rect 1089 31213 1105 31238
rect 1157 31213 1173 31238
rect 1225 31213 1241 31238
rect 885 31201 887 31213
rect 953 31201 967 31213
rect 1023 31201 1037 31213
rect 1103 31201 1105 31213
rect 1293 31201 1295 31253
rect 695 31189 727 31201
rect 783 31189 807 31201
rect 863 31189 887 31201
rect 943 31189 967 31201
rect 1023 31189 1047 31201
rect 1103 31189 1127 31201
rect 1183 31189 1207 31201
rect 1263 31189 1295 31201
rect 695 31137 697 31189
rect 885 31157 887 31189
rect 953 31157 967 31189
rect 1023 31157 1037 31189
rect 1103 31157 1105 31189
rect 749 31137 765 31157
rect 817 31137 833 31157
rect 885 31137 901 31157
rect 953 31137 969 31157
rect 1021 31137 1037 31157
rect 1089 31137 1105 31157
rect 1157 31137 1173 31157
rect 1225 31137 1241 31157
rect 1293 31137 1295 31189
rect 695 31132 1295 31137
rect 695 31125 727 31132
rect 783 31125 807 31132
rect 863 31125 887 31132
rect 943 31125 967 31132
rect 1023 31125 1047 31132
rect 1103 31125 1127 31132
rect 1183 31125 1207 31132
rect 1263 31125 1295 31132
rect 695 31073 697 31125
rect 885 31076 887 31125
rect 953 31076 967 31125
rect 1023 31076 1037 31125
rect 1103 31076 1105 31125
rect 749 31073 765 31076
rect 817 31073 833 31076
rect 885 31073 901 31076
rect 953 31073 969 31076
rect 1021 31073 1037 31076
rect 1089 31073 1105 31076
rect 1157 31073 1173 31076
rect 1225 31073 1241 31076
rect 1293 31073 1295 31125
rect 695 29872 1295 31073
rect 695 29820 697 29872
rect 749 29869 765 29872
rect 817 29869 833 29872
rect 885 29869 901 29872
rect 953 29869 969 29872
rect 1021 29869 1037 29872
rect 1089 29869 1105 29872
rect 1157 29869 1173 29872
rect 1225 29869 1241 29872
rect 1293 29820 1295 29872
rect 695 29808 727 29820
rect 1263 29808 1295 29820
rect 695 29756 697 29808
rect 1293 29756 1295 29808
rect 695 29744 727 29756
rect 1263 29744 1295 29756
rect 695 29692 697 29744
rect 1293 29692 1295 29744
rect 695 29680 727 29692
rect 1263 29680 1295 29692
rect 695 29628 697 29680
rect 1293 29628 1295 29680
rect 695 29616 727 29628
rect 1263 29616 1295 29628
rect 695 29564 697 29616
rect 1293 29564 1295 29616
rect 695 29552 727 29564
rect 1263 29552 1295 29564
rect 695 29500 697 29552
rect 1293 29500 1295 29552
rect 695 29488 727 29500
rect 1263 29488 1295 29500
rect 695 29436 697 29488
rect 1293 29436 1295 29488
rect 695 29424 727 29436
rect 1263 29424 1295 29436
rect 695 29372 697 29424
rect 749 29388 765 29413
rect 817 29388 833 29413
rect 885 29388 901 29413
rect 953 29388 969 29413
rect 1021 29388 1037 29413
rect 1089 29388 1105 29413
rect 1157 29388 1173 29413
rect 1225 29388 1241 29413
rect 885 29372 887 29388
rect 953 29372 967 29388
rect 1023 29372 1037 29388
rect 1103 29372 1105 29388
rect 1293 29372 1295 29424
rect 695 29360 727 29372
rect 783 29360 807 29372
rect 863 29360 887 29372
rect 943 29360 967 29372
rect 1023 29360 1047 29372
rect 1103 29360 1127 29372
rect 1183 29360 1207 29372
rect 1263 29360 1295 29372
rect 695 29308 697 29360
rect 885 29332 887 29360
rect 953 29332 967 29360
rect 1023 29332 1037 29360
rect 1103 29332 1105 29360
rect 749 29308 765 29332
rect 817 29308 833 29332
rect 885 29308 901 29332
rect 953 29308 969 29332
rect 1021 29308 1037 29332
rect 1089 29308 1105 29332
rect 1157 29308 1173 29332
rect 1225 29308 1241 29332
rect 1293 29308 1295 29360
rect 695 29307 1295 29308
rect 695 29296 727 29307
rect 783 29296 807 29307
rect 863 29296 887 29307
rect 943 29296 967 29307
rect 1023 29296 1047 29307
rect 1103 29296 1127 29307
rect 1183 29296 1207 29307
rect 1263 29296 1295 29307
rect 695 29244 697 29296
rect 885 29251 887 29296
rect 953 29251 967 29296
rect 1023 29251 1037 29296
rect 1103 29251 1105 29296
rect 749 29244 765 29251
rect 817 29244 833 29251
rect 885 29244 901 29251
rect 953 29244 969 29251
rect 1021 29244 1037 29251
rect 1089 29244 1105 29251
rect 1157 29244 1173 29251
rect 1225 29244 1241 29251
rect 1293 29244 1295 29296
rect 695 29232 1295 29244
rect 695 29180 697 29232
rect 749 29226 765 29232
rect 817 29226 833 29232
rect 885 29226 901 29232
rect 953 29226 969 29232
rect 1021 29226 1037 29232
rect 1089 29226 1105 29232
rect 1157 29226 1173 29232
rect 1225 29226 1241 29232
rect 885 29180 887 29226
rect 953 29180 967 29226
rect 1023 29180 1037 29226
rect 1103 29180 1105 29226
rect 1293 29180 1295 29232
rect 695 29170 727 29180
rect 783 29170 807 29180
rect 863 29170 887 29180
rect 943 29170 967 29180
rect 1023 29170 1047 29180
rect 1103 29170 1127 29180
rect 1183 29170 1207 29180
rect 1263 29170 1295 29180
rect 695 29168 1295 29170
rect 695 29116 697 29168
rect 749 29145 765 29168
rect 817 29145 833 29168
rect 885 29145 901 29168
rect 953 29145 969 29168
rect 1021 29145 1037 29168
rect 1089 29145 1105 29168
rect 1157 29145 1173 29168
rect 1225 29145 1241 29168
rect 885 29116 887 29145
rect 953 29116 967 29145
rect 1023 29116 1037 29145
rect 1103 29116 1105 29145
rect 1293 29116 1295 29168
rect 695 29104 727 29116
rect 783 29104 807 29116
rect 863 29104 887 29116
rect 943 29104 967 29116
rect 1023 29104 1047 29116
rect 1103 29104 1127 29116
rect 1183 29104 1207 29116
rect 1263 29104 1295 29116
rect 695 29052 697 29104
rect 885 29089 887 29104
rect 953 29089 967 29104
rect 1023 29089 1037 29104
rect 1103 29089 1105 29104
rect 749 29064 765 29089
rect 817 29064 833 29089
rect 885 29064 901 29089
rect 953 29064 969 29089
rect 1021 29064 1037 29089
rect 1089 29064 1105 29089
rect 1157 29064 1173 29089
rect 1225 29064 1241 29089
rect 885 29052 887 29064
rect 953 29052 967 29064
rect 1023 29052 1037 29064
rect 1103 29052 1105 29064
rect 1293 29052 1295 29104
rect 695 29040 727 29052
rect 783 29040 807 29052
rect 863 29040 887 29052
rect 943 29040 967 29052
rect 1023 29040 1047 29052
rect 1103 29040 1127 29052
rect 1183 29040 1207 29052
rect 1263 29040 1295 29052
rect 695 28988 697 29040
rect 885 29008 887 29040
rect 953 29008 967 29040
rect 1023 29008 1037 29040
rect 1103 29008 1105 29040
rect 749 28988 765 29008
rect 817 28988 833 29008
rect 885 28988 901 29008
rect 953 28988 969 29008
rect 1021 28988 1037 29008
rect 1089 28988 1105 29008
rect 1157 28988 1173 29008
rect 1225 28988 1241 29008
rect 1293 28988 1295 29040
rect 695 28983 1295 28988
rect 695 28976 727 28983
rect 783 28976 807 28983
rect 863 28976 887 28983
rect 943 28976 967 28983
rect 1023 28976 1047 28983
rect 1103 28976 1127 28983
rect 1183 28976 1207 28983
rect 1263 28976 1295 28983
rect 695 28924 697 28976
rect 885 28927 887 28976
rect 953 28927 967 28976
rect 1023 28927 1037 28976
rect 1103 28927 1105 28976
rect 749 28924 765 28927
rect 817 28924 833 28927
rect 885 28924 901 28927
rect 953 28924 969 28927
rect 1021 28924 1037 28927
rect 1089 28924 1105 28927
rect 1157 28924 1173 28927
rect 1225 28924 1241 28927
rect 1293 28924 1295 28976
rect 695 27865 1295 28924
rect 695 27813 697 27865
rect 749 27862 765 27865
rect 817 27862 833 27865
rect 885 27862 901 27865
rect 953 27862 969 27865
rect 1021 27862 1037 27865
rect 1089 27862 1105 27865
rect 1157 27862 1173 27865
rect 1225 27862 1241 27865
rect 1293 27813 1295 27865
rect 695 27801 727 27813
rect 1263 27801 1295 27813
rect 695 27749 697 27801
rect 1293 27749 1295 27801
rect 695 27737 727 27749
rect 1263 27737 1295 27749
rect 695 27685 697 27737
rect 1293 27685 1295 27737
rect 695 27673 727 27685
rect 1263 27673 1295 27685
rect 695 27621 697 27673
rect 1293 27621 1295 27673
rect 695 27609 727 27621
rect 1263 27609 1295 27621
rect 695 27557 697 27609
rect 1293 27557 1295 27609
rect 695 27545 727 27557
rect 1263 27545 1295 27557
rect 695 27493 697 27545
rect 1293 27493 1295 27545
rect 695 27481 727 27493
rect 1263 27481 1295 27493
rect 695 27429 697 27481
rect 1293 27429 1295 27481
rect 695 27417 727 27429
rect 1263 27417 1295 27429
rect 695 27365 697 27417
rect 749 27381 765 27406
rect 817 27381 833 27406
rect 885 27381 901 27406
rect 953 27381 969 27406
rect 1021 27381 1037 27406
rect 1089 27381 1105 27406
rect 1157 27381 1173 27406
rect 1225 27381 1241 27406
rect 885 27365 887 27381
rect 953 27365 967 27381
rect 1023 27365 1037 27381
rect 1103 27365 1105 27381
rect 1293 27365 1295 27417
rect 695 27353 727 27365
rect 783 27353 807 27365
rect 863 27353 887 27365
rect 943 27353 967 27365
rect 1023 27353 1047 27365
rect 1103 27353 1127 27365
rect 1183 27353 1207 27365
rect 1263 27353 1295 27365
rect 695 27301 697 27353
rect 885 27325 887 27353
rect 953 27325 967 27353
rect 1023 27325 1037 27353
rect 1103 27325 1105 27353
rect 749 27301 765 27325
rect 817 27301 833 27325
rect 885 27301 901 27325
rect 953 27301 969 27325
rect 1021 27301 1037 27325
rect 1089 27301 1105 27325
rect 1157 27301 1173 27325
rect 1225 27301 1241 27325
rect 1293 27301 1295 27353
rect 695 27300 1295 27301
rect 695 27289 727 27300
rect 783 27289 807 27300
rect 863 27289 887 27300
rect 943 27289 967 27300
rect 1023 27289 1047 27300
rect 1103 27289 1127 27300
rect 1183 27289 1207 27300
rect 1263 27289 1295 27300
rect 695 27237 697 27289
rect 885 27244 887 27289
rect 953 27244 967 27289
rect 1023 27244 1037 27289
rect 1103 27244 1105 27289
rect 749 27237 765 27244
rect 817 27237 833 27244
rect 885 27237 901 27244
rect 953 27237 969 27244
rect 1021 27237 1037 27244
rect 1089 27237 1105 27244
rect 1157 27237 1173 27244
rect 1225 27237 1241 27244
rect 1293 27237 1295 27289
rect 695 27225 1295 27237
rect 695 27173 697 27225
rect 749 27219 765 27225
rect 817 27219 833 27225
rect 885 27219 901 27225
rect 953 27219 969 27225
rect 1021 27219 1037 27225
rect 1089 27219 1105 27225
rect 1157 27219 1173 27225
rect 1225 27219 1241 27225
rect 885 27173 887 27219
rect 953 27173 967 27219
rect 1023 27173 1037 27219
rect 1103 27173 1105 27219
rect 1293 27173 1295 27225
rect 695 27163 727 27173
rect 783 27163 807 27173
rect 863 27163 887 27173
rect 943 27163 967 27173
rect 1023 27163 1047 27173
rect 1103 27163 1127 27173
rect 1183 27163 1207 27173
rect 1263 27163 1295 27173
rect 695 27161 1295 27163
rect 695 27109 697 27161
rect 749 27138 765 27161
rect 817 27138 833 27161
rect 885 27138 901 27161
rect 953 27138 969 27161
rect 1021 27138 1037 27161
rect 1089 27138 1105 27161
rect 1157 27138 1173 27161
rect 1225 27138 1241 27161
rect 885 27109 887 27138
rect 953 27109 967 27138
rect 1023 27109 1037 27138
rect 1103 27109 1105 27138
rect 1293 27109 1295 27161
rect 695 27097 727 27109
rect 783 27097 807 27109
rect 863 27097 887 27109
rect 943 27097 967 27109
rect 1023 27097 1047 27109
rect 1103 27097 1127 27109
rect 1183 27097 1207 27109
rect 1263 27097 1295 27109
rect 695 27045 697 27097
rect 885 27082 887 27097
rect 953 27082 967 27097
rect 1023 27082 1037 27097
rect 1103 27082 1105 27097
rect 749 27057 765 27082
rect 817 27057 833 27082
rect 885 27057 901 27082
rect 953 27057 969 27082
rect 1021 27057 1037 27082
rect 1089 27057 1105 27082
rect 1157 27057 1173 27082
rect 1225 27057 1241 27082
rect 885 27045 887 27057
rect 953 27045 967 27057
rect 1023 27045 1037 27057
rect 1103 27045 1105 27057
rect 1293 27045 1295 27097
rect 695 27033 727 27045
rect 783 27033 807 27045
rect 863 27033 887 27045
rect 943 27033 967 27045
rect 1023 27033 1047 27045
rect 1103 27033 1127 27045
rect 1183 27033 1207 27045
rect 1263 27033 1295 27045
rect 695 26981 697 27033
rect 885 27001 887 27033
rect 953 27001 967 27033
rect 1023 27001 1037 27033
rect 1103 27001 1105 27033
rect 749 26981 765 27001
rect 817 26981 833 27001
rect 885 26981 901 27001
rect 953 26981 969 27001
rect 1021 26981 1037 27001
rect 1089 26981 1105 27001
rect 1157 26981 1173 27001
rect 1225 26981 1241 27001
rect 1293 26981 1295 27033
rect 695 26976 1295 26981
rect 695 26969 727 26976
rect 783 26969 807 26976
rect 863 26969 887 26976
rect 943 26969 967 26976
rect 1023 26969 1047 26976
rect 1103 26969 1127 26976
rect 1183 26969 1207 26976
rect 1263 26969 1295 26976
rect 695 26917 697 26969
rect 885 26920 887 26969
rect 953 26920 967 26969
rect 1023 26920 1037 26969
rect 1103 26920 1105 26969
rect 749 26917 765 26920
rect 817 26917 833 26920
rect 885 26917 901 26920
rect 953 26917 969 26920
rect 1021 26917 1037 26920
rect 1089 26917 1105 26920
rect 1157 26917 1173 26920
rect 1225 26917 1241 26920
rect 1293 26917 1295 26969
rect 695 25679 1295 26917
rect 695 25627 697 25679
rect 749 25676 765 25679
rect 817 25676 833 25679
rect 885 25676 901 25679
rect 953 25676 969 25679
rect 1021 25676 1037 25679
rect 1089 25676 1105 25679
rect 1157 25676 1173 25679
rect 1225 25676 1241 25679
rect 1293 25627 1295 25679
rect 695 25615 727 25627
rect 1263 25615 1295 25627
rect 695 25563 697 25615
rect 1293 25563 1295 25615
rect 695 25551 727 25563
rect 1263 25551 1295 25563
rect 695 25499 697 25551
rect 1293 25499 1295 25551
rect 695 25487 727 25499
rect 1263 25487 1295 25499
rect 695 25435 697 25487
rect 1293 25435 1295 25487
rect 695 25423 727 25435
rect 1263 25423 1295 25435
rect 695 25371 697 25423
rect 1293 25371 1295 25423
rect 695 25359 727 25371
rect 1263 25359 1295 25371
rect 695 25307 697 25359
rect 1293 25307 1295 25359
rect 695 25295 727 25307
rect 1263 25295 1295 25307
rect 695 25243 697 25295
rect 1293 25243 1295 25295
rect 695 25231 727 25243
rect 1263 25231 1295 25243
rect 695 25179 697 25231
rect 749 25195 765 25220
rect 817 25195 833 25220
rect 885 25195 901 25220
rect 953 25195 969 25220
rect 1021 25195 1037 25220
rect 1089 25195 1105 25220
rect 1157 25195 1173 25220
rect 1225 25195 1241 25220
rect 885 25179 887 25195
rect 953 25179 967 25195
rect 1023 25179 1037 25195
rect 1103 25179 1105 25195
rect 1293 25179 1295 25231
rect 695 25167 727 25179
rect 783 25167 807 25179
rect 863 25167 887 25179
rect 943 25167 967 25179
rect 1023 25167 1047 25179
rect 1103 25167 1127 25179
rect 1183 25167 1207 25179
rect 1263 25167 1295 25179
rect 695 25115 697 25167
rect 885 25139 887 25167
rect 953 25139 967 25167
rect 1023 25139 1037 25167
rect 1103 25139 1105 25167
rect 749 25115 765 25139
rect 817 25115 833 25139
rect 885 25115 901 25139
rect 953 25115 969 25139
rect 1021 25115 1037 25139
rect 1089 25115 1105 25139
rect 1157 25115 1173 25139
rect 1225 25115 1241 25139
rect 1293 25115 1295 25167
rect 695 25114 1295 25115
rect 695 25103 727 25114
rect 783 25103 807 25114
rect 863 25103 887 25114
rect 943 25103 967 25114
rect 1023 25103 1047 25114
rect 1103 25103 1127 25114
rect 1183 25103 1207 25114
rect 1263 25103 1295 25114
rect 695 25051 697 25103
rect 885 25058 887 25103
rect 953 25058 967 25103
rect 1023 25058 1037 25103
rect 1103 25058 1105 25103
rect 749 25051 765 25058
rect 817 25051 833 25058
rect 885 25051 901 25058
rect 953 25051 969 25058
rect 1021 25051 1037 25058
rect 1089 25051 1105 25058
rect 1157 25051 1173 25058
rect 1225 25051 1241 25058
rect 1293 25051 1295 25103
rect 695 25039 1295 25051
rect 695 24987 697 25039
rect 749 25033 765 25039
rect 817 25033 833 25039
rect 885 25033 901 25039
rect 953 25033 969 25039
rect 1021 25033 1037 25039
rect 1089 25033 1105 25039
rect 1157 25033 1173 25039
rect 1225 25033 1241 25039
rect 885 24987 887 25033
rect 953 24987 967 25033
rect 1023 24987 1037 25033
rect 1103 24987 1105 25033
rect 1293 24987 1295 25039
rect 695 24977 727 24987
rect 783 24977 807 24987
rect 863 24977 887 24987
rect 943 24977 967 24987
rect 1023 24977 1047 24987
rect 1103 24977 1127 24987
rect 1183 24977 1207 24987
rect 1263 24977 1295 24987
rect 695 24975 1295 24977
rect 695 24923 697 24975
rect 749 24952 765 24975
rect 817 24952 833 24975
rect 885 24952 901 24975
rect 953 24952 969 24975
rect 1021 24952 1037 24975
rect 1089 24952 1105 24975
rect 1157 24952 1173 24975
rect 1225 24952 1241 24975
rect 885 24923 887 24952
rect 953 24923 967 24952
rect 1023 24923 1037 24952
rect 1103 24923 1105 24952
rect 1293 24923 1295 24975
rect 695 24911 727 24923
rect 783 24911 807 24923
rect 863 24911 887 24923
rect 943 24911 967 24923
rect 1023 24911 1047 24923
rect 1103 24911 1127 24923
rect 1183 24911 1207 24923
rect 1263 24911 1295 24923
rect 695 24859 697 24911
rect 885 24896 887 24911
rect 953 24896 967 24911
rect 1023 24896 1037 24911
rect 1103 24896 1105 24911
rect 749 24871 765 24896
rect 817 24871 833 24896
rect 885 24871 901 24896
rect 953 24871 969 24896
rect 1021 24871 1037 24896
rect 1089 24871 1105 24896
rect 1157 24871 1173 24896
rect 1225 24871 1241 24896
rect 885 24859 887 24871
rect 953 24859 967 24871
rect 1023 24859 1037 24871
rect 1103 24859 1105 24871
rect 1293 24859 1295 24911
rect 695 24847 727 24859
rect 783 24847 807 24859
rect 863 24847 887 24859
rect 943 24847 967 24859
rect 1023 24847 1047 24859
rect 1103 24847 1127 24859
rect 1183 24847 1207 24859
rect 1263 24847 1295 24859
rect 695 24795 697 24847
rect 885 24815 887 24847
rect 953 24815 967 24847
rect 1023 24815 1037 24847
rect 1103 24815 1105 24847
rect 749 24795 765 24815
rect 817 24795 833 24815
rect 885 24795 901 24815
rect 953 24795 969 24815
rect 1021 24795 1037 24815
rect 1089 24795 1105 24815
rect 1157 24795 1173 24815
rect 1225 24795 1241 24815
rect 1293 24795 1295 24847
rect 695 24790 1295 24795
rect 695 24783 727 24790
rect 783 24783 807 24790
rect 863 24783 887 24790
rect 943 24783 967 24790
rect 1023 24783 1047 24790
rect 1103 24783 1127 24790
rect 1183 24783 1207 24790
rect 1263 24783 1295 24790
rect 695 24731 697 24783
rect 885 24734 887 24783
rect 953 24734 967 24783
rect 1023 24734 1037 24783
rect 1103 24734 1105 24783
rect 749 24731 765 24734
rect 817 24731 833 24734
rect 885 24731 901 24734
rect 953 24731 969 24734
rect 1021 24731 1037 24734
rect 1089 24731 1105 24734
rect 1157 24731 1173 24734
rect 1225 24731 1241 24734
rect 1293 24731 1295 24783
rect 695 23531 1295 24731
rect 695 23479 697 23531
rect 749 23528 765 23531
rect 817 23528 833 23531
rect 885 23528 901 23531
rect 953 23528 969 23531
rect 1021 23528 1037 23531
rect 1089 23528 1105 23531
rect 1157 23528 1173 23531
rect 1225 23528 1241 23531
rect 1293 23479 1295 23531
rect 695 23467 727 23479
rect 1263 23467 1295 23479
rect 695 23415 697 23467
rect 1293 23415 1295 23467
rect 695 23403 727 23415
rect 1263 23403 1295 23415
rect 695 23351 697 23403
rect 1293 23351 1295 23403
rect 695 23339 727 23351
rect 1263 23339 1295 23351
rect 695 23287 697 23339
rect 1293 23287 1295 23339
rect 695 23275 727 23287
rect 1263 23275 1295 23287
rect 695 23223 697 23275
rect 1293 23223 1295 23275
rect 695 23211 727 23223
rect 1263 23211 1295 23223
rect 695 23159 697 23211
rect 1293 23159 1295 23211
rect 695 23147 727 23159
rect 1263 23147 1295 23159
rect 695 23095 697 23147
rect 1293 23095 1295 23147
rect 695 23083 727 23095
rect 1263 23083 1295 23095
rect 695 23031 697 23083
rect 749 23047 765 23072
rect 817 23047 833 23072
rect 885 23047 901 23072
rect 953 23047 969 23072
rect 1021 23047 1037 23072
rect 1089 23047 1105 23072
rect 1157 23047 1173 23072
rect 1225 23047 1241 23072
rect 885 23031 887 23047
rect 953 23031 967 23047
rect 1023 23031 1037 23047
rect 1103 23031 1105 23047
rect 1293 23031 1295 23083
rect 695 23019 727 23031
rect 783 23019 807 23031
rect 863 23019 887 23031
rect 943 23019 967 23031
rect 1023 23019 1047 23031
rect 1103 23019 1127 23031
rect 1183 23019 1207 23031
rect 1263 23019 1295 23031
rect 695 22967 697 23019
rect 885 22991 887 23019
rect 953 22991 967 23019
rect 1023 22991 1037 23019
rect 1103 22991 1105 23019
rect 749 22967 765 22991
rect 817 22967 833 22991
rect 885 22967 901 22991
rect 953 22967 969 22991
rect 1021 22967 1037 22991
rect 1089 22967 1105 22991
rect 1157 22967 1173 22991
rect 1225 22967 1241 22991
rect 1293 22967 1295 23019
rect 695 22966 1295 22967
rect 695 22955 727 22966
rect 783 22955 807 22966
rect 863 22955 887 22966
rect 943 22955 967 22966
rect 1023 22955 1047 22966
rect 1103 22955 1127 22966
rect 1183 22955 1207 22966
rect 1263 22955 1295 22966
rect 695 22903 697 22955
rect 885 22910 887 22955
rect 953 22910 967 22955
rect 1023 22910 1037 22955
rect 1103 22910 1105 22955
rect 749 22903 765 22910
rect 817 22903 833 22910
rect 885 22903 901 22910
rect 953 22903 969 22910
rect 1021 22903 1037 22910
rect 1089 22903 1105 22910
rect 1157 22903 1173 22910
rect 1225 22903 1241 22910
rect 1293 22903 1295 22955
rect 695 22891 1295 22903
rect 695 22839 697 22891
rect 749 22885 765 22891
rect 817 22885 833 22891
rect 885 22885 901 22891
rect 953 22885 969 22891
rect 1021 22885 1037 22891
rect 1089 22885 1105 22891
rect 1157 22885 1173 22891
rect 1225 22885 1241 22891
rect 885 22839 887 22885
rect 953 22839 967 22885
rect 1023 22839 1037 22885
rect 1103 22839 1105 22885
rect 1293 22839 1295 22891
rect 695 22829 727 22839
rect 783 22829 807 22839
rect 863 22829 887 22839
rect 943 22829 967 22839
rect 1023 22829 1047 22839
rect 1103 22829 1127 22839
rect 1183 22829 1207 22839
rect 1263 22829 1295 22839
rect 695 22827 1295 22829
rect 695 22775 697 22827
rect 749 22804 765 22827
rect 817 22804 833 22827
rect 885 22804 901 22827
rect 953 22804 969 22827
rect 1021 22804 1037 22827
rect 1089 22804 1105 22827
rect 1157 22804 1173 22827
rect 1225 22804 1241 22827
rect 885 22775 887 22804
rect 953 22775 967 22804
rect 1023 22775 1037 22804
rect 1103 22775 1105 22804
rect 1293 22775 1295 22827
rect 695 22763 727 22775
rect 783 22763 807 22775
rect 863 22763 887 22775
rect 943 22763 967 22775
rect 1023 22763 1047 22775
rect 1103 22763 1127 22775
rect 1183 22763 1207 22775
rect 1263 22763 1295 22775
rect 695 22711 697 22763
rect 885 22748 887 22763
rect 953 22748 967 22763
rect 1023 22748 1037 22763
rect 1103 22748 1105 22763
rect 749 22723 765 22748
rect 817 22723 833 22748
rect 885 22723 901 22748
rect 953 22723 969 22748
rect 1021 22723 1037 22748
rect 1089 22723 1105 22748
rect 1157 22723 1173 22748
rect 1225 22723 1241 22748
rect 885 22711 887 22723
rect 953 22711 967 22723
rect 1023 22711 1037 22723
rect 1103 22711 1105 22723
rect 1293 22711 1295 22763
rect 695 22699 727 22711
rect 783 22699 807 22711
rect 863 22699 887 22711
rect 943 22699 967 22711
rect 1023 22699 1047 22711
rect 1103 22699 1127 22711
rect 1183 22699 1207 22711
rect 1263 22699 1295 22711
rect 695 22647 697 22699
rect 885 22667 887 22699
rect 953 22667 967 22699
rect 1023 22667 1037 22699
rect 1103 22667 1105 22699
rect 749 22647 765 22667
rect 817 22647 833 22667
rect 885 22647 901 22667
rect 953 22647 969 22667
rect 1021 22647 1037 22667
rect 1089 22647 1105 22667
rect 1157 22647 1173 22667
rect 1225 22647 1241 22667
rect 1293 22647 1295 22699
rect 695 22642 1295 22647
rect 695 22635 727 22642
rect 783 22635 807 22642
rect 863 22635 887 22642
rect 943 22635 967 22642
rect 1023 22635 1047 22642
rect 1103 22635 1127 22642
rect 1183 22635 1207 22642
rect 1263 22635 1295 22642
rect 695 22583 697 22635
rect 885 22586 887 22635
rect 953 22586 967 22635
rect 1023 22586 1037 22635
rect 1103 22586 1105 22635
rect 749 22583 765 22586
rect 817 22583 833 22586
rect 885 22583 901 22586
rect 953 22583 969 22586
rect 1021 22583 1037 22586
rect 1089 22583 1105 22586
rect 1157 22583 1173 22586
rect 1225 22583 1241 22586
rect 1293 22583 1295 22635
rect 695 21361 1295 22583
rect 695 21309 697 21361
rect 749 21358 765 21361
rect 817 21358 833 21361
rect 885 21358 901 21361
rect 953 21358 969 21361
rect 1021 21358 1037 21361
rect 1089 21358 1105 21361
rect 1157 21358 1173 21361
rect 1225 21358 1241 21361
rect 1293 21309 1295 21361
rect 695 21297 727 21309
rect 1263 21297 1295 21309
rect 695 21245 697 21297
rect 1293 21245 1295 21297
rect 695 21233 727 21245
rect 1263 21233 1295 21245
rect 695 21181 697 21233
rect 1293 21181 1295 21233
rect 695 21169 727 21181
rect 1263 21169 1295 21181
rect 695 21117 697 21169
rect 1293 21117 1295 21169
rect 695 21105 727 21117
rect 1263 21105 1295 21117
rect 695 21053 697 21105
rect 1293 21053 1295 21105
rect 695 21041 727 21053
rect 1263 21041 1295 21053
rect 695 20989 697 21041
rect 1293 20989 1295 21041
rect 695 20977 727 20989
rect 1263 20977 1295 20989
rect 695 20925 697 20977
rect 1293 20925 1295 20977
rect 695 20913 727 20925
rect 1263 20913 1295 20925
rect 695 20861 697 20913
rect 749 20877 765 20902
rect 817 20877 833 20902
rect 885 20877 901 20902
rect 953 20877 969 20902
rect 1021 20877 1037 20902
rect 1089 20877 1105 20902
rect 1157 20877 1173 20902
rect 1225 20877 1241 20902
rect 885 20861 887 20877
rect 953 20861 967 20877
rect 1023 20861 1037 20877
rect 1103 20861 1105 20877
rect 1293 20861 1295 20913
rect 695 20849 727 20861
rect 783 20849 807 20861
rect 863 20849 887 20861
rect 943 20849 967 20861
rect 1023 20849 1047 20861
rect 1103 20849 1127 20861
rect 1183 20849 1207 20861
rect 1263 20849 1295 20861
rect 695 20797 697 20849
rect 885 20821 887 20849
rect 953 20821 967 20849
rect 1023 20821 1037 20849
rect 1103 20821 1105 20849
rect 749 20797 765 20821
rect 817 20797 833 20821
rect 885 20797 901 20821
rect 953 20797 969 20821
rect 1021 20797 1037 20821
rect 1089 20797 1105 20821
rect 1157 20797 1173 20821
rect 1225 20797 1241 20821
rect 1293 20797 1295 20849
rect 695 20796 1295 20797
rect 695 20785 727 20796
rect 783 20785 807 20796
rect 863 20785 887 20796
rect 943 20785 967 20796
rect 1023 20785 1047 20796
rect 1103 20785 1127 20796
rect 1183 20785 1207 20796
rect 1263 20785 1295 20796
rect 695 20733 697 20785
rect 885 20740 887 20785
rect 953 20740 967 20785
rect 1023 20740 1037 20785
rect 1103 20740 1105 20785
rect 749 20733 765 20740
rect 817 20733 833 20740
rect 885 20733 901 20740
rect 953 20733 969 20740
rect 1021 20733 1037 20740
rect 1089 20733 1105 20740
rect 1157 20733 1173 20740
rect 1225 20733 1241 20740
rect 1293 20733 1295 20785
rect 695 20721 1295 20733
rect 695 20669 697 20721
rect 749 20715 765 20721
rect 817 20715 833 20721
rect 885 20715 901 20721
rect 953 20715 969 20721
rect 1021 20715 1037 20721
rect 1089 20715 1105 20721
rect 1157 20715 1173 20721
rect 1225 20715 1241 20721
rect 885 20669 887 20715
rect 953 20669 967 20715
rect 1023 20669 1037 20715
rect 1103 20669 1105 20715
rect 1293 20669 1295 20721
rect 695 20659 727 20669
rect 783 20659 807 20669
rect 863 20659 887 20669
rect 943 20659 967 20669
rect 1023 20659 1047 20669
rect 1103 20659 1127 20669
rect 1183 20659 1207 20669
rect 1263 20659 1295 20669
rect 695 20657 1295 20659
rect 695 20605 697 20657
rect 749 20634 765 20657
rect 817 20634 833 20657
rect 885 20634 901 20657
rect 953 20634 969 20657
rect 1021 20634 1037 20657
rect 1089 20634 1105 20657
rect 1157 20634 1173 20657
rect 1225 20634 1241 20657
rect 885 20605 887 20634
rect 953 20605 967 20634
rect 1023 20605 1037 20634
rect 1103 20605 1105 20634
rect 1293 20605 1295 20657
rect 695 20593 727 20605
rect 783 20593 807 20605
rect 863 20593 887 20605
rect 943 20593 967 20605
rect 1023 20593 1047 20605
rect 1103 20593 1127 20605
rect 1183 20593 1207 20605
rect 1263 20593 1295 20605
rect 695 20541 697 20593
rect 885 20578 887 20593
rect 953 20578 967 20593
rect 1023 20578 1037 20593
rect 1103 20578 1105 20593
rect 749 20553 765 20578
rect 817 20553 833 20578
rect 885 20553 901 20578
rect 953 20553 969 20578
rect 1021 20553 1037 20578
rect 1089 20553 1105 20578
rect 1157 20553 1173 20578
rect 1225 20553 1241 20578
rect 885 20541 887 20553
rect 953 20541 967 20553
rect 1023 20541 1037 20553
rect 1103 20541 1105 20553
rect 1293 20541 1295 20593
rect 695 20529 727 20541
rect 783 20529 807 20541
rect 863 20529 887 20541
rect 943 20529 967 20541
rect 1023 20529 1047 20541
rect 1103 20529 1127 20541
rect 1183 20529 1207 20541
rect 1263 20529 1295 20541
rect 695 20477 697 20529
rect 885 20497 887 20529
rect 953 20497 967 20529
rect 1023 20497 1037 20529
rect 1103 20497 1105 20529
rect 749 20477 765 20497
rect 817 20477 833 20497
rect 885 20477 901 20497
rect 953 20477 969 20497
rect 1021 20477 1037 20497
rect 1089 20477 1105 20497
rect 1157 20477 1173 20497
rect 1225 20477 1241 20497
rect 1293 20477 1295 20529
rect 695 20472 1295 20477
rect 695 20465 727 20472
rect 783 20465 807 20472
rect 863 20465 887 20472
rect 943 20465 967 20472
rect 1023 20465 1047 20472
rect 1103 20465 1127 20472
rect 1183 20465 1207 20472
rect 1263 20465 1295 20472
rect 695 20413 697 20465
rect 885 20416 887 20465
rect 953 20416 967 20465
rect 1023 20416 1037 20465
rect 1103 20416 1105 20465
rect 749 20413 765 20416
rect 817 20413 833 20416
rect 885 20413 901 20416
rect 953 20413 969 20416
rect 1021 20413 1037 20416
rect 1089 20413 1105 20416
rect 1157 20413 1173 20416
rect 1225 20413 1241 20416
rect 1293 20413 1295 20465
rect 695 19257 1295 20413
rect 695 19205 697 19257
rect 749 19254 765 19257
rect 817 19254 833 19257
rect 885 19254 901 19257
rect 953 19254 969 19257
rect 1021 19254 1037 19257
rect 1089 19254 1105 19257
rect 1157 19254 1173 19257
rect 1225 19254 1241 19257
rect 1293 19205 1295 19257
rect 695 19193 727 19205
rect 1263 19193 1295 19205
rect 695 19141 697 19193
rect 1293 19141 1295 19193
rect 695 19129 727 19141
rect 1263 19129 1295 19141
rect 695 19077 697 19129
rect 1293 19077 1295 19129
rect 695 19065 727 19077
rect 1263 19065 1295 19077
rect 695 19013 697 19065
rect 1293 19013 1295 19065
rect 695 19001 727 19013
rect 1263 19001 1295 19013
rect 695 18949 697 19001
rect 1293 18949 1295 19001
rect 695 18937 727 18949
rect 1263 18937 1295 18949
rect 695 18885 697 18937
rect 1293 18885 1295 18937
rect 695 18873 727 18885
rect 1263 18873 1295 18885
rect 695 18821 697 18873
rect 1293 18821 1295 18873
rect 695 18809 727 18821
rect 1263 18809 1295 18821
rect 695 18757 697 18809
rect 749 18773 765 18798
rect 817 18773 833 18798
rect 885 18773 901 18798
rect 953 18773 969 18798
rect 1021 18773 1037 18798
rect 1089 18773 1105 18798
rect 1157 18773 1173 18798
rect 1225 18773 1241 18798
rect 885 18757 887 18773
rect 953 18757 967 18773
rect 1023 18757 1037 18773
rect 1103 18757 1105 18773
rect 1293 18757 1295 18809
rect 695 18745 727 18757
rect 783 18745 807 18757
rect 863 18745 887 18757
rect 943 18745 967 18757
rect 1023 18745 1047 18757
rect 1103 18745 1127 18757
rect 1183 18745 1207 18757
rect 1263 18745 1295 18757
rect 695 18693 697 18745
rect 885 18717 887 18745
rect 953 18717 967 18745
rect 1023 18717 1037 18745
rect 1103 18717 1105 18745
rect 749 18693 765 18717
rect 817 18693 833 18717
rect 885 18693 901 18717
rect 953 18693 969 18717
rect 1021 18693 1037 18717
rect 1089 18693 1105 18717
rect 1157 18693 1173 18717
rect 1225 18693 1241 18717
rect 1293 18693 1295 18745
rect 695 18692 1295 18693
rect 695 18681 727 18692
rect 783 18681 807 18692
rect 863 18681 887 18692
rect 943 18681 967 18692
rect 1023 18681 1047 18692
rect 1103 18681 1127 18692
rect 1183 18681 1207 18692
rect 1263 18681 1295 18692
rect 695 18629 697 18681
rect 885 18636 887 18681
rect 953 18636 967 18681
rect 1023 18636 1037 18681
rect 1103 18636 1105 18681
rect 749 18629 765 18636
rect 817 18629 833 18636
rect 885 18629 901 18636
rect 953 18629 969 18636
rect 1021 18629 1037 18636
rect 1089 18629 1105 18636
rect 1157 18629 1173 18636
rect 1225 18629 1241 18636
rect 1293 18629 1295 18681
rect 695 18617 1295 18629
rect 695 18565 697 18617
rect 749 18611 765 18617
rect 817 18611 833 18617
rect 885 18611 901 18617
rect 953 18611 969 18617
rect 1021 18611 1037 18617
rect 1089 18611 1105 18617
rect 1157 18611 1173 18617
rect 1225 18611 1241 18617
rect 885 18565 887 18611
rect 953 18565 967 18611
rect 1023 18565 1037 18611
rect 1103 18565 1105 18611
rect 1293 18565 1295 18617
rect 695 18555 727 18565
rect 783 18555 807 18565
rect 863 18555 887 18565
rect 943 18555 967 18565
rect 1023 18555 1047 18565
rect 1103 18555 1127 18565
rect 1183 18555 1207 18565
rect 1263 18555 1295 18565
rect 695 18553 1295 18555
rect 695 18501 697 18553
rect 749 18530 765 18553
rect 817 18530 833 18553
rect 885 18530 901 18553
rect 953 18530 969 18553
rect 1021 18530 1037 18553
rect 1089 18530 1105 18553
rect 1157 18530 1173 18553
rect 1225 18530 1241 18553
rect 885 18501 887 18530
rect 953 18501 967 18530
rect 1023 18501 1037 18530
rect 1103 18501 1105 18530
rect 1293 18501 1295 18553
rect 695 18489 727 18501
rect 783 18489 807 18501
rect 863 18489 887 18501
rect 943 18489 967 18501
rect 1023 18489 1047 18501
rect 1103 18489 1127 18501
rect 1183 18489 1207 18501
rect 1263 18489 1295 18501
rect 695 18437 697 18489
rect 885 18474 887 18489
rect 953 18474 967 18489
rect 1023 18474 1037 18489
rect 1103 18474 1105 18489
rect 749 18449 765 18474
rect 817 18449 833 18474
rect 885 18449 901 18474
rect 953 18449 969 18474
rect 1021 18449 1037 18474
rect 1089 18449 1105 18474
rect 1157 18449 1173 18474
rect 1225 18449 1241 18474
rect 885 18437 887 18449
rect 953 18437 967 18449
rect 1023 18437 1037 18449
rect 1103 18437 1105 18449
rect 1293 18437 1295 18489
rect 695 18425 727 18437
rect 783 18425 807 18437
rect 863 18425 887 18437
rect 943 18425 967 18437
rect 1023 18425 1047 18437
rect 1103 18425 1127 18437
rect 1183 18425 1207 18437
rect 1263 18425 1295 18437
rect 695 18373 697 18425
rect 885 18393 887 18425
rect 953 18393 967 18425
rect 1023 18393 1037 18425
rect 1103 18393 1105 18425
rect 749 18373 765 18393
rect 817 18373 833 18393
rect 885 18373 901 18393
rect 953 18373 969 18393
rect 1021 18373 1037 18393
rect 1089 18373 1105 18393
rect 1157 18373 1173 18393
rect 1225 18373 1241 18393
rect 1293 18373 1295 18425
rect 695 18368 1295 18373
rect 695 18361 727 18368
rect 783 18361 807 18368
rect 863 18361 887 18368
rect 943 18361 967 18368
rect 1023 18361 1047 18368
rect 1103 18361 1127 18368
rect 1183 18361 1207 18368
rect 1263 18361 1295 18368
rect 695 18309 697 18361
rect 885 18312 887 18361
rect 953 18312 967 18361
rect 1023 18312 1037 18361
rect 1103 18312 1105 18361
rect 749 18309 765 18312
rect 817 18309 833 18312
rect 885 18309 901 18312
rect 953 18309 969 18312
rect 1021 18309 1037 18312
rect 1089 18309 1105 18312
rect 1157 18309 1173 18312
rect 1225 18309 1241 18312
rect 1293 18309 1295 18361
rect 695 17146 1295 18309
rect 695 17094 697 17146
rect 749 17143 765 17146
rect 817 17143 833 17146
rect 885 17143 901 17146
rect 953 17143 969 17146
rect 1021 17143 1037 17146
rect 1089 17143 1105 17146
rect 1157 17143 1173 17146
rect 1225 17143 1241 17146
rect 1293 17094 1295 17146
rect 695 17082 727 17094
rect 1263 17082 1295 17094
rect 695 17030 697 17082
rect 1293 17030 1295 17082
rect 695 17018 727 17030
rect 1263 17018 1295 17030
rect 695 16966 697 17018
rect 1293 16966 1295 17018
rect 695 16954 727 16966
rect 1263 16954 1295 16966
rect 695 16902 697 16954
rect 1293 16902 1295 16954
rect 695 16890 727 16902
rect 1263 16890 1295 16902
rect 695 16838 697 16890
rect 1293 16838 1295 16890
rect 695 16826 727 16838
rect 1263 16826 1295 16838
rect 695 16774 697 16826
rect 1293 16774 1295 16826
rect 695 16762 727 16774
rect 1263 16762 1295 16774
rect 695 16710 697 16762
rect 1293 16710 1295 16762
rect 695 16698 727 16710
rect 1263 16698 1295 16710
rect 695 16646 697 16698
rect 749 16662 765 16687
rect 817 16662 833 16687
rect 885 16662 901 16687
rect 953 16662 969 16687
rect 1021 16662 1037 16687
rect 1089 16662 1105 16687
rect 1157 16662 1173 16687
rect 1225 16662 1241 16687
rect 885 16646 887 16662
rect 953 16646 967 16662
rect 1023 16646 1037 16662
rect 1103 16646 1105 16662
rect 1293 16646 1295 16698
rect 695 16634 727 16646
rect 783 16634 807 16646
rect 863 16634 887 16646
rect 943 16634 967 16646
rect 1023 16634 1047 16646
rect 1103 16634 1127 16646
rect 1183 16634 1207 16646
rect 1263 16634 1295 16646
rect 695 16582 697 16634
rect 885 16606 887 16634
rect 953 16606 967 16634
rect 1023 16606 1037 16634
rect 1103 16606 1105 16634
rect 749 16582 765 16606
rect 817 16582 833 16606
rect 885 16582 901 16606
rect 953 16582 969 16606
rect 1021 16582 1037 16606
rect 1089 16582 1105 16606
rect 1157 16582 1173 16606
rect 1225 16582 1241 16606
rect 1293 16582 1295 16634
rect 695 16581 1295 16582
rect 695 16570 727 16581
rect 783 16570 807 16581
rect 863 16570 887 16581
rect 943 16570 967 16581
rect 1023 16570 1047 16581
rect 1103 16570 1127 16581
rect 1183 16570 1207 16581
rect 1263 16570 1295 16581
rect 695 16518 697 16570
rect 885 16525 887 16570
rect 953 16525 967 16570
rect 1023 16525 1037 16570
rect 1103 16525 1105 16570
rect 749 16518 765 16525
rect 817 16518 833 16525
rect 885 16518 901 16525
rect 953 16518 969 16525
rect 1021 16518 1037 16525
rect 1089 16518 1105 16525
rect 1157 16518 1173 16525
rect 1225 16518 1241 16525
rect 1293 16518 1295 16570
rect 695 16506 1295 16518
rect 695 16454 697 16506
rect 749 16500 765 16506
rect 817 16500 833 16506
rect 885 16500 901 16506
rect 953 16500 969 16506
rect 1021 16500 1037 16506
rect 1089 16500 1105 16506
rect 1157 16500 1173 16506
rect 1225 16500 1241 16506
rect 885 16454 887 16500
rect 953 16454 967 16500
rect 1023 16454 1037 16500
rect 1103 16454 1105 16500
rect 1293 16454 1295 16506
rect 695 16444 727 16454
rect 783 16444 807 16454
rect 863 16444 887 16454
rect 943 16444 967 16454
rect 1023 16444 1047 16454
rect 1103 16444 1127 16454
rect 1183 16444 1207 16454
rect 1263 16444 1295 16454
rect 695 16442 1295 16444
rect 695 16390 697 16442
rect 749 16419 765 16442
rect 817 16419 833 16442
rect 885 16419 901 16442
rect 953 16419 969 16442
rect 1021 16419 1037 16442
rect 1089 16419 1105 16442
rect 1157 16419 1173 16442
rect 1225 16419 1241 16442
rect 885 16390 887 16419
rect 953 16390 967 16419
rect 1023 16390 1037 16419
rect 1103 16390 1105 16419
rect 1293 16390 1295 16442
rect 695 16378 727 16390
rect 783 16378 807 16390
rect 863 16378 887 16390
rect 943 16378 967 16390
rect 1023 16378 1047 16390
rect 1103 16378 1127 16390
rect 1183 16378 1207 16390
rect 1263 16378 1295 16390
rect 695 16326 697 16378
rect 885 16363 887 16378
rect 953 16363 967 16378
rect 1023 16363 1037 16378
rect 1103 16363 1105 16378
rect 749 16338 765 16363
rect 817 16338 833 16363
rect 885 16338 901 16363
rect 953 16338 969 16363
rect 1021 16338 1037 16363
rect 1089 16338 1105 16363
rect 1157 16338 1173 16363
rect 1225 16338 1241 16363
rect 885 16326 887 16338
rect 953 16326 967 16338
rect 1023 16326 1037 16338
rect 1103 16326 1105 16338
rect 1293 16326 1295 16378
rect 695 16314 727 16326
rect 783 16314 807 16326
rect 863 16314 887 16326
rect 943 16314 967 16326
rect 1023 16314 1047 16326
rect 1103 16314 1127 16326
rect 1183 16314 1207 16326
rect 1263 16314 1295 16326
rect 695 16262 697 16314
rect 885 16282 887 16314
rect 953 16282 967 16314
rect 1023 16282 1037 16314
rect 1103 16282 1105 16314
rect 749 16262 765 16282
rect 817 16262 833 16282
rect 885 16262 901 16282
rect 953 16262 969 16282
rect 1021 16262 1037 16282
rect 1089 16262 1105 16282
rect 1157 16262 1173 16282
rect 1225 16262 1241 16282
rect 1293 16262 1295 16314
rect 695 16257 1295 16262
rect 695 16250 727 16257
rect 783 16250 807 16257
rect 863 16250 887 16257
rect 943 16250 967 16257
rect 1023 16250 1047 16257
rect 1103 16250 1127 16257
rect 1183 16250 1207 16257
rect 1263 16250 1295 16257
rect 695 16198 697 16250
rect 885 16201 887 16250
rect 953 16201 967 16250
rect 1023 16201 1037 16250
rect 1103 16201 1105 16250
rect 749 16198 765 16201
rect 817 16198 833 16201
rect 885 16198 901 16201
rect 953 16198 969 16201
rect 1021 16198 1037 16201
rect 1089 16198 1105 16201
rect 1157 16198 1173 16201
rect 1225 16198 1241 16201
rect 1293 16198 1295 16250
rect 695 15009 1295 16198
rect 695 14957 697 15009
rect 749 15006 765 15009
rect 817 15006 833 15009
rect 885 15006 901 15009
rect 953 15006 969 15009
rect 1021 15006 1037 15009
rect 1089 15006 1105 15009
rect 1157 15006 1173 15009
rect 1225 15006 1241 15009
rect 1293 14957 1295 15009
rect 695 14945 727 14957
rect 1263 14945 1295 14957
rect 695 14893 697 14945
rect 1293 14893 1295 14945
rect 695 14881 727 14893
rect 1263 14881 1295 14893
rect 695 14829 697 14881
rect 1293 14829 1295 14881
rect 695 14817 727 14829
rect 1263 14817 1295 14829
rect 695 14765 697 14817
rect 1293 14765 1295 14817
rect 695 14753 727 14765
rect 1263 14753 1295 14765
rect 695 14701 697 14753
rect 1293 14701 1295 14753
rect 695 14689 727 14701
rect 1263 14689 1295 14701
rect 695 14637 697 14689
rect 1293 14637 1295 14689
rect 695 14625 727 14637
rect 1263 14625 1295 14637
rect 695 14573 697 14625
rect 1293 14573 1295 14625
rect 695 14561 727 14573
rect 1263 14561 1295 14573
rect 695 14509 697 14561
rect 749 14525 765 14550
rect 817 14525 833 14550
rect 885 14525 901 14550
rect 953 14525 969 14550
rect 1021 14525 1037 14550
rect 1089 14525 1105 14550
rect 1157 14525 1173 14550
rect 1225 14525 1241 14550
rect 885 14509 887 14525
rect 953 14509 967 14525
rect 1023 14509 1037 14525
rect 1103 14509 1105 14525
rect 1293 14509 1295 14561
rect 695 14497 727 14509
rect 783 14497 807 14509
rect 863 14497 887 14509
rect 943 14497 967 14509
rect 1023 14497 1047 14509
rect 1103 14497 1127 14509
rect 1183 14497 1207 14509
rect 1263 14497 1295 14509
rect 695 14445 697 14497
rect 885 14469 887 14497
rect 953 14469 967 14497
rect 1023 14469 1037 14497
rect 1103 14469 1105 14497
rect 749 14445 765 14469
rect 817 14445 833 14469
rect 885 14445 901 14469
rect 953 14445 969 14469
rect 1021 14445 1037 14469
rect 1089 14445 1105 14469
rect 1157 14445 1173 14469
rect 1225 14445 1241 14469
rect 1293 14445 1295 14497
rect 695 14444 1295 14445
rect 695 14433 727 14444
rect 783 14433 807 14444
rect 863 14433 887 14444
rect 943 14433 967 14444
rect 1023 14433 1047 14444
rect 1103 14433 1127 14444
rect 1183 14433 1207 14444
rect 1263 14433 1295 14444
rect 695 14381 697 14433
rect 885 14388 887 14433
rect 953 14388 967 14433
rect 1023 14388 1037 14433
rect 1103 14388 1105 14433
rect 749 14381 765 14388
rect 817 14381 833 14388
rect 885 14381 901 14388
rect 953 14381 969 14388
rect 1021 14381 1037 14388
rect 1089 14381 1105 14388
rect 1157 14381 1173 14388
rect 1225 14381 1241 14388
rect 1293 14381 1295 14433
rect 695 14369 1295 14381
rect 695 14317 697 14369
rect 749 14363 765 14369
rect 817 14363 833 14369
rect 885 14363 901 14369
rect 953 14363 969 14369
rect 1021 14363 1037 14369
rect 1089 14363 1105 14369
rect 1157 14363 1173 14369
rect 1225 14363 1241 14369
rect 885 14317 887 14363
rect 953 14317 967 14363
rect 1023 14317 1037 14363
rect 1103 14317 1105 14363
rect 1293 14317 1295 14369
rect 695 14307 727 14317
rect 783 14307 807 14317
rect 863 14307 887 14317
rect 943 14307 967 14317
rect 1023 14307 1047 14317
rect 1103 14307 1127 14317
rect 1183 14307 1207 14317
rect 1263 14307 1295 14317
rect 695 14305 1295 14307
rect 695 14253 697 14305
rect 749 14282 765 14305
rect 817 14282 833 14305
rect 885 14282 901 14305
rect 953 14282 969 14305
rect 1021 14282 1037 14305
rect 1089 14282 1105 14305
rect 1157 14282 1173 14305
rect 1225 14282 1241 14305
rect 885 14253 887 14282
rect 953 14253 967 14282
rect 1023 14253 1037 14282
rect 1103 14253 1105 14282
rect 1293 14253 1295 14305
rect 695 14241 727 14253
rect 783 14241 807 14253
rect 863 14241 887 14253
rect 943 14241 967 14253
rect 1023 14241 1047 14253
rect 1103 14241 1127 14253
rect 1183 14241 1207 14253
rect 1263 14241 1295 14253
rect 695 14189 697 14241
rect 885 14226 887 14241
rect 953 14226 967 14241
rect 1023 14226 1037 14241
rect 1103 14226 1105 14241
rect 749 14201 765 14226
rect 817 14201 833 14226
rect 885 14201 901 14226
rect 953 14201 969 14226
rect 1021 14201 1037 14226
rect 1089 14201 1105 14226
rect 1157 14201 1173 14226
rect 1225 14201 1241 14226
rect 885 14189 887 14201
rect 953 14189 967 14201
rect 1023 14189 1037 14201
rect 1103 14189 1105 14201
rect 1293 14189 1295 14241
rect 695 14177 727 14189
rect 783 14177 807 14189
rect 863 14177 887 14189
rect 943 14177 967 14189
rect 1023 14177 1047 14189
rect 1103 14177 1127 14189
rect 1183 14177 1207 14189
rect 1263 14177 1295 14189
rect 695 14125 697 14177
rect 885 14145 887 14177
rect 953 14145 967 14177
rect 1023 14145 1037 14177
rect 1103 14145 1105 14177
rect 749 14125 765 14145
rect 817 14125 833 14145
rect 885 14125 901 14145
rect 953 14125 969 14145
rect 1021 14125 1037 14145
rect 1089 14125 1105 14145
rect 1157 14125 1173 14145
rect 1225 14125 1241 14145
rect 1293 14125 1295 14177
rect 695 14120 1295 14125
rect 695 14113 727 14120
rect 783 14113 807 14120
rect 863 14113 887 14120
rect 943 14113 967 14120
rect 1023 14113 1047 14120
rect 1103 14113 1127 14120
rect 1183 14113 1207 14120
rect 1263 14113 1295 14120
rect 695 14061 697 14113
rect 885 14064 887 14113
rect 953 14064 967 14113
rect 1023 14064 1037 14113
rect 1103 14064 1105 14113
rect 749 14061 765 14064
rect 817 14061 833 14064
rect 885 14061 901 14064
rect 953 14061 969 14064
rect 1021 14061 1037 14064
rect 1089 14061 1105 14064
rect 1157 14061 1173 14064
rect 1225 14061 1241 14064
rect 1293 14061 1295 14113
rect 115 13701 171 13707
rect 115 13698 117 13701
rect 169 13698 171 13701
rect 115 13633 171 13642
rect 115 13617 117 13633
rect 169 13617 171 13633
rect 115 13536 117 13561
rect 169 13536 171 13561
rect 115 13455 117 13480
rect 169 13455 171 13480
rect 115 13375 117 13399
rect 169 13375 171 13399
rect 115 13374 171 13375
rect 115 13306 117 13318
rect 169 13306 171 13318
rect 115 13292 171 13306
rect 115 13220 171 13236
rect 115 13210 117 13220
rect 169 13210 171 13220
rect 115 13151 171 13154
rect 115 13128 117 13151
rect 169 13128 171 13151
rect 115 13046 117 13072
rect 169 13046 171 13072
rect 115 12964 117 12990
rect 169 12964 171 12990
rect 115 12892 117 12908
rect 169 12892 171 12908
rect 115 12882 171 12892
rect 115 12823 117 12826
rect 169 12823 171 12826
rect 115 12817 171 12823
rect 695 12907 1295 14061
rect 695 12855 697 12907
rect 749 12904 765 12907
rect 817 12904 833 12907
rect 885 12904 901 12907
rect 953 12904 969 12907
rect 1021 12904 1037 12907
rect 1089 12904 1105 12907
rect 1157 12904 1173 12907
rect 1225 12904 1241 12907
rect 1293 12855 1295 12907
rect 695 12843 727 12855
rect 1263 12843 1295 12855
rect 695 12791 697 12843
rect 1293 12791 1295 12843
rect 695 12779 727 12791
rect 1263 12779 1295 12791
rect 695 12727 697 12779
rect 1293 12727 1295 12779
rect 695 12715 727 12727
rect 1263 12715 1295 12727
rect 695 12663 697 12715
rect 1293 12663 1295 12715
rect 695 12651 727 12663
rect 1263 12651 1295 12663
rect 695 12599 697 12651
rect 1293 12599 1295 12651
rect 695 12587 727 12599
rect 1263 12587 1295 12599
rect 695 12535 697 12587
rect 1293 12535 1295 12587
rect 695 12523 727 12535
rect 1263 12523 1295 12535
rect 695 12471 697 12523
rect 1293 12471 1295 12523
rect 695 12459 727 12471
rect 1263 12459 1295 12471
rect 695 12407 697 12459
rect 749 12423 765 12448
rect 817 12423 833 12448
rect 885 12423 901 12448
rect 953 12423 969 12448
rect 1021 12423 1037 12448
rect 1089 12423 1105 12448
rect 1157 12423 1173 12448
rect 1225 12423 1241 12448
rect 885 12407 887 12423
rect 953 12407 967 12423
rect 1023 12407 1037 12423
rect 1103 12407 1105 12423
rect 1293 12407 1295 12459
rect 695 12395 727 12407
rect 783 12395 807 12407
rect 863 12395 887 12407
rect 943 12395 967 12407
rect 1023 12395 1047 12407
rect 1103 12395 1127 12407
rect 1183 12395 1207 12407
rect 1263 12395 1295 12407
rect 695 12343 697 12395
rect 885 12367 887 12395
rect 953 12367 967 12395
rect 1023 12367 1037 12395
rect 1103 12367 1105 12395
rect 749 12343 765 12367
rect 817 12343 833 12367
rect 885 12343 901 12367
rect 953 12343 969 12367
rect 1021 12343 1037 12367
rect 1089 12343 1105 12367
rect 1157 12343 1173 12367
rect 1225 12343 1241 12367
rect 1293 12343 1295 12395
rect 695 12342 1295 12343
rect 695 12331 727 12342
rect 783 12331 807 12342
rect 863 12331 887 12342
rect 943 12331 967 12342
rect 1023 12331 1047 12342
rect 1103 12331 1127 12342
rect 1183 12331 1207 12342
rect 1263 12331 1295 12342
rect 695 12279 697 12331
rect 885 12286 887 12331
rect 953 12286 967 12331
rect 1023 12286 1037 12331
rect 1103 12286 1105 12331
rect 749 12279 765 12286
rect 817 12279 833 12286
rect 885 12279 901 12286
rect 953 12279 969 12286
rect 1021 12279 1037 12286
rect 1089 12279 1105 12286
rect 1157 12279 1173 12286
rect 1225 12279 1241 12286
rect 1293 12279 1295 12331
rect 695 12267 1295 12279
rect 695 12215 697 12267
rect 749 12261 765 12267
rect 817 12261 833 12267
rect 885 12261 901 12267
rect 953 12261 969 12267
rect 1021 12261 1037 12267
rect 1089 12261 1105 12267
rect 1157 12261 1173 12267
rect 1225 12261 1241 12267
rect 885 12215 887 12261
rect 953 12215 967 12261
rect 1023 12215 1037 12261
rect 1103 12215 1105 12261
rect 1293 12215 1295 12267
rect 695 12205 727 12215
rect 783 12205 807 12215
rect 863 12205 887 12215
rect 943 12205 967 12215
rect 1023 12205 1047 12215
rect 1103 12205 1127 12215
rect 1183 12205 1207 12215
rect 1263 12205 1295 12215
rect 695 12203 1295 12205
rect 695 12151 697 12203
rect 749 12180 765 12203
rect 817 12180 833 12203
rect 885 12180 901 12203
rect 953 12180 969 12203
rect 1021 12180 1037 12203
rect 1089 12180 1105 12203
rect 1157 12180 1173 12203
rect 1225 12180 1241 12203
rect 885 12151 887 12180
rect 953 12151 967 12180
rect 1023 12151 1037 12180
rect 1103 12151 1105 12180
rect 1293 12151 1295 12203
rect 695 12139 727 12151
rect 783 12139 807 12151
rect 863 12139 887 12151
rect 943 12139 967 12151
rect 1023 12139 1047 12151
rect 1103 12139 1127 12151
rect 1183 12139 1207 12151
rect 1263 12139 1295 12151
rect 695 12087 697 12139
rect 885 12124 887 12139
rect 953 12124 967 12139
rect 1023 12124 1037 12139
rect 1103 12124 1105 12139
rect 749 12099 765 12124
rect 817 12099 833 12124
rect 885 12099 901 12124
rect 953 12099 969 12124
rect 1021 12099 1037 12124
rect 1089 12099 1105 12124
rect 1157 12099 1173 12124
rect 1225 12099 1241 12124
rect 885 12087 887 12099
rect 953 12087 967 12099
rect 1023 12087 1037 12099
rect 1103 12087 1105 12099
rect 1293 12087 1295 12139
rect 695 12075 727 12087
rect 783 12075 807 12087
rect 863 12075 887 12087
rect 943 12075 967 12087
rect 1023 12075 1047 12087
rect 1103 12075 1127 12087
rect 1183 12075 1207 12087
rect 1263 12075 1295 12087
rect 695 12023 697 12075
rect 885 12043 887 12075
rect 953 12043 967 12075
rect 1023 12043 1037 12075
rect 1103 12043 1105 12075
rect 749 12023 765 12043
rect 817 12023 833 12043
rect 885 12023 901 12043
rect 953 12023 969 12043
rect 1021 12023 1037 12043
rect 1089 12023 1105 12043
rect 1157 12023 1173 12043
rect 1225 12023 1241 12043
rect 1293 12023 1295 12075
rect 695 12018 1295 12023
rect 695 12011 727 12018
rect 783 12011 807 12018
rect 863 12011 887 12018
rect 943 12011 967 12018
rect 1023 12011 1047 12018
rect 1103 12011 1127 12018
rect 1183 12011 1207 12018
rect 1263 12011 1295 12018
rect 695 11959 697 12011
rect 885 11962 887 12011
rect 953 11962 967 12011
rect 1023 11962 1037 12011
rect 1103 11962 1105 12011
rect 749 11959 765 11962
rect 817 11959 833 11962
rect 885 11959 901 11962
rect 953 11959 969 11962
rect 1021 11959 1037 11962
rect 1089 11959 1105 11962
rect 1157 11959 1173 11962
rect 1225 11959 1241 11962
rect 1293 11959 1295 12011
rect 695 10813 1295 11959
rect 695 10761 697 10813
rect 749 10810 765 10813
rect 817 10810 833 10813
rect 885 10810 901 10813
rect 953 10810 969 10813
rect 1021 10810 1037 10813
rect 1089 10810 1105 10813
rect 1157 10810 1173 10813
rect 1225 10810 1241 10813
rect 1293 10761 1295 10813
rect 695 10749 727 10761
rect 1263 10749 1295 10761
rect 695 10697 697 10749
rect 1293 10697 1295 10749
rect 695 10685 727 10697
rect 1263 10685 1295 10697
rect 695 10633 697 10685
rect 1293 10633 1295 10685
rect 695 10621 727 10633
rect 1263 10621 1295 10633
rect 695 10569 697 10621
rect 1293 10569 1295 10621
rect 695 10557 727 10569
rect 1263 10557 1295 10569
rect 695 10505 697 10557
rect 1293 10505 1295 10557
rect 695 10493 727 10505
rect 1263 10493 1295 10505
rect 695 10441 697 10493
rect 1293 10441 1295 10493
rect 695 10429 727 10441
rect 1263 10429 1295 10441
rect 695 10377 697 10429
rect 1293 10377 1295 10429
rect 695 10365 727 10377
rect 1263 10365 1295 10377
rect 695 10313 697 10365
rect 749 10329 765 10354
rect 817 10329 833 10354
rect 885 10329 901 10354
rect 953 10329 969 10354
rect 1021 10329 1037 10354
rect 1089 10329 1105 10354
rect 1157 10329 1173 10354
rect 1225 10329 1241 10354
rect 885 10313 887 10329
rect 953 10313 967 10329
rect 1023 10313 1037 10329
rect 1103 10313 1105 10329
rect 1293 10313 1295 10365
rect 695 10301 727 10313
rect 783 10301 807 10313
rect 863 10301 887 10313
rect 943 10301 967 10313
rect 1023 10301 1047 10313
rect 1103 10301 1127 10313
rect 1183 10301 1207 10313
rect 1263 10301 1295 10313
rect 695 10249 697 10301
rect 885 10273 887 10301
rect 953 10273 967 10301
rect 1023 10273 1037 10301
rect 1103 10273 1105 10301
rect 749 10249 765 10273
rect 817 10249 833 10273
rect 885 10249 901 10273
rect 953 10249 969 10273
rect 1021 10249 1037 10273
rect 1089 10249 1105 10273
rect 1157 10249 1173 10273
rect 1225 10249 1241 10273
rect 1293 10249 1295 10301
rect 695 10248 1295 10249
rect 695 10237 727 10248
rect 783 10237 807 10248
rect 863 10237 887 10248
rect 943 10237 967 10248
rect 1023 10237 1047 10248
rect 1103 10237 1127 10248
rect 1183 10237 1207 10248
rect 1263 10237 1295 10248
rect 695 10185 697 10237
rect 885 10192 887 10237
rect 953 10192 967 10237
rect 1023 10192 1037 10237
rect 1103 10192 1105 10237
rect 749 10185 765 10192
rect 817 10185 833 10192
rect 885 10185 901 10192
rect 953 10185 969 10192
rect 1021 10185 1037 10192
rect 1089 10185 1105 10192
rect 1157 10185 1173 10192
rect 1225 10185 1241 10192
rect 1293 10185 1295 10237
rect 695 10173 1295 10185
rect 695 10121 697 10173
rect 749 10167 765 10173
rect 817 10167 833 10173
rect 885 10167 901 10173
rect 953 10167 969 10173
rect 1021 10167 1037 10173
rect 1089 10167 1105 10173
rect 1157 10167 1173 10173
rect 1225 10167 1241 10173
rect 885 10121 887 10167
rect 953 10121 967 10167
rect 1023 10121 1037 10167
rect 1103 10121 1105 10167
rect 1293 10121 1295 10173
rect 695 10111 727 10121
rect 783 10111 807 10121
rect 863 10111 887 10121
rect 943 10111 967 10121
rect 1023 10111 1047 10121
rect 1103 10111 1127 10121
rect 1183 10111 1207 10121
rect 1263 10111 1295 10121
rect 695 10109 1295 10111
rect 695 10057 697 10109
rect 749 10086 765 10109
rect 817 10086 833 10109
rect 885 10086 901 10109
rect 953 10086 969 10109
rect 1021 10086 1037 10109
rect 1089 10086 1105 10109
rect 1157 10086 1173 10109
rect 1225 10086 1241 10109
rect 885 10057 887 10086
rect 953 10057 967 10086
rect 1023 10057 1037 10086
rect 1103 10057 1105 10086
rect 1293 10057 1295 10109
rect 695 10045 727 10057
rect 783 10045 807 10057
rect 863 10045 887 10057
rect 943 10045 967 10057
rect 1023 10045 1047 10057
rect 1103 10045 1127 10057
rect 1183 10045 1207 10057
rect 1263 10045 1295 10057
rect 695 9993 697 10045
rect 885 10030 887 10045
rect 953 10030 967 10045
rect 1023 10030 1037 10045
rect 1103 10030 1105 10045
rect 749 10005 765 10030
rect 817 10005 833 10030
rect 885 10005 901 10030
rect 953 10005 969 10030
rect 1021 10005 1037 10030
rect 1089 10005 1105 10030
rect 1157 10005 1173 10030
rect 1225 10005 1241 10030
rect 885 9993 887 10005
rect 953 9993 967 10005
rect 1023 9993 1037 10005
rect 1103 9993 1105 10005
rect 1293 9993 1295 10045
rect 695 9981 727 9993
rect 783 9981 807 9993
rect 863 9981 887 9993
rect 943 9981 967 9993
rect 1023 9981 1047 9993
rect 1103 9981 1127 9993
rect 1183 9981 1207 9993
rect 1263 9981 1295 9993
rect 695 9929 697 9981
rect 885 9949 887 9981
rect 953 9949 967 9981
rect 1023 9949 1037 9981
rect 1103 9949 1105 9981
rect 749 9929 765 9949
rect 817 9929 833 9949
rect 885 9929 901 9949
rect 953 9929 969 9949
rect 1021 9929 1037 9949
rect 1089 9929 1105 9949
rect 1157 9929 1173 9949
rect 1225 9929 1241 9949
rect 1293 9929 1295 9981
rect 695 9924 1295 9929
rect 695 9917 727 9924
rect 783 9917 807 9924
rect 863 9917 887 9924
rect 943 9917 967 9924
rect 1023 9917 1047 9924
rect 1103 9917 1127 9924
rect 1183 9917 1207 9924
rect 1263 9917 1295 9924
rect 695 9865 697 9917
rect 885 9868 887 9917
rect 953 9868 967 9917
rect 1023 9868 1037 9917
rect 1103 9868 1105 9917
rect 749 9865 765 9868
rect 817 9865 833 9868
rect 885 9865 901 9868
rect 953 9865 969 9868
rect 1021 9865 1037 9868
rect 1089 9865 1105 9868
rect 1157 9865 1173 9868
rect 1225 9865 1241 9868
rect 1293 9865 1295 9917
rect 695 8611 1295 9865
rect 695 8559 697 8611
rect 749 8608 765 8611
rect 817 8608 833 8611
rect 885 8608 901 8611
rect 953 8608 969 8611
rect 1021 8608 1037 8611
rect 1089 8608 1105 8611
rect 1157 8608 1173 8611
rect 1225 8608 1241 8611
rect 1293 8559 1295 8611
rect 695 8547 727 8559
rect 1263 8547 1295 8559
rect 695 8495 697 8547
rect 1293 8495 1295 8547
rect 695 8483 727 8495
rect 1263 8483 1295 8495
rect 695 8431 697 8483
rect 1293 8431 1295 8483
rect 695 8419 727 8431
rect 1263 8419 1295 8431
rect 695 8367 697 8419
rect 1293 8367 1295 8419
rect 695 8355 727 8367
rect 1263 8355 1295 8367
rect 695 8303 697 8355
rect 1293 8303 1295 8355
rect 695 8291 727 8303
rect 1263 8291 1295 8303
rect 695 8239 697 8291
rect 1293 8239 1295 8291
rect 695 8227 727 8239
rect 1263 8227 1295 8239
rect 695 8175 697 8227
rect 1293 8175 1295 8227
rect 695 8163 727 8175
rect 1263 8163 1295 8175
rect 695 8111 697 8163
rect 749 8127 765 8152
rect 817 8127 833 8152
rect 885 8127 901 8152
rect 953 8127 969 8152
rect 1021 8127 1037 8152
rect 1089 8127 1105 8152
rect 1157 8127 1173 8152
rect 1225 8127 1241 8152
rect 885 8111 887 8127
rect 953 8111 967 8127
rect 1023 8111 1037 8127
rect 1103 8111 1105 8127
rect 1293 8111 1295 8163
rect 695 8099 727 8111
rect 783 8099 807 8111
rect 863 8099 887 8111
rect 943 8099 967 8111
rect 1023 8099 1047 8111
rect 1103 8099 1127 8111
rect 1183 8099 1207 8111
rect 1263 8099 1295 8111
rect 695 8047 697 8099
rect 885 8071 887 8099
rect 953 8071 967 8099
rect 1023 8071 1037 8099
rect 1103 8071 1105 8099
rect 749 8047 765 8071
rect 817 8047 833 8071
rect 885 8047 901 8071
rect 953 8047 969 8071
rect 1021 8047 1037 8071
rect 1089 8047 1105 8071
rect 1157 8047 1173 8071
rect 1225 8047 1241 8071
rect 1293 8047 1295 8099
rect 695 8046 1295 8047
rect 695 8035 727 8046
rect 783 8035 807 8046
rect 863 8035 887 8046
rect 943 8035 967 8046
rect 1023 8035 1047 8046
rect 1103 8035 1127 8046
rect 1183 8035 1207 8046
rect 1263 8035 1295 8046
rect 695 7983 697 8035
rect 885 7990 887 8035
rect 953 7990 967 8035
rect 1023 7990 1037 8035
rect 1103 7990 1105 8035
rect 749 7983 765 7990
rect 817 7983 833 7990
rect 885 7983 901 7990
rect 953 7983 969 7990
rect 1021 7983 1037 7990
rect 1089 7983 1105 7990
rect 1157 7983 1173 7990
rect 1225 7983 1241 7990
rect 1293 7983 1295 8035
rect 695 7971 1295 7983
rect 695 7919 697 7971
rect 749 7965 765 7971
rect 817 7965 833 7971
rect 885 7965 901 7971
rect 953 7965 969 7971
rect 1021 7965 1037 7971
rect 1089 7965 1105 7971
rect 1157 7965 1173 7971
rect 1225 7965 1241 7971
rect 885 7919 887 7965
rect 953 7919 967 7965
rect 1023 7919 1037 7965
rect 1103 7919 1105 7965
rect 1293 7919 1295 7971
rect 695 7909 727 7919
rect 783 7909 807 7919
rect 863 7909 887 7919
rect 943 7909 967 7919
rect 1023 7909 1047 7919
rect 1103 7909 1127 7919
rect 1183 7909 1207 7919
rect 1263 7909 1295 7919
rect 695 7907 1295 7909
rect 695 7855 697 7907
rect 749 7884 765 7907
rect 817 7884 833 7907
rect 885 7884 901 7907
rect 953 7884 969 7907
rect 1021 7884 1037 7907
rect 1089 7884 1105 7907
rect 1157 7884 1173 7907
rect 1225 7884 1241 7907
rect 885 7855 887 7884
rect 953 7855 967 7884
rect 1023 7855 1037 7884
rect 1103 7855 1105 7884
rect 1293 7855 1295 7907
rect 695 7843 727 7855
rect 783 7843 807 7855
rect 863 7843 887 7855
rect 943 7843 967 7855
rect 1023 7843 1047 7855
rect 1103 7843 1127 7855
rect 1183 7843 1207 7855
rect 1263 7843 1295 7855
rect 695 7791 697 7843
rect 885 7828 887 7843
rect 953 7828 967 7843
rect 1023 7828 1037 7843
rect 1103 7828 1105 7843
rect 749 7803 765 7828
rect 817 7803 833 7828
rect 885 7803 901 7828
rect 953 7803 969 7828
rect 1021 7803 1037 7828
rect 1089 7803 1105 7828
rect 1157 7803 1173 7828
rect 1225 7803 1241 7828
rect 885 7791 887 7803
rect 953 7791 967 7803
rect 1023 7791 1037 7803
rect 1103 7791 1105 7803
rect 1293 7791 1295 7843
rect 695 7779 727 7791
rect 783 7779 807 7791
rect 863 7779 887 7791
rect 943 7779 967 7791
rect 1023 7779 1047 7791
rect 1103 7779 1127 7791
rect 1183 7779 1207 7791
rect 1263 7779 1295 7791
rect 695 7727 697 7779
rect 885 7747 887 7779
rect 953 7747 967 7779
rect 1023 7747 1037 7779
rect 1103 7747 1105 7779
rect 749 7727 765 7747
rect 817 7727 833 7747
rect 885 7727 901 7747
rect 953 7727 969 7747
rect 1021 7727 1037 7747
rect 1089 7727 1105 7747
rect 1157 7727 1173 7747
rect 1225 7727 1241 7747
rect 1293 7727 1295 7779
rect 695 7722 1295 7727
rect 695 7715 727 7722
rect 783 7715 807 7722
rect 863 7715 887 7722
rect 943 7715 967 7722
rect 1023 7715 1047 7722
rect 1103 7715 1127 7722
rect 1183 7715 1207 7722
rect 1263 7715 1295 7722
rect 695 7663 697 7715
rect 885 7666 887 7715
rect 953 7666 967 7715
rect 1023 7666 1037 7715
rect 1103 7666 1105 7715
rect 749 7663 765 7666
rect 817 7663 833 7666
rect 885 7663 901 7666
rect 953 7663 969 7666
rect 1021 7663 1037 7666
rect 1089 7663 1105 7666
rect 1157 7663 1173 7666
rect 1225 7663 1241 7666
rect 1293 7663 1295 7715
rect 695 6501 1295 7663
rect 695 6449 697 6501
rect 749 6498 765 6501
rect 817 6498 833 6501
rect 885 6498 901 6501
rect 953 6498 969 6501
rect 1021 6498 1037 6501
rect 1089 6498 1105 6501
rect 1157 6498 1173 6501
rect 1225 6498 1241 6501
rect 1293 6449 1295 6501
rect 695 6437 727 6449
rect 1263 6437 1295 6449
rect 695 6385 697 6437
rect 1293 6385 1295 6437
rect 695 6373 727 6385
rect 1263 6373 1295 6385
rect 695 6321 697 6373
rect 1293 6321 1295 6373
rect 695 6309 727 6321
rect 1263 6309 1295 6321
rect 695 6257 697 6309
rect 1293 6257 1295 6309
rect 695 6245 727 6257
rect 1263 6245 1295 6257
rect 695 6193 697 6245
rect 1293 6193 1295 6245
rect 695 6181 727 6193
rect 1263 6181 1295 6193
rect 695 6129 697 6181
rect 1293 6129 1295 6181
rect 695 6117 727 6129
rect 1263 6117 1295 6129
rect 695 6065 697 6117
rect 1293 6065 1295 6117
rect 695 6053 727 6065
rect 1263 6053 1295 6065
rect 695 6001 697 6053
rect 749 6017 765 6042
rect 817 6017 833 6042
rect 885 6017 901 6042
rect 953 6017 969 6042
rect 1021 6017 1037 6042
rect 1089 6017 1105 6042
rect 1157 6017 1173 6042
rect 1225 6017 1241 6042
rect 885 6001 887 6017
rect 953 6001 967 6017
rect 1023 6001 1037 6017
rect 1103 6001 1105 6017
rect 1293 6001 1295 6053
rect 695 5989 727 6001
rect 783 5989 807 6001
rect 863 5989 887 6001
rect 943 5989 967 6001
rect 1023 5989 1047 6001
rect 1103 5989 1127 6001
rect 1183 5989 1207 6001
rect 1263 5989 1295 6001
rect 695 5937 697 5989
rect 885 5961 887 5989
rect 953 5961 967 5989
rect 1023 5961 1037 5989
rect 1103 5961 1105 5989
rect 749 5937 765 5961
rect 817 5937 833 5961
rect 885 5937 901 5961
rect 953 5937 969 5961
rect 1021 5937 1037 5961
rect 1089 5937 1105 5961
rect 1157 5937 1173 5961
rect 1225 5937 1241 5961
rect 1293 5937 1295 5989
rect 695 5936 1295 5937
rect 695 5925 727 5936
rect 783 5925 807 5936
rect 863 5925 887 5936
rect 943 5925 967 5936
rect 1023 5925 1047 5936
rect 1103 5925 1127 5936
rect 1183 5925 1207 5936
rect 1263 5925 1295 5936
rect 695 5873 697 5925
rect 885 5880 887 5925
rect 953 5880 967 5925
rect 1023 5880 1037 5925
rect 1103 5880 1105 5925
rect 749 5873 765 5880
rect 817 5873 833 5880
rect 885 5873 901 5880
rect 953 5873 969 5880
rect 1021 5873 1037 5880
rect 1089 5873 1105 5880
rect 1157 5873 1173 5880
rect 1225 5873 1241 5880
rect 1293 5873 1295 5925
rect 695 5861 1295 5873
rect 695 5809 697 5861
rect 749 5855 765 5861
rect 817 5855 833 5861
rect 885 5855 901 5861
rect 953 5855 969 5861
rect 1021 5855 1037 5861
rect 1089 5855 1105 5861
rect 1157 5855 1173 5861
rect 1225 5855 1241 5861
rect 885 5809 887 5855
rect 953 5809 967 5855
rect 1023 5809 1037 5855
rect 1103 5809 1105 5855
rect 1293 5809 1295 5861
rect 695 5799 727 5809
rect 783 5799 807 5809
rect 863 5799 887 5809
rect 943 5799 967 5809
rect 1023 5799 1047 5809
rect 1103 5799 1127 5809
rect 1183 5799 1207 5809
rect 1263 5799 1295 5809
rect 695 5797 1295 5799
rect 695 5745 697 5797
rect 749 5774 765 5797
rect 817 5774 833 5797
rect 885 5774 901 5797
rect 953 5774 969 5797
rect 1021 5774 1037 5797
rect 1089 5774 1105 5797
rect 1157 5774 1173 5797
rect 1225 5774 1241 5797
rect 885 5745 887 5774
rect 953 5745 967 5774
rect 1023 5745 1037 5774
rect 1103 5745 1105 5774
rect 1293 5745 1295 5797
rect 695 5733 727 5745
rect 783 5733 807 5745
rect 863 5733 887 5745
rect 943 5733 967 5745
rect 1023 5733 1047 5745
rect 1103 5733 1127 5745
rect 1183 5733 1207 5745
rect 1263 5733 1295 5745
rect 695 5681 697 5733
rect 885 5718 887 5733
rect 953 5718 967 5733
rect 1023 5718 1037 5733
rect 1103 5718 1105 5733
rect 749 5693 765 5718
rect 817 5693 833 5718
rect 885 5693 901 5718
rect 953 5693 969 5718
rect 1021 5693 1037 5718
rect 1089 5693 1105 5718
rect 1157 5693 1173 5718
rect 1225 5693 1241 5718
rect 885 5681 887 5693
rect 953 5681 967 5693
rect 1023 5681 1037 5693
rect 1103 5681 1105 5693
rect 1293 5681 1295 5733
rect 695 5669 727 5681
rect 783 5669 807 5681
rect 863 5669 887 5681
rect 943 5669 967 5681
rect 1023 5669 1047 5681
rect 1103 5669 1127 5681
rect 1183 5669 1207 5681
rect 1263 5669 1295 5681
rect 695 5617 697 5669
rect 885 5637 887 5669
rect 953 5637 967 5669
rect 1023 5637 1037 5669
rect 1103 5637 1105 5669
rect 749 5617 765 5637
rect 817 5617 833 5637
rect 885 5617 901 5637
rect 953 5617 969 5637
rect 1021 5617 1037 5637
rect 1089 5617 1105 5637
rect 1157 5617 1173 5637
rect 1225 5617 1241 5637
rect 1293 5617 1295 5669
rect 695 5612 1295 5617
rect 695 5605 727 5612
rect 783 5605 807 5612
rect 863 5605 887 5612
rect 943 5605 967 5612
rect 1023 5605 1047 5612
rect 1103 5605 1127 5612
rect 1183 5605 1207 5612
rect 1263 5605 1295 5612
rect 695 5553 697 5605
rect 885 5556 887 5605
rect 953 5556 967 5605
rect 1023 5556 1037 5605
rect 1103 5556 1105 5605
rect 749 5553 765 5556
rect 817 5553 833 5556
rect 885 5553 901 5556
rect 953 5553 969 5556
rect 1021 5553 1037 5556
rect 1089 5553 1105 5556
rect 1157 5553 1173 5556
rect 1225 5553 1241 5556
rect 1293 5553 1295 5605
rect 695 4437 1295 5553
rect 695 4385 697 4437
rect 749 4434 765 4437
rect 817 4434 833 4437
rect 885 4434 901 4437
rect 953 4434 969 4437
rect 1021 4434 1037 4437
rect 1089 4434 1105 4437
rect 1157 4434 1173 4437
rect 1225 4434 1241 4437
rect 1293 4385 1295 4437
rect 695 4373 727 4385
rect 1263 4373 1295 4385
rect 695 4321 697 4373
rect 1293 4321 1295 4373
rect 695 4309 727 4321
rect 1263 4309 1295 4321
rect 695 4257 697 4309
rect 1293 4257 1295 4309
rect 695 4245 727 4257
rect 1263 4245 1295 4257
rect 695 4193 697 4245
rect 1293 4193 1295 4245
rect 695 4181 727 4193
rect 1263 4181 1295 4193
rect 695 4129 697 4181
rect 1293 4129 1295 4181
rect 695 4117 727 4129
rect 1263 4117 1295 4129
rect 695 4065 697 4117
rect 1293 4065 1295 4117
rect 695 4053 727 4065
rect 1263 4053 1295 4065
rect 695 4001 697 4053
rect 1293 4001 1295 4053
rect 695 3989 727 4001
rect 1263 3989 1295 4001
rect 695 3937 697 3989
rect 749 3953 765 3978
rect 817 3953 833 3978
rect 885 3953 901 3978
rect 953 3953 969 3978
rect 1021 3953 1037 3978
rect 1089 3953 1105 3978
rect 1157 3953 1173 3978
rect 1225 3953 1241 3978
rect 885 3937 887 3953
rect 953 3937 967 3953
rect 1023 3937 1037 3953
rect 1103 3937 1105 3953
rect 1293 3937 1295 3989
rect 695 3925 727 3937
rect 783 3925 807 3937
rect 863 3925 887 3937
rect 943 3925 967 3937
rect 1023 3925 1047 3937
rect 1103 3925 1127 3937
rect 1183 3925 1207 3937
rect 1263 3925 1295 3937
rect 695 3873 697 3925
rect 885 3897 887 3925
rect 953 3897 967 3925
rect 1023 3897 1037 3925
rect 1103 3897 1105 3925
rect 749 3873 765 3897
rect 817 3873 833 3897
rect 885 3873 901 3897
rect 953 3873 969 3897
rect 1021 3873 1037 3897
rect 1089 3873 1105 3897
rect 1157 3873 1173 3897
rect 1225 3873 1241 3897
rect 1293 3873 1295 3925
rect 695 3872 1295 3873
rect 695 3861 727 3872
rect 783 3861 807 3872
rect 863 3861 887 3872
rect 943 3861 967 3872
rect 1023 3861 1047 3872
rect 1103 3861 1127 3872
rect 1183 3861 1207 3872
rect 1263 3861 1295 3872
rect 695 3809 697 3861
rect 885 3816 887 3861
rect 953 3816 967 3861
rect 1023 3816 1037 3861
rect 1103 3816 1105 3861
rect 749 3809 765 3816
rect 817 3809 833 3816
rect 885 3809 901 3816
rect 953 3809 969 3816
rect 1021 3809 1037 3816
rect 1089 3809 1105 3816
rect 1157 3809 1173 3816
rect 1225 3809 1241 3816
rect 1293 3809 1295 3861
rect 695 3797 1295 3809
rect 695 3745 697 3797
rect 749 3791 765 3797
rect 817 3791 833 3797
rect 885 3791 901 3797
rect 953 3791 969 3797
rect 1021 3791 1037 3797
rect 1089 3791 1105 3797
rect 1157 3791 1173 3797
rect 1225 3791 1241 3797
rect 885 3745 887 3791
rect 953 3745 967 3791
rect 1023 3745 1037 3791
rect 1103 3745 1105 3791
rect 1293 3745 1295 3797
rect 695 3735 727 3745
rect 783 3735 807 3745
rect 863 3735 887 3745
rect 943 3735 967 3745
rect 1023 3735 1047 3745
rect 1103 3735 1127 3745
rect 1183 3735 1207 3745
rect 1263 3735 1295 3745
rect 695 3733 1295 3735
rect 695 3681 697 3733
rect 749 3710 765 3733
rect 817 3710 833 3733
rect 885 3710 901 3733
rect 953 3710 969 3733
rect 1021 3710 1037 3733
rect 1089 3710 1105 3733
rect 1157 3710 1173 3733
rect 1225 3710 1241 3733
rect 885 3681 887 3710
rect 953 3681 967 3710
rect 1023 3681 1037 3710
rect 1103 3681 1105 3710
rect 1293 3681 1295 3733
rect 695 3669 727 3681
rect 783 3669 807 3681
rect 863 3669 887 3681
rect 943 3669 967 3681
rect 1023 3669 1047 3681
rect 1103 3669 1127 3681
rect 1183 3669 1207 3681
rect 1263 3669 1295 3681
rect 695 3617 697 3669
rect 885 3654 887 3669
rect 953 3654 967 3669
rect 1023 3654 1037 3669
rect 1103 3654 1105 3669
rect 749 3629 765 3654
rect 817 3629 833 3654
rect 885 3629 901 3654
rect 953 3629 969 3654
rect 1021 3629 1037 3654
rect 1089 3629 1105 3654
rect 1157 3629 1173 3654
rect 1225 3629 1241 3654
rect 885 3617 887 3629
rect 953 3617 967 3629
rect 1023 3617 1037 3629
rect 1103 3617 1105 3629
rect 1293 3617 1295 3669
rect 695 3605 727 3617
rect 783 3605 807 3617
rect 863 3605 887 3617
rect 943 3605 967 3617
rect 1023 3605 1047 3617
rect 1103 3605 1127 3617
rect 1183 3605 1207 3617
rect 1263 3605 1295 3617
rect 695 3553 697 3605
rect 885 3573 887 3605
rect 953 3573 967 3605
rect 1023 3573 1037 3605
rect 1103 3573 1105 3605
rect 749 3553 765 3573
rect 817 3553 833 3573
rect 885 3553 901 3573
rect 953 3553 969 3573
rect 1021 3553 1037 3573
rect 1089 3553 1105 3573
rect 1157 3553 1173 3573
rect 1225 3553 1241 3573
rect 1293 3553 1295 3605
rect 695 3548 1295 3553
rect 695 3541 727 3548
rect 783 3541 807 3548
rect 863 3541 887 3548
rect 943 3541 967 3548
rect 1023 3541 1047 3548
rect 1103 3541 1127 3548
rect 1183 3541 1207 3548
rect 1263 3541 1295 3548
rect 695 3489 697 3541
rect 885 3492 887 3541
rect 953 3492 967 3541
rect 1023 3492 1037 3541
rect 1103 3492 1105 3541
rect 749 3489 765 3492
rect 817 3489 833 3492
rect 885 3489 901 3492
rect 953 3489 969 3492
rect 1021 3489 1037 3492
rect 1089 3489 1105 3492
rect 1157 3489 1173 3492
rect 1225 3489 1241 3492
rect 1293 3489 1295 3541
rect 695 2243 1295 3489
rect 695 2191 697 2243
rect 749 2240 765 2243
rect 817 2240 833 2243
rect 885 2240 901 2243
rect 953 2240 969 2243
rect 1021 2240 1037 2243
rect 1089 2240 1105 2243
rect 1157 2240 1173 2243
rect 1225 2240 1241 2243
rect 1293 2191 1295 2243
rect 695 2179 727 2191
rect 1263 2179 1295 2191
rect 695 2127 697 2179
rect 1293 2127 1295 2179
rect 695 2115 727 2127
rect 1263 2115 1295 2127
rect 695 2063 697 2115
rect 1293 2063 1295 2115
rect 695 2051 727 2063
rect 1263 2051 1295 2063
rect 695 1999 697 2051
rect 1293 1999 1295 2051
rect 695 1987 727 1999
rect 1263 1987 1295 1999
rect 695 1935 697 1987
rect 1293 1935 1295 1987
rect 695 1923 727 1935
rect 1263 1923 1295 1935
rect 695 1871 697 1923
rect 1293 1871 1295 1923
rect 695 1859 727 1871
rect 1263 1859 1295 1871
rect 695 1807 697 1859
rect 1293 1807 1295 1859
rect 695 1795 727 1807
rect 1263 1795 1295 1807
rect 695 1743 697 1795
rect 749 1759 765 1784
rect 817 1759 833 1784
rect 885 1759 901 1784
rect 953 1759 969 1784
rect 1021 1759 1037 1784
rect 1089 1759 1105 1784
rect 1157 1759 1173 1784
rect 1225 1759 1241 1784
rect 885 1743 887 1759
rect 953 1743 967 1759
rect 1023 1743 1037 1759
rect 1103 1743 1105 1759
rect 1293 1743 1295 1795
rect 695 1731 727 1743
rect 783 1731 807 1743
rect 863 1731 887 1743
rect 943 1731 967 1743
rect 1023 1731 1047 1743
rect 1103 1731 1127 1743
rect 1183 1731 1207 1743
rect 1263 1731 1295 1743
rect 695 1679 697 1731
rect 885 1703 887 1731
rect 953 1703 967 1731
rect 1023 1703 1037 1731
rect 1103 1703 1105 1731
rect 749 1679 765 1703
rect 817 1679 833 1703
rect 885 1679 901 1703
rect 953 1679 969 1703
rect 1021 1679 1037 1703
rect 1089 1679 1105 1703
rect 1157 1679 1173 1703
rect 1225 1679 1241 1703
rect 1293 1679 1295 1731
rect 695 1678 1295 1679
rect 695 1667 727 1678
rect 783 1667 807 1678
rect 863 1667 887 1678
rect 943 1667 967 1678
rect 1023 1667 1047 1678
rect 1103 1667 1127 1678
rect 1183 1667 1207 1678
rect 1263 1667 1295 1678
rect 695 1615 697 1667
rect 885 1622 887 1667
rect 953 1622 967 1667
rect 1023 1622 1037 1667
rect 1103 1622 1105 1667
rect 749 1615 765 1622
rect 817 1615 833 1622
rect 885 1615 901 1622
rect 953 1615 969 1622
rect 1021 1615 1037 1622
rect 1089 1615 1105 1622
rect 1157 1615 1173 1622
rect 1225 1615 1241 1622
rect 1293 1615 1295 1667
rect 695 1603 1295 1615
rect 695 1551 697 1603
rect 749 1597 765 1603
rect 817 1597 833 1603
rect 885 1597 901 1603
rect 953 1597 969 1603
rect 1021 1597 1037 1603
rect 1089 1597 1105 1603
rect 1157 1597 1173 1603
rect 1225 1597 1241 1603
rect 885 1551 887 1597
rect 953 1551 967 1597
rect 1023 1551 1037 1597
rect 1103 1551 1105 1597
rect 1293 1551 1295 1603
rect 695 1541 727 1551
rect 783 1541 807 1551
rect 863 1541 887 1551
rect 943 1541 967 1551
rect 1023 1541 1047 1551
rect 1103 1541 1127 1551
rect 1183 1541 1207 1551
rect 1263 1541 1295 1551
rect 695 1539 1295 1541
rect 695 1487 697 1539
rect 749 1516 765 1539
rect 817 1516 833 1539
rect 885 1516 901 1539
rect 953 1516 969 1539
rect 1021 1516 1037 1539
rect 1089 1516 1105 1539
rect 1157 1516 1173 1539
rect 1225 1516 1241 1539
rect 885 1487 887 1516
rect 953 1487 967 1516
rect 1023 1487 1037 1516
rect 1103 1487 1105 1516
rect 1293 1487 1295 1539
rect 695 1475 727 1487
rect 783 1475 807 1487
rect 863 1475 887 1487
rect 943 1475 967 1487
rect 1023 1475 1047 1487
rect 1103 1475 1127 1487
rect 1183 1475 1207 1487
rect 1263 1475 1295 1487
rect 695 1423 697 1475
rect 885 1460 887 1475
rect 953 1460 967 1475
rect 1023 1460 1037 1475
rect 1103 1460 1105 1475
rect 749 1435 765 1460
rect 817 1435 833 1460
rect 885 1435 901 1460
rect 953 1435 969 1460
rect 1021 1435 1037 1460
rect 1089 1435 1105 1460
rect 1157 1435 1173 1460
rect 1225 1435 1241 1460
rect 885 1423 887 1435
rect 953 1423 967 1435
rect 1023 1423 1037 1435
rect 1103 1423 1105 1435
rect 1293 1423 1295 1475
rect 695 1411 727 1423
rect 783 1411 807 1423
rect 863 1411 887 1423
rect 943 1411 967 1423
rect 1023 1411 1047 1423
rect 1103 1411 1127 1423
rect 1183 1411 1207 1423
rect 1263 1411 1295 1423
rect 695 1359 697 1411
rect 885 1379 887 1411
rect 953 1379 967 1411
rect 1023 1379 1037 1411
rect 1103 1379 1105 1411
rect 749 1359 765 1379
rect 817 1359 833 1379
rect 885 1359 901 1379
rect 953 1359 969 1379
rect 1021 1359 1037 1379
rect 1089 1359 1105 1379
rect 1157 1359 1173 1379
rect 1225 1359 1241 1379
rect 1293 1359 1295 1411
rect 695 1354 1295 1359
rect 695 1347 727 1354
rect 783 1347 807 1354
rect 863 1347 887 1354
rect 943 1347 967 1354
rect 1023 1347 1047 1354
rect 1103 1347 1127 1354
rect 1183 1347 1207 1354
rect 1263 1347 1295 1354
rect 695 1295 697 1347
rect 885 1298 887 1347
rect 953 1298 967 1347
rect 1023 1298 1037 1347
rect 1103 1298 1105 1347
rect 749 1295 765 1298
rect 817 1295 833 1298
rect 885 1295 901 1298
rect 953 1295 969 1298
rect 1021 1295 1037 1298
rect 1089 1295 1105 1298
rect 1157 1295 1173 1298
rect 1225 1295 1241 1298
rect 1293 1295 1295 1347
rect 695 141 1295 1295
rect 695 85 704 141
rect 760 85 792 141
rect 848 85 880 141
rect 936 85 968 141
rect 1024 85 1056 141
rect 1112 85 1143 141
rect 1199 85 1230 141
rect 1286 85 1295 141
rect 695 61 1295 85
rect 695 5 704 61
rect 760 5 792 61
rect 848 5 880 61
rect 936 5 968 61
rect 1024 5 1056 61
rect 1112 5 1143 61
rect 1199 5 1230 61
rect 1286 5 1295 61
rect 695 0 1295 5
rect 1495 39011 1501 39063
rect 1553 39011 1569 39063
rect 1621 39011 1636 39063
rect 1688 39011 1703 39063
rect 1755 39011 1770 39063
rect 1822 39011 1837 39063
rect 1889 39011 1895 39063
rect 1495 36933 1895 39011
rect 1495 36881 1501 36933
rect 1553 36881 1569 36933
rect 1621 36881 1636 36933
rect 1688 36881 1703 36933
rect 1755 36881 1770 36933
rect 1822 36881 1837 36933
rect 1889 36881 1895 36933
rect 1495 34803 1895 36881
rect 1495 34751 1501 34803
rect 1553 34751 1569 34803
rect 1621 34751 1636 34803
rect 1688 34751 1703 34803
rect 1755 34751 1770 34803
rect 1822 34751 1837 34803
rect 1889 34751 1895 34803
rect 1495 32673 1895 34751
rect 1495 32621 1501 32673
rect 1553 32621 1569 32673
rect 1621 32621 1636 32673
rect 1688 32621 1703 32673
rect 1755 32621 1770 32673
rect 1822 32621 1837 32673
rect 1889 32621 1895 32673
rect 1495 30543 1895 32621
rect 1495 30491 1501 30543
rect 1553 30491 1569 30543
rect 1621 30491 1636 30543
rect 1688 30491 1703 30543
rect 1755 30491 1770 30543
rect 1822 30491 1837 30543
rect 1889 30491 1895 30543
rect 1495 28413 1895 30491
rect 1495 28361 1501 28413
rect 1553 28361 1569 28413
rect 1621 28361 1636 28413
rect 1688 28361 1703 28413
rect 1755 28361 1770 28413
rect 1822 28361 1837 28413
rect 1889 28361 1895 28413
rect 1495 26283 1895 28361
rect 1495 26231 1501 26283
rect 1553 26231 1569 26283
rect 1621 26231 1636 26283
rect 1688 26231 1703 26283
rect 1755 26231 1770 26283
rect 1822 26231 1837 26283
rect 1889 26231 1895 26283
rect 1495 24153 1895 26231
rect 1495 24101 1501 24153
rect 1553 24101 1569 24153
rect 1621 24101 1636 24153
rect 1688 24101 1703 24153
rect 1755 24101 1770 24153
rect 1822 24101 1837 24153
rect 1889 24101 1895 24153
rect 1495 22023 1895 24101
rect 1495 21971 1501 22023
rect 1553 21971 1569 22023
rect 1621 21971 1636 22023
rect 1688 21971 1703 22023
rect 1755 21971 1770 22023
rect 1822 21971 1837 22023
rect 1889 21971 1895 22023
rect 1495 19893 1895 21971
rect 1495 19841 1501 19893
rect 1553 19841 1569 19893
rect 1621 19841 1636 19893
rect 1688 19841 1703 19893
rect 1755 19841 1770 19893
rect 1822 19841 1837 19893
rect 1889 19841 1895 19893
rect 1495 17763 1895 19841
rect 1495 17711 1501 17763
rect 1553 17711 1569 17763
rect 1621 17711 1636 17763
rect 1688 17711 1703 17763
rect 1755 17711 1770 17763
rect 1822 17711 1837 17763
rect 1889 17711 1895 17763
rect 1495 15633 1895 17711
rect 1495 15581 1501 15633
rect 1553 15581 1569 15633
rect 1621 15581 1636 15633
rect 1688 15581 1703 15633
rect 1755 15581 1770 15633
rect 1822 15581 1837 15633
rect 1889 15581 1895 15633
rect 1495 13503 1895 15581
rect 1495 13451 1501 13503
rect 1553 13451 1569 13503
rect 1621 13451 1636 13503
rect 1688 13451 1703 13503
rect 1755 13451 1770 13503
rect 1822 13451 1837 13503
rect 1889 13451 1895 13503
rect 1495 11373 1895 13451
rect 1495 11321 1501 11373
rect 1553 11321 1569 11373
rect 1621 11321 1636 11373
rect 1688 11321 1703 11373
rect 1755 11321 1770 11373
rect 1822 11321 1837 11373
rect 1889 11321 1895 11373
rect 1495 9243 1895 11321
rect 1495 9191 1501 9243
rect 1553 9191 1569 9243
rect 1621 9191 1636 9243
rect 1688 9191 1703 9243
rect 1755 9191 1770 9243
rect 1822 9191 1837 9243
rect 1889 9191 1895 9243
rect 1495 7113 1895 9191
rect 1495 7061 1501 7113
rect 1553 7061 1569 7113
rect 1621 7061 1636 7113
rect 1688 7061 1703 7113
rect 1755 7061 1770 7113
rect 1822 7061 1837 7113
rect 1889 7061 1895 7113
rect 1495 4983 1895 7061
rect 1495 4931 1501 4983
rect 1553 4931 1569 4983
rect 1621 4931 1636 4983
rect 1688 4931 1703 4983
rect 1755 4931 1770 4983
rect 1822 4931 1837 4983
rect 1889 4931 1895 4983
rect 1495 2853 1895 4931
rect 1495 2801 1501 2853
rect 1553 2801 1569 2853
rect 1621 2801 1636 2853
rect 1688 2801 1703 2853
rect 1755 2801 1770 2853
rect 1822 2801 1837 2853
rect 1889 2801 1895 2853
rect 1495 723 1895 2801
rect 1495 671 1501 723
rect 1553 671 1569 723
rect 1621 671 1636 723
rect 1688 671 1703 723
rect 1755 671 1770 723
rect 1822 671 1837 723
rect 1889 671 1895 723
rect 1495 141 1895 671
rect 1495 85 1504 141
rect 1560 85 1585 141
rect 1641 85 1666 141
rect 1722 85 1747 141
rect 1495 61 1747 85
rect 1495 5 1504 61
rect 1560 5 1585 61
rect 1641 5 1666 61
rect 1722 5 1747 61
rect 1883 5 1895 141
rect 1495 0 1895 5
rect 2095 38423 2695 39341
rect 2095 38371 2097 38423
rect 2149 38420 2165 38423
rect 2217 38420 2233 38423
rect 2285 38420 2301 38423
rect 2353 38420 2369 38423
rect 2421 38420 2437 38423
rect 2489 38420 2505 38423
rect 2557 38420 2573 38423
rect 2625 38420 2641 38423
rect 2693 38371 2695 38423
rect 2095 38359 2127 38371
rect 2663 38359 2695 38371
rect 2095 38307 2097 38359
rect 2693 38307 2695 38359
rect 2095 38295 2127 38307
rect 2663 38295 2695 38307
rect 2095 38243 2097 38295
rect 2693 38243 2695 38295
rect 2095 38231 2127 38243
rect 2663 38231 2695 38243
rect 2095 38179 2097 38231
rect 2693 38179 2695 38231
rect 2095 38167 2127 38179
rect 2663 38167 2695 38179
rect 2095 38115 2097 38167
rect 2693 38115 2695 38167
rect 2095 38103 2127 38115
rect 2663 38103 2695 38115
rect 2095 38051 2097 38103
rect 2693 38051 2695 38103
rect 2095 38039 2127 38051
rect 2663 38039 2695 38051
rect 2095 37987 2097 38039
rect 2693 37987 2695 38039
rect 2095 37975 2127 37987
rect 2663 37975 2695 37987
rect 2095 37923 2097 37975
rect 2149 37939 2165 37964
rect 2217 37939 2233 37964
rect 2285 37939 2301 37964
rect 2353 37939 2369 37964
rect 2421 37939 2437 37964
rect 2489 37939 2505 37964
rect 2557 37939 2573 37964
rect 2625 37939 2641 37964
rect 2285 37923 2287 37939
rect 2353 37923 2367 37939
rect 2423 37923 2437 37939
rect 2503 37923 2505 37939
rect 2693 37923 2695 37975
rect 2095 37911 2127 37923
rect 2183 37911 2207 37923
rect 2263 37911 2287 37923
rect 2343 37911 2367 37923
rect 2423 37911 2447 37923
rect 2503 37911 2527 37923
rect 2583 37911 2607 37923
rect 2663 37911 2695 37923
rect 2095 37859 2097 37911
rect 2285 37883 2287 37911
rect 2353 37883 2367 37911
rect 2423 37883 2437 37911
rect 2503 37883 2505 37911
rect 2149 37859 2165 37883
rect 2217 37859 2233 37883
rect 2285 37859 2301 37883
rect 2353 37859 2369 37883
rect 2421 37859 2437 37883
rect 2489 37859 2505 37883
rect 2557 37859 2573 37883
rect 2625 37859 2641 37883
rect 2693 37859 2695 37911
rect 2095 37858 2695 37859
rect 2095 37847 2127 37858
rect 2183 37847 2207 37858
rect 2263 37847 2287 37858
rect 2343 37847 2367 37858
rect 2423 37847 2447 37858
rect 2503 37847 2527 37858
rect 2583 37847 2607 37858
rect 2663 37847 2695 37858
rect 2095 37795 2097 37847
rect 2285 37802 2287 37847
rect 2353 37802 2367 37847
rect 2423 37802 2437 37847
rect 2503 37802 2505 37847
rect 2149 37795 2165 37802
rect 2217 37795 2233 37802
rect 2285 37795 2301 37802
rect 2353 37795 2369 37802
rect 2421 37795 2437 37802
rect 2489 37795 2505 37802
rect 2557 37795 2573 37802
rect 2625 37795 2641 37802
rect 2693 37795 2695 37847
rect 2095 37783 2695 37795
rect 2095 37731 2097 37783
rect 2149 37777 2165 37783
rect 2217 37777 2233 37783
rect 2285 37777 2301 37783
rect 2353 37777 2369 37783
rect 2421 37777 2437 37783
rect 2489 37777 2505 37783
rect 2557 37777 2573 37783
rect 2625 37777 2641 37783
rect 2285 37731 2287 37777
rect 2353 37731 2367 37777
rect 2423 37731 2437 37777
rect 2503 37731 2505 37777
rect 2693 37731 2695 37783
rect 2095 37721 2127 37731
rect 2183 37721 2207 37731
rect 2263 37721 2287 37731
rect 2343 37721 2367 37731
rect 2423 37721 2447 37731
rect 2503 37721 2527 37731
rect 2583 37721 2607 37731
rect 2663 37721 2695 37731
rect 2095 37719 2695 37721
rect 2095 37667 2097 37719
rect 2149 37696 2165 37719
rect 2217 37696 2233 37719
rect 2285 37696 2301 37719
rect 2353 37696 2369 37719
rect 2421 37696 2437 37719
rect 2489 37696 2505 37719
rect 2557 37696 2573 37719
rect 2625 37696 2641 37719
rect 2285 37667 2287 37696
rect 2353 37667 2367 37696
rect 2423 37667 2437 37696
rect 2503 37667 2505 37696
rect 2693 37667 2695 37719
rect 2095 37655 2127 37667
rect 2183 37655 2207 37667
rect 2263 37655 2287 37667
rect 2343 37655 2367 37667
rect 2423 37655 2447 37667
rect 2503 37655 2527 37667
rect 2583 37655 2607 37667
rect 2663 37655 2695 37667
rect 2095 37603 2097 37655
rect 2285 37640 2287 37655
rect 2353 37640 2367 37655
rect 2423 37640 2437 37655
rect 2503 37640 2505 37655
rect 2149 37615 2165 37640
rect 2217 37615 2233 37640
rect 2285 37615 2301 37640
rect 2353 37615 2369 37640
rect 2421 37615 2437 37640
rect 2489 37615 2505 37640
rect 2557 37615 2573 37640
rect 2625 37615 2641 37640
rect 2285 37603 2287 37615
rect 2353 37603 2367 37615
rect 2423 37603 2437 37615
rect 2503 37603 2505 37615
rect 2693 37603 2695 37655
rect 2095 37591 2127 37603
rect 2183 37591 2207 37603
rect 2263 37591 2287 37603
rect 2343 37591 2367 37603
rect 2423 37591 2447 37603
rect 2503 37591 2527 37603
rect 2583 37591 2607 37603
rect 2663 37591 2695 37603
rect 2095 37539 2097 37591
rect 2285 37559 2287 37591
rect 2353 37559 2367 37591
rect 2423 37559 2437 37591
rect 2503 37559 2505 37591
rect 2149 37539 2165 37559
rect 2217 37539 2233 37559
rect 2285 37539 2301 37559
rect 2353 37539 2369 37559
rect 2421 37539 2437 37559
rect 2489 37539 2505 37559
rect 2557 37539 2573 37559
rect 2625 37539 2641 37559
rect 2693 37539 2695 37591
rect 2095 37534 2695 37539
rect 2095 37527 2127 37534
rect 2183 37527 2207 37534
rect 2263 37527 2287 37534
rect 2343 37527 2367 37534
rect 2423 37527 2447 37534
rect 2503 37527 2527 37534
rect 2583 37527 2607 37534
rect 2663 37527 2695 37534
rect 2095 37475 2097 37527
rect 2285 37478 2287 37527
rect 2353 37478 2367 37527
rect 2423 37478 2437 37527
rect 2503 37478 2505 37527
rect 2149 37475 2165 37478
rect 2217 37475 2233 37478
rect 2285 37475 2301 37478
rect 2353 37475 2369 37478
rect 2421 37475 2437 37478
rect 2489 37475 2505 37478
rect 2557 37475 2573 37478
rect 2625 37475 2641 37478
rect 2693 37475 2695 37527
rect 2095 36369 2695 37475
rect 2095 36317 2097 36369
rect 2149 36366 2165 36369
rect 2217 36366 2233 36369
rect 2285 36366 2301 36369
rect 2353 36366 2369 36369
rect 2421 36366 2437 36369
rect 2489 36366 2505 36369
rect 2557 36366 2573 36369
rect 2625 36366 2641 36369
rect 2693 36317 2695 36369
rect 2095 36305 2127 36317
rect 2663 36305 2695 36317
rect 2095 36253 2097 36305
rect 2693 36253 2695 36305
rect 2095 36241 2127 36253
rect 2663 36241 2695 36253
rect 2095 36189 2097 36241
rect 2693 36189 2695 36241
rect 2095 36177 2127 36189
rect 2663 36177 2695 36189
rect 2095 36125 2097 36177
rect 2693 36125 2695 36177
rect 2095 36113 2127 36125
rect 2663 36113 2695 36125
rect 2095 36061 2097 36113
rect 2693 36061 2695 36113
rect 2095 36049 2127 36061
rect 2663 36049 2695 36061
rect 2095 35997 2097 36049
rect 2693 35997 2695 36049
rect 2095 35985 2127 35997
rect 2663 35985 2695 35997
rect 2095 35933 2097 35985
rect 2693 35933 2695 35985
rect 2095 35921 2127 35933
rect 2663 35921 2695 35933
rect 2095 35869 2097 35921
rect 2149 35885 2165 35910
rect 2217 35885 2233 35910
rect 2285 35885 2301 35910
rect 2353 35885 2369 35910
rect 2421 35885 2437 35910
rect 2489 35885 2505 35910
rect 2557 35885 2573 35910
rect 2625 35885 2641 35910
rect 2285 35869 2287 35885
rect 2353 35869 2367 35885
rect 2423 35869 2437 35885
rect 2503 35869 2505 35885
rect 2693 35869 2695 35921
rect 2095 35857 2127 35869
rect 2183 35857 2207 35869
rect 2263 35857 2287 35869
rect 2343 35857 2367 35869
rect 2423 35857 2447 35869
rect 2503 35857 2527 35869
rect 2583 35857 2607 35869
rect 2663 35857 2695 35869
rect 2095 35805 2097 35857
rect 2285 35829 2287 35857
rect 2353 35829 2367 35857
rect 2423 35829 2437 35857
rect 2503 35829 2505 35857
rect 2149 35805 2165 35829
rect 2217 35805 2233 35829
rect 2285 35805 2301 35829
rect 2353 35805 2369 35829
rect 2421 35805 2437 35829
rect 2489 35805 2505 35829
rect 2557 35805 2573 35829
rect 2625 35805 2641 35829
rect 2693 35805 2695 35857
rect 2095 35804 2695 35805
rect 2095 35793 2127 35804
rect 2183 35793 2207 35804
rect 2263 35793 2287 35804
rect 2343 35793 2367 35804
rect 2423 35793 2447 35804
rect 2503 35793 2527 35804
rect 2583 35793 2607 35804
rect 2663 35793 2695 35804
rect 2095 35741 2097 35793
rect 2285 35748 2287 35793
rect 2353 35748 2367 35793
rect 2423 35748 2437 35793
rect 2503 35748 2505 35793
rect 2149 35741 2165 35748
rect 2217 35741 2233 35748
rect 2285 35741 2301 35748
rect 2353 35741 2369 35748
rect 2421 35741 2437 35748
rect 2489 35741 2505 35748
rect 2557 35741 2573 35748
rect 2625 35741 2641 35748
rect 2693 35741 2695 35793
rect 2095 35729 2695 35741
rect 2095 35677 2097 35729
rect 2149 35723 2165 35729
rect 2217 35723 2233 35729
rect 2285 35723 2301 35729
rect 2353 35723 2369 35729
rect 2421 35723 2437 35729
rect 2489 35723 2505 35729
rect 2557 35723 2573 35729
rect 2625 35723 2641 35729
rect 2285 35677 2287 35723
rect 2353 35677 2367 35723
rect 2423 35677 2437 35723
rect 2503 35677 2505 35723
rect 2693 35677 2695 35729
rect 2095 35667 2127 35677
rect 2183 35667 2207 35677
rect 2263 35667 2287 35677
rect 2343 35667 2367 35677
rect 2423 35667 2447 35677
rect 2503 35667 2527 35677
rect 2583 35667 2607 35677
rect 2663 35667 2695 35677
rect 2095 35665 2695 35667
rect 2095 35613 2097 35665
rect 2149 35642 2165 35665
rect 2217 35642 2233 35665
rect 2285 35642 2301 35665
rect 2353 35642 2369 35665
rect 2421 35642 2437 35665
rect 2489 35642 2505 35665
rect 2557 35642 2573 35665
rect 2625 35642 2641 35665
rect 2285 35613 2287 35642
rect 2353 35613 2367 35642
rect 2423 35613 2437 35642
rect 2503 35613 2505 35642
rect 2693 35613 2695 35665
rect 2095 35601 2127 35613
rect 2183 35601 2207 35613
rect 2263 35601 2287 35613
rect 2343 35601 2367 35613
rect 2423 35601 2447 35613
rect 2503 35601 2527 35613
rect 2583 35601 2607 35613
rect 2663 35601 2695 35613
rect 2095 35549 2097 35601
rect 2285 35586 2287 35601
rect 2353 35586 2367 35601
rect 2423 35586 2437 35601
rect 2503 35586 2505 35601
rect 2149 35561 2165 35586
rect 2217 35561 2233 35586
rect 2285 35561 2301 35586
rect 2353 35561 2369 35586
rect 2421 35561 2437 35586
rect 2489 35561 2505 35586
rect 2557 35561 2573 35586
rect 2625 35561 2641 35586
rect 2285 35549 2287 35561
rect 2353 35549 2367 35561
rect 2423 35549 2437 35561
rect 2503 35549 2505 35561
rect 2693 35549 2695 35601
rect 2095 35537 2127 35549
rect 2183 35537 2207 35549
rect 2263 35537 2287 35549
rect 2343 35537 2367 35549
rect 2423 35537 2447 35549
rect 2503 35537 2527 35549
rect 2583 35537 2607 35549
rect 2663 35537 2695 35549
rect 2095 35485 2097 35537
rect 2285 35505 2287 35537
rect 2353 35505 2367 35537
rect 2423 35505 2437 35537
rect 2503 35505 2505 35537
rect 2149 35485 2165 35505
rect 2217 35485 2233 35505
rect 2285 35485 2301 35505
rect 2353 35485 2369 35505
rect 2421 35485 2437 35505
rect 2489 35485 2505 35505
rect 2557 35485 2573 35505
rect 2625 35485 2641 35505
rect 2693 35485 2695 35537
rect 2095 35480 2695 35485
rect 2095 35473 2127 35480
rect 2183 35473 2207 35480
rect 2263 35473 2287 35480
rect 2343 35473 2367 35480
rect 2423 35473 2447 35480
rect 2503 35473 2527 35480
rect 2583 35473 2607 35480
rect 2663 35473 2695 35480
rect 2095 35421 2097 35473
rect 2285 35424 2287 35473
rect 2353 35424 2367 35473
rect 2423 35424 2437 35473
rect 2503 35424 2505 35473
rect 2149 35421 2165 35424
rect 2217 35421 2233 35424
rect 2285 35421 2301 35424
rect 2353 35421 2369 35424
rect 2421 35421 2437 35424
rect 2489 35421 2505 35424
rect 2557 35421 2573 35424
rect 2625 35421 2641 35424
rect 2693 35421 2695 35473
rect 2095 34150 2695 35421
rect 2095 34098 2097 34150
rect 2149 34147 2165 34150
rect 2217 34147 2233 34150
rect 2285 34147 2301 34150
rect 2353 34147 2369 34150
rect 2421 34147 2437 34150
rect 2489 34147 2505 34150
rect 2557 34147 2573 34150
rect 2625 34147 2641 34150
rect 2693 34098 2695 34150
rect 2095 34086 2127 34098
rect 2663 34086 2695 34098
rect 2095 34034 2097 34086
rect 2693 34034 2695 34086
rect 2095 34022 2127 34034
rect 2663 34022 2695 34034
rect 2095 33970 2097 34022
rect 2693 33970 2695 34022
rect 2095 33958 2127 33970
rect 2663 33958 2695 33970
rect 2095 33906 2097 33958
rect 2693 33906 2695 33958
rect 2095 33894 2127 33906
rect 2663 33894 2695 33906
rect 2095 33842 2097 33894
rect 2693 33842 2695 33894
rect 2095 33830 2127 33842
rect 2663 33830 2695 33842
rect 2095 33778 2097 33830
rect 2693 33778 2695 33830
rect 2095 33766 2127 33778
rect 2663 33766 2695 33778
rect 2095 33714 2097 33766
rect 2693 33714 2695 33766
rect 2095 33702 2127 33714
rect 2663 33702 2695 33714
rect 2095 33650 2097 33702
rect 2149 33666 2165 33691
rect 2217 33666 2233 33691
rect 2285 33666 2301 33691
rect 2353 33666 2369 33691
rect 2421 33666 2437 33691
rect 2489 33666 2505 33691
rect 2557 33666 2573 33691
rect 2625 33666 2641 33691
rect 2285 33650 2287 33666
rect 2353 33650 2367 33666
rect 2423 33650 2437 33666
rect 2503 33650 2505 33666
rect 2693 33650 2695 33702
rect 2095 33638 2127 33650
rect 2183 33638 2207 33650
rect 2263 33638 2287 33650
rect 2343 33638 2367 33650
rect 2423 33638 2447 33650
rect 2503 33638 2527 33650
rect 2583 33638 2607 33650
rect 2663 33638 2695 33650
rect 2095 33586 2097 33638
rect 2285 33610 2287 33638
rect 2353 33610 2367 33638
rect 2423 33610 2437 33638
rect 2503 33610 2505 33638
rect 2149 33586 2165 33610
rect 2217 33586 2233 33610
rect 2285 33586 2301 33610
rect 2353 33586 2369 33610
rect 2421 33586 2437 33610
rect 2489 33586 2505 33610
rect 2557 33586 2573 33610
rect 2625 33586 2641 33610
rect 2693 33586 2695 33638
rect 2095 33585 2695 33586
rect 2095 33574 2127 33585
rect 2183 33574 2207 33585
rect 2263 33574 2287 33585
rect 2343 33574 2367 33585
rect 2423 33574 2447 33585
rect 2503 33574 2527 33585
rect 2583 33574 2607 33585
rect 2663 33574 2695 33585
rect 2095 33522 2097 33574
rect 2285 33529 2287 33574
rect 2353 33529 2367 33574
rect 2423 33529 2437 33574
rect 2503 33529 2505 33574
rect 2149 33522 2165 33529
rect 2217 33522 2233 33529
rect 2285 33522 2301 33529
rect 2353 33522 2369 33529
rect 2421 33522 2437 33529
rect 2489 33522 2505 33529
rect 2557 33522 2573 33529
rect 2625 33522 2641 33529
rect 2693 33522 2695 33574
rect 2095 33510 2695 33522
rect 2095 33458 2097 33510
rect 2149 33504 2165 33510
rect 2217 33504 2233 33510
rect 2285 33504 2301 33510
rect 2353 33504 2369 33510
rect 2421 33504 2437 33510
rect 2489 33504 2505 33510
rect 2557 33504 2573 33510
rect 2625 33504 2641 33510
rect 2285 33458 2287 33504
rect 2353 33458 2367 33504
rect 2423 33458 2437 33504
rect 2503 33458 2505 33504
rect 2693 33458 2695 33510
rect 2095 33448 2127 33458
rect 2183 33448 2207 33458
rect 2263 33448 2287 33458
rect 2343 33448 2367 33458
rect 2423 33448 2447 33458
rect 2503 33448 2527 33458
rect 2583 33448 2607 33458
rect 2663 33448 2695 33458
rect 2095 33446 2695 33448
rect 2095 33394 2097 33446
rect 2149 33423 2165 33446
rect 2217 33423 2233 33446
rect 2285 33423 2301 33446
rect 2353 33423 2369 33446
rect 2421 33423 2437 33446
rect 2489 33423 2505 33446
rect 2557 33423 2573 33446
rect 2625 33423 2641 33446
rect 2285 33394 2287 33423
rect 2353 33394 2367 33423
rect 2423 33394 2437 33423
rect 2503 33394 2505 33423
rect 2693 33394 2695 33446
rect 2095 33382 2127 33394
rect 2183 33382 2207 33394
rect 2263 33382 2287 33394
rect 2343 33382 2367 33394
rect 2423 33382 2447 33394
rect 2503 33382 2527 33394
rect 2583 33382 2607 33394
rect 2663 33382 2695 33394
rect 2095 33330 2097 33382
rect 2285 33367 2287 33382
rect 2353 33367 2367 33382
rect 2423 33367 2437 33382
rect 2503 33367 2505 33382
rect 2149 33342 2165 33367
rect 2217 33342 2233 33367
rect 2285 33342 2301 33367
rect 2353 33342 2369 33367
rect 2421 33342 2437 33367
rect 2489 33342 2505 33367
rect 2557 33342 2573 33367
rect 2625 33342 2641 33367
rect 2285 33330 2287 33342
rect 2353 33330 2367 33342
rect 2423 33330 2437 33342
rect 2503 33330 2505 33342
rect 2693 33330 2695 33382
rect 2095 33318 2127 33330
rect 2183 33318 2207 33330
rect 2263 33318 2287 33330
rect 2343 33318 2367 33330
rect 2423 33318 2447 33330
rect 2503 33318 2527 33330
rect 2583 33318 2607 33330
rect 2663 33318 2695 33330
rect 2095 33266 2097 33318
rect 2285 33286 2287 33318
rect 2353 33286 2367 33318
rect 2423 33286 2437 33318
rect 2503 33286 2505 33318
rect 2149 33266 2165 33286
rect 2217 33266 2233 33286
rect 2285 33266 2301 33286
rect 2353 33266 2369 33286
rect 2421 33266 2437 33286
rect 2489 33266 2505 33286
rect 2557 33266 2573 33286
rect 2625 33266 2641 33286
rect 2693 33266 2695 33318
rect 2095 33261 2695 33266
rect 2095 33254 2127 33261
rect 2183 33254 2207 33261
rect 2263 33254 2287 33261
rect 2343 33254 2367 33261
rect 2423 33254 2447 33261
rect 2503 33254 2527 33261
rect 2583 33254 2607 33261
rect 2663 33254 2695 33261
rect 2095 33202 2097 33254
rect 2285 33205 2287 33254
rect 2353 33205 2367 33254
rect 2423 33205 2437 33254
rect 2503 33205 2505 33254
rect 2149 33202 2165 33205
rect 2217 33202 2233 33205
rect 2285 33202 2301 33205
rect 2353 33202 2369 33205
rect 2421 33202 2437 33205
rect 2489 33202 2505 33205
rect 2557 33202 2573 33205
rect 2625 33202 2641 33205
rect 2693 33202 2695 33254
rect 2095 32021 2695 33202
rect 2095 31969 2097 32021
rect 2149 32018 2165 32021
rect 2217 32018 2233 32021
rect 2285 32018 2301 32021
rect 2353 32018 2369 32021
rect 2421 32018 2437 32021
rect 2489 32018 2505 32021
rect 2557 32018 2573 32021
rect 2625 32018 2641 32021
rect 2693 31969 2695 32021
rect 2095 31957 2127 31969
rect 2663 31957 2695 31969
rect 2095 31905 2097 31957
rect 2693 31905 2695 31957
rect 2095 31893 2127 31905
rect 2663 31893 2695 31905
rect 2095 31841 2097 31893
rect 2693 31841 2695 31893
rect 2095 31829 2127 31841
rect 2663 31829 2695 31841
rect 2095 31777 2097 31829
rect 2693 31777 2695 31829
rect 2095 31765 2127 31777
rect 2663 31765 2695 31777
rect 2095 31713 2097 31765
rect 2693 31713 2695 31765
rect 2095 31701 2127 31713
rect 2663 31701 2695 31713
rect 2095 31649 2097 31701
rect 2693 31649 2695 31701
rect 2095 31637 2127 31649
rect 2663 31637 2695 31649
rect 2095 31585 2097 31637
rect 2693 31585 2695 31637
rect 2095 31573 2127 31585
rect 2663 31573 2695 31585
rect 2095 31521 2097 31573
rect 2149 31537 2165 31562
rect 2217 31537 2233 31562
rect 2285 31537 2301 31562
rect 2353 31537 2369 31562
rect 2421 31537 2437 31562
rect 2489 31537 2505 31562
rect 2557 31537 2573 31562
rect 2625 31537 2641 31562
rect 2285 31521 2287 31537
rect 2353 31521 2367 31537
rect 2423 31521 2437 31537
rect 2503 31521 2505 31537
rect 2693 31521 2695 31573
rect 2095 31509 2127 31521
rect 2183 31509 2207 31521
rect 2263 31509 2287 31521
rect 2343 31509 2367 31521
rect 2423 31509 2447 31521
rect 2503 31509 2527 31521
rect 2583 31509 2607 31521
rect 2663 31509 2695 31521
rect 2095 31457 2097 31509
rect 2285 31481 2287 31509
rect 2353 31481 2367 31509
rect 2423 31481 2437 31509
rect 2503 31481 2505 31509
rect 2149 31457 2165 31481
rect 2217 31457 2233 31481
rect 2285 31457 2301 31481
rect 2353 31457 2369 31481
rect 2421 31457 2437 31481
rect 2489 31457 2505 31481
rect 2557 31457 2573 31481
rect 2625 31457 2641 31481
rect 2693 31457 2695 31509
rect 2095 31456 2695 31457
rect 2095 31445 2127 31456
rect 2183 31445 2207 31456
rect 2263 31445 2287 31456
rect 2343 31445 2367 31456
rect 2423 31445 2447 31456
rect 2503 31445 2527 31456
rect 2583 31445 2607 31456
rect 2663 31445 2695 31456
rect 2095 31393 2097 31445
rect 2285 31400 2287 31445
rect 2353 31400 2367 31445
rect 2423 31400 2437 31445
rect 2503 31400 2505 31445
rect 2149 31393 2165 31400
rect 2217 31393 2233 31400
rect 2285 31393 2301 31400
rect 2353 31393 2369 31400
rect 2421 31393 2437 31400
rect 2489 31393 2505 31400
rect 2557 31393 2573 31400
rect 2625 31393 2641 31400
rect 2693 31393 2695 31445
rect 2095 31381 2695 31393
rect 2095 31329 2097 31381
rect 2149 31375 2165 31381
rect 2217 31375 2233 31381
rect 2285 31375 2301 31381
rect 2353 31375 2369 31381
rect 2421 31375 2437 31381
rect 2489 31375 2505 31381
rect 2557 31375 2573 31381
rect 2625 31375 2641 31381
rect 2285 31329 2287 31375
rect 2353 31329 2367 31375
rect 2423 31329 2437 31375
rect 2503 31329 2505 31375
rect 2693 31329 2695 31381
rect 2095 31319 2127 31329
rect 2183 31319 2207 31329
rect 2263 31319 2287 31329
rect 2343 31319 2367 31329
rect 2423 31319 2447 31329
rect 2503 31319 2527 31329
rect 2583 31319 2607 31329
rect 2663 31319 2695 31329
rect 2095 31317 2695 31319
rect 2095 31265 2097 31317
rect 2149 31294 2165 31317
rect 2217 31294 2233 31317
rect 2285 31294 2301 31317
rect 2353 31294 2369 31317
rect 2421 31294 2437 31317
rect 2489 31294 2505 31317
rect 2557 31294 2573 31317
rect 2625 31294 2641 31317
rect 2285 31265 2287 31294
rect 2353 31265 2367 31294
rect 2423 31265 2437 31294
rect 2503 31265 2505 31294
rect 2693 31265 2695 31317
rect 2095 31253 2127 31265
rect 2183 31253 2207 31265
rect 2263 31253 2287 31265
rect 2343 31253 2367 31265
rect 2423 31253 2447 31265
rect 2503 31253 2527 31265
rect 2583 31253 2607 31265
rect 2663 31253 2695 31265
rect 2095 31201 2097 31253
rect 2285 31238 2287 31253
rect 2353 31238 2367 31253
rect 2423 31238 2437 31253
rect 2503 31238 2505 31253
rect 2149 31213 2165 31238
rect 2217 31213 2233 31238
rect 2285 31213 2301 31238
rect 2353 31213 2369 31238
rect 2421 31213 2437 31238
rect 2489 31213 2505 31238
rect 2557 31213 2573 31238
rect 2625 31213 2641 31238
rect 2285 31201 2287 31213
rect 2353 31201 2367 31213
rect 2423 31201 2437 31213
rect 2503 31201 2505 31213
rect 2693 31201 2695 31253
rect 2095 31189 2127 31201
rect 2183 31189 2207 31201
rect 2263 31189 2287 31201
rect 2343 31189 2367 31201
rect 2423 31189 2447 31201
rect 2503 31189 2527 31201
rect 2583 31189 2607 31201
rect 2663 31189 2695 31201
rect 2095 31137 2097 31189
rect 2285 31157 2287 31189
rect 2353 31157 2367 31189
rect 2423 31157 2437 31189
rect 2503 31157 2505 31189
rect 2149 31137 2165 31157
rect 2217 31137 2233 31157
rect 2285 31137 2301 31157
rect 2353 31137 2369 31157
rect 2421 31137 2437 31157
rect 2489 31137 2505 31157
rect 2557 31137 2573 31157
rect 2625 31137 2641 31157
rect 2693 31137 2695 31189
rect 2095 31132 2695 31137
rect 2095 31125 2127 31132
rect 2183 31125 2207 31132
rect 2263 31125 2287 31132
rect 2343 31125 2367 31132
rect 2423 31125 2447 31132
rect 2503 31125 2527 31132
rect 2583 31125 2607 31132
rect 2663 31125 2695 31132
rect 2095 31073 2097 31125
rect 2285 31076 2287 31125
rect 2353 31076 2367 31125
rect 2423 31076 2437 31125
rect 2503 31076 2505 31125
rect 2149 31073 2165 31076
rect 2217 31073 2233 31076
rect 2285 31073 2301 31076
rect 2353 31073 2369 31076
rect 2421 31073 2437 31076
rect 2489 31073 2505 31076
rect 2557 31073 2573 31076
rect 2625 31073 2641 31076
rect 2693 31073 2695 31125
rect 2095 29872 2695 31073
rect 2095 29820 2097 29872
rect 2149 29869 2165 29872
rect 2217 29869 2233 29872
rect 2285 29869 2301 29872
rect 2353 29869 2369 29872
rect 2421 29869 2437 29872
rect 2489 29869 2505 29872
rect 2557 29869 2573 29872
rect 2625 29869 2641 29872
rect 2693 29820 2695 29872
rect 2095 29808 2127 29820
rect 2663 29808 2695 29820
rect 2095 29756 2097 29808
rect 2693 29756 2695 29808
rect 2095 29744 2127 29756
rect 2663 29744 2695 29756
rect 2095 29692 2097 29744
rect 2693 29692 2695 29744
rect 2095 29680 2127 29692
rect 2663 29680 2695 29692
rect 2095 29628 2097 29680
rect 2693 29628 2695 29680
rect 2095 29616 2127 29628
rect 2663 29616 2695 29628
rect 2095 29564 2097 29616
rect 2693 29564 2695 29616
rect 2095 29552 2127 29564
rect 2663 29552 2695 29564
rect 2095 29500 2097 29552
rect 2693 29500 2695 29552
rect 2095 29488 2127 29500
rect 2663 29488 2695 29500
rect 2095 29436 2097 29488
rect 2693 29436 2695 29488
rect 2095 29424 2127 29436
rect 2663 29424 2695 29436
rect 2095 29372 2097 29424
rect 2149 29388 2165 29413
rect 2217 29388 2233 29413
rect 2285 29388 2301 29413
rect 2353 29388 2369 29413
rect 2421 29388 2437 29413
rect 2489 29388 2505 29413
rect 2557 29388 2573 29413
rect 2625 29388 2641 29413
rect 2285 29372 2287 29388
rect 2353 29372 2367 29388
rect 2423 29372 2437 29388
rect 2503 29372 2505 29388
rect 2693 29372 2695 29424
rect 2095 29360 2127 29372
rect 2183 29360 2207 29372
rect 2263 29360 2287 29372
rect 2343 29360 2367 29372
rect 2423 29360 2447 29372
rect 2503 29360 2527 29372
rect 2583 29360 2607 29372
rect 2663 29360 2695 29372
rect 2095 29308 2097 29360
rect 2285 29332 2287 29360
rect 2353 29332 2367 29360
rect 2423 29332 2437 29360
rect 2503 29332 2505 29360
rect 2149 29308 2165 29332
rect 2217 29308 2233 29332
rect 2285 29308 2301 29332
rect 2353 29308 2369 29332
rect 2421 29308 2437 29332
rect 2489 29308 2505 29332
rect 2557 29308 2573 29332
rect 2625 29308 2641 29332
rect 2693 29308 2695 29360
rect 2095 29307 2695 29308
rect 2095 29296 2127 29307
rect 2183 29296 2207 29307
rect 2263 29296 2287 29307
rect 2343 29296 2367 29307
rect 2423 29296 2447 29307
rect 2503 29296 2527 29307
rect 2583 29296 2607 29307
rect 2663 29296 2695 29307
rect 2095 29244 2097 29296
rect 2285 29251 2287 29296
rect 2353 29251 2367 29296
rect 2423 29251 2437 29296
rect 2503 29251 2505 29296
rect 2149 29244 2165 29251
rect 2217 29244 2233 29251
rect 2285 29244 2301 29251
rect 2353 29244 2369 29251
rect 2421 29244 2437 29251
rect 2489 29244 2505 29251
rect 2557 29244 2573 29251
rect 2625 29244 2641 29251
rect 2693 29244 2695 29296
rect 2095 29232 2695 29244
rect 2095 29180 2097 29232
rect 2149 29226 2165 29232
rect 2217 29226 2233 29232
rect 2285 29226 2301 29232
rect 2353 29226 2369 29232
rect 2421 29226 2437 29232
rect 2489 29226 2505 29232
rect 2557 29226 2573 29232
rect 2625 29226 2641 29232
rect 2285 29180 2287 29226
rect 2353 29180 2367 29226
rect 2423 29180 2437 29226
rect 2503 29180 2505 29226
rect 2693 29180 2695 29232
rect 2095 29170 2127 29180
rect 2183 29170 2207 29180
rect 2263 29170 2287 29180
rect 2343 29170 2367 29180
rect 2423 29170 2447 29180
rect 2503 29170 2527 29180
rect 2583 29170 2607 29180
rect 2663 29170 2695 29180
rect 2095 29168 2695 29170
rect 2095 29116 2097 29168
rect 2149 29145 2165 29168
rect 2217 29145 2233 29168
rect 2285 29145 2301 29168
rect 2353 29145 2369 29168
rect 2421 29145 2437 29168
rect 2489 29145 2505 29168
rect 2557 29145 2573 29168
rect 2625 29145 2641 29168
rect 2285 29116 2287 29145
rect 2353 29116 2367 29145
rect 2423 29116 2437 29145
rect 2503 29116 2505 29145
rect 2693 29116 2695 29168
rect 2095 29104 2127 29116
rect 2183 29104 2207 29116
rect 2263 29104 2287 29116
rect 2343 29104 2367 29116
rect 2423 29104 2447 29116
rect 2503 29104 2527 29116
rect 2583 29104 2607 29116
rect 2663 29104 2695 29116
rect 2095 29052 2097 29104
rect 2285 29089 2287 29104
rect 2353 29089 2367 29104
rect 2423 29089 2437 29104
rect 2503 29089 2505 29104
rect 2149 29064 2165 29089
rect 2217 29064 2233 29089
rect 2285 29064 2301 29089
rect 2353 29064 2369 29089
rect 2421 29064 2437 29089
rect 2489 29064 2505 29089
rect 2557 29064 2573 29089
rect 2625 29064 2641 29089
rect 2285 29052 2287 29064
rect 2353 29052 2367 29064
rect 2423 29052 2437 29064
rect 2503 29052 2505 29064
rect 2693 29052 2695 29104
rect 2095 29040 2127 29052
rect 2183 29040 2207 29052
rect 2263 29040 2287 29052
rect 2343 29040 2367 29052
rect 2423 29040 2447 29052
rect 2503 29040 2527 29052
rect 2583 29040 2607 29052
rect 2663 29040 2695 29052
rect 2095 28988 2097 29040
rect 2285 29008 2287 29040
rect 2353 29008 2367 29040
rect 2423 29008 2437 29040
rect 2503 29008 2505 29040
rect 2149 28988 2165 29008
rect 2217 28988 2233 29008
rect 2285 28988 2301 29008
rect 2353 28988 2369 29008
rect 2421 28988 2437 29008
rect 2489 28988 2505 29008
rect 2557 28988 2573 29008
rect 2625 28988 2641 29008
rect 2693 28988 2695 29040
rect 2095 28983 2695 28988
rect 2095 28976 2127 28983
rect 2183 28976 2207 28983
rect 2263 28976 2287 28983
rect 2343 28976 2367 28983
rect 2423 28976 2447 28983
rect 2503 28976 2527 28983
rect 2583 28976 2607 28983
rect 2663 28976 2695 28983
rect 2095 28924 2097 28976
rect 2285 28927 2287 28976
rect 2353 28927 2367 28976
rect 2423 28927 2437 28976
rect 2503 28927 2505 28976
rect 2149 28924 2165 28927
rect 2217 28924 2233 28927
rect 2285 28924 2301 28927
rect 2353 28924 2369 28927
rect 2421 28924 2437 28927
rect 2489 28924 2505 28927
rect 2557 28924 2573 28927
rect 2625 28924 2641 28927
rect 2693 28924 2695 28976
rect 2095 27865 2695 28924
rect 2095 27813 2097 27865
rect 2149 27862 2165 27865
rect 2217 27862 2233 27865
rect 2285 27862 2301 27865
rect 2353 27862 2369 27865
rect 2421 27862 2437 27865
rect 2489 27862 2505 27865
rect 2557 27862 2573 27865
rect 2625 27862 2641 27865
rect 2693 27813 2695 27865
rect 2095 27801 2127 27813
rect 2663 27801 2695 27813
rect 2095 27749 2097 27801
rect 2693 27749 2695 27801
rect 2095 27737 2127 27749
rect 2663 27737 2695 27749
rect 2095 27685 2097 27737
rect 2693 27685 2695 27737
rect 2095 27673 2127 27685
rect 2663 27673 2695 27685
rect 2095 27621 2097 27673
rect 2693 27621 2695 27673
rect 2095 27609 2127 27621
rect 2663 27609 2695 27621
rect 2095 27557 2097 27609
rect 2693 27557 2695 27609
rect 2095 27545 2127 27557
rect 2663 27545 2695 27557
rect 2095 27493 2097 27545
rect 2693 27493 2695 27545
rect 2095 27481 2127 27493
rect 2663 27481 2695 27493
rect 2095 27429 2097 27481
rect 2693 27429 2695 27481
rect 2095 27417 2127 27429
rect 2663 27417 2695 27429
rect 2095 27365 2097 27417
rect 2149 27381 2165 27406
rect 2217 27381 2233 27406
rect 2285 27381 2301 27406
rect 2353 27381 2369 27406
rect 2421 27381 2437 27406
rect 2489 27381 2505 27406
rect 2557 27381 2573 27406
rect 2625 27381 2641 27406
rect 2285 27365 2287 27381
rect 2353 27365 2367 27381
rect 2423 27365 2437 27381
rect 2503 27365 2505 27381
rect 2693 27365 2695 27417
rect 2095 27353 2127 27365
rect 2183 27353 2207 27365
rect 2263 27353 2287 27365
rect 2343 27353 2367 27365
rect 2423 27353 2447 27365
rect 2503 27353 2527 27365
rect 2583 27353 2607 27365
rect 2663 27353 2695 27365
rect 2095 27301 2097 27353
rect 2285 27325 2287 27353
rect 2353 27325 2367 27353
rect 2423 27325 2437 27353
rect 2503 27325 2505 27353
rect 2149 27301 2165 27325
rect 2217 27301 2233 27325
rect 2285 27301 2301 27325
rect 2353 27301 2369 27325
rect 2421 27301 2437 27325
rect 2489 27301 2505 27325
rect 2557 27301 2573 27325
rect 2625 27301 2641 27325
rect 2693 27301 2695 27353
rect 2095 27300 2695 27301
rect 2095 27289 2127 27300
rect 2183 27289 2207 27300
rect 2263 27289 2287 27300
rect 2343 27289 2367 27300
rect 2423 27289 2447 27300
rect 2503 27289 2527 27300
rect 2583 27289 2607 27300
rect 2663 27289 2695 27300
rect 2095 27237 2097 27289
rect 2285 27244 2287 27289
rect 2353 27244 2367 27289
rect 2423 27244 2437 27289
rect 2503 27244 2505 27289
rect 2149 27237 2165 27244
rect 2217 27237 2233 27244
rect 2285 27237 2301 27244
rect 2353 27237 2369 27244
rect 2421 27237 2437 27244
rect 2489 27237 2505 27244
rect 2557 27237 2573 27244
rect 2625 27237 2641 27244
rect 2693 27237 2695 27289
rect 2095 27225 2695 27237
rect 2095 27173 2097 27225
rect 2149 27219 2165 27225
rect 2217 27219 2233 27225
rect 2285 27219 2301 27225
rect 2353 27219 2369 27225
rect 2421 27219 2437 27225
rect 2489 27219 2505 27225
rect 2557 27219 2573 27225
rect 2625 27219 2641 27225
rect 2285 27173 2287 27219
rect 2353 27173 2367 27219
rect 2423 27173 2437 27219
rect 2503 27173 2505 27219
rect 2693 27173 2695 27225
rect 2095 27163 2127 27173
rect 2183 27163 2207 27173
rect 2263 27163 2287 27173
rect 2343 27163 2367 27173
rect 2423 27163 2447 27173
rect 2503 27163 2527 27173
rect 2583 27163 2607 27173
rect 2663 27163 2695 27173
rect 2095 27161 2695 27163
rect 2095 27109 2097 27161
rect 2149 27138 2165 27161
rect 2217 27138 2233 27161
rect 2285 27138 2301 27161
rect 2353 27138 2369 27161
rect 2421 27138 2437 27161
rect 2489 27138 2505 27161
rect 2557 27138 2573 27161
rect 2625 27138 2641 27161
rect 2285 27109 2287 27138
rect 2353 27109 2367 27138
rect 2423 27109 2437 27138
rect 2503 27109 2505 27138
rect 2693 27109 2695 27161
rect 2095 27097 2127 27109
rect 2183 27097 2207 27109
rect 2263 27097 2287 27109
rect 2343 27097 2367 27109
rect 2423 27097 2447 27109
rect 2503 27097 2527 27109
rect 2583 27097 2607 27109
rect 2663 27097 2695 27109
rect 2095 27045 2097 27097
rect 2285 27082 2287 27097
rect 2353 27082 2367 27097
rect 2423 27082 2437 27097
rect 2503 27082 2505 27097
rect 2149 27057 2165 27082
rect 2217 27057 2233 27082
rect 2285 27057 2301 27082
rect 2353 27057 2369 27082
rect 2421 27057 2437 27082
rect 2489 27057 2505 27082
rect 2557 27057 2573 27082
rect 2625 27057 2641 27082
rect 2285 27045 2287 27057
rect 2353 27045 2367 27057
rect 2423 27045 2437 27057
rect 2503 27045 2505 27057
rect 2693 27045 2695 27097
rect 2095 27033 2127 27045
rect 2183 27033 2207 27045
rect 2263 27033 2287 27045
rect 2343 27033 2367 27045
rect 2423 27033 2447 27045
rect 2503 27033 2527 27045
rect 2583 27033 2607 27045
rect 2663 27033 2695 27045
rect 2095 26981 2097 27033
rect 2285 27001 2287 27033
rect 2353 27001 2367 27033
rect 2423 27001 2437 27033
rect 2503 27001 2505 27033
rect 2149 26981 2165 27001
rect 2217 26981 2233 27001
rect 2285 26981 2301 27001
rect 2353 26981 2369 27001
rect 2421 26981 2437 27001
rect 2489 26981 2505 27001
rect 2557 26981 2573 27001
rect 2625 26981 2641 27001
rect 2693 26981 2695 27033
rect 2095 26976 2695 26981
rect 2095 26969 2127 26976
rect 2183 26969 2207 26976
rect 2263 26969 2287 26976
rect 2343 26969 2367 26976
rect 2423 26969 2447 26976
rect 2503 26969 2527 26976
rect 2583 26969 2607 26976
rect 2663 26969 2695 26976
rect 2095 26917 2097 26969
rect 2285 26920 2287 26969
rect 2353 26920 2367 26969
rect 2423 26920 2437 26969
rect 2503 26920 2505 26969
rect 2149 26917 2165 26920
rect 2217 26917 2233 26920
rect 2285 26917 2301 26920
rect 2353 26917 2369 26920
rect 2421 26917 2437 26920
rect 2489 26917 2505 26920
rect 2557 26917 2573 26920
rect 2625 26917 2641 26920
rect 2693 26917 2695 26969
rect 2095 25679 2695 26917
rect 2095 25627 2097 25679
rect 2149 25676 2165 25679
rect 2217 25676 2233 25679
rect 2285 25676 2301 25679
rect 2353 25676 2369 25679
rect 2421 25676 2437 25679
rect 2489 25676 2505 25679
rect 2557 25676 2573 25679
rect 2625 25676 2641 25679
rect 2693 25627 2695 25679
rect 2095 25615 2127 25627
rect 2663 25615 2695 25627
rect 2095 25563 2097 25615
rect 2693 25563 2695 25615
rect 2095 25551 2127 25563
rect 2663 25551 2695 25563
rect 2095 25499 2097 25551
rect 2693 25499 2695 25551
rect 2095 25487 2127 25499
rect 2663 25487 2695 25499
rect 2095 25435 2097 25487
rect 2693 25435 2695 25487
rect 2095 25423 2127 25435
rect 2663 25423 2695 25435
rect 2095 25371 2097 25423
rect 2693 25371 2695 25423
rect 2095 25359 2127 25371
rect 2663 25359 2695 25371
rect 2095 25307 2097 25359
rect 2693 25307 2695 25359
rect 2095 25295 2127 25307
rect 2663 25295 2695 25307
rect 2095 25243 2097 25295
rect 2693 25243 2695 25295
rect 2095 25231 2127 25243
rect 2663 25231 2695 25243
rect 2095 25179 2097 25231
rect 2149 25195 2165 25220
rect 2217 25195 2233 25220
rect 2285 25195 2301 25220
rect 2353 25195 2369 25220
rect 2421 25195 2437 25220
rect 2489 25195 2505 25220
rect 2557 25195 2573 25220
rect 2625 25195 2641 25220
rect 2285 25179 2287 25195
rect 2353 25179 2367 25195
rect 2423 25179 2437 25195
rect 2503 25179 2505 25195
rect 2693 25179 2695 25231
rect 2095 25167 2127 25179
rect 2183 25167 2207 25179
rect 2263 25167 2287 25179
rect 2343 25167 2367 25179
rect 2423 25167 2447 25179
rect 2503 25167 2527 25179
rect 2583 25167 2607 25179
rect 2663 25167 2695 25179
rect 2095 25115 2097 25167
rect 2285 25139 2287 25167
rect 2353 25139 2367 25167
rect 2423 25139 2437 25167
rect 2503 25139 2505 25167
rect 2149 25115 2165 25139
rect 2217 25115 2233 25139
rect 2285 25115 2301 25139
rect 2353 25115 2369 25139
rect 2421 25115 2437 25139
rect 2489 25115 2505 25139
rect 2557 25115 2573 25139
rect 2625 25115 2641 25139
rect 2693 25115 2695 25167
rect 2095 25114 2695 25115
rect 2095 25103 2127 25114
rect 2183 25103 2207 25114
rect 2263 25103 2287 25114
rect 2343 25103 2367 25114
rect 2423 25103 2447 25114
rect 2503 25103 2527 25114
rect 2583 25103 2607 25114
rect 2663 25103 2695 25114
rect 2095 25051 2097 25103
rect 2285 25058 2287 25103
rect 2353 25058 2367 25103
rect 2423 25058 2437 25103
rect 2503 25058 2505 25103
rect 2149 25051 2165 25058
rect 2217 25051 2233 25058
rect 2285 25051 2301 25058
rect 2353 25051 2369 25058
rect 2421 25051 2437 25058
rect 2489 25051 2505 25058
rect 2557 25051 2573 25058
rect 2625 25051 2641 25058
rect 2693 25051 2695 25103
rect 2095 25039 2695 25051
rect 2095 24987 2097 25039
rect 2149 25033 2165 25039
rect 2217 25033 2233 25039
rect 2285 25033 2301 25039
rect 2353 25033 2369 25039
rect 2421 25033 2437 25039
rect 2489 25033 2505 25039
rect 2557 25033 2573 25039
rect 2625 25033 2641 25039
rect 2285 24987 2287 25033
rect 2353 24987 2367 25033
rect 2423 24987 2437 25033
rect 2503 24987 2505 25033
rect 2693 24987 2695 25039
rect 2095 24977 2127 24987
rect 2183 24977 2207 24987
rect 2263 24977 2287 24987
rect 2343 24977 2367 24987
rect 2423 24977 2447 24987
rect 2503 24977 2527 24987
rect 2583 24977 2607 24987
rect 2663 24977 2695 24987
rect 2095 24975 2695 24977
rect 2095 24923 2097 24975
rect 2149 24952 2165 24975
rect 2217 24952 2233 24975
rect 2285 24952 2301 24975
rect 2353 24952 2369 24975
rect 2421 24952 2437 24975
rect 2489 24952 2505 24975
rect 2557 24952 2573 24975
rect 2625 24952 2641 24975
rect 2285 24923 2287 24952
rect 2353 24923 2367 24952
rect 2423 24923 2437 24952
rect 2503 24923 2505 24952
rect 2693 24923 2695 24975
rect 2095 24911 2127 24923
rect 2183 24911 2207 24923
rect 2263 24911 2287 24923
rect 2343 24911 2367 24923
rect 2423 24911 2447 24923
rect 2503 24911 2527 24923
rect 2583 24911 2607 24923
rect 2663 24911 2695 24923
rect 2095 24859 2097 24911
rect 2285 24896 2287 24911
rect 2353 24896 2367 24911
rect 2423 24896 2437 24911
rect 2503 24896 2505 24911
rect 2149 24871 2165 24896
rect 2217 24871 2233 24896
rect 2285 24871 2301 24896
rect 2353 24871 2369 24896
rect 2421 24871 2437 24896
rect 2489 24871 2505 24896
rect 2557 24871 2573 24896
rect 2625 24871 2641 24896
rect 2285 24859 2287 24871
rect 2353 24859 2367 24871
rect 2423 24859 2437 24871
rect 2503 24859 2505 24871
rect 2693 24859 2695 24911
rect 2095 24847 2127 24859
rect 2183 24847 2207 24859
rect 2263 24847 2287 24859
rect 2343 24847 2367 24859
rect 2423 24847 2447 24859
rect 2503 24847 2527 24859
rect 2583 24847 2607 24859
rect 2663 24847 2695 24859
rect 2095 24795 2097 24847
rect 2285 24815 2287 24847
rect 2353 24815 2367 24847
rect 2423 24815 2437 24847
rect 2503 24815 2505 24847
rect 2149 24795 2165 24815
rect 2217 24795 2233 24815
rect 2285 24795 2301 24815
rect 2353 24795 2369 24815
rect 2421 24795 2437 24815
rect 2489 24795 2505 24815
rect 2557 24795 2573 24815
rect 2625 24795 2641 24815
rect 2693 24795 2695 24847
rect 2095 24790 2695 24795
rect 2095 24783 2127 24790
rect 2183 24783 2207 24790
rect 2263 24783 2287 24790
rect 2343 24783 2367 24790
rect 2423 24783 2447 24790
rect 2503 24783 2527 24790
rect 2583 24783 2607 24790
rect 2663 24783 2695 24790
rect 2095 24731 2097 24783
rect 2285 24734 2287 24783
rect 2353 24734 2367 24783
rect 2423 24734 2437 24783
rect 2503 24734 2505 24783
rect 2149 24731 2165 24734
rect 2217 24731 2233 24734
rect 2285 24731 2301 24734
rect 2353 24731 2369 24734
rect 2421 24731 2437 24734
rect 2489 24731 2505 24734
rect 2557 24731 2573 24734
rect 2625 24731 2641 24734
rect 2693 24731 2695 24783
rect 2095 23531 2695 24731
rect 2095 23479 2097 23531
rect 2149 23528 2165 23531
rect 2217 23528 2233 23531
rect 2285 23528 2301 23531
rect 2353 23528 2369 23531
rect 2421 23528 2437 23531
rect 2489 23528 2505 23531
rect 2557 23528 2573 23531
rect 2625 23528 2641 23531
rect 2693 23479 2695 23531
rect 2095 23467 2127 23479
rect 2663 23467 2695 23479
rect 2095 23415 2097 23467
rect 2693 23415 2695 23467
rect 2095 23403 2127 23415
rect 2663 23403 2695 23415
rect 2095 23351 2097 23403
rect 2693 23351 2695 23403
rect 2095 23339 2127 23351
rect 2663 23339 2695 23351
rect 2095 23287 2097 23339
rect 2693 23287 2695 23339
rect 2095 23275 2127 23287
rect 2663 23275 2695 23287
rect 2095 23223 2097 23275
rect 2693 23223 2695 23275
rect 2095 23211 2127 23223
rect 2663 23211 2695 23223
rect 2095 23159 2097 23211
rect 2693 23159 2695 23211
rect 2095 23147 2127 23159
rect 2663 23147 2695 23159
rect 2095 23095 2097 23147
rect 2693 23095 2695 23147
rect 2095 23083 2127 23095
rect 2663 23083 2695 23095
rect 2095 23031 2097 23083
rect 2149 23047 2165 23072
rect 2217 23047 2233 23072
rect 2285 23047 2301 23072
rect 2353 23047 2369 23072
rect 2421 23047 2437 23072
rect 2489 23047 2505 23072
rect 2557 23047 2573 23072
rect 2625 23047 2641 23072
rect 2285 23031 2287 23047
rect 2353 23031 2367 23047
rect 2423 23031 2437 23047
rect 2503 23031 2505 23047
rect 2693 23031 2695 23083
rect 2095 23019 2127 23031
rect 2183 23019 2207 23031
rect 2263 23019 2287 23031
rect 2343 23019 2367 23031
rect 2423 23019 2447 23031
rect 2503 23019 2527 23031
rect 2583 23019 2607 23031
rect 2663 23019 2695 23031
rect 2095 22967 2097 23019
rect 2285 22991 2287 23019
rect 2353 22991 2367 23019
rect 2423 22991 2437 23019
rect 2503 22991 2505 23019
rect 2149 22967 2165 22991
rect 2217 22967 2233 22991
rect 2285 22967 2301 22991
rect 2353 22967 2369 22991
rect 2421 22967 2437 22991
rect 2489 22967 2505 22991
rect 2557 22967 2573 22991
rect 2625 22967 2641 22991
rect 2693 22967 2695 23019
rect 2095 22966 2695 22967
rect 2095 22955 2127 22966
rect 2183 22955 2207 22966
rect 2263 22955 2287 22966
rect 2343 22955 2367 22966
rect 2423 22955 2447 22966
rect 2503 22955 2527 22966
rect 2583 22955 2607 22966
rect 2663 22955 2695 22966
rect 2095 22903 2097 22955
rect 2285 22910 2287 22955
rect 2353 22910 2367 22955
rect 2423 22910 2437 22955
rect 2503 22910 2505 22955
rect 2149 22903 2165 22910
rect 2217 22903 2233 22910
rect 2285 22903 2301 22910
rect 2353 22903 2369 22910
rect 2421 22903 2437 22910
rect 2489 22903 2505 22910
rect 2557 22903 2573 22910
rect 2625 22903 2641 22910
rect 2693 22903 2695 22955
rect 2095 22891 2695 22903
rect 2095 22839 2097 22891
rect 2149 22885 2165 22891
rect 2217 22885 2233 22891
rect 2285 22885 2301 22891
rect 2353 22885 2369 22891
rect 2421 22885 2437 22891
rect 2489 22885 2505 22891
rect 2557 22885 2573 22891
rect 2625 22885 2641 22891
rect 2285 22839 2287 22885
rect 2353 22839 2367 22885
rect 2423 22839 2437 22885
rect 2503 22839 2505 22885
rect 2693 22839 2695 22891
rect 2095 22829 2127 22839
rect 2183 22829 2207 22839
rect 2263 22829 2287 22839
rect 2343 22829 2367 22839
rect 2423 22829 2447 22839
rect 2503 22829 2527 22839
rect 2583 22829 2607 22839
rect 2663 22829 2695 22839
rect 2095 22827 2695 22829
rect 2095 22775 2097 22827
rect 2149 22804 2165 22827
rect 2217 22804 2233 22827
rect 2285 22804 2301 22827
rect 2353 22804 2369 22827
rect 2421 22804 2437 22827
rect 2489 22804 2505 22827
rect 2557 22804 2573 22827
rect 2625 22804 2641 22827
rect 2285 22775 2287 22804
rect 2353 22775 2367 22804
rect 2423 22775 2437 22804
rect 2503 22775 2505 22804
rect 2693 22775 2695 22827
rect 2095 22763 2127 22775
rect 2183 22763 2207 22775
rect 2263 22763 2287 22775
rect 2343 22763 2367 22775
rect 2423 22763 2447 22775
rect 2503 22763 2527 22775
rect 2583 22763 2607 22775
rect 2663 22763 2695 22775
rect 2095 22711 2097 22763
rect 2285 22748 2287 22763
rect 2353 22748 2367 22763
rect 2423 22748 2437 22763
rect 2503 22748 2505 22763
rect 2149 22723 2165 22748
rect 2217 22723 2233 22748
rect 2285 22723 2301 22748
rect 2353 22723 2369 22748
rect 2421 22723 2437 22748
rect 2489 22723 2505 22748
rect 2557 22723 2573 22748
rect 2625 22723 2641 22748
rect 2285 22711 2287 22723
rect 2353 22711 2367 22723
rect 2423 22711 2437 22723
rect 2503 22711 2505 22723
rect 2693 22711 2695 22763
rect 2095 22699 2127 22711
rect 2183 22699 2207 22711
rect 2263 22699 2287 22711
rect 2343 22699 2367 22711
rect 2423 22699 2447 22711
rect 2503 22699 2527 22711
rect 2583 22699 2607 22711
rect 2663 22699 2695 22711
rect 2095 22647 2097 22699
rect 2285 22667 2287 22699
rect 2353 22667 2367 22699
rect 2423 22667 2437 22699
rect 2503 22667 2505 22699
rect 2149 22647 2165 22667
rect 2217 22647 2233 22667
rect 2285 22647 2301 22667
rect 2353 22647 2369 22667
rect 2421 22647 2437 22667
rect 2489 22647 2505 22667
rect 2557 22647 2573 22667
rect 2625 22647 2641 22667
rect 2693 22647 2695 22699
rect 2095 22642 2695 22647
rect 2095 22635 2127 22642
rect 2183 22635 2207 22642
rect 2263 22635 2287 22642
rect 2343 22635 2367 22642
rect 2423 22635 2447 22642
rect 2503 22635 2527 22642
rect 2583 22635 2607 22642
rect 2663 22635 2695 22642
rect 2095 22583 2097 22635
rect 2285 22586 2287 22635
rect 2353 22586 2367 22635
rect 2423 22586 2437 22635
rect 2503 22586 2505 22635
rect 2149 22583 2165 22586
rect 2217 22583 2233 22586
rect 2285 22583 2301 22586
rect 2353 22583 2369 22586
rect 2421 22583 2437 22586
rect 2489 22583 2505 22586
rect 2557 22583 2573 22586
rect 2625 22583 2641 22586
rect 2693 22583 2695 22635
rect 2095 21361 2695 22583
rect 2095 21309 2097 21361
rect 2149 21358 2165 21361
rect 2217 21358 2233 21361
rect 2285 21358 2301 21361
rect 2353 21358 2369 21361
rect 2421 21358 2437 21361
rect 2489 21358 2505 21361
rect 2557 21358 2573 21361
rect 2625 21358 2641 21361
rect 2693 21309 2695 21361
rect 2095 21297 2127 21309
rect 2663 21297 2695 21309
rect 2095 21245 2097 21297
rect 2693 21245 2695 21297
rect 2095 21233 2127 21245
rect 2663 21233 2695 21245
rect 2095 21181 2097 21233
rect 2693 21181 2695 21233
rect 2095 21169 2127 21181
rect 2663 21169 2695 21181
rect 2095 21117 2097 21169
rect 2693 21117 2695 21169
rect 2095 21105 2127 21117
rect 2663 21105 2695 21117
rect 2095 21053 2097 21105
rect 2693 21053 2695 21105
rect 2095 21041 2127 21053
rect 2663 21041 2695 21053
rect 2095 20989 2097 21041
rect 2693 20989 2695 21041
rect 2095 20977 2127 20989
rect 2663 20977 2695 20989
rect 2095 20925 2097 20977
rect 2693 20925 2695 20977
rect 2095 20913 2127 20925
rect 2663 20913 2695 20925
rect 2095 20861 2097 20913
rect 2149 20877 2165 20902
rect 2217 20877 2233 20902
rect 2285 20877 2301 20902
rect 2353 20877 2369 20902
rect 2421 20877 2437 20902
rect 2489 20877 2505 20902
rect 2557 20877 2573 20902
rect 2625 20877 2641 20902
rect 2285 20861 2287 20877
rect 2353 20861 2367 20877
rect 2423 20861 2437 20877
rect 2503 20861 2505 20877
rect 2693 20861 2695 20913
rect 2095 20849 2127 20861
rect 2183 20849 2207 20861
rect 2263 20849 2287 20861
rect 2343 20849 2367 20861
rect 2423 20849 2447 20861
rect 2503 20849 2527 20861
rect 2583 20849 2607 20861
rect 2663 20849 2695 20861
rect 2095 20797 2097 20849
rect 2285 20821 2287 20849
rect 2353 20821 2367 20849
rect 2423 20821 2437 20849
rect 2503 20821 2505 20849
rect 2149 20797 2165 20821
rect 2217 20797 2233 20821
rect 2285 20797 2301 20821
rect 2353 20797 2369 20821
rect 2421 20797 2437 20821
rect 2489 20797 2505 20821
rect 2557 20797 2573 20821
rect 2625 20797 2641 20821
rect 2693 20797 2695 20849
rect 2095 20796 2695 20797
rect 2095 20785 2127 20796
rect 2183 20785 2207 20796
rect 2263 20785 2287 20796
rect 2343 20785 2367 20796
rect 2423 20785 2447 20796
rect 2503 20785 2527 20796
rect 2583 20785 2607 20796
rect 2663 20785 2695 20796
rect 2095 20733 2097 20785
rect 2285 20740 2287 20785
rect 2353 20740 2367 20785
rect 2423 20740 2437 20785
rect 2503 20740 2505 20785
rect 2149 20733 2165 20740
rect 2217 20733 2233 20740
rect 2285 20733 2301 20740
rect 2353 20733 2369 20740
rect 2421 20733 2437 20740
rect 2489 20733 2505 20740
rect 2557 20733 2573 20740
rect 2625 20733 2641 20740
rect 2693 20733 2695 20785
rect 2095 20721 2695 20733
rect 2095 20669 2097 20721
rect 2149 20715 2165 20721
rect 2217 20715 2233 20721
rect 2285 20715 2301 20721
rect 2353 20715 2369 20721
rect 2421 20715 2437 20721
rect 2489 20715 2505 20721
rect 2557 20715 2573 20721
rect 2625 20715 2641 20721
rect 2285 20669 2287 20715
rect 2353 20669 2367 20715
rect 2423 20669 2437 20715
rect 2503 20669 2505 20715
rect 2693 20669 2695 20721
rect 2095 20659 2127 20669
rect 2183 20659 2207 20669
rect 2263 20659 2287 20669
rect 2343 20659 2367 20669
rect 2423 20659 2447 20669
rect 2503 20659 2527 20669
rect 2583 20659 2607 20669
rect 2663 20659 2695 20669
rect 2095 20657 2695 20659
rect 2095 20605 2097 20657
rect 2149 20634 2165 20657
rect 2217 20634 2233 20657
rect 2285 20634 2301 20657
rect 2353 20634 2369 20657
rect 2421 20634 2437 20657
rect 2489 20634 2505 20657
rect 2557 20634 2573 20657
rect 2625 20634 2641 20657
rect 2285 20605 2287 20634
rect 2353 20605 2367 20634
rect 2423 20605 2437 20634
rect 2503 20605 2505 20634
rect 2693 20605 2695 20657
rect 2095 20593 2127 20605
rect 2183 20593 2207 20605
rect 2263 20593 2287 20605
rect 2343 20593 2367 20605
rect 2423 20593 2447 20605
rect 2503 20593 2527 20605
rect 2583 20593 2607 20605
rect 2663 20593 2695 20605
rect 2095 20541 2097 20593
rect 2285 20578 2287 20593
rect 2353 20578 2367 20593
rect 2423 20578 2437 20593
rect 2503 20578 2505 20593
rect 2149 20553 2165 20578
rect 2217 20553 2233 20578
rect 2285 20553 2301 20578
rect 2353 20553 2369 20578
rect 2421 20553 2437 20578
rect 2489 20553 2505 20578
rect 2557 20553 2573 20578
rect 2625 20553 2641 20578
rect 2285 20541 2287 20553
rect 2353 20541 2367 20553
rect 2423 20541 2437 20553
rect 2503 20541 2505 20553
rect 2693 20541 2695 20593
rect 2095 20529 2127 20541
rect 2183 20529 2207 20541
rect 2263 20529 2287 20541
rect 2343 20529 2367 20541
rect 2423 20529 2447 20541
rect 2503 20529 2527 20541
rect 2583 20529 2607 20541
rect 2663 20529 2695 20541
rect 2095 20477 2097 20529
rect 2285 20497 2287 20529
rect 2353 20497 2367 20529
rect 2423 20497 2437 20529
rect 2503 20497 2505 20529
rect 2149 20477 2165 20497
rect 2217 20477 2233 20497
rect 2285 20477 2301 20497
rect 2353 20477 2369 20497
rect 2421 20477 2437 20497
rect 2489 20477 2505 20497
rect 2557 20477 2573 20497
rect 2625 20477 2641 20497
rect 2693 20477 2695 20529
rect 2095 20472 2695 20477
rect 2095 20465 2127 20472
rect 2183 20465 2207 20472
rect 2263 20465 2287 20472
rect 2343 20465 2367 20472
rect 2423 20465 2447 20472
rect 2503 20465 2527 20472
rect 2583 20465 2607 20472
rect 2663 20465 2695 20472
rect 2095 20413 2097 20465
rect 2285 20416 2287 20465
rect 2353 20416 2367 20465
rect 2423 20416 2437 20465
rect 2503 20416 2505 20465
rect 2149 20413 2165 20416
rect 2217 20413 2233 20416
rect 2285 20413 2301 20416
rect 2353 20413 2369 20416
rect 2421 20413 2437 20416
rect 2489 20413 2505 20416
rect 2557 20413 2573 20416
rect 2625 20413 2641 20416
rect 2693 20413 2695 20465
rect 2095 19257 2695 20413
rect 2095 19205 2097 19257
rect 2149 19254 2165 19257
rect 2217 19254 2233 19257
rect 2285 19254 2301 19257
rect 2353 19254 2369 19257
rect 2421 19254 2437 19257
rect 2489 19254 2505 19257
rect 2557 19254 2573 19257
rect 2625 19254 2641 19257
rect 2693 19205 2695 19257
rect 2095 19193 2127 19205
rect 2663 19193 2695 19205
rect 2095 19141 2097 19193
rect 2693 19141 2695 19193
rect 2095 19129 2127 19141
rect 2663 19129 2695 19141
rect 2095 19077 2097 19129
rect 2693 19077 2695 19129
rect 2095 19065 2127 19077
rect 2663 19065 2695 19077
rect 2095 19013 2097 19065
rect 2693 19013 2695 19065
rect 2095 19001 2127 19013
rect 2663 19001 2695 19013
rect 2095 18949 2097 19001
rect 2693 18949 2695 19001
rect 2095 18937 2127 18949
rect 2663 18937 2695 18949
rect 2095 18885 2097 18937
rect 2693 18885 2695 18937
rect 2095 18873 2127 18885
rect 2663 18873 2695 18885
rect 2095 18821 2097 18873
rect 2693 18821 2695 18873
rect 2095 18809 2127 18821
rect 2663 18809 2695 18821
rect 2095 18757 2097 18809
rect 2149 18773 2165 18798
rect 2217 18773 2233 18798
rect 2285 18773 2301 18798
rect 2353 18773 2369 18798
rect 2421 18773 2437 18798
rect 2489 18773 2505 18798
rect 2557 18773 2573 18798
rect 2625 18773 2641 18798
rect 2285 18757 2287 18773
rect 2353 18757 2367 18773
rect 2423 18757 2437 18773
rect 2503 18757 2505 18773
rect 2693 18757 2695 18809
rect 2095 18745 2127 18757
rect 2183 18745 2207 18757
rect 2263 18745 2287 18757
rect 2343 18745 2367 18757
rect 2423 18745 2447 18757
rect 2503 18745 2527 18757
rect 2583 18745 2607 18757
rect 2663 18745 2695 18757
rect 2095 18693 2097 18745
rect 2285 18717 2287 18745
rect 2353 18717 2367 18745
rect 2423 18717 2437 18745
rect 2503 18717 2505 18745
rect 2149 18693 2165 18717
rect 2217 18693 2233 18717
rect 2285 18693 2301 18717
rect 2353 18693 2369 18717
rect 2421 18693 2437 18717
rect 2489 18693 2505 18717
rect 2557 18693 2573 18717
rect 2625 18693 2641 18717
rect 2693 18693 2695 18745
rect 2095 18692 2695 18693
rect 2095 18681 2127 18692
rect 2183 18681 2207 18692
rect 2263 18681 2287 18692
rect 2343 18681 2367 18692
rect 2423 18681 2447 18692
rect 2503 18681 2527 18692
rect 2583 18681 2607 18692
rect 2663 18681 2695 18692
rect 2095 18629 2097 18681
rect 2285 18636 2287 18681
rect 2353 18636 2367 18681
rect 2423 18636 2437 18681
rect 2503 18636 2505 18681
rect 2149 18629 2165 18636
rect 2217 18629 2233 18636
rect 2285 18629 2301 18636
rect 2353 18629 2369 18636
rect 2421 18629 2437 18636
rect 2489 18629 2505 18636
rect 2557 18629 2573 18636
rect 2625 18629 2641 18636
rect 2693 18629 2695 18681
rect 2095 18617 2695 18629
rect 2095 18565 2097 18617
rect 2149 18611 2165 18617
rect 2217 18611 2233 18617
rect 2285 18611 2301 18617
rect 2353 18611 2369 18617
rect 2421 18611 2437 18617
rect 2489 18611 2505 18617
rect 2557 18611 2573 18617
rect 2625 18611 2641 18617
rect 2285 18565 2287 18611
rect 2353 18565 2367 18611
rect 2423 18565 2437 18611
rect 2503 18565 2505 18611
rect 2693 18565 2695 18617
rect 2095 18555 2127 18565
rect 2183 18555 2207 18565
rect 2263 18555 2287 18565
rect 2343 18555 2367 18565
rect 2423 18555 2447 18565
rect 2503 18555 2527 18565
rect 2583 18555 2607 18565
rect 2663 18555 2695 18565
rect 2095 18553 2695 18555
rect 2095 18501 2097 18553
rect 2149 18530 2165 18553
rect 2217 18530 2233 18553
rect 2285 18530 2301 18553
rect 2353 18530 2369 18553
rect 2421 18530 2437 18553
rect 2489 18530 2505 18553
rect 2557 18530 2573 18553
rect 2625 18530 2641 18553
rect 2285 18501 2287 18530
rect 2353 18501 2367 18530
rect 2423 18501 2437 18530
rect 2503 18501 2505 18530
rect 2693 18501 2695 18553
rect 2095 18489 2127 18501
rect 2183 18489 2207 18501
rect 2263 18489 2287 18501
rect 2343 18489 2367 18501
rect 2423 18489 2447 18501
rect 2503 18489 2527 18501
rect 2583 18489 2607 18501
rect 2663 18489 2695 18501
rect 2095 18437 2097 18489
rect 2285 18474 2287 18489
rect 2353 18474 2367 18489
rect 2423 18474 2437 18489
rect 2503 18474 2505 18489
rect 2149 18449 2165 18474
rect 2217 18449 2233 18474
rect 2285 18449 2301 18474
rect 2353 18449 2369 18474
rect 2421 18449 2437 18474
rect 2489 18449 2505 18474
rect 2557 18449 2573 18474
rect 2625 18449 2641 18474
rect 2285 18437 2287 18449
rect 2353 18437 2367 18449
rect 2423 18437 2437 18449
rect 2503 18437 2505 18449
rect 2693 18437 2695 18489
rect 2095 18425 2127 18437
rect 2183 18425 2207 18437
rect 2263 18425 2287 18437
rect 2343 18425 2367 18437
rect 2423 18425 2447 18437
rect 2503 18425 2527 18437
rect 2583 18425 2607 18437
rect 2663 18425 2695 18437
rect 2095 18373 2097 18425
rect 2285 18393 2287 18425
rect 2353 18393 2367 18425
rect 2423 18393 2437 18425
rect 2503 18393 2505 18425
rect 2149 18373 2165 18393
rect 2217 18373 2233 18393
rect 2285 18373 2301 18393
rect 2353 18373 2369 18393
rect 2421 18373 2437 18393
rect 2489 18373 2505 18393
rect 2557 18373 2573 18393
rect 2625 18373 2641 18393
rect 2693 18373 2695 18425
rect 2095 18368 2695 18373
rect 2095 18361 2127 18368
rect 2183 18361 2207 18368
rect 2263 18361 2287 18368
rect 2343 18361 2367 18368
rect 2423 18361 2447 18368
rect 2503 18361 2527 18368
rect 2583 18361 2607 18368
rect 2663 18361 2695 18368
rect 2095 18309 2097 18361
rect 2285 18312 2287 18361
rect 2353 18312 2367 18361
rect 2423 18312 2437 18361
rect 2503 18312 2505 18361
rect 2149 18309 2165 18312
rect 2217 18309 2233 18312
rect 2285 18309 2301 18312
rect 2353 18309 2369 18312
rect 2421 18309 2437 18312
rect 2489 18309 2505 18312
rect 2557 18309 2573 18312
rect 2625 18309 2641 18312
rect 2693 18309 2695 18361
rect 2095 17146 2695 18309
rect 2095 17094 2097 17146
rect 2149 17143 2165 17146
rect 2217 17143 2233 17146
rect 2285 17143 2301 17146
rect 2353 17143 2369 17146
rect 2421 17143 2437 17146
rect 2489 17143 2505 17146
rect 2557 17143 2573 17146
rect 2625 17143 2641 17146
rect 2693 17094 2695 17146
rect 2095 17082 2127 17094
rect 2663 17082 2695 17094
rect 2095 17030 2097 17082
rect 2693 17030 2695 17082
rect 2095 17018 2127 17030
rect 2663 17018 2695 17030
rect 2095 16966 2097 17018
rect 2693 16966 2695 17018
rect 2095 16954 2127 16966
rect 2663 16954 2695 16966
rect 2095 16902 2097 16954
rect 2693 16902 2695 16954
rect 2095 16890 2127 16902
rect 2663 16890 2695 16902
rect 2095 16838 2097 16890
rect 2693 16838 2695 16890
rect 2095 16826 2127 16838
rect 2663 16826 2695 16838
rect 2095 16774 2097 16826
rect 2693 16774 2695 16826
rect 2095 16762 2127 16774
rect 2663 16762 2695 16774
rect 2095 16710 2097 16762
rect 2693 16710 2695 16762
rect 2095 16698 2127 16710
rect 2663 16698 2695 16710
rect 2095 16646 2097 16698
rect 2149 16662 2165 16687
rect 2217 16662 2233 16687
rect 2285 16662 2301 16687
rect 2353 16662 2369 16687
rect 2421 16662 2437 16687
rect 2489 16662 2505 16687
rect 2557 16662 2573 16687
rect 2625 16662 2641 16687
rect 2285 16646 2287 16662
rect 2353 16646 2367 16662
rect 2423 16646 2437 16662
rect 2503 16646 2505 16662
rect 2693 16646 2695 16698
rect 2095 16634 2127 16646
rect 2183 16634 2207 16646
rect 2263 16634 2287 16646
rect 2343 16634 2367 16646
rect 2423 16634 2447 16646
rect 2503 16634 2527 16646
rect 2583 16634 2607 16646
rect 2663 16634 2695 16646
rect 2095 16582 2097 16634
rect 2285 16606 2287 16634
rect 2353 16606 2367 16634
rect 2423 16606 2437 16634
rect 2503 16606 2505 16634
rect 2149 16582 2165 16606
rect 2217 16582 2233 16606
rect 2285 16582 2301 16606
rect 2353 16582 2369 16606
rect 2421 16582 2437 16606
rect 2489 16582 2505 16606
rect 2557 16582 2573 16606
rect 2625 16582 2641 16606
rect 2693 16582 2695 16634
rect 2095 16581 2695 16582
rect 2095 16570 2127 16581
rect 2183 16570 2207 16581
rect 2263 16570 2287 16581
rect 2343 16570 2367 16581
rect 2423 16570 2447 16581
rect 2503 16570 2527 16581
rect 2583 16570 2607 16581
rect 2663 16570 2695 16581
rect 2095 16518 2097 16570
rect 2285 16525 2287 16570
rect 2353 16525 2367 16570
rect 2423 16525 2437 16570
rect 2503 16525 2505 16570
rect 2149 16518 2165 16525
rect 2217 16518 2233 16525
rect 2285 16518 2301 16525
rect 2353 16518 2369 16525
rect 2421 16518 2437 16525
rect 2489 16518 2505 16525
rect 2557 16518 2573 16525
rect 2625 16518 2641 16525
rect 2693 16518 2695 16570
rect 2095 16506 2695 16518
rect 2095 16454 2097 16506
rect 2149 16500 2165 16506
rect 2217 16500 2233 16506
rect 2285 16500 2301 16506
rect 2353 16500 2369 16506
rect 2421 16500 2437 16506
rect 2489 16500 2505 16506
rect 2557 16500 2573 16506
rect 2625 16500 2641 16506
rect 2285 16454 2287 16500
rect 2353 16454 2367 16500
rect 2423 16454 2437 16500
rect 2503 16454 2505 16500
rect 2693 16454 2695 16506
rect 2095 16444 2127 16454
rect 2183 16444 2207 16454
rect 2263 16444 2287 16454
rect 2343 16444 2367 16454
rect 2423 16444 2447 16454
rect 2503 16444 2527 16454
rect 2583 16444 2607 16454
rect 2663 16444 2695 16454
rect 2095 16442 2695 16444
rect 2095 16390 2097 16442
rect 2149 16419 2165 16442
rect 2217 16419 2233 16442
rect 2285 16419 2301 16442
rect 2353 16419 2369 16442
rect 2421 16419 2437 16442
rect 2489 16419 2505 16442
rect 2557 16419 2573 16442
rect 2625 16419 2641 16442
rect 2285 16390 2287 16419
rect 2353 16390 2367 16419
rect 2423 16390 2437 16419
rect 2503 16390 2505 16419
rect 2693 16390 2695 16442
rect 2095 16378 2127 16390
rect 2183 16378 2207 16390
rect 2263 16378 2287 16390
rect 2343 16378 2367 16390
rect 2423 16378 2447 16390
rect 2503 16378 2527 16390
rect 2583 16378 2607 16390
rect 2663 16378 2695 16390
rect 2095 16326 2097 16378
rect 2285 16363 2287 16378
rect 2353 16363 2367 16378
rect 2423 16363 2437 16378
rect 2503 16363 2505 16378
rect 2149 16338 2165 16363
rect 2217 16338 2233 16363
rect 2285 16338 2301 16363
rect 2353 16338 2369 16363
rect 2421 16338 2437 16363
rect 2489 16338 2505 16363
rect 2557 16338 2573 16363
rect 2625 16338 2641 16363
rect 2285 16326 2287 16338
rect 2353 16326 2367 16338
rect 2423 16326 2437 16338
rect 2503 16326 2505 16338
rect 2693 16326 2695 16378
rect 2095 16314 2127 16326
rect 2183 16314 2207 16326
rect 2263 16314 2287 16326
rect 2343 16314 2367 16326
rect 2423 16314 2447 16326
rect 2503 16314 2527 16326
rect 2583 16314 2607 16326
rect 2663 16314 2695 16326
rect 2095 16262 2097 16314
rect 2285 16282 2287 16314
rect 2353 16282 2367 16314
rect 2423 16282 2437 16314
rect 2503 16282 2505 16314
rect 2149 16262 2165 16282
rect 2217 16262 2233 16282
rect 2285 16262 2301 16282
rect 2353 16262 2369 16282
rect 2421 16262 2437 16282
rect 2489 16262 2505 16282
rect 2557 16262 2573 16282
rect 2625 16262 2641 16282
rect 2693 16262 2695 16314
rect 2095 16257 2695 16262
rect 2095 16250 2127 16257
rect 2183 16250 2207 16257
rect 2263 16250 2287 16257
rect 2343 16250 2367 16257
rect 2423 16250 2447 16257
rect 2503 16250 2527 16257
rect 2583 16250 2607 16257
rect 2663 16250 2695 16257
rect 2095 16198 2097 16250
rect 2285 16201 2287 16250
rect 2353 16201 2367 16250
rect 2423 16201 2437 16250
rect 2503 16201 2505 16250
rect 2149 16198 2165 16201
rect 2217 16198 2233 16201
rect 2285 16198 2301 16201
rect 2353 16198 2369 16201
rect 2421 16198 2437 16201
rect 2489 16198 2505 16201
rect 2557 16198 2573 16201
rect 2625 16198 2641 16201
rect 2693 16198 2695 16250
rect 2095 15009 2695 16198
rect 2095 14957 2097 15009
rect 2149 15006 2165 15009
rect 2217 15006 2233 15009
rect 2285 15006 2301 15009
rect 2353 15006 2369 15009
rect 2421 15006 2437 15009
rect 2489 15006 2505 15009
rect 2557 15006 2573 15009
rect 2625 15006 2641 15009
rect 2693 14957 2695 15009
rect 2095 14945 2127 14957
rect 2663 14945 2695 14957
rect 2095 14893 2097 14945
rect 2693 14893 2695 14945
rect 2095 14881 2127 14893
rect 2663 14881 2695 14893
rect 2095 14829 2097 14881
rect 2693 14829 2695 14881
rect 2095 14817 2127 14829
rect 2663 14817 2695 14829
rect 2095 14765 2097 14817
rect 2693 14765 2695 14817
rect 2095 14753 2127 14765
rect 2663 14753 2695 14765
rect 2095 14701 2097 14753
rect 2693 14701 2695 14753
rect 2095 14689 2127 14701
rect 2663 14689 2695 14701
rect 2095 14637 2097 14689
rect 2693 14637 2695 14689
rect 2095 14625 2127 14637
rect 2663 14625 2695 14637
rect 2095 14573 2097 14625
rect 2693 14573 2695 14625
rect 2095 14561 2127 14573
rect 2663 14561 2695 14573
rect 2095 14509 2097 14561
rect 2149 14525 2165 14550
rect 2217 14525 2233 14550
rect 2285 14525 2301 14550
rect 2353 14525 2369 14550
rect 2421 14525 2437 14550
rect 2489 14525 2505 14550
rect 2557 14525 2573 14550
rect 2625 14525 2641 14550
rect 2285 14509 2287 14525
rect 2353 14509 2367 14525
rect 2423 14509 2437 14525
rect 2503 14509 2505 14525
rect 2693 14509 2695 14561
rect 2095 14497 2127 14509
rect 2183 14497 2207 14509
rect 2263 14497 2287 14509
rect 2343 14497 2367 14509
rect 2423 14497 2447 14509
rect 2503 14497 2527 14509
rect 2583 14497 2607 14509
rect 2663 14497 2695 14509
rect 2095 14445 2097 14497
rect 2285 14469 2287 14497
rect 2353 14469 2367 14497
rect 2423 14469 2437 14497
rect 2503 14469 2505 14497
rect 2149 14445 2165 14469
rect 2217 14445 2233 14469
rect 2285 14445 2301 14469
rect 2353 14445 2369 14469
rect 2421 14445 2437 14469
rect 2489 14445 2505 14469
rect 2557 14445 2573 14469
rect 2625 14445 2641 14469
rect 2693 14445 2695 14497
rect 2095 14444 2695 14445
rect 2095 14433 2127 14444
rect 2183 14433 2207 14444
rect 2263 14433 2287 14444
rect 2343 14433 2367 14444
rect 2423 14433 2447 14444
rect 2503 14433 2527 14444
rect 2583 14433 2607 14444
rect 2663 14433 2695 14444
rect 2095 14381 2097 14433
rect 2285 14388 2287 14433
rect 2353 14388 2367 14433
rect 2423 14388 2437 14433
rect 2503 14388 2505 14433
rect 2149 14381 2165 14388
rect 2217 14381 2233 14388
rect 2285 14381 2301 14388
rect 2353 14381 2369 14388
rect 2421 14381 2437 14388
rect 2489 14381 2505 14388
rect 2557 14381 2573 14388
rect 2625 14381 2641 14388
rect 2693 14381 2695 14433
rect 2095 14369 2695 14381
rect 2095 14317 2097 14369
rect 2149 14363 2165 14369
rect 2217 14363 2233 14369
rect 2285 14363 2301 14369
rect 2353 14363 2369 14369
rect 2421 14363 2437 14369
rect 2489 14363 2505 14369
rect 2557 14363 2573 14369
rect 2625 14363 2641 14369
rect 2285 14317 2287 14363
rect 2353 14317 2367 14363
rect 2423 14317 2437 14363
rect 2503 14317 2505 14363
rect 2693 14317 2695 14369
rect 2095 14307 2127 14317
rect 2183 14307 2207 14317
rect 2263 14307 2287 14317
rect 2343 14307 2367 14317
rect 2423 14307 2447 14317
rect 2503 14307 2527 14317
rect 2583 14307 2607 14317
rect 2663 14307 2695 14317
rect 2095 14305 2695 14307
rect 2095 14253 2097 14305
rect 2149 14282 2165 14305
rect 2217 14282 2233 14305
rect 2285 14282 2301 14305
rect 2353 14282 2369 14305
rect 2421 14282 2437 14305
rect 2489 14282 2505 14305
rect 2557 14282 2573 14305
rect 2625 14282 2641 14305
rect 2285 14253 2287 14282
rect 2353 14253 2367 14282
rect 2423 14253 2437 14282
rect 2503 14253 2505 14282
rect 2693 14253 2695 14305
rect 2095 14241 2127 14253
rect 2183 14241 2207 14253
rect 2263 14241 2287 14253
rect 2343 14241 2367 14253
rect 2423 14241 2447 14253
rect 2503 14241 2527 14253
rect 2583 14241 2607 14253
rect 2663 14241 2695 14253
rect 2095 14189 2097 14241
rect 2285 14226 2287 14241
rect 2353 14226 2367 14241
rect 2423 14226 2437 14241
rect 2503 14226 2505 14241
rect 2149 14201 2165 14226
rect 2217 14201 2233 14226
rect 2285 14201 2301 14226
rect 2353 14201 2369 14226
rect 2421 14201 2437 14226
rect 2489 14201 2505 14226
rect 2557 14201 2573 14226
rect 2625 14201 2641 14226
rect 2285 14189 2287 14201
rect 2353 14189 2367 14201
rect 2423 14189 2437 14201
rect 2503 14189 2505 14201
rect 2693 14189 2695 14241
rect 2095 14177 2127 14189
rect 2183 14177 2207 14189
rect 2263 14177 2287 14189
rect 2343 14177 2367 14189
rect 2423 14177 2447 14189
rect 2503 14177 2527 14189
rect 2583 14177 2607 14189
rect 2663 14177 2695 14189
rect 2095 14125 2097 14177
rect 2285 14145 2287 14177
rect 2353 14145 2367 14177
rect 2423 14145 2437 14177
rect 2503 14145 2505 14177
rect 2149 14125 2165 14145
rect 2217 14125 2233 14145
rect 2285 14125 2301 14145
rect 2353 14125 2369 14145
rect 2421 14125 2437 14145
rect 2489 14125 2505 14145
rect 2557 14125 2573 14145
rect 2625 14125 2641 14145
rect 2693 14125 2695 14177
rect 2095 14120 2695 14125
rect 2095 14113 2127 14120
rect 2183 14113 2207 14120
rect 2263 14113 2287 14120
rect 2343 14113 2367 14120
rect 2423 14113 2447 14120
rect 2503 14113 2527 14120
rect 2583 14113 2607 14120
rect 2663 14113 2695 14120
rect 2095 14061 2097 14113
rect 2285 14064 2287 14113
rect 2353 14064 2367 14113
rect 2423 14064 2437 14113
rect 2503 14064 2505 14113
rect 2149 14061 2165 14064
rect 2217 14061 2233 14064
rect 2285 14061 2301 14064
rect 2353 14061 2369 14064
rect 2421 14061 2437 14064
rect 2489 14061 2505 14064
rect 2557 14061 2573 14064
rect 2625 14061 2641 14064
rect 2693 14061 2695 14113
rect 2095 12907 2695 14061
rect 2095 12855 2097 12907
rect 2149 12904 2165 12907
rect 2217 12904 2233 12907
rect 2285 12904 2301 12907
rect 2353 12904 2369 12907
rect 2421 12904 2437 12907
rect 2489 12904 2505 12907
rect 2557 12904 2573 12907
rect 2625 12904 2641 12907
rect 2693 12855 2695 12907
rect 2095 12843 2127 12855
rect 2663 12843 2695 12855
rect 2095 12791 2097 12843
rect 2693 12791 2695 12843
rect 3285 13701 3341 13707
rect 3285 13698 3287 13701
rect 3339 13698 3341 13701
rect 3285 13633 3341 13642
rect 3285 13617 3287 13633
rect 3339 13617 3341 13633
rect 3285 13536 3287 13561
rect 3339 13536 3341 13561
rect 3285 13455 3287 13480
rect 3339 13455 3341 13480
rect 3285 13375 3287 13399
rect 3339 13375 3341 13399
rect 3285 13374 3341 13375
rect 3285 13306 3287 13318
rect 3339 13306 3341 13318
rect 3285 13292 3341 13306
rect 3285 13220 3341 13236
rect 3285 13210 3287 13220
rect 3339 13210 3341 13220
rect 3285 13151 3341 13154
rect 3285 13128 3287 13151
rect 3339 13128 3341 13151
rect 3285 13046 3287 13072
rect 3339 13046 3341 13072
rect 3285 12964 3287 12990
rect 3339 12964 3341 12990
rect 3285 12892 3287 12908
rect 3339 12892 3341 12908
rect 3285 12882 3341 12892
rect 3285 12823 3287 12826
rect 3339 12823 3341 12826
rect 3285 12817 3341 12823
rect 2095 12779 2127 12791
rect 2663 12779 2695 12791
rect 2095 12727 2097 12779
rect 2693 12727 2695 12779
rect 2095 12715 2127 12727
rect 2663 12715 2695 12727
rect 2095 12663 2097 12715
rect 2693 12663 2695 12715
rect 2095 12651 2127 12663
rect 2663 12651 2695 12663
rect 2095 12599 2097 12651
rect 2693 12599 2695 12651
rect 2095 12587 2127 12599
rect 2663 12587 2695 12599
rect 2095 12535 2097 12587
rect 2693 12535 2695 12587
rect 2095 12523 2127 12535
rect 2663 12523 2695 12535
rect 2095 12471 2097 12523
rect 2693 12471 2695 12523
rect 2095 12459 2127 12471
rect 2663 12459 2695 12471
rect 2095 12407 2097 12459
rect 2149 12423 2165 12448
rect 2217 12423 2233 12448
rect 2285 12423 2301 12448
rect 2353 12423 2369 12448
rect 2421 12423 2437 12448
rect 2489 12423 2505 12448
rect 2557 12423 2573 12448
rect 2625 12423 2641 12448
rect 2285 12407 2287 12423
rect 2353 12407 2367 12423
rect 2423 12407 2437 12423
rect 2503 12407 2505 12423
rect 2693 12407 2695 12459
rect 2095 12395 2127 12407
rect 2183 12395 2207 12407
rect 2263 12395 2287 12407
rect 2343 12395 2367 12407
rect 2423 12395 2447 12407
rect 2503 12395 2527 12407
rect 2583 12395 2607 12407
rect 2663 12395 2695 12407
rect 2095 12343 2097 12395
rect 2285 12367 2287 12395
rect 2353 12367 2367 12395
rect 2423 12367 2437 12395
rect 2503 12367 2505 12395
rect 2149 12343 2165 12367
rect 2217 12343 2233 12367
rect 2285 12343 2301 12367
rect 2353 12343 2369 12367
rect 2421 12343 2437 12367
rect 2489 12343 2505 12367
rect 2557 12343 2573 12367
rect 2625 12343 2641 12367
rect 2693 12343 2695 12395
rect 2095 12342 2695 12343
rect 2095 12331 2127 12342
rect 2183 12331 2207 12342
rect 2263 12331 2287 12342
rect 2343 12331 2367 12342
rect 2423 12331 2447 12342
rect 2503 12331 2527 12342
rect 2583 12331 2607 12342
rect 2663 12331 2695 12342
rect 2095 12279 2097 12331
rect 2285 12286 2287 12331
rect 2353 12286 2367 12331
rect 2423 12286 2437 12331
rect 2503 12286 2505 12331
rect 2149 12279 2165 12286
rect 2217 12279 2233 12286
rect 2285 12279 2301 12286
rect 2353 12279 2369 12286
rect 2421 12279 2437 12286
rect 2489 12279 2505 12286
rect 2557 12279 2573 12286
rect 2625 12279 2641 12286
rect 2693 12279 2695 12331
rect 2095 12267 2695 12279
rect 2095 12215 2097 12267
rect 2149 12261 2165 12267
rect 2217 12261 2233 12267
rect 2285 12261 2301 12267
rect 2353 12261 2369 12267
rect 2421 12261 2437 12267
rect 2489 12261 2505 12267
rect 2557 12261 2573 12267
rect 2625 12261 2641 12267
rect 2285 12215 2287 12261
rect 2353 12215 2367 12261
rect 2423 12215 2437 12261
rect 2503 12215 2505 12261
rect 2693 12215 2695 12267
rect 2095 12205 2127 12215
rect 2183 12205 2207 12215
rect 2263 12205 2287 12215
rect 2343 12205 2367 12215
rect 2423 12205 2447 12215
rect 2503 12205 2527 12215
rect 2583 12205 2607 12215
rect 2663 12205 2695 12215
rect 2095 12203 2695 12205
rect 2095 12151 2097 12203
rect 2149 12180 2165 12203
rect 2217 12180 2233 12203
rect 2285 12180 2301 12203
rect 2353 12180 2369 12203
rect 2421 12180 2437 12203
rect 2489 12180 2505 12203
rect 2557 12180 2573 12203
rect 2625 12180 2641 12203
rect 2285 12151 2287 12180
rect 2353 12151 2367 12180
rect 2423 12151 2437 12180
rect 2503 12151 2505 12180
rect 2693 12151 2695 12203
rect 2095 12139 2127 12151
rect 2183 12139 2207 12151
rect 2263 12139 2287 12151
rect 2343 12139 2367 12151
rect 2423 12139 2447 12151
rect 2503 12139 2527 12151
rect 2583 12139 2607 12151
rect 2663 12139 2695 12151
rect 2095 12087 2097 12139
rect 2285 12124 2287 12139
rect 2353 12124 2367 12139
rect 2423 12124 2437 12139
rect 2503 12124 2505 12139
rect 2149 12099 2165 12124
rect 2217 12099 2233 12124
rect 2285 12099 2301 12124
rect 2353 12099 2369 12124
rect 2421 12099 2437 12124
rect 2489 12099 2505 12124
rect 2557 12099 2573 12124
rect 2625 12099 2641 12124
rect 2285 12087 2287 12099
rect 2353 12087 2367 12099
rect 2423 12087 2437 12099
rect 2503 12087 2505 12099
rect 2693 12087 2695 12139
rect 2095 12075 2127 12087
rect 2183 12075 2207 12087
rect 2263 12075 2287 12087
rect 2343 12075 2367 12087
rect 2423 12075 2447 12087
rect 2503 12075 2527 12087
rect 2583 12075 2607 12087
rect 2663 12075 2695 12087
rect 2095 12023 2097 12075
rect 2285 12043 2287 12075
rect 2353 12043 2367 12075
rect 2423 12043 2437 12075
rect 2503 12043 2505 12075
rect 2149 12023 2165 12043
rect 2217 12023 2233 12043
rect 2285 12023 2301 12043
rect 2353 12023 2369 12043
rect 2421 12023 2437 12043
rect 2489 12023 2505 12043
rect 2557 12023 2573 12043
rect 2625 12023 2641 12043
rect 2693 12023 2695 12075
rect 2095 12018 2695 12023
rect 2095 12011 2127 12018
rect 2183 12011 2207 12018
rect 2263 12011 2287 12018
rect 2343 12011 2367 12018
rect 2423 12011 2447 12018
rect 2503 12011 2527 12018
rect 2583 12011 2607 12018
rect 2663 12011 2695 12018
rect 2095 11959 2097 12011
rect 2285 11962 2287 12011
rect 2353 11962 2367 12011
rect 2423 11962 2437 12011
rect 2503 11962 2505 12011
rect 2149 11959 2165 11962
rect 2217 11959 2233 11962
rect 2285 11959 2301 11962
rect 2353 11959 2369 11962
rect 2421 11959 2437 11962
rect 2489 11959 2505 11962
rect 2557 11959 2573 11962
rect 2625 11959 2641 11962
rect 2693 11959 2695 12011
rect 2095 10813 2695 11959
rect 2095 10761 2097 10813
rect 2149 10810 2165 10813
rect 2217 10810 2233 10813
rect 2285 10810 2301 10813
rect 2353 10810 2369 10813
rect 2421 10810 2437 10813
rect 2489 10810 2505 10813
rect 2557 10810 2573 10813
rect 2625 10810 2641 10813
rect 2693 10761 2695 10813
rect 2095 10749 2127 10761
rect 2663 10749 2695 10761
rect 2095 10697 2097 10749
rect 2693 10697 2695 10749
rect 2095 10685 2127 10697
rect 2663 10685 2695 10697
rect 2095 10633 2097 10685
rect 2693 10633 2695 10685
rect 2095 10621 2127 10633
rect 2663 10621 2695 10633
rect 2095 10569 2097 10621
rect 2693 10569 2695 10621
rect 2095 10557 2127 10569
rect 2663 10557 2695 10569
rect 2095 10505 2097 10557
rect 2693 10505 2695 10557
rect 2095 10493 2127 10505
rect 2663 10493 2695 10505
rect 2095 10441 2097 10493
rect 2693 10441 2695 10493
rect 2095 10429 2127 10441
rect 2663 10429 2695 10441
rect 2095 10377 2097 10429
rect 2693 10377 2695 10429
rect 2095 10365 2127 10377
rect 2663 10365 2695 10377
rect 2095 10313 2097 10365
rect 2149 10329 2165 10354
rect 2217 10329 2233 10354
rect 2285 10329 2301 10354
rect 2353 10329 2369 10354
rect 2421 10329 2437 10354
rect 2489 10329 2505 10354
rect 2557 10329 2573 10354
rect 2625 10329 2641 10354
rect 2285 10313 2287 10329
rect 2353 10313 2367 10329
rect 2423 10313 2437 10329
rect 2503 10313 2505 10329
rect 2693 10313 2695 10365
rect 2095 10301 2127 10313
rect 2183 10301 2207 10313
rect 2263 10301 2287 10313
rect 2343 10301 2367 10313
rect 2423 10301 2447 10313
rect 2503 10301 2527 10313
rect 2583 10301 2607 10313
rect 2663 10301 2695 10313
rect 2095 10249 2097 10301
rect 2285 10273 2287 10301
rect 2353 10273 2367 10301
rect 2423 10273 2437 10301
rect 2503 10273 2505 10301
rect 2149 10249 2165 10273
rect 2217 10249 2233 10273
rect 2285 10249 2301 10273
rect 2353 10249 2369 10273
rect 2421 10249 2437 10273
rect 2489 10249 2505 10273
rect 2557 10249 2573 10273
rect 2625 10249 2641 10273
rect 2693 10249 2695 10301
rect 2095 10248 2695 10249
rect 2095 10237 2127 10248
rect 2183 10237 2207 10248
rect 2263 10237 2287 10248
rect 2343 10237 2367 10248
rect 2423 10237 2447 10248
rect 2503 10237 2527 10248
rect 2583 10237 2607 10248
rect 2663 10237 2695 10248
rect 2095 10185 2097 10237
rect 2285 10192 2287 10237
rect 2353 10192 2367 10237
rect 2423 10192 2437 10237
rect 2503 10192 2505 10237
rect 2149 10185 2165 10192
rect 2217 10185 2233 10192
rect 2285 10185 2301 10192
rect 2353 10185 2369 10192
rect 2421 10185 2437 10192
rect 2489 10185 2505 10192
rect 2557 10185 2573 10192
rect 2625 10185 2641 10192
rect 2693 10185 2695 10237
rect 2095 10173 2695 10185
rect 2095 10121 2097 10173
rect 2149 10167 2165 10173
rect 2217 10167 2233 10173
rect 2285 10167 2301 10173
rect 2353 10167 2369 10173
rect 2421 10167 2437 10173
rect 2489 10167 2505 10173
rect 2557 10167 2573 10173
rect 2625 10167 2641 10173
rect 2285 10121 2287 10167
rect 2353 10121 2367 10167
rect 2423 10121 2437 10167
rect 2503 10121 2505 10167
rect 2693 10121 2695 10173
rect 2095 10111 2127 10121
rect 2183 10111 2207 10121
rect 2263 10111 2287 10121
rect 2343 10111 2367 10121
rect 2423 10111 2447 10121
rect 2503 10111 2527 10121
rect 2583 10111 2607 10121
rect 2663 10111 2695 10121
rect 2095 10109 2695 10111
rect 2095 10057 2097 10109
rect 2149 10086 2165 10109
rect 2217 10086 2233 10109
rect 2285 10086 2301 10109
rect 2353 10086 2369 10109
rect 2421 10086 2437 10109
rect 2489 10086 2505 10109
rect 2557 10086 2573 10109
rect 2625 10086 2641 10109
rect 2285 10057 2287 10086
rect 2353 10057 2367 10086
rect 2423 10057 2437 10086
rect 2503 10057 2505 10086
rect 2693 10057 2695 10109
rect 2095 10045 2127 10057
rect 2183 10045 2207 10057
rect 2263 10045 2287 10057
rect 2343 10045 2367 10057
rect 2423 10045 2447 10057
rect 2503 10045 2527 10057
rect 2583 10045 2607 10057
rect 2663 10045 2695 10057
rect 2095 9993 2097 10045
rect 2285 10030 2287 10045
rect 2353 10030 2367 10045
rect 2423 10030 2437 10045
rect 2503 10030 2505 10045
rect 2149 10005 2165 10030
rect 2217 10005 2233 10030
rect 2285 10005 2301 10030
rect 2353 10005 2369 10030
rect 2421 10005 2437 10030
rect 2489 10005 2505 10030
rect 2557 10005 2573 10030
rect 2625 10005 2641 10030
rect 2285 9993 2287 10005
rect 2353 9993 2367 10005
rect 2423 9993 2437 10005
rect 2503 9993 2505 10005
rect 2693 9993 2695 10045
rect 2095 9981 2127 9993
rect 2183 9981 2207 9993
rect 2263 9981 2287 9993
rect 2343 9981 2367 9993
rect 2423 9981 2447 9993
rect 2503 9981 2527 9993
rect 2583 9981 2607 9993
rect 2663 9981 2695 9993
rect 2095 9929 2097 9981
rect 2285 9949 2287 9981
rect 2353 9949 2367 9981
rect 2423 9949 2437 9981
rect 2503 9949 2505 9981
rect 2149 9929 2165 9949
rect 2217 9929 2233 9949
rect 2285 9929 2301 9949
rect 2353 9929 2369 9949
rect 2421 9929 2437 9949
rect 2489 9929 2505 9949
rect 2557 9929 2573 9949
rect 2625 9929 2641 9949
rect 2693 9929 2695 9981
rect 2095 9924 2695 9929
rect 2095 9917 2127 9924
rect 2183 9917 2207 9924
rect 2263 9917 2287 9924
rect 2343 9917 2367 9924
rect 2423 9917 2447 9924
rect 2503 9917 2527 9924
rect 2583 9917 2607 9924
rect 2663 9917 2695 9924
rect 2095 9865 2097 9917
rect 2285 9868 2287 9917
rect 2353 9868 2367 9917
rect 2423 9868 2437 9917
rect 2503 9868 2505 9917
rect 2149 9865 2165 9868
rect 2217 9865 2233 9868
rect 2285 9865 2301 9868
rect 2353 9865 2369 9868
rect 2421 9865 2437 9868
rect 2489 9865 2505 9868
rect 2557 9865 2573 9868
rect 2625 9865 2641 9868
rect 2693 9865 2695 9917
rect 2095 8611 2695 9865
rect 2095 8559 2097 8611
rect 2149 8608 2165 8611
rect 2217 8608 2233 8611
rect 2285 8608 2301 8611
rect 2353 8608 2369 8611
rect 2421 8608 2437 8611
rect 2489 8608 2505 8611
rect 2557 8608 2573 8611
rect 2625 8608 2641 8611
rect 2693 8559 2695 8611
rect 2095 8547 2127 8559
rect 2663 8547 2695 8559
rect 2095 8495 2097 8547
rect 2693 8495 2695 8547
rect 2095 8483 2127 8495
rect 2663 8483 2695 8495
rect 2095 8431 2097 8483
rect 2693 8431 2695 8483
rect 2095 8419 2127 8431
rect 2663 8419 2695 8431
rect 2095 8367 2097 8419
rect 2693 8367 2695 8419
rect 2095 8355 2127 8367
rect 2663 8355 2695 8367
rect 2095 8303 2097 8355
rect 2693 8303 2695 8355
rect 2095 8291 2127 8303
rect 2663 8291 2695 8303
rect 2095 8239 2097 8291
rect 2693 8239 2695 8291
rect 2095 8227 2127 8239
rect 2663 8227 2695 8239
rect 2095 8175 2097 8227
rect 2693 8175 2695 8227
rect 2095 8163 2127 8175
rect 2663 8163 2695 8175
rect 2095 8111 2097 8163
rect 2149 8127 2165 8152
rect 2217 8127 2233 8152
rect 2285 8127 2301 8152
rect 2353 8127 2369 8152
rect 2421 8127 2437 8152
rect 2489 8127 2505 8152
rect 2557 8127 2573 8152
rect 2625 8127 2641 8152
rect 2285 8111 2287 8127
rect 2353 8111 2367 8127
rect 2423 8111 2437 8127
rect 2503 8111 2505 8127
rect 2693 8111 2695 8163
rect 2095 8099 2127 8111
rect 2183 8099 2207 8111
rect 2263 8099 2287 8111
rect 2343 8099 2367 8111
rect 2423 8099 2447 8111
rect 2503 8099 2527 8111
rect 2583 8099 2607 8111
rect 2663 8099 2695 8111
rect 2095 8047 2097 8099
rect 2285 8071 2287 8099
rect 2353 8071 2367 8099
rect 2423 8071 2437 8099
rect 2503 8071 2505 8099
rect 2149 8047 2165 8071
rect 2217 8047 2233 8071
rect 2285 8047 2301 8071
rect 2353 8047 2369 8071
rect 2421 8047 2437 8071
rect 2489 8047 2505 8071
rect 2557 8047 2573 8071
rect 2625 8047 2641 8071
rect 2693 8047 2695 8099
rect 2095 8046 2695 8047
rect 2095 8035 2127 8046
rect 2183 8035 2207 8046
rect 2263 8035 2287 8046
rect 2343 8035 2367 8046
rect 2423 8035 2447 8046
rect 2503 8035 2527 8046
rect 2583 8035 2607 8046
rect 2663 8035 2695 8046
rect 2095 7983 2097 8035
rect 2285 7990 2287 8035
rect 2353 7990 2367 8035
rect 2423 7990 2437 8035
rect 2503 7990 2505 8035
rect 2149 7983 2165 7990
rect 2217 7983 2233 7990
rect 2285 7983 2301 7990
rect 2353 7983 2369 7990
rect 2421 7983 2437 7990
rect 2489 7983 2505 7990
rect 2557 7983 2573 7990
rect 2625 7983 2641 7990
rect 2693 7983 2695 8035
rect 2095 7971 2695 7983
rect 2095 7919 2097 7971
rect 2149 7965 2165 7971
rect 2217 7965 2233 7971
rect 2285 7965 2301 7971
rect 2353 7965 2369 7971
rect 2421 7965 2437 7971
rect 2489 7965 2505 7971
rect 2557 7965 2573 7971
rect 2625 7965 2641 7971
rect 2285 7919 2287 7965
rect 2353 7919 2367 7965
rect 2423 7919 2437 7965
rect 2503 7919 2505 7965
rect 2693 7919 2695 7971
rect 2095 7909 2127 7919
rect 2183 7909 2207 7919
rect 2263 7909 2287 7919
rect 2343 7909 2367 7919
rect 2423 7909 2447 7919
rect 2503 7909 2527 7919
rect 2583 7909 2607 7919
rect 2663 7909 2695 7919
rect 2095 7907 2695 7909
rect 2095 7855 2097 7907
rect 2149 7884 2165 7907
rect 2217 7884 2233 7907
rect 2285 7884 2301 7907
rect 2353 7884 2369 7907
rect 2421 7884 2437 7907
rect 2489 7884 2505 7907
rect 2557 7884 2573 7907
rect 2625 7884 2641 7907
rect 2285 7855 2287 7884
rect 2353 7855 2367 7884
rect 2423 7855 2437 7884
rect 2503 7855 2505 7884
rect 2693 7855 2695 7907
rect 2095 7843 2127 7855
rect 2183 7843 2207 7855
rect 2263 7843 2287 7855
rect 2343 7843 2367 7855
rect 2423 7843 2447 7855
rect 2503 7843 2527 7855
rect 2583 7843 2607 7855
rect 2663 7843 2695 7855
rect 2095 7791 2097 7843
rect 2285 7828 2287 7843
rect 2353 7828 2367 7843
rect 2423 7828 2437 7843
rect 2503 7828 2505 7843
rect 2149 7803 2165 7828
rect 2217 7803 2233 7828
rect 2285 7803 2301 7828
rect 2353 7803 2369 7828
rect 2421 7803 2437 7828
rect 2489 7803 2505 7828
rect 2557 7803 2573 7828
rect 2625 7803 2641 7828
rect 2285 7791 2287 7803
rect 2353 7791 2367 7803
rect 2423 7791 2437 7803
rect 2503 7791 2505 7803
rect 2693 7791 2695 7843
rect 2095 7779 2127 7791
rect 2183 7779 2207 7791
rect 2263 7779 2287 7791
rect 2343 7779 2367 7791
rect 2423 7779 2447 7791
rect 2503 7779 2527 7791
rect 2583 7779 2607 7791
rect 2663 7779 2695 7791
rect 2095 7727 2097 7779
rect 2285 7747 2287 7779
rect 2353 7747 2367 7779
rect 2423 7747 2437 7779
rect 2503 7747 2505 7779
rect 2149 7727 2165 7747
rect 2217 7727 2233 7747
rect 2285 7727 2301 7747
rect 2353 7727 2369 7747
rect 2421 7727 2437 7747
rect 2489 7727 2505 7747
rect 2557 7727 2573 7747
rect 2625 7727 2641 7747
rect 2693 7727 2695 7779
rect 2095 7722 2695 7727
rect 2095 7715 2127 7722
rect 2183 7715 2207 7722
rect 2263 7715 2287 7722
rect 2343 7715 2367 7722
rect 2423 7715 2447 7722
rect 2503 7715 2527 7722
rect 2583 7715 2607 7722
rect 2663 7715 2695 7722
rect 2095 7663 2097 7715
rect 2285 7666 2287 7715
rect 2353 7666 2367 7715
rect 2423 7666 2437 7715
rect 2503 7666 2505 7715
rect 2149 7663 2165 7666
rect 2217 7663 2233 7666
rect 2285 7663 2301 7666
rect 2353 7663 2369 7666
rect 2421 7663 2437 7666
rect 2489 7663 2505 7666
rect 2557 7663 2573 7666
rect 2625 7663 2641 7666
rect 2693 7663 2695 7715
rect 2095 6501 2695 7663
rect 2095 6449 2097 6501
rect 2149 6498 2165 6501
rect 2217 6498 2233 6501
rect 2285 6498 2301 6501
rect 2353 6498 2369 6501
rect 2421 6498 2437 6501
rect 2489 6498 2505 6501
rect 2557 6498 2573 6501
rect 2625 6498 2641 6501
rect 2693 6449 2695 6501
rect 2095 6437 2127 6449
rect 2663 6437 2695 6449
rect 2095 6385 2097 6437
rect 2693 6385 2695 6437
rect 2095 6373 2127 6385
rect 2663 6373 2695 6385
rect 2095 6321 2097 6373
rect 2693 6321 2695 6373
rect 2095 6309 2127 6321
rect 2663 6309 2695 6321
rect 2095 6257 2097 6309
rect 2693 6257 2695 6309
rect 2095 6245 2127 6257
rect 2663 6245 2695 6257
rect 2095 6193 2097 6245
rect 2693 6193 2695 6245
rect 2095 6181 2127 6193
rect 2663 6181 2695 6193
rect 2095 6129 2097 6181
rect 2693 6129 2695 6181
rect 2095 6117 2127 6129
rect 2663 6117 2695 6129
rect 2095 6065 2097 6117
rect 2693 6065 2695 6117
rect 2095 6053 2127 6065
rect 2663 6053 2695 6065
rect 2095 6001 2097 6053
rect 2149 6017 2165 6042
rect 2217 6017 2233 6042
rect 2285 6017 2301 6042
rect 2353 6017 2369 6042
rect 2421 6017 2437 6042
rect 2489 6017 2505 6042
rect 2557 6017 2573 6042
rect 2625 6017 2641 6042
rect 2285 6001 2287 6017
rect 2353 6001 2367 6017
rect 2423 6001 2437 6017
rect 2503 6001 2505 6017
rect 2693 6001 2695 6053
rect 2095 5989 2127 6001
rect 2183 5989 2207 6001
rect 2263 5989 2287 6001
rect 2343 5989 2367 6001
rect 2423 5989 2447 6001
rect 2503 5989 2527 6001
rect 2583 5989 2607 6001
rect 2663 5989 2695 6001
rect 2095 5937 2097 5989
rect 2285 5961 2287 5989
rect 2353 5961 2367 5989
rect 2423 5961 2437 5989
rect 2503 5961 2505 5989
rect 2149 5937 2165 5961
rect 2217 5937 2233 5961
rect 2285 5937 2301 5961
rect 2353 5937 2369 5961
rect 2421 5937 2437 5961
rect 2489 5937 2505 5961
rect 2557 5937 2573 5961
rect 2625 5937 2641 5961
rect 2693 5937 2695 5989
rect 2095 5936 2695 5937
rect 2095 5925 2127 5936
rect 2183 5925 2207 5936
rect 2263 5925 2287 5936
rect 2343 5925 2367 5936
rect 2423 5925 2447 5936
rect 2503 5925 2527 5936
rect 2583 5925 2607 5936
rect 2663 5925 2695 5936
rect 2095 5873 2097 5925
rect 2285 5880 2287 5925
rect 2353 5880 2367 5925
rect 2423 5880 2437 5925
rect 2503 5880 2505 5925
rect 2149 5873 2165 5880
rect 2217 5873 2233 5880
rect 2285 5873 2301 5880
rect 2353 5873 2369 5880
rect 2421 5873 2437 5880
rect 2489 5873 2505 5880
rect 2557 5873 2573 5880
rect 2625 5873 2641 5880
rect 2693 5873 2695 5925
rect 2095 5861 2695 5873
rect 2095 5809 2097 5861
rect 2149 5855 2165 5861
rect 2217 5855 2233 5861
rect 2285 5855 2301 5861
rect 2353 5855 2369 5861
rect 2421 5855 2437 5861
rect 2489 5855 2505 5861
rect 2557 5855 2573 5861
rect 2625 5855 2641 5861
rect 2285 5809 2287 5855
rect 2353 5809 2367 5855
rect 2423 5809 2437 5855
rect 2503 5809 2505 5855
rect 2693 5809 2695 5861
rect 2095 5799 2127 5809
rect 2183 5799 2207 5809
rect 2263 5799 2287 5809
rect 2343 5799 2367 5809
rect 2423 5799 2447 5809
rect 2503 5799 2527 5809
rect 2583 5799 2607 5809
rect 2663 5799 2695 5809
rect 2095 5797 2695 5799
rect 2095 5745 2097 5797
rect 2149 5774 2165 5797
rect 2217 5774 2233 5797
rect 2285 5774 2301 5797
rect 2353 5774 2369 5797
rect 2421 5774 2437 5797
rect 2489 5774 2505 5797
rect 2557 5774 2573 5797
rect 2625 5774 2641 5797
rect 2285 5745 2287 5774
rect 2353 5745 2367 5774
rect 2423 5745 2437 5774
rect 2503 5745 2505 5774
rect 2693 5745 2695 5797
rect 2095 5733 2127 5745
rect 2183 5733 2207 5745
rect 2263 5733 2287 5745
rect 2343 5733 2367 5745
rect 2423 5733 2447 5745
rect 2503 5733 2527 5745
rect 2583 5733 2607 5745
rect 2663 5733 2695 5745
rect 2095 5681 2097 5733
rect 2285 5718 2287 5733
rect 2353 5718 2367 5733
rect 2423 5718 2437 5733
rect 2503 5718 2505 5733
rect 2149 5693 2165 5718
rect 2217 5693 2233 5718
rect 2285 5693 2301 5718
rect 2353 5693 2369 5718
rect 2421 5693 2437 5718
rect 2489 5693 2505 5718
rect 2557 5693 2573 5718
rect 2625 5693 2641 5718
rect 2285 5681 2287 5693
rect 2353 5681 2367 5693
rect 2423 5681 2437 5693
rect 2503 5681 2505 5693
rect 2693 5681 2695 5733
rect 2095 5669 2127 5681
rect 2183 5669 2207 5681
rect 2263 5669 2287 5681
rect 2343 5669 2367 5681
rect 2423 5669 2447 5681
rect 2503 5669 2527 5681
rect 2583 5669 2607 5681
rect 2663 5669 2695 5681
rect 2095 5617 2097 5669
rect 2285 5637 2287 5669
rect 2353 5637 2367 5669
rect 2423 5637 2437 5669
rect 2503 5637 2505 5669
rect 2149 5617 2165 5637
rect 2217 5617 2233 5637
rect 2285 5617 2301 5637
rect 2353 5617 2369 5637
rect 2421 5617 2437 5637
rect 2489 5617 2505 5637
rect 2557 5617 2573 5637
rect 2625 5617 2641 5637
rect 2693 5617 2695 5669
rect 2095 5612 2695 5617
rect 2095 5605 2127 5612
rect 2183 5605 2207 5612
rect 2263 5605 2287 5612
rect 2343 5605 2367 5612
rect 2423 5605 2447 5612
rect 2503 5605 2527 5612
rect 2583 5605 2607 5612
rect 2663 5605 2695 5612
rect 2095 5553 2097 5605
rect 2285 5556 2287 5605
rect 2353 5556 2367 5605
rect 2423 5556 2437 5605
rect 2503 5556 2505 5605
rect 2149 5553 2165 5556
rect 2217 5553 2233 5556
rect 2285 5553 2301 5556
rect 2353 5553 2369 5556
rect 2421 5553 2437 5556
rect 2489 5553 2505 5556
rect 2557 5553 2573 5556
rect 2625 5553 2641 5556
rect 2693 5553 2695 5605
rect 2095 4437 2695 5553
rect 2095 4385 2097 4437
rect 2149 4434 2165 4437
rect 2217 4434 2233 4437
rect 2285 4434 2301 4437
rect 2353 4434 2369 4437
rect 2421 4434 2437 4437
rect 2489 4434 2505 4437
rect 2557 4434 2573 4437
rect 2625 4434 2641 4437
rect 2693 4385 2695 4437
rect 2095 4373 2127 4385
rect 2663 4373 2695 4385
rect 2095 4321 2097 4373
rect 2693 4321 2695 4373
rect 2095 4309 2127 4321
rect 2663 4309 2695 4321
rect 2095 4257 2097 4309
rect 2693 4257 2695 4309
rect 2095 4245 2127 4257
rect 2663 4245 2695 4257
rect 2095 4193 2097 4245
rect 2693 4193 2695 4245
rect 2095 4181 2127 4193
rect 2663 4181 2695 4193
rect 2095 4129 2097 4181
rect 2693 4129 2695 4181
rect 2095 4117 2127 4129
rect 2663 4117 2695 4129
rect 2095 4065 2097 4117
rect 2693 4065 2695 4117
rect 2095 4053 2127 4065
rect 2663 4053 2695 4065
rect 2095 4001 2097 4053
rect 2693 4001 2695 4053
rect 2095 3989 2127 4001
rect 2663 3989 2695 4001
rect 2095 3937 2097 3989
rect 2149 3953 2165 3978
rect 2217 3953 2233 3978
rect 2285 3953 2301 3978
rect 2353 3953 2369 3978
rect 2421 3953 2437 3978
rect 2489 3953 2505 3978
rect 2557 3953 2573 3978
rect 2625 3953 2641 3978
rect 2285 3937 2287 3953
rect 2353 3937 2367 3953
rect 2423 3937 2437 3953
rect 2503 3937 2505 3953
rect 2693 3937 2695 3989
rect 2095 3925 2127 3937
rect 2183 3925 2207 3937
rect 2263 3925 2287 3937
rect 2343 3925 2367 3937
rect 2423 3925 2447 3937
rect 2503 3925 2527 3937
rect 2583 3925 2607 3937
rect 2663 3925 2695 3937
rect 2095 3873 2097 3925
rect 2285 3897 2287 3925
rect 2353 3897 2367 3925
rect 2423 3897 2437 3925
rect 2503 3897 2505 3925
rect 2149 3873 2165 3897
rect 2217 3873 2233 3897
rect 2285 3873 2301 3897
rect 2353 3873 2369 3897
rect 2421 3873 2437 3897
rect 2489 3873 2505 3897
rect 2557 3873 2573 3897
rect 2625 3873 2641 3897
rect 2693 3873 2695 3925
rect 2095 3872 2695 3873
rect 2095 3861 2127 3872
rect 2183 3861 2207 3872
rect 2263 3861 2287 3872
rect 2343 3861 2367 3872
rect 2423 3861 2447 3872
rect 2503 3861 2527 3872
rect 2583 3861 2607 3872
rect 2663 3861 2695 3872
rect 2095 3809 2097 3861
rect 2285 3816 2287 3861
rect 2353 3816 2367 3861
rect 2423 3816 2437 3861
rect 2503 3816 2505 3861
rect 2149 3809 2165 3816
rect 2217 3809 2233 3816
rect 2285 3809 2301 3816
rect 2353 3809 2369 3816
rect 2421 3809 2437 3816
rect 2489 3809 2505 3816
rect 2557 3809 2573 3816
rect 2625 3809 2641 3816
rect 2693 3809 2695 3861
rect 2095 3797 2695 3809
rect 2095 3745 2097 3797
rect 2149 3791 2165 3797
rect 2217 3791 2233 3797
rect 2285 3791 2301 3797
rect 2353 3791 2369 3797
rect 2421 3791 2437 3797
rect 2489 3791 2505 3797
rect 2557 3791 2573 3797
rect 2625 3791 2641 3797
rect 2285 3745 2287 3791
rect 2353 3745 2367 3791
rect 2423 3745 2437 3791
rect 2503 3745 2505 3791
rect 2693 3745 2695 3797
rect 2095 3735 2127 3745
rect 2183 3735 2207 3745
rect 2263 3735 2287 3745
rect 2343 3735 2367 3745
rect 2423 3735 2447 3745
rect 2503 3735 2527 3745
rect 2583 3735 2607 3745
rect 2663 3735 2695 3745
rect 2095 3733 2695 3735
rect 2095 3681 2097 3733
rect 2149 3710 2165 3733
rect 2217 3710 2233 3733
rect 2285 3710 2301 3733
rect 2353 3710 2369 3733
rect 2421 3710 2437 3733
rect 2489 3710 2505 3733
rect 2557 3710 2573 3733
rect 2625 3710 2641 3733
rect 2285 3681 2287 3710
rect 2353 3681 2367 3710
rect 2423 3681 2437 3710
rect 2503 3681 2505 3710
rect 2693 3681 2695 3733
rect 2095 3669 2127 3681
rect 2183 3669 2207 3681
rect 2263 3669 2287 3681
rect 2343 3669 2367 3681
rect 2423 3669 2447 3681
rect 2503 3669 2527 3681
rect 2583 3669 2607 3681
rect 2663 3669 2695 3681
rect 2095 3617 2097 3669
rect 2285 3654 2287 3669
rect 2353 3654 2367 3669
rect 2423 3654 2437 3669
rect 2503 3654 2505 3669
rect 2149 3629 2165 3654
rect 2217 3629 2233 3654
rect 2285 3629 2301 3654
rect 2353 3629 2369 3654
rect 2421 3629 2437 3654
rect 2489 3629 2505 3654
rect 2557 3629 2573 3654
rect 2625 3629 2641 3654
rect 2285 3617 2287 3629
rect 2353 3617 2367 3629
rect 2423 3617 2437 3629
rect 2503 3617 2505 3629
rect 2693 3617 2695 3669
rect 2095 3605 2127 3617
rect 2183 3605 2207 3617
rect 2263 3605 2287 3617
rect 2343 3605 2367 3617
rect 2423 3605 2447 3617
rect 2503 3605 2527 3617
rect 2583 3605 2607 3617
rect 2663 3605 2695 3617
rect 2095 3553 2097 3605
rect 2285 3573 2287 3605
rect 2353 3573 2367 3605
rect 2423 3573 2437 3605
rect 2503 3573 2505 3605
rect 2149 3553 2165 3573
rect 2217 3553 2233 3573
rect 2285 3553 2301 3573
rect 2353 3553 2369 3573
rect 2421 3553 2437 3573
rect 2489 3553 2505 3573
rect 2557 3553 2573 3573
rect 2625 3553 2641 3573
rect 2693 3553 2695 3605
rect 2095 3548 2695 3553
rect 2095 3541 2127 3548
rect 2183 3541 2207 3548
rect 2263 3541 2287 3548
rect 2343 3541 2367 3548
rect 2423 3541 2447 3548
rect 2503 3541 2527 3548
rect 2583 3541 2607 3548
rect 2663 3541 2695 3548
rect 2095 3489 2097 3541
rect 2285 3492 2287 3541
rect 2353 3492 2367 3541
rect 2423 3492 2437 3541
rect 2503 3492 2505 3541
rect 2149 3489 2165 3492
rect 2217 3489 2233 3492
rect 2285 3489 2301 3492
rect 2353 3489 2369 3492
rect 2421 3489 2437 3492
rect 2489 3489 2505 3492
rect 2557 3489 2573 3492
rect 2625 3489 2641 3492
rect 2693 3489 2695 3541
rect 2095 2243 2695 3489
rect 2095 2191 2097 2243
rect 2149 2240 2165 2243
rect 2217 2240 2233 2243
rect 2285 2240 2301 2243
rect 2353 2240 2369 2243
rect 2421 2240 2437 2243
rect 2489 2240 2505 2243
rect 2557 2240 2573 2243
rect 2625 2240 2641 2243
rect 2693 2191 2695 2243
rect 2095 2179 2127 2191
rect 2663 2179 2695 2191
rect 2095 2127 2097 2179
rect 2693 2127 2695 2179
rect 2095 2115 2127 2127
rect 2663 2115 2695 2127
rect 2095 2063 2097 2115
rect 2693 2063 2695 2115
rect 2095 2051 2127 2063
rect 2663 2051 2695 2063
rect 2095 1999 2097 2051
rect 2693 1999 2695 2051
rect 2095 1987 2127 1999
rect 2663 1987 2695 1999
rect 2095 1935 2097 1987
rect 2693 1935 2695 1987
rect 2095 1923 2127 1935
rect 2663 1923 2695 1935
rect 2095 1871 2097 1923
rect 2693 1871 2695 1923
rect 2095 1859 2127 1871
rect 2663 1859 2695 1871
rect 2095 1807 2097 1859
rect 2693 1807 2695 1859
rect 2095 1795 2127 1807
rect 2663 1795 2695 1807
rect 2095 1743 2097 1795
rect 2149 1759 2165 1784
rect 2217 1759 2233 1784
rect 2285 1759 2301 1784
rect 2353 1759 2369 1784
rect 2421 1759 2437 1784
rect 2489 1759 2505 1784
rect 2557 1759 2573 1784
rect 2625 1759 2641 1784
rect 2285 1743 2287 1759
rect 2353 1743 2367 1759
rect 2423 1743 2437 1759
rect 2503 1743 2505 1759
rect 2693 1743 2695 1795
rect 2095 1731 2127 1743
rect 2183 1731 2207 1743
rect 2263 1731 2287 1743
rect 2343 1731 2367 1743
rect 2423 1731 2447 1743
rect 2503 1731 2527 1743
rect 2583 1731 2607 1743
rect 2663 1731 2695 1743
rect 2095 1679 2097 1731
rect 2285 1703 2287 1731
rect 2353 1703 2367 1731
rect 2423 1703 2437 1731
rect 2503 1703 2505 1731
rect 2149 1679 2165 1703
rect 2217 1679 2233 1703
rect 2285 1679 2301 1703
rect 2353 1679 2369 1703
rect 2421 1679 2437 1703
rect 2489 1679 2505 1703
rect 2557 1679 2573 1703
rect 2625 1679 2641 1703
rect 2693 1679 2695 1731
rect 2095 1678 2695 1679
rect 2095 1667 2127 1678
rect 2183 1667 2207 1678
rect 2263 1667 2287 1678
rect 2343 1667 2367 1678
rect 2423 1667 2447 1678
rect 2503 1667 2527 1678
rect 2583 1667 2607 1678
rect 2663 1667 2695 1678
rect 2095 1615 2097 1667
rect 2285 1622 2287 1667
rect 2353 1622 2367 1667
rect 2423 1622 2437 1667
rect 2503 1622 2505 1667
rect 2149 1615 2165 1622
rect 2217 1615 2233 1622
rect 2285 1615 2301 1622
rect 2353 1615 2369 1622
rect 2421 1615 2437 1622
rect 2489 1615 2505 1622
rect 2557 1615 2573 1622
rect 2625 1615 2641 1622
rect 2693 1615 2695 1667
rect 2095 1603 2695 1615
rect 2095 1551 2097 1603
rect 2149 1597 2165 1603
rect 2217 1597 2233 1603
rect 2285 1597 2301 1603
rect 2353 1597 2369 1603
rect 2421 1597 2437 1603
rect 2489 1597 2505 1603
rect 2557 1597 2573 1603
rect 2625 1597 2641 1603
rect 2285 1551 2287 1597
rect 2353 1551 2367 1597
rect 2423 1551 2437 1597
rect 2503 1551 2505 1597
rect 2693 1551 2695 1603
rect 2095 1541 2127 1551
rect 2183 1541 2207 1551
rect 2263 1541 2287 1551
rect 2343 1541 2367 1551
rect 2423 1541 2447 1551
rect 2503 1541 2527 1551
rect 2583 1541 2607 1551
rect 2663 1541 2695 1551
rect 2095 1539 2695 1541
rect 2095 1487 2097 1539
rect 2149 1516 2165 1539
rect 2217 1516 2233 1539
rect 2285 1516 2301 1539
rect 2353 1516 2369 1539
rect 2421 1516 2437 1539
rect 2489 1516 2505 1539
rect 2557 1516 2573 1539
rect 2625 1516 2641 1539
rect 2285 1487 2287 1516
rect 2353 1487 2367 1516
rect 2423 1487 2437 1516
rect 2503 1487 2505 1516
rect 2693 1487 2695 1539
rect 2095 1475 2127 1487
rect 2183 1475 2207 1487
rect 2263 1475 2287 1487
rect 2343 1475 2367 1487
rect 2423 1475 2447 1487
rect 2503 1475 2527 1487
rect 2583 1475 2607 1487
rect 2663 1475 2695 1487
rect 2095 1423 2097 1475
rect 2285 1460 2287 1475
rect 2353 1460 2367 1475
rect 2423 1460 2437 1475
rect 2503 1460 2505 1475
rect 2149 1435 2165 1460
rect 2217 1435 2233 1460
rect 2285 1435 2301 1460
rect 2353 1435 2369 1460
rect 2421 1435 2437 1460
rect 2489 1435 2505 1460
rect 2557 1435 2573 1460
rect 2625 1435 2641 1460
rect 2285 1423 2287 1435
rect 2353 1423 2367 1435
rect 2423 1423 2437 1435
rect 2503 1423 2505 1435
rect 2693 1423 2695 1475
rect 2095 1411 2127 1423
rect 2183 1411 2207 1423
rect 2263 1411 2287 1423
rect 2343 1411 2367 1423
rect 2423 1411 2447 1423
rect 2503 1411 2527 1423
rect 2583 1411 2607 1423
rect 2663 1411 2695 1423
rect 2095 1359 2097 1411
rect 2285 1379 2287 1411
rect 2353 1379 2367 1411
rect 2423 1379 2437 1411
rect 2503 1379 2505 1411
rect 2149 1359 2165 1379
rect 2217 1359 2233 1379
rect 2285 1359 2301 1379
rect 2353 1359 2369 1379
rect 2421 1359 2437 1379
rect 2489 1359 2505 1379
rect 2557 1359 2573 1379
rect 2625 1359 2641 1379
rect 2693 1359 2695 1411
rect 2095 1354 2695 1359
rect 2095 1347 2127 1354
rect 2183 1347 2207 1354
rect 2263 1347 2287 1354
rect 2343 1347 2367 1354
rect 2423 1347 2447 1354
rect 2503 1347 2527 1354
rect 2583 1347 2607 1354
rect 2663 1347 2695 1354
rect 2095 1295 2097 1347
rect 2285 1298 2287 1347
rect 2353 1298 2367 1347
rect 2423 1298 2437 1347
rect 2503 1298 2505 1347
rect 2149 1295 2165 1298
rect 2217 1295 2233 1298
rect 2285 1295 2301 1298
rect 2353 1295 2369 1298
rect 2421 1295 2437 1298
rect 2489 1295 2505 1298
rect 2557 1295 2573 1298
rect 2625 1295 2641 1298
rect 2693 1295 2695 1347
rect 2095 141 2695 1295
rect 2095 85 2104 141
rect 2160 85 2192 141
rect 2248 85 2280 141
rect 2336 85 2368 141
rect 2424 85 2456 141
rect 2512 85 2543 141
rect 2599 85 2630 141
rect 2686 85 2695 141
rect 2095 61 2695 85
rect 2095 5 2104 61
rect 2160 5 2192 61
rect 2248 5 2280 61
rect 2336 5 2368 61
rect 2424 5 2456 61
rect 2512 5 2543 61
rect 2599 5 2630 61
rect 2686 5 2695 61
rect 2095 0 2695 5
<< via2 >>
rect 727 38371 749 38420
rect 749 38371 765 38420
rect 765 38371 817 38420
rect 817 38371 833 38420
rect 833 38371 885 38420
rect 885 38371 901 38420
rect 901 38371 953 38420
rect 953 38371 969 38420
rect 969 38371 1021 38420
rect 1021 38371 1037 38420
rect 1037 38371 1089 38420
rect 1089 38371 1105 38420
rect 1105 38371 1157 38420
rect 1157 38371 1173 38420
rect 1173 38371 1225 38420
rect 1225 38371 1241 38420
rect 1241 38371 1263 38420
rect 727 38359 1263 38371
rect 727 38307 749 38359
rect 749 38307 765 38359
rect 765 38307 817 38359
rect 817 38307 833 38359
rect 833 38307 885 38359
rect 885 38307 901 38359
rect 901 38307 953 38359
rect 953 38307 969 38359
rect 969 38307 1021 38359
rect 1021 38307 1037 38359
rect 1037 38307 1089 38359
rect 1089 38307 1105 38359
rect 1105 38307 1157 38359
rect 1157 38307 1173 38359
rect 1173 38307 1225 38359
rect 1225 38307 1241 38359
rect 1241 38307 1263 38359
rect 727 38295 1263 38307
rect 727 38243 749 38295
rect 749 38243 765 38295
rect 765 38243 817 38295
rect 817 38243 833 38295
rect 833 38243 885 38295
rect 885 38243 901 38295
rect 901 38243 953 38295
rect 953 38243 969 38295
rect 969 38243 1021 38295
rect 1021 38243 1037 38295
rect 1037 38243 1089 38295
rect 1089 38243 1105 38295
rect 1105 38243 1157 38295
rect 1157 38243 1173 38295
rect 1173 38243 1225 38295
rect 1225 38243 1241 38295
rect 1241 38243 1263 38295
rect 727 38231 1263 38243
rect 727 38179 749 38231
rect 749 38179 765 38231
rect 765 38179 817 38231
rect 817 38179 833 38231
rect 833 38179 885 38231
rect 885 38179 901 38231
rect 901 38179 953 38231
rect 953 38179 969 38231
rect 969 38179 1021 38231
rect 1021 38179 1037 38231
rect 1037 38179 1089 38231
rect 1089 38179 1105 38231
rect 1105 38179 1157 38231
rect 1157 38179 1173 38231
rect 1173 38179 1225 38231
rect 1225 38179 1241 38231
rect 1241 38179 1263 38231
rect 727 38167 1263 38179
rect 727 38115 749 38167
rect 749 38115 765 38167
rect 765 38115 817 38167
rect 817 38115 833 38167
rect 833 38115 885 38167
rect 885 38115 901 38167
rect 901 38115 953 38167
rect 953 38115 969 38167
rect 969 38115 1021 38167
rect 1021 38115 1037 38167
rect 1037 38115 1089 38167
rect 1089 38115 1105 38167
rect 1105 38115 1157 38167
rect 1157 38115 1173 38167
rect 1173 38115 1225 38167
rect 1225 38115 1241 38167
rect 1241 38115 1263 38167
rect 727 38103 1263 38115
rect 727 38051 749 38103
rect 749 38051 765 38103
rect 765 38051 817 38103
rect 817 38051 833 38103
rect 833 38051 885 38103
rect 885 38051 901 38103
rect 901 38051 953 38103
rect 953 38051 969 38103
rect 969 38051 1021 38103
rect 1021 38051 1037 38103
rect 1037 38051 1089 38103
rect 1089 38051 1105 38103
rect 1105 38051 1157 38103
rect 1157 38051 1173 38103
rect 1173 38051 1225 38103
rect 1225 38051 1241 38103
rect 1241 38051 1263 38103
rect 727 38039 1263 38051
rect 727 37987 749 38039
rect 749 37987 765 38039
rect 765 37987 817 38039
rect 817 37987 833 38039
rect 833 37987 885 38039
rect 885 37987 901 38039
rect 901 37987 953 38039
rect 953 37987 969 38039
rect 969 37987 1021 38039
rect 1021 37987 1037 38039
rect 1037 37987 1089 38039
rect 1089 37987 1105 38039
rect 1105 37987 1157 38039
rect 1157 37987 1173 38039
rect 1173 37987 1225 38039
rect 1225 37987 1241 38039
rect 1241 37987 1263 38039
rect 727 37975 1263 37987
rect 727 37964 749 37975
rect 749 37964 765 37975
rect 765 37964 817 37975
rect 817 37964 833 37975
rect 833 37964 885 37975
rect 885 37964 901 37975
rect 901 37964 953 37975
rect 953 37964 969 37975
rect 969 37964 1021 37975
rect 1021 37964 1037 37975
rect 1037 37964 1089 37975
rect 1089 37964 1105 37975
rect 1105 37964 1157 37975
rect 1157 37964 1173 37975
rect 1173 37964 1225 37975
rect 1225 37964 1241 37975
rect 1241 37964 1263 37975
rect 727 37923 749 37939
rect 749 37923 765 37939
rect 765 37923 783 37939
rect 807 37923 817 37939
rect 817 37923 833 37939
rect 833 37923 863 37939
rect 887 37923 901 37939
rect 901 37923 943 37939
rect 967 37923 969 37939
rect 969 37923 1021 37939
rect 1021 37923 1023 37939
rect 1047 37923 1089 37939
rect 1089 37923 1103 37939
rect 1127 37923 1157 37939
rect 1157 37923 1173 37939
rect 1173 37923 1183 37939
rect 1207 37923 1225 37939
rect 1225 37923 1241 37939
rect 1241 37923 1263 37939
rect 727 37911 783 37923
rect 807 37911 863 37923
rect 887 37911 943 37923
rect 967 37911 1023 37923
rect 1047 37911 1103 37923
rect 1127 37911 1183 37923
rect 1207 37911 1263 37923
rect 727 37883 749 37911
rect 749 37883 765 37911
rect 765 37883 783 37911
rect 807 37883 817 37911
rect 817 37883 833 37911
rect 833 37883 863 37911
rect 887 37883 901 37911
rect 901 37883 943 37911
rect 967 37883 969 37911
rect 969 37883 1021 37911
rect 1021 37883 1023 37911
rect 1047 37883 1089 37911
rect 1089 37883 1103 37911
rect 1127 37883 1157 37911
rect 1157 37883 1173 37911
rect 1173 37883 1183 37911
rect 1207 37883 1225 37911
rect 1225 37883 1241 37911
rect 1241 37883 1263 37911
rect 727 37847 783 37858
rect 807 37847 863 37858
rect 887 37847 943 37858
rect 967 37847 1023 37858
rect 1047 37847 1103 37858
rect 1127 37847 1183 37858
rect 1207 37847 1263 37858
rect 727 37802 749 37847
rect 749 37802 765 37847
rect 765 37802 783 37847
rect 807 37802 817 37847
rect 817 37802 833 37847
rect 833 37802 863 37847
rect 887 37802 901 37847
rect 901 37802 943 37847
rect 967 37802 969 37847
rect 969 37802 1021 37847
rect 1021 37802 1023 37847
rect 1047 37802 1089 37847
rect 1089 37802 1103 37847
rect 1127 37802 1157 37847
rect 1157 37802 1173 37847
rect 1173 37802 1183 37847
rect 1207 37802 1225 37847
rect 1225 37802 1241 37847
rect 1241 37802 1263 37847
rect 727 37731 749 37777
rect 749 37731 765 37777
rect 765 37731 783 37777
rect 807 37731 817 37777
rect 817 37731 833 37777
rect 833 37731 863 37777
rect 887 37731 901 37777
rect 901 37731 943 37777
rect 967 37731 969 37777
rect 969 37731 1021 37777
rect 1021 37731 1023 37777
rect 1047 37731 1089 37777
rect 1089 37731 1103 37777
rect 1127 37731 1157 37777
rect 1157 37731 1173 37777
rect 1173 37731 1183 37777
rect 1207 37731 1225 37777
rect 1225 37731 1241 37777
rect 1241 37731 1263 37777
rect 727 37721 783 37731
rect 807 37721 863 37731
rect 887 37721 943 37731
rect 967 37721 1023 37731
rect 1047 37721 1103 37731
rect 1127 37721 1183 37731
rect 1207 37721 1263 37731
rect 727 37667 749 37696
rect 749 37667 765 37696
rect 765 37667 783 37696
rect 807 37667 817 37696
rect 817 37667 833 37696
rect 833 37667 863 37696
rect 887 37667 901 37696
rect 901 37667 943 37696
rect 967 37667 969 37696
rect 969 37667 1021 37696
rect 1021 37667 1023 37696
rect 1047 37667 1089 37696
rect 1089 37667 1103 37696
rect 1127 37667 1157 37696
rect 1157 37667 1173 37696
rect 1173 37667 1183 37696
rect 1207 37667 1225 37696
rect 1225 37667 1241 37696
rect 1241 37667 1263 37696
rect 727 37655 783 37667
rect 807 37655 863 37667
rect 887 37655 943 37667
rect 967 37655 1023 37667
rect 1047 37655 1103 37667
rect 1127 37655 1183 37667
rect 1207 37655 1263 37667
rect 727 37640 749 37655
rect 749 37640 765 37655
rect 765 37640 783 37655
rect 807 37640 817 37655
rect 817 37640 833 37655
rect 833 37640 863 37655
rect 887 37640 901 37655
rect 901 37640 943 37655
rect 967 37640 969 37655
rect 969 37640 1021 37655
rect 1021 37640 1023 37655
rect 1047 37640 1089 37655
rect 1089 37640 1103 37655
rect 1127 37640 1157 37655
rect 1157 37640 1173 37655
rect 1173 37640 1183 37655
rect 1207 37640 1225 37655
rect 1225 37640 1241 37655
rect 1241 37640 1263 37655
rect 727 37603 749 37615
rect 749 37603 765 37615
rect 765 37603 783 37615
rect 807 37603 817 37615
rect 817 37603 833 37615
rect 833 37603 863 37615
rect 887 37603 901 37615
rect 901 37603 943 37615
rect 967 37603 969 37615
rect 969 37603 1021 37615
rect 1021 37603 1023 37615
rect 1047 37603 1089 37615
rect 1089 37603 1103 37615
rect 1127 37603 1157 37615
rect 1157 37603 1173 37615
rect 1173 37603 1183 37615
rect 1207 37603 1225 37615
rect 1225 37603 1241 37615
rect 1241 37603 1263 37615
rect 727 37591 783 37603
rect 807 37591 863 37603
rect 887 37591 943 37603
rect 967 37591 1023 37603
rect 1047 37591 1103 37603
rect 1127 37591 1183 37603
rect 1207 37591 1263 37603
rect 727 37559 749 37591
rect 749 37559 765 37591
rect 765 37559 783 37591
rect 807 37559 817 37591
rect 817 37559 833 37591
rect 833 37559 863 37591
rect 887 37559 901 37591
rect 901 37559 943 37591
rect 967 37559 969 37591
rect 969 37559 1021 37591
rect 1021 37559 1023 37591
rect 1047 37559 1089 37591
rect 1089 37559 1103 37591
rect 1127 37559 1157 37591
rect 1157 37559 1173 37591
rect 1173 37559 1183 37591
rect 1207 37559 1225 37591
rect 1225 37559 1241 37591
rect 1241 37559 1263 37591
rect 727 37527 783 37534
rect 807 37527 863 37534
rect 887 37527 943 37534
rect 967 37527 1023 37534
rect 1047 37527 1103 37534
rect 1127 37527 1183 37534
rect 1207 37527 1263 37534
rect 727 37478 749 37527
rect 749 37478 765 37527
rect 765 37478 783 37527
rect 807 37478 817 37527
rect 817 37478 833 37527
rect 833 37478 863 37527
rect 887 37478 901 37527
rect 901 37478 943 37527
rect 967 37478 969 37527
rect 969 37478 1021 37527
rect 1021 37478 1023 37527
rect 1047 37478 1089 37527
rect 1089 37478 1103 37527
rect 1127 37478 1157 37527
rect 1157 37478 1173 37527
rect 1173 37478 1183 37527
rect 1207 37478 1225 37527
rect 1225 37478 1241 37527
rect 1241 37478 1263 37527
rect 727 36317 749 36366
rect 749 36317 765 36366
rect 765 36317 817 36366
rect 817 36317 833 36366
rect 833 36317 885 36366
rect 885 36317 901 36366
rect 901 36317 953 36366
rect 953 36317 969 36366
rect 969 36317 1021 36366
rect 1021 36317 1037 36366
rect 1037 36317 1089 36366
rect 1089 36317 1105 36366
rect 1105 36317 1157 36366
rect 1157 36317 1173 36366
rect 1173 36317 1225 36366
rect 1225 36317 1241 36366
rect 1241 36317 1263 36366
rect 727 36305 1263 36317
rect 727 36253 749 36305
rect 749 36253 765 36305
rect 765 36253 817 36305
rect 817 36253 833 36305
rect 833 36253 885 36305
rect 885 36253 901 36305
rect 901 36253 953 36305
rect 953 36253 969 36305
rect 969 36253 1021 36305
rect 1021 36253 1037 36305
rect 1037 36253 1089 36305
rect 1089 36253 1105 36305
rect 1105 36253 1157 36305
rect 1157 36253 1173 36305
rect 1173 36253 1225 36305
rect 1225 36253 1241 36305
rect 1241 36253 1263 36305
rect 727 36241 1263 36253
rect 727 36189 749 36241
rect 749 36189 765 36241
rect 765 36189 817 36241
rect 817 36189 833 36241
rect 833 36189 885 36241
rect 885 36189 901 36241
rect 901 36189 953 36241
rect 953 36189 969 36241
rect 969 36189 1021 36241
rect 1021 36189 1037 36241
rect 1037 36189 1089 36241
rect 1089 36189 1105 36241
rect 1105 36189 1157 36241
rect 1157 36189 1173 36241
rect 1173 36189 1225 36241
rect 1225 36189 1241 36241
rect 1241 36189 1263 36241
rect 727 36177 1263 36189
rect 727 36125 749 36177
rect 749 36125 765 36177
rect 765 36125 817 36177
rect 817 36125 833 36177
rect 833 36125 885 36177
rect 885 36125 901 36177
rect 901 36125 953 36177
rect 953 36125 969 36177
rect 969 36125 1021 36177
rect 1021 36125 1037 36177
rect 1037 36125 1089 36177
rect 1089 36125 1105 36177
rect 1105 36125 1157 36177
rect 1157 36125 1173 36177
rect 1173 36125 1225 36177
rect 1225 36125 1241 36177
rect 1241 36125 1263 36177
rect 727 36113 1263 36125
rect 727 36061 749 36113
rect 749 36061 765 36113
rect 765 36061 817 36113
rect 817 36061 833 36113
rect 833 36061 885 36113
rect 885 36061 901 36113
rect 901 36061 953 36113
rect 953 36061 969 36113
rect 969 36061 1021 36113
rect 1021 36061 1037 36113
rect 1037 36061 1089 36113
rect 1089 36061 1105 36113
rect 1105 36061 1157 36113
rect 1157 36061 1173 36113
rect 1173 36061 1225 36113
rect 1225 36061 1241 36113
rect 1241 36061 1263 36113
rect 727 36049 1263 36061
rect 727 35997 749 36049
rect 749 35997 765 36049
rect 765 35997 817 36049
rect 817 35997 833 36049
rect 833 35997 885 36049
rect 885 35997 901 36049
rect 901 35997 953 36049
rect 953 35997 969 36049
rect 969 35997 1021 36049
rect 1021 35997 1037 36049
rect 1037 35997 1089 36049
rect 1089 35997 1105 36049
rect 1105 35997 1157 36049
rect 1157 35997 1173 36049
rect 1173 35997 1225 36049
rect 1225 35997 1241 36049
rect 1241 35997 1263 36049
rect 727 35985 1263 35997
rect 727 35933 749 35985
rect 749 35933 765 35985
rect 765 35933 817 35985
rect 817 35933 833 35985
rect 833 35933 885 35985
rect 885 35933 901 35985
rect 901 35933 953 35985
rect 953 35933 969 35985
rect 969 35933 1021 35985
rect 1021 35933 1037 35985
rect 1037 35933 1089 35985
rect 1089 35933 1105 35985
rect 1105 35933 1157 35985
rect 1157 35933 1173 35985
rect 1173 35933 1225 35985
rect 1225 35933 1241 35985
rect 1241 35933 1263 35985
rect 727 35921 1263 35933
rect 727 35910 749 35921
rect 749 35910 765 35921
rect 765 35910 817 35921
rect 817 35910 833 35921
rect 833 35910 885 35921
rect 885 35910 901 35921
rect 901 35910 953 35921
rect 953 35910 969 35921
rect 969 35910 1021 35921
rect 1021 35910 1037 35921
rect 1037 35910 1089 35921
rect 1089 35910 1105 35921
rect 1105 35910 1157 35921
rect 1157 35910 1173 35921
rect 1173 35910 1225 35921
rect 1225 35910 1241 35921
rect 1241 35910 1263 35921
rect 727 35869 749 35885
rect 749 35869 765 35885
rect 765 35869 783 35885
rect 807 35869 817 35885
rect 817 35869 833 35885
rect 833 35869 863 35885
rect 887 35869 901 35885
rect 901 35869 943 35885
rect 967 35869 969 35885
rect 969 35869 1021 35885
rect 1021 35869 1023 35885
rect 1047 35869 1089 35885
rect 1089 35869 1103 35885
rect 1127 35869 1157 35885
rect 1157 35869 1173 35885
rect 1173 35869 1183 35885
rect 1207 35869 1225 35885
rect 1225 35869 1241 35885
rect 1241 35869 1263 35885
rect 727 35857 783 35869
rect 807 35857 863 35869
rect 887 35857 943 35869
rect 967 35857 1023 35869
rect 1047 35857 1103 35869
rect 1127 35857 1183 35869
rect 1207 35857 1263 35869
rect 727 35829 749 35857
rect 749 35829 765 35857
rect 765 35829 783 35857
rect 807 35829 817 35857
rect 817 35829 833 35857
rect 833 35829 863 35857
rect 887 35829 901 35857
rect 901 35829 943 35857
rect 967 35829 969 35857
rect 969 35829 1021 35857
rect 1021 35829 1023 35857
rect 1047 35829 1089 35857
rect 1089 35829 1103 35857
rect 1127 35829 1157 35857
rect 1157 35829 1173 35857
rect 1173 35829 1183 35857
rect 1207 35829 1225 35857
rect 1225 35829 1241 35857
rect 1241 35829 1263 35857
rect 727 35793 783 35804
rect 807 35793 863 35804
rect 887 35793 943 35804
rect 967 35793 1023 35804
rect 1047 35793 1103 35804
rect 1127 35793 1183 35804
rect 1207 35793 1263 35804
rect 727 35748 749 35793
rect 749 35748 765 35793
rect 765 35748 783 35793
rect 807 35748 817 35793
rect 817 35748 833 35793
rect 833 35748 863 35793
rect 887 35748 901 35793
rect 901 35748 943 35793
rect 967 35748 969 35793
rect 969 35748 1021 35793
rect 1021 35748 1023 35793
rect 1047 35748 1089 35793
rect 1089 35748 1103 35793
rect 1127 35748 1157 35793
rect 1157 35748 1173 35793
rect 1173 35748 1183 35793
rect 1207 35748 1225 35793
rect 1225 35748 1241 35793
rect 1241 35748 1263 35793
rect 727 35677 749 35723
rect 749 35677 765 35723
rect 765 35677 783 35723
rect 807 35677 817 35723
rect 817 35677 833 35723
rect 833 35677 863 35723
rect 887 35677 901 35723
rect 901 35677 943 35723
rect 967 35677 969 35723
rect 969 35677 1021 35723
rect 1021 35677 1023 35723
rect 1047 35677 1089 35723
rect 1089 35677 1103 35723
rect 1127 35677 1157 35723
rect 1157 35677 1173 35723
rect 1173 35677 1183 35723
rect 1207 35677 1225 35723
rect 1225 35677 1241 35723
rect 1241 35677 1263 35723
rect 727 35667 783 35677
rect 807 35667 863 35677
rect 887 35667 943 35677
rect 967 35667 1023 35677
rect 1047 35667 1103 35677
rect 1127 35667 1183 35677
rect 1207 35667 1263 35677
rect 727 35613 749 35642
rect 749 35613 765 35642
rect 765 35613 783 35642
rect 807 35613 817 35642
rect 817 35613 833 35642
rect 833 35613 863 35642
rect 887 35613 901 35642
rect 901 35613 943 35642
rect 967 35613 969 35642
rect 969 35613 1021 35642
rect 1021 35613 1023 35642
rect 1047 35613 1089 35642
rect 1089 35613 1103 35642
rect 1127 35613 1157 35642
rect 1157 35613 1173 35642
rect 1173 35613 1183 35642
rect 1207 35613 1225 35642
rect 1225 35613 1241 35642
rect 1241 35613 1263 35642
rect 727 35601 783 35613
rect 807 35601 863 35613
rect 887 35601 943 35613
rect 967 35601 1023 35613
rect 1047 35601 1103 35613
rect 1127 35601 1183 35613
rect 1207 35601 1263 35613
rect 727 35586 749 35601
rect 749 35586 765 35601
rect 765 35586 783 35601
rect 807 35586 817 35601
rect 817 35586 833 35601
rect 833 35586 863 35601
rect 887 35586 901 35601
rect 901 35586 943 35601
rect 967 35586 969 35601
rect 969 35586 1021 35601
rect 1021 35586 1023 35601
rect 1047 35586 1089 35601
rect 1089 35586 1103 35601
rect 1127 35586 1157 35601
rect 1157 35586 1173 35601
rect 1173 35586 1183 35601
rect 1207 35586 1225 35601
rect 1225 35586 1241 35601
rect 1241 35586 1263 35601
rect 727 35549 749 35561
rect 749 35549 765 35561
rect 765 35549 783 35561
rect 807 35549 817 35561
rect 817 35549 833 35561
rect 833 35549 863 35561
rect 887 35549 901 35561
rect 901 35549 943 35561
rect 967 35549 969 35561
rect 969 35549 1021 35561
rect 1021 35549 1023 35561
rect 1047 35549 1089 35561
rect 1089 35549 1103 35561
rect 1127 35549 1157 35561
rect 1157 35549 1173 35561
rect 1173 35549 1183 35561
rect 1207 35549 1225 35561
rect 1225 35549 1241 35561
rect 1241 35549 1263 35561
rect 727 35537 783 35549
rect 807 35537 863 35549
rect 887 35537 943 35549
rect 967 35537 1023 35549
rect 1047 35537 1103 35549
rect 1127 35537 1183 35549
rect 1207 35537 1263 35549
rect 727 35505 749 35537
rect 749 35505 765 35537
rect 765 35505 783 35537
rect 807 35505 817 35537
rect 817 35505 833 35537
rect 833 35505 863 35537
rect 887 35505 901 35537
rect 901 35505 943 35537
rect 967 35505 969 35537
rect 969 35505 1021 35537
rect 1021 35505 1023 35537
rect 1047 35505 1089 35537
rect 1089 35505 1103 35537
rect 1127 35505 1157 35537
rect 1157 35505 1173 35537
rect 1173 35505 1183 35537
rect 1207 35505 1225 35537
rect 1225 35505 1241 35537
rect 1241 35505 1263 35537
rect 727 35473 783 35480
rect 807 35473 863 35480
rect 887 35473 943 35480
rect 967 35473 1023 35480
rect 1047 35473 1103 35480
rect 1127 35473 1183 35480
rect 1207 35473 1263 35480
rect 727 35424 749 35473
rect 749 35424 765 35473
rect 765 35424 783 35473
rect 807 35424 817 35473
rect 817 35424 833 35473
rect 833 35424 863 35473
rect 887 35424 901 35473
rect 901 35424 943 35473
rect 967 35424 969 35473
rect 969 35424 1021 35473
rect 1021 35424 1023 35473
rect 1047 35424 1089 35473
rect 1089 35424 1103 35473
rect 1127 35424 1157 35473
rect 1157 35424 1173 35473
rect 1173 35424 1183 35473
rect 1207 35424 1225 35473
rect 1225 35424 1241 35473
rect 1241 35424 1263 35473
rect 727 34098 749 34147
rect 749 34098 765 34147
rect 765 34098 817 34147
rect 817 34098 833 34147
rect 833 34098 885 34147
rect 885 34098 901 34147
rect 901 34098 953 34147
rect 953 34098 969 34147
rect 969 34098 1021 34147
rect 1021 34098 1037 34147
rect 1037 34098 1089 34147
rect 1089 34098 1105 34147
rect 1105 34098 1157 34147
rect 1157 34098 1173 34147
rect 1173 34098 1225 34147
rect 1225 34098 1241 34147
rect 1241 34098 1263 34147
rect 727 34086 1263 34098
rect 727 34034 749 34086
rect 749 34034 765 34086
rect 765 34034 817 34086
rect 817 34034 833 34086
rect 833 34034 885 34086
rect 885 34034 901 34086
rect 901 34034 953 34086
rect 953 34034 969 34086
rect 969 34034 1021 34086
rect 1021 34034 1037 34086
rect 1037 34034 1089 34086
rect 1089 34034 1105 34086
rect 1105 34034 1157 34086
rect 1157 34034 1173 34086
rect 1173 34034 1225 34086
rect 1225 34034 1241 34086
rect 1241 34034 1263 34086
rect 727 34022 1263 34034
rect 727 33970 749 34022
rect 749 33970 765 34022
rect 765 33970 817 34022
rect 817 33970 833 34022
rect 833 33970 885 34022
rect 885 33970 901 34022
rect 901 33970 953 34022
rect 953 33970 969 34022
rect 969 33970 1021 34022
rect 1021 33970 1037 34022
rect 1037 33970 1089 34022
rect 1089 33970 1105 34022
rect 1105 33970 1157 34022
rect 1157 33970 1173 34022
rect 1173 33970 1225 34022
rect 1225 33970 1241 34022
rect 1241 33970 1263 34022
rect 727 33958 1263 33970
rect 727 33906 749 33958
rect 749 33906 765 33958
rect 765 33906 817 33958
rect 817 33906 833 33958
rect 833 33906 885 33958
rect 885 33906 901 33958
rect 901 33906 953 33958
rect 953 33906 969 33958
rect 969 33906 1021 33958
rect 1021 33906 1037 33958
rect 1037 33906 1089 33958
rect 1089 33906 1105 33958
rect 1105 33906 1157 33958
rect 1157 33906 1173 33958
rect 1173 33906 1225 33958
rect 1225 33906 1241 33958
rect 1241 33906 1263 33958
rect 727 33894 1263 33906
rect 727 33842 749 33894
rect 749 33842 765 33894
rect 765 33842 817 33894
rect 817 33842 833 33894
rect 833 33842 885 33894
rect 885 33842 901 33894
rect 901 33842 953 33894
rect 953 33842 969 33894
rect 969 33842 1021 33894
rect 1021 33842 1037 33894
rect 1037 33842 1089 33894
rect 1089 33842 1105 33894
rect 1105 33842 1157 33894
rect 1157 33842 1173 33894
rect 1173 33842 1225 33894
rect 1225 33842 1241 33894
rect 1241 33842 1263 33894
rect 727 33830 1263 33842
rect 727 33778 749 33830
rect 749 33778 765 33830
rect 765 33778 817 33830
rect 817 33778 833 33830
rect 833 33778 885 33830
rect 885 33778 901 33830
rect 901 33778 953 33830
rect 953 33778 969 33830
rect 969 33778 1021 33830
rect 1021 33778 1037 33830
rect 1037 33778 1089 33830
rect 1089 33778 1105 33830
rect 1105 33778 1157 33830
rect 1157 33778 1173 33830
rect 1173 33778 1225 33830
rect 1225 33778 1241 33830
rect 1241 33778 1263 33830
rect 727 33766 1263 33778
rect 727 33714 749 33766
rect 749 33714 765 33766
rect 765 33714 817 33766
rect 817 33714 833 33766
rect 833 33714 885 33766
rect 885 33714 901 33766
rect 901 33714 953 33766
rect 953 33714 969 33766
rect 969 33714 1021 33766
rect 1021 33714 1037 33766
rect 1037 33714 1089 33766
rect 1089 33714 1105 33766
rect 1105 33714 1157 33766
rect 1157 33714 1173 33766
rect 1173 33714 1225 33766
rect 1225 33714 1241 33766
rect 1241 33714 1263 33766
rect 727 33702 1263 33714
rect 727 33691 749 33702
rect 749 33691 765 33702
rect 765 33691 817 33702
rect 817 33691 833 33702
rect 833 33691 885 33702
rect 885 33691 901 33702
rect 901 33691 953 33702
rect 953 33691 969 33702
rect 969 33691 1021 33702
rect 1021 33691 1037 33702
rect 1037 33691 1089 33702
rect 1089 33691 1105 33702
rect 1105 33691 1157 33702
rect 1157 33691 1173 33702
rect 1173 33691 1225 33702
rect 1225 33691 1241 33702
rect 1241 33691 1263 33702
rect 727 33650 749 33666
rect 749 33650 765 33666
rect 765 33650 783 33666
rect 807 33650 817 33666
rect 817 33650 833 33666
rect 833 33650 863 33666
rect 887 33650 901 33666
rect 901 33650 943 33666
rect 967 33650 969 33666
rect 969 33650 1021 33666
rect 1021 33650 1023 33666
rect 1047 33650 1089 33666
rect 1089 33650 1103 33666
rect 1127 33650 1157 33666
rect 1157 33650 1173 33666
rect 1173 33650 1183 33666
rect 1207 33650 1225 33666
rect 1225 33650 1241 33666
rect 1241 33650 1263 33666
rect 727 33638 783 33650
rect 807 33638 863 33650
rect 887 33638 943 33650
rect 967 33638 1023 33650
rect 1047 33638 1103 33650
rect 1127 33638 1183 33650
rect 1207 33638 1263 33650
rect 727 33610 749 33638
rect 749 33610 765 33638
rect 765 33610 783 33638
rect 807 33610 817 33638
rect 817 33610 833 33638
rect 833 33610 863 33638
rect 887 33610 901 33638
rect 901 33610 943 33638
rect 967 33610 969 33638
rect 969 33610 1021 33638
rect 1021 33610 1023 33638
rect 1047 33610 1089 33638
rect 1089 33610 1103 33638
rect 1127 33610 1157 33638
rect 1157 33610 1173 33638
rect 1173 33610 1183 33638
rect 1207 33610 1225 33638
rect 1225 33610 1241 33638
rect 1241 33610 1263 33638
rect 727 33574 783 33585
rect 807 33574 863 33585
rect 887 33574 943 33585
rect 967 33574 1023 33585
rect 1047 33574 1103 33585
rect 1127 33574 1183 33585
rect 1207 33574 1263 33585
rect 727 33529 749 33574
rect 749 33529 765 33574
rect 765 33529 783 33574
rect 807 33529 817 33574
rect 817 33529 833 33574
rect 833 33529 863 33574
rect 887 33529 901 33574
rect 901 33529 943 33574
rect 967 33529 969 33574
rect 969 33529 1021 33574
rect 1021 33529 1023 33574
rect 1047 33529 1089 33574
rect 1089 33529 1103 33574
rect 1127 33529 1157 33574
rect 1157 33529 1173 33574
rect 1173 33529 1183 33574
rect 1207 33529 1225 33574
rect 1225 33529 1241 33574
rect 1241 33529 1263 33574
rect 727 33458 749 33504
rect 749 33458 765 33504
rect 765 33458 783 33504
rect 807 33458 817 33504
rect 817 33458 833 33504
rect 833 33458 863 33504
rect 887 33458 901 33504
rect 901 33458 943 33504
rect 967 33458 969 33504
rect 969 33458 1021 33504
rect 1021 33458 1023 33504
rect 1047 33458 1089 33504
rect 1089 33458 1103 33504
rect 1127 33458 1157 33504
rect 1157 33458 1173 33504
rect 1173 33458 1183 33504
rect 1207 33458 1225 33504
rect 1225 33458 1241 33504
rect 1241 33458 1263 33504
rect 727 33448 783 33458
rect 807 33448 863 33458
rect 887 33448 943 33458
rect 967 33448 1023 33458
rect 1047 33448 1103 33458
rect 1127 33448 1183 33458
rect 1207 33448 1263 33458
rect 727 33394 749 33423
rect 749 33394 765 33423
rect 765 33394 783 33423
rect 807 33394 817 33423
rect 817 33394 833 33423
rect 833 33394 863 33423
rect 887 33394 901 33423
rect 901 33394 943 33423
rect 967 33394 969 33423
rect 969 33394 1021 33423
rect 1021 33394 1023 33423
rect 1047 33394 1089 33423
rect 1089 33394 1103 33423
rect 1127 33394 1157 33423
rect 1157 33394 1173 33423
rect 1173 33394 1183 33423
rect 1207 33394 1225 33423
rect 1225 33394 1241 33423
rect 1241 33394 1263 33423
rect 727 33382 783 33394
rect 807 33382 863 33394
rect 887 33382 943 33394
rect 967 33382 1023 33394
rect 1047 33382 1103 33394
rect 1127 33382 1183 33394
rect 1207 33382 1263 33394
rect 727 33367 749 33382
rect 749 33367 765 33382
rect 765 33367 783 33382
rect 807 33367 817 33382
rect 817 33367 833 33382
rect 833 33367 863 33382
rect 887 33367 901 33382
rect 901 33367 943 33382
rect 967 33367 969 33382
rect 969 33367 1021 33382
rect 1021 33367 1023 33382
rect 1047 33367 1089 33382
rect 1089 33367 1103 33382
rect 1127 33367 1157 33382
rect 1157 33367 1173 33382
rect 1173 33367 1183 33382
rect 1207 33367 1225 33382
rect 1225 33367 1241 33382
rect 1241 33367 1263 33382
rect 727 33330 749 33342
rect 749 33330 765 33342
rect 765 33330 783 33342
rect 807 33330 817 33342
rect 817 33330 833 33342
rect 833 33330 863 33342
rect 887 33330 901 33342
rect 901 33330 943 33342
rect 967 33330 969 33342
rect 969 33330 1021 33342
rect 1021 33330 1023 33342
rect 1047 33330 1089 33342
rect 1089 33330 1103 33342
rect 1127 33330 1157 33342
rect 1157 33330 1173 33342
rect 1173 33330 1183 33342
rect 1207 33330 1225 33342
rect 1225 33330 1241 33342
rect 1241 33330 1263 33342
rect 727 33318 783 33330
rect 807 33318 863 33330
rect 887 33318 943 33330
rect 967 33318 1023 33330
rect 1047 33318 1103 33330
rect 1127 33318 1183 33330
rect 1207 33318 1263 33330
rect 727 33286 749 33318
rect 749 33286 765 33318
rect 765 33286 783 33318
rect 807 33286 817 33318
rect 817 33286 833 33318
rect 833 33286 863 33318
rect 887 33286 901 33318
rect 901 33286 943 33318
rect 967 33286 969 33318
rect 969 33286 1021 33318
rect 1021 33286 1023 33318
rect 1047 33286 1089 33318
rect 1089 33286 1103 33318
rect 1127 33286 1157 33318
rect 1157 33286 1173 33318
rect 1173 33286 1183 33318
rect 1207 33286 1225 33318
rect 1225 33286 1241 33318
rect 1241 33286 1263 33318
rect 727 33254 783 33261
rect 807 33254 863 33261
rect 887 33254 943 33261
rect 967 33254 1023 33261
rect 1047 33254 1103 33261
rect 1127 33254 1183 33261
rect 1207 33254 1263 33261
rect 727 33205 749 33254
rect 749 33205 765 33254
rect 765 33205 783 33254
rect 807 33205 817 33254
rect 817 33205 833 33254
rect 833 33205 863 33254
rect 887 33205 901 33254
rect 901 33205 943 33254
rect 967 33205 969 33254
rect 969 33205 1021 33254
rect 1021 33205 1023 33254
rect 1047 33205 1089 33254
rect 1089 33205 1103 33254
rect 1127 33205 1157 33254
rect 1157 33205 1173 33254
rect 1173 33205 1183 33254
rect 1207 33205 1225 33254
rect 1225 33205 1241 33254
rect 1241 33205 1263 33254
rect 727 31969 749 32018
rect 749 31969 765 32018
rect 765 31969 817 32018
rect 817 31969 833 32018
rect 833 31969 885 32018
rect 885 31969 901 32018
rect 901 31969 953 32018
rect 953 31969 969 32018
rect 969 31969 1021 32018
rect 1021 31969 1037 32018
rect 1037 31969 1089 32018
rect 1089 31969 1105 32018
rect 1105 31969 1157 32018
rect 1157 31969 1173 32018
rect 1173 31969 1225 32018
rect 1225 31969 1241 32018
rect 1241 31969 1263 32018
rect 727 31957 1263 31969
rect 727 31905 749 31957
rect 749 31905 765 31957
rect 765 31905 817 31957
rect 817 31905 833 31957
rect 833 31905 885 31957
rect 885 31905 901 31957
rect 901 31905 953 31957
rect 953 31905 969 31957
rect 969 31905 1021 31957
rect 1021 31905 1037 31957
rect 1037 31905 1089 31957
rect 1089 31905 1105 31957
rect 1105 31905 1157 31957
rect 1157 31905 1173 31957
rect 1173 31905 1225 31957
rect 1225 31905 1241 31957
rect 1241 31905 1263 31957
rect 727 31893 1263 31905
rect 727 31841 749 31893
rect 749 31841 765 31893
rect 765 31841 817 31893
rect 817 31841 833 31893
rect 833 31841 885 31893
rect 885 31841 901 31893
rect 901 31841 953 31893
rect 953 31841 969 31893
rect 969 31841 1021 31893
rect 1021 31841 1037 31893
rect 1037 31841 1089 31893
rect 1089 31841 1105 31893
rect 1105 31841 1157 31893
rect 1157 31841 1173 31893
rect 1173 31841 1225 31893
rect 1225 31841 1241 31893
rect 1241 31841 1263 31893
rect 727 31829 1263 31841
rect 727 31777 749 31829
rect 749 31777 765 31829
rect 765 31777 817 31829
rect 817 31777 833 31829
rect 833 31777 885 31829
rect 885 31777 901 31829
rect 901 31777 953 31829
rect 953 31777 969 31829
rect 969 31777 1021 31829
rect 1021 31777 1037 31829
rect 1037 31777 1089 31829
rect 1089 31777 1105 31829
rect 1105 31777 1157 31829
rect 1157 31777 1173 31829
rect 1173 31777 1225 31829
rect 1225 31777 1241 31829
rect 1241 31777 1263 31829
rect 727 31765 1263 31777
rect 727 31713 749 31765
rect 749 31713 765 31765
rect 765 31713 817 31765
rect 817 31713 833 31765
rect 833 31713 885 31765
rect 885 31713 901 31765
rect 901 31713 953 31765
rect 953 31713 969 31765
rect 969 31713 1021 31765
rect 1021 31713 1037 31765
rect 1037 31713 1089 31765
rect 1089 31713 1105 31765
rect 1105 31713 1157 31765
rect 1157 31713 1173 31765
rect 1173 31713 1225 31765
rect 1225 31713 1241 31765
rect 1241 31713 1263 31765
rect 727 31701 1263 31713
rect 727 31649 749 31701
rect 749 31649 765 31701
rect 765 31649 817 31701
rect 817 31649 833 31701
rect 833 31649 885 31701
rect 885 31649 901 31701
rect 901 31649 953 31701
rect 953 31649 969 31701
rect 969 31649 1021 31701
rect 1021 31649 1037 31701
rect 1037 31649 1089 31701
rect 1089 31649 1105 31701
rect 1105 31649 1157 31701
rect 1157 31649 1173 31701
rect 1173 31649 1225 31701
rect 1225 31649 1241 31701
rect 1241 31649 1263 31701
rect 727 31637 1263 31649
rect 727 31585 749 31637
rect 749 31585 765 31637
rect 765 31585 817 31637
rect 817 31585 833 31637
rect 833 31585 885 31637
rect 885 31585 901 31637
rect 901 31585 953 31637
rect 953 31585 969 31637
rect 969 31585 1021 31637
rect 1021 31585 1037 31637
rect 1037 31585 1089 31637
rect 1089 31585 1105 31637
rect 1105 31585 1157 31637
rect 1157 31585 1173 31637
rect 1173 31585 1225 31637
rect 1225 31585 1241 31637
rect 1241 31585 1263 31637
rect 727 31573 1263 31585
rect 727 31562 749 31573
rect 749 31562 765 31573
rect 765 31562 817 31573
rect 817 31562 833 31573
rect 833 31562 885 31573
rect 885 31562 901 31573
rect 901 31562 953 31573
rect 953 31562 969 31573
rect 969 31562 1021 31573
rect 1021 31562 1037 31573
rect 1037 31562 1089 31573
rect 1089 31562 1105 31573
rect 1105 31562 1157 31573
rect 1157 31562 1173 31573
rect 1173 31562 1225 31573
rect 1225 31562 1241 31573
rect 1241 31562 1263 31573
rect 727 31521 749 31537
rect 749 31521 765 31537
rect 765 31521 783 31537
rect 807 31521 817 31537
rect 817 31521 833 31537
rect 833 31521 863 31537
rect 887 31521 901 31537
rect 901 31521 943 31537
rect 967 31521 969 31537
rect 969 31521 1021 31537
rect 1021 31521 1023 31537
rect 1047 31521 1089 31537
rect 1089 31521 1103 31537
rect 1127 31521 1157 31537
rect 1157 31521 1173 31537
rect 1173 31521 1183 31537
rect 1207 31521 1225 31537
rect 1225 31521 1241 31537
rect 1241 31521 1263 31537
rect 727 31509 783 31521
rect 807 31509 863 31521
rect 887 31509 943 31521
rect 967 31509 1023 31521
rect 1047 31509 1103 31521
rect 1127 31509 1183 31521
rect 1207 31509 1263 31521
rect 727 31481 749 31509
rect 749 31481 765 31509
rect 765 31481 783 31509
rect 807 31481 817 31509
rect 817 31481 833 31509
rect 833 31481 863 31509
rect 887 31481 901 31509
rect 901 31481 943 31509
rect 967 31481 969 31509
rect 969 31481 1021 31509
rect 1021 31481 1023 31509
rect 1047 31481 1089 31509
rect 1089 31481 1103 31509
rect 1127 31481 1157 31509
rect 1157 31481 1173 31509
rect 1173 31481 1183 31509
rect 1207 31481 1225 31509
rect 1225 31481 1241 31509
rect 1241 31481 1263 31509
rect 727 31445 783 31456
rect 807 31445 863 31456
rect 887 31445 943 31456
rect 967 31445 1023 31456
rect 1047 31445 1103 31456
rect 1127 31445 1183 31456
rect 1207 31445 1263 31456
rect 727 31400 749 31445
rect 749 31400 765 31445
rect 765 31400 783 31445
rect 807 31400 817 31445
rect 817 31400 833 31445
rect 833 31400 863 31445
rect 887 31400 901 31445
rect 901 31400 943 31445
rect 967 31400 969 31445
rect 969 31400 1021 31445
rect 1021 31400 1023 31445
rect 1047 31400 1089 31445
rect 1089 31400 1103 31445
rect 1127 31400 1157 31445
rect 1157 31400 1173 31445
rect 1173 31400 1183 31445
rect 1207 31400 1225 31445
rect 1225 31400 1241 31445
rect 1241 31400 1263 31445
rect 727 31329 749 31375
rect 749 31329 765 31375
rect 765 31329 783 31375
rect 807 31329 817 31375
rect 817 31329 833 31375
rect 833 31329 863 31375
rect 887 31329 901 31375
rect 901 31329 943 31375
rect 967 31329 969 31375
rect 969 31329 1021 31375
rect 1021 31329 1023 31375
rect 1047 31329 1089 31375
rect 1089 31329 1103 31375
rect 1127 31329 1157 31375
rect 1157 31329 1173 31375
rect 1173 31329 1183 31375
rect 1207 31329 1225 31375
rect 1225 31329 1241 31375
rect 1241 31329 1263 31375
rect 727 31319 783 31329
rect 807 31319 863 31329
rect 887 31319 943 31329
rect 967 31319 1023 31329
rect 1047 31319 1103 31329
rect 1127 31319 1183 31329
rect 1207 31319 1263 31329
rect 727 31265 749 31294
rect 749 31265 765 31294
rect 765 31265 783 31294
rect 807 31265 817 31294
rect 817 31265 833 31294
rect 833 31265 863 31294
rect 887 31265 901 31294
rect 901 31265 943 31294
rect 967 31265 969 31294
rect 969 31265 1021 31294
rect 1021 31265 1023 31294
rect 1047 31265 1089 31294
rect 1089 31265 1103 31294
rect 1127 31265 1157 31294
rect 1157 31265 1173 31294
rect 1173 31265 1183 31294
rect 1207 31265 1225 31294
rect 1225 31265 1241 31294
rect 1241 31265 1263 31294
rect 727 31253 783 31265
rect 807 31253 863 31265
rect 887 31253 943 31265
rect 967 31253 1023 31265
rect 1047 31253 1103 31265
rect 1127 31253 1183 31265
rect 1207 31253 1263 31265
rect 727 31238 749 31253
rect 749 31238 765 31253
rect 765 31238 783 31253
rect 807 31238 817 31253
rect 817 31238 833 31253
rect 833 31238 863 31253
rect 887 31238 901 31253
rect 901 31238 943 31253
rect 967 31238 969 31253
rect 969 31238 1021 31253
rect 1021 31238 1023 31253
rect 1047 31238 1089 31253
rect 1089 31238 1103 31253
rect 1127 31238 1157 31253
rect 1157 31238 1173 31253
rect 1173 31238 1183 31253
rect 1207 31238 1225 31253
rect 1225 31238 1241 31253
rect 1241 31238 1263 31253
rect 727 31201 749 31213
rect 749 31201 765 31213
rect 765 31201 783 31213
rect 807 31201 817 31213
rect 817 31201 833 31213
rect 833 31201 863 31213
rect 887 31201 901 31213
rect 901 31201 943 31213
rect 967 31201 969 31213
rect 969 31201 1021 31213
rect 1021 31201 1023 31213
rect 1047 31201 1089 31213
rect 1089 31201 1103 31213
rect 1127 31201 1157 31213
rect 1157 31201 1173 31213
rect 1173 31201 1183 31213
rect 1207 31201 1225 31213
rect 1225 31201 1241 31213
rect 1241 31201 1263 31213
rect 727 31189 783 31201
rect 807 31189 863 31201
rect 887 31189 943 31201
rect 967 31189 1023 31201
rect 1047 31189 1103 31201
rect 1127 31189 1183 31201
rect 1207 31189 1263 31201
rect 727 31157 749 31189
rect 749 31157 765 31189
rect 765 31157 783 31189
rect 807 31157 817 31189
rect 817 31157 833 31189
rect 833 31157 863 31189
rect 887 31157 901 31189
rect 901 31157 943 31189
rect 967 31157 969 31189
rect 969 31157 1021 31189
rect 1021 31157 1023 31189
rect 1047 31157 1089 31189
rect 1089 31157 1103 31189
rect 1127 31157 1157 31189
rect 1157 31157 1173 31189
rect 1173 31157 1183 31189
rect 1207 31157 1225 31189
rect 1225 31157 1241 31189
rect 1241 31157 1263 31189
rect 727 31125 783 31132
rect 807 31125 863 31132
rect 887 31125 943 31132
rect 967 31125 1023 31132
rect 1047 31125 1103 31132
rect 1127 31125 1183 31132
rect 1207 31125 1263 31132
rect 727 31076 749 31125
rect 749 31076 765 31125
rect 765 31076 783 31125
rect 807 31076 817 31125
rect 817 31076 833 31125
rect 833 31076 863 31125
rect 887 31076 901 31125
rect 901 31076 943 31125
rect 967 31076 969 31125
rect 969 31076 1021 31125
rect 1021 31076 1023 31125
rect 1047 31076 1089 31125
rect 1089 31076 1103 31125
rect 1127 31076 1157 31125
rect 1157 31076 1173 31125
rect 1173 31076 1183 31125
rect 1207 31076 1225 31125
rect 1225 31076 1241 31125
rect 1241 31076 1263 31125
rect 727 29820 749 29869
rect 749 29820 765 29869
rect 765 29820 817 29869
rect 817 29820 833 29869
rect 833 29820 885 29869
rect 885 29820 901 29869
rect 901 29820 953 29869
rect 953 29820 969 29869
rect 969 29820 1021 29869
rect 1021 29820 1037 29869
rect 1037 29820 1089 29869
rect 1089 29820 1105 29869
rect 1105 29820 1157 29869
rect 1157 29820 1173 29869
rect 1173 29820 1225 29869
rect 1225 29820 1241 29869
rect 1241 29820 1263 29869
rect 727 29808 1263 29820
rect 727 29756 749 29808
rect 749 29756 765 29808
rect 765 29756 817 29808
rect 817 29756 833 29808
rect 833 29756 885 29808
rect 885 29756 901 29808
rect 901 29756 953 29808
rect 953 29756 969 29808
rect 969 29756 1021 29808
rect 1021 29756 1037 29808
rect 1037 29756 1089 29808
rect 1089 29756 1105 29808
rect 1105 29756 1157 29808
rect 1157 29756 1173 29808
rect 1173 29756 1225 29808
rect 1225 29756 1241 29808
rect 1241 29756 1263 29808
rect 727 29744 1263 29756
rect 727 29692 749 29744
rect 749 29692 765 29744
rect 765 29692 817 29744
rect 817 29692 833 29744
rect 833 29692 885 29744
rect 885 29692 901 29744
rect 901 29692 953 29744
rect 953 29692 969 29744
rect 969 29692 1021 29744
rect 1021 29692 1037 29744
rect 1037 29692 1089 29744
rect 1089 29692 1105 29744
rect 1105 29692 1157 29744
rect 1157 29692 1173 29744
rect 1173 29692 1225 29744
rect 1225 29692 1241 29744
rect 1241 29692 1263 29744
rect 727 29680 1263 29692
rect 727 29628 749 29680
rect 749 29628 765 29680
rect 765 29628 817 29680
rect 817 29628 833 29680
rect 833 29628 885 29680
rect 885 29628 901 29680
rect 901 29628 953 29680
rect 953 29628 969 29680
rect 969 29628 1021 29680
rect 1021 29628 1037 29680
rect 1037 29628 1089 29680
rect 1089 29628 1105 29680
rect 1105 29628 1157 29680
rect 1157 29628 1173 29680
rect 1173 29628 1225 29680
rect 1225 29628 1241 29680
rect 1241 29628 1263 29680
rect 727 29616 1263 29628
rect 727 29564 749 29616
rect 749 29564 765 29616
rect 765 29564 817 29616
rect 817 29564 833 29616
rect 833 29564 885 29616
rect 885 29564 901 29616
rect 901 29564 953 29616
rect 953 29564 969 29616
rect 969 29564 1021 29616
rect 1021 29564 1037 29616
rect 1037 29564 1089 29616
rect 1089 29564 1105 29616
rect 1105 29564 1157 29616
rect 1157 29564 1173 29616
rect 1173 29564 1225 29616
rect 1225 29564 1241 29616
rect 1241 29564 1263 29616
rect 727 29552 1263 29564
rect 727 29500 749 29552
rect 749 29500 765 29552
rect 765 29500 817 29552
rect 817 29500 833 29552
rect 833 29500 885 29552
rect 885 29500 901 29552
rect 901 29500 953 29552
rect 953 29500 969 29552
rect 969 29500 1021 29552
rect 1021 29500 1037 29552
rect 1037 29500 1089 29552
rect 1089 29500 1105 29552
rect 1105 29500 1157 29552
rect 1157 29500 1173 29552
rect 1173 29500 1225 29552
rect 1225 29500 1241 29552
rect 1241 29500 1263 29552
rect 727 29488 1263 29500
rect 727 29436 749 29488
rect 749 29436 765 29488
rect 765 29436 817 29488
rect 817 29436 833 29488
rect 833 29436 885 29488
rect 885 29436 901 29488
rect 901 29436 953 29488
rect 953 29436 969 29488
rect 969 29436 1021 29488
rect 1021 29436 1037 29488
rect 1037 29436 1089 29488
rect 1089 29436 1105 29488
rect 1105 29436 1157 29488
rect 1157 29436 1173 29488
rect 1173 29436 1225 29488
rect 1225 29436 1241 29488
rect 1241 29436 1263 29488
rect 727 29424 1263 29436
rect 727 29413 749 29424
rect 749 29413 765 29424
rect 765 29413 817 29424
rect 817 29413 833 29424
rect 833 29413 885 29424
rect 885 29413 901 29424
rect 901 29413 953 29424
rect 953 29413 969 29424
rect 969 29413 1021 29424
rect 1021 29413 1037 29424
rect 1037 29413 1089 29424
rect 1089 29413 1105 29424
rect 1105 29413 1157 29424
rect 1157 29413 1173 29424
rect 1173 29413 1225 29424
rect 1225 29413 1241 29424
rect 1241 29413 1263 29424
rect 727 29372 749 29388
rect 749 29372 765 29388
rect 765 29372 783 29388
rect 807 29372 817 29388
rect 817 29372 833 29388
rect 833 29372 863 29388
rect 887 29372 901 29388
rect 901 29372 943 29388
rect 967 29372 969 29388
rect 969 29372 1021 29388
rect 1021 29372 1023 29388
rect 1047 29372 1089 29388
rect 1089 29372 1103 29388
rect 1127 29372 1157 29388
rect 1157 29372 1173 29388
rect 1173 29372 1183 29388
rect 1207 29372 1225 29388
rect 1225 29372 1241 29388
rect 1241 29372 1263 29388
rect 727 29360 783 29372
rect 807 29360 863 29372
rect 887 29360 943 29372
rect 967 29360 1023 29372
rect 1047 29360 1103 29372
rect 1127 29360 1183 29372
rect 1207 29360 1263 29372
rect 727 29332 749 29360
rect 749 29332 765 29360
rect 765 29332 783 29360
rect 807 29332 817 29360
rect 817 29332 833 29360
rect 833 29332 863 29360
rect 887 29332 901 29360
rect 901 29332 943 29360
rect 967 29332 969 29360
rect 969 29332 1021 29360
rect 1021 29332 1023 29360
rect 1047 29332 1089 29360
rect 1089 29332 1103 29360
rect 1127 29332 1157 29360
rect 1157 29332 1173 29360
rect 1173 29332 1183 29360
rect 1207 29332 1225 29360
rect 1225 29332 1241 29360
rect 1241 29332 1263 29360
rect 727 29296 783 29307
rect 807 29296 863 29307
rect 887 29296 943 29307
rect 967 29296 1023 29307
rect 1047 29296 1103 29307
rect 1127 29296 1183 29307
rect 1207 29296 1263 29307
rect 727 29251 749 29296
rect 749 29251 765 29296
rect 765 29251 783 29296
rect 807 29251 817 29296
rect 817 29251 833 29296
rect 833 29251 863 29296
rect 887 29251 901 29296
rect 901 29251 943 29296
rect 967 29251 969 29296
rect 969 29251 1021 29296
rect 1021 29251 1023 29296
rect 1047 29251 1089 29296
rect 1089 29251 1103 29296
rect 1127 29251 1157 29296
rect 1157 29251 1173 29296
rect 1173 29251 1183 29296
rect 1207 29251 1225 29296
rect 1225 29251 1241 29296
rect 1241 29251 1263 29296
rect 727 29180 749 29226
rect 749 29180 765 29226
rect 765 29180 783 29226
rect 807 29180 817 29226
rect 817 29180 833 29226
rect 833 29180 863 29226
rect 887 29180 901 29226
rect 901 29180 943 29226
rect 967 29180 969 29226
rect 969 29180 1021 29226
rect 1021 29180 1023 29226
rect 1047 29180 1089 29226
rect 1089 29180 1103 29226
rect 1127 29180 1157 29226
rect 1157 29180 1173 29226
rect 1173 29180 1183 29226
rect 1207 29180 1225 29226
rect 1225 29180 1241 29226
rect 1241 29180 1263 29226
rect 727 29170 783 29180
rect 807 29170 863 29180
rect 887 29170 943 29180
rect 967 29170 1023 29180
rect 1047 29170 1103 29180
rect 1127 29170 1183 29180
rect 1207 29170 1263 29180
rect 727 29116 749 29145
rect 749 29116 765 29145
rect 765 29116 783 29145
rect 807 29116 817 29145
rect 817 29116 833 29145
rect 833 29116 863 29145
rect 887 29116 901 29145
rect 901 29116 943 29145
rect 967 29116 969 29145
rect 969 29116 1021 29145
rect 1021 29116 1023 29145
rect 1047 29116 1089 29145
rect 1089 29116 1103 29145
rect 1127 29116 1157 29145
rect 1157 29116 1173 29145
rect 1173 29116 1183 29145
rect 1207 29116 1225 29145
rect 1225 29116 1241 29145
rect 1241 29116 1263 29145
rect 727 29104 783 29116
rect 807 29104 863 29116
rect 887 29104 943 29116
rect 967 29104 1023 29116
rect 1047 29104 1103 29116
rect 1127 29104 1183 29116
rect 1207 29104 1263 29116
rect 727 29089 749 29104
rect 749 29089 765 29104
rect 765 29089 783 29104
rect 807 29089 817 29104
rect 817 29089 833 29104
rect 833 29089 863 29104
rect 887 29089 901 29104
rect 901 29089 943 29104
rect 967 29089 969 29104
rect 969 29089 1021 29104
rect 1021 29089 1023 29104
rect 1047 29089 1089 29104
rect 1089 29089 1103 29104
rect 1127 29089 1157 29104
rect 1157 29089 1173 29104
rect 1173 29089 1183 29104
rect 1207 29089 1225 29104
rect 1225 29089 1241 29104
rect 1241 29089 1263 29104
rect 727 29052 749 29064
rect 749 29052 765 29064
rect 765 29052 783 29064
rect 807 29052 817 29064
rect 817 29052 833 29064
rect 833 29052 863 29064
rect 887 29052 901 29064
rect 901 29052 943 29064
rect 967 29052 969 29064
rect 969 29052 1021 29064
rect 1021 29052 1023 29064
rect 1047 29052 1089 29064
rect 1089 29052 1103 29064
rect 1127 29052 1157 29064
rect 1157 29052 1173 29064
rect 1173 29052 1183 29064
rect 1207 29052 1225 29064
rect 1225 29052 1241 29064
rect 1241 29052 1263 29064
rect 727 29040 783 29052
rect 807 29040 863 29052
rect 887 29040 943 29052
rect 967 29040 1023 29052
rect 1047 29040 1103 29052
rect 1127 29040 1183 29052
rect 1207 29040 1263 29052
rect 727 29008 749 29040
rect 749 29008 765 29040
rect 765 29008 783 29040
rect 807 29008 817 29040
rect 817 29008 833 29040
rect 833 29008 863 29040
rect 887 29008 901 29040
rect 901 29008 943 29040
rect 967 29008 969 29040
rect 969 29008 1021 29040
rect 1021 29008 1023 29040
rect 1047 29008 1089 29040
rect 1089 29008 1103 29040
rect 1127 29008 1157 29040
rect 1157 29008 1173 29040
rect 1173 29008 1183 29040
rect 1207 29008 1225 29040
rect 1225 29008 1241 29040
rect 1241 29008 1263 29040
rect 727 28976 783 28983
rect 807 28976 863 28983
rect 887 28976 943 28983
rect 967 28976 1023 28983
rect 1047 28976 1103 28983
rect 1127 28976 1183 28983
rect 1207 28976 1263 28983
rect 727 28927 749 28976
rect 749 28927 765 28976
rect 765 28927 783 28976
rect 807 28927 817 28976
rect 817 28927 833 28976
rect 833 28927 863 28976
rect 887 28927 901 28976
rect 901 28927 943 28976
rect 967 28927 969 28976
rect 969 28927 1021 28976
rect 1021 28927 1023 28976
rect 1047 28927 1089 28976
rect 1089 28927 1103 28976
rect 1127 28927 1157 28976
rect 1157 28927 1173 28976
rect 1173 28927 1183 28976
rect 1207 28927 1225 28976
rect 1225 28927 1241 28976
rect 1241 28927 1263 28976
rect 727 27813 749 27862
rect 749 27813 765 27862
rect 765 27813 817 27862
rect 817 27813 833 27862
rect 833 27813 885 27862
rect 885 27813 901 27862
rect 901 27813 953 27862
rect 953 27813 969 27862
rect 969 27813 1021 27862
rect 1021 27813 1037 27862
rect 1037 27813 1089 27862
rect 1089 27813 1105 27862
rect 1105 27813 1157 27862
rect 1157 27813 1173 27862
rect 1173 27813 1225 27862
rect 1225 27813 1241 27862
rect 1241 27813 1263 27862
rect 727 27801 1263 27813
rect 727 27749 749 27801
rect 749 27749 765 27801
rect 765 27749 817 27801
rect 817 27749 833 27801
rect 833 27749 885 27801
rect 885 27749 901 27801
rect 901 27749 953 27801
rect 953 27749 969 27801
rect 969 27749 1021 27801
rect 1021 27749 1037 27801
rect 1037 27749 1089 27801
rect 1089 27749 1105 27801
rect 1105 27749 1157 27801
rect 1157 27749 1173 27801
rect 1173 27749 1225 27801
rect 1225 27749 1241 27801
rect 1241 27749 1263 27801
rect 727 27737 1263 27749
rect 727 27685 749 27737
rect 749 27685 765 27737
rect 765 27685 817 27737
rect 817 27685 833 27737
rect 833 27685 885 27737
rect 885 27685 901 27737
rect 901 27685 953 27737
rect 953 27685 969 27737
rect 969 27685 1021 27737
rect 1021 27685 1037 27737
rect 1037 27685 1089 27737
rect 1089 27685 1105 27737
rect 1105 27685 1157 27737
rect 1157 27685 1173 27737
rect 1173 27685 1225 27737
rect 1225 27685 1241 27737
rect 1241 27685 1263 27737
rect 727 27673 1263 27685
rect 727 27621 749 27673
rect 749 27621 765 27673
rect 765 27621 817 27673
rect 817 27621 833 27673
rect 833 27621 885 27673
rect 885 27621 901 27673
rect 901 27621 953 27673
rect 953 27621 969 27673
rect 969 27621 1021 27673
rect 1021 27621 1037 27673
rect 1037 27621 1089 27673
rect 1089 27621 1105 27673
rect 1105 27621 1157 27673
rect 1157 27621 1173 27673
rect 1173 27621 1225 27673
rect 1225 27621 1241 27673
rect 1241 27621 1263 27673
rect 727 27609 1263 27621
rect 727 27557 749 27609
rect 749 27557 765 27609
rect 765 27557 817 27609
rect 817 27557 833 27609
rect 833 27557 885 27609
rect 885 27557 901 27609
rect 901 27557 953 27609
rect 953 27557 969 27609
rect 969 27557 1021 27609
rect 1021 27557 1037 27609
rect 1037 27557 1089 27609
rect 1089 27557 1105 27609
rect 1105 27557 1157 27609
rect 1157 27557 1173 27609
rect 1173 27557 1225 27609
rect 1225 27557 1241 27609
rect 1241 27557 1263 27609
rect 727 27545 1263 27557
rect 727 27493 749 27545
rect 749 27493 765 27545
rect 765 27493 817 27545
rect 817 27493 833 27545
rect 833 27493 885 27545
rect 885 27493 901 27545
rect 901 27493 953 27545
rect 953 27493 969 27545
rect 969 27493 1021 27545
rect 1021 27493 1037 27545
rect 1037 27493 1089 27545
rect 1089 27493 1105 27545
rect 1105 27493 1157 27545
rect 1157 27493 1173 27545
rect 1173 27493 1225 27545
rect 1225 27493 1241 27545
rect 1241 27493 1263 27545
rect 727 27481 1263 27493
rect 727 27429 749 27481
rect 749 27429 765 27481
rect 765 27429 817 27481
rect 817 27429 833 27481
rect 833 27429 885 27481
rect 885 27429 901 27481
rect 901 27429 953 27481
rect 953 27429 969 27481
rect 969 27429 1021 27481
rect 1021 27429 1037 27481
rect 1037 27429 1089 27481
rect 1089 27429 1105 27481
rect 1105 27429 1157 27481
rect 1157 27429 1173 27481
rect 1173 27429 1225 27481
rect 1225 27429 1241 27481
rect 1241 27429 1263 27481
rect 727 27417 1263 27429
rect 727 27406 749 27417
rect 749 27406 765 27417
rect 765 27406 817 27417
rect 817 27406 833 27417
rect 833 27406 885 27417
rect 885 27406 901 27417
rect 901 27406 953 27417
rect 953 27406 969 27417
rect 969 27406 1021 27417
rect 1021 27406 1037 27417
rect 1037 27406 1089 27417
rect 1089 27406 1105 27417
rect 1105 27406 1157 27417
rect 1157 27406 1173 27417
rect 1173 27406 1225 27417
rect 1225 27406 1241 27417
rect 1241 27406 1263 27417
rect 727 27365 749 27381
rect 749 27365 765 27381
rect 765 27365 783 27381
rect 807 27365 817 27381
rect 817 27365 833 27381
rect 833 27365 863 27381
rect 887 27365 901 27381
rect 901 27365 943 27381
rect 967 27365 969 27381
rect 969 27365 1021 27381
rect 1021 27365 1023 27381
rect 1047 27365 1089 27381
rect 1089 27365 1103 27381
rect 1127 27365 1157 27381
rect 1157 27365 1173 27381
rect 1173 27365 1183 27381
rect 1207 27365 1225 27381
rect 1225 27365 1241 27381
rect 1241 27365 1263 27381
rect 727 27353 783 27365
rect 807 27353 863 27365
rect 887 27353 943 27365
rect 967 27353 1023 27365
rect 1047 27353 1103 27365
rect 1127 27353 1183 27365
rect 1207 27353 1263 27365
rect 727 27325 749 27353
rect 749 27325 765 27353
rect 765 27325 783 27353
rect 807 27325 817 27353
rect 817 27325 833 27353
rect 833 27325 863 27353
rect 887 27325 901 27353
rect 901 27325 943 27353
rect 967 27325 969 27353
rect 969 27325 1021 27353
rect 1021 27325 1023 27353
rect 1047 27325 1089 27353
rect 1089 27325 1103 27353
rect 1127 27325 1157 27353
rect 1157 27325 1173 27353
rect 1173 27325 1183 27353
rect 1207 27325 1225 27353
rect 1225 27325 1241 27353
rect 1241 27325 1263 27353
rect 727 27289 783 27300
rect 807 27289 863 27300
rect 887 27289 943 27300
rect 967 27289 1023 27300
rect 1047 27289 1103 27300
rect 1127 27289 1183 27300
rect 1207 27289 1263 27300
rect 727 27244 749 27289
rect 749 27244 765 27289
rect 765 27244 783 27289
rect 807 27244 817 27289
rect 817 27244 833 27289
rect 833 27244 863 27289
rect 887 27244 901 27289
rect 901 27244 943 27289
rect 967 27244 969 27289
rect 969 27244 1021 27289
rect 1021 27244 1023 27289
rect 1047 27244 1089 27289
rect 1089 27244 1103 27289
rect 1127 27244 1157 27289
rect 1157 27244 1173 27289
rect 1173 27244 1183 27289
rect 1207 27244 1225 27289
rect 1225 27244 1241 27289
rect 1241 27244 1263 27289
rect 727 27173 749 27219
rect 749 27173 765 27219
rect 765 27173 783 27219
rect 807 27173 817 27219
rect 817 27173 833 27219
rect 833 27173 863 27219
rect 887 27173 901 27219
rect 901 27173 943 27219
rect 967 27173 969 27219
rect 969 27173 1021 27219
rect 1021 27173 1023 27219
rect 1047 27173 1089 27219
rect 1089 27173 1103 27219
rect 1127 27173 1157 27219
rect 1157 27173 1173 27219
rect 1173 27173 1183 27219
rect 1207 27173 1225 27219
rect 1225 27173 1241 27219
rect 1241 27173 1263 27219
rect 727 27163 783 27173
rect 807 27163 863 27173
rect 887 27163 943 27173
rect 967 27163 1023 27173
rect 1047 27163 1103 27173
rect 1127 27163 1183 27173
rect 1207 27163 1263 27173
rect 727 27109 749 27138
rect 749 27109 765 27138
rect 765 27109 783 27138
rect 807 27109 817 27138
rect 817 27109 833 27138
rect 833 27109 863 27138
rect 887 27109 901 27138
rect 901 27109 943 27138
rect 967 27109 969 27138
rect 969 27109 1021 27138
rect 1021 27109 1023 27138
rect 1047 27109 1089 27138
rect 1089 27109 1103 27138
rect 1127 27109 1157 27138
rect 1157 27109 1173 27138
rect 1173 27109 1183 27138
rect 1207 27109 1225 27138
rect 1225 27109 1241 27138
rect 1241 27109 1263 27138
rect 727 27097 783 27109
rect 807 27097 863 27109
rect 887 27097 943 27109
rect 967 27097 1023 27109
rect 1047 27097 1103 27109
rect 1127 27097 1183 27109
rect 1207 27097 1263 27109
rect 727 27082 749 27097
rect 749 27082 765 27097
rect 765 27082 783 27097
rect 807 27082 817 27097
rect 817 27082 833 27097
rect 833 27082 863 27097
rect 887 27082 901 27097
rect 901 27082 943 27097
rect 967 27082 969 27097
rect 969 27082 1021 27097
rect 1021 27082 1023 27097
rect 1047 27082 1089 27097
rect 1089 27082 1103 27097
rect 1127 27082 1157 27097
rect 1157 27082 1173 27097
rect 1173 27082 1183 27097
rect 1207 27082 1225 27097
rect 1225 27082 1241 27097
rect 1241 27082 1263 27097
rect 727 27045 749 27057
rect 749 27045 765 27057
rect 765 27045 783 27057
rect 807 27045 817 27057
rect 817 27045 833 27057
rect 833 27045 863 27057
rect 887 27045 901 27057
rect 901 27045 943 27057
rect 967 27045 969 27057
rect 969 27045 1021 27057
rect 1021 27045 1023 27057
rect 1047 27045 1089 27057
rect 1089 27045 1103 27057
rect 1127 27045 1157 27057
rect 1157 27045 1173 27057
rect 1173 27045 1183 27057
rect 1207 27045 1225 27057
rect 1225 27045 1241 27057
rect 1241 27045 1263 27057
rect 727 27033 783 27045
rect 807 27033 863 27045
rect 887 27033 943 27045
rect 967 27033 1023 27045
rect 1047 27033 1103 27045
rect 1127 27033 1183 27045
rect 1207 27033 1263 27045
rect 727 27001 749 27033
rect 749 27001 765 27033
rect 765 27001 783 27033
rect 807 27001 817 27033
rect 817 27001 833 27033
rect 833 27001 863 27033
rect 887 27001 901 27033
rect 901 27001 943 27033
rect 967 27001 969 27033
rect 969 27001 1021 27033
rect 1021 27001 1023 27033
rect 1047 27001 1089 27033
rect 1089 27001 1103 27033
rect 1127 27001 1157 27033
rect 1157 27001 1173 27033
rect 1173 27001 1183 27033
rect 1207 27001 1225 27033
rect 1225 27001 1241 27033
rect 1241 27001 1263 27033
rect 727 26969 783 26976
rect 807 26969 863 26976
rect 887 26969 943 26976
rect 967 26969 1023 26976
rect 1047 26969 1103 26976
rect 1127 26969 1183 26976
rect 1207 26969 1263 26976
rect 727 26920 749 26969
rect 749 26920 765 26969
rect 765 26920 783 26969
rect 807 26920 817 26969
rect 817 26920 833 26969
rect 833 26920 863 26969
rect 887 26920 901 26969
rect 901 26920 943 26969
rect 967 26920 969 26969
rect 969 26920 1021 26969
rect 1021 26920 1023 26969
rect 1047 26920 1089 26969
rect 1089 26920 1103 26969
rect 1127 26920 1157 26969
rect 1157 26920 1173 26969
rect 1173 26920 1183 26969
rect 1207 26920 1225 26969
rect 1225 26920 1241 26969
rect 1241 26920 1263 26969
rect 727 25627 749 25676
rect 749 25627 765 25676
rect 765 25627 817 25676
rect 817 25627 833 25676
rect 833 25627 885 25676
rect 885 25627 901 25676
rect 901 25627 953 25676
rect 953 25627 969 25676
rect 969 25627 1021 25676
rect 1021 25627 1037 25676
rect 1037 25627 1089 25676
rect 1089 25627 1105 25676
rect 1105 25627 1157 25676
rect 1157 25627 1173 25676
rect 1173 25627 1225 25676
rect 1225 25627 1241 25676
rect 1241 25627 1263 25676
rect 727 25615 1263 25627
rect 727 25563 749 25615
rect 749 25563 765 25615
rect 765 25563 817 25615
rect 817 25563 833 25615
rect 833 25563 885 25615
rect 885 25563 901 25615
rect 901 25563 953 25615
rect 953 25563 969 25615
rect 969 25563 1021 25615
rect 1021 25563 1037 25615
rect 1037 25563 1089 25615
rect 1089 25563 1105 25615
rect 1105 25563 1157 25615
rect 1157 25563 1173 25615
rect 1173 25563 1225 25615
rect 1225 25563 1241 25615
rect 1241 25563 1263 25615
rect 727 25551 1263 25563
rect 727 25499 749 25551
rect 749 25499 765 25551
rect 765 25499 817 25551
rect 817 25499 833 25551
rect 833 25499 885 25551
rect 885 25499 901 25551
rect 901 25499 953 25551
rect 953 25499 969 25551
rect 969 25499 1021 25551
rect 1021 25499 1037 25551
rect 1037 25499 1089 25551
rect 1089 25499 1105 25551
rect 1105 25499 1157 25551
rect 1157 25499 1173 25551
rect 1173 25499 1225 25551
rect 1225 25499 1241 25551
rect 1241 25499 1263 25551
rect 727 25487 1263 25499
rect 727 25435 749 25487
rect 749 25435 765 25487
rect 765 25435 817 25487
rect 817 25435 833 25487
rect 833 25435 885 25487
rect 885 25435 901 25487
rect 901 25435 953 25487
rect 953 25435 969 25487
rect 969 25435 1021 25487
rect 1021 25435 1037 25487
rect 1037 25435 1089 25487
rect 1089 25435 1105 25487
rect 1105 25435 1157 25487
rect 1157 25435 1173 25487
rect 1173 25435 1225 25487
rect 1225 25435 1241 25487
rect 1241 25435 1263 25487
rect 727 25423 1263 25435
rect 727 25371 749 25423
rect 749 25371 765 25423
rect 765 25371 817 25423
rect 817 25371 833 25423
rect 833 25371 885 25423
rect 885 25371 901 25423
rect 901 25371 953 25423
rect 953 25371 969 25423
rect 969 25371 1021 25423
rect 1021 25371 1037 25423
rect 1037 25371 1089 25423
rect 1089 25371 1105 25423
rect 1105 25371 1157 25423
rect 1157 25371 1173 25423
rect 1173 25371 1225 25423
rect 1225 25371 1241 25423
rect 1241 25371 1263 25423
rect 727 25359 1263 25371
rect 727 25307 749 25359
rect 749 25307 765 25359
rect 765 25307 817 25359
rect 817 25307 833 25359
rect 833 25307 885 25359
rect 885 25307 901 25359
rect 901 25307 953 25359
rect 953 25307 969 25359
rect 969 25307 1021 25359
rect 1021 25307 1037 25359
rect 1037 25307 1089 25359
rect 1089 25307 1105 25359
rect 1105 25307 1157 25359
rect 1157 25307 1173 25359
rect 1173 25307 1225 25359
rect 1225 25307 1241 25359
rect 1241 25307 1263 25359
rect 727 25295 1263 25307
rect 727 25243 749 25295
rect 749 25243 765 25295
rect 765 25243 817 25295
rect 817 25243 833 25295
rect 833 25243 885 25295
rect 885 25243 901 25295
rect 901 25243 953 25295
rect 953 25243 969 25295
rect 969 25243 1021 25295
rect 1021 25243 1037 25295
rect 1037 25243 1089 25295
rect 1089 25243 1105 25295
rect 1105 25243 1157 25295
rect 1157 25243 1173 25295
rect 1173 25243 1225 25295
rect 1225 25243 1241 25295
rect 1241 25243 1263 25295
rect 727 25231 1263 25243
rect 727 25220 749 25231
rect 749 25220 765 25231
rect 765 25220 817 25231
rect 817 25220 833 25231
rect 833 25220 885 25231
rect 885 25220 901 25231
rect 901 25220 953 25231
rect 953 25220 969 25231
rect 969 25220 1021 25231
rect 1021 25220 1037 25231
rect 1037 25220 1089 25231
rect 1089 25220 1105 25231
rect 1105 25220 1157 25231
rect 1157 25220 1173 25231
rect 1173 25220 1225 25231
rect 1225 25220 1241 25231
rect 1241 25220 1263 25231
rect 727 25179 749 25195
rect 749 25179 765 25195
rect 765 25179 783 25195
rect 807 25179 817 25195
rect 817 25179 833 25195
rect 833 25179 863 25195
rect 887 25179 901 25195
rect 901 25179 943 25195
rect 967 25179 969 25195
rect 969 25179 1021 25195
rect 1021 25179 1023 25195
rect 1047 25179 1089 25195
rect 1089 25179 1103 25195
rect 1127 25179 1157 25195
rect 1157 25179 1173 25195
rect 1173 25179 1183 25195
rect 1207 25179 1225 25195
rect 1225 25179 1241 25195
rect 1241 25179 1263 25195
rect 727 25167 783 25179
rect 807 25167 863 25179
rect 887 25167 943 25179
rect 967 25167 1023 25179
rect 1047 25167 1103 25179
rect 1127 25167 1183 25179
rect 1207 25167 1263 25179
rect 727 25139 749 25167
rect 749 25139 765 25167
rect 765 25139 783 25167
rect 807 25139 817 25167
rect 817 25139 833 25167
rect 833 25139 863 25167
rect 887 25139 901 25167
rect 901 25139 943 25167
rect 967 25139 969 25167
rect 969 25139 1021 25167
rect 1021 25139 1023 25167
rect 1047 25139 1089 25167
rect 1089 25139 1103 25167
rect 1127 25139 1157 25167
rect 1157 25139 1173 25167
rect 1173 25139 1183 25167
rect 1207 25139 1225 25167
rect 1225 25139 1241 25167
rect 1241 25139 1263 25167
rect 727 25103 783 25114
rect 807 25103 863 25114
rect 887 25103 943 25114
rect 967 25103 1023 25114
rect 1047 25103 1103 25114
rect 1127 25103 1183 25114
rect 1207 25103 1263 25114
rect 727 25058 749 25103
rect 749 25058 765 25103
rect 765 25058 783 25103
rect 807 25058 817 25103
rect 817 25058 833 25103
rect 833 25058 863 25103
rect 887 25058 901 25103
rect 901 25058 943 25103
rect 967 25058 969 25103
rect 969 25058 1021 25103
rect 1021 25058 1023 25103
rect 1047 25058 1089 25103
rect 1089 25058 1103 25103
rect 1127 25058 1157 25103
rect 1157 25058 1173 25103
rect 1173 25058 1183 25103
rect 1207 25058 1225 25103
rect 1225 25058 1241 25103
rect 1241 25058 1263 25103
rect 727 24987 749 25033
rect 749 24987 765 25033
rect 765 24987 783 25033
rect 807 24987 817 25033
rect 817 24987 833 25033
rect 833 24987 863 25033
rect 887 24987 901 25033
rect 901 24987 943 25033
rect 967 24987 969 25033
rect 969 24987 1021 25033
rect 1021 24987 1023 25033
rect 1047 24987 1089 25033
rect 1089 24987 1103 25033
rect 1127 24987 1157 25033
rect 1157 24987 1173 25033
rect 1173 24987 1183 25033
rect 1207 24987 1225 25033
rect 1225 24987 1241 25033
rect 1241 24987 1263 25033
rect 727 24977 783 24987
rect 807 24977 863 24987
rect 887 24977 943 24987
rect 967 24977 1023 24987
rect 1047 24977 1103 24987
rect 1127 24977 1183 24987
rect 1207 24977 1263 24987
rect 727 24923 749 24952
rect 749 24923 765 24952
rect 765 24923 783 24952
rect 807 24923 817 24952
rect 817 24923 833 24952
rect 833 24923 863 24952
rect 887 24923 901 24952
rect 901 24923 943 24952
rect 967 24923 969 24952
rect 969 24923 1021 24952
rect 1021 24923 1023 24952
rect 1047 24923 1089 24952
rect 1089 24923 1103 24952
rect 1127 24923 1157 24952
rect 1157 24923 1173 24952
rect 1173 24923 1183 24952
rect 1207 24923 1225 24952
rect 1225 24923 1241 24952
rect 1241 24923 1263 24952
rect 727 24911 783 24923
rect 807 24911 863 24923
rect 887 24911 943 24923
rect 967 24911 1023 24923
rect 1047 24911 1103 24923
rect 1127 24911 1183 24923
rect 1207 24911 1263 24923
rect 727 24896 749 24911
rect 749 24896 765 24911
rect 765 24896 783 24911
rect 807 24896 817 24911
rect 817 24896 833 24911
rect 833 24896 863 24911
rect 887 24896 901 24911
rect 901 24896 943 24911
rect 967 24896 969 24911
rect 969 24896 1021 24911
rect 1021 24896 1023 24911
rect 1047 24896 1089 24911
rect 1089 24896 1103 24911
rect 1127 24896 1157 24911
rect 1157 24896 1173 24911
rect 1173 24896 1183 24911
rect 1207 24896 1225 24911
rect 1225 24896 1241 24911
rect 1241 24896 1263 24911
rect 727 24859 749 24871
rect 749 24859 765 24871
rect 765 24859 783 24871
rect 807 24859 817 24871
rect 817 24859 833 24871
rect 833 24859 863 24871
rect 887 24859 901 24871
rect 901 24859 943 24871
rect 967 24859 969 24871
rect 969 24859 1021 24871
rect 1021 24859 1023 24871
rect 1047 24859 1089 24871
rect 1089 24859 1103 24871
rect 1127 24859 1157 24871
rect 1157 24859 1173 24871
rect 1173 24859 1183 24871
rect 1207 24859 1225 24871
rect 1225 24859 1241 24871
rect 1241 24859 1263 24871
rect 727 24847 783 24859
rect 807 24847 863 24859
rect 887 24847 943 24859
rect 967 24847 1023 24859
rect 1047 24847 1103 24859
rect 1127 24847 1183 24859
rect 1207 24847 1263 24859
rect 727 24815 749 24847
rect 749 24815 765 24847
rect 765 24815 783 24847
rect 807 24815 817 24847
rect 817 24815 833 24847
rect 833 24815 863 24847
rect 887 24815 901 24847
rect 901 24815 943 24847
rect 967 24815 969 24847
rect 969 24815 1021 24847
rect 1021 24815 1023 24847
rect 1047 24815 1089 24847
rect 1089 24815 1103 24847
rect 1127 24815 1157 24847
rect 1157 24815 1173 24847
rect 1173 24815 1183 24847
rect 1207 24815 1225 24847
rect 1225 24815 1241 24847
rect 1241 24815 1263 24847
rect 727 24783 783 24790
rect 807 24783 863 24790
rect 887 24783 943 24790
rect 967 24783 1023 24790
rect 1047 24783 1103 24790
rect 1127 24783 1183 24790
rect 1207 24783 1263 24790
rect 727 24734 749 24783
rect 749 24734 765 24783
rect 765 24734 783 24783
rect 807 24734 817 24783
rect 817 24734 833 24783
rect 833 24734 863 24783
rect 887 24734 901 24783
rect 901 24734 943 24783
rect 967 24734 969 24783
rect 969 24734 1021 24783
rect 1021 24734 1023 24783
rect 1047 24734 1089 24783
rect 1089 24734 1103 24783
rect 1127 24734 1157 24783
rect 1157 24734 1173 24783
rect 1173 24734 1183 24783
rect 1207 24734 1225 24783
rect 1225 24734 1241 24783
rect 1241 24734 1263 24783
rect 727 23479 749 23528
rect 749 23479 765 23528
rect 765 23479 817 23528
rect 817 23479 833 23528
rect 833 23479 885 23528
rect 885 23479 901 23528
rect 901 23479 953 23528
rect 953 23479 969 23528
rect 969 23479 1021 23528
rect 1021 23479 1037 23528
rect 1037 23479 1089 23528
rect 1089 23479 1105 23528
rect 1105 23479 1157 23528
rect 1157 23479 1173 23528
rect 1173 23479 1225 23528
rect 1225 23479 1241 23528
rect 1241 23479 1263 23528
rect 727 23467 1263 23479
rect 727 23415 749 23467
rect 749 23415 765 23467
rect 765 23415 817 23467
rect 817 23415 833 23467
rect 833 23415 885 23467
rect 885 23415 901 23467
rect 901 23415 953 23467
rect 953 23415 969 23467
rect 969 23415 1021 23467
rect 1021 23415 1037 23467
rect 1037 23415 1089 23467
rect 1089 23415 1105 23467
rect 1105 23415 1157 23467
rect 1157 23415 1173 23467
rect 1173 23415 1225 23467
rect 1225 23415 1241 23467
rect 1241 23415 1263 23467
rect 727 23403 1263 23415
rect 727 23351 749 23403
rect 749 23351 765 23403
rect 765 23351 817 23403
rect 817 23351 833 23403
rect 833 23351 885 23403
rect 885 23351 901 23403
rect 901 23351 953 23403
rect 953 23351 969 23403
rect 969 23351 1021 23403
rect 1021 23351 1037 23403
rect 1037 23351 1089 23403
rect 1089 23351 1105 23403
rect 1105 23351 1157 23403
rect 1157 23351 1173 23403
rect 1173 23351 1225 23403
rect 1225 23351 1241 23403
rect 1241 23351 1263 23403
rect 727 23339 1263 23351
rect 727 23287 749 23339
rect 749 23287 765 23339
rect 765 23287 817 23339
rect 817 23287 833 23339
rect 833 23287 885 23339
rect 885 23287 901 23339
rect 901 23287 953 23339
rect 953 23287 969 23339
rect 969 23287 1021 23339
rect 1021 23287 1037 23339
rect 1037 23287 1089 23339
rect 1089 23287 1105 23339
rect 1105 23287 1157 23339
rect 1157 23287 1173 23339
rect 1173 23287 1225 23339
rect 1225 23287 1241 23339
rect 1241 23287 1263 23339
rect 727 23275 1263 23287
rect 727 23223 749 23275
rect 749 23223 765 23275
rect 765 23223 817 23275
rect 817 23223 833 23275
rect 833 23223 885 23275
rect 885 23223 901 23275
rect 901 23223 953 23275
rect 953 23223 969 23275
rect 969 23223 1021 23275
rect 1021 23223 1037 23275
rect 1037 23223 1089 23275
rect 1089 23223 1105 23275
rect 1105 23223 1157 23275
rect 1157 23223 1173 23275
rect 1173 23223 1225 23275
rect 1225 23223 1241 23275
rect 1241 23223 1263 23275
rect 727 23211 1263 23223
rect 727 23159 749 23211
rect 749 23159 765 23211
rect 765 23159 817 23211
rect 817 23159 833 23211
rect 833 23159 885 23211
rect 885 23159 901 23211
rect 901 23159 953 23211
rect 953 23159 969 23211
rect 969 23159 1021 23211
rect 1021 23159 1037 23211
rect 1037 23159 1089 23211
rect 1089 23159 1105 23211
rect 1105 23159 1157 23211
rect 1157 23159 1173 23211
rect 1173 23159 1225 23211
rect 1225 23159 1241 23211
rect 1241 23159 1263 23211
rect 727 23147 1263 23159
rect 727 23095 749 23147
rect 749 23095 765 23147
rect 765 23095 817 23147
rect 817 23095 833 23147
rect 833 23095 885 23147
rect 885 23095 901 23147
rect 901 23095 953 23147
rect 953 23095 969 23147
rect 969 23095 1021 23147
rect 1021 23095 1037 23147
rect 1037 23095 1089 23147
rect 1089 23095 1105 23147
rect 1105 23095 1157 23147
rect 1157 23095 1173 23147
rect 1173 23095 1225 23147
rect 1225 23095 1241 23147
rect 1241 23095 1263 23147
rect 727 23083 1263 23095
rect 727 23072 749 23083
rect 749 23072 765 23083
rect 765 23072 817 23083
rect 817 23072 833 23083
rect 833 23072 885 23083
rect 885 23072 901 23083
rect 901 23072 953 23083
rect 953 23072 969 23083
rect 969 23072 1021 23083
rect 1021 23072 1037 23083
rect 1037 23072 1089 23083
rect 1089 23072 1105 23083
rect 1105 23072 1157 23083
rect 1157 23072 1173 23083
rect 1173 23072 1225 23083
rect 1225 23072 1241 23083
rect 1241 23072 1263 23083
rect 727 23031 749 23047
rect 749 23031 765 23047
rect 765 23031 783 23047
rect 807 23031 817 23047
rect 817 23031 833 23047
rect 833 23031 863 23047
rect 887 23031 901 23047
rect 901 23031 943 23047
rect 967 23031 969 23047
rect 969 23031 1021 23047
rect 1021 23031 1023 23047
rect 1047 23031 1089 23047
rect 1089 23031 1103 23047
rect 1127 23031 1157 23047
rect 1157 23031 1173 23047
rect 1173 23031 1183 23047
rect 1207 23031 1225 23047
rect 1225 23031 1241 23047
rect 1241 23031 1263 23047
rect 727 23019 783 23031
rect 807 23019 863 23031
rect 887 23019 943 23031
rect 967 23019 1023 23031
rect 1047 23019 1103 23031
rect 1127 23019 1183 23031
rect 1207 23019 1263 23031
rect 727 22991 749 23019
rect 749 22991 765 23019
rect 765 22991 783 23019
rect 807 22991 817 23019
rect 817 22991 833 23019
rect 833 22991 863 23019
rect 887 22991 901 23019
rect 901 22991 943 23019
rect 967 22991 969 23019
rect 969 22991 1021 23019
rect 1021 22991 1023 23019
rect 1047 22991 1089 23019
rect 1089 22991 1103 23019
rect 1127 22991 1157 23019
rect 1157 22991 1173 23019
rect 1173 22991 1183 23019
rect 1207 22991 1225 23019
rect 1225 22991 1241 23019
rect 1241 22991 1263 23019
rect 727 22955 783 22966
rect 807 22955 863 22966
rect 887 22955 943 22966
rect 967 22955 1023 22966
rect 1047 22955 1103 22966
rect 1127 22955 1183 22966
rect 1207 22955 1263 22966
rect 727 22910 749 22955
rect 749 22910 765 22955
rect 765 22910 783 22955
rect 807 22910 817 22955
rect 817 22910 833 22955
rect 833 22910 863 22955
rect 887 22910 901 22955
rect 901 22910 943 22955
rect 967 22910 969 22955
rect 969 22910 1021 22955
rect 1021 22910 1023 22955
rect 1047 22910 1089 22955
rect 1089 22910 1103 22955
rect 1127 22910 1157 22955
rect 1157 22910 1173 22955
rect 1173 22910 1183 22955
rect 1207 22910 1225 22955
rect 1225 22910 1241 22955
rect 1241 22910 1263 22955
rect 727 22839 749 22885
rect 749 22839 765 22885
rect 765 22839 783 22885
rect 807 22839 817 22885
rect 817 22839 833 22885
rect 833 22839 863 22885
rect 887 22839 901 22885
rect 901 22839 943 22885
rect 967 22839 969 22885
rect 969 22839 1021 22885
rect 1021 22839 1023 22885
rect 1047 22839 1089 22885
rect 1089 22839 1103 22885
rect 1127 22839 1157 22885
rect 1157 22839 1173 22885
rect 1173 22839 1183 22885
rect 1207 22839 1225 22885
rect 1225 22839 1241 22885
rect 1241 22839 1263 22885
rect 727 22829 783 22839
rect 807 22829 863 22839
rect 887 22829 943 22839
rect 967 22829 1023 22839
rect 1047 22829 1103 22839
rect 1127 22829 1183 22839
rect 1207 22829 1263 22839
rect 727 22775 749 22804
rect 749 22775 765 22804
rect 765 22775 783 22804
rect 807 22775 817 22804
rect 817 22775 833 22804
rect 833 22775 863 22804
rect 887 22775 901 22804
rect 901 22775 943 22804
rect 967 22775 969 22804
rect 969 22775 1021 22804
rect 1021 22775 1023 22804
rect 1047 22775 1089 22804
rect 1089 22775 1103 22804
rect 1127 22775 1157 22804
rect 1157 22775 1173 22804
rect 1173 22775 1183 22804
rect 1207 22775 1225 22804
rect 1225 22775 1241 22804
rect 1241 22775 1263 22804
rect 727 22763 783 22775
rect 807 22763 863 22775
rect 887 22763 943 22775
rect 967 22763 1023 22775
rect 1047 22763 1103 22775
rect 1127 22763 1183 22775
rect 1207 22763 1263 22775
rect 727 22748 749 22763
rect 749 22748 765 22763
rect 765 22748 783 22763
rect 807 22748 817 22763
rect 817 22748 833 22763
rect 833 22748 863 22763
rect 887 22748 901 22763
rect 901 22748 943 22763
rect 967 22748 969 22763
rect 969 22748 1021 22763
rect 1021 22748 1023 22763
rect 1047 22748 1089 22763
rect 1089 22748 1103 22763
rect 1127 22748 1157 22763
rect 1157 22748 1173 22763
rect 1173 22748 1183 22763
rect 1207 22748 1225 22763
rect 1225 22748 1241 22763
rect 1241 22748 1263 22763
rect 727 22711 749 22723
rect 749 22711 765 22723
rect 765 22711 783 22723
rect 807 22711 817 22723
rect 817 22711 833 22723
rect 833 22711 863 22723
rect 887 22711 901 22723
rect 901 22711 943 22723
rect 967 22711 969 22723
rect 969 22711 1021 22723
rect 1021 22711 1023 22723
rect 1047 22711 1089 22723
rect 1089 22711 1103 22723
rect 1127 22711 1157 22723
rect 1157 22711 1173 22723
rect 1173 22711 1183 22723
rect 1207 22711 1225 22723
rect 1225 22711 1241 22723
rect 1241 22711 1263 22723
rect 727 22699 783 22711
rect 807 22699 863 22711
rect 887 22699 943 22711
rect 967 22699 1023 22711
rect 1047 22699 1103 22711
rect 1127 22699 1183 22711
rect 1207 22699 1263 22711
rect 727 22667 749 22699
rect 749 22667 765 22699
rect 765 22667 783 22699
rect 807 22667 817 22699
rect 817 22667 833 22699
rect 833 22667 863 22699
rect 887 22667 901 22699
rect 901 22667 943 22699
rect 967 22667 969 22699
rect 969 22667 1021 22699
rect 1021 22667 1023 22699
rect 1047 22667 1089 22699
rect 1089 22667 1103 22699
rect 1127 22667 1157 22699
rect 1157 22667 1173 22699
rect 1173 22667 1183 22699
rect 1207 22667 1225 22699
rect 1225 22667 1241 22699
rect 1241 22667 1263 22699
rect 727 22635 783 22642
rect 807 22635 863 22642
rect 887 22635 943 22642
rect 967 22635 1023 22642
rect 1047 22635 1103 22642
rect 1127 22635 1183 22642
rect 1207 22635 1263 22642
rect 727 22586 749 22635
rect 749 22586 765 22635
rect 765 22586 783 22635
rect 807 22586 817 22635
rect 817 22586 833 22635
rect 833 22586 863 22635
rect 887 22586 901 22635
rect 901 22586 943 22635
rect 967 22586 969 22635
rect 969 22586 1021 22635
rect 1021 22586 1023 22635
rect 1047 22586 1089 22635
rect 1089 22586 1103 22635
rect 1127 22586 1157 22635
rect 1157 22586 1173 22635
rect 1173 22586 1183 22635
rect 1207 22586 1225 22635
rect 1225 22586 1241 22635
rect 1241 22586 1263 22635
rect 727 21309 749 21358
rect 749 21309 765 21358
rect 765 21309 817 21358
rect 817 21309 833 21358
rect 833 21309 885 21358
rect 885 21309 901 21358
rect 901 21309 953 21358
rect 953 21309 969 21358
rect 969 21309 1021 21358
rect 1021 21309 1037 21358
rect 1037 21309 1089 21358
rect 1089 21309 1105 21358
rect 1105 21309 1157 21358
rect 1157 21309 1173 21358
rect 1173 21309 1225 21358
rect 1225 21309 1241 21358
rect 1241 21309 1263 21358
rect 727 21297 1263 21309
rect 727 21245 749 21297
rect 749 21245 765 21297
rect 765 21245 817 21297
rect 817 21245 833 21297
rect 833 21245 885 21297
rect 885 21245 901 21297
rect 901 21245 953 21297
rect 953 21245 969 21297
rect 969 21245 1021 21297
rect 1021 21245 1037 21297
rect 1037 21245 1089 21297
rect 1089 21245 1105 21297
rect 1105 21245 1157 21297
rect 1157 21245 1173 21297
rect 1173 21245 1225 21297
rect 1225 21245 1241 21297
rect 1241 21245 1263 21297
rect 727 21233 1263 21245
rect 727 21181 749 21233
rect 749 21181 765 21233
rect 765 21181 817 21233
rect 817 21181 833 21233
rect 833 21181 885 21233
rect 885 21181 901 21233
rect 901 21181 953 21233
rect 953 21181 969 21233
rect 969 21181 1021 21233
rect 1021 21181 1037 21233
rect 1037 21181 1089 21233
rect 1089 21181 1105 21233
rect 1105 21181 1157 21233
rect 1157 21181 1173 21233
rect 1173 21181 1225 21233
rect 1225 21181 1241 21233
rect 1241 21181 1263 21233
rect 727 21169 1263 21181
rect 727 21117 749 21169
rect 749 21117 765 21169
rect 765 21117 817 21169
rect 817 21117 833 21169
rect 833 21117 885 21169
rect 885 21117 901 21169
rect 901 21117 953 21169
rect 953 21117 969 21169
rect 969 21117 1021 21169
rect 1021 21117 1037 21169
rect 1037 21117 1089 21169
rect 1089 21117 1105 21169
rect 1105 21117 1157 21169
rect 1157 21117 1173 21169
rect 1173 21117 1225 21169
rect 1225 21117 1241 21169
rect 1241 21117 1263 21169
rect 727 21105 1263 21117
rect 727 21053 749 21105
rect 749 21053 765 21105
rect 765 21053 817 21105
rect 817 21053 833 21105
rect 833 21053 885 21105
rect 885 21053 901 21105
rect 901 21053 953 21105
rect 953 21053 969 21105
rect 969 21053 1021 21105
rect 1021 21053 1037 21105
rect 1037 21053 1089 21105
rect 1089 21053 1105 21105
rect 1105 21053 1157 21105
rect 1157 21053 1173 21105
rect 1173 21053 1225 21105
rect 1225 21053 1241 21105
rect 1241 21053 1263 21105
rect 727 21041 1263 21053
rect 727 20989 749 21041
rect 749 20989 765 21041
rect 765 20989 817 21041
rect 817 20989 833 21041
rect 833 20989 885 21041
rect 885 20989 901 21041
rect 901 20989 953 21041
rect 953 20989 969 21041
rect 969 20989 1021 21041
rect 1021 20989 1037 21041
rect 1037 20989 1089 21041
rect 1089 20989 1105 21041
rect 1105 20989 1157 21041
rect 1157 20989 1173 21041
rect 1173 20989 1225 21041
rect 1225 20989 1241 21041
rect 1241 20989 1263 21041
rect 727 20977 1263 20989
rect 727 20925 749 20977
rect 749 20925 765 20977
rect 765 20925 817 20977
rect 817 20925 833 20977
rect 833 20925 885 20977
rect 885 20925 901 20977
rect 901 20925 953 20977
rect 953 20925 969 20977
rect 969 20925 1021 20977
rect 1021 20925 1037 20977
rect 1037 20925 1089 20977
rect 1089 20925 1105 20977
rect 1105 20925 1157 20977
rect 1157 20925 1173 20977
rect 1173 20925 1225 20977
rect 1225 20925 1241 20977
rect 1241 20925 1263 20977
rect 727 20913 1263 20925
rect 727 20902 749 20913
rect 749 20902 765 20913
rect 765 20902 817 20913
rect 817 20902 833 20913
rect 833 20902 885 20913
rect 885 20902 901 20913
rect 901 20902 953 20913
rect 953 20902 969 20913
rect 969 20902 1021 20913
rect 1021 20902 1037 20913
rect 1037 20902 1089 20913
rect 1089 20902 1105 20913
rect 1105 20902 1157 20913
rect 1157 20902 1173 20913
rect 1173 20902 1225 20913
rect 1225 20902 1241 20913
rect 1241 20902 1263 20913
rect 727 20861 749 20877
rect 749 20861 765 20877
rect 765 20861 783 20877
rect 807 20861 817 20877
rect 817 20861 833 20877
rect 833 20861 863 20877
rect 887 20861 901 20877
rect 901 20861 943 20877
rect 967 20861 969 20877
rect 969 20861 1021 20877
rect 1021 20861 1023 20877
rect 1047 20861 1089 20877
rect 1089 20861 1103 20877
rect 1127 20861 1157 20877
rect 1157 20861 1173 20877
rect 1173 20861 1183 20877
rect 1207 20861 1225 20877
rect 1225 20861 1241 20877
rect 1241 20861 1263 20877
rect 727 20849 783 20861
rect 807 20849 863 20861
rect 887 20849 943 20861
rect 967 20849 1023 20861
rect 1047 20849 1103 20861
rect 1127 20849 1183 20861
rect 1207 20849 1263 20861
rect 727 20821 749 20849
rect 749 20821 765 20849
rect 765 20821 783 20849
rect 807 20821 817 20849
rect 817 20821 833 20849
rect 833 20821 863 20849
rect 887 20821 901 20849
rect 901 20821 943 20849
rect 967 20821 969 20849
rect 969 20821 1021 20849
rect 1021 20821 1023 20849
rect 1047 20821 1089 20849
rect 1089 20821 1103 20849
rect 1127 20821 1157 20849
rect 1157 20821 1173 20849
rect 1173 20821 1183 20849
rect 1207 20821 1225 20849
rect 1225 20821 1241 20849
rect 1241 20821 1263 20849
rect 727 20785 783 20796
rect 807 20785 863 20796
rect 887 20785 943 20796
rect 967 20785 1023 20796
rect 1047 20785 1103 20796
rect 1127 20785 1183 20796
rect 1207 20785 1263 20796
rect 727 20740 749 20785
rect 749 20740 765 20785
rect 765 20740 783 20785
rect 807 20740 817 20785
rect 817 20740 833 20785
rect 833 20740 863 20785
rect 887 20740 901 20785
rect 901 20740 943 20785
rect 967 20740 969 20785
rect 969 20740 1021 20785
rect 1021 20740 1023 20785
rect 1047 20740 1089 20785
rect 1089 20740 1103 20785
rect 1127 20740 1157 20785
rect 1157 20740 1173 20785
rect 1173 20740 1183 20785
rect 1207 20740 1225 20785
rect 1225 20740 1241 20785
rect 1241 20740 1263 20785
rect 727 20669 749 20715
rect 749 20669 765 20715
rect 765 20669 783 20715
rect 807 20669 817 20715
rect 817 20669 833 20715
rect 833 20669 863 20715
rect 887 20669 901 20715
rect 901 20669 943 20715
rect 967 20669 969 20715
rect 969 20669 1021 20715
rect 1021 20669 1023 20715
rect 1047 20669 1089 20715
rect 1089 20669 1103 20715
rect 1127 20669 1157 20715
rect 1157 20669 1173 20715
rect 1173 20669 1183 20715
rect 1207 20669 1225 20715
rect 1225 20669 1241 20715
rect 1241 20669 1263 20715
rect 727 20659 783 20669
rect 807 20659 863 20669
rect 887 20659 943 20669
rect 967 20659 1023 20669
rect 1047 20659 1103 20669
rect 1127 20659 1183 20669
rect 1207 20659 1263 20669
rect 727 20605 749 20634
rect 749 20605 765 20634
rect 765 20605 783 20634
rect 807 20605 817 20634
rect 817 20605 833 20634
rect 833 20605 863 20634
rect 887 20605 901 20634
rect 901 20605 943 20634
rect 967 20605 969 20634
rect 969 20605 1021 20634
rect 1021 20605 1023 20634
rect 1047 20605 1089 20634
rect 1089 20605 1103 20634
rect 1127 20605 1157 20634
rect 1157 20605 1173 20634
rect 1173 20605 1183 20634
rect 1207 20605 1225 20634
rect 1225 20605 1241 20634
rect 1241 20605 1263 20634
rect 727 20593 783 20605
rect 807 20593 863 20605
rect 887 20593 943 20605
rect 967 20593 1023 20605
rect 1047 20593 1103 20605
rect 1127 20593 1183 20605
rect 1207 20593 1263 20605
rect 727 20578 749 20593
rect 749 20578 765 20593
rect 765 20578 783 20593
rect 807 20578 817 20593
rect 817 20578 833 20593
rect 833 20578 863 20593
rect 887 20578 901 20593
rect 901 20578 943 20593
rect 967 20578 969 20593
rect 969 20578 1021 20593
rect 1021 20578 1023 20593
rect 1047 20578 1089 20593
rect 1089 20578 1103 20593
rect 1127 20578 1157 20593
rect 1157 20578 1173 20593
rect 1173 20578 1183 20593
rect 1207 20578 1225 20593
rect 1225 20578 1241 20593
rect 1241 20578 1263 20593
rect 727 20541 749 20553
rect 749 20541 765 20553
rect 765 20541 783 20553
rect 807 20541 817 20553
rect 817 20541 833 20553
rect 833 20541 863 20553
rect 887 20541 901 20553
rect 901 20541 943 20553
rect 967 20541 969 20553
rect 969 20541 1021 20553
rect 1021 20541 1023 20553
rect 1047 20541 1089 20553
rect 1089 20541 1103 20553
rect 1127 20541 1157 20553
rect 1157 20541 1173 20553
rect 1173 20541 1183 20553
rect 1207 20541 1225 20553
rect 1225 20541 1241 20553
rect 1241 20541 1263 20553
rect 727 20529 783 20541
rect 807 20529 863 20541
rect 887 20529 943 20541
rect 967 20529 1023 20541
rect 1047 20529 1103 20541
rect 1127 20529 1183 20541
rect 1207 20529 1263 20541
rect 727 20497 749 20529
rect 749 20497 765 20529
rect 765 20497 783 20529
rect 807 20497 817 20529
rect 817 20497 833 20529
rect 833 20497 863 20529
rect 887 20497 901 20529
rect 901 20497 943 20529
rect 967 20497 969 20529
rect 969 20497 1021 20529
rect 1021 20497 1023 20529
rect 1047 20497 1089 20529
rect 1089 20497 1103 20529
rect 1127 20497 1157 20529
rect 1157 20497 1173 20529
rect 1173 20497 1183 20529
rect 1207 20497 1225 20529
rect 1225 20497 1241 20529
rect 1241 20497 1263 20529
rect 727 20465 783 20472
rect 807 20465 863 20472
rect 887 20465 943 20472
rect 967 20465 1023 20472
rect 1047 20465 1103 20472
rect 1127 20465 1183 20472
rect 1207 20465 1263 20472
rect 727 20416 749 20465
rect 749 20416 765 20465
rect 765 20416 783 20465
rect 807 20416 817 20465
rect 817 20416 833 20465
rect 833 20416 863 20465
rect 887 20416 901 20465
rect 901 20416 943 20465
rect 967 20416 969 20465
rect 969 20416 1021 20465
rect 1021 20416 1023 20465
rect 1047 20416 1089 20465
rect 1089 20416 1103 20465
rect 1127 20416 1157 20465
rect 1157 20416 1173 20465
rect 1173 20416 1183 20465
rect 1207 20416 1225 20465
rect 1225 20416 1241 20465
rect 1241 20416 1263 20465
rect 727 19205 749 19254
rect 749 19205 765 19254
rect 765 19205 817 19254
rect 817 19205 833 19254
rect 833 19205 885 19254
rect 885 19205 901 19254
rect 901 19205 953 19254
rect 953 19205 969 19254
rect 969 19205 1021 19254
rect 1021 19205 1037 19254
rect 1037 19205 1089 19254
rect 1089 19205 1105 19254
rect 1105 19205 1157 19254
rect 1157 19205 1173 19254
rect 1173 19205 1225 19254
rect 1225 19205 1241 19254
rect 1241 19205 1263 19254
rect 727 19193 1263 19205
rect 727 19141 749 19193
rect 749 19141 765 19193
rect 765 19141 817 19193
rect 817 19141 833 19193
rect 833 19141 885 19193
rect 885 19141 901 19193
rect 901 19141 953 19193
rect 953 19141 969 19193
rect 969 19141 1021 19193
rect 1021 19141 1037 19193
rect 1037 19141 1089 19193
rect 1089 19141 1105 19193
rect 1105 19141 1157 19193
rect 1157 19141 1173 19193
rect 1173 19141 1225 19193
rect 1225 19141 1241 19193
rect 1241 19141 1263 19193
rect 727 19129 1263 19141
rect 727 19077 749 19129
rect 749 19077 765 19129
rect 765 19077 817 19129
rect 817 19077 833 19129
rect 833 19077 885 19129
rect 885 19077 901 19129
rect 901 19077 953 19129
rect 953 19077 969 19129
rect 969 19077 1021 19129
rect 1021 19077 1037 19129
rect 1037 19077 1089 19129
rect 1089 19077 1105 19129
rect 1105 19077 1157 19129
rect 1157 19077 1173 19129
rect 1173 19077 1225 19129
rect 1225 19077 1241 19129
rect 1241 19077 1263 19129
rect 727 19065 1263 19077
rect 727 19013 749 19065
rect 749 19013 765 19065
rect 765 19013 817 19065
rect 817 19013 833 19065
rect 833 19013 885 19065
rect 885 19013 901 19065
rect 901 19013 953 19065
rect 953 19013 969 19065
rect 969 19013 1021 19065
rect 1021 19013 1037 19065
rect 1037 19013 1089 19065
rect 1089 19013 1105 19065
rect 1105 19013 1157 19065
rect 1157 19013 1173 19065
rect 1173 19013 1225 19065
rect 1225 19013 1241 19065
rect 1241 19013 1263 19065
rect 727 19001 1263 19013
rect 727 18949 749 19001
rect 749 18949 765 19001
rect 765 18949 817 19001
rect 817 18949 833 19001
rect 833 18949 885 19001
rect 885 18949 901 19001
rect 901 18949 953 19001
rect 953 18949 969 19001
rect 969 18949 1021 19001
rect 1021 18949 1037 19001
rect 1037 18949 1089 19001
rect 1089 18949 1105 19001
rect 1105 18949 1157 19001
rect 1157 18949 1173 19001
rect 1173 18949 1225 19001
rect 1225 18949 1241 19001
rect 1241 18949 1263 19001
rect 727 18937 1263 18949
rect 727 18885 749 18937
rect 749 18885 765 18937
rect 765 18885 817 18937
rect 817 18885 833 18937
rect 833 18885 885 18937
rect 885 18885 901 18937
rect 901 18885 953 18937
rect 953 18885 969 18937
rect 969 18885 1021 18937
rect 1021 18885 1037 18937
rect 1037 18885 1089 18937
rect 1089 18885 1105 18937
rect 1105 18885 1157 18937
rect 1157 18885 1173 18937
rect 1173 18885 1225 18937
rect 1225 18885 1241 18937
rect 1241 18885 1263 18937
rect 727 18873 1263 18885
rect 727 18821 749 18873
rect 749 18821 765 18873
rect 765 18821 817 18873
rect 817 18821 833 18873
rect 833 18821 885 18873
rect 885 18821 901 18873
rect 901 18821 953 18873
rect 953 18821 969 18873
rect 969 18821 1021 18873
rect 1021 18821 1037 18873
rect 1037 18821 1089 18873
rect 1089 18821 1105 18873
rect 1105 18821 1157 18873
rect 1157 18821 1173 18873
rect 1173 18821 1225 18873
rect 1225 18821 1241 18873
rect 1241 18821 1263 18873
rect 727 18809 1263 18821
rect 727 18798 749 18809
rect 749 18798 765 18809
rect 765 18798 817 18809
rect 817 18798 833 18809
rect 833 18798 885 18809
rect 885 18798 901 18809
rect 901 18798 953 18809
rect 953 18798 969 18809
rect 969 18798 1021 18809
rect 1021 18798 1037 18809
rect 1037 18798 1089 18809
rect 1089 18798 1105 18809
rect 1105 18798 1157 18809
rect 1157 18798 1173 18809
rect 1173 18798 1225 18809
rect 1225 18798 1241 18809
rect 1241 18798 1263 18809
rect 727 18757 749 18773
rect 749 18757 765 18773
rect 765 18757 783 18773
rect 807 18757 817 18773
rect 817 18757 833 18773
rect 833 18757 863 18773
rect 887 18757 901 18773
rect 901 18757 943 18773
rect 967 18757 969 18773
rect 969 18757 1021 18773
rect 1021 18757 1023 18773
rect 1047 18757 1089 18773
rect 1089 18757 1103 18773
rect 1127 18757 1157 18773
rect 1157 18757 1173 18773
rect 1173 18757 1183 18773
rect 1207 18757 1225 18773
rect 1225 18757 1241 18773
rect 1241 18757 1263 18773
rect 727 18745 783 18757
rect 807 18745 863 18757
rect 887 18745 943 18757
rect 967 18745 1023 18757
rect 1047 18745 1103 18757
rect 1127 18745 1183 18757
rect 1207 18745 1263 18757
rect 727 18717 749 18745
rect 749 18717 765 18745
rect 765 18717 783 18745
rect 807 18717 817 18745
rect 817 18717 833 18745
rect 833 18717 863 18745
rect 887 18717 901 18745
rect 901 18717 943 18745
rect 967 18717 969 18745
rect 969 18717 1021 18745
rect 1021 18717 1023 18745
rect 1047 18717 1089 18745
rect 1089 18717 1103 18745
rect 1127 18717 1157 18745
rect 1157 18717 1173 18745
rect 1173 18717 1183 18745
rect 1207 18717 1225 18745
rect 1225 18717 1241 18745
rect 1241 18717 1263 18745
rect 727 18681 783 18692
rect 807 18681 863 18692
rect 887 18681 943 18692
rect 967 18681 1023 18692
rect 1047 18681 1103 18692
rect 1127 18681 1183 18692
rect 1207 18681 1263 18692
rect 727 18636 749 18681
rect 749 18636 765 18681
rect 765 18636 783 18681
rect 807 18636 817 18681
rect 817 18636 833 18681
rect 833 18636 863 18681
rect 887 18636 901 18681
rect 901 18636 943 18681
rect 967 18636 969 18681
rect 969 18636 1021 18681
rect 1021 18636 1023 18681
rect 1047 18636 1089 18681
rect 1089 18636 1103 18681
rect 1127 18636 1157 18681
rect 1157 18636 1173 18681
rect 1173 18636 1183 18681
rect 1207 18636 1225 18681
rect 1225 18636 1241 18681
rect 1241 18636 1263 18681
rect 727 18565 749 18611
rect 749 18565 765 18611
rect 765 18565 783 18611
rect 807 18565 817 18611
rect 817 18565 833 18611
rect 833 18565 863 18611
rect 887 18565 901 18611
rect 901 18565 943 18611
rect 967 18565 969 18611
rect 969 18565 1021 18611
rect 1021 18565 1023 18611
rect 1047 18565 1089 18611
rect 1089 18565 1103 18611
rect 1127 18565 1157 18611
rect 1157 18565 1173 18611
rect 1173 18565 1183 18611
rect 1207 18565 1225 18611
rect 1225 18565 1241 18611
rect 1241 18565 1263 18611
rect 727 18555 783 18565
rect 807 18555 863 18565
rect 887 18555 943 18565
rect 967 18555 1023 18565
rect 1047 18555 1103 18565
rect 1127 18555 1183 18565
rect 1207 18555 1263 18565
rect 727 18501 749 18530
rect 749 18501 765 18530
rect 765 18501 783 18530
rect 807 18501 817 18530
rect 817 18501 833 18530
rect 833 18501 863 18530
rect 887 18501 901 18530
rect 901 18501 943 18530
rect 967 18501 969 18530
rect 969 18501 1021 18530
rect 1021 18501 1023 18530
rect 1047 18501 1089 18530
rect 1089 18501 1103 18530
rect 1127 18501 1157 18530
rect 1157 18501 1173 18530
rect 1173 18501 1183 18530
rect 1207 18501 1225 18530
rect 1225 18501 1241 18530
rect 1241 18501 1263 18530
rect 727 18489 783 18501
rect 807 18489 863 18501
rect 887 18489 943 18501
rect 967 18489 1023 18501
rect 1047 18489 1103 18501
rect 1127 18489 1183 18501
rect 1207 18489 1263 18501
rect 727 18474 749 18489
rect 749 18474 765 18489
rect 765 18474 783 18489
rect 807 18474 817 18489
rect 817 18474 833 18489
rect 833 18474 863 18489
rect 887 18474 901 18489
rect 901 18474 943 18489
rect 967 18474 969 18489
rect 969 18474 1021 18489
rect 1021 18474 1023 18489
rect 1047 18474 1089 18489
rect 1089 18474 1103 18489
rect 1127 18474 1157 18489
rect 1157 18474 1173 18489
rect 1173 18474 1183 18489
rect 1207 18474 1225 18489
rect 1225 18474 1241 18489
rect 1241 18474 1263 18489
rect 727 18437 749 18449
rect 749 18437 765 18449
rect 765 18437 783 18449
rect 807 18437 817 18449
rect 817 18437 833 18449
rect 833 18437 863 18449
rect 887 18437 901 18449
rect 901 18437 943 18449
rect 967 18437 969 18449
rect 969 18437 1021 18449
rect 1021 18437 1023 18449
rect 1047 18437 1089 18449
rect 1089 18437 1103 18449
rect 1127 18437 1157 18449
rect 1157 18437 1173 18449
rect 1173 18437 1183 18449
rect 1207 18437 1225 18449
rect 1225 18437 1241 18449
rect 1241 18437 1263 18449
rect 727 18425 783 18437
rect 807 18425 863 18437
rect 887 18425 943 18437
rect 967 18425 1023 18437
rect 1047 18425 1103 18437
rect 1127 18425 1183 18437
rect 1207 18425 1263 18437
rect 727 18393 749 18425
rect 749 18393 765 18425
rect 765 18393 783 18425
rect 807 18393 817 18425
rect 817 18393 833 18425
rect 833 18393 863 18425
rect 887 18393 901 18425
rect 901 18393 943 18425
rect 967 18393 969 18425
rect 969 18393 1021 18425
rect 1021 18393 1023 18425
rect 1047 18393 1089 18425
rect 1089 18393 1103 18425
rect 1127 18393 1157 18425
rect 1157 18393 1173 18425
rect 1173 18393 1183 18425
rect 1207 18393 1225 18425
rect 1225 18393 1241 18425
rect 1241 18393 1263 18425
rect 727 18361 783 18368
rect 807 18361 863 18368
rect 887 18361 943 18368
rect 967 18361 1023 18368
rect 1047 18361 1103 18368
rect 1127 18361 1183 18368
rect 1207 18361 1263 18368
rect 727 18312 749 18361
rect 749 18312 765 18361
rect 765 18312 783 18361
rect 807 18312 817 18361
rect 817 18312 833 18361
rect 833 18312 863 18361
rect 887 18312 901 18361
rect 901 18312 943 18361
rect 967 18312 969 18361
rect 969 18312 1021 18361
rect 1021 18312 1023 18361
rect 1047 18312 1089 18361
rect 1089 18312 1103 18361
rect 1127 18312 1157 18361
rect 1157 18312 1173 18361
rect 1173 18312 1183 18361
rect 1207 18312 1225 18361
rect 1225 18312 1241 18361
rect 1241 18312 1263 18361
rect 727 17094 749 17143
rect 749 17094 765 17143
rect 765 17094 817 17143
rect 817 17094 833 17143
rect 833 17094 885 17143
rect 885 17094 901 17143
rect 901 17094 953 17143
rect 953 17094 969 17143
rect 969 17094 1021 17143
rect 1021 17094 1037 17143
rect 1037 17094 1089 17143
rect 1089 17094 1105 17143
rect 1105 17094 1157 17143
rect 1157 17094 1173 17143
rect 1173 17094 1225 17143
rect 1225 17094 1241 17143
rect 1241 17094 1263 17143
rect 727 17082 1263 17094
rect 727 17030 749 17082
rect 749 17030 765 17082
rect 765 17030 817 17082
rect 817 17030 833 17082
rect 833 17030 885 17082
rect 885 17030 901 17082
rect 901 17030 953 17082
rect 953 17030 969 17082
rect 969 17030 1021 17082
rect 1021 17030 1037 17082
rect 1037 17030 1089 17082
rect 1089 17030 1105 17082
rect 1105 17030 1157 17082
rect 1157 17030 1173 17082
rect 1173 17030 1225 17082
rect 1225 17030 1241 17082
rect 1241 17030 1263 17082
rect 727 17018 1263 17030
rect 727 16966 749 17018
rect 749 16966 765 17018
rect 765 16966 817 17018
rect 817 16966 833 17018
rect 833 16966 885 17018
rect 885 16966 901 17018
rect 901 16966 953 17018
rect 953 16966 969 17018
rect 969 16966 1021 17018
rect 1021 16966 1037 17018
rect 1037 16966 1089 17018
rect 1089 16966 1105 17018
rect 1105 16966 1157 17018
rect 1157 16966 1173 17018
rect 1173 16966 1225 17018
rect 1225 16966 1241 17018
rect 1241 16966 1263 17018
rect 727 16954 1263 16966
rect 727 16902 749 16954
rect 749 16902 765 16954
rect 765 16902 817 16954
rect 817 16902 833 16954
rect 833 16902 885 16954
rect 885 16902 901 16954
rect 901 16902 953 16954
rect 953 16902 969 16954
rect 969 16902 1021 16954
rect 1021 16902 1037 16954
rect 1037 16902 1089 16954
rect 1089 16902 1105 16954
rect 1105 16902 1157 16954
rect 1157 16902 1173 16954
rect 1173 16902 1225 16954
rect 1225 16902 1241 16954
rect 1241 16902 1263 16954
rect 727 16890 1263 16902
rect 727 16838 749 16890
rect 749 16838 765 16890
rect 765 16838 817 16890
rect 817 16838 833 16890
rect 833 16838 885 16890
rect 885 16838 901 16890
rect 901 16838 953 16890
rect 953 16838 969 16890
rect 969 16838 1021 16890
rect 1021 16838 1037 16890
rect 1037 16838 1089 16890
rect 1089 16838 1105 16890
rect 1105 16838 1157 16890
rect 1157 16838 1173 16890
rect 1173 16838 1225 16890
rect 1225 16838 1241 16890
rect 1241 16838 1263 16890
rect 727 16826 1263 16838
rect 727 16774 749 16826
rect 749 16774 765 16826
rect 765 16774 817 16826
rect 817 16774 833 16826
rect 833 16774 885 16826
rect 885 16774 901 16826
rect 901 16774 953 16826
rect 953 16774 969 16826
rect 969 16774 1021 16826
rect 1021 16774 1037 16826
rect 1037 16774 1089 16826
rect 1089 16774 1105 16826
rect 1105 16774 1157 16826
rect 1157 16774 1173 16826
rect 1173 16774 1225 16826
rect 1225 16774 1241 16826
rect 1241 16774 1263 16826
rect 727 16762 1263 16774
rect 727 16710 749 16762
rect 749 16710 765 16762
rect 765 16710 817 16762
rect 817 16710 833 16762
rect 833 16710 885 16762
rect 885 16710 901 16762
rect 901 16710 953 16762
rect 953 16710 969 16762
rect 969 16710 1021 16762
rect 1021 16710 1037 16762
rect 1037 16710 1089 16762
rect 1089 16710 1105 16762
rect 1105 16710 1157 16762
rect 1157 16710 1173 16762
rect 1173 16710 1225 16762
rect 1225 16710 1241 16762
rect 1241 16710 1263 16762
rect 727 16698 1263 16710
rect 727 16687 749 16698
rect 749 16687 765 16698
rect 765 16687 817 16698
rect 817 16687 833 16698
rect 833 16687 885 16698
rect 885 16687 901 16698
rect 901 16687 953 16698
rect 953 16687 969 16698
rect 969 16687 1021 16698
rect 1021 16687 1037 16698
rect 1037 16687 1089 16698
rect 1089 16687 1105 16698
rect 1105 16687 1157 16698
rect 1157 16687 1173 16698
rect 1173 16687 1225 16698
rect 1225 16687 1241 16698
rect 1241 16687 1263 16698
rect 727 16646 749 16662
rect 749 16646 765 16662
rect 765 16646 783 16662
rect 807 16646 817 16662
rect 817 16646 833 16662
rect 833 16646 863 16662
rect 887 16646 901 16662
rect 901 16646 943 16662
rect 967 16646 969 16662
rect 969 16646 1021 16662
rect 1021 16646 1023 16662
rect 1047 16646 1089 16662
rect 1089 16646 1103 16662
rect 1127 16646 1157 16662
rect 1157 16646 1173 16662
rect 1173 16646 1183 16662
rect 1207 16646 1225 16662
rect 1225 16646 1241 16662
rect 1241 16646 1263 16662
rect 727 16634 783 16646
rect 807 16634 863 16646
rect 887 16634 943 16646
rect 967 16634 1023 16646
rect 1047 16634 1103 16646
rect 1127 16634 1183 16646
rect 1207 16634 1263 16646
rect 727 16606 749 16634
rect 749 16606 765 16634
rect 765 16606 783 16634
rect 807 16606 817 16634
rect 817 16606 833 16634
rect 833 16606 863 16634
rect 887 16606 901 16634
rect 901 16606 943 16634
rect 967 16606 969 16634
rect 969 16606 1021 16634
rect 1021 16606 1023 16634
rect 1047 16606 1089 16634
rect 1089 16606 1103 16634
rect 1127 16606 1157 16634
rect 1157 16606 1173 16634
rect 1173 16606 1183 16634
rect 1207 16606 1225 16634
rect 1225 16606 1241 16634
rect 1241 16606 1263 16634
rect 727 16570 783 16581
rect 807 16570 863 16581
rect 887 16570 943 16581
rect 967 16570 1023 16581
rect 1047 16570 1103 16581
rect 1127 16570 1183 16581
rect 1207 16570 1263 16581
rect 727 16525 749 16570
rect 749 16525 765 16570
rect 765 16525 783 16570
rect 807 16525 817 16570
rect 817 16525 833 16570
rect 833 16525 863 16570
rect 887 16525 901 16570
rect 901 16525 943 16570
rect 967 16525 969 16570
rect 969 16525 1021 16570
rect 1021 16525 1023 16570
rect 1047 16525 1089 16570
rect 1089 16525 1103 16570
rect 1127 16525 1157 16570
rect 1157 16525 1173 16570
rect 1173 16525 1183 16570
rect 1207 16525 1225 16570
rect 1225 16525 1241 16570
rect 1241 16525 1263 16570
rect 727 16454 749 16500
rect 749 16454 765 16500
rect 765 16454 783 16500
rect 807 16454 817 16500
rect 817 16454 833 16500
rect 833 16454 863 16500
rect 887 16454 901 16500
rect 901 16454 943 16500
rect 967 16454 969 16500
rect 969 16454 1021 16500
rect 1021 16454 1023 16500
rect 1047 16454 1089 16500
rect 1089 16454 1103 16500
rect 1127 16454 1157 16500
rect 1157 16454 1173 16500
rect 1173 16454 1183 16500
rect 1207 16454 1225 16500
rect 1225 16454 1241 16500
rect 1241 16454 1263 16500
rect 727 16444 783 16454
rect 807 16444 863 16454
rect 887 16444 943 16454
rect 967 16444 1023 16454
rect 1047 16444 1103 16454
rect 1127 16444 1183 16454
rect 1207 16444 1263 16454
rect 727 16390 749 16419
rect 749 16390 765 16419
rect 765 16390 783 16419
rect 807 16390 817 16419
rect 817 16390 833 16419
rect 833 16390 863 16419
rect 887 16390 901 16419
rect 901 16390 943 16419
rect 967 16390 969 16419
rect 969 16390 1021 16419
rect 1021 16390 1023 16419
rect 1047 16390 1089 16419
rect 1089 16390 1103 16419
rect 1127 16390 1157 16419
rect 1157 16390 1173 16419
rect 1173 16390 1183 16419
rect 1207 16390 1225 16419
rect 1225 16390 1241 16419
rect 1241 16390 1263 16419
rect 727 16378 783 16390
rect 807 16378 863 16390
rect 887 16378 943 16390
rect 967 16378 1023 16390
rect 1047 16378 1103 16390
rect 1127 16378 1183 16390
rect 1207 16378 1263 16390
rect 727 16363 749 16378
rect 749 16363 765 16378
rect 765 16363 783 16378
rect 807 16363 817 16378
rect 817 16363 833 16378
rect 833 16363 863 16378
rect 887 16363 901 16378
rect 901 16363 943 16378
rect 967 16363 969 16378
rect 969 16363 1021 16378
rect 1021 16363 1023 16378
rect 1047 16363 1089 16378
rect 1089 16363 1103 16378
rect 1127 16363 1157 16378
rect 1157 16363 1173 16378
rect 1173 16363 1183 16378
rect 1207 16363 1225 16378
rect 1225 16363 1241 16378
rect 1241 16363 1263 16378
rect 727 16326 749 16338
rect 749 16326 765 16338
rect 765 16326 783 16338
rect 807 16326 817 16338
rect 817 16326 833 16338
rect 833 16326 863 16338
rect 887 16326 901 16338
rect 901 16326 943 16338
rect 967 16326 969 16338
rect 969 16326 1021 16338
rect 1021 16326 1023 16338
rect 1047 16326 1089 16338
rect 1089 16326 1103 16338
rect 1127 16326 1157 16338
rect 1157 16326 1173 16338
rect 1173 16326 1183 16338
rect 1207 16326 1225 16338
rect 1225 16326 1241 16338
rect 1241 16326 1263 16338
rect 727 16314 783 16326
rect 807 16314 863 16326
rect 887 16314 943 16326
rect 967 16314 1023 16326
rect 1047 16314 1103 16326
rect 1127 16314 1183 16326
rect 1207 16314 1263 16326
rect 727 16282 749 16314
rect 749 16282 765 16314
rect 765 16282 783 16314
rect 807 16282 817 16314
rect 817 16282 833 16314
rect 833 16282 863 16314
rect 887 16282 901 16314
rect 901 16282 943 16314
rect 967 16282 969 16314
rect 969 16282 1021 16314
rect 1021 16282 1023 16314
rect 1047 16282 1089 16314
rect 1089 16282 1103 16314
rect 1127 16282 1157 16314
rect 1157 16282 1173 16314
rect 1173 16282 1183 16314
rect 1207 16282 1225 16314
rect 1225 16282 1241 16314
rect 1241 16282 1263 16314
rect 727 16250 783 16257
rect 807 16250 863 16257
rect 887 16250 943 16257
rect 967 16250 1023 16257
rect 1047 16250 1103 16257
rect 1127 16250 1183 16257
rect 1207 16250 1263 16257
rect 727 16201 749 16250
rect 749 16201 765 16250
rect 765 16201 783 16250
rect 807 16201 817 16250
rect 817 16201 833 16250
rect 833 16201 863 16250
rect 887 16201 901 16250
rect 901 16201 943 16250
rect 967 16201 969 16250
rect 969 16201 1021 16250
rect 1021 16201 1023 16250
rect 1047 16201 1089 16250
rect 1089 16201 1103 16250
rect 1127 16201 1157 16250
rect 1157 16201 1173 16250
rect 1173 16201 1183 16250
rect 1207 16201 1225 16250
rect 1225 16201 1241 16250
rect 1241 16201 1263 16250
rect 727 14957 749 15006
rect 749 14957 765 15006
rect 765 14957 817 15006
rect 817 14957 833 15006
rect 833 14957 885 15006
rect 885 14957 901 15006
rect 901 14957 953 15006
rect 953 14957 969 15006
rect 969 14957 1021 15006
rect 1021 14957 1037 15006
rect 1037 14957 1089 15006
rect 1089 14957 1105 15006
rect 1105 14957 1157 15006
rect 1157 14957 1173 15006
rect 1173 14957 1225 15006
rect 1225 14957 1241 15006
rect 1241 14957 1263 15006
rect 727 14945 1263 14957
rect 727 14893 749 14945
rect 749 14893 765 14945
rect 765 14893 817 14945
rect 817 14893 833 14945
rect 833 14893 885 14945
rect 885 14893 901 14945
rect 901 14893 953 14945
rect 953 14893 969 14945
rect 969 14893 1021 14945
rect 1021 14893 1037 14945
rect 1037 14893 1089 14945
rect 1089 14893 1105 14945
rect 1105 14893 1157 14945
rect 1157 14893 1173 14945
rect 1173 14893 1225 14945
rect 1225 14893 1241 14945
rect 1241 14893 1263 14945
rect 727 14881 1263 14893
rect 727 14829 749 14881
rect 749 14829 765 14881
rect 765 14829 817 14881
rect 817 14829 833 14881
rect 833 14829 885 14881
rect 885 14829 901 14881
rect 901 14829 953 14881
rect 953 14829 969 14881
rect 969 14829 1021 14881
rect 1021 14829 1037 14881
rect 1037 14829 1089 14881
rect 1089 14829 1105 14881
rect 1105 14829 1157 14881
rect 1157 14829 1173 14881
rect 1173 14829 1225 14881
rect 1225 14829 1241 14881
rect 1241 14829 1263 14881
rect 727 14817 1263 14829
rect 727 14765 749 14817
rect 749 14765 765 14817
rect 765 14765 817 14817
rect 817 14765 833 14817
rect 833 14765 885 14817
rect 885 14765 901 14817
rect 901 14765 953 14817
rect 953 14765 969 14817
rect 969 14765 1021 14817
rect 1021 14765 1037 14817
rect 1037 14765 1089 14817
rect 1089 14765 1105 14817
rect 1105 14765 1157 14817
rect 1157 14765 1173 14817
rect 1173 14765 1225 14817
rect 1225 14765 1241 14817
rect 1241 14765 1263 14817
rect 727 14753 1263 14765
rect 727 14701 749 14753
rect 749 14701 765 14753
rect 765 14701 817 14753
rect 817 14701 833 14753
rect 833 14701 885 14753
rect 885 14701 901 14753
rect 901 14701 953 14753
rect 953 14701 969 14753
rect 969 14701 1021 14753
rect 1021 14701 1037 14753
rect 1037 14701 1089 14753
rect 1089 14701 1105 14753
rect 1105 14701 1157 14753
rect 1157 14701 1173 14753
rect 1173 14701 1225 14753
rect 1225 14701 1241 14753
rect 1241 14701 1263 14753
rect 727 14689 1263 14701
rect 727 14637 749 14689
rect 749 14637 765 14689
rect 765 14637 817 14689
rect 817 14637 833 14689
rect 833 14637 885 14689
rect 885 14637 901 14689
rect 901 14637 953 14689
rect 953 14637 969 14689
rect 969 14637 1021 14689
rect 1021 14637 1037 14689
rect 1037 14637 1089 14689
rect 1089 14637 1105 14689
rect 1105 14637 1157 14689
rect 1157 14637 1173 14689
rect 1173 14637 1225 14689
rect 1225 14637 1241 14689
rect 1241 14637 1263 14689
rect 727 14625 1263 14637
rect 727 14573 749 14625
rect 749 14573 765 14625
rect 765 14573 817 14625
rect 817 14573 833 14625
rect 833 14573 885 14625
rect 885 14573 901 14625
rect 901 14573 953 14625
rect 953 14573 969 14625
rect 969 14573 1021 14625
rect 1021 14573 1037 14625
rect 1037 14573 1089 14625
rect 1089 14573 1105 14625
rect 1105 14573 1157 14625
rect 1157 14573 1173 14625
rect 1173 14573 1225 14625
rect 1225 14573 1241 14625
rect 1241 14573 1263 14625
rect 727 14561 1263 14573
rect 727 14550 749 14561
rect 749 14550 765 14561
rect 765 14550 817 14561
rect 817 14550 833 14561
rect 833 14550 885 14561
rect 885 14550 901 14561
rect 901 14550 953 14561
rect 953 14550 969 14561
rect 969 14550 1021 14561
rect 1021 14550 1037 14561
rect 1037 14550 1089 14561
rect 1089 14550 1105 14561
rect 1105 14550 1157 14561
rect 1157 14550 1173 14561
rect 1173 14550 1225 14561
rect 1225 14550 1241 14561
rect 1241 14550 1263 14561
rect 727 14509 749 14525
rect 749 14509 765 14525
rect 765 14509 783 14525
rect 807 14509 817 14525
rect 817 14509 833 14525
rect 833 14509 863 14525
rect 887 14509 901 14525
rect 901 14509 943 14525
rect 967 14509 969 14525
rect 969 14509 1021 14525
rect 1021 14509 1023 14525
rect 1047 14509 1089 14525
rect 1089 14509 1103 14525
rect 1127 14509 1157 14525
rect 1157 14509 1173 14525
rect 1173 14509 1183 14525
rect 1207 14509 1225 14525
rect 1225 14509 1241 14525
rect 1241 14509 1263 14525
rect 727 14497 783 14509
rect 807 14497 863 14509
rect 887 14497 943 14509
rect 967 14497 1023 14509
rect 1047 14497 1103 14509
rect 1127 14497 1183 14509
rect 1207 14497 1263 14509
rect 727 14469 749 14497
rect 749 14469 765 14497
rect 765 14469 783 14497
rect 807 14469 817 14497
rect 817 14469 833 14497
rect 833 14469 863 14497
rect 887 14469 901 14497
rect 901 14469 943 14497
rect 967 14469 969 14497
rect 969 14469 1021 14497
rect 1021 14469 1023 14497
rect 1047 14469 1089 14497
rect 1089 14469 1103 14497
rect 1127 14469 1157 14497
rect 1157 14469 1173 14497
rect 1173 14469 1183 14497
rect 1207 14469 1225 14497
rect 1225 14469 1241 14497
rect 1241 14469 1263 14497
rect 727 14433 783 14444
rect 807 14433 863 14444
rect 887 14433 943 14444
rect 967 14433 1023 14444
rect 1047 14433 1103 14444
rect 1127 14433 1183 14444
rect 1207 14433 1263 14444
rect 727 14388 749 14433
rect 749 14388 765 14433
rect 765 14388 783 14433
rect 807 14388 817 14433
rect 817 14388 833 14433
rect 833 14388 863 14433
rect 887 14388 901 14433
rect 901 14388 943 14433
rect 967 14388 969 14433
rect 969 14388 1021 14433
rect 1021 14388 1023 14433
rect 1047 14388 1089 14433
rect 1089 14388 1103 14433
rect 1127 14388 1157 14433
rect 1157 14388 1173 14433
rect 1173 14388 1183 14433
rect 1207 14388 1225 14433
rect 1225 14388 1241 14433
rect 1241 14388 1263 14433
rect 727 14317 749 14363
rect 749 14317 765 14363
rect 765 14317 783 14363
rect 807 14317 817 14363
rect 817 14317 833 14363
rect 833 14317 863 14363
rect 887 14317 901 14363
rect 901 14317 943 14363
rect 967 14317 969 14363
rect 969 14317 1021 14363
rect 1021 14317 1023 14363
rect 1047 14317 1089 14363
rect 1089 14317 1103 14363
rect 1127 14317 1157 14363
rect 1157 14317 1173 14363
rect 1173 14317 1183 14363
rect 1207 14317 1225 14363
rect 1225 14317 1241 14363
rect 1241 14317 1263 14363
rect 727 14307 783 14317
rect 807 14307 863 14317
rect 887 14307 943 14317
rect 967 14307 1023 14317
rect 1047 14307 1103 14317
rect 1127 14307 1183 14317
rect 1207 14307 1263 14317
rect 727 14253 749 14282
rect 749 14253 765 14282
rect 765 14253 783 14282
rect 807 14253 817 14282
rect 817 14253 833 14282
rect 833 14253 863 14282
rect 887 14253 901 14282
rect 901 14253 943 14282
rect 967 14253 969 14282
rect 969 14253 1021 14282
rect 1021 14253 1023 14282
rect 1047 14253 1089 14282
rect 1089 14253 1103 14282
rect 1127 14253 1157 14282
rect 1157 14253 1173 14282
rect 1173 14253 1183 14282
rect 1207 14253 1225 14282
rect 1225 14253 1241 14282
rect 1241 14253 1263 14282
rect 727 14241 783 14253
rect 807 14241 863 14253
rect 887 14241 943 14253
rect 967 14241 1023 14253
rect 1047 14241 1103 14253
rect 1127 14241 1183 14253
rect 1207 14241 1263 14253
rect 727 14226 749 14241
rect 749 14226 765 14241
rect 765 14226 783 14241
rect 807 14226 817 14241
rect 817 14226 833 14241
rect 833 14226 863 14241
rect 887 14226 901 14241
rect 901 14226 943 14241
rect 967 14226 969 14241
rect 969 14226 1021 14241
rect 1021 14226 1023 14241
rect 1047 14226 1089 14241
rect 1089 14226 1103 14241
rect 1127 14226 1157 14241
rect 1157 14226 1173 14241
rect 1173 14226 1183 14241
rect 1207 14226 1225 14241
rect 1225 14226 1241 14241
rect 1241 14226 1263 14241
rect 727 14189 749 14201
rect 749 14189 765 14201
rect 765 14189 783 14201
rect 807 14189 817 14201
rect 817 14189 833 14201
rect 833 14189 863 14201
rect 887 14189 901 14201
rect 901 14189 943 14201
rect 967 14189 969 14201
rect 969 14189 1021 14201
rect 1021 14189 1023 14201
rect 1047 14189 1089 14201
rect 1089 14189 1103 14201
rect 1127 14189 1157 14201
rect 1157 14189 1173 14201
rect 1173 14189 1183 14201
rect 1207 14189 1225 14201
rect 1225 14189 1241 14201
rect 1241 14189 1263 14201
rect 727 14177 783 14189
rect 807 14177 863 14189
rect 887 14177 943 14189
rect 967 14177 1023 14189
rect 1047 14177 1103 14189
rect 1127 14177 1183 14189
rect 1207 14177 1263 14189
rect 727 14145 749 14177
rect 749 14145 765 14177
rect 765 14145 783 14177
rect 807 14145 817 14177
rect 817 14145 833 14177
rect 833 14145 863 14177
rect 887 14145 901 14177
rect 901 14145 943 14177
rect 967 14145 969 14177
rect 969 14145 1021 14177
rect 1021 14145 1023 14177
rect 1047 14145 1089 14177
rect 1089 14145 1103 14177
rect 1127 14145 1157 14177
rect 1157 14145 1173 14177
rect 1173 14145 1183 14177
rect 1207 14145 1225 14177
rect 1225 14145 1241 14177
rect 1241 14145 1263 14177
rect 727 14113 783 14120
rect 807 14113 863 14120
rect 887 14113 943 14120
rect 967 14113 1023 14120
rect 1047 14113 1103 14120
rect 1127 14113 1183 14120
rect 1207 14113 1263 14120
rect 727 14064 749 14113
rect 749 14064 765 14113
rect 765 14064 783 14113
rect 807 14064 817 14113
rect 817 14064 833 14113
rect 833 14064 863 14113
rect 887 14064 901 14113
rect 901 14064 943 14113
rect 967 14064 969 14113
rect 969 14064 1021 14113
rect 1021 14064 1023 14113
rect 1047 14064 1089 14113
rect 1089 14064 1103 14113
rect 1127 14064 1157 14113
rect 1157 14064 1173 14113
rect 1173 14064 1183 14113
rect 1207 14064 1225 14113
rect 1225 14064 1241 14113
rect 1241 14064 1263 14113
rect 115 13649 117 13698
rect 117 13649 169 13698
rect 169 13649 171 13698
rect 115 13642 171 13649
rect 115 13581 117 13617
rect 117 13581 169 13617
rect 169 13581 171 13617
rect 115 13565 171 13581
rect 115 13561 117 13565
rect 117 13561 169 13565
rect 169 13561 171 13565
rect 115 13513 117 13536
rect 117 13513 169 13536
rect 169 13513 171 13536
rect 115 13496 171 13513
rect 115 13480 117 13496
rect 117 13480 169 13496
rect 169 13480 171 13496
rect 115 13444 117 13455
rect 117 13444 169 13455
rect 169 13444 171 13455
rect 115 13427 171 13444
rect 115 13399 117 13427
rect 117 13399 169 13427
rect 169 13399 171 13427
rect 115 13358 171 13374
rect 115 13318 117 13358
rect 117 13318 169 13358
rect 169 13318 171 13358
rect 115 13289 171 13292
rect 115 13237 117 13289
rect 117 13237 169 13289
rect 169 13237 171 13289
rect 115 13236 171 13237
rect 115 13168 117 13210
rect 117 13168 169 13210
rect 169 13168 171 13210
rect 115 13154 171 13168
rect 115 13099 117 13128
rect 117 13099 169 13128
rect 169 13099 171 13128
rect 115 13082 171 13099
rect 115 13072 117 13082
rect 117 13072 169 13082
rect 169 13072 171 13082
rect 115 13030 117 13046
rect 117 13030 169 13046
rect 169 13030 171 13046
rect 115 13013 171 13030
rect 115 12990 117 13013
rect 117 12990 169 13013
rect 169 12990 171 13013
rect 115 12961 117 12964
rect 117 12961 169 12964
rect 169 12961 171 12964
rect 115 12944 171 12961
rect 115 12908 117 12944
rect 117 12908 169 12944
rect 169 12908 171 12944
rect 115 12875 171 12882
rect 115 12826 117 12875
rect 117 12826 169 12875
rect 169 12826 171 12875
rect 727 12855 749 12904
rect 749 12855 765 12904
rect 765 12855 817 12904
rect 817 12855 833 12904
rect 833 12855 885 12904
rect 885 12855 901 12904
rect 901 12855 953 12904
rect 953 12855 969 12904
rect 969 12855 1021 12904
rect 1021 12855 1037 12904
rect 1037 12855 1089 12904
rect 1089 12855 1105 12904
rect 1105 12855 1157 12904
rect 1157 12855 1173 12904
rect 1173 12855 1225 12904
rect 1225 12855 1241 12904
rect 1241 12855 1263 12904
rect 727 12843 1263 12855
rect 727 12791 749 12843
rect 749 12791 765 12843
rect 765 12791 817 12843
rect 817 12791 833 12843
rect 833 12791 885 12843
rect 885 12791 901 12843
rect 901 12791 953 12843
rect 953 12791 969 12843
rect 969 12791 1021 12843
rect 1021 12791 1037 12843
rect 1037 12791 1089 12843
rect 1089 12791 1105 12843
rect 1105 12791 1157 12843
rect 1157 12791 1173 12843
rect 1173 12791 1225 12843
rect 1225 12791 1241 12843
rect 1241 12791 1263 12843
rect 727 12779 1263 12791
rect 727 12727 749 12779
rect 749 12727 765 12779
rect 765 12727 817 12779
rect 817 12727 833 12779
rect 833 12727 885 12779
rect 885 12727 901 12779
rect 901 12727 953 12779
rect 953 12727 969 12779
rect 969 12727 1021 12779
rect 1021 12727 1037 12779
rect 1037 12727 1089 12779
rect 1089 12727 1105 12779
rect 1105 12727 1157 12779
rect 1157 12727 1173 12779
rect 1173 12727 1225 12779
rect 1225 12727 1241 12779
rect 1241 12727 1263 12779
rect 727 12715 1263 12727
rect 727 12663 749 12715
rect 749 12663 765 12715
rect 765 12663 817 12715
rect 817 12663 833 12715
rect 833 12663 885 12715
rect 885 12663 901 12715
rect 901 12663 953 12715
rect 953 12663 969 12715
rect 969 12663 1021 12715
rect 1021 12663 1037 12715
rect 1037 12663 1089 12715
rect 1089 12663 1105 12715
rect 1105 12663 1157 12715
rect 1157 12663 1173 12715
rect 1173 12663 1225 12715
rect 1225 12663 1241 12715
rect 1241 12663 1263 12715
rect 727 12651 1263 12663
rect 727 12599 749 12651
rect 749 12599 765 12651
rect 765 12599 817 12651
rect 817 12599 833 12651
rect 833 12599 885 12651
rect 885 12599 901 12651
rect 901 12599 953 12651
rect 953 12599 969 12651
rect 969 12599 1021 12651
rect 1021 12599 1037 12651
rect 1037 12599 1089 12651
rect 1089 12599 1105 12651
rect 1105 12599 1157 12651
rect 1157 12599 1173 12651
rect 1173 12599 1225 12651
rect 1225 12599 1241 12651
rect 1241 12599 1263 12651
rect 727 12587 1263 12599
rect 727 12535 749 12587
rect 749 12535 765 12587
rect 765 12535 817 12587
rect 817 12535 833 12587
rect 833 12535 885 12587
rect 885 12535 901 12587
rect 901 12535 953 12587
rect 953 12535 969 12587
rect 969 12535 1021 12587
rect 1021 12535 1037 12587
rect 1037 12535 1089 12587
rect 1089 12535 1105 12587
rect 1105 12535 1157 12587
rect 1157 12535 1173 12587
rect 1173 12535 1225 12587
rect 1225 12535 1241 12587
rect 1241 12535 1263 12587
rect 727 12523 1263 12535
rect 727 12471 749 12523
rect 749 12471 765 12523
rect 765 12471 817 12523
rect 817 12471 833 12523
rect 833 12471 885 12523
rect 885 12471 901 12523
rect 901 12471 953 12523
rect 953 12471 969 12523
rect 969 12471 1021 12523
rect 1021 12471 1037 12523
rect 1037 12471 1089 12523
rect 1089 12471 1105 12523
rect 1105 12471 1157 12523
rect 1157 12471 1173 12523
rect 1173 12471 1225 12523
rect 1225 12471 1241 12523
rect 1241 12471 1263 12523
rect 727 12459 1263 12471
rect 727 12448 749 12459
rect 749 12448 765 12459
rect 765 12448 817 12459
rect 817 12448 833 12459
rect 833 12448 885 12459
rect 885 12448 901 12459
rect 901 12448 953 12459
rect 953 12448 969 12459
rect 969 12448 1021 12459
rect 1021 12448 1037 12459
rect 1037 12448 1089 12459
rect 1089 12448 1105 12459
rect 1105 12448 1157 12459
rect 1157 12448 1173 12459
rect 1173 12448 1225 12459
rect 1225 12448 1241 12459
rect 1241 12448 1263 12459
rect 727 12407 749 12423
rect 749 12407 765 12423
rect 765 12407 783 12423
rect 807 12407 817 12423
rect 817 12407 833 12423
rect 833 12407 863 12423
rect 887 12407 901 12423
rect 901 12407 943 12423
rect 967 12407 969 12423
rect 969 12407 1021 12423
rect 1021 12407 1023 12423
rect 1047 12407 1089 12423
rect 1089 12407 1103 12423
rect 1127 12407 1157 12423
rect 1157 12407 1173 12423
rect 1173 12407 1183 12423
rect 1207 12407 1225 12423
rect 1225 12407 1241 12423
rect 1241 12407 1263 12423
rect 727 12395 783 12407
rect 807 12395 863 12407
rect 887 12395 943 12407
rect 967 12395 1023 12407
rect 1047 12395 1103 12407
rect 1127 12395 1183 12407
rect 1207 12395 1263 12407
rect 727 12367 749 12395
rect 749 12367 765 12395
rect 765 12367 783 12395
rect 807 12367 817 12395
rect 817 12367 833 12395
rect 833 12367 863 12395
rect 887 12367 901 12395
rect 901 12367 943 12395
rect 967 12367 969 12395
rect 969 12367 1021 12395
rect 1021 12367 1023 12395
rect 1047 12367 1089 12395
rect 1089 12367 1103 12395
rect 1127 12367 1157 12395
rect 1157 12367 1173 12395
rect 1173 12367 1183 12395
rect 1207 12367 1225 12395
rect 1225 12367 1241 12395
rect 1241 12367 1263 12395
rect 727 12331 783 12342
rect 807 12331 863 12342
rect 887 12331 943 12342
rect 967 12331 1023 12342
rect 1047 12331 1103 12342
rect 1127 12331 1183 12342
rect 1207 12331 1263 12342
rect 727 12286 749 12331
rect 749 12286 765 12331
rect 765 12286 783 12331
rect 807 12286 817 12331
rect 817 12286 833 12331
rect 833 12286 863 12331
rect 887 12286 901 12331
rect 901 12286 943 12331
rect 967 12286 969 12331
rect 969 12286 1021 12331
rect 1021 12286 1023 12331
rect 1047 12286 1089 12331
rect 1089 12286 1103 12331
rect 1127 12286 1157 12331
rect 1157 12286 1173 12331
rect 1173 12286 1183 12331
rect 1207 12286 1225 12331
rect 1225 12286 1241 12331
rect 1241 12286 1263 12331
rect 727 12215 749 12261
rect 749 12215 765 12261
rect 765 12215 783 12261
rect 807 12215 817 12261
rect 817 12215 833 12261
rect 833 12215 863 12261
rect 887 12215 901 12261
rect 901 12215 943 12261
rect 967 12215 969 12261
rect 969 12215 1021 12261
rect 1021 12215 1023 12261
rect 1047 12215 1089 12261
rect 1089 12215 1103 12261
rect 1127 12215 1157 12261
rect 1157 12215 1173 12261
rect 1173 12215 1183 12261
rect 1207 12215 1225 12261
rect 1225 12215 1241 12261
rect 1241 12215 1263 12261
rect 727 12205 783 12215
rect 807 12205 863 12215
rect 887 12205 943 12215
rect 967 12205 1023 12215
rect 1047 12205 1103 12215
rect 1127 12205 1183 12215
rect 1207 12205 1263 12215
rect 727 12151 749 12180
rect 749 12151 765 12180
rect 765 12151 783 12180
rect 807 12151 817 12180
rect 817 12151 833 12180
rect 833 12151 863 12180
rect 887 12151 901 12180
rect 901 12151 943 12180
rect 967 12151 969 12180
rect 969 12151 1021 12180
rect 1021 12151 1023 12180
rect 1047 12151 1089 12180
rect 1089 12151 1103 12180
rect 1127 12151 1157 12180
rect 1157 12151 1173 12180
rect 1173 12151 1183 12180
rect 1207 12151 1225 12180
rect 1225 12151 1241 12180
rect 1241 12151 1263 12180
rect 727 12139 783 12151
rect 807 12139 863 12151
rect 887 12139 943 12151
rect 967 12139 1023 12151
rect 1047 12139 1103 12151
rect 1127 12139 1183 12151
rect 1207 12139 1263 12151
rect 727 12124 749 12139
rect 749 12124 765 12139
rect 765 12124 783 12139
rect 807 12124 817 12139
rect 817 12124 833 12139
rect 833 12124 863 12139
rect 887 12124 901 12139
rect 901 12124 943 12139
rect 967 12124 969 12139
rect 969 12124 1021 12139
rect 1021 12124 1023 12139
rect 1047 12124 1089 12139
rect 1089 12124 1103 12139
rect 1127 12124 1157 12139
rect 1157 12124 1173 12139
rect 1173 12124 1183 12139
rect 1207 12124 1225 12139
rect 1225 12124 1241 12139
rect 1241 12124 1263 12139
rect 727 12087 749 12099
rect 749 12087 765 12099
rect 765 12087 783 12099
rect 807 12087 817 12099
rect 817 12087 833 12099
rect 833 12087 863 12099
rect 887 12087 901 12099
rect 901 12087 943 12099
rect 967 12087 969 12099
rect 969 12087 1021 12099
rect 1021 12087 1023 12099
rect 1047 12087 1089 12099
rect 1089 12087 1103 12099
rect 1127 12087 1157 12099
rect 1157 12087 1173 12099
rect 1173 12087 1183 12099
rect 1207 12087 1225 12099
rect 1225 12087 1241 12099
rect 1241 12087 1263 12099
rect 727 12075 783 12087
rect 807 12075 863 12087
rect 887 12075 943 12087
rect 967 12075 1023 12087
rect 1047 12075 1103 12087
rect 1127 12075 1183 12087
rect 1207 12075 1263 12087
rect 727 12043 749 12075
rect 749 12043 765 12075
rect 765 12043 783 12075
rect 807 12043 817 12075
rect 817 12043 833 12075
rect 833 12043 863 12075
rect 887 12043 901 12075
rect 901 12043 943 12075
rect 967 12043 969 12075
rect 969 12043 1021 12075
rect 1021 12043 1023 12075
rect 1047 12043 1089 12075
rect 1089 12043 1103 12075
rect 1127 12043 1157 12075
rect 1157 12043 1173 12075
rect 1173 12043 1183 12075
rect 1207 12043 1225 12075
rect 1225 12043 1241 12075
rect 1241 12043 1263 12075
rect 727 12011 783 12018
rect 807 12011 863 12018
rect 887 12011 943 12018
rect 967 12011 1023 12018
rect 1047 12011 1103 12018
rect 1127 12011 1183 12018
rect 1207 12011 1263 12018
rect 727 11962 749 12011
rect 749 11962 765 12011
rect 765 11962 783 12011
rect 807 11962 817 12011
rect 817 11962 833 12011
rect 833 11962 863 12011
rect 887 11962 901 12011
rect 901 11962 943 12011
rect 967 11962 969 12011
rect 969 11962 1021 12011
rect 1021 11962 1023 12011
rect 1047 11962 1089 12011
rect 1089 11962 1103 12011
rect 1127 11962 1157 12011
rect 1157 11962 1173 12011
rect 1173 11962 1183 12011
rect 1207 11962 1225 12011
rect 1225 11962 1241 12011
rect 1241 11962 1263 12011
rect 727 10761 749 10810
rect 749 10761 765 10810
rect 765 10761 817 10810
rect 817 10761 833 10810
rect 833 10761 885 10810
rect 885 10761 901 10810
rect 901 10761 953 10810
rect 953 10761 969 10810
rect 969 10761 1021 10810
rect 1021 10761 1037 10810
rect 1037 10761 1089 10810
rect 1089 10761 1105 10810
rect 1105 10761 1157 10810
rect 1157 10761 1173 10810
rect 1173 10761 1225 10810
rect 1225 10761 1241 10810
rect 1241 10761 1263 10810
rect 727 10749 1263 10761
rect 727 10697 749 10749
rect 749 10697 765 10749
rect 765 10697 817 10749
rect 817 10697 833 10749
rect 833 10697 885 10749
rect 885 10697 901 10749
rect 901 10697 953 10749
rect 953 10697 969 10749
rect 969 10697 1021 10749
rect 1021 10697 1037 10749
rect 1037 10697 1089 10749
rect 1089 10697 1105 10749
rect 1105 10697 1157 10749
rect 1157 10697 1173 10749
rect 1173 10697 1225 10749
rect 1225 10697 1241 10749
rect 1241 10697 1263 10749
rect 727 10685 1263 10697
rect 727 10633 749 10685
rect 749 10633 765 10685
rect 765 10633 817 10685
rect 817 10633 833 10685
rect 833 10633 885 10685
rect 885 10633 901 10685
rect 901 10633 953 10685
rect 953 10633 969 10685
rect 969 10633 1021 10685
rect 1021 10633 1037 10685
rect 1037 10633 1089 10685
rect 1089 10633 1105 10685
rect 1105 10633 1157 10685
rect 1157 10633 1173 10685
rect 1173 10633 1225 10685
rect 1225 10633 1241 10685
rect 1241 10633 1263 10685
rect 727 10621 1263 10633
rect 727 10569 749 10621
rect 749 10569 765 10621
rect 765 10569 817 10621
rect 817 10569 833 10621
rect 833 10569 885 10621
rect 885 10569 901 10621
rect 901 10569 953 10621
rect 953 10569 969 10621
rect 969 10569 1021 10621
rect 1021 10569 1037 10621
rect 1037 10569 1089 10621
rect 1089 10569 1105 10621
rect 1105 10569 1157 10621
rect 1157 10569 1173 10621
rect 1173 10569 1225 10621
rect 1225 10569 1241 10621
rect 1241 10569 1263 10621
rect 727 10557 1263 10569
rect 727 10505 749 10557
rect 749 10505 765 10557
rect 765 10505 817 10557
rect 817 10505 833 10557
rect 833 10505 885 10557
rect 885 10505 901 10557
rect 901 10505 953 10557
rect 953 10505 969 10557
rect 969 10505 1021 10557
rect 1021 10505 1037 10557
rect 1037 10505 1089 10557
rect 1089 10505 1105 10557
rect 1105 10505 1157 10557
rect 1157 10505 1173 10557
rect 1173 10505 1225 10557
rect 1225 10505 1241 10557
rect 1241 10505 1263 10557
rect 727 10493 1263 10505
rect 727 10441 749 10493
rect 749 10441 765 10493
rect 765 10441 817 10493
rect 817 10441 833 10493
rect 833 10441 885 10493
rect 885 10441 901 10493
rect 901 10441 953 10493
rect 953 10441 969 10493
rect 969 10441 1021 10493
rect 1021 10441 1037 10493
rect 1037 10441 1089 10493
rect 1089 10441 1105 10493
rect 1105 10441 1157 10493
rect 1157 10441 1173 10493
rect 1173 10441 1225 10493
rect 1225 10441 1241 10493
rect 1241 10441 1263 10493
rect 727 10429 1263 10441
rect 727 10377 749 10429
rect 749 10377 765 10429
rect 765 10377 817 10429
rect 817 10377 833 10429
rect 833 10377 885 10429
rect 885 10377 901 10429
rect 901 10377 953 10429
rect 953 10377 969 10429
rect 969 10377 1021 10429
rect 1021 10377 1037 10429
rect 1037 10377 1089 10429
rect 1089 10377 1105 10429
rect 1105 10377 1157 10429
rect 1157 10377 1173 10429
rect 1173 10377 1225 10429
rect 1225 10377 1241 10429
rect 1241 10377 1263 10429
rect 727 10365 1263 10377
rect 727 10354 749 10365
rect 749 10354 765 10365
rect 765 10354 817 10365
rect 817 10354 833 10365
rect 833 10354 885 10365
rect 885 10354 901 10365
rect 901 10354 953 10365
rect 953 10354 969 10365
rect 969 10354 1021 10365
rect 1021 10354 1037 10365
rect 1037 10354 1089 10365
rect 1089 10354 1105 10365
rect 1105 10354 1157 10365
rect 1157 10354 1173 10365
rect 1173 10354 1225 10365
rect 1225 10354 1241 10365
rect 1241 10354 1263 10365
rect 727 10313 749 10329
rect 749 10313 765 10329
rect 765 10313 783 10329
rect 807 10313 817 10329
rect 817 10313 833 10329
rect 833 10313 863 10329
rect 887 10313 901 10329
rect 901 10313 943 10329
rect 967 10313 969 10329
rect 969 10313 1021 10329
rect 1021 10313 1023 10329
rect 1047 10313 1089 10329
rect 1089 10313 1103 10329
rect 1127 10313 1157 10329
rect 1157 10313 1173 10329
rect 1173 10313 1183 10329
rect 1207 10313 1225 10329
rect 1225 10313 1241 10329
rect 1241 10313 1263 10329
rect 727 10301 783 10313
rect 807 10301 863 10313
rect 887 10301 943 10313
rect 967 10301 1023 10313
rect 1047 10301 1103 10313
rect 1127 10301 1183 10313
rect 1207 10301 1263 10313
rect 727 10273 749 10301
rect 749 10273 765 10301
rect 765 10273 783 10301
rect 807 10273 817 10301
rect 817 10273 833 10301
rect 833 10273 863 10301
rect 887 10273 901 10301
rect 901 10273 943 10301
rect 967 10273 969 10301
rect 969 10273 1021 10301
rect 1021 10273 1023 10301
rect 1047 10273 1089 10301
rect 1089 10273 1103 10301
rect 1127 10273 1157 10301
rect 1157 10273 1173 10301
rect 1173 10273 1183 10301
rect 1207 10273 1225 10301
rect 1225 10273 1241 10301
rect 1241 10273 1263 10301
rect 727 10237 783 10248
rect 807 10237 863 10248
rect 887 10237 943 10248
rect 967 10237 1023 10248
rect 1047 10237 1103 10248
rect 1127 10237 1183 10248
rect 1207 10237 1263 10248
rect 727 10192 749 10237
rect 749 10192 765 10237
rect 765 10192 783 10237
rect 807 10192 817 10237
rect 817 10192 833 10237
rect 833 10192 863 10237
rect 887 10192 901 10237
rect 901 10192 943 10237
rect 967 10192 969 10237
rect 969 10192 1021 10237
rect 1021 10192 1023 10237
rect 1047 10192 1089 10237
rect 1089 10192 1103 10237
rect 1127 10192 1157 10237
rect 1157 10192 1173 10237
rect 1173 10192 1183 10237
rect 1207 10192 1225 10237
rect 1225 10192 1241 10237
rect 1241 10192 1263 10237
rect 727 10121 749 10167
rect 749 10121 765 10167
rect 765 10121 783 10167
rect 807 10121 817 10167
rect 817 10121 833 10167
rect 833 10121 863 10167
rect 887 10121 901 10167
rect 901 10121 943 10167
rect 967 10121 969 10167
rect 969 10121 1021 10167
rect 1021 10121 1023 10167
rect 1047 10121 1089 10167
rect 1089 10121 1103 10167
rect 1127 10121 1157 10167
rect 1157 10121 1173 10167
rect 1173 10121 1183 10167
rect 1207 10121 1225 10167
rect 1225 10121 1241 10167
rect 1241 10121 1263 10167
rect 727 10111 783 10121
rect 807 10111 863 10121
rect 887 10111 943 10121
rect 967 10111 1023 10121
rect 1047 10111 1103 10121
rect 1127 10111 1183 10121
rect 1207 10111 1263 10121
rect 727 10057 749 10086
rect 749 10057 765 10086
rect 765 10057 783 10086
rect 807 10057 817 10086
rect 817 10057 833 10086
rect 833 10057 863 10086
rect 887 10057 901 10086
rect 901 10057 943 10086
rect 967 10057 969 10086
rect 969 10057 1021 10086
rect 1021 10057 1023 10086
rect 1047 10057 1089 10086
rect 1089 10057 1103 10086
rect 1127 10057 1157 10086
rect 1157 10057 1173 10086
rect 1173 10057 1183 10086
rect 1207 10057 1225 10086
rect 1225 10057 1241 10086
rect 1241 10057 1263 10086
rect 727 10045 783 10057
rect 807 10045 863 10057
rect 887 10045 943 10057
rect 967 10045 1023 10057
rect 1047 10045 1103 10057
rect 1127 10045 1183 10057
rect 1207 10045 1263 10057
rect 727 10030 749 10045
rect 749 10030 765 10045
rect 765 10030 783 10045
rect 807 10030 817 10045
rect 817 10030 833 10045
rect 833 10030 863 10045
rect 887 10030 901 10045
rect 901 10030 943 10045
rect 967 10030 969 10045
rect 969 10030 1021 10045
rect 1021 10030 1023 10045
rect 1047 10030 1089 10045
rect 1089 10030 1103 10045
rect 1127 10030 1157 10045
rect 1157 10030 1173 10045
rect 1173 10030 1183 10045
rect 1207 10030 1225 10045
rect 1225 10030 1241 10045
rect 1241 10030 1263 10045
rect 727 9993 749 10005
rect 749 9993 765 10005
rect 765 9993 783 10005
rect 807 9993 817 10005
rect 817 9993 833 10005
rect 833 9993 863 10005
rect 887 9993 901 10005
rect 901 9993 943 10005
rect 967 9993 969 10005
rect 969 9993 1021 10005
rect 1021 9993 1023 10005
rect 1047 9993 1089 10005
rect 1089 9993 1103 10005
rect 1127 9993 1157 10005
rect 1157 9993 1173 10005
rect 1173 9993 1183 10005
rect 1207 9993 1225 10005
rect 1225 9993 1241 10005
rect 1241 9993 1263 10005
rect 727 9981 783 9993
rect 807 9981 863 9993
rect 887 9981 943 9993
rect 967 9981 1023 9993
rect 1047 9981 1103 9993
rect 1127 9981 1183 9993
rect 1207 9981 1263 9993
rect 727 9949 749 9981
rect 749 9949 765 9981
rect 765 9949 783 9981
rect 807 9949 817 9981
rect 817 9949 833 9981
rect 833 9949 863 9981
rect 887 9949 901 9981
rect 901 9949 943 9981
rect 967 9949 969 9981
rect 969 9949 1021 9981
rect 1021 9949 1023 9981
rect 1047 9949 1089 9981
rect 1089 9949 1103 9981
rect 1127 9949 1157 9981
rect 1157 9949 1173 9981
rect 1173 9949 1183 9981
rect 1207 9949 1225 9981
rect 1225 9949 1241 9981
rect 1241 9949 1263 9981
rect 727 9917 783 9924
rect 807 9917 863 9924
rect 887 9917 943 9924
rect 967 9917 1023 9924
rect 1047 9917 1103 9924
rect 1127 9917 1183 9924
rect 1207 9917 1263 9924
rect 727 9868 749 9917
rect 749 9868 765 9917
rect 765 9868 783 9917
rect 807 9868 817 9917
rect 817 9868 833 9917
rect 833 9868 863 9917
rect 887 9868 901 9917
rect 901 9868 943 9917
rect 967 9868 969 9917
rect 969 9868 1021 9917
rect 1021 9868 1023 9917
rect 1047 9868 1089 9917
rect 1089 9868 1103 9917
rect 1127 9868 1157 9917
rect 1157 9868 1173 9917
rect 1173 9868 1183 9917
rect 1207 9868 1225 9917
rect 1225 9868 1241 9917
rect 1241 9868 1263 9917
rect 727 8559 749 8608
rect 749 8559 765 8608
rect 765 8559 817 8608
rect 817 8559 833 8608
rect 833 8559 885 8608
rect 885 8559 901 8608
rect 901 8559 953 8608
rect 953 8559 969 8608
rect 969 8559 1021 8608
rect 1021 8559 1037 8608
rect 1037 8559 1089 8608
rect 1089 8559 1105 8608
rect 1105 8559 1157 8608
rect 1157 8559 1173 8608
rect 1173 8559 1225 8608
rect 1225 8559 1241 8608
rect 1241 8559 1263 8608
rect 727 8547 1263 8559
rect 727 8495 749 8547
rect 749 8495 765 8547
rect 765 8495 817 8547
rect 817 8495 833 8547
rect 833 8495 885 8547
rect 885 8495 901 8547
rect 901 8495 953 8547
rect 953 8495 969 8547
rect 969 8495 1021 8547
rect 1021 8495 1037 8547
rect 1037 8495 1089 8547
rect 1089 8495 1105 8547
rect 1105 8495 1157 8547
rect 1157 8495 1173 8547
rect 1173 8495 1225 8547
rect 1225 8495 1241 8547
rect 1241 8495 1263 8547
rect 727 8483 1263 8495
rect 727 8431 749 8483
rect 749 8431 765 8483
rect 765 8431 817 8483
rect 817 8431 833 8483
rect 833 8431 885 8483
rect 885 8431 901 8483
rect 901 8431 953 8483
rect 953 8431 969 8483
rect 969 8431 1021 8483
rect 1021 8431 1037 8483
rect 1037 8431 1089 8483
rect 1089 8431 1105 8483
rect 1105 8431 1157 8483
rect 1157 8431 1173 8483
rect 1173 8431 1225 8483
rect 1225 8431 1241 8483
rect 1241 8431 1263 8483
rect 727 8419 1263 8431
rect 727 8367 749 8419
rect 749 8367 765 8419
rect 765 8367 817 8419
rect 817 8367 833 8419
rect 833 8367 885 8419
rect 885 8367 901 8419
rect 901 8367 953 8419
rect 953 8367 969 8419
rect 969 8367 1021 8419
rect 1021 8367 1037 8419
rect 1037 8367 1089 8419
rect 1089 8367 1105 8419
rect 1105 8367 1157 8419
rect 1157 8367 1173 8419
rect 1173 8367 1225 8419
rect 1225 8367 1241 8419
rect 1241 8367 1263 8419
rect 727 8355 1263 8367
rect 727 8303 749 8355
rect 749 8303 765 8355
rect 765 8303 817 8355
rect 817 8303 833 8355
rect 833 8303 885 8355
rect 885 8303 901 8355
rect 901 8303 953 8355
rect 953 8303 969 8355
rect 969 8303 1021 8355
rect 1021 8303 1037 8355
rect 1037 8303 1089 8355
rect 1089 8303 1105 8355
rect 1105 8303 1157 8355
rect 1157 8303 1173 8355
rect 1173 8303 1225 8355
rect 1225 8303 1241 8355
rect 1241 8303 1263 8355
rect 727 8291 1263 8303
rect 727 8239 749 8291
rect 749 8239 765 8291
rect 765 8239 817 8291
rect 817 8239 833 8291
rect 833 8239 885 8291
rect 885 8239 901 8291
rect 901 8239 953 8291
rect 953 8239 969 8291
rect 969 8239 1021 8291
rect 1021 8239 1037 8291
rect 1037 8239 1089 8291
rect 1089 8239 1105 8291
rect 1105 8239 1157 8291
rect 1157 8239 1173 8291
rect 1173 8239 1225 8291
rect 1225 8239 1241 8291
rect 1241 8239 1263 8291
rect 727 8227 1263 8239
rect 727 8175 749 8227
rect 749 8175 765 8227
rect 765 8175 817 8227
rect 817 8175 833 8227
rect 833 8175 885 8227
rect 885 8175 901 8227
rect 901 8175 953 8227
rect 953 8175 969 8227
rect 969 8175 1021 8227
rect 1021 8175 1037 8227
rect 1037 8175 1089 8227
rect 1089 8175 1105 8227
rect 1105 8175 1157 8227
rect 1157 8175 1173 8227
rect 1173 8175 1225 8227
rect 1225 8175 1241 8227
rect 1241 8175 1263 8227
rect 727 8163 1263 8175
rect 727 8152 749 8163
rect 749 8152 765 8163
rect 765 8152 817 8163
rect 817 8152 833 8163
rect 833 8152 885 8163
rect 885 8152 901 8163
rect 901 8152 953 8163
rect 953 8152 969 8163
rect 969 8152 1021 8163
rect 1021 8152 1037 8163
rect 1037 8152 1089 8163
rect 1089 8152 1105 8163
rect 1105 8152 1157 8163
rect 1157 8152 1173 8163
rect 1173 8152 1225 8163
rect 1225 8152 1241 8163
rect 1241 8152 1263 8163
rect 727 8111 749 8127
rect 749 8111 765 8127
rect 765 8111 783 8127
rect 807 8111 817 8127
rect 817 8111 833 8127
rect 833 8111 863 8127
rect 887 8111 901 8127
rect 901 8111 943 8127
rect 967 8111 969 8127
rect 969 8111 1021 8127
rect 1021 8111 1023 8127
rect 1047 8111 1089 8127
rect 1089 8111 1103 8127
rect 1127 8111 1157 8127
rect 1157 8111 1173 8127
rect 1173 8111 1183 8127
rect 1207 8111 1225 8127
rect 1225 8111 1241 8127
rect 1241 8111 1263 8127
rect 727 8099 783 8111
rect 807 8099 863 8111
rect 887 8099 943 8111
rect 967 8099 1023 8111
rect 1047 8099 1103 8111
rect 1127 8099 1183 8111
rect 1207 8099 1263 8111
rect 727 8071 749 8099
rect 749 8071 765 8099
rect 765 8071 783 8099
rect 807 8071 817 8099
rect 817 8071 833 8099
rect 833 8071 863 8099
rect 887 8071 901 8099
rect 901 8071 943 8099
rect 967 8071 969 8099
rect 969 8071 1021 8099
rect 1021 8071 1023 8099
rect 1047 8071 1089 8099
rect 1089 8071 1103 8099
rect 1127 8071 1157 8099
rect 1157 8071 1173 8099
rect 1173 8071 1183 8099
rect 1207 8071 1225 8099
rect 1225 8071 1241 8099
rect 1241 8071 1263 8099
rect 727 8035 783 8046
rect 807 8035 863 8046
rect 887 8035 943 8046
rect 967 8035 1023 8046
rect 1047 8035 1103 8046
rect 1127 8035 1183 8046
rect 1207 8035 1263 8046
rect 727 7990 749 8035
rect 749 7990 765 8035
rect 765 7990 783 8035
rect 807 7990 817 8035
rect 817 7990 833 8035
rect 833 7990 863 8035
rect 887 7990 901 8035
rect 901 7990 943 8035
rect 967 7990 969 8035
rect 969 7990 1021 8035
rect 1021 7990 1023 8035
rect 1047 7990 1089 8035
rect 1089 7990 1103 8035
rect 1127 7990 1157 8035
rect 1157 7990 1173 8035
rect 1173 7990 1183 8035
rect 1207 7990 1225 8035
rect 1225 7990 1241 8035
rect 1241 7990 1263 8035
rect 727 7919 749 7965
rect 749 7919 765 7965
rect 765 7919 783 7965
rect 807 7919 817 7965
rect 817 7919 833 7965
rect 833 7919 863 7965
rect 887 7919 901 7965
rect 901 7919 943 7965
rect 967 7919 969 7965
rect 969 7919 1021 7965
rect 1021 7919 1023 7965
rect 1047 7919 1089 7965
rect 1089 7919 1103 7965
rect 1127 7919 1157 7965
rect 1157 7919 1173 7965
rect 1173 7919 1183 7965
rect 1207 7919 1225 7965
rect 1225 7919 1241 7965
rect 1241 7919 1263 7965
rect 727 7909 783 7919
rect 807 7909 863 7919
rect 887 7909 943 7919
rect 967 7909 1023 7919
rect 1047 7909 1103 7919
rect 1127 7909 1183 7919
rect 1207 7909 1263 7919
rect 727 7855 749 7884
rect 749 7855 765 7884
rect 765 7855 783 7884
rect 807 7855 817 7884
rect 817 7855 833 7884
rect 833 7855 863 7884
rect 887 7855 901 7884
rect 901 7855 943 7884
rect 967 7855 969 7884
rect 969 7855 1021 7884
rect 1021 7855 1023 7884
rect 1047 7855 1089 7884
rect 1089 7855 1103 7884
rect 1127 7855 1157 7884
rect 1157 7855 1173 7884
rect 1173 7855 1183 7884
rect 1207 7855 1225 7884
rect 1225 7855 1241 7884
rect 1241 7855 1263 7884
rect 727 7843 783 7855
rect 807 7843 863 7855
rect 887 7843 943 7855
rect 967 7843 1023 7855
rect 1047 7843 1103 7855
rect 1127 7843 1183 7855
rect 1207 7843 1263 7855
rect 727 7828 749 7843
rect 749 7828 765 7843
rect 765 7828 783 7843
rect 807 7828 817 7843
rect 817 7828 833 7843
rect 833 7828 863 7843
rect 887 7828 901 7843
rect 901 7828 943 7843
rect 967 7828 969 7843
rect 969 7828 1021 7843
rect 1021 7828 1023 7843
rect 1047 7828 1089 7843
rect 1089 7828 1103 7843
rect 1127 7828 1157 7843
rect 1157 7828 1173 7843
rect 1173 7828 1183 7843
rect 1207 7828 1225 7843
rect 1225 7828 1241 7843
rect 1241 7828 1263 7843
rect 727 7791 749 7803
rect 749 7791 765 7803
rect 765 7791 783 7803
rect 807 7791 817 7803
rect 817 7791 833 7803
rect 833 7791 863 7803
rect 887 7791 901 7803
rect 901 7791 943 7803
rect 967 7791 969 7803
rect 969 7791 1021 7803
rect 1021 7791 1023 7803
rect 1047 7791 1089 7803
rect 1089 7791 1103 7803
rect 1127 7791 1157 7803
rect 1157 7791 1173 7803
rect 1173 7791 1183 7803
rect 1207 7791 1225 7803
rect 1225 7791 1241 7803
rect 1241 7791 1263 7803
rect 727 7779 783 7791
rect 807 7779 863 7791
rect 887 7779 943 7791
rect 967 7779 1023 7791
rect 1047 7779 1103 7791
rect 1127 7779 1183 7791
rect 1207 7779 1263 7791
rect 727 7747 749 7779
rect 749 7747 765 7779
rect 765 7747 783 7779
rect 807 7747 817 7779
rect 817 7747 833 7779
rect 833 7747 863 7779
rect 887 7747 901 7779
rect 901 7747 943 7779
rect 967 7747 969 7779
rect 969 7747 1021 7779
rect 1021 7747 1023 7779
rect 1047 7747 1089 7779
rect 1089 7747 1103 7779
rect 1127 7747 1157 7779
rect 1157 7747 1173 7779
rect 1173 7747 1183 7779
rect 1207 7747 1225 7779
rect 1225 7747 1241 7779
rect 1241 7747 1263 7779
rect 727 7715 783 7722
rect 807 7715 863 7722
rect 887 7715 943 7722
rect 967 7715 1023 7722
rect 1047 7715 1103 7722
rect 1127 7715 1183 7722
rect 1207 7715 1263 7722
rect 727 7666 749 7715
rect 749 7666 765 7715
rect 765 7666 783 7715
rect 807 7666 817 7715
rect 817 7666 833 7715
rect 833 7666 863 7715
rect 887 7666 901 7715
rect 901 7666 943 7715
rect 967 7666 969 7715
rect 969 7666 1021 7715
rect 1021 7666 1023 7715
rect 1047 7666 1089 7715
rect 1089 7666 1103 7715
rect 1127 7666 1157 7715
rect 1157 7666 1173 7715
rect 1173 7666 1183 7715
rect 1207 7666 1225 7715
rect 1225 7666 1241 7715
rect 1241 7666 1263 7715
rect 727 6449 749 6498
rect 749 6449 765 6498
rect 765 6449 817 6498
rect 817 6449 833 6498
rect 833 6449 885 6498
rect 885 6449 901 6498
rect 901 6449 953 6498
rect 953 6449 969 6498
rect 969 6449 1021 6498
rect 1021 6449 1037 6498
rect 1037 6449 1089 6498
rect 1089 6449 1105 6498
rect 1105 6449 1157 6498
rect 1157 6449 1173 6498
rect 1173 6449 1225 6498
rect 1225 6449 1241 6498
rect 1241 6449 1263 6498
rect 727 6437 1263 6449
rect 727 6385 749 6437
rect 749 6385 765 6437
rect 765 6385 817 6437
rect 817 6385 833 6437
rect 833 6385 885 6437
rect 885 6385 901 6437
rect 901 6385 953 6437
rect 953 6385 969 6437
rect 969 6385 1021 6437
rect 1021 6385 1037 6437
rect 1037 6385 1089 6437
rect 1089 6385 1105 6437
rect 1105 6385 1157 6437
rect 1157 6385 1173 6437
rect 1173 6385 1225 6437
rect 1225 6385 1241 6437
rect 1241 6385 1263 6437
rect 727 6373 1263 6385
rect 727 6321 749 6373
rect 749 6321 765 6373
rect 765 6321 817 6373
rect 817 6321 833 6373
rect 833 6321 885 6373
rect 885 6321 901 6373
rect 901 6321 953 6373
rect 953 6321 969 6373
rect 969 6321 1021 6373
rect 1021 6321 1037 6373
rect 1037 6321 1089 6373
rect 1089 6321 1105 6373
rect 1105 6321 1157 6373
rect 1157 6321 1173 6373
rect 1173 6321 1225 6373
rect 1225 6321 1241 6373
rect 1241 6321 1263 6373
rect 727 6309 1263 6321
rect 727 6257 749 6309
rect 749 6257 765 6309
rect 765 6257 817 6309
rect 817 6257 833 6309
rect 833 6257 885 6309
rect 885 6257 901 6309
rect 901 6257 953 6309
rect 953 6257 969 6309
rect 969 6257 1021 6309
rect 1021 6257 1037 6309
rect 1037 6257 1089 6309
rect 1089 6257 1105 6309
rect 1105 6257 1157 6309
rect 1157 6257 1173 6309
rect 1173 6257 1225 6309
rect 1225 6257 1241 6309
rect 1241 6257 1263 6309
rect 727 6245 1263 6257
rect 727 6193 749 6245
rect 749 6193 765 6245
rect 765 6193 817 6245
rect 817 6193 833 6245
rect 833 6193 885 6245
rect 885 6193 901 6245
rect 901 6193 953 6245
rect 953 6193 969 6245
rect 969 6193 1021 6245
rect 1021 6193 1037 6245
rect 1037 6193 1089 6245
rect 1089 6193 1105 6245
rect 1105 6193 1157 6245
rect 1157 6193 1173 6245
rect 1173 6193 1225 6245
rect 1225 6193 1241 6245
rect 1241 6193 1263 6245
rect 727 6181 1263 6193
rect 727 6129 749 6181
rect 749 6129 765 6181
rect 765 6129 817 6181
rect 817 6129 833 6181
rect 833 6129 885 6181
rect 885 6129 901 6181
rect 901 6129 953 6181
rect 953 6129 969 6181
rect 969 6129 1021 6181
rect 1021 6129 1037 6181
rect 1037 6129 1089 6181
rect 1089 6129 1105 6181
rect 1105 6129 1157 6181
rect 1157 6129 1173 6181
rect 1173 6129 1225 6181
rect 1225 6129 1241 6181
rect 1241 6129 1263 6181
rect 727 6117 1263 6129
rect 727 6065 749 6117
rect 749 6065 765 6117
rect 765 6065 817 6117
rect 817 6065 833 6117
rect 833 6065 885 6117
rect 885 6065 901 6117
rect 901 6065 953 6117
rect 953 6065 969 6117
rect 969 6065 1021 6117
rect 1021 6065 1037 6117
rect 1037 6065 1089 6117
rect 1089 6065 1105 6117
rect 1105 6065 1157 6117
rect 1157 6065 1173 6117
rect 1173 6065 1225 6117
rect 1225 6065 1241 6117
rect 1241 6065 1263 6117
rect 727 6053 1263 6065
rect 727 6042 749 6053
rect 749 6042 765 6053
rect 765 6042 817 6053
rect 817 6042 833 6053
rect 833 6042 885 6053
rect 885 6042 901 6053
rect 901 6042 953 6053
rect 953 6042 969 6053
rect 969 6042 1021 6053
rect 1021 6042 1037 6053
rect 1037 6042 1089 6053
rect 1089 6042 1105 6053
rect 1105 6042 1157 6053
rect 1157 6042 1173 6053
rect 1173 6042 1225 6053
rect 1225 6042 1241 6053
rect 1241 6042 1263 6053
rect 727 6001 749 6017
rect 749 6001 765 6017
rect 765 6001 783 6017
rect 807 6001 817 6017
rect 817 6001 833 6017
rect 833 6001 863 6017
rect 887 6001 901 6017
rect 901 6001 943 6017
rect 967 6001 969 6017
rect 969 6001 1021 6017
rect 1021 6001 1023 6017
rect 1047 6001 1089 6017
rect 1089 6001 1103 6017
rect 1127 6001 1157 6017
rect 1157 6001 1173 6017
rect 1173 6001 1183 6017
rect 1207 6001 1225 6017
rect 1225 6001 1241 6017
rect 1241 6001 1263 6017
rect 727 5989 783 6001
rect 807 5989 863 6001
rect 887 5989 943 6001
rect 967 5989 1023 6001
rect 1047 5989 1103 6001
rect 1127 5989 1183 6001
rect 1207 5989 1263 6001
rect 727 5961 749 5989
rect 749 5961 765 5989
rect 765 5961 783 5989
rect 807 5961 817 5989
rect 817 5961 833 5989
rect 833 5961 863 5989
rect 887 5961 901 5989
rect 901 5961 943 5989
rect 967 5961 969 5989
rect 969 5961 1021 5989
rect 1021 5961 1023 5989
rect 1047 5961 1089 5989
rect 1089 5961 1103 5989
rect 1127 5961 1157 5989
rect 1157 5961 1173 5989
rect 1173 5961 1183 5989
rect 1207 5961 1225 5989
rect 1225 5961 1241 5989
rect 1241 5961 1263 5989
rect 727 5925 783 5936
rect 807 5925 863 5936
rect 887 5925 943 5936
rect 967 5925 1023 5936
rect 1047 5925 1103 5936
rect 1127 5925 1183 5936
rect 1207 5925 1263 5936
rect 727 5880 749 5925
rect 749 5880 765 5925
rect 765 5880 783 5925
rect 807 5880 817 5925
rect 817 5880 833 5925
rect 833 5880 863 5925
rect 887 5880 901 5925
rect 901 5880 943 5925
rect 967 5880 969 5925
rect 969 5880 1021 5925
rect 1021 5880 1023 5925
rect 1047 5880 1089 5925
rect 1089 5880 1103 5925
rect 1127 5880 1157 5925
rect 1157 5880 1173 5925
rect 1173 5880 1183 5925
rect 1207 5880 1225 5925
rect 1225 5880 1241 5925
rect 1241 5880 1263 5925
rect 727 5809 749 5855
rect 749 5809 765 5855
rect 765 5809 783 5855
rect 807 5809 817 5855
rect 817 5809 833 5855
rect 833 5809 863 5855
rect 887 5809 901 5855
rect 901 5809 943 5855
rect 967 5809 969 5855
rect 969 5809 1021 5855
rect 1021 5809 1023 5855
rect 1047 5809 1089 5855
rect 1089 5809 1103 5855
rect 1127 5809 1157 5855
rect 1157 5809 1173 5855
rect 1173 5809 1183 5855
rect 1207 5809 1225 5855
rect 1225 5809 1241 5855
rect 1241 5809 1263 5855
rect 727 5799 783 5809
rect 807 5799 863 5809
rect 887 5799 943 5809
rect 967 5799 1023 5809
rect 1047 5799 1103 5809
rect 1127 5799 1183 5809
rect 1207 5799 1263 5809
rect 727 5745 749 5774
rect 749 5745 765 5774
rect 765 5745 783 5774
rect 807 5745 817 5774
rect 817 5745 833 5774
rect 833 5745 863 5774
rect 887 5745 901 5774
rect 901 5745 943 5774
rect 967 5745 969 5774
rect 969 5745 1021 5774
rect 1021 5745 1023 5774
rect 1047 5745 1089 5774
rect 1089 5745 1103 5774
rect 1127 5745 1157 5774
rect 1157 5745 1173 5774
rect 1173 5745 1183 5774
rect 1207 5745 1225 5774
rect 1225 5745 1241 5774
rect 1241 5745 1263 5774
rect 727 5733 783 5745
rect 807 5733 863 5745
rect 887 5733 943 5745
rect 967 5733 1023 5745
rect 1047 5733 1103 5745
rect 1127 5733 1183 5745
rect 1207 5733 1263 5745
rect 727 5718 749 5733
rect 749 5718 765 5733
rect 765 5718 783 5733
rect 807 5718 817 5733
rect 817 5718 833 5733
rect 833 5718 863 5733
rect 887 5718 901 5733
rect 901 5718 943 5733
rect 967 5718 969 5733
rect 969 5718 1021 5733
rect 1021 5718 1023 5733
rect 1047 5718 1089 5733
rect 1089 5718 1103 5733
rect 1127 5718 1157 5733
rect 1157 5718 1173 5733
rect 1173 5718 1183 5733
rect 1207 5718 1225 5733
rect 1225 5718 1241 5733
rect 1241 5718 1263 5733
rect 727 5681 749 5693
rect 749 5681 765 5693
rect 765 5681 783 5693
rect 807 5681 817 5693
rect 817 5681 833 5693
rect 833 5681 863 5693
rect 887 5681 901 5693
rect 901 5681 943 5693
rect 967 5681 969 5693
rect 969 5681 1021 5693
rect 1021 5681 1023 5693
rect 1047 5681 1089 5693
rect 1089 5681 1103 5693
rect 1127 5681 1157 5693
rect 1157 5681 1173 5693
rect 1173 5681 1183 5693
rect 1207 5681 1225 5693
rect 1225 5681 1241 5693
rect 1241 5681 1263 5693
rect 727 5669 783 5681
rect 807 5669 863 5681
rect 887 5669 943 5681
rect 967 5669 1023 5681
rect 1047 5669 1103 5681
rect 1127 5669 1183 5681
rect 1207 5669 1263 5681
rect 727 5637 749 5669
rect 749 5637 765 5669
rect 765 5637 783 5669
rect 807 5637 817 5669
rect 817 5637 833 5669
rect 833 5637 863 5669
rect 887 5637 901 5669
rect 901 5637 943 5669
rect 967 5637 969 5669
rect 969 5637 1021 5669
rect 1021 5637 1023 5669
rect 1047 5637 1089 5669
rect 1089 5637 1103 5669
rect 1127 5637 1157 5669
rect 1157 5637 1173 5669
rect 1173 5637 1183 5669
rect 1207 5637 1225 5669
rect 1225 5637 1241 5669
rect 1241 5637 1263 5669
rect 727 5605 783 5612
rect 807 5605 863 5612
rect 887 5605 943 5612
rect 967 5605 1023 5612
rect 1047 5605 1103 5612
rect 1127 5605 1183 5612
rect 1207 5605 1263 5612
rect 727 5556 749 5605
rect 749 5556 765 5605
rect 765 5556 783 5605
rect 807 5556 817 5605
rect 817 5556 833 5605
rect 833 5556 863 5605
rect 887 5556 901 5605
rect 901 5556 943 5605
rect 967 5556 969 5605
rect 969 5556 1021 5605
rect 1021 5556 1023 5605
rect 1047 5556 1089 5605
rect 1089 5556 1103 5605
rect 1127 5556 1157 5605
rect 1157 5556 1173 5605
rect 1173 5556 1183 5605
rect 1207 5556 1225 5605
rect 1225 5556 1241 5605
rect 1241 5556 1263 5605
rect 727 4385 749 4434
rect 749 4385 765 4434
rect 765 4385 817 4434
rect 817 4385 833 4434
rect 833 4385 885 4434
rect 885 4385 901 4434
rect 901 4385 953 4434
rect 953 4385 969 4434
rect 969 4385 1021 4434
rect 1021 4385 1037 4434
rect 1037 4385 1089 4434
rect 1089 4385 1105 4434
rect 1105 4385 1157 4434
rect 1157 4385 1173 4434
rect 1173 4385 1225 4434
rect 1225 4385 1241 4434
rect 1241 4385 1263 4434
rect 727 4373 1263 4385
rect 727 4321 749 4373
rect 749 4321 765 4373
rect 765 4321 817 4373
rect 817 4321 833 4373
rect 833 4321 885 4373
rect 885 4321 901 4373
rect 901 4321 953 4373
rect 953 4321 969 4373
rect 969 4321 1021 4373
rect 1021 4321 1037 4373
rect 1037 4321 1089 4373
rect 1089 4321 1105 4373
rect 1105 4321 1157 4373
rect 1157 4321 1173 4373
rect 1173 4321 1225 4373
rect 1225 4321 1241 4373
rect 1241 4321 1263 4373
rect 727 4309 1263 4321
rect 727 4257 749 4309
rect 749 4257 765 4309
rect 765 4257 817 4309
rect 817 4257 833 4309
rect 833 4257 885 4309
rect 885 4257 901 4309
rect 901 4257 953 4309
rect 953 4257 969 4309
rect 969 4257 1021 4309
rect 1021 4257 1037 4309
rect 1037 4257 1089 4309
rect 1089 4257 1105 4309
rect 1105 4257 1157 4309
rect 1157 4257 1173 4309
rect 1173 4257 1225 4309
rect 1225 4257 1241 4309
rect 1241 4257 1263 4309
rect 727 4245 1263 4257
rect 727 4193 749 4245
rect 749 4193 765 4245
rect 765 4193 817 4245
rect 817 4193 833 4245
rect 833 4193 885 4245
rect 885 4193 901 4245
rect 901 4193 953 4245
rect 953 4193 969 4245
rect 969 4193 1021 4245
rect 1021 4193 1037 4245
rect 1037 4193 1089 4245
rect 1089 4193 1105 4245
rect 1105 4193 1157 4245
rect 1157 4193 1173 4245
rect 1173 4193 1225 4245
rect 1225 4193 1241 4245
rect 1241 4193 1263 4245
rect 727 4181 1263 4193
rect 727 4129 749 4181
rect 749 4129 765 4181
rect 765 4129 817 4181
rect 817 4129 833 4181
rect 833 4129 885 4181
rect 885 4129 901 4181
rect 901 4129 953 4181
rect 953 4129 969 4181
rect 969 4129 1021 4181
rect 1021 4129 1037 4181
rect 1037 4129 1089 4181
rect 1089 4129 1105 4181
rect 1105 4129 1157 4181
rect 1157 4129 1173 4181
rect 1173 4129 1225 4181
rect 1225 4129 1241 4181
rect 1241 4129 1263 4181
rect 727 4117 1263 4129
rect 727 4065 749 4117
rect 749 4065 765 4117
rect 765 4065 817 4117
rect 817 4065 833 4117
rect 833 4065 885 4117
rect 885 4065 901 4117
rect 901 4065 953 4117
rect 953 4065 969 4117
rect 969 4065 1021 4117
rect 1021 4065 1037 4117
rect 1037 4065 1089 4117
rect 1089 4065 1105 4117
rect 1105 4065 1157 4117
rect 1157 4065 1173 4117
rect 1173 4065 1225 4117
rect 1225 4065 1241 4117
rect 1241 4065 1263 4117
rect 727 4053 1263 4065
rect 727 4001 749 4053
rect 749 4001 765 4053
rect 765 4001 817 4053
rect 817 4001 833 4053
rect 833 4001 885 4053
rect 885 4001 901 4053
rect 901 4001 953 4053
rect 953 4001 969 4053
rect 969 4001 1021 4053
rect 1021 4001 1037 4053
rect 1037 4001 1089 4053
rect 1089 4001 1105 4053
rect 1105 4001 1157 4053
rect 1157 4001 1173 4053
rect 1173 4001 1225 4053
rect 1225 4001 1241 4053
rect 1241 4001 1263 4053
rect 727 3989 1263 4001
rect 727 3978 749 3989
rect 749 3978 765 3989
rect 765 3978 817 3989
rect 817 3978 833 3989
rect 833 3978 885 3989
rect 885 3978 901 3989
rect 901 3978 953 3989
rect 953 3978 969 3989
rect 969 3978 1021 3989
rect 1021 3978 1037 3989
rect 1037 3978 1089 3989
rect 1089 3978 1105 3989
rect 1105 3978 1157 3989
rect 1157 3978 1173 3989
rect 1173 3978 1225 3989
rect 1225 3978 1241 3989
rect 1241 3978 1263 3989
rect 727 3937 749 3953
rect 749 3937 765 3953
rect 765 3937 783 3953
rect 807 3937 817 3953
rect 817 3937 833 3953
rect 833 3937 863 3953
rect 887 3937 901 3953
rect 901 3937 943 3953
rect 967 3937 969 3953
rect 969 3937 1021 3953
rect 1021 3937 1023 3953
rect 1047 3937 1089 3953
rect 1089 3937 1103 3953
rect 1127 3937 1157 3953
rect 1157 3937 1173 3953
rect 1173 3937 1183 3953
rect 1207 3937 1225 3953
rect 1225 3937 1241 3953
rect 1241 3937 1263 3953
rect 727 3925 783 3937
rect 807 3925 863 3937
rect 887 3925 943 3937
rect 967 3925 1023 3937
rect 1047 3925 1103 3937
rect 1127 3925 1183 3937
rect 1207 3925 1263 3937
rect 727 3897 749 3925
rect 749 3897 765 3925
rect 765 3897 783 3925
rect 807 3897 817 3925
rect 817 3897 833 3925
rect 833 3897 863 3925
rect 887 3897 901 3925
rect 901 3897 943 3925
rect 967 3897 969 3925
rect 969 3897 1021 3925
rect 1021 3897 1023 3925
rect 1047 3897 1089 3925
rect 1089 3897 1103 3925
rect 1127 3897 1157 3925
rect 1157 3897 1173 3925
rect 1173 3897 1183 3925
rect 1207 3897 1225 3925
rect 1225 3897 1241 3925
rect 1241 3897 1263 3925
rect 727 3861 783 3872
rect 807 3861 863 3872
rect 887 3861 943 3872
rect 967 3861 1023 3872
rect 1047 3861 1103 3872
rect 1127 3861 1183 3872
rect 1207 3861 1263 3872
rect 727 3816 749 3861
rect 749 3816 765 3861
rect 765 3816 783 3861
rect 807 3816 817 3861
rect 817 3816 833 3861
rect 833 3816 863 3861
rect 887 3816 901 3861
rect 901 3816 943 3861
rect 967 3816 969 3861
rect 969 3816 1021 3861
rect 1021 3816 1023 3861
rect 1047 3816 1089 3861
rect 1089 3816 1103 3861
rect 1127 3816 1157 3861
rect 1157 3816 1173 3861
rect 1173 3816 1183 3861
rect 1207 3816 1225 3861
rect 1225 3816 1241 3861
rect 1241 3816 1263 3861
rect 727 3745 749 3791
rect 749 3745 765 3791
rect 765 3745 783 3791
rect 807 3745 817 3791
rect 817 3745 833 3791
rect 833 3745 863 3791
rect 887 3745 901 3791
rect 901 3745 943 3791
rect 967 3745 969 3791
rect 969 3745 1021 3791
rect 1021 3745 1023 3791
rect 1047 3745 1089 3791
rect 1089 3745 1103 3791
rect 1127 3745 1157 3791
rect 1157 3745 1173 3791
rect 1173 3745 1183 3791
rect 1207 3745 1225 3791
rect 1225 3745 1241 3791
rect 1241 3745 1263 3791
rect 727 3735 783 3745
rect 807 3735 863 3745
rect 887 3735 943 3745
rect 967 3735 1023 3745
rect 1047 3735 1103 3745
rect 1127 3735 1183 3745
rect 1207 3735 1263 3745
rect 727 3681 749 3710
rect 749 3681 765 3710
rect 765 3681 783 3710
rect 807 3681 817 3710
rect 817 3681 833 3710
rect 833 3681 863 3710
rect 887 3681 901 3710
rect 901 3681 943 3710
rect 967 3681 969 3710
rect 969 3681 1021 3710
rect 1021 3681 1023 3710
rect 1047 3681 1089 3710
rect 1089 3681 1103 3710
rect 1127 3681 1157 3710
rect 1157 3681 1173 3710
rect 1173 3681 1183 3710
rect 1207 3681 1225 3710
rect 1225 3681 1241 3710
rect 1241 3681 1263 3710
rect 727 3669 783 3681
rect 807 3669 863 3681
rect 887 3669 943 3681
rect 967 3669 1023 3681
rect 1047 3669 1103 3681
rect 1127 3669 1183 3681
rect 1207 3669 1263 3681
rect 727 3654 749 3669
rect 749 3654 765 3669
rect 765 3654 783 3669
rect 807 3654 817 3669
rect 817 3654 833 3669
rect 833 3654 863 3669
rect 887 3654 901 3669
rect 901 3654 943 3669
rect 967 3654 969 3669
rect 969 3654 1021 3669
rect 1021 3654 1023 3669
rect 1047 3654 1089 3669
rect 1089 3654 1103 3669
rect 1127 3654 1157 3669
rect 1157 3654 1173 3669
rect 1173 3654 1183 3669
rect 1207 3654 1225 3669
rect 1225 3654 1241 3669
rect 1241 3654 1263 3669
rect 727 3617 749 3629
rect 749 3617 765 3629
rect 765 3617 783 3629
rect 807 3617 817 3629
rect 817 3617 833 3629
rect 833 3617 863 3629
rect 887 3617 901 3629
rect 901 3617 943 3629
rect 967 3617 969 3629
rect 969 3617 1021 3629
rect 1021 3617 1023 3629
rect 1047 3617 1089 3629
rect 1089 3617 1103 3629
rect 1127 3617 1157 3629
rect 1157 3617 1173 3629
rect 1173 3617 1183 3629
rect 1207 3617 1225 3629
rect 1225 3617 1241 3629
rect 1241 3617 1263 3629
rect 727 3605 783 3617
rect 807 3605 863 3617
rect 887 3605 943 3617
rect 967 3605 1023 3617
rect 1047 3605 1103 3617
rect 1127 3605 1183 3617
rect 1207 3605 1263 3617
rect 727 3573 749 3605
rect 749 3573 765 3605
rect 765 3573 783 3605
rect 807 3573 817 3605
rect 817 3573 833 3605
rect 833 3573 863 3605
rect 887 3573 901 3605
rect 901 3573 943 3605
rect 967 3573 969 3605
rect 969 3573 1021 3605
rect 1021 3573 1023 3605
rect 1047 3573 1089 3605
rect 1089 3573 1103 3605
rect 1127 3573 1157 3605
rect 1157 3573 1173 3605
rect 1173 3573 1183 3605
rect 1207 3573 1225 3605
rect 1225 3573 1241 3605
rect 1241 3573 1263 3605
rect 727 3541 783 3548
rect 807 3541 863 3548
rect 887 3541 943 3548
rect 967 3541 1023 3548
rect 1047 3541 1103 3548
rect 1127 3541 1183 3548
rect 1207 3541 1263 3548
rect 727 3492 749 3541
rect 749 3492 765 3541
rect 765 3492 783 3541
rect 807 3492 817 3541
rect 817 3492 833 3541
rect 833 3492 863 3541
rect 887 3492 901 3541
rect 901 3492 943 3541
rect 967 3492 969 3541
rect 969 3492 1021 3541
rect 1021 3492 1023 3541
rect 1047 3492 1089 3541
rect 1089 3492 1103 3541
rect 1127 3492 1157 3541
rect 1157 3492 1173 3541
rect 1173 3492 1183 3541
rect 1207 3492 1225 3541
rect 1225 3492 1241 3541
rect 1241 3492 1263 3541
rect 727 2191 749 2240
rect 749 2191 765 2240
rect 765 2191 817 2240
rect 817 2191 833 2240
rect 833 2191 885 2240
rect 885 2191 901 2240
rect 901 2191 953 2240
rect 953 2191 969 2240
rect 969 2191 1021 2240
rect 1021 2191 1037 2240
rect 1037 2191 1089 2240
rect 1089 2191 1105 2240
rect 1105 2191 1157 2240
rect 1157 2191 1173 2240
rect 1173 2191 1225 2240
rect 1225 2191 1241 2240
rect 1241 2191 1263 2240
rect 727 2179 1263 2191
rect 727 2127 749 2179
rect 749 2127 765 2179
rect 765 2127 817 2179
rect 817 2127 833 2179
rect 833 2127 885 2179
rect 885 2127 901 2179
rect 901 2127 953 2179
rect 953 2127 969 2179
rect 969 2127 1021 2179
rect 1021 2127 1037 2179
rect 1037 2127 1089 2179
rect 1089 2127 1105 2179
rect 1105 2127 1157 2179
rect 1157 2127 1173 2179
rect 1173 2127 1225 2179
rect 1225 2127 1241 2179
rect 1241 2127 1263 2179
rect 727 2115 1263 2127
rect 727 2063 749 2115
rect 749 2063 765 2115
rect 765 2063 817 2115
rect 817 2063 833 2115
rect 833 2063 885 2115
rect 885 2063 901 2115
rect 901 2063 953 2115
rect 953 2063 969 2115
rect 969 2063 1021 2115
rect 1021 2063 1037 2115
rect 1037 2063 1089 2115
rect 1089 2063 1105 2115
rect 1105 2063 1157 2115
rect 1157 2063 1173 2115
rect 1173 2063 1225 2115
rect 1225 2063 1241 2115
rect 1241 2063 1263 2115
rect 727 2051 1263 2063
rect 727 1999 749 2051
rect 749 1999 765 2051
rect 765 1999 817 2051
rect 817 1999 833 2051
rect 833 1999 885 2051
rect 885 1999 901 2051
rect 901 1999 953 2051
rect 953 1999 969 2051
rect 969 1999 1021 2051
rect 1021 1999 1037 2051
rect 1037 1999 1089 2051
rect 1089 1999 1105 2051
rect 1105 1999 1157 2051
rect 1157 1999 1173 2051
rect 1173 1999 1225 2051
rect 1225 1999 1241 2051
rect 1241 1999 1263 2051
rect 727 1987 1263 1999
rect 727 1935 749 1987
rect 749 1935 765 1987
rect 765 1935 817 1987
rect 817 1935 833 1987
rect 833 1935 885 1987
rect 885 1935 901 1987
rect 901 1935 953 1987
rect 953 1935 969 1987
rect 969 1935 1021 1987
rect 1021 1935 1037 1987
rect 1037 1935 1089 1987
rect 1089 1935 1105 1987
rect 1105 1935 1157 1987
rect 1157 1935 1173 1987
rect 1173 1935 1225 1987
rect 1225 1935 1241 1987
rect 1241 1935 1263 1987
rect 727 1923 1263 1935
rect 727 1871 749 1923
rect 749 1871 765 1923
rect 765 1871 817 1923
rect 817 1871 833 1923
rect 833 1871 885 1923
rect 885 1871 901 1923
rect 901 1871 953 1923
rect 953 1871 969 1923
rect 969 1871 1021 1923
rect 1021 1871 1037 1923
rect 1037 1871 1089 1923
rect 1089 1871 1105 1923
rect 1105 1871 1157 1923
rect 1157 1871 1173 1923
rect 1173 1871 1225 1923
rect 1225 1871 1241 1923
rect 1241 1871 1263 1923
rect 727 1859 1263 1871
rect 727 1807 749 1859
rect 749 1807 765 1859
rect 765 1807 817 1859
rect 817 1807 833 1859
rect 833 1807 885 1859
rect 885 1807 901 1859
rect 901 1807 953 1859
rect 953 1807 969 1859
rect 969 1807 1021 1859
rect 1021 1807 1037 1859
rect 1037 1807 1089 1859
rect 1089 1807 1105 1859
rect 1105 1807 1157 1859
rect 1157 1807 1173 1859
rect 1173 1807 1225 1859
rect 1225 1807 1241 1859
rect 1241 1807 1263 1859
rect 727 1795 1263 1807
rect 727 1784 749 1795
rect 749 1784 765 1795
rect 765 1784 817 1795
rect 817 1784 833 1795
rect 833 1784 885 1795
rect 885 1784 901 1795
rect 901 1784 953 1795
rect 953 1784 969 1795
rect 969 1784 1021 1795
rect 1021 1784 1037 1795
rect 1037 1784 1089 1795
rect 1089 1784 1105 1795
rect 1105 1784 1157 1795
rect 1157 1784 1173 1795
rect 1173 1784 1225 1795
rect 1225 1784 1241 1795
rect 1241 1784 1263 1795
rect 727 1743 749 1759
rect 749 1743 765 1759
rect 765 1743 783 1759
rect 807 1743 817 1759
rect 817 1743 833 1759
rect 833 1743 863 1759
rect 887 1743 901 1759
rect 901 1743 943 1759
rect 967 1743 969 1759
rect 969 1743 1021 1759
rect 1021 1743 1023 1759
rect 1047 1743 1089 1759
rect 1089 1743 1103 1759
rect 1127 1743 1157 1759
rect 1157 1743 1173 1759
rect 1173 1743 1183 1759
rect 1207 1743 1225 1759
rect 1225 1743 1241 1759
rect 1241 1743 1263 1759
rect 727 1731 783 1743
rect 807 1731 863 1743
rect 887 1731 943 1743
rect 967 1731 1023 1743
rect 1047 1731 1103 1743
rect 1127 1731 1183 1743
rect 1207 1731 1263 1743
rect 727 1703 749 1731
rect 749 1703 765 1731
rect 765 1703 783 1731
rect 807 1703 817 1731
rect 817 1703 833 1731
rect 833 1703 863 1731
rect 887 1703 901 1731
rect 901 1703 943 1731
rect 967 1703 969 1731
rect 969 1703 1021 1731
rect 1021 1703 1023 1731
rect 1047 1703 1089 1731
rect 1089 1703 1103 1731
rect 1127 1703 1157 1731
rect 1157 1703 1173 1731
rect 1173 1703 1183 1731
rect 1207 1703 1225 1731
rect 1225 1703 1241 1731
rect 1241 1703 1263 1731
rect 727 1667 783 1678
rect 807 1667 863 1678
rect 887 1667 943 1678
rect 967 1667 1023 1678
rect 1047 1667 1103 1678
rect 1127 1667 1183 1678
rect 1207 1667 1263 1678
rect 727 1622 749 1667
rect 749 1622 765 1667
rect 765 1622 783 1667
rect 807 1622 817 1667
rect 817 1622 833 1667
rect 833 1622 863 1667
rect 887 1622 901 1667
rect 901 1622 943 1667
rect 967 1622 969 1667
rect 969 1622 1021 1667
rect 1021 1622 1023 1667
rect 1047 1622 1089 1667
rect 1089 1622 1103 1667
rect 1127 1622 1157 1667
rect 1157 1622 1173 1667
rect 1173 1622 1183 1667
rect 1207 1622 1225 1667
rect 1225 1622 1241 1667
rect 1241 1622 1263 1667
rect 727 1551 749 1597
rect 749 1551 765 1597
rect 765 1551 783 1597
rect 807 1551 817 1597
rect 817 1551 833 1597
rect 833 1551 863 1597
rect 887 1551 901 1597
rect 901 1551 943 1597
rect 967 1551 969 1597
rect 969 1551 1021 1597
rect 1021 1551 1023 1597
rect 1047 1551 1089 1597
rect 1089 1551 1103 1597
rect 1127 1551 1157 1597
rect 1157 1551 1173 1597
rect 1173 1551 1183 1597
rect 1207 1551 1225 1597
rect 1225 1551 1241 1597
rect 1241 1551 1263 1597
rect 727 1541 783 1551
rect 807 1541 863 1551
rect 887 1541 943 1551
rect 967 1541 1023 1551
rect 1047 1541 1103 1551
rect 1127 1541 1183 1551
rect 1207 1541 1263 1551
rect 727 1487 749 1516
rect 749 1487 765 1516
rect 765 1487 783 1516
rect 807 1487 817 1516
rect 817 1487 833 1516
rect 833 1487 863 1516
rect 887 1487 901 1516
rect 901 1487 943 1516
rect 967 1487 969 1516
rect 969 1487 1021 1516
rect 1021 1487 1023 1516
rect 1047 1487 1089 1516
rect 1089 1487 1103 1516
rect 1127 1487 1157 1516
rect 1157 1487 1173 1516
rect 1173 1487 1183 1516
rect 1207 1487 1225 1516
rect 1225 1487 1241 1516
rect 1241 1487 1263 1516
rect 727 1475 783 1487
rect 807 1475 863 1487
rect 887 1475 943 1487
rect 967 1475 1023 1487
rect 1047 1475 1103 1487
rect 1127 1475 1183 1487
rect 1207 1475 1263 1487
rect 727 1460 749 1475
rect 749 1460 765 1475
rect 765 1460 783 1475
rect 807 1460 817 1475
rect 817 1460 833 1475
rect 833 1460 863 1475
rect 887 1460 901 1475
rect 901 1460 943 1475
rect 967 1460 969 1475
rect 969 1460 1021 1475
rect 1021 1460 1023 1475
rect 1047 1460 1089 1475
rect 1089 1460 1103 1475
rect 1127 1460 1157 1475
rect 1157 1460 1173 1475
rect 1173 1460 1183 1475
rect 1207 1460 1225 1475
rect 1225 1460 1241 1475
rect 1241 1460 1263 1475
rect 727 1423 749 1435
rect 749 1423 765 1435
rect 765 1423 783 1435
rect 807 1423 817 1435
rect 817 1423 833 1435
rect 833 1423 863 1435
rect 887 1423 901 1435
rect 901 1423 943 1435
rect 967 1423 969 1435
rect 969 1423 1021 1435
rect 1021 1423 1023 1435
rect 1047 1423 1089 1435
rect 1089 1423 1103 1435
rect 1127 1423 1157 1435
rect 1157 1423 1173 1435
rect 1173 1423 1183 1435
rect 1207 1423 1225 1435
rect 1225 1423 1241 1435
rect 1241 1423 1263 1435
rect 727 1411 783 1423
rect 807 1411 863 1423
rect 887 1411 943 1423
rect 967 1411 1023 1423
rect 1047 1411 1103 1423
rect 1127 1411 1183 1423
rect 1207 1411 1263 1423
rect 727 1379 749 1411
rect 749 1379 765 1411
rect 765 1379 783 1411
rect 807 1379 817 1411
rect 817 1379 833 1411
rect 833 1379 863 1411
rect 887 1379 901 1411
rect 901 1379 943 1411
rect 967 1379 969 1411
rect 969 1379 1021 1411
rect 1021 1379 1023 1411
rect 1047 1379 1089 1411
rect 1089 1379 1103 1411
rect 1127 1379 1157 1411
rect 1157 1379 1173 1411
rect 1173 1379 1183 1411
rect 1207 1379 1225 1411
rect 1225 1379 1241 1411
rect 1241 1379 1263 1411
rect 727 1347 783 1354
rect 807 1347 863 1354
rect 887 1347 943 1354
rect 967 1347 1023 1354
rect 1047 1347 1103 1354
rect 1127 1347 1183 1354
rect 1207 1347 1263 1354
rect 727 1298 749 1347
rect 749 1298 765 1347
rect 765 1298 783 1347
rect 807 1298 817 1347
rect 817 1298 833 1347
rect 833 1298 863 1347
rect 887 1298 901 1347
rect 901 1298 943 1347
rect 967 1298 969 1347
rect 969 1298 1021 1347
rect 1021 1298 1023 1347
rect 1047 1298 1089 1347
rect 1089 1298 1103 1347
rect 1127 1298 1157 1347
rect 1157 1298 1173 1347
rect 1173 1298 1183 1347
rect 1207 1298 1225 1347
rect 1225 1298 1241 1347
rect 1241 1298 1263 1347
rect 704 85 760 141
rect 792 85 848 141
rect 880 85 936 141
rect 968 85 1024 141
rect 1056 85 1112 141
rect 1143 85 1199 141
rect 1230 85 1286 141
rect 704 5 760 61
rect 792 5 848 61
rect 880 5 936 61
rect 968 5 1024 61
rect 1056 5 1112 61
rect 1143 5 1199 61
rect 1230 5 1286 61
rect 1504 85 1560 141
rect 1585 85 1641 141
rect 1666 85 1722 141
rect 1504 5 1560 61
rect 1585 5 1641 61
rect 1666 5 1722 61
rect 1747 5 1883 141
rect 2127 38371 2149 38420
rect 2149 38371 2165 38420
rect 2165 38371 2217 38420
rect 2217 38371 2233 38420
rect 2233 38371 2285 38420
rect 2285 38371 2301 38420
rect 2301 38371 2353 38420
rect 2353 38371 2369 38420
rect 2369 38371 2421 38420
rect 2421 38371 2437 38420
rect 2437 38371 2489 38420
rect 2489 38371 2505 38420
rect 2505 38371 2557 38420
rect 2557 38371 2573 38420
rect 2573 38371 2625 38420
rect 2625 38371 2641 38420
rect 2641 38371 2663 38420
rect 2127 38359 2663 38371
rect 2127 38307 2149 38359
rect 2149 38307 2165 38359
rect 2165 38307 2217 38359
rect 2217 38307 2233 38359
rect 2233 38307 2285 38359
rect 2285 38307 2301 38359
rect 2301 38307 2353 38359
rect 2353 38307 2369 38359
rect 2369 38307 2421 38359
rect 2421 38307 2437 38359
rect 2437 38307 2489 38359
rect 2489 38307 2505 38359
rect 2505 38307 2557 38359
rect 2557 38307 2573 38359
rect 2573 38307 2625 38359
rect 2625 38307 2641 38359
rect 2641 38307 2663 38359
rect 2127 38295 2663 38307
rect 2127 38243 2149 38295
rect 2149 38243 2165 38295
rect 2165 38243 2217 38295
rect 2217 38243 2233 38295
rect 2233 38243 2285 38295
rect 2285 38243 2301 38295
rect 2301 38243 2353 38295
rect 2353 38243 2369 38295
rect 2369 38243 2421 38295
rect 2421 38243 2437 38295
rect 2437 38243 2489 38295
rect 2489 38243 2505 38295
rect 2505 38243 2557 38295
rect 2557 38243 2573 38295
rect 2573 38243 2625 38295
rect 2625 38243 2641 38295
rect 2641 38243 2663 38295
rect 2127 38231 2663 38243
rect 2127 38179 2149 38231
rect 2149 38179 2165 38231
rect 2165 38179 2217 38231
rect 2217 38179 2233 38231
rect 2233 38179 2285 38231
rect 2285 38179 2301 38231
rect 2301 38179 2353 38231
rect 2353 38179 2369 38231
rect 2369 38179 2421 38231
rect 2421 38179 2437 38231
rect 2437 38179 2489 38231
rect 2489 38179 2505 38231
rect 2505 38179 2557 38231
rect 2557 38179 2573 38231
rect 2573 38179 2625 38231
rect 2625 38179 2641 38231
rect 2641 38179 2663 38231
rect 2127 38167 2663 38179
rect 2127 38115 2149 38167
rect 2149 38115 2165 38167
rect 2165 38115 2217 38167
rect 2217 38115 2233 38167
rect 2233 38115 2285 38167
rect 2285 38115 2301 38167
rect 2301 38115 2353 38167
rect 2353 38115 2369 38167
rect 2369 38115 2421 38167
rect 2421 38115 2437 38167
rect 2437 38115 2489 38167
rect 2489 38115 2505 38167
rect 2505 38115 2557 38167
rect 2557 38115 2573 38167
rect 2573 38115 2625 38167
rect 2625 38115 2641 38167
rect 2641 38115 2663 38167
rect 2127 38103 2663 38115
rect 2127 38051 2149 38103
rect 2149 38051 2165 38103
rect 2165 38051 2217 38103
rect 2217 38051 2233 38103
rect 2233 38051 2285 38103
rect 2285 38051 2301 38103
rect 2301 38051 2353 38103
rect 2353 38051 2369 38103
rect 2369 38051 2421 38103
rect 2421 38051 2437 38103
rect 2437 38051 2489 38103
rect 2489 38051 2505 38103
rect 2505 38051 2557 38103
rect 2557 38051 2573 38103
rect 2573 38051 2625 38103
rect 2625 38051 2641 38103
rect 2641 38051 2663 38103
rect 2127 38039 2663 38051
rect 2127 37987 2149 38039
rect 2149 37987 2165 38039
rect 2165 37987 2217 38039
rect 2217 37987 2233 38039
rect 2233 37987 2285 38039
rect 2285 37987 2301 38039
rect 2301 37987 2353 38039
rect 2353 37987 2369 38039
rect 2369 37987 2421 38039
rect 2421 37987 2437 38039
rect 2437 37987 2489 38039
rect 2489 37987 2505 38039
rect 2505 37987 2557 38039
rect 2557 37987 2573 38039
rect 2573 37987 2625 38039
rect 2625 37987 2641 38039
rect 2641 37987 2663 38039
rect 2127 37975 2663 37987
rect 2127 37964 2149 37975
rect 2149 37964 2165 37975
rect 2165 37964 2217 37975
rect 2217 37964 2233 37975
rect 2233 37964 2285 37975
rect 2285 37964 2301 37975
rect 2301 37964 2353 37975
rect 2353 37964 2369 37975
rect 2369 37964 2421 37975
rect 2421 37964 2437 37975
rect 2437 37964 2489 37975
rect 2489 37964 2505 37975
rect 2505 37964 2557 37975
rect 2557 37964 2573 37975
rect 2573 37964 2625 37975
rect 2625 37964 2641 37975
rect 2641 37964 2663 37975
rect 2127 37923 2149 37939
rect 2149 37923 2165 37939
rect 2165 37923 2183 37939
rect 2207 37923 2217 37939
rect 2217 37923 2233 37939
rect 2233 37923 2263 37939
rect 2287 37923 2301 37939
rect 2301 37923 2343 37939
rect 2367 37923 2369 37939
rect 2369 37923 2421 37939
rect 2421 37923 2423 37939
rect 2447 37923 2489 37939
rect 2489 37923 2503 37939
rect 2527 37923 2557 37939
rect 2557 37923 2573 37939
rect 2573 37923 2583 37939
rect 2607 37923 2625 37939
rect 2625 37923 2641 37939
rect 2641 37923 2663 37939
rect 2127 37911 2183 37923
rect 2207 37911 2263 37923
rect 2287 37911 2343 37923
rect 2367 37911 2423 37923
rect 2447 37911 2503 37923
rect 2527 37911 2583 37923
rect 2607 37911 2663 37923
rect 2127 37883 2149 37911
rect 2149 37883 2165 37911
rect 2165 37883 2183 37911
rect 2207 37883 2217 37911
rect 2217 37883 2233 37911
rect 2233 37883 2263 37911
rect 2287 37883 2301 37911
rect 2301 37883 2343 37911
rect 2367 37883 2369 37911
rect 2369 37883 2421 37911
rect 2421 37883 2423 37911
rect 2447 37883 2489 37911
rect 2489 37883 2503 37911
rect 2527 37883 2557 37911
rect 2557 37883 2573 37911
rect 2573 37883 2583 37911
rect 2607 37883 2625 37911
rect 2625 37883 2641 37911
rect 2641 37883 2663 37911
rect 2127 37847 2183 37858
rect 2207 37847 2263 37858
rect 2287 37847 2343 37858
rect 2367 37847 2423 37858
rect 2447 37847 2503 37858
rect 2527 37847 2583 37858
rect 2607 37847 2663 37858
rect 2127 37802 2149 37847
rect 2149 37802 2165 37847
rect 2165 37802 2183 37847
rect 2207 37802 2217 37847
rect 2217 37802 2233 37847
rect 2233 37802 2263 37847
rect 2287 37802 2301 37847
rect 2301 37802 2343 37847
rect 2367 37802 2369 37847
rect 2369 37802 2421 37847
rect 2421 37802 2423 37847
rect 2447 37802 2489 37847
rect 2489 37802 2503 37847
rect 2527 37802 2557 37847
rect 2557 37802 2573 37847
rect 2573 37802 2583 37847
rect 2607 37802 2625 37847
rect 2625 37802 2641 37847
rect 2641 37802 2663 37847
rect 2127 37731 2149 37777
rect 2149 37731 2165 37777
rect 2165 37731 2183 37777
rect 2207 37731 2217 37777
rect 2217 37731 2233 37777
rect 2233 37731 2263 37777
rect 2287 37731 2301 37777
rect 2301 37731 2343 37777
rect 2367 37731 2369 37777
rect 2369 37731 2421 37777
rect 2421 37731 2423 37777
rect 2447 37731 2489 37777
rect 2489 37731 2503 37777
rect 2527 37731 2557 37777
rect 2557 37731 2573 37777
rect 2573 37731 2583 37777
rect 2607 37731 2625 37777
rect 2625 37731 2641 37777
rect 2641 37731 2663 37777
rect 2127 37721 2183 37731
rect 2207 37721 2263 37731
rect 2287 37721 2343 37731
rect 2367 37721 2423 37731
rect 2447 37721 2503 37731
rect 2527 37721 2583 37731
rect 2607 37721 2663 37731
rect 2127 37667 2149 37696
rect 2149 37667 2165 37696
rect 2165 37667 2183 37696
rect 2207 37667 2217 37696
rect 2217 37667 2233 37696
rect 2233 37667 2263 37696
rect 2287 37667 2301 37696
rect 2301 37667 2343 37696
rect 2367 37667 2369 37696
rect 2369 37667 2421 37696
rect 2421 37667 2423 37696
rect 2447 37667 2489 37696
rect 2489 37667 2503 37696
rect 2527 37667 2557 37696
rect 2557 37667 2573 37696
rect 2573 37667 2583 37696
rect 2607 37667 2625 37696
rect 2625 37667 2641 37696
rect 2641 37667 2663 37696
rect 2127 37655 2183 37667
rect 2207 37655 2263 37667
rect 2287 37655 2343 37667
rect 2367 37655 2423 37667
rect 2447 37655 2503 37667
rect 2527 37655 2583 37667
rect 2607 37655 2663 37667
rect 2127 37640 2149 37655
rect 2149 37640 2165 37655
rect 2165 37640 2183 37655
rect 2207 37640 2217 37655
rect 2217 37640 2233 37655
rect 2233 37640 2263 37655
rect 2287 37640 2301 37655
rect 2301 37640 2343 37655
rect 2367 37640 2369 37655
rect 2369 37640 2421 37655
rect 2421 37640 2423 37655
rect 2447 37640 2489 37655
rect 2489 37640 2503 37655
rect 2527 37640 2557 37655
rect 2557 37640 2573 37655
rect 2573 37640 2583 37655
rect 2607 37640 2625 37655
rect 2625 37640 2641 37655
rect 2641 37640 2663 37655
rect 2127 37603 2149 37615
rect 2149 37603 2165 37615
rect 2165 37603 2183 37615
rect 2207 37603 2217 37615
rect 2217 37603 2233 37615
rect 2233 37603 2263 37615
rect 2287 37603 2301 37615
rect 2301 37603 2343 37615
rect 2367 37603 2369 37615
rect 2369 37603 2421 37615
rect 2421 37603 2423 37615
rect 2447 37603 2489 37615
rect 2489 37603 2503 37615
rect 2527 37603 2557 37615
rect 2557 37603 2573 37615
rect 2573 37603 2583 37615
rect 2607 37603 2625 37615
rect 2625 37603 2641 37615
rect 2641 37603 2663 37615
rect 2127 37591 2183 37603
rect 2207 37591 2263 37603
rect 2287 37591 2343 37603
rect 2367 37591 2423 37603
rect 2447 37591 2503 37603
rect 2527 37591 2583 37603
rect 2607 37591 2663 37603
rect 2127 37559 2149 37591
rect 2149 37559 2165 37591
rect 2165 37559 2183 37591
rect 2207 37559 2217 37591
rect 2217 37559 2233 37591
rect 2233 37559 2263 37591
rect 2287 37559 2301 37591
rect 2301 37559 2343 37591
rect 2367 37559 2369 37591
rect 2369 37559 2421 37591
rect 2421 37559 2423 37591
rect 2447 37559 2489 37591
rect 2489 37559 2503 37591
rect 2527 37559 2557 37591
rect 2557 37559 2573 37591
rect 2573 37559 2583 37591
rect 2607 37559 2625 37591
rect 2625 37559 2641 37591
rect 2641 37559 2663 37591
rect 2127 37527 2183 37534
rect 2207 37527 2263 37534
rect 2287 37527 2343 37534
rect 2367 37527 2423 37534
rect 2447 37527 2503 37534
rect 2527 37527 2583 37534
rect 2607 37527 2663 37534
rect 2127 37478 2149 37527
rect 2149 37478 2165 37527
rect 2165 37478 2183 37527
rect 2207 37478 2217 37527
rect 2217 37478 2233 37527
rect 2233 37478 2263 37527
rect 2287 37478 2301 37527
rect 2301 37478 2343 37527
rect 2367 37478 2369 37527
rect 2369 37478 2421 37527
rect 2421 37478 2423 37527
rect 2447 37478 2489 37527
rect 2489 37478 2503 37527
rect 2527 37478 2557 37527
rect 2557 37478 2573 37527
rect 2573 37478 2583 37527
rect 2607 37478 2625 37527
rect 2625 37478 2641 37527
rect 2641 37478 2663 37527
rect 2127 36317 2149 36366
rect 2149 36317 2165 36366
rect 2165 36317 2217 36366
rect 2217 36317 2233 36366
rect 2233 36317 2285 36366
rect 2285 36317 2301 36366
rect 2301 36317 2353 36366
rect 2353 36317 2369 36366
rect 2369 36317 2421 36366
rect 2421 36317 2437 36366
rect 2437 36317 2489 36366
rect 2489 36317 2505 36366
rect 2505 36317 2557 36366
rect 2557 36317 2573 36366
rect 2573 36317 2625 36366
rect 2625 36317 2641 36366
rect 2641 36317 2663 36366
rect 2127 36305 2663 36317
rect 2127 36253 2149 36305
rect 2149 36253 2165 36305
rect 2165 36253 2217 36305
rect 2217 36253 2233 36305
rect 2233 36253 2285 36305
rect 2285 36253 2301 36305
rect 2301 36253 2353 36305
rect 2353 36253 2369 36305
rect 2369 36253 2421 36305
rect 2421 36253 2437 36305
rect 2437 36253 2489 36305
rect 2489 36253 2505 36305
rect 2505 36253 2557 36305
rect 2557 36253 2573 36305
rect 2573 36253 2625 36305
rect 2625 36253 2641 36305
rect 2641 36253 2663 36305
rect 2127 36241 2663 36253
rect 2127 36189 2149 36241
rect 2149 36189 2165 36241
rect 2165 36189 2217 36241
rect 2217 36189 2233 36241
rect 2233 36189 2285 36241
rect 2285 36189 2301 36241
rect 2301 36189 2353 36241
rect 2353 36189 2369 36241
rect 2369 36189 2421 36241
rect 2421 36189 2437 36241
rect 2437 36189 2489 36241
rect 2489 36189 2505 36241
rect 2505 36189 2557 36241
rect 2557 36189 2573 36241
rect 2573 36189 2625 36241
rect 2625 36189 2641 36241
rect 2641 36189 2663 36241
rect 2127 36177 2663 36189
rect 2127 36125 2149 36177
rect 2149 36125 2165 36177
rect 2165 36125 2217 36177
rect 2217 36125 2233 36177
rect 2233 36125 2285 36177
rect 2285 36125 2301 36177
rect 2301 36125 2353 36177
rect 2353 36125 2369 36177
rect 2369 36125 2421 36177
rect 2421 36125 2437 36177
rect 2437 36125 2489 36177
rect 2489 36125 2505 36177
rect 2505 36125 2557 36177
rect 2557 36125 2573 36177
rect 2573 36125 2625 36177
rect 2625 36125 2641 36177
rect 2641 36125 2663 36177
rect 2127 36113 2663 36125
rect 2127 36061 2149 36113
rect 2149 36061 2165 36113
rect 2165 36061 2217 36113
rect 2217 36061 2233 36113
rect 2233 36061 2285 36113
rect 2285 36061 2301 36113
rect 2301 36061 2353 36113
rect 2353 36061 2369 36113
rect 2369 36061 2421 36113
rect 2421 36061 2437 36113
rect 2437 36061 2489 36113
rect 2489 36061 2505 36113
rect 2505 36061 2557 36113
rect 2557 36061 2573 36113
rect 2573 36061 2625 36113
rect 2625 36061 2641 36113
rect 2641 36061 2663 36113
rect 2127 36049 2663 36061
rect 2127 35997 2149 36049
rect 2149 35997 2165 36049
rect 2165 35997 2217 36049
rect 2217 35997 2233 36049
rect 2233 35997 2285 36049
rect 2285 35997 2301 36049
rect 2301 35997 2353 36049
rect 2353 35997 2369 36049
rect 2369 35997 2421 36049
rect 2421 35997 2437 36049
rect 2437 35997 2489 36049
rect 2489 35997 2505 36049
rect 2505 35997 2557 36049
rect 2557 35997 2573 36049
rect 2573 35997 2625 36049
rect 2625 35997 2641 36049
rect 2641 35997 2663 36049
rect 2127 35985 2663 35997
rect 2127 35933 2149 35985
rect 2149 35933 2165 35985
rect 2165 35933 2217 35985
rect 2217 35933 2233 35985
rect 2233 35933 2285 35985
rect 2285 35933 2301 35985
rect 2301 35933 2353 35985
rect 2353 35933 2369 35985
rect 2369 35933 2421 35985
rect 2421 35933 2437 35985
rect 2437 35933 2489 35985
rect 2489 35933 2505 35985
rect 2505 35933 2557 35985
rect 2557 35933 2573 35985
rect 2573 35933 2625 35985
rect 2625 35933 2641 35985
rect 2641 35933 2663 35985
rect 2127 35921 2663 35933
rect 2127 35910 2149 35921
rect 2149 35910 2165 35921
rect 2165 35910 2217 35921
rect 2217 35910 2233 35921
rect 2233 35910 2285 35921
rect 2285 35910 2301 35921
rect 2301 35910 2353 35921
rect 2353 35910 2369 35921
rect 2369 35910 2421 35921
rect 2421 35910 2437 35921
rect 2437 35910 2489 35921
rect 2489 35910 2505 35921
rect 2505 35910 2557 35921
rect 2557 35910 2573 35921
rect 2573 35910 2625 35921
rect 2625 35910 2641 35921
rect 2641 35910 2663 35921
rect 2127 35869 2149 35885
rect 2149 35869 2165 35885
rect 2165 35869 2183 35885
rect 2207 35869 2217 35885
rect 2217 35869 2233 35885
rect 2233 35869 2263 35885
rect 2287 35869 2301 35885
rect 2301 35869 2343 35885
rect 2367 35869 2369 35885
rect 2369 35869 2421 35885
rect 2421 35869 2423 35885
rect 2447 35869 2489 35885
rect 2489 35869 2503 35885
rect 2527 35869 2557 35885
rect 2557 35869 2573 35885
rect 2573 35869 2583 35885
rect 2607 35869 2625 35885
rect 2625 35869 2641 35885
rect 2641 35869 2663 35885
rect 2127 35857 2183 35869
rect 2207 35857 2263 35869
rect 2287 35857 2343 35869
rect 2367 35857 2423 35869
rect 2447 35857 2503 35869
rect 2527 35857 2583 35869
rect 2607 35857 2663 35869
rect 2127 35829 2149 35857
rect 2149 35829 2165 35857
rect 2165 35829 2183 35857
rect 2207 35829 2217 35857
rect 2217 35829 2233 35857
rect 2233 35829 2263 35857
rect 2287 35829 2301 35857
rect 2301 35829 2343 35857
rect 2367 35829 2369 35857
rect 2369 35829 2421 35857
rect 2421 35829 2423 35857
rect 2447 35829 2489 35857
rect 2489 35829 2503 35857
rect 2527 35829 2557 35857
rect 2557 35829 2573 35857
rect 2573 35829 2583 35857
rect 2607 35829 2625 35857
rect 2625 35829 2641 35857
rect 2641 35829 2663 35857
rect 2127 35793 2183 35804
rect 2207 35793 2263 35804
rect 2287 35793 2343 35804
rect 2367 35793 2423 35804
rect 2447 35793 2503 35804
rect 2527 35793 2583 35804
rect 2607 35793 2663 35804
rect 2127 35748 2149 35793
rect 2149 35748 2165 35793
rect 2165 35748 2183 35793
rect 2207 35748 2217 35793
rect 2217 35748 2233 35793
rect 2233 35748 2263 35793
rect 2287 35748 2301 35793
rect 2301 35748 2343 35793
rect 2367 35748 2369 35793
rect 2369 35748 2421 35793
rect 2421 35748 2423 35793
rect 2447 35748 2489 35793
rect 2489 35748 2503 35793
rect 2527 35748 2557 35793
rect 2557 35748 2573 35793
rect 2573 35748 2583 35793
rect 2607 35748 2625 35793
rect 2625 35748 2641 35793
rect 2641 35748 2663 35793
rect 2127 35677 2149 35723
rect 2149 35677 2165 35723
rect 2165 35677 2183 35723
rect 2207 35677 2217 35723
rect 2217 35677 2233 35723
rect 2233 35677 2263 35723
rect 2287 35677 2301 35723
rect 2301 35677 2343 35723
rect 2367 35677 2369 35723
rect 2369 35677 2421 35723
rect 2421 35677 2423 35723
rect 2447 35677 2489 35723
rect 2489 35677 2503 35723
rect 2527 35677 2557 35723
rect 2557 35677 2573 35723
rect 2573 35677 2583 35723
rect 2607 35677 2625 35723
rect 2625 35677 2641 35723
rect 2641 35677 2663 35723
rect 2127 35667 2183 35677
rect 2207 35667 2263 35677
rect 2287 35667 2343 35677
rect 2367 35667 2423 35677
rect 2447 35667 2503 35677
rect 2527 35667 2583 35677
rect 2607 35667 2663 35677
rect 2127 35613 2149 35642
rect 2149 35613 2165 35642
rect 2165 35613 2183 35642
rect 2207 35613 2217 35642
rect 2217 35613 2233 35642
rect 2233 35613 2263 35642
rect 2287 35613 2301 35642
rect 2301 35613 2343 35642
rect 2367 35613 2369 35642
rect 2369 35613 2421 35642
rect 2421 35613 2423 35642
rect 2447 35613 2489 35642
rect 2489 35613 2503 35642
rect 2527 35613 2557 35642
rect 2557 35613 2573 35642
rect 2573 35613 2583 35642
rect 2607 35613 2625 35642
rect 2625 35613 2641 35642
rect 2641 35613 2663 35642
rect 2127 35601 2183 35613
rect 2207 35601 2263 35613
rect 2287 35601 2343 35613
rect 2367 35601 2423 35613
rect 2447 35601 2503 35613
rect 2527 35601 2583 35613
rect 2607 35601 2663 35613
rect 2127 35586 2149 35601
rect 2149 35586 2165 35601
rect 2165 35586 2183 35601
rect 2207 35586 2217 35601
rect 2217 35586 2233 35601
rect 2233 35586 2263 35601
rect 2287 35586 2301 35601
rect 2301 35586 2343 35601
rect 2367 35586 2369 35601
rect 2369 35586 2421 35601
rect 2421 35586 2423 35601
rect 2447 35586 2489 35601
rect 2489 35586 2503 35601
rect 2527 35586 2557 35601
rect 2557 35586 2573 35601
rect 2573 35586 2583 35601
rect 2607 35586 2625 35601
rect 2625 35586 2641 35601
rect 2641 35586 2663 35601
rect 2127 35549 2149 35561
rect 2149 35549 2165 35561
rect 2165 35549 2183 35561
rect 2207 35549 2217 35561
rect 2217 35549 2233 35561
rect 2233 35549 2263 35561
rect 2287 35549 2301 35561
rect 2301 35549 2343 35561
rect 2367 35549 2369 35561
rect 2369 35549 2421 35561
rect 2421 35549 2423 35561
rect 2447 35549 2489 35561
rect 2489 35549 2503 35561
rect 2527 35549 2557 35561
rect 2557 35549 2573 35561
rect 2573 35549 2583 35561
rect 2607 35549 2625 35561
rect 2625 35549 2641 35561
rect 2641 35549 2663 35561
rect 2127 35537 2183 35549
rect 2207 35537 2263 35549
rect 2287 35537 2343 35549
rect 2367 35537 2423 35549
rect 2447 35537 2503 35549
rect 2527 35537 2583 35549
rect 2607 35537 2663 35549
rect 2127 35505 2149 35537
rect 2149 35505 2165 35537
rect 2165 35505 2183 35537
rect 2207 35505 2217 35537
rect 2217 35505 2233 35537
rect 2233 35505 2263 35537
rect 2287 35505 2301 35537
rect 2301 35505 2343 35537
rect 2367 35505 2369 35537
rect 2369 35505 2421 35537
rect 2421 35505 2423 35537
rect 2447 35505 2489 35537
rect 2489 35505 2503 35537
rect 2527 35505 2557 35537
rect 2557 35505 2573 35537
rect 2573 35505 2583 35537
rect 2607 35505 2625 35537
rect 2625 35505 2641 35537
rect 2641 35505 2663 35537
rect 2127 35473 2183 35480
rect 2207 35473 2263 35480
rect 2287 35473 2343 35480
rect 2367 35473 2423 35480
rect 2447 35473 2503 35480
rect 2527 35473 2583 35480
rect 2607 35473 2663 35480
rect 2127 35424 2149 35473
rect 2149 35424 2165 35473
rect 2165 35424 2183 35473
rect 2207 35424 2217 35473
rect 2217 35424 2233 35473
rect 2233 35424 2263 35473
rect 2287 35424 2301 35473
rect 2301 35424 2343 35473
rect 2367 35424 2369 35473
rect 2369 35424 2421 35473
rect 2421 35424 2423 35473
rect 2447 35424 2489 35473
rect 2489 35424 2503 35473
rect 2527 35424 2557 35473
rect 2557 35424 2573 35473
rect 2573 35424 2583 35473
rect 2607 35424 2625 35473
rect 2625 35424 2641 35473
rect 2641 35424 2663 35473
rect 2127 34098 2149 34147
rect 2149 34098 2165 34147
rect 2165 34098 2217 34147
rect 2217 34098 2233 34147
rect 2233 34098 2285 34147
rect 2285 34098 2301 34147
rect 2301 34098 2353 34147
rect 2353 34098 2369 34147
rect 2369 34098 2421 34147
rect 2421 34098 2437 34147
rect 2437 34098 2489 34147
rect 2489 34098 2505 34147
rect 2505 34098 2557 34147
rect 2557 34098 2573 34147
rect 2573 34098 2625 34147
rect 2625 34098 2641 34147
rect 2641 34098 2663 34147
rect 2127 34086 2663 34098
rect 2127 34034 2149 34086
rect 2149 34034 2165 34086
rect 2165 34034 2217 34086
rect 2217 34034 2233 34086
rect 2233 34034 2285 34086
rect 2285 34034 2301 34086
rect 2301 34034 2353 34086
rect 2353 34034 2369 34086
rect 2369 34034 2421 34086
rect 2421 34034 2437 34086
rect 2437 34034 2489 34086
rect 2489 34034 2505 34086
rect 2505 34034 2557 34086
rect 2557 34034 2573 34086
rect 2573 34034 2625 34086
rect 2625 34034 2641 34086
rect 2641 34034 2663 34086
rect 2127 34022 2663 34034
rect 2127 33970 2149 34022
rect 2149 33970 2165 34022
rect 2165 33970 2217 34022
rect 2217 33970 2233 34022
rect 2233 33970 2285 34022
rect 2285 33970 2301 34022
rect 2301 33970 2353 34022
rect 2353 33970 2369 34022
rect 2369 33970 2421 34022
rect 2421 33970 2437 34022
rect 2437 33970 2489 34022
rect 2489 33970 2505 34022
rect 2505 33970 2557 34022
rect 2557 33970 2573 34022
rect 2573 33970 2625 34022
rect 2625 33970 2641 34022
rect 2641 33970 2663 34022
rect 2127 33958 2663 33970
rect 2127 33906 2149 33958
rect 2149 33906 2165 33958
rect 2165 33906 2217 33958
rect 2217 33906 2233 33958
rect 2233 33906 2285 33958
rect 2285 33906 2301 33958
rect 2301 33906 2353 33958
rect 2353 33906 2369 33958
rect 2369 33906 2421 33958
rect 2421 33906 2437 33958
rect 2437 33906 2489 33958
rect 2489 33906 2505 33958
rect 2505 33906 2557 33958
rect 2557 33906 2573 33958
rect 2573 33906 2625 33958
rect 2625 33906 2641 33958
rect 2641 33906 2663 33958
rect 2127 33894 2663 33906
rect 2127 33842 2149 33894
rect 2149 33842 2165 33894
rect 2165 33842 2217 33894
rect 2217 33842 2233 33894
rect 2233 33842 2285 33894
rect 2285 33842 2301 33894
rect 2301 33842 2353 33894
rect 2353 33842 2369 33894
rect 2369 33842 2421 33894
rect 2421 33842 2437 33894
rect 2437 33842 2489 33894
rect 2489 33842 2505 33894
rect 2505 33842 2557 33894
rect 2557 33842 2573 33894
rect 2573 33842 2625 33894
rect 2625 33842 2641 33894
rect 2641 33842 2663 33894
rect 2127 33830 2663 33842
rect 2127 33778 2149 33830
rect 2149 33778 2165 33830
rect 2165 33778 2217 33830
rect 2217 33778 2233 33830
rect 2233 33778 2285 33830
rect 2285 33778 2301 33830
rect 2301 33778 2353 33830
rect 2353 33778 2369 33830
rect 2369 33778 2421 33830
rect 2421 33778 2437 33830
rect 2437 33778 2489 33830
rect 2489 33778 2505 33830
rect 2505 33778 2557 33830
rect 2557 33778 2573 33830
rect 2573 33778 2625 33830
rect 2625 33778 2641 33830
rect 2641 33778 2663 33830
rect 2127 33766 2663 33778
rect 2127 33714 2149 33766
rect 2149 33714 2165 33766
rect 2165 33714 2217 33766
rect 2217 33714 2233 33766
rect 2233 33714 2285 33766
rect 2285 33714 2301 33766
rect 2301 33714 2353 33766
rect 2353 33714 2369 33766
rect 2369 33714 2421 33766
rect 2421 33714 2437 33766
rect 2437 33714 2489 33766
rect 2489 33714 2505 33766
rect 2505 33714 2557 33766
rect 2557 33714 2573 33766
rect 2573 33714 2625 33766
rect 2625 33714 2641 33766
rect 2641 33714 2663 33766
rect 2127 33702 2663 33714
rect 2127 33691 2149 33702
rect 2149 33691 2165 33702
rect 2165 33691 2217 33702
rect 2217 33691 2233 33702
rect 2233 33691 2285 33702
rect 2285 33691 2301 33702
rect 2301 33691 2353 33702
rect 2353 33691 2369 33702
rect 2369 33691 2421 33702
rect 2421 33691 2437 33702
rect 2437 33691 2489 33702
rect 2489 33691 2505 33702
rect 2505 33691 2557 33702
rect 2557 33691 2573 33702
rect 2573 33691 2625 33702
rect 2625 33691 2641 33702
rect 2641 33691 2663 33702
rect 2127 33650 2149 33666
rect 2149 33650 2165 33666
rect 2165 33650 2183 33666
rect 2207 33650 2217 33666
rect 2217 33650 2233 33666
rect 2233 33650 2263 33666
rect 2287 33650 2301 33666
rect 2301 33650 2343 33666
rect 2367 33650 2369 33666
rect 2369 33650 2421 33666
rect 2421 33650 2423 33666
rect 2447 33650 2489 33666
rect 2489 33650 2503 33666
rect 2527 33650 2557 33666
rect 2557 33650 2573 33666
rect 2573 33650 2583 33666
rect 2607 33650 2625 33666
rect 2625 33650 2641 33666
rect 2641 33650 2663 33666
rect 2127 33638 2183 33650
rect 2207 33638 2263 33650
rect 2287 33638 2343 33650
rect 2367 33638 2423 33650
rect 2447 33638 2503 33650
rect 2527 33638 2583 33650
rect 2607 33638 2663 33650
rect 2127 33610 2149 33638
rect 2149 33610 2165 33638
rect 2165 33610 2183 33638
rect 2207 33610 2217 33638
rect 2217 33610 2233 33638
rect 2233 33610 2263 33638
rect 2287 33610 2301 33638
rect 2301 33610 2343 33638
rect 2367 33610 2369 33638
rect 2369 33610 2421 33638
rect 2421 33610 2423 33638
rect 2447 33610 2489 33638
rect 2489 33610 2503 33638
rect 2527 33610 2557 33638
rect 2557 33610 2573 33638
rect 2573 33610 2583 33638
rect 2607 33610 2625 33638
rect 2625 33610 2641 33638
rect 2641 33610 2663 33638
rect 2127 33574 2183 33585
rect 2207 33574 2263 33585
rect 2287 33574 2343 33585
rect 2367 33574 2423 33585
rect 2447 33574 2503 33585
rect 2527 33574 2583 33585
rect 2607 33574 2663 33585
rect 2127 33529 2149 33574
rect 2149 33529 2165 33574
rect 2165 33529 2183 33574
rect 2207 33529 2217 33574
rect 2217 33529 2233 33574
rect 2233 33529 2263 33574
rect 2287 33529 2301 33574
rect 2301 33529 2343 33574
rect 2367 33529 2369 33574
rect 2369 33529 2421 33574
rect 2421 33529 2423 33574
rect 2447 33529 2489 33574
rect 2489 33529 2503 33574
rect 2527 33529 2557 33574
rect 2557 33529 2573 33574
rect 2573 33529 2583 33574
rect 2607 33529 2625 33574
rect 2625 33529 2641 33574
rect 2641 33529 2663 33574
rect 2127 33458 2149 33504
rect 2149 33458 2165 33504
rect 2165 33458 2183 33504
rect 2207 33458 2217 33504
rect 2217 33458 2233 33504
rect 2233 33458 2263 33504
rect 2287 33458 2301 33504
rect 2301 33458 2343 33504
rect 2367 33458 2369 33504
rect 2369 33458 2421 33504
rect 2421 33458 2423 33504
rect 2447 33458 2489 33504
rect 2489 33458 2503 33504
rect 2527 33458 2557 33504
rect 2557 33458 2573 33504
rect 2573 33458 2583 33504
rect 2607 33458 2625 33504
rect 2625 33458 2641 33504
rect 2641 33458 2663 33504
rect 2127 33448 2183 33458
rect 2207 33448 2263 33458
rect 2287 33448 2343 33458
rect 2367 33448 2423 33458
rect 2447 33448 2503 33458
rect 2527 33448 2583 33458
rect 2607 33448 2663 33458
rect 2127 33394 2149 33423
rect 2149 33394 2165 33423
rect 2165 33394 2183 33423
rect 2207 33394 2217 33423
rect 2217 33394 2233 33423
rect 2233 33394 2263 33423
rect 2287 33394 2301 33423
rect 2301 33394 2343 33423
rect 2367 33394 2369 33423
rect 2369 33394 2421 33423
rect 2421 33394 2423 33423
rect 2447 33394 2489 33423
rect 2489 33394 2503 33423
rect 2527 33394 2557 33423
rect 2557 33394 2573 33423
rect 2573 33394 2583 33423
rect 2607 33394 2625 33423
rect 2625 33394 2641 33423
rect 2641 33394 2663 33423
rect 2127 33382 2183 33394
rect 2207 33382 2263 33394
rect 2287 33382 2343 33394
rect 2367 33382 2423 33394
rect 2447 33382 2503 33394
rect 2527 33382 2583 33394
rect 2607 33382 2663 33394
rect 2127 33367 2149 33382
rect 2149 33367 2165 33382
rect 2165 33367 2183 33382
rect 2207 33367 2217 33382
rect 2217 33367 2233 33382
rect 2233 33367 2263 33382
rect 2287 33367 2301 33382
rect 2301 33367 2343 33382
rect 2367 33367 2369 33382
rect 2369 33367 2421 33382
rect 2421 33367 2423 33382
rect 2447 33367 2489 33382
rect 2489 33367 2503 33382
rect 2527 33367 2557 33382
rect 2557 33367 2573 33382
rect 2573 33367 2583 33382
rect 2607 33367 2625 33382
rect 2625 33367 2641 33382
rect 2641 33367 2663 33382
rect 2127 33330 2149 33342
rect 2149 33330 2165 33342
rect 2165 33330 2183 33342
rect 2207 33330 2217 33342
rect 2217 33330 2233 33342
rect 2233 33330 2263 33342
rect 2287 33330 2301 33342
rect 2301 33330 2343 33342
rect 2367 33330 2369 33342
rect 2369 33330 2421 33342
rect 2421 33330 2423 33342
rect 2447 33330 2489 33342
rect 2489 33330 2503 33342
rect 2527 33330 2557 33342
rect 2557 33330 2573 33342
rect 2573 33330 2583 33342
rect 2607 33330 2625 33342
rect 2625 33330 2641 33342
rect 2641 33330 2663 33342
rect 2127 33318 2183 33330
rect 2207 33318 2263 33330
rect 2287 33318 2343 33330
rect 2367 33318 2423 33330
rect 2447 33318 2503 33330
rect 2527 33318 2583 33330
rect 2607 33318 2663 33330
rect 2127 33286 2149 33318
rect 2149 33286 2165 33318
rect 2165 33286 2183 33318
rect 2207 33286 2217 33318
rect 2217 33286 2233 33318
rect 2233 33286 2263 33318
rect 2287 33286 2301 33318
rect 2301 33286 2343 33318
rect 2367 33286 2369 33318
rect 2369 33286 2421 33318
rect 2421 33286 2423 33318
rect 2447 33286 2489 33318
rect 2489 33286 2503 33318
rect 2527 33286 2557 33318
rect 2557 33286 2573 33318
rect 2573 33286 2583 33318
rect 2607 33286 2625 33318
rect 2625 33286 2641 33318
rect 2641 33286 2663 33318
rect 2127 33254 2183 33261
rect 2207 33254 2263 33261
rect 2287 33254 2343 33261
rect 2367 33254 2423 33261
rect 2447 33254 2503 33261
rect 2527 33254 2583 33261
rect 2607 33254 2663 33261
rect 2127 33205 2149 33254
rect 2149 33205 2165 33254
rect 2165 33205 2183 33254
rect 2207 33205 2217 33254
rect 2217 33205 2233 33254
rect 2233 33205 2263 33254
rect 2287 33205 2301 33254
rect 2301 33205 2343 33254
rect 2367 33205 2369 33254
rect 2369 33205 2421 33254
rect 2421 33205 2423 33254
rect 2447 33205 2489 33254
rect 2489 33205 2503 33254
rect 2527 33205 2557 33254
rect 2557 33205 2573 33254
rect 2573 33205 2583 33254
rect 2607 33205 2625 33254
rect 2625 33205 2641 33254
rect 2641 33205 2663 33254
rect 2127 31969 2149 32018
rect 2149 31969 2165 32018
rect 2165 31969 2217 32018
rect 2217 31969 2233 32018
rect 2233 31969 2285 32018
rect 2285 31969 2301 32018
rect 2301 31969 2353 32018
rect 2353 31969 2369 32018
rect 2369 31969 2421 32018
rect 2421 31969 2437 32018
rect 2437 31969 2489 32018
rect 2489 31969 2505 32018
rect 2505 31969 2557 32018
rect 2557 31969 2573 32018
rect 2573 31969 2625 32018
rect 2625 31969 2641 32018
rect 2641 31969 2663 32018
rect 2127 31957 2663 31969
rect 2127 31905 2149 31957
rect 2149 31905 2165 31957
rect 2165 31905 2217 31957
rect 2217 31905 2233 31957
rect 2233 31905 2285 31957
rect 2285 31905 2301 31957
rect 2301 31905 2353 31957
rect 2353 31905 2369 31957
rect 2369 31905 2421 31957
rect 2421 31905 2437 31957
rect 2437 31905 2489 31957
rect 2489 31905 2505 31957
rect 2505 31905 2557 31957
rect 2557 31905 2573 31957
rect 2573 31905 2625 31957
rect 2625 31905 2641 31957
rect 2641 31905 2663 31957
rect 2127 31893 2663 31905
rect 2127 31841 2149 31893
rect 2149 31841 2165 31893
rect 2165 31841 2217 31893
rect 2217 31841 2233 31893
rect 2233 31841 2285 31893
rect 2285 31841 2301 31893
rect 2301 31841 2353 31893
rect 2353 31841 2369 31893
rect 2369 31841 2421 31893
rect 2421 31841 2437 31893
rect 2437 31841 2489 31893
rect 2489 31841 2505 31893
rect 2505 31841 2557 31893
rect 2557 31841 2573 31893
rect 2573 31841 2625 31893
rect 2625 31841 2641 31893
rect 2641 31841 2663 31893
rect 2127 31829 2663 31841
rect 2127 31777 2149 31829
rect 2149 31777 2165 31829
rect 2165 31777 2217 31829
rect 2217 31777 2233 31829
rect 2233 31777 2285 31829
rect 2285 31777 2301 31829
rect 2301 31777 2353 31829
rect 2353 31777 2369 31829
rect 2369 31777 2421 31829
rect 2421 31777 2437 31829
rect 2437 31777 2489 31829
rect 2489 31777 2505 31829
rect 2505 31777 2557 31829
rect 2557 31777 2573 31829
rect 2573 31777 2625 31829
rect 2625 31777 2641 31829
rect 2641 31777 2663 31829
rect 2127 31765 2663 31777
rect 2127 31713 2149 31765
rect 2149 31713 2165 31765
rect 2165 31713 2217 31765
rect 2217 31713 2233 31765
rect 2233 31713 2285 31765
rect 2285 31713 2301 31765
rect 2301 31713 2353 31765
rect 2353 31713 2369 31765
rect 2369 31713 2421 31765
rect 2421 31713 2437 31765
rect 2437 31713 2489 31765
rect 2489 31713 2505 31765
rect 2505 31713 2557 31765
rect 2557 31713 2573 31765
rect 2573 31713 2625 31765
rect 2625 31713 2641 31765
rect 2641 31713 2663 31765
rect 2127 31701 2663 31713
rect 2127 31649 2149 31701
rect 2149 31649 2165 31701
rect 2165 31649 2217 31701
rect 2217 31649 2233 31701
rect 2233 31649 2285 31701
rect 2285 31649 2301 31701
rect 2301 31649 2353 31701
rect 2353 31649 2369 31701
rect 2369 31649 2421 31701
rect 2421 31649 2437 31701
rect 2437 31649 2489 31701
rect 2489 31649 2505 31701
rect 2505 31649 2557 31701
rect 2557 31649 2573 31701
rect 2573 31649 2625 31701
rect 2625 31649 2641 31701
rect 2641 31649 2663 31701
rect 2127 31637 2663 31649
rect 2127 31585 2149 31637
rect 2149 31585 2165 31637
rect 2165 31585 2217 31637
rect 2217 31585 2233 31637
rect 2233 31585 2285 31637
rect 2285 31585 2301 31637
rect 2301 31585 2353 31637
rect 2353 31585 2369 31637
rect 2369 31585 2421 31637
rect 2421 31585 2437 31637
rect 2437 31585 2489 31637
rect 2489 31585 2505 31637
rect 2505 31585 2557 31637
rect 2557 31585 2573 31637
rect 2573 31585 2625 31637
rect 2625 31585 2641 31637
rect 2641 31585 2663 31637
rect 2127 31573 2663 31585
rect 2127 31562 2149 31573
rect 2149 31562 2165 31573
rect 2165 31562 2217 31573
rect 2217 31562 2233 31573
rect 2233 31562 2285 31573
rect 2285 31562 2301 31573
rect 2301 31562 2353 31573
rect 2353 31562 2369 31573
rect 2369 31562 2421 31573
rect 2421 31562 2437 31573
rect 2437 31562 2489 31573
rect 2489 31562 2505 31573
rect 2505 31562 2557 31573
rect 2557 31562 2573 31573
rect 2573 31562 2625 31573
rect 2625 31562 2641 31573
rect 2641 31562 2663 31573
rect 2127 31521 2149 31537
rect 2149 31521 2165 31537
rect 2165 31521 2183 31537
rect 2207 31521 2217 31537
rect 2217 31521 2233 31537
rect 2233 31521 2263 31537
rect 2287 31521 2301 31537
rect 2301 31521 2343 31537
rect 2367 31521 2369 31537
rect 2369 31521 2421 31537
rect 2421 31521 2423 31537
rect 2447 31521 2489 31537
rect 2489 31521 2503 31537
rect 2527 31521 2557 31537
rect 2557 31521 2573 31537
rect 2573 31521 2583 31537
rect 2607 31521 2625 31537
rect 2625 31521 2641 31537
rect 2641 31521 2663 31537
rect 2127 31509 2183 31521
rect 2207 31509 2263 31521
rect 2287 31509 2343 31521
rect 2367 31509 2423 31521
rect 2447 31509 2503 31521
rect 2527 31509 2583 31521
rect 2607 31509 2663 31521
rect 2127 31481 2149 31509
rect 2149 31481 2165 31509
rect 2165 31481 2183 31509
rect 2207 31481 2217 31509
rect 2217 31481 2233 31509
rect 2233 31481 2263 31509
rect 2287 31481 2301 31509
rect 2301 31481 2343 31509
rect 2367 31481 2369 31509
rect 2369 31481 2421 31509
rect 2421 31481 2423 31509
rect 2447 31481 2489 31509
rect 2489 31481 2503 31509
rect 2527 31481 2557 31509
rect 2557 31481 2573 31509
rect 2573 31481 2583 31509
rect 2607 31481 2625 31509
rect 2625 31481 2641 31509
rect 2641 31481 2663 31509
rect 2127 31445 2183 31456
rect 2207 31445 2263 31456
rect 2287 31445 2343 31456
rect 2367 31445 2423 31456
rect 2447 31445 2503 31456
rect 2527 31445 2583 31456
rect 2607 31445 2663 31456
rect 2127 31400 2149 31445
rect 2149 31400 2165 31445
rect 2165 31400 2183 31445
rect 2207 31400 2217 31445
rect 2217 31400 2233 31445
rect 2233 31400 2263 31445
rect 2287 31400 2301 31445
rect 2301 31400 2343 31445
rect 2367 31400 2369 31445
rect 2369 31400 2421 31445
rect 2421 31400 2423 31445
rect 2447 31400 2489 31445
rect 2489 31400 2503 31445
rect 2527 31400 2557 31445
rect 2557 31400 2573 31445
rect 2573 31400 2583 31445
rect 2607 31400 2625 31445
rect 2625 31400 2641 31445
rect 2641 31400 2663 31445
rect 2127 31329 2149 31375
rect 2149 31329 2165 31375
rect 2165 31329 2183 31375
rect 2207 31329 2217 31375
rect 2217 31329 2233 31375
rect 2233 31329 2263 31375
rect 2287 31329 2301 31375
rect 2301 31329 2343 31375
rect 2367 31329 2369 31375
rect 2369 31329 2421 31375
rect 2421 31329 2423 31375
rect 2447 31329 2489 31375
rect 2489 31329 2503 31375
rect 2527 31329 2557 31375
rect 2557 31329 2573 31375
rect 2573 31329 2583 31375
rect 2607 31329 2625 31375
rect 2625 31329 2641 31375
rect 2641 31329 2663 31375
rect 2127 31319 2183 31329
rect 2207 31319 2263 31329
rect 2287 31319 2343 31329
rect 2367 31319 2423 31329
rect 2447 31319 2503 31329
rect 2527 31319 2583 31329
rect 2607 31319 2663 31329
rect 2127 31265 2149 31294
rect 2149 31265 2165 31294
rect 2165 31265 2183 31294
rect 2207 31265 2217 31294
rect 2217 31265 2233 31294
rect 2233 31265 2263 31294
rect 2287 31265 2301 31294
rect 2301 31265 2343 31294
rect 2367 31265 2369 31294
rect 2369 31265 2421 31294
rect 2421 31265 2423 31294
rect 2447 31265 2489 31294
rect 2489 31265 2503 31294
rect 2527 31265 2557 31294
rect 2557 31265 2573 31294
rect 2573 31265 2583 31294
rect 2607 31265 2625 31294
rect 2625 31265 2641 31294
rect 2641 31265 2663 31294
rect 2127 31253 2183 31265
rect 2207 31253 2263 31265
rect 2287 31253 2343 31265
rect 2367 31253 2423 31265
rect 2447 31253 2503 31265
rect 2527 31253 2583 31265
rect 2607 31253 2663 31265
rect 2127 31238 2149 31253
rect 2149 31238 2165 31253
rect 2165 31238 2183 31253
rect 2207 31238 2217 31253
rect 2217 31238 2233 31253
rect 2233 31238 2263 31253
rect 2287 31238 2301 31253
rect 2301 31238 2343 31253
rect 2367 31238 2369 31253
rect 2369 31238 2421 31253
rect 2421 31238 2423 31253
rect 2447 31238 2489 31253
rect 2489 31238 2503 31253
rect 2527 31238 2557 31253
rect 2557 31238 2573 31253
rect 2573 31238 2583 31253
rect 2607 31238 2625 31253
rect 2625 31238 2641 31253
rect 2641 31238 2663 31253
rect 2127 31201 2149 31213
rect 2149 31201 2165 31213
rect 2165 31201 2183 31213
rect 2207 31201 2217 31213
rect 2217 31201 2233 31213
rect 2233 31201 2263 31213
rect 2287 31201 2301 31213
rect 2301 31201 2343 31213
rect 2367 31201 2369 31213
rect 2369 31201 2421 31213
rect 2421 31201 2423 31213
rect 2447 31201 2489 31213
rect 2489 31201 2503 31213
rect 2527 31201 2557 31213
rect 2557 31201 2573 31213
rect 2573 31201 2583 31213
rect 2607 31201 2625 31213
rect 2625 31201 2641 31213
rect 2641 31201 2663 31213
rect 2127 31189 2183 31201
rect 2207 31189 2263 31201
rect 2287 31189 2343 31201
rect 2367 31189 2423 31201
rect 2447 31189 2503 31201
rect 2527 31189 2583 31201
rect 2607 31189 2663 31201
rect 2127 31157 2149 31189
rect 2149 31157 2165 31189
rect 2165 31157 2183 31189
rect 2207 31157 2217 31189
rect 2217 31157 2233 31189
rect 2233 31157 2263 31189
rect 2287 31157 2301 31189
rect 2301 31157 2343 31189
rect 2367 31157 2369 31189
rect 2369 31157 2421 31189
rect 2421 31157 2423 31189
rect 2447 31157 2489 31189
rect 2489 31157 2503 31189
rect 2527 31157 2557 31189
rect 2557 31157 2573 31189
rect 2573 31157 2583 31189
rect 2607 31157 2625 31189
rect 2625 31157 2641 31189
rect 2641 31157 2663 31189
rect 2127 31125 2183 31132
rect 2207 31125 2263 31132
rect 2287 31125 2343 31132
rect 2367 31125 2423 31132
rect 2447 31125 2503 31132
rect 2527 31125 2583 31132
rect 2607 31125 2663 31132
rect 2127 31076 2149 31125
rect 2149 31076 2165 31125
rect 2165 31076 2183 31125
rect 2207 31076 2217 31125
rect 2217 31076 2233 31125
rect 2233 31076 2263 31125
rect 2287 31076 2301 31125
rect 2301 31076 2343 31125
rect 2367 31076 2369 31125
rect 2369 31076 2421 31125
rect 2421 31076 2423 31125
rect 2447 31076 2489 31125
rect 2489 31076 2503 31125
rect 2527 31076 2557 31125
rect 2557 31076 2573 31125
rect 2573 31076 2583 31125
rect 2607 31076 2625 31125
rect 2625 31076 2641 31125
rect 2641 31076 2663 31125
rect 2127 29820 2149 29869
rect 2149 29820 2165 29869
rect 2165 29820 2217 29869
rect 2217 29820 2233 29869
rect 2233 29820 2285 29869
rect 2285 29820 2301 29869
rect 2301 29820 2353 29869
rect 2353 29820 2369 29869
rect 2369 29820 2421 29869
rect 2421 29820 2437 29869
rect 2437 29820 2489 29869
rect 2489 29820 2505 29869
rect 2505 29820 2557 29869
rect 2557 29820 2573 29869
rect 2573 29820 2625 29869
rect 2625 29820 2641 29869
rect 2641 29820 2663 29869
rect 2127 29808 2663 29820
rect 2127 29756 2149 29808
rect 2149 29756 2165 29808
rect 2165 29756 2217 29808
rect 2217 29756 2233 29808
rect 2233 29756 2285 29808
rect 2285 29756 2301 29808
rect 2301 29756 2353 29808
rect 2353 29756 2369 29808
rect 2369 29756 2421 29808
rect 2421 29756 2437 29808
rect 2437 29756 2489 29808
rect 2489 29756 2505 29808
rect 2505 29756 2557 29808
rect 2557 29756 2573 29808
rect 2573 29756 2625 29808
rect 2625 29756 2641 29808
rect 2641 29756 2663 29808
rect 2127 29744 2663 29756
rect 2127 29692 2149 29744
rect 2149 29692 2165 29744
rect 2165 29692 2217 29744
rect 2217 29692 2233 29744
rect 2233 29692 2285 29744
rect 2285 29692 2301 29744
rect 2301 29692 2353 29744
rect 2353 29692 2369 29744
rect 2369 29692 2421 29744
rect 2421 29692 2437 29744
rect 2437 29692 2489 29744
rect 2489 29692 2505 29744
rect 2505 29692 2557 29744
rect 2557 29692 2573 29744
rect 2573 29692 2625 29744
rect 2625 29692 2641 29744
rect 2641 29692 2663 29744
rect 2127 29680 2663 29692
rect 2127 29628 2149 29680
rect 2149 29628 2165 29680
rect 2165 29628 2217 29680
rect 2217 29628 2233 29680
rect 2233 29628 2285 29680
rect 2285 29628 2301 29680
rect 2301 29628 2353 29680
rect 2353 29628 2369 29680
rect 2369 29628 2421 29680
rect 2421 29628 2437 29680
rect 2437 29628 2489 29680
rect 2489 29628 2505 29680
rect 2505 29628 2557 29680
rect 2557 29628 2573 29680
rect 2573 29628 2625 29680
rect 2625 29628 2641 29680
rect 2641 29628 2663 29680
rect 2127 29616 2663 29628
rect 2127 29564 2149 29616
rect 2149 29564 2165 29616
rect 2165 29564 2217 29616
rect 2217 29564 2233 29616
rect 2233 29564 2285 29616
rect 2285 29564 2301 29616
rect 2301 29564 2353 29616
rect 2353 29564 2369 29616
rect 2369 29564 2421 29616
rect 2421 29564 2437 29616
rect 2437 29564 2489 29616
rect 2489 29564 2505 29616
rect 2505 29564 2557 29616
rect 2557 29564 2573 29616
rect 2573 29564 2625 29616
rect 2625 29564 2641 29616
rect 2641 29564 2663 29616
rect 2127 29552 2663 29564
rect 2127 29500 2149 29552
rect 2149 29500 2165 29552
rect 2165 29500 2217 29552
rect 2217 29500 2233 29552
rect 2233 29500 2285 29552
rect 2285 29500 2301 29552
rect 2301 29500 2353 29552
rect 2353 29500 2369 29552
rect 2369 29500 2421 29552
rect 2421 29500 2437 29552
rect 2437 29500 2489 29552
rect 2489 29500 2505 29552
rect 2505 29500 2557 29552
rect 2557 29500 2573 29552
rect 2573 29500 2625 29552
rect 2625 29500 2641 29552
rect 2641 29500 2663 29552
rect 2127 29488 2663 29500
rect 2127 29436 2149 29488
rect 2149 29436 2165 29488
rect 2165 29436 2217 29488
rect 2217 29436 2233 29488
rect 2233 29436 2285 29488
rect 2285 29436 2301 29488
rect 2301 29436 2353 29488
rect 2353 29436 2369 29488
rect 2369 29436 2421 29488
rect 2421 29436 2437 29488
rect 2437 29436 2489 29488
rect 2489 29436 2505 29488
rect 2505 29436 2557 29488
rect 2557 29436 2573 29488
rect 2573 29436 2625 29488
rect 2625 29436 2641 29488
rect 2641 29436 2663 29488
rect 2127 29424 2663 29436
rect 2127 29413 2149 29424
rect 2149 29413 2165 29424
rect 2165 29413 2217 29424
rect 2217 29413 2233 29424
rect 2233 29413 2285 29424
rect 2285 29413 2301 29424
rect 2301 29413 2353 29424
rect 2353 29413 2369 29424
rect 2369 29413 2421 29424
rect 2421 29413 2437 29424
rect 2437 29413 2489 29424
rect 2489 29413 2505 29424
rect 2505 29413 2557 29424
rect 2557 29413 2573 29424
rect 2573 29413 2625 29424
rect 2625 29413 2641 29424
rect 2641 29413 2663 29424
rect 2127 29372 2149 29388
rect 2149 29372 2165 29388
rect 2165 29372 2183 29388
rect 2207 29372 2217 29388
rect 2217 29372 2233 29388
rect 2233 29372 2263 29388
rect 2287 29372 2301 29388
rect 2301 29372 2343 29388
rect 2367 29372 2369 29388
rect 2369 29372 2421 29388
rect 2421 29372 2423 29388
rect 2447 29372 2489 29388
rect 2489 29372 2503 29388
rect 2527 29372 2557 29388
rect 2557 29372 2573 29388
rect 2573 29372 2583 29388
rect 2607 29372 2625 29388
rect 2625 29372 2641 29388
rect 2641 29372 2663 29388
rect 2127 29360 2183 29372
rect 2207 29360 2263 29372
rect 2287 29360 2343 29372
rect 2367 29360 2423 29372
rect 2447 29360 2503 29372
rect 2527 29360 2583 29372
rect 2607 29360 2663 29372
rect 2127 29332 2149 29360
rect 2149 29332 2165 29360
rect 2165 29332 2183 29360
rect 2207 29332 2217 29360
rect 2217 29332 2233 29360
rect 2233 29332 2263 29360
rect 2287 29332 2301 29360
rect 2301 29332 2343 29360
rect 2367 29332 2369 29360
rect 2369 29332 2421 29360
rect 2421 29332 2423 29360
rect 2447 29332 2489 29360
rect 2489 29332 2503 29360
rect 2527 29332 2557 29360
rect 2557 29332 2573 29360
rect 2573 29332 2583 29360
rect 2607 29332 2625 29360
rect 2625 29332 2641 29360
rect 2641 29332 2663 29360
rect 2127 29296 2183 29307
rect 2207 29296 2263 29307
rect 2287 29296 2343 29307
rect 2367 29296 2423 29307
rect 2447 29296 2503 29307
rect 2527 29296 2583 29307
rect 2607 29296 2663 29307
rect 2127 29251 2149 29296
rect 2149 29251 2165 29296
rect 2165 29251 2183 29296
rect 2207 29251 2217 29296
rect 2217 29251 2233 29296
rect 2233 29251 2263 29296
rect 2287 29251 2301 29296
rect 2301 29251 2343 29296
rect 2367 29251 2369 29296
rect 2369 29251 2421 29296
rect 2421 29251 2423 29296
rect 2447 29251 2489 29296
rect 2489 29251 2503 29296
rect 2527 29251 2557 29296
rect 2557 29251 2573 29296
rect 2573 29251 2583 29296
rect 2607 29251 2625 29296
rect 2625 29251 2641 29296
rect 2641 29251 2663 29296
rect 2127 29180 2149 29226
rect 2149 29180 2165 29226
rect 2165 29180 2183 29226
rect 2207 29180 2217 29226
rect 2217 29180 2233 29226
rect 2233 29180 2263 29226
rect 2287 29180 2301 29226
rect 2301 29180 2343 29226
rect 2367 29180 2369 29226
rect 2369 29180 2421 29226
rect 2421 29180 2423 29226
rect 2447 29180 2489 29226
rect 2489 29180 2503 29226
rect 2527 29180 2557 29226
rect 2557 29180 2573 29226
rect 2573 29180 2583 29226
rect 2607 29180 2625 29226
rect 2625 29180 2641 29226
rect 2641 29180 2663 29226
rect 2127 29170 2183 29180
rect 2207 29170 2263 29180
rect 2287 29170 2343 29180
rect 2367 29170 2423 29180
rect 2447 29170 2503 29180
rect 2527 29170 2583 29180
rect 2607 29170 2663 29180
rect 2127 29116 2149 29145
rect 2149 29116 2165 29145
rect 2165 29116 2183 29145
rect 2207 29116 2217 29145
rect 2217 29116 2233 29145
rect 2233 29116 2263 29145
rect 2287 29116 2301 29145
rect 2301 29116 2343 29145
rect 2367 29116 2369 29145
rect 2369 29116 2421 29145
rect 2421 29116 2423 29145
rect 2447 29116 2489 29145
rect 2489 29116 2503 29145
rect 2527 29116 2557 29145
rect 2557 29116 2573 29145
rect 2573 29116 2583 29145
rect 2607 29116 2625 29145
rect 2625 29116 2641 29145
rect 2641 29116 2663 29145
rect 2127 29104 2183 29116
rect 2207 29104 2263 29116
rect 2287 29104 2343 29116
rect 2367 29104 2423 29116
rect 2447 29104 2503 29116
rect 2527 29104 2583 29116
rect 2607 29104 2663 29116
rect 2127 29089 2149 29104
rect 2149 29089 2165 29104
rect 2165 29089 2183 29104
rect 2207 29089 2217 29104
rect 2217 29089 2233 29104
rect 2233 29089 2263 29104
rect 2287 29089 2301 29104
rect 2301 29089 2343 29104
rect 2367 29089 2369 29104
rect 2369 29089 2421 29104
rect 2421 29089 2423 29104
rect 2447 29089 2489 29104
rect 2489 29089 2503 29104
rect 2527 29089 2557 29104
rect 2557 29089 2573 29104
rect 2573 29089 2583 29104
rect 2607 29089 2625 29104
rect 2625 29089 2641 29104
rect 2641 29089 2663 29104
rect 2127 29052 2149 29064
rect 2149 29052 2165 29064
rect 2165 29052 2183 29064
rect 2207 29052 2217 29064
rect 2217 29052 2233 29064
rect 2233 29052 2263 29064
rect 2287 29052 2301 29064
rect 2301 29052 2343 29064
rect 2367 29052 2369 29064
rect 2369 29052 2421 29064
rect 2421 29052 2423 29064
rect 2447 29052 2489 29064
rect 2489 29052 2503 29064
rect 2527 29052 2557 29064
rect 2557 29052 2573 29064
rect 2573 29052 2583 29064
rect 2607 29052 2625 29064
rect 2625 29052 2641 29064
rect 2641 29052 2663 29064
rect 2127 29040 2183 29052
rect 2207 29040 2263 29052
rect 2287 29040 2343 29052
rect 2367 29040 2423 29052
rect 2447 29040 2503 29052
rect 2527 29040 2583 29052
rect 2607 29040 2663 29052
rect 2127 29008 2149 29040
rect 2149 29008 2165 29040
rect 2165 29008 2183 29040
rect 2207 29008 2217 29040
rect 2217 29008 2233 29040
rect 2233 29008 2263 29040
rect 2287 29008 2301 29040
rect 2301 29008 2343 29040
rect 2367 29008 2369 29040
rect 2369 29008 2421 29040
rect 2421 29008 2423 29040
rect 2447 29008 2489 29040
rect 2489 29008 2503 29040
rect 2527 29008 2557 29040
rect 2557 29008 2573 29040
rect 2573 29008 2583 29040
rect 2607 29008 2625 29040
rect 2625 29008 2641 29040
rect 2641 29008 2663 29040
rect 2127 28976 2183 28983
rect 2207 28976 2263 28983
rect 2287 28976 2343 28983
rect 2367 28976 2423 28983
rect 2447 28976 2503 28983
rect 2527 28976 2583 28983
rect 2607 28976 2663 28983
rect 2127 28927 2149 28976
rect 2149 28927 2165 28976
rect 2165 28927 2183 28976
rect 2207 28927 2217 28976
rect 2217 28927 2233 28976
rect 2233 28927 2263 28976
rect 2287 28927 2301 28976
rect 2301 28927 2343 28976
rect 2367 28927 2369 28976
rect 2369 28927 2421 28976
rect 2421 28927 2423 28976
rect 2447 28927 2489 28976
rect 2489 28927 2503 28976
rect 2527 28927 2557 28976
rect 2557 28927 2573 28976
rect 2573 28927 2583 28976
rect 2607 28927 2625 28976
rect 2625 28927 2641 28976
rect 2641 28927 2663 28976
rect 2127 27813 2149 27862
rect 2149 27813 2165 27862
rect 2165 27813 2217 27862
rect 2217 27813 2233 27862
rect 2233 27813 2285 27862
rect 2285 27813 2301 27862
rect 2301 27813 2353 27862
rect 2353 27813 2369 27862
rect 2369 27813 2421 27862
rect 2421 27813 2437 27862
rect 2437 27813 2489 27862
rect 2489 27813 2505 27862
rect 2505 27813 2557 27862
rect 2557 27813 2573 27862
rect 2573 27813 2625 27862
rect 2625 27813 2641 27862
rect 2641 27813 2663 27862
rect 2127 27801 2663 27813
rect 2127 27749 2149 27801
rect 2149 27749 2165 27801
rect 2165 27749 2217 27801
rect 2217 27749 2233 27801
rect 2233 27749 2285 27801
rect 2285 27749 2301 27801
rect 2301 27749 2353 27801
rect 2353 27749 2369 27801
rect 2369 27749 2421 27801
rect 2421 27749 2437 27801
rect 2437 27749 2489 27801
rect 2489 27749 2505 27801
rect 2505 27749 2557 27801
rect 2557 27749 2573 27801
rect 2573 27749 2625 27801
rect 2625 27749 2641 27801
rect 2641 27749 2663 27801
rect 2127 27737 2663 27749
rect 2127 27685 2149 27737
rect 2149 27685 2165 27737
rect 2165 27685 2217 27737
rect 2217 27685 2233 27737
rect 2233 27685 2285 27737
rect 2285 27685 2301 27737
rect 2301 27685 2353 27737
rect 2353 27685 2369 27737
rect 2369 27685 2421 27737
rect 2421 27685 2437 27737
rect 2437 27685 2489 27737
rect 2489 27685 2505 27737
rect 2505 27685 2557 27737
rect 2557 27685 2573 27737
rect 2573 27685 2625 27737
rect 2625 27685 2641 27737
rect 2641 27685 2663 27737
rect 2127 27673 2663 27685
rect 2127 27621 2149 27673
rect 2149 27621 2165 27673
rect 2165 27621 2217 27673
rect 2217 27621 2233 27673
rect 2233 27621 2285 27673
rect 2285 27621 2301 27673
rect 2301 27621 2353 27673
rect 2353 27621 2369 27673
rect 2369 27621 2421 27673
rect 2421 27621 2437 27673
rect 2437 27621 2489 27673
rect 2489 27621 2505 27673
rect 2505 27621 2557 27673
rect 2557 27621 2573 27673
rect 2573 27621 2625 27673
rect 2625 27621 2641 27673
rect 2641 27621 2663 27673
rect 2127 27609 2663 27621
rect 2127 27557 2149 27609
rect 2149 27557 2165 27609
rect 2165 27557 2217 27609
rect 2217 27557 2233 27609
rect 2233 27557 2285 27609
rect 2285 27557 2301 27609
rect 2301 27557 2353 27609
rect 2353 27557 2369 27609
rect 2369 27557 2421 27609
rect 2421 27557 2437 27609
rect 2437 27557 2489 27609
rect 2489 27557 2505 27609
rect 2505 27557 2557 27609
rect 2557 27557 2573 27609
rect 2573 27557 2625 27609
rect 2625 27557 2641 27609
rect 2641 27557 2663 27609
rect 2127 27545 2663 27557
rect 2127 27493 2149 27545
rect 2149 27493 2165 27545
rect 2165 27493 2217 27545
rect 2217 27493 2233 27545
rect 2233 27493 2285 27545
rect 2285 27493 2301 27545
rect 2301 27493 2353 27545
rect 2353 27493 2369 27545
rect 2369 27493 2421 27545
rect 2421 27493 2437 27545
rect 2437 27493 2489 27545
rect 2489 27493 2505 27545
rect 2505 27493 2557 27545
rect 2557 27493 2573 27545
rect 2573 27493 2625 27545
rect 2625 27493 2641 27545
rect 2641 27493 2663 27545
rect 2127 27481 2663 27493
rect 2127 27429 2149 27481
rect 2149 27429 2165 27481
rect 2165 27429 2217 27481
rect 2217 27429 2233 27481
rect 2233 27429 2285 27481
rect 2285 27429 2301 27481
rect 2301 27429 2353 27481
rect 2353 27429 2369 27481
rect 2369 27429 2421 27481
rect 2421 27429 2437 27481
rect 2437 27429 2489 27481
rect 2489 27429 2505 27481
rect 2505 27429 2557 27481
rect 2557 27429 2573 27481
rect 2573 27429 2625 27481
rect 2625 27429 2641 27481
rect 2641 27429 2663 27481
rect 2127 27417 2663 27429
rect 2127 27406 2149 27417
rect 2149 27406 2165 27417
rect 2165 27406 2217 27417
rect 2217 27406 2233 27417
rect 2233 27406 2285 27417
rect 2285 27406 2301 27417
rect 2301 27406 2353 27417
rect 2353 27406 2369 27417
rect 2369 27406 2421 27417
rect 2421 27406 2437 27417
rect 2437 27406 2489 27417
rect 2489 27406 2505 27417
rect 2505 27406 2557 27417
rect 2557 27406 2573 27417
rect 2573 27406 2625 27417
rect 2625 27406 2641 27417
rect 2641 27406 2663 27417
rect 2127 27365 2149 27381
rect 2149 27365 2165 27381
rect 2165 27365 2183 27381
rect 2207 27365 2217 27381
rect 2217 27365 2233 27381
rect 2233 27365 2263 27381
rect 2287 27365 2301 27381
rect 2301 27365 2343 27381
rect 2367 27365 2369 27381
rect 2369 27365 2421 27381
rect 2421 27365 2423 27381
rect 2447 27365 2489 27381
rect 2489 27365 2503 27381
rect 2527 27365 2557 27381
rect 2557 27365 2573 27381
rect 2573 27365 2583 27381
rect 2607 27365 2625 27381
rect 2625 27365 2641 27381
rect 2641 27365 2663 27381
rect 2127 27353 2183 27365
rect 2207 27353 2263 27365
rect 2287 27353 2343 27365
rect 2367 27353 2423 27365
rect 2447 27353 2503 27365
rect 2527 27353 2583 27365
rect 2607 27353 2663 27365
rect 2127 27325 2149 27353
rect 2149 27325 2165 27353
rect 2165 27325 2183 27353
rect 2207 27325 2217 27353
rect 2217 27325 2233 27353
rect 2233 27325 2263 27353
rect 2287 27325 2301 27353
rect 2301 27325 2343 27353
rect 2367 27325 2369 27353
rect 2369 27325 2421 27353
rect 2421 27325 2423 27353
rect 2447 27325 2489 27353
rect 2489 27325 2503 27353
rect 2527 27325 2557 27353
rect 2557 27325 2573 27353
rect 2573 27325 2583 27353
rect 2607 27325 2625 27353
rect 2625 27325 2641 27353
rect 2641 27325 2663 27353
rect 2127 27289 2183 27300
rect 2207 27289 2263 27300
rect 2287 27289 2343 27300
rect 2367 27289 2423 27300
rect 2447 27289 2503 27300
rect 2527 27289 2583 27300
rect 2607 27289 2663 27300
rect 2127 27244 2149 27289
rect 2149 27244 2165 27289
rect 2165 27244 2183 27289
rect 2207 27244 2217 27289
rect 2217 27244 2233 27289
rect 2233 27244 2263 27289
rect 2287 27244 2301 27289
rect 2301 27244 2343 27289
rect 2367 27244 2369 27289
rect 2369 27244 2421 27289
rect 2421 27244 2423 27289
rect 2447 27244 2489 27289
rect 2489 27244 2503 27289
rect 2527 27244 2557 27289
rect 2557 27244 2573 27289
rect 2573 27244 2583 27289
rect 2607 27244 2625 27289
rect 2625 27244 2641 27289
rect 2641 27244 2663 27289
rect 2127 27173 2149 27219
rect 2149 27173 2165 27219
rect 2165 27173 2183 27219
rect 2207 27173 2217 27219
rect 2217 27173 2233 27219
rect 2233 27173 2263 27219
rect 2287 27173 2301 27219
rect 2301 27173 2343 27219
rect 2367 27173 2369 27219
rect 2369 27173 2421 27219
rect 2421 27173 2423 27219
rect 2447 27173 2489 27219
rect 2489 27173 2503 27219
rect 2527 27173 2557 27219
rect 2557 27173 2573 27219
rect 2573 27173 2583 27219
rect 2607 27173 2625 27219
rect 2625 27173 2641 27219
rect 2641 27173 2663 27219
rect 2127 27163 2183 27173
rect 2207 27163 2263 27173
rect 2287 27163 2343 27173
rect 2367 27163 2423 27173
rect 2447 27163 2503 27173
rect 2527 27163 2583 27173
rect 2607 27163 2663 27173
rect 2127 27109 2149 27138
rect 2149 27109 2165 27138
rect 2165 27109 2183 27138
rect 2207 27109 2217 27138
rect 2217 27109 2233 27138
rect 2233 27109 2263 27138
rect 2287 27109 2301 27138
rect 2301 27109 2343 27138
rect 2367 27109 2369 27138
rect 2369 27109 2421 27138
rect 2421 27109 2423 27138
rect 2447 27109 2489 27138
rect 2489 27109 2503 27138
rect 2527 27109 2557 27138
rect 2557 27109 2573 27138
rect 2573 27109 2583 27138
rect 2607 27109 2625 27138
rect 2625 27109 2641 27138
rect 2641 27109 2663 27138
rect 2127 27097 2183 27109
rect 2207 27097 2263 27109
rect 2287 27097 2343 27109
rect 2367 27097 2423 27109
rect 2447 27097 2503 27109
rect 2527 27097 2583 27109
rect 2607 27097 2663 27109
rect 2127 27082 2149 27097
rect 2149 27082 2165 27097
rect 2165 27082 2183 27097
rect 2207 27082 2217 27097
rect 2217 27082 2233 27097
rect 2233 27082 2263 27097
rect 2287 27082 2301 27097
rect 2301 27082 2343 27097
rect 2367 27082 2369 27097
rect 2369 27082 2421 27097
rect 2421 27082 2423 27097
rect 2447 27082 2489 27097
rect 2489 27082 2503 27097
rect 2527 27082 2557 27097
rect 2557 27082 2573 27097
rect 2573 27082 2583 27097
rect 2607 27082 2625 27097
rect 2625 27082 2641 27097
rect 2641 27082 2663 27097
rect 2127 27045 2149 27057
rect 2149 27045 2165 27057
rect 2165 27045 2183 27057
rect 2207 27045 2217 27057
rect 2217 27045 2233 27057
rect 2233 27045 2263 27057
rect 2287 27045 2301 27057
rect 2301 27045 2343 27057
rect 2367 27045 2369 27057
rect 2369 27045 2421 27057
rect 2421 27045 2423 27057
rect 2447 27045 2489 27057
rect 2489 27045 2503 27057
rect 2527 27045 2557 27057
rect 2557 27045 2573 27057
rect 2573 27045 2583 27057
rect 2607 27045 2625 27057
rect 2625 27045 2641 27057
rect 2641 27045 2663 27057
rect 2127 27033 2183 27045
rect 2207 27033 2263 27045
rect 2287 27033 2343 27045
rect 2367 27033 2423 27045
rect 2447 27033 2503 27045
rect 2527 27033 2583 27045
rect 2607 27033 2663 27045
rect 2127 27001 2149 27033
rect 2149 27001 2165 27033
rect 2165 27001 2183 27033
rect 2207 27001 2217 27033
rect 2217 27001 2233 27033
rect 2233 27001 2263 27033
rect 2287 27001 2301 27033
rect 2301 27001 2343 27033
rect 2367 27001 2369 27033
rect 2369 27001 2421 27033
rect 2421 27001 2423 27033
rect 2447 27001 2489 27033
rect 2489 27001 2503 27033
rect 2527 27001 2557 27033
rect 2557 27001 2573 27033
rect 2573 27001 2583 27033
rect 2607 27001 2625 27033
rect 2625 27001 2641 27033
rect 2641 27001 2663 27033
rect 2127 26969 2183 26976
rect 2207 26969 2263 26976
rect 2287 26969 2343 26976
rect 2367 26969 2423 26976
rect 2447 26969 2503 26976
rect 2527 26969 2583 26976
rect 2607 26969 2663 26976
rect 2127 26920 2149 26969
rect 2149 26920 2165 26969
rect 2165 26920 2183 26969
rect 2207 26920 2217 26969
rect 2217 26920 2233 26969
rect 2233 26920 2263 26969
rect 2287 26920 2301 26969
rect 2301 26920 2343 26969
rect 2367 26920 2369 26969
rect 2369 26920 2421 26969
rect 2421 26920 2423 26969
rect 2447 26920 2489 26969
rect 2489 26920 2503 26969
rect 2527 26920 2557 26969
rect 2557 26920 2573 26969
rect 2573 26920 2583 26969
rect 2607 26920 2625 26969
rect 2625 26920 2641 26969
rect 2641 26920 2663 26969
rect 2127 25627 2149 25676
rect 2149 25627 2165 25676
rect 2165 25627 2217 25676
rect 2217 25627 2233 25676
rect 2233 25627 2285 25676
rect 2285 25627 2301 25676
rect 2301 25627 2353 25676
rect 2353 25627 2369 25676
rect 2369 25627 2421 25676
rect 2421 25627 2437 25676
rect 2437 25627 2489 25676
rect 2489 25627 2505 25676
rect 2505 25627 2557 25676
rect 2557 25627 2573 25676
rect 2573 25627 2625 25676
rect 2625 25627 2641 25676
rect 2641 25627 2663 25676
rect 2127 25615 2663 25627
rect 2127 25563 2149 25615
rect 2149 25563 2165 25615
rect 2165 25563 2217 25615
rect 2217 25563 2233 25615
rect 2233 25563 2285 25615
rect 2285 25563 2301 25615
rect 2301 25563 2353 25615
rect 2353 25563 2369 25615
rect 2369 25563 2421 25615
rect 2421 25563 2437 25615
rect 2437 25563 2489 25615
rect 2489 25563 2505 25615
rect 2505 25563 2557 25615
rect 2557 25563 2573 25615
rect 2573 25563 2625 25615
rect 2625 25563 2641 25615
rect 2641 25563 2663 25615
rect 2127 25551 2663 25563
rect 2127 25499 2149 25551
rect 2149 25499 2165 25551
rect 2165 25499 2217 25551
rect 2217 25499 2233 25551
rect 2233 25499 2285 25551
rect 2285 25499 2301 25551
rect 2301 25499 2353 25551
rect 2353 25499 2369 25551
rect 2369 25499 2421 25551
rect 2421 25499 2437 25551
rect 2437 25499 2489 25551
rect 2489 25499 2505 25551
rect 2505 25499 2557 25551
rect 2557 25499 2573 25551
rect 2573 25499 2625 25551
rect 2625 25499 2641 25551
rect 2641 25499 2663 25551
rect 2127 25487 2663 25499
rect 2127 25435 2149 25487
rect 2149 25435 2165 25487
rect 2165 25435 2217 25487
rect 2217 25435 2233 25487
rect 2233 25435 2285 25487
rect 2285 25435 2301 25487
rect 2301 25435 2353 25487
rect 2353 25435 2369 25487
rect 2369 25435 2421 25487
rect 2421 25435 2437 25487
rect 2437 25435 2489 25487
rect 2489 25435 2505 25487
rect 2505 25435 2557 25487
rect 2557 25435 2573 25487
rect 2573 25435 2625 25487
rect 2625 25435 2641 25487
rect 2641 25435 2663 25487
rect 2127 25423 2663 25435
rect 2127 25371 2149 25423
rect 2149 25371 2165 25423
rect 2165 25371 2217 25423
rect 2217 25371 2233 25423
rect 2233 25371 2285 25423
rect 2285 25371 2301 25423
rect 2301 25371 2353 25423
rect 2353 25371 2369 25423
rect 2369 25371 2421 25423
rect 2421 25371 2437 25423
rect 2437 25371 2489 25423
rect 2489 25371 2505 25423
rect 2505 25371 2557 25423
rect 2557 25371 2573 25423
rect 2573 25371 2625 25423
rect 2625 25371 2641 25423
rect 2641 25371 2663 25423
rect 2127 25359 2663 25371
rect 2127 25307 2149 25359
rect 2149 25307 2165 25359
rect 2165 25307 2217 25359
rect 2217 25307 2233 25359
rect 2233 25307 2285 25359
rect 2285 25307 2301 25359
rect 2301 25307 2353 25359
rect 2353 25307 2369 25359
rect 2369 25307 2421 25359
rect 2421 25307 2437 25359
rect 2437 25307 2489 25359
rect 2489 25307 2505 25359
rect 2505 25307 2557 25359
rect 2557 25307 2573 25359
rect 2573 25307 2625 25359
rect 2625 25307 2641 25359
rect 2641 25307 2663 25359
rect 2127 25295 2663 25307
rect 2127 25243 2149 25295
rect 2149 25243 2165 25295
rect 2165 25243 2217 25295
rect 2217 25243 2233 25295
rect 2233 25243 2285 25295
rect 2285 25243 2301 25295
rect 2301 25243 2353 25295
rect 2353 25243 2369 25295
rect 2369 25243 2421 25295
rect 2421 25243 2437 25295
rect 2437 25243 2489 25295
rect 2489 25243 2505 25295
rect 2505 25243 2557 25295
rect 2557 25243 2573 25295
rect 2573 25243 2625 25295
rect 2625 25243 2641 25295
rect 2641 25243 2663 25295
rect 2127 25231 2663 25243
rect 2127 25220 2149 25231
rect 2149 25220 2165 25231
rect 2165 25220 2217 25231
rect 2217 25220 2233 25231
rect 2233 25220 2285 25231
rect 2285 25220 2301 25231
rect 2301 25220 2353 25231
rect 2353 25220 2369 25231
rect 2369 25220 2421 25231
rect 2421 25220 2437 25231
rect 2437 25220 2489 25231
rect 2489 25220 2505 25231
rect 2505 25220 2557 25231
rect 2557 25220 2573 25231
rect 2573 25220 2625 25231
rect 2625 25220 2641 25231
rect 2641 25220 2663 25231
rect 2127 25179 2149 25195
rect 2149 25179 2165 25195
rect 2165 25179 2183 25195
rect 2207 25179 2217 25195
rect 2217 25179 2233 25195
rect 2233 25179 2263 25195
rect 2287 25179 2301 25195
rect 2301 25179 2343 25195
rect 2367 25179 2369 25195
rect 2369 25179 2421 25195
rect 2421 25179 2423 25195
rect 2447 25179 2489 25195
rect 2489 25179 2503 25195
rect 2527 25179 2557 25195
rect 2557 25179 2573 25195
rect 2573 25179 2583 25195
rect 2607 25179 2625 25195
rect 2625 25179 2641 25195
rect 2641 25179 2663 25195
rect 2127 25167 2183 25179
rect 2207 25167 2263 25179
rect 2287 25167 2343 25179
rect 2367 25167 2423 25179
rect 2447 25167 2503 25179
rect 2527 25167 2583 25179
rect 2607 25167 2663 25179
rect 2127 25139 2149 25167
rect 2149 25139 2165 25167
rect 2165 25139 2183 25167
rect 2207 25139 2217 25167
rect 2217 25139 2233 25167
rect 2233 25139 2263 25167
rect 2287 25139 2301 25167
rect 2301 25139 2343 25167
rect 2367 25139 2369 25167
rect 2369 25139 2421 25167
rect 2421 25139 2423 25167
rect 2447 25139 2489 25167
rect 2489 25139 2503 25167
rect 2527 25139 2557 25167
rect 2557 25139 2573 25167
rect 2573 25139 2583 25167
rect 2607 25139 2625 25167
rect 2625 25139 2641 25167
rect 2641 25139 2663 25167
rect 2127 25103 2183 25114
rect 2207 25103 2263 25114
rect 2287 25103 2343 25114
rect 2367 25103 2423 25114
rect 2447 25103 2503 25114
rect 2527 25103 2583 25114
rect 2607 25103 2663 25114
rect 2127 25058 2149 25103
rect 2149 25058 2165 25103
rect 2165 25058 2183 25103
rect 2207 25058 2217 25103
rect 2217 25058 2233 25103
rect 2233 25058 2263 25103
rect 2287 25058 2301 25103
rect 2301 25058 2343 25103
rect 2367 25058 2369 25103
rect 2369 25058 2421 25103
rect 2421 25058 2423 25103
rect 2447 25058 2489 25103
rect 2489 25058 2503 25103
rect 2527 25058 2557 25103
rect 2557 25058 2573 25103
rect 2573 25058 2583 25103
rect 2607 25058 2625 25103
rect 2625 25058 2641 25103
rect 2641 25058 2663 25103
rect 2127 24987 2149 25033
rect 2149 24987 2165 25033
rect 2165 24987 2183 25033
rect 2207 24987 2217 25033
rect 2217 24987 2233 25033
rect 2233 24987 2263 25033
rect 2287 24987 2301 25033
rect 2301 24987 2343 25033
rect 2367 24987 2369 25033
rect 2369 24987 2421 25033
rect 2421 24987 2423 25033
rect 2447 24987 2489 25033
rect 2489 24987 2503 25033
rect 2527 24987 2557 25033
rect 2557 24987 2573 25033
rect 2573 24987 2583 25033
rect 2607 24987 2625 25033
rect 2625 24987 2641 25033
rect 2641 24987 2663 25033
rect 2127 24977 2183 24987
rect 2207 24977 2263 24987
rect 2287 24977 2343 24987
rect 2367 24977 2423 24987
rect 2447 24977 2503 24987
rect 2527 24977 2583 24987
rect 2607 24977 2663 24987
rect 2127 24923 2149 24952
rect 2149 24923 2165 24952
rect 2165 24923 2183 24952
rect 2207 24923 2217 24952
rect 2217 24923 2233 24952
rect 2233 24923 2263 24952
rect 2287 24923 2301 24952
rect 2301 24923 2343 24952
rect 2367 24923 2369 24952
rect 2369 24923 2421 24952
rect 2421 24923 2423 24952
rect 2447 24923 2489 24952
rect 2489 24923 2503 24952
rect 2527 24923 2557 24952
rect 2557 24923 2573 24952
rect 2573 24923 2583 24952
rect 2607 24923 2625 24952
rect 2625 24923 2641 24952
rect 2641 24923 2663 24952
rect 2127 24911 2183 24923
rect 2207 24911 2263 24923
rect 2287 24911 2343 24923
rect 2367 24911 2423 24923
rect 2447 24911 2503 24923
rect 2527 24911 2583 24923
rect 2607 24911 2663 24923
rect 2127 24896 2149 24911
rect 2149 24896 2165 24911
rect 2165 24896 2183 24911
rect 2207 24896 2217 24911
rect 2217 24896 2233 24911
rect 2233 24896 2263 24911
rect 2287 24896 2301 24911
rect 2301 24896 2343 24911
rect 2367 24896 2369 24911
rect 2369 24896 2421 24911
rect 2421 24896 2423 24911
rect 2447 24896 2489 24911
rect 2489 24896 2503 24911
rect 2527 24896 2557 24911
rect 2557 24896 2573 24911
rect 2573 24896 2583 24911
rect 2607 24896 2625 24911
rect 2625 24896 2641 24911
rect 2641 24896 2663 24911
rect 2127 24859 2149 24871
rect 2149 24859 2165 24871
rect 2165 24859 2183 24871
rect 2207 24859 2217 24871
rect 2217 24859 2233 24871
rect 2233 24859 2263 24871
rect 2287 24859 2301 24871
rect 2301 24859 2343 24871
rect 2367 24859 2369 24871
rect 2369 24859 2421 24871
rect 2421 24859 2423 24871
rect 2447 24859 2489 24871
rect 2489 24859 2503 24871
rect 2527 24859 2557 24871
rect 2557 24859 2573 24871
rect 2573 24859 2583 24871
rect 2607 24859 2625 24871
rect 2625 24859 2641 24871
rect 2641 24859 2663 24871
rect 2127 24847 2183 24859
rect 2207 24847 2263 24859
rect 2287 24847 2343 24859
rect 2367 24847 2423 24859
rect 2447 24847 2503 24859
rect 2527 24847 2583 24859
rect 2607 24847 2663 24859
rect 2127 24815 2149 24847
rect 2149 24815 2165 24847
rect 2165 24815 2183 24847
rect 2207 24815 2217 24847
rect 2217 24815 2233 24847
rect 2233 24815 2263 24847
rect 2287 24815 2301 24847
rect 2301 24815 2343 24847
rect 2367 24815 2369 24847
rect 2369 24815 2421 24847
rect 2421 24815 2423 24847
rect 2447 24815 2489 24847
rect 2489 24815 2503 24847
rect 2527 24815 2557 24847
rect 2557 24815 2573 24847
rect 2573 24815 2583 24847
rect 2607 24815 2625 24847
rect 2625 24815 2641 24847
rect 2641 24815 2663 24847
rect 2127 24783 2183 24790
rect 2207 24783 2263 24790
rect 2287 24783 2343 24790
rect 2367 24783 2423 24790
rect 2447 24783 2503 24790
rect 2527 24783 2583 24790
rect 2607 24783 2663 24790
rect 2127 24734 2149 24783
rect 2149 24734 2165 24783
rect 2165 24734 2183 24783
rect 2207 24734 2217 24783
rect 2217 24734 2233 24783
rect 2233 24734 2263 24783
rect 2287 24734 2301 24783
rect 2301 24734 2343 24783
rect 2367 24734 2369 24783
rect 2369 24734 2421 24783
rect 2421 24734 2423 24783
rect 2447 24734 2489 24783
rect 2489 24734 2503 24783
rect 2527 24734 2557 24783
rect 2557 24734 2573 24783
rect 2573 24734 2583 24783
rect 2607 24734 2625 24783
rect 2625 24734 2641 24783
rect 2641 24734 2663 24783
rect 2127 23479 2149 23528
rect 2149 23479 2165 23528
rect 2165 23479 2217 23528
rect 2217 23479 2233 23528
rect 2233 23479 2285 23528
rect 2285 23479 2301 23528
rect 2301 23479 2353 23528
rect 2353 23479 2369 23528
rect 2369 23479 2421 23528
rect 2421 23479 2437 23528
rect 2437 23479 2489 23528
rect 2489 23479 2505 23528
rect 2505 23479 2557 23528
rect 2557 23479 2573 23528
rect 2573 23479 2625 23528
rect 2625 23479 2641 23528
rect 2641 23479 2663 23528
rect 2127 23467 2663 23479
rect 2127 23415 2149 23467
rect 2149 23415 2165 23467
rect 2165 23415 2217 23467
rect 2217 23415 2233 23467
rect 2233 23415 2285 23467
rect 2285 23415 2301 23467
rect 2301 23415 2353 23467
rect 2353 23415 2369 23467
rect 2369 23415 2421 23467
rect 2421 23415 2437 23467
rect 2437 23415 2489 23467
rect 2489 23415 2505 23467
rect 2505 23415 2557 23467
rect 2557 23415 2573 23467
rect 2573 23415 2625 23467
rect 2625 23415 2641 23467
rect 2641 23415 2663 23467
rect 2127 23403 2663 23415
rect 2127 23351 2149 23403
rect 2149 23351 2165 23403
rect 2165 23351 2217 23403
rect 2217 23351 2233 23403
rect 2233 23351 2285 23403
rect 2285 23351 2301 23403
rect 2301 23351 2353 23403
rect 2353 23351 2369 23403
rect 2369 23351 2421 23403
rect 2421 23351 2437 23403
rect 2437 23351 2489 23403
rect 2489 23351 2505 23403
rect 2505 23351 2557 23403
rect 2557 23351 2573 23403
rect 2573 23351 2625 23403
rect 2625 23351 2641 23403
rect 2641 23351 2663 23403
rect 2127 23339 2663 23351
rect 2127 23287 2149 23339
rect 2149 23287 2165 23339
rect 2165 23287 2217 23339
rect 2217 23287 2233 23339
rect 2233 23287 2285 23339
rect 2285 23287 2301 23339
rect 2301 23287 2353 23339
rect 2353 23287 2369 23339
rect 2369 23287 2421 23339
rect 2421 23287 2437 23339
rect 2437 23287 2489 23339
rect 2489 23287 2505 23339
rect 2505 23287 2557 23339
rect 2557 23287 2573 23339
rect 2573 23287 2625 23339
rect 2625 23287 2641 23339
rect 2641 23287 2663 23339
rect 2127 23275 2663 23287
rect 2127 23223 2149 23275
rect 2149 23223 2165 23275
rect 2165 23223 2217 23275
rect 2217 23223 2233 23275
rect 2233 23223 2285 23275
rect 2285 23223 2301 23275
rect 2301 23223 2353 23275
rect 2353 23223 2369 23275
rect 2369 23223 2421 23275
rect 2421 23223 2437 23275
rect 2437 23223 2489 23275
rect 2489 23223 2505 23275
rect 2505 23223 2557 23275
rect 2557 23223 2573 23275
rect 2573 23223 2625 23275
rect 2625 23223 2641 23275
rect 2641 23223 2663 23275
rect 2127 23211 2663 23223
rect 2127 23159 2149 23211
rect 2149 23159 2165 23211
rect 2165 23159 2217 23211
rect 2217 23159 2233 23211
rect 2233 23159 2285 23211
rect 2285 23159 2301 23211
rect 2301 23159 2353 23211
rect 2353 23159 2369 23211
rect 2369 23159 2421 23211
rect 2421 23159 2437 23211
rect 2437 23159 2489 23211
rect 2489 23159 2505 23211
rect 2505 23159 2557 23211
rect 2557 23159 2573 23211
rect 2573 23159 2625 23211
rect 2625 23159 2641 23211
rect 2641 23159 2663 23211
rect 2127 23147 2663 23159
rect 2127 23095 2149 23147
rect 2149 23095 2165 23147
rect 2165 23095 2217 23147
rect 2217 23095 2233 23147
rect 2233 23095 2285 23147
rect 2285 23095 2301 23147
rect 2301 23095 2353 23147
rect 2353 23095 2369 23147
rect 2369 23095 2421 23147
rect 2421 23095 2437 23147
rect 2437 23095 2489 23147
rect 2489 23095 2505 23147
rect 2505 23095 2557 23147
rect 2557 23095 2573 23147
rect 2573 23095 2625 23147
rect 2625 23095 2641 23147
rect 2641 23095 2663 23147
rect 2127 23083 2663 23095
rect 2127 23072 2149 23083
rect 2149 23072 2165 23083
rect 2165 23072 2217 23083
rect 2217 23072 2233 23083
rect 2233 23072 2285 23083
rect 2285 23072 2301 23083
rect 2301 23072 2353 23083
rect 2353 23072 2369 23083
rect 2369 23072 2421 23083
rect 2421 23072 2437 23083
rect 2437 23072 2489 23083
rect 2489 23072 2505 23083
rect 2505 23072 2557 23083
rect 2557 23072 2573 23083
rect 2573 23072 2625 23083
rect 2625 23072 2641 23083
rect 2641 23072 2663 23083
rect 2127 23031 2149 23047
rect 2149 23031 2165 23047
rect 2165 23031 2183 23047
rect 2207 23031 2217 23047
rect 2217 23031 2233 23047
rect 2233 23031 2263 23047
rect 2287 23031 2301 23047
rect 2301 23031 2343 23047
rect 2367 23031 2369 23047
rect 2369 23031 2421 23047
rect 2421 23031 2423 23047
rect 2447 23031 2489 23047
rect 2489 23031 2503 23047
rect 2527 23031 2557 23047
rect 2557 23031 2573 23047
rect 2573 23031 2583 23047
rect 2607 23031 2625 23047
rect 2625 23031 2641 23047
rect 2641 23031 2663 23047
rect 2127 23019 2183 23031
rect 2207 23019 2263 23031
rect 2287 23019 2343 23031
rect 2367 23019 2423 23031
rect 2447 23019 2503 23031
rect 2527 23019 2583 23031
rect 2607 23019 2663 23031
rect 2127 22991 2149 23019
rect 2149 22991 2165 23019
rect 2165 22991 2183 23019
rect 2207 22991 2217 23019
rect 2217 22991 2233 23019
rect 2233 22991 2263 23019
rect 2287 22991 2301 23019
rect 2301 22991 2343 23019
rect 2367 22991 2369 23019
rect 2369 22991 2421 23019
rect 2421 22991 2423 23019
rect 2447 22991 2489 23019
rect 2489 22991 2503 23019
rect 2527 22991 2557 23019
rect 2557 22991 2573 23019
rect 2573 22991 2583 23019
rect 2607 22991 2625 23019
rect 2625 22991 2641 23019
rect 2641 22991 2663 23019
rect 2127 22955 2183 22966
rect 2207 22955 2263 22966
rect 2287 22955 2343 22966
rect 2367 22955 2423 22966
rect 2447 22955 2503 22966
rect 2527 22955 2583 22966
rect 2607 22955 2663 22966
rect 2127 22910 2149 22955
rect 2149 22910 2165 22955
rect 2165 22910 2183 22955
rect 2207 22910 2217 22955
rect 2217 22910 2233 22955
rect 2233 22910 2263 22955
rect 2287 22910 2301 22955
rect 2301 22910 2343 22955
rect 2367 22910 2369 22955
rect 2369 22910 2421 22955
rect 2421 22910 2423 22955
rect 2447 22910 2489 22955
rect 2489 22910 2503 22955
rect 2527 22910 2557 22955
rect 2557 22910 2573 22955
rect 2573 22910 2583 22955
rect 2607 22910 2625 22955
rect 2625 22910 2641 22955
rect 2641 22910 2663 22955
rect 2127 22839 2149 22885
rect 2149 22839 2165 22885
rect 2165 22839 2183 22885
rect 2207 22839 2217 22885
rect 2217 22839 2233 22885
rect 2233 22839 2263 22885
rect 2287 22839 2301 22885
rect 2301 22839 2343 22885
rect 2367 22839 2369 22885
rect 2369 22839 2421 22885
rect 2421 22839 2423 22885
rect 2447 22839 2489 22885
rect 2489 22839 2503 22885
rect 2527 22839 2557 22885
rect 2557 22839 2573 22885
rect 2573 22839 2583 22885
rect 2607 22839 2625 22885
rect 2625 22839 2641 22885
rect 2641 22839 2663 22885
rect 2127 22829 2183 22839
rect 2207 22829 2263 22839
rect 2287 22829 2343 22839
rect 2367 22829 2423 22839
rect 2447 22829 2503 22839
rect 2527 22829 2583 22839
rect 2607 22829 2663 22839
rect 2127 22775 2149 22804
rect 2149 22775 2165 22804
rect 2165 22775 2183 22804
rect 2207 22775 2217 22804
rect 2217 22775 2233 22804
rect 2233 22775 2263 22804
rect 2287 22775 2301 22804
rect 2301 22775 2343 22804
rect 2367 22775 2369 22804
rect 2369 22775 2421 22804
rect 2421 22775 2423 22804
rect 2447 22775 2489 22804
rect 2489 22775 2503 22804
rect 2527 22775 2557 22804
rect 2557 22775 2573 22804
rect 2573 22775 2583 22804
rect 2607 22775 2625 22804
rect 2625 22775 2641 22804
rect 2641 22775 2663 22804
rect 2127 22763 2183 22775
rect 2207 22763 2263 22775
rect 2287 22763 2343 22775
rect 2367 22763 2423 22775
rect 2447 22763 2503 22775
rect 2527 22763 2583 22775
rect 2607 22763 2663 22775
rect 2127 22748 2149 22763
rect 2149 22748 2165 22763
rect 2165 22748 2183 22763
rect 2207 22748 2217 22763
rect 2217 22748 2233 22763
rect 2233 22748 2263 22763
rect 2287 22748 2301 22763
rect 2301 22748 2343 22763
rect 2367 22748 2369 22763
rect 2369 22748 2421 22763
rect 2421 22748 2423 22763
rect 2447 22748 2489 22763
rect 2489 22748 2503 22763
rect 2527 22748 2557 22763
rect 2557 22748 2573 22763
rect 2573 22748 2583 22763
rect 2607 22748 2625 22763
rect 2625 22748 2641 22763
rect 2641 22748 2663 22763
rect 2127 22711 2149 22723
rect 2149 22711 2165 22723
rect 2165 22711 2183 22723
rect 2207 22711 2217 22723
rect 2217 22711 2233 22723
rect 2233 22711 2263 22723
rect 2287 22711 2301 22723
rect 2301 22711 2343 22723
rect 2367 22711 2369 22723
rect 2369 22711 2421 22723
rect 2421 22711 2423 22723
rect 2447 22711 2489 22723
rect 2489 22711 2503 22723
rect 2527 22711 2557 22723
rect 2557 22711 2573 22723
rect 2573 22711 2583 22723
rect 2607 22711 2625 22723
rect 2625 22711 2641 22723
rect 2641 22711 2663 22723
rect 2127 22699 2183 22711
rect 2207 22699 2263 22711
rect 2287 22699 2343 22711
rect 2367 22699 2423 22711
rect 2447 22699 2503 22711
rect 2527 22699 2583 22711
rect 2607 22699 2663 22711
rect 2127 22667 2149 22699
rect 2149 22667 2165 22699
rect 2165 22667 2183 22699
rect 2207 22667 2217 22699
rect 2217 22667 2233 22699
rect 2233 22667 2263 22699
rect 2287 22667 2301 22699
rect 2301 22667 2343 22699
rect 2367 22667 2369 22699
rect 2369 22667 2421 22699
rect 2421 22667 2423 22699
rect 2447 22667 2489 22699
rect 2489 22667 2503 22699
rect 2527 22667 2557 22699
rect 2557 22667 2573 22699
rect 2573 22667 2583 22699
rect 2607 22667 2625 22699
rect 2625 22667 2641 22699
rect 2641 22667 2663 22699
rect 2127 22635 2183 22642
rect 2207 22635 2263 22642
rect 2287 22635 2343 22642
rect 2367 22635 2423 22642
rect 2447 22635 2503 22642
rect 2527 22635 2583 22642
rect 2607 22635 2663 22642
rect 2127 22586 2149 22635
rect 2149 22586 2165 22635
rect 2165 22586 2183 22635
rect 2207 22586 2217 22635
rect 2217 22586 2233 22635
rect 2233 22586 2263 22635
rect 2287 22586 2301 22635
rect 2301 22586 2343 22635
rect 2367 22586 2369 22635
rect 2369 22586 2421 22635
rect 2421 22586 2423 22635
rect 2447 22586 2489 22635
rect 2489 22586 2503 22635
rect 2527 22586 2557 22635
rect 2557 22586 2573 22635
rect 2573 22586 2583 22635
rect 2607 22586 2625 22635
rect 2625 22586 2641 22635
rect 2641 22586 2663 22635
rect 2127 21309 2149 21358
rect 2149 21309 2165 21358
rect 2165 21309 2217 21358
rect 2217 21309 2233 21358
rect 2233 21309 2285 21358
rect 2285 21309 2301 21358
rect 2301 21309 2353 21358
rect 2353 21309 2369 21358
rect 2369 21309 2421 21358
rect 2421 21309 2437 21358
rect 2437 21309 2489 21358
rect 2489 21309 2505 21358
rect 2505 21309 2557 21358
rect 2557 21309 2573 21358
rect 2573 21309 2625 21358
rect 2625 21309 2641 21358
rect 2641 21309 2663 21358
rect 2127 21297 2663 21309
rect 2127 21245 2149 21297
rect 2149 21245 2165 21297
rect 2165 21245 2217 21297
rect 2217 21245 2233 21297
rect 2233 21245 2285 21297
rect 2285 21245 2301 21297
rect 2301 21245 2353 21297
rect 2353 21245 2369 21297
rect 2369 21245 2421 21297
rect 2421 21245 2437 21297
rect 2437 21245 2489 21297
rect 2489 21245 2505 21297
rect 2505 21245 2557 21297
rect 2557 21245 2573 21297
rect 2573 21245 2625 21297
rect 2625 21245 2641 21297
rect 2641 21245 2663 21297
rect 2127 21233 2663 21245
rect 2127 21181 2149 21233
rect 2149 21181 2165 21233
rect 2165 21181 2217 21233
rect 2217 21181 2233 21233
rect 2233 21181 2285 21233
rect 2285 21181 2301 21233
rect 2301 21181 2353 21233
rect 2353 21181 2369 21233
rect 2369 21181 2421 21233
rect 2421 21181 2437 21233
rect 2437 21181 2489 21233
rect 2489 21181 2505 21233
rect 2505 21181 2557 21233
rect 2557 21181 2573 21233
rect 2573 21181 2625 21233
rect 2625 21181 2641 21233
rect 2641 21181 2663 21233
rect 2127 21169 2663 21181
rect 2127 21117 2149 21169
rect 2149 21117 2165 21169
rect 2165 21117 2217 21169
rect 2217 21117 2233 21169
rect 2233 21117 2285 21169
rect 2285 21117 2301 21169
rect 2301 21117 2353 21169
rect 2353 21117 2369 21169
rect 2369 21117 2421 21169
rect 2421 21117 2437 21169
rect 2437 21117 2489 21169
rect 2489 21117 2505 21169
rect 2505 21117 2557 21169
rect 2557 21117 2573 21169
rect 2573 21117 2625 21169
rect 2625 21117 2641 21169
rect 2641 21117 2663 21169
rect 2127 21105 2663 21117
rect 2127 21053 2149 21105
rect 2149 21053 2165 21105
rect 2165 21053 2217 21105
rect 2217 21053 2233 21105
rect 2233 21053 2285 21105
rect 2285 21053 2301 21105
rect 2301 21053 2353 21105
rect 2353 21053 2369 21105
rect 2369 21053 2421 21105
rect 2421 21053 2437 21105
rect 2437 21053 2489 21105
rect 2489 21053 2505 21105
rect 2505 21053 2557 21105
rect 2557 21053 2573 21105
rect 2573 21053 2625 21105
rect 2625 21053 2641 21105
rect 2641 21053 2663 21105
rect 2127 21041 2663 21053
rect 2127 20989 2149 21041
rect 2149 20989 2165 21041
rect 2165 20989 2217 21041
rect 2217 20989 2233 21041
rect 2233 20989 2285 21041
rect 2285 20989 2301 21041
rect 2301 20989 2353 21041
rect 2353 20989 2369 21041
rect 2369 20989 2421 21041
rect 2421 20989 2437 21041
rect 2437 20989 2489 21041
rect 2489 20989 2505 21041
rect 2505 20989 2557 21041
rect 2557 20989 2573 21041
rect 2573 20989 2625 21041
rect 2625 20989 2641 21041
rect 2641 20989 2663 21041
rect 2127 20977 2663 20989
rect 2127 20925 2149 20977
rect 2149 20925 2165 20977
rect 2165 20925 2217 20977
rect 2217 20925 2233 20977
rect 2233 20925 2285 20977
rect 2285 20925 2301 20977
rect 2301 20925 2353 20977
rect 2353 20925 2369 20977
rect 2369 20925 2421 20977
rect 2421 20925 2437 20977
rect 2437 20925 2489 20977
rect 2489 20925 2505 20977
rect 2505 20925 2557 20977
rect 2557 20925 2573 20977
rect 2573 20925 2625 20977
rect 2625 20925 2641 20977
rect 2641 20925 2663 20977
rect 2127 20913 2663 20925
rect 2127 20902 2149 20913
rect 2149 20902 2165 20913
rect 2165 20902 2217 20913
rect 2217 20902 2233 20913
rect 2233 20902 2285 20913
rect 2285 20902 2301 20913
rect 2301 20902 2353 20913
rect 2353 20902 2369 20913
rect 2369 20902 2421 20913
rect 2421 20902 2437 20913
rect 2437 20902 2489 20913
rect 2489 20902 2505 20913
rect 2505 20902 2557 20913
rect 2557 20902 2573 20913
rect 2573 20902 2625 20913
rect 2625 20902 2641 20913
rect 2641 20902 2663 20913
rect 2127 20861 2149 20877
rect 2149 20861 2165 20877
rect 2165 20861 2183 20877
rect 2207 20861 2217 20877
rect 2217 20861 2233 20877
rect 2233 20861 2263 20877
rect 2287 20861 2301 20877
rect 2301 20861 2343 20877
rect 2367 20861 2369 20877
rect 2369 20861 2421 20877
rect 2421 20861 2423 20877
rect 2447 20861 2489 20877
rect 2489 20861 2503 20877
rect 2527 20861 2557 20877
rect 2557 20861 2573 20877
rect 2573 20861 2583 20877
rect 2607 20861 2625 20877
rect 2625 20861 2641 20877
rect 2641 20861 2663 20877
rect 2127 20849 2183 20861
rect 2207 20849 2263 20861
rect 2287 20849 2343 20861
rect 2367 20849 2423 20861
rect 2447 20849 2503 20861
rect 2527 20849 2583 20861
rect 2607 20849 2663 20861
rect 2127 20821 2149 20849
rect 2149 20821 2165 20849
rect 2165 20821 2183 20849
rect 2207 20821 2217 20849
rect 2217 20821 2233 20849
rect 2233 20821 2263 20849
rect 2287 20821 2301 20849
rect 2301 20821 2343 20849
rect 2367 20821 2369 20849
rect 2369 20821 2421 20849
rect 2421 20821 2423 20849
rect 2447 20821 2489 20849
rect 2489 20821 2503 20849
rect 2527 20821 2557 20849
rect 2557 20821 2573 20849
rect 2573 20821 2583 20849
rect 2607 20821 2625 20849
rect 2625 20821 2641 20849
rect 2641 20821 2663 20849
rect 2127 20785 2183 20796
rect 2207 20785 2263 20796
rect 2287 20785 2343 20796
rect 2367 20785 2423 20796
rect 2447 20785 2503 20796
rect 2527 20785 2583 20796
rect 2607 20785 2663 20796
rect 2127 20740 2149 20785
rect 2149 20740 2165 20785
rect 2165 20740 2183 20785
rect 2207 20740 2217 20785
rect 2217 20740 2233 20785
rect 2233 20740 2263 20785
rect 2287 20740 2301 20785
rect 2301 20740 2343 20785
rect 2367 20740 2369 20785
rect 2369 20740 2421 20785
rect 2421 20740 2423 20785
rect 2447 20740 2489 20785
rect 2489 20740 2503 20785
rect 2527 20740 2557 20785
rect 2557 20740 2573 20785
rect 2573 20740 2583 20785
rect 2607 20740 2625 20785
rect 2625 20740 2641 20785
rect 2641 20740 2663 20785
rect 2127 20669 2149 20715
rect 2149 20669 2165 20715
rect 2165 20669 2183 20715
rect 2207 20669 2217 20715
rect 2217 20669 2233 20715
rect 2233 20669 2263 20715
rect 2287 20669 2301 20715
rect 2301 20669 2343 20715
rect 2367 20669 2369 20715
rect 2369 20669 2421 20715
rect 2421 20669 2423 20715
rect 2447 20669 2489 20715
rect 2489 20669 2503 20715
rect 2527 20669 2557 20715
rect 2557 20669 2573 20715
rect 2573 20669 2583 20715
rect 2607 20669 2625 20715
rect 2625 20669 2641 20715
rect 2641 20669 2663 20715
rect 2127 20659 2183 20669
rect 2207 20659 2263 20669
rect 2287 20659 2343 20669
rect 2367 20659 2423 20669
rect 2447 20659 2503 20669
rect 2527 20659 2583 20669
rect 2607 20659 2663 20669
rect 2127 20605 2149 20634
rect 2149 20605 2165 20634
rect 2165 20605 2183 20634
rect 2207 20605 2217 20634
rect 2217 20605 2233 20634
rect 2233 20605 2263 20634
rect 2287 20605 2301 20634
rect 2301 20605 2343 20634
rect 2367 20605 2369 20634
rect 2369 20605 2421 20634
rect 2421 20605 2423 20634
rect 2447 20605 2489 20634
rect 2489 20605 2503 20634
rect 2527 20605 2557 20634
rect 2557 20605 2573 20634
rect 2573 20605 2583 20634
rect 2607 20605 2625 20634
rect 2625 20605 2641 20634
rect 2641 20605 2663 20634
rect 2127 20593 2183 20605
rect 2207 20593 2263 20605
rect 2287 20593 2343 20605
rect 2367 20593 2423 20605
rect 2447 20593 2503 20605
rect 2527 20593 2583 20605
rect 2607 20593 2663 20605
rect 2127 20578 2149 20593
rect 2149 20578 2165 20593
rect 2165 20578 2183 20593
rect 2207 20578 2217 20593
rect 2217 20578 2233 20593
rect 2233 20578 2263 20593
rect 2287 20578 2301 20593
rect 2301 20578 2343 20593
rect 2367 20578 2369 20593
rect 2369 20578 2421 20593
rect 2421 20578 2423 20593
rect 2447 20578 2489 20593
rect 2489 20578 2503 20593
rect 2527 20578 2557 20593
rect 2557 20578 2573 20593
rect 2573 20578 2583 20593
rect 2607 20578 2625 20593
rect 2625 20578 2641 20593
rect 2641 20578 2663 20593
rect 2127 20541 2149 20553
rect 2149 20541 2165 20553
rect 2165 20541 2183 20553
rect 2207 20541 2217 20553
rect 2217 20541 2233 20553
rect 2233 20541 2263 20553
rect 2287 20541 2301 20553
rect 2301 20541 2343 20553
rect 2367 20541 2369 20553
rect 2369 20541 2421 20553
rect 2421 20541 2423 20553
rect 2447 20541 2489 20553
rect 2489 20541 2503 20553
rect 2527 20541 2557 20553
rect 2557 20541 2573 20553
rect 2573 20541 2583 20553
rect 2607 20541 2625 20553
rect 2625 20541 2641 20553
rect 2641 20541 2663 20553
rect 2127 20529 2183 20541
rect 2207 20529 2263 20541
rect 2287 20529 2343 20541
rect 2367 20529 2423 20541
rect 2447 20529 2503 20541
rect 2527 20529 2583 20541
rect 2607 20529 2663 20541
rect 2127 20497 2149 20529
rect 2149 20497 2165 20529
rect 2165 20497 2183 20529
rect 2207 20497 2217 20529
rect 2217 20497 2233 20529
rect 2233 20497 2263 20529
rect 2287 20497 2301 20529
rect 2301 20497 2343 20529
rect 2367 20497 2369 20529
rect 2369 20497 2421 20529
rect 2421 20497 2423 20529
rect 2447 20497 2489 20529
rect 2489 20497 2503 20529
rect 2527 20497 2557 20529
rect 2557 20497 2573 20529
rect 2573 20497 2583 20529
rect 2607 20497 2625 20529
rect 2625 20497 2641 20529
rect 2641 20497 2663 20529
rect 2127 20465 2183 20472
rect 2207 20465 2263 20472
rect 2287 20465 2343 20472
rect 2367 20465 2423 20472
rect 2447 20465 2503 20472
rect 2527 20465 2583 20472
rect 2607 20465 2663 20472
rect 2127 20416 2149 20465
rect 2149 20416 2165 20465
rect 2165 20416 2183 20465
rect 2207 20416 2217 20465
rect 2217 20416 2233 20465
rect 2233 20416 2263 20465
rect 2287 20416 2301 20465
rect 2301 20416 2343 20465
rect 2367 20416 2369 20465
rect 2369 20416 2421 20465
rect 2421 20416 2423 20465
rect 2447 20416 2489 20465
rect 2489 20416 2503 20465
rect 2527 20416 2557 20465
rect 2557 20416 2573 20465
rect 2573 20416 2583 20465
rect 2607 20416 2625 20465
rect 2625 20416 2641 20465
rect 2641 20416 2663 20465
rect 2127 19205 2149 19254
rect 2149 19205 2165 19254
rect 2165 19205 2217 19254
rect 2217 19205 2233 19254
rect 2233 19205 2285 19254
rect 2285 19205 2301 19254
rect 2301 19205 2353 19254
rect 2353 19205 2369 19254
rect 2369 19205 2421 19254
rect 2421 19205 2437 19254
rect 2437 19205 2489 19254
rect 2489 19205 2505 19254
rect 2505 19205 2557 19254
rect 2557 19205 2573 19254
rect 2573 19205 2625 19254
rect 2625 19205 2641 19254
rect 2641 19205 2663 19254
rect 2127 19193 2663 19205
rect 2127 19141 2149 19193
rect 2149 19141 2165 19193
rect 2165 19141 2217 19193
rect 2217 19141 2233 19193
rect 2233 19141 2285 19193
rect 2285 19141 2301 19193
rect 2301 19141 2353 19193
rect 2353 19141 2369 19193
rect 2369 19141 2421 19193
rect 2421 19141 2437 19193
rect 2437 19141 2489 19193
rect 2489 19141 2505 19193
rect 2505 19141 2557 19193
rect 2557 19141 2573 19193
rect 2573 19141 2625 19193
rect 2625 19141 2641 19193
rect 2641 19141 2663 19193
rect 2127 19129 2663 19141
rect 2127 19077 2149 19129
rect 2149 19077 2165 19129
rect 2165 19077 2217 19129
rect 2217 19077 2233 19129
rect 2233 19077 2285 19129
rect 2285 19077 2301 19129
rect 2301 19077 2353 19129
rect 2353 19077 2369 19129
rect 2369 19077 2421 19129
rect 2421 19077 2437 19129
rect 2437 19077 2489 19129
rect 2489 19077 2505 19129
rect 2505 19077 2557 19129
rect 2557 19077 2573 19129
rect 2573 19077 2625 19129
rect 2625 19077 2641 19129
rect 2641 19077 2663 19129
rect 2127 19065 2663 19077
rect 2127 19013 2149 19065
rect 2149 19013 2165 19065
rect 2165 19013 2217 19065
rect 2217 19013 2233 19065
rect 2233 19013 2285 19065
rect 2285 19013 2301 19065
rect 2301 19013 2353 19065
rect 2353 19013 2369 19065
rect 2369 19013 2421 19065
rect 2421 19013 2437 19065
rect 2437 19013 2489 19065
rect 2489 19013 2505 19065
rect 2505 19013 2557 19065
rect 2557 19013 2573 19065
rect 2573 19013 2625 19065
rect 2625 19013 2641 19065
rect 2641 19013 2663 19065
rect 2127 19001 2663 19013
rect 2127 18949 2149 19001
rect 2149 18949 2165 19001
rect 2165 18949 2217 19001
rect 2217 18949 2233 19001
rect 2233 18949 2285 19001
rect 2285 18949 2301 19001
rect 2301 18949 2353 19001
rect 2353 18949 2369 19001
rect 2369 18949 2421 19001
rect 2421 18949 2437 19001
rect 2437 18949 2489 19001
rect 2489 18949 2505 19001
rect 2505 18949 2557 19001
rect 2557 18949 2573 19001
rect 2573 18949 2625 19001
rect 2625 18949 2641 19001
rect 2641 18949 2663 19001
rect 2127 18937 2663 18949
rect 2127 18885 2149 18937
rect 2149 18885 2165 18937
rect 2165 18885 2217 18937
rect 2217 18885 2233 18937
rect 2233 18885 2285 18937
rect 2285 18885 2301 18937
rect 2301 18885 2353 18937
rect 2353 18885 2369 18937
rect 2369 18885 2421 18937
rect 2421 18885 2437 18937
rect 2437 18885 2489 18937
rect 2489 18885 2505 18937
rect 2505 18885 2557 18937
rect 2557 18885 2573 18937
rect 2573 18885 2625 18937
rect 2625 18885 2641 18937
rect 2641 18885 2663 18937
rect 2127 18873 2663 18885
rect 2127 18821 2149 18873
rect 2149 18821 2165 18873
rect 2165 18821 2217 18873
rect 2217 18821 2233 18873
rect 2233 18821 2285 18873
rect 2285 18821 2301 18873
rect 2301 18821 2353 18873
rect 2353 18821 2369 18873
rect 2369 18821 2421 18873
rect 2421 18821 2437 18873
rect 2437 18821 2489 18873
rect 2489 18821 2505 18873
rect 2505 18821 2557 18873
rect 2557 18821 2573 18873
rect 2573 18821 2625 18873
rect 2625 18821 2641 18873
rect 2641 18821 2663 18873
rect 2127 18809 2663 18821
rect 2127 18798 2149 18809
rect 2149 18798 2165 18809
rect 2165 18798 2217 18809
rect 2217 18798 2233 18809
rect 2233 18798 2285 18809
rect 2285 18798 2301 18809
rect 2301 18798 2353 18809
rect 2353 18798 2369 18809
rect 2369 18798 2421 18809
rect 2421 18798 2437 18809
rect 2437 18798 2489 18809
rect 2489 18798 2505 18809
rect 2505 18798 2557 18809
rect 2557 18798 2573 18809
rect 2573 18798 2625 18809
rect 2625 18798 2641 18809
rect 2641 18798 2663 18809
rect 2127 18757 2149 18773
rect 2149 18757 2165 18773
rect 2165 18757 2183 18773
rect 2207 18757 2217 18773
rect 2217 18757 2233 18773
rect 2233 18757 2263 18773
rect 2287 18757 2301 18773
rect 2301 18757 2343 18773
rect 2367 18757 2369 18773
rect 2369 18757 2421 18773
rect 2421 18757 2423 18773
rect 2447 18757 2489 18773
rect 2489 18757 2503 18773
rect 2527 18757 2557 18773
rect 2557 18757 2573 18773
rect 2573 18757 2583 18773
rect 2607 18757 2625 18773
rect 2625 18757 2641 18773
rect 2641 18757 2663 18773
rect 2127 18745 2183 18757
rect 2207 18745 2263 18757
rect 2287 18745 2343 18757
rect 2367 18745 2423 18757
rect 2447 18745 2503 18757
rect 2527 18745 2583 18757
rect 2607 18745 2663 18757
rect 2127 18717 2149 18745
rect 2149 18717 2165 18745
rect 2165 18717 2183 18745
rect 2207 18717 2217 18745
rect 2217 18717 2233 18745
rect 2233 18717 2263 18745
rect 2287 18717 2301 18745
rect 2301 18717 2343 18745
rect 2367 18717 2369 18745
rect 2369 18717 2421 18745
rect 2421 18717 2423 18745
rect 2447 18717 2489 18745
rect 2489 18717 2503 18745
rect 2527 18717 2557 18745
rect 2557 18717 2573 18745
rect 2573 18717 2583 18745
rect 2607 18717 2625 18745
rect 2625 18717 2641 18745
rect 2641 18717 2663 18745
rect 2127 18681 2183 18692
rect 2207 18681 2263 18692
rect 2287 18681 2343 18692
rect 2367 18681 2423 18692
rect 2447 18681 2503 18692
rect 2527 18681 2583 18692
rect 2607 18681 2663 18692
rect 2127 18636 2149 18681
rect 2149 18636 2165 18681
rect 2165 18636 2183 18681
rect 2207 18636 2217 18681
rect 2217 18636 2233 18681
rect 2233 18636 2263 18681
rect 2287 18636 2301 18681
rect 2301 18636 2343 18681
rect 2367 18636 2369 18681
rect 2369 18636 2421 18681
rect 2421 18636 2423 18681
rect 2447 18636 2489 18681
rect 2489 18636 2503 18681
rect 2527 18636 2557 18681
rect 2557 18636 2573 18681
rect 2573 18636 2583 18681
rect 2607 18636 2625 18681
rect 2625 18636 2641 18681
rect 2641 18636 2663 18681
rect 2127 18565 2149 18611
rect 2149 18565 2165 18611
rect 2165 18565 2183 18611
rect 2207 18565 2217 18611
rect 2217 18565 2233 18611
rect 2233 18565 2263 18611
rect 2287 18565 2301 18611
rect 2301 18565 2343 18611
rect 2367 18565 2369 18611
rect 2369 18565 2421 18611
rect 2421 18565 2423 18611
rect 2447 18565 2489 18611
rect 2489 18565 2503 18611
rect 2527 18565 2557 18611
rect 2557 18565 2573 18611
rect 2573 18565 2583 18611
rect 2607 18565 2625 18611
rect 2625 18565 2641 18611
rect 2641 18565 2663 18611
rect 2127 18555 2183 18565
rect 2207 18555 2263 18565
rect 2287 18555 2343 18565
rect 2367 18555 2423 18565
rect 2447 18555 2503 18565
rect 2527 18555 2583 18565
rect 2607 18555 2663 18565
rect 2127 18501 2149 18530
rect 2149 18501 2165 18530
rect 2165 18501 2183 18530
rect 2207 18501 2217 18530
rect 2217 18501 2233 18530
rect 2233 18501 2263 18530
rect 2287 18501 2301 18530
rect 2301 18501 2343 18530
rect 2367 18501 2369 18530
rect 2369 18501 2421 18530
rect 2421 18501 2423 18530
rect 2447 18501 2489 18530
rect 2489 18501 2503 18530
rect 2527 18501 2557 18530
rect 2557 18501 2573 18530
rect 2573 18501 2583 18530
rect 2607 18501 2625 18530
rect 2625 18501 2641 18530
rect 2641 18501 2663 18530
rect 2127 18489 2183 18501
rect 2207 18489 2263 18501
rect 2287 18489 2343 18501
rect 2367 18489 2423 18501
rect 2447 18489 2503 18501
rect 2527 18489 2583 18501
rect 2607 18489 2663 18501
rect 2127 18474 2149 18489
rect 2149 18474 2165 18489
rect 2165 18474 2183 18489
rect 2207 18474 2217 18489
rect 2217 18474 2233 18489
rect 2233 18474 2263 18489
rect 2287 18474 2301 18489
rect 2301 18474 2343 18489
rect 2367 18474 2369 18489
rect 2369 18474 2421 18489
rect 2421 18474 2423 18489
rect 2447 18474 2489 18489
rect 2489 18474 2503 18489
rect 2527 18474 2557 18489
rect 2557 18474 2573 18489
rect 2573 18474 2583 18489
rect 2607 18474 2625 18489
rect 2625 18474 2641 18489
rect 2641 18474 2663 18489
rect 2127 18437 2149 18449
rect 2149 18437 2165 18449
rect 2165 18437 2183 18449
rect 2207 18437 2217 18449
rect 2217 18437 2233 18449
rect 2233 18437 2263 18449
rect 2287 18437 2301 18449
rect 2301 18437 2343 18449
rect 2367 18437 2369 18449
rect 2369 18437 2421 18449
rect 2421 18437 2423 18449
rect 2447 18437 2489 18449
rect 2489 18437 2503 18449
rect 2527 18437 2557 18449
rect 2557 18437 2573 18449
rect 2573 18437 2583 18449
rect 2607 18437 2625 18449
rect 2625 18437 2641 18449
rect 2641 18437 2663 18449
rect 2127 18425 2183 18437
rect 2207 18425 2263 18437
rect 2287 18425 2343 18437
rect 2367 18425 2423 18437
rect 2447 18425 2503 18437
rect 2527 18425 2583 18437
rect 2607 18425 2663 18437
rect 2127 18393 2149 18425
rect 2149 18393 2165 18425
rect 2165 18393 2183 18425
rect 2207 18393 2217 18425
rect 2217 18393 2233 18425
rect 2233 18393 2263 18425
rect 2287 18393 2301 18425
rect 2301 18393 2343 18425
rect 2367 18393 2369 18425
rect 2369 18393 2421 18425
rect 2421 18393 2423 18425
rect 2447 18393 2489 18425
rect 2489 18393 2503 18425
rect 2527 18393 2557 18425
rect 2557 18393 2573 18425
rect 2573 18393 2583 18425
rect 2607 18393 2625 18425
rect 2625 18393 2641 18425
rect 2641 18393 2663 18425
rect 2127 18361 2183 18368
rect 2207 18361 2263 18368
rect 2287 18361 2343 18368
rect 2367 18361 2423 18368
rect 2447 18361 2503 18368
rect 2527 18361 2583 18368
rect 2607 18361 2663 18368
rect 2127 18312 2149 18361
rect 2149 18312 2165 18361
rect 2165 18312 2183 18361
rect 2207 18312 2217 18361
rect 2217 18312 2233 18361
rect 2233 18312 2263 18361
rect 2287 18312 2301 18361
rect 2301 18312 2343 18361
rect 2367 18312 2369 18361
rect 2369 18312 2421 18361
rect 2421 18312 2423 18361
rect 2447 18312 2489 18361
rect 2489 18312 2503 18361
rect 2527 18312 2557 18361
rect 2557 18312 2573 18361
rect 2573 18312 2583 18361
rect 2607 18312 2625 18361
rect 2625 18312 2641 18361
rect 2641 18312 2663 18361
rect 2127 17094 2149 17143
rect 2149 17094 2165 17143
rect 2165 17094 2217 17143
rect 2217 17094 2233 17143
rect 2233 17094 2285 17143
rect 2285 17094 2301 17143
rect 2301 17094 2353 17143
rect 2353 17094 2369 17143
rect 2369 17094 2421 17143
rect 2421 17094 2437 17143
rect 2437 17094 2489 17143
rect 2489 17094 2505 17143
rect 2505 17094 2557 17143
rect 2557 17094 2573 17143
rect 2573 17094 2625 17143
rect 2625 17094 2641 17143
rect 2641 17094 2663 17143
rect 2127 17082 2663 17094
rect 2127 17030 2149 17082
rect 2149 17030 2165 17082
rect 2165 17030 2217 17082
rect 2217 17030 2233 17082
rect 2233 17030 2285 17082
rect 2285 17030 2301 17082
rect 2301 17030 2353 17082
rect 2353 17030 2369 17082
rect 2369 17030 2421 17082
rect 2421 17030 2437 17082
rect 2437 17030 2489 17082
rect 2489 17030 2505 17082
rect 2505 17030 2557 17082
rect 2557 17030 2573 17082
rect 2573 17030 2625 17082
rect 2625 17030 2641 17082
rect 2641 17030 2663 17082
rect 2127 17018 2663 17030
rect 2127 16966 2149 17018
rect 2149 16966 2165 17018
rect 2165 16966 2217 17018
rect 2217 16966 2233 17018
rect 2233 16966 2285 17018
rect 2285 16966 2301 17018
rect 2301 16966 2353 17018
rect 2353 16966 2369 17018
rect 2369 16966 2421 17018
rect 2421 16966 2437 17018
rect 2437 16966 2489 17018
rect 2489 16966 2505 17018
rect 2505 16966 2557 17018
rect 2557 16966 2573 17018
rect 2573 16966 2625 17018
rect 2625 16966 2641 17018
rect 2641 16966 2663 17018
rect 2127 16954 2663 16966
rect 2127 16902 2149 16954
rect 2149 16902 2165 16954
rect 2165 16902 2217 16954
rect 2217 16902 2233 16954
rect 2233 16902 2285 16954
rect 2285 16902 2301 16954
rect 2301 16902 2353 16954
rect 2353 16902 2369 16954
rect 2369 16902 2421 16954
rect 2421 16902 2437 16954
rect 2437 16902 2489 16954
rect 2489 16902 2505 16954
rect 2505 16902 2557 16954
rect 2557 16902 2573 16954
rect 2573 16902 2625 16954
rect 2625 16902 2641 16954
rect 2641 16902 2663 16954
rect 2127 16890 2663 16902
rect 2127 16838 2149 16890
rect 2149 16838 2165 16890
rect 2165 16838 2217 16890
rect 2217 16838 2233 16890
rect 2233 16838 2285 16890
rect 2285 16838 2301 16890
rect 2301 16838 2353 16890
rect 2353 16838 2369 16890
rect 2369 16838 2421 16890
rect 2421 16838 2437 16890
rect 2437 16838 2489 16890
rect 2489 16838 2505 16890
rect 2505 16838 2557 16890
rect 2557 16838 2573 16890
rect 2573 16838 2625 16890
rect 2625 16838 2641 16890
rect 2641 16838 2663 16890
rect 2127 16826 2663 16838
rect 2127 16774 2149 16826
rect 2149 16774 2165 16826
rect 2165 16774 2217 16826
rect 2217 16774 2233 16826
rect 2233 16774 2285 16826
rect 2285 16774 2301 16826
rect 2301 16774 2353 16826
rect 2353 16774 2369 16826
rect 2369 16774 2421 16826
rect 2421 16774 2437 16826
rect 2437 16774 2489 16826
rect 2489 16774 2505 16826
rect 2505 16774 2557 16826
rect 2557 16774 2573 16826
rect 2573 16774 2625 16826
rect 2625 16774 2641 16826
rect 2641 16774 2663 16826
rect 2127 16762 2663 16774
rect 2127 16710 2149 16762
rect 2149 16710 2165 16762
rect 2165 16710 2217 16762
rect 2217 16710 2233 16762
rect 2233 16710 2285 16762
rect 2285 16710 2301 16762
rect 2301 16710 2353 16762
rect 2353 16710 2369 16762
rect 2369 16710 2421 16762
rect 2421 16710 2437 16762
rect 2437 16710 2489 16762
rect 2489 16710 2505 16762
rect 2505 16710 2557 16762
rect 2557 16710 2573 16762
rect 2573 16710 2625 16762
rect 2625 16710 2641 16762
rect 2641 16710 2663 16762
rect 2127 16698 2663 16710
rect 2127 16687 2149 16698
rect 2149 16687 2165 16698
rect 2165 16687 2217 16698
rect 2217 16687 2233 16698
rect 2233 16687 2285 16698
rect 2285 16687 2301 16698
rect 2301 16687 2353 16698
rect 2353 16687 2369 16698
rect 2369 16687 2421 16698
rect 2421 16687 2437 16698
rect 2437 16687 2489 16698
rect 2489 16687 2505 16698
rect 2505 16687 2557 16698
rect 2557 16687 2573 16698
rect 2573 16687 2625 16698
rect 2625 16687 2641 16698
rect 2641 16687 2663 16698
rect 2127 16646 2149 16662
rect 2149 16646 2165 16662
rect 2165 16646 2183 16662
rect 2207 16646 2217 16662
rect 2217 16646 2233 16662
rect 2233 16646 2263 16662
rect 2287 16646 2301 16662
rect 2301 16646 2343 16662
rect 2367 16646 2369 16662
rect 2369 16646 2421 16662
rect 2421 16646 2423 16662
rect 2447 16646 2489 16662
rect 2489 16646 2503 16662
rect 2527 16646 2557 16662
rect 2557 16646 2573 16662
rect 2573 16646 2583 16662
rect 2607 16646 2625 16662
rect 2625 16646 2641 16662
rect 2641 16646 2663 16662
rect 2127 16634 2183 16646
rect 2207 16634 2263 16646
rect 2287 16634 2343 16646
rect 2367 16634 2423 16646
rect 2447 16634 2503 16646
rect 2527 16634 2583 16646
rect 2607 16634 2663 16646
rect 2127 16606 2149 16634
rect 2149 16606 2165 16634
rect 2165 16606 2183 16634
rect 2207 16606 2217 16634
rect 2217 16606 2233 16634
rect 2233 16606 2263 16634
rect 2287 16606 2301 16634
rect 2301 16606 2343 16634
rect 2367 16606 2369 16634
rect 2369 16606 2421 16634
rect 2421 16606 2423 16634
rect 2447 16606 2489 16634
rect 2489 16606 2503 16634
rect 2527 16606 2557 16634
rect 2557 16606 2573 16634
rect 2573 16606 2583 16634
rect 2607 16606 2625 16634
rect 2625 16606 2641 16634
rect 2641 16606 2663 16634
rect 2127 16570 2183 16581
rect 2207 16570 2263 16581
rect 2287 16570 2343 16581
rect 2367 16570 2423 16581
rect 2447 16570 2503 16581
rect 2527 16570 2583 16581
rect 2607 16570 2663 16581
rect 2127 16525 2149 16570
rect 2149 16525 2165 16570
rect 2165 16525 2183 16570
rect 2207 16525 2217 16570
rect 2217 16525 2233 16570
rect 2233 16525 2263 16570
rect 2287 16525 2301 16570
rect 2301 16525 2343 16570
rect 2367 16525 2369 16570
rect 2369 16525 2421 16570
rect 2421 16525 2423 16570
rect 2447 16525 2489 16570
rect 2489 16525 2503 16570
rect 2527 16525 2557 16570
rect 2557 16525 2573 16570
rect 2573 16525 2583 16570
rect 2607 16525 2625 16570
rect 2625 16525 2641 16570
rect 2641 16525 2663 16570
rect 2127 16454 2149 16500
rect 2149 16454 2165 16500
rect 2165 16454 2183 16500
rect 2207 16454 2217 16500
rect 2217 16454 2233 16500
rect 2233 16454 2263 16500
rect 2287 16454 2301 16500
rect 2301 16454 2343 16500
rect 2367 16454 2369 16500
rect 2369 16454 2421 16500
rect 2421 16454 2423 16500
rect 2447 16454 2489 16500
rect 2489 16454 2503 16500
rect 2527 16454 2557 16500
rect 2557 16454 2573 16500
rect 2573 16454 2583 16500
rect 2607 16454 2625 16500
rect 2625 16454 2641 16500
rect 2641 16454 2663 16500
rect 2127 16444 2183 16454
rect 2207 16444 2263 16454
rect 2287 16444 2343 16454
rect 2367 16444 2423 16454
rect 2447 16444 2503 16454
rect 2527 16444 2583 16454
rect 2607 16444 2663 16454
rect 2127 16390 2149 16419
rect 2149 16390 2165 16419
rect 2165 16390 2183 16419
rect 2207 16390 2217 16419
rect 2217 16390 2233 16419
rect 2233 16390 2263 16419
rect 2287 16390 2301 16419
rect 2301 16390 2343 16419
rect 2367 16390 2369 16419
rect 2369 16390 2421 16419
rect 2421 16390 2423 16419
rect 2447 16390 2489 16419
rect 2489 16390 2503 16419
rect 2527 16390 2557 16419
rect 2557 16390 2573 16419
rect 2573 16390 2583 16419
rect 2607 16390 2625 16419
rect 2625 16390 2641 16419
rect 2641 16390 2663 16419
rect 2127 16378 2183 16390
rect 2207 16378 2263 16390
rect 2287 16378 2343 16390
rect 2367 16378 2423 16390
rect 2447 16378 2503 16390
rect 2527 16378 2583 16390
rect 2607 16378 2663 16390
rect 2127 16363 2149 16378
rect 2149 16363 2165 16378
rect 2165 16363 2183 16378
rect 2207 16363 2217 16378
rect 2217 16363 2233 16378
rect 2233 16363 2263 16378
rect 2287 16363 2301 16378
rect 2301 16363 2343 16378
rect 2367 16363 2369 16378
rect 2369 16363 2421 16378
rect 2421 16363 2423 16378
rect 2447 16363 2489 16378
rect 2489 16363 2503 16378
rect 2527 16363 2557 16378
rect 2557 16363 2573 16378
rect 2573 16363 2583 16378
rect 2607 16363 2625 16378
rect 2625 16363 2641 16378
rect 2641 16363 2663 16378
rect 2127 16326 2149 16338
rect 2149 16326 2165 16338
rect 2165 16326 2183 16338
rect 2207 16326 2217 16338
rect 2217 16326 2233 16338
rect 2233 16326 2263 16338
rect 2287 16326 2301 16338
rect 2301 16326 2343 16338
rect 2367 16326 2369 16338
rect 2369 16326 2421 16338
rect 2421 16326 2423 16338
rect 2447 16326 2489 16338
rect 2489 16326 2503 16338
rect 2527 16326 2557 16338
rect 2557 16326 2573 16338
rect 2573 16326 2583 16338
rect 2607 16326 2625 16338
rect 2625 16326 2641 16338
rect 2641 16326 2663 16338
rect 2127 16314 2183 16326
rect 2207 16314 2263 16326
rect 2287 16314 2343 16326
rect 2367 16314 2423 16326
rect 2447 16314 2503 16326
rect 2527 16314 2583 16326
rect 2607 16314 2663 16326
rect 2127 16282 2149 16314
rect 2149 16282 2165 16314
rect 2165 16282 2183 16314
rect 2207 16282 2217 16314
rect 2217 16282 2233 16314
rect 2233 16282 2263 16314
rect 2287 16282 2301 16314
rect 2301 16282 2343 16314
rect 2367 16282 2369 16314
rect 2369 16282 2421 16314
rect 2421 16282 2423 16314
rect 2447 16282 2489 16314
rect 2489 16282 2503 16314
rect 2527 16282 2557 16314
rect 2557 16282 2573 16314
rect 2573 16282 2583 16314
rect 2607 16282 2625 16314
rect 2625 16282 2641 16314
rect 2641 16282 2663 16314
rect 2127 16250 2183 16257
rect 2207 16250 2263 16257
rect 2287 16250 2343 16257
rect 2367 16250 2423 16257
rect 2447 16250 2503 16257
rect 2527 16250 2583 16257
rect 2607 16250 2663 16257
rect 2127 16201 2149 16250
rect 2149 16201 2165 16250
rect 2165 16201 2183 16250
rect 2207 16201 2217 16250
rect 2217 16201 2233 16250
rect 2233 16201 2263 16250
rect 2287 16201 2301 16250
rect 2301 16201 2343 16250
rect 2367 16201 2369 16250
rect 2369 16201 2421 16250
rect 2421 16201 2423 16250
rect 2447 16201 2489 16250
rect 2489 16201 2503 16250
rect 2527 16201 2557 16250
rect 2557 16201 2573 16250
rect 2573 16201 2583 16250
rect 2607 16201 2625 16250
rect 2625 16201 2641 16250
rect 2641 16201 2663 16250
rect 2127 14957 2149 15006
rect 2149 14957 2165 15006
rect 2165 14957 2217 15006
rect 2217 14957 2233 15006
rect 2233 14957 2285 15006
rect 2285 14957 2301 15006
rect 2301 14957 2353 15006
rect 2353 14957 2369 15006
rect 2369 14957 2421 15006
rect 2421 14957 2437 15006
rect 2437 14957 2489 15006
rect 2489 14957 2505 15006
rect 2505 14957 2557 15006
rect 2557 14957 2573 15006
rect 2573 14957 2625 15006
rect 2625 14957 2641 15006
rect 2641 14957 2663 15006
rect 2127 14945 2663 14957
rect 2127 14893 2149 14945
rect 2149 14893 2165 14945
rect 2165 14893 2217 14945
rect 2217 14893 2233 14945
rect 2233 14893 2285 14945
rect 2285 14893 2301 14945
rect 2301 14893 2353 14945
rect 2353 14893 2369 14945
rect 2369 14893 2421 14945
rect 2421 14893 2437 14945
rect 2437 14893 2489 14945
rect 2489 14893 2505 14945
rect 2505 14893 2557 14945
rect 2557 14893 2573 14945
rect 2573 14893 2625 14945
rect 2625 14893 2641 14945
rect 2641 14893 2663 14945
rect 2127 14881 2663 14893
rect 2127 14829 2149 14881
rect 2149 14829 2165 14881
rect 2165 14829 2217 14881
rect 2217 14829 2233 14881
rect 2233 14829 2285 14881
rect 2285 14829 2301 14881
rect 2301 14829 2353 14881
rect 2353 14829 2369 14881
rect 2369 14829 2421 14881
rect 2421 14829 2437 14881
rect 2437 14829 2489 14881
rect 2489 14829 2505 14881
rect 2505 14829 2557 14881
rect 2557 14829 2573 14881
rect 2573 14829 2625 14881
rect 2625 14829 2641 14881
rect 2641 14829 2663 14881
rect 2127 14817 2663 14829
rect 2127 14765 2149 14817
rect 2149 14765 2165 14817
rect 2165 14765 2217 14817
rect 2217 14765 2233 14817
rect 2233 14765 2285 14817
rect 2285 14765 2301 14817
rect 2301 14765 2353 14817
rect 2353 14765 2369 14817
rect 2369 14765 2421 14817
rect 2421 14765 2437 14817
rect 2437 14765 2489 14817
rect 2489 14765 2505 14817
rect 2505 14765 2557 14817
rect 2557 14765 2573 14817
rect 2573 14765 2625 14817
rect 2625 14765 2641 14817
rect 2641 14765 2663 14817
rect 2127 14753 2663 14765
rect 2127 14701 2149 14753
rect 2149 14701 2165 14753
rect 2165 14701 2217 14753
rect 2217 14701 2233 14753
rect 2233 14701 2285 14753
rect 2285 14701 2301 14753
rect 2301 14701 2353 14753
rect 2353 14701 2369 14753
rect 2369 14701 2421 14753
rect 2421 14701 2437 14753
rect 2437 14701 2489 14753
rect 2489 14701 2505 14753
rect 2505 14701 2557 14753
rect 2557 14701 2573 14753
rect 2573 14701 2625 14753
rect 2625 14701 2641 14753
rect 2641 14701 2663 14753
rect 2127 14689 2663 14701
rect 2127 14637 2149 14689
rect 2149 14637 2165 14689
rect 2165 14637 2217 14689
rect 2217 14637 2233 14689
rect 2233 14637 2285 14689
rect 2285 14637 2301 14689
rect 2301 14637 2353 14689
rect 2353 14637 2369 14689
rect 2369 14637 2421 14689
rect 2421 14637 2437 14689
rect 2437 14637 2489 14689
rect 2489 14637 2505 14689
rect 2505 14637 2557 14689
rect 2557 14637 2573 14689
rect 2573 14637 2625 14689
rect 2625 14637 2641 14689
rect 2641 14637 2663 14689
rect 2127 14625 2663 14637
rect 2127 14573 2149 14625
rect 2149 14573 2165 14625
rect 2165 14573 2217 14625
rect 2217 14573 2233 14625
rect 2233 14573 2285 14625
rect 2285 14573 2301 14625
rect 2301 14573 2353 14625
rect 2353 14573 2369 14625
rect 2369 14573 2421 14625
rect 2421 14573 2437 14625
rect 2437 14573 2489 14625
rect 2489 14573 2505 14625
rect 2505 14573 2557 14625
rect 2557 14573 2573 14625
rect 2573 14573 2625 14625
rect 2625 14573 2641 14625
rect 2641 14573 2663 14625
rect 2127 14561 2663 14573
rect 2127 14550 2149 14561
rect 2149 14550 2165 14561
rect 2165 14550 2217 14561
rect 2217 14550 2233 14561
rect 2233 14550 2285 14561
rect 2285 14550 2301 14561
rect 2301 14550 2353 14561
rect 2353 14550 2369 14561
rect 2369 14550 2421 14561
rect 2421 14550 2437 14561
rect 2437 14550 2489 14561
rect 2489 14550 2505 14561
rect 2505 14550 2557 14561
rect 2557 14550 2573 14561
rect 2573 14550 2625 14561
rect 2625 14550 2641 14561
rect 2641 14550 2663 14561
rect 2127 14509 2149 14525
rect 2149 14509 2165 14525
rect 2165 14509 2183 14525
rect 2207 14509 2217 14525
rect 2217 14509 2233 14525
rect 2233 14509 2263 14525
rect 2287 14509 2301 14525
rect 2301 14509 2343 14525
rect 2367 14509 2369 14525
rect 2369 14509 2421 14525
rect 2421 14509 2423 14525
rect 2447 14509 2489 14525
rect 2489 14509 2503 14525
rect 2527 14509 2557 14525
rect 2557 14509 2573 14525
rect 2573 14509 2583 14525
rect 2607 14509 2625 14525
rect 2625 14509 2641 14525
rect 2641 14509 2663 14525
rect 2127 14497 2183 14509
rect 2207 14497 2263 14509
rect 2287 14497 2343 14509
rect 2367 14497 2423 14509
rect 2447 14497 2503 14509
rect 2527 14497 2583 14509
rect 2607 14497 2663 14509
rect 2127 14469 2149 14497
rect 2149 14469 2165 14497
rect 2165 14469 2183 14497
rect 2207 14469 2217 14497
rect 2217 14469 2233 14497
rect 2233 14469 2263 14497
rect 2287 14469 2301 14497
rect 2301 14469 2343 14497
rect 2367 14469 2369 14497
rect 2369 14469 2421 14497
rect 2421 14469 2423 14497
rect 2447 14469 2489 14497
rect 2489 14469 2503 14497
rect 2527 14469 2557 14497
rect 2557 14469 2573 14497
rect 2573 14469 2583 14497
rect 2607 14469 2625 14497
rect 2625 14469 2641 14497
rect 2641 14469 2663 14497
rect 2127 14433 2183 14444
rect 2207 14433 2263 14444
rect 2287 14433 2343 14444
rect 2367 14433 2423 14444
rect 2447 14433 2503 14444
rect 2527 14433 2583 14444
rect 2607 14433 2663 14444
rect 2127 14388 2149 14433
rect 2149 14388 2165 14433
rect 2165 14388 2183 14433
rect 2207 14388 2217 14433
rect 2217 14388 2233 14433
rect 2233 14388 2263 14433
rect 2287 14388 2301 14433
rect 2301 14388 2343 14433
rect 2367 14388 2369 14433
rect 2369 14388 2421 14433
rect 2421 14388 2423 14433
rect 2447 14388 2489 14433
rect 2489 14388 2503 14433
rect 2527 14388 2557 14433
rect 2557 14388 2573 14433
rect 2573 14388 2583 14433
rect 2607 14388 2625 14433
rect 2625 14388 2641 14433
rect 2641 14388 2663 14433
rect 2127 14317 2149 14363
rect 2149 14317 2165 14363
rect 2165 14317 2183 14363
rect 2207 14317 2217 14363
rect 2217 14317 2233 14363
rect 2233 14317 2263 14363
rect 2287 14317 2301 14363
rect 2301 14317 2343 14363
rect 2367 14317 2369 14363
rect 2369 14317 2421 14363
rect 2421 14317 2423 14363
rect 2447 14317 2489 14363
rect 2489 14317 2503 14363
rect 2527 14317 2557 14363
rect 2557 14317 2573 14363
rect 2573 14317 2583 14363
rect 2607 14317 2625 14363
rect 2625 14317 2641 14363
rect 2641 14317 2663 14363
rect 2127 14307 2183 14317
rect 2207 14307 2263 14317
rect 2287 14307 2343 14317
rect 2367 14307 2423 14317
rect 2447 14307 2503 14317
rect 2527 14307 2583 14317
rect 2607 14307 2663 14317
rect 2127 14253 2149 14282
rect 2149 14253 2165 14282
rect 2165 14253 2183 14282
rect 2207 14253 2217 14282
rect 2217 14253 2233 14282
rect 2233 14253 2263 14282
rect 2287 14253 2301 14282
rect 2301 14253 2343 14282
rect 2367 14253 2369 14282
rect 2369 14253 2421 14282
rect 2421 14253 2423 14282
rect 2447 14253 2489 14282
rect 2489 14253 2503 14282
rect 2527 14253 2557 14282
rect 2557 14253 2573 14282
rect 2573 14253 2583 14282
rect 2607 14253 2625 14282
rect 2625 14253 2641 14282
rect 2641 14253 2663 14282
rect 2127 14241 2183 14253
rect 2207 14241 2263 14253
rect 2287 14241 2343 14253
rect 2367 14241 2423 14253
rect 2447 14241 2503 14253
rect 2527 14241 2583 14253
rect 2607 14241 2663 14253
rect 2127 14226 2149 14241
rect 2149 14226 2165 14241
rect 2165 14226 2183 14241
rect 2207 14226 2217 14241
rect 2217 14226 2233 14241
rect 2233 14226 2263 14241
rect 2287 14226 2301 14241
rect 2301 14226 2343 14241
rect 2367 14226 2369 14241
rect 2369 14226 2421 14241
rect 2421 14226 2423 14241
rect 2447 14226 2489 14241
rect 2489 14226 2503 14241
rect 2527 14226 2557 14241
rect 2557 14226 2573 14241
rect 2573 14226 2583 14241
rect 2607 14226 2625 14241
rect 2625 14226 2641 14241
rect 2641 14226 2663 14241
rect 2127 14189 2149 14201
rect 2149 14189 2165 14201
rect 2165 14189 2183 14201
rect 2207 14189 2217 14201
rect 2217 14189 2233 14201
rect 2233 14189 2263 14201
rect 2287 14189 2301 14201
rect 2301 14189 2343 14201
rect 2367 14189 2369 14201
rect 2369 14189 2421 14201
rect 2421 14189 2423 14201
rect 2447 14189 2489 14201
rect 2489 14189 2503 14201
rect 2527 14189 2557 14201
rect 2557 14189 2573 14201
rect 2573 14189 2583 14201
rect 2607 14189 2625 14201
rect 2625 14189 2641 14201
rect 2641 14189 2663 14201
rect 2127 14177 2183 14189
rect 2207 14177 2263 14189
rect 2287 14177 2343 14189
rect 2367 14177 2423 14189
rect 2447 14177 2503 14189
rect 2527 14177 2583 14189
rect 2607 14177 2663 14189
rect 2127 14145 2149 14177
rect 2149 14145 2165 14177
rect 2165 14145 2183 14177
rect 2207 14145 2217 14177
rect 2217 14145 2233 14177
rect 2233 14145 2263 14177
rect 2287 14145 2301 14177
rect 2301 14145 2343 14177
rect 2367 14145 2369 14177
rect 2369 14145 2421 14177
rect 2421 14145 2423 14177
rect 2447 14145 2489 14177
rect 2489 14145 2503 14177
rect 2527 14145 2557 14177
rect 2557 14145 2573 14177
rect 2573 14145 2583 14177
rect 2607 14145 2625 14177
rect 2625 14145 2641 14177
rect 2641 14145 2663 14177
rect 2127 14113 2183 14120
rect 2207 14113 2263 14120
rect 2287 14113 2343 14120
rect 2367 14113 2423 14120
rect 2447 14113 2503 14120
rect 2527 14113 2583 14120
rect 2607 14113 2663 14120
rect 2127 14064 2149 14113
rect 2149 14064 2165 14113
rect 2165 14064 2183 14113
rect 2207 14064 2217 14113
rect 2217 14064 2233 14113
rect 2233 14064 2263 14113
rect 2287 14064 2301 14113
rect 2301 14064 2343 14113
rect 2367 14064 2369 14113
rect 2369 14064 2421 14113
rect 2421 14064 2423 14113
rect 2447 14064 2489 14113
rect 2489 14064 2503 14113
rect 2527 14064 2557 14113
rect 2557 14064 2573 14113
rect 2573 14064 2583 14113
rect 2607 14064 2625 14113
rect 2625 14064 2641 14113
rect 2641 14064 2663 14113
rect 2127 12855 2149 12904
rect 2149 12855 2165 12904
rect 2165 12855 2217 12904
rect 2217 12855 2233 12904
rect 2233 12855 2285 12904
rect 2285 12855 2301 12904
rect 2301 12855 2353 12904
rect 2353 12855 2369 12904
rect 2369 12855 2421 12904
rect 2421 12855 2437 12904
rect 2437 12855 2489 12904
rect 2489 12855 2505 12904
rect 2505 12855 2557 12904
rect 2557 12855 2573 12904
rect 2573 12855 2625 12904
rect 2625 12855 2641 12904
rect 2641 12855 2663 12904
rect 2127 12843 2663 12855
rect 2127 12791 2149 12843
rect 2149 12791 2165 12843
rect 2165 12791 2217 12843
rect 2217 12791 2233 12843
rect 2233 12791 2285 12843
rect 2285 12791 2301 12843
rect 2301 12791 2353 12843
rect 2353 12791 2369 12843
rect 2369 12791 2421 12843
rect 2421 12791 2437 12843
rect 2437 12791 2489 12843
rect 2489 12791 2505 12843
rect 2505 12791 2557 12843
rect 2557 12791 2573 12843
rect 2573 12791 2625 12843
rect 2625 12791 2641 12843
rect 2641 12791 2663 12843
rect 3285 13649 3287 13698
rect 3287 13649 3339 13698
rect 3339 13649 3341 13698
rect 3285 13642 3341 13649
rect 3285 13581 3287 13617
rect 3287 13581 3339 13617
rect 3339 13581 3341 13617
rect 3285 13565 3341 13581
rect 3285 13561 3287 13565
rect 3287 13561 3339 13565
rect 3339 13561 3341 13565
rect 3285 13513 3287 13536
rect 3287 13513 3339 13536
rect 3339 13513 3341 13536
rect 3285 13496 3341 13513
rect 3285 13480 3287 13496
rect 3287 13480 3339 13496
rect 3339 13480 3341 13496
rect 3285 13444 3287 13455
rect 3287 13444 3339 13455
rect 3339 13444 3341 13455
rect 3285 13427 3341 13444
rect 3285 13399 3287 13427
rect 3287 13399 3339 13427
rect 3339 13399 3341 13427
rect 3285 13358 3341 13374
rect 3285 13318 3287 13358
rect 3287 13318 3339 13358
rect 3339 13318 3341 13358
rect 3285 13289 3341 13292
rect 3285 13237 3287 13289
rect 3287 13237 3339 13289
rect 3339 13237 3341 13289
rect 3285 13236 3341 13237
rect 3285 13168 3287 13210
rect 3287 13168 3339 13210
rect 3339 13168 3341 13210
rect 3285 13154 3341 13168
rect 3285 13099 3287 13128
rect 3287 13099 3339 13128
rect 3339 13099 3341 13128
rect 3285 13082 3341 13099
rect 3285 13072 3287 13082
rect 3287 13072 3339 13082
rect 3339 13072 3341 13082
rect 3285 13030 3287 13046
rect 3287 13030 3339 13046
rect 3339 13030 3341 13046
rect 3285 13013 3341 13030
rect 3285 12990 3287 13013
rect 3287 12990 3339 13013
rect 3339 12990 3341 13013
rect 3285 12961 3287 12964
rect 3287 12961 3339 12964
rect 3339 12961 3341 12964
rect 3285 12944 3341 12961
rect 3285 12908 3287 12944
rect 3287 12908 3339 12944
rect 3339 12908 3341 12944
rect 3285 12875 3341 12882
rect 3285 12826 3287 12875
rect 3287 12826 3339 12875
rect 3339 12826 3341 12875
rect 2127 12779 2663 12791
rect 2127 12727 2149 12779
rect 2149 12727 2165 12779
rect 2165 12727 2217 12779
rect 2217 12727 2233 12779
rect 2233 12727 2285 12779
rect 2285 12727 2301 12779
rect 2301 12727 2353 12779
rect 2353 12727 2369 12779
rect 2369 12727 2421 12779
rect 2421 12727 2437 12779
rect 2437 12727 2489 12779
rect 2489 12727 2505 12779
rect 2505 12727 2557 12779
rect 2557 12727 2573 12779
rect 2573 12727 2625 12779
rect 2625 12727 2641 12779
rect 2641 12727 2663 12779
rect 2127 12715 2663 12727
rect 2127 12663 2149 12715
rect 2149 12663 2165 12715
rect 2165 12663 2217 12715
rect 2217 12663 2233 12715
rect 2233 12663 2285 12715
rect 2285 12663 2301 12715
rect 2301 12663 2353 12715
rect 2353 12663 2369 12715
rect 2369 12663 2421 12715
rect 2421 12663 2437 12715
rect 2437 12663 2489 12715
rect 2489 12663 2505 12715
rect 2505 12663 2557 12715
rect 2557 12663 2573 12715
rect 2573 12663 2625 12715
rect 2625 12663 2641 12715
rect 2641 12663 2663 12715
rect 2127 12651 2663 12663
rect 2127 12599 2149 12651
rect 2149 12599 2165 12651
rect 2165 12599 2217 12651
rect 2217 12599 2233 12651
rect 2233 12599 2285 12651
rect 2285 12599 2301 12651
rect 2301 12599 2353 12651
rect 2353 12599 2369 12651
rect 2369 12599 2421 12651
rect 2421 12599 2437 12651
rect 2437 12599 2489 12651
rect 2489 12599 2505 12651
rect 2505 12599 2557 12651
rect 2557 12599 2573 12651
rect 2573 12599 2625 12651
rect 2625 12599 2641 12651
rect 2641 12599 2663 12651
rect 2127 12587 2663 12599
rect 2127 12535 2149 12587
rect 2149 12535 2165 12587
rect 2165 12535 2217 12587
rect 2217 12535 2233 12587
rect 2233 12535 2285 12587
rect 2285 12535 2301 12587
rect 2301 12535 2353 12587
rect 2353 12535 2369 12587
rect 2369 12535 2421 12587
rect 2421 12535 2437 12587
rect 2437 12535 2489 12587
rect 2489 12535 2505 12587
rect 2505 12535 2557 12587
rect 2557 12535 2573 12587
rect 2573 12535 2625 12587
rect 2625 12535 2641 12587
rect 2641 12535 2663 12587
rect 2127 12523 2663 12535
rect 2127 12471 2149 12523
rect 2149 12471 2165 12523
rect 2165 12471 2217 12523
rect 2217 12471 2233 12523
rect 2233 12471 2285 12523
rect 2285 12471 2301 12523
rect 2301 12471 2353 12523
rect 2353 12471 2369 12523
rect 2369 12471 2421 12523
rect 2421 12471 2437 12523
rect 2437 12471 2489 12523
rect 2489 12471 2505 12523
rect 2505 12471 2557 12523
rect 2557 12471 2573 12523
rect 2573 12471 2625 12523
rect 2625 12471 2641 12523
rect 2641 12471 2663 12523
rect 2127 12459 2663 12471
rect 2127 12448 2149 12459
rect 2149 12448 2165 12459
rect 2165 12448 2217 12459
rect 2217 12448 2233 12459
rect 2233 12448 2285 12459
rect 2285 12448 2301 12459
rect 2301 12448 2353 12459
rect 2353 12448 2369 12459
rect 2369 12448 2421 12459
rect 2421 12448 2437 12459
rect 2437 12448 2489 12459
rect 2489 12448 2505 12459
rect 2505 12448 2557 12459
rect 2557 12448 2573 12459
rect 2573 12448 2625 12459
rect 2625 12448 2641 12459
rect 2641 12448 2663 12459
rect 2127 12407 2149 12423
rect 2149 12407 2165 12423
rect 2165 12407 2183 12423
rect 2207 12407 2217 12423
rect 2217 12407 2233 12423
rect 2233 12407 2263 12423
rect 2287 12407 2301 12423
rect 2301 12407 2343 12423
rect 2367 12407 2369 12423
rect 2369 12407 2421 12423
rect 2421 12407 2423 12423
rect 2447 12407 2489 12423
rect 2489 12407 2503 12423
rect 2527 12407 2557 12423
rect 2557 12407 2573 12423
rect 2573 12407 2583 12423
rect 2607 12407 2625 12423
rect 2625 12407 2641 12423
rect 2641 12407 2663 12423
rect 2127 12395 2183 12407
rect 2207 12395 2263 12407
rect 2287 12395 2343 12407
rect 2367 12395 2423 12407
rect 2447 12395 2503 12407
rect 2527 12395 2583 12407
rect 2607 12395 2663 12407
rect 2127 12367 2149 12395
rect 2149 12367 2165 12395
rect 2165 12367 2183 12395
rect 2207 12367 2217 12395
rect 2217 12367 2233 12395
rect 2233 12367 2263 12395
rect 2287 12367 2301 12395
rect 2301 12367 2343 12395
rect 2367 12367 2369 12395
rect 2369 12367 2421 12395
rect 2421 12367 2423 12395
rect 2447 12367 2489 12395
rect 2489 12367 2503 12395
rect 2527 12367 2557 12395
rect 2557 12367 2573 12395
rect 2573 12367 2583 12395
rect 2607 12367 2625 12395
rect 2625 12367 2641 12395
rect 2641 12367 2663 12395
rect 2127 12331 2183 12342
rect 2207 12331 2263 12342
rect 2287 12331 2343 12342
rect 2367 12331 2423 12342
rect 2447 12331 2503 12342
rect 2527 12331 2583 12342
rect 2607 12331 2663 12342
rect 2127 12286 2149 12331
rect 2149 12286 2165 12331
rect 2165 12286 2183 12331
rect 2207 12286 2217 12331
rect 2217 12286 2233 12331
rect 2233 12286 2263 12331
rect 2287 12286 2301 12331
rect 2301 12286 2343 12331
rect 2367 12286 2369 12331
rect 2369 12286 2421 12331
rect 2421 12286 2423 12331
rect 2447 12286 2489 12331
rect 2489 12286 2503 12331
rect 2527 12286 2557 12331
rect 2557 12286 2573 12331
rect 2573 12286 2583 12331
rect 2607 12286 2625 12331
rect 2625 12286 2641 12331
rect 2641 12286 2663 12331
rect 2127 12215 2149 12261
rect 2149 12215 2165 12261
rect 2165 12215 2183 12261
rect 2207 12215 2217 12261
rect 2217 12215 2233 12261
rect 2233 12215 2263 12261
rect 2287 12215 2301 12261
rect 2301 12215 2343 12261
rect 2367 12215 2369 12261
rect 2369 12215 2421 12261
rect 2421 12215 2423 12261
rect 2447 12215 2489 12261
rect 2489 12215 2503 12261
rect 2527 12215 2557 12261
rect 2557 12215 2573 12261
rect 2573 12215 2583 12261
rect 2607 12215 2625 12261
rect 2625 12215 2641 12261
rect 2641 12215 2663 12261
rect 2127 12205 2183 12215
rect 2207 12205 2263 12215
rect 2287 12205 2343 12215
rect 2367 12205 2423 12215
rect 2447 12205 2503 12215
rect 2527 12205 2583 12215
rect 2607 12205 2663 12215
rect 2127 12151 2149 12180
rect 2149 12151 2165 12180
rect 2165 12151 2183 12180
rect 2207 12151 2217 12180
rect 2217 12151 2233 12180
rect 2233 12151 2263 12180
rect 2287 12151 2301 12180
rect 2301 12151 2343 12180
rect 2367 12151 2369 12180
rect 2369 12151 2421 12180
rect 2421 12151 2423 12180
rect 2447 12151 2489 12180
rect 2489 12151 2503 12180
rect 2527 12151 2557 12180
rect 2557 12151 2573 12180
rect 2573 12151 2583 12180
rect 2607 12151 2625 12180
rect 2625 12151 2641 12180
rect 2641 12151 2663 12180
rect 2127 12139 2183 12151
rect 2207 12139 2263 12151
rect 2287 12139 2343 12151
rect 2367 12139 2423 12151
rect 2447 12139 2503 12151
rect 2527 12139 2583 12151
rect 2607 12139 2663 12151
rect 2127 12124 2149 12139
rect 2149 12124 2165 12139
rect 2165 12124 2183 12139
rect 2207 12124 2217 12139
rect 2217 12124 2233 12139
rect 2233 12124 2263 12139
rect 2287 12124 2301 12139
rect 2301 12124 2343 12139
rect 2367 12124 2369 12139
rect 2369 12124 2421 12139
rect 2421 12124 2423 12139
rect 2447 12124 2489 12139
rect 2489 12124 2503 12139
rect 2527 12124 2557 12139
rect 2557 12124 2573 12139
rect 2573 12124 2583 12139
rect 2607 12124 2625 12139
rect 2625 12124 2641 12139
rect 2641 12124 2663 12139
rect 2127 12087 2149 12099
rect 2149 12087 2165 12099
rect 2165 12087 2183 12099
rect 2207 12087 2217 12099
rect 2217 12087 2233 12099
rect 2233 12087 2263 12099
rect 2287 12087 2301 12099
rect 2301 12087 2343 12099
rect 2367 12087 2369 12099
rect 2369 12087 2421 12099
rect 2421 12087 2423 12099
rect 2447 12087 2489 12099
rect 2489 12087 2503 12099
rect 2527 12087 2557 12099
rect 2557 12087 2573 12099
rect 2573 12087 2583 12099
rect 2607 12087 2625 12099
rect 2625 12087 2641 12099
rect 2641 12087 2663 12099
rect 2127 12075 2183 12087
rect 2207 12075 2263 12087
rect 2287 12075 2343 12087
rect 2367 12075 2423 12087
rect 2447 12075 2503 12087
rect 2527 12075 2583 12087
rect 2607 12075 2663 12087
rect 2127 12043 2149 12075
rect 2149 12043 2165 12075
rect 2165 12043 2183 12075
rect 2207 12043 2217 12075
rect 2217 12043 2233 12075
rect 2233 12043 2263 12075
rect 2287 12043 2301 12075
rect 2301 12043 2343 12075
rect 2367 12043 2369 12075
rect 2369 12043 2421 12075
rect 2421 12043 2423 12075
rect 2447 12043 2489 12075
rect 2489 12043 2503 12075
rect 2527 12043 2557 12075
rect 2557 12043 2573 12075
rect 2573 12043 2583 12075
rect 2607 12043 2625 12075
rect 2625 12043 2641 12075
rect 2641 12043 2663 12075
rect 2127 12011 2183 12018
rect 2207 12011 2263 12018
rect 2287 12011 2343 12018
rect 2367 12011 2423 12018
rect 2447 12011 2503 12018
rect 2527 12011 2583 12018
rect 2607 12011 2663 12018
rect 2127 11962 2149 12011
rect 2149 11962 2165 12011
rect 2165 11962 2183 12011
rect 2207 11962 2217 12011
rect 2217 11962 2233 12011
rect 2233 11962 2263 12011
rect 2287 11962 2301 12011
rect 2301 11962 2343 12011
rect 2367 11962 2369 12011
rect 2369 11962 2421 12011
rect 2421 11962 2423 12011
rect 2447 11962 2489 12011
rect 2489 11962 2503 12011
rect 2527 11962 2557 12011
rect 2557 11962 2573 12011
rect 2573 11962 2583 12011
rect 2607 11962 2625 12011
rect 2625 11962 2641 12011
rect 2641 11962 2663 12011
rect 2127 10761 2149 10810
rect 2149 10761 2165 10810
rect 2165 10761 2217 10810
rect 2217 10761 2233 10810
rect 2233 10761 2285 10810
rect 2285 10761 2301 10810
rect 2301 10761 2353 10810
rect 2353 10761 2369 10810
rect 2369 10761 2421 10810
rect 2421 10761 2437 10810
rect 2437 10761 2489 10810
rect 2489 10761 2505 10810
rect 2505 10761 2557 10810
rect 2557 10761 2573 10810
rect 2573 10761 2625 10810
rect 2625 10761 2641 10810
rect 2641 10761 2663 10810
rect 2127 10749 2663 10761
rect 2127 10697 2149 10749
rect 2149 10697 2165 10749
rect 2165 10697 2217 10749
rect 2217 10697 2233 10749
rect 2233 10697 2285 10749
rect 2285 10697 2301 10749
rect 2301 10697 2353 10749
rect 2353 10697 2369 10749
rect 2369 10697 2421 10749
rect 2421 10697 2437 10749
rect 2437 10697 2489 10749
rect 2489 10697 2505 10749
rect 2505 10697 2557 10749
rect 2557 10697 2573 10749
rect 2573 10697 2625 10749
rect 2625 10697 2641 10749
rect 2641 10697 2663 10749
rect 2127 10685 2663 10697
rect 2127 10633 2149 10685
rect 2149 10633 2165 10685
rect 2165 10633 2217 10685
rect 2217 10633 2233 10685
rect 2233 10633 2285 10685
rect 2285 10633 2301 10685
rect 2301 10633 2353 10685
rect 2353 10633 2369 10685
rect 2369 10633 2421 10685
rect 2421 10633 2437 10685
rect 2437 10633 2489 10685
rect 2489 10633 2505 10685
rect 2505 10633 2557 10685
rect 2557 10633 2573 10685
rect 2573 10633 2625 10685
rect 2625 10633 2641 10685
rect 2641 10633 2663 10685
rect 2127 10621 2663 10633
rect 2127 10569 2149 10621
rect 2149 10569 2165 10621
rect 2165 10569 2217 10621
rect 2217 10569 2233 10621
rect 2233 10569 2285 10621
rect 2285 10569 2301 10621
rect 2301 10569 2353 10621
rect 2353 10569 2369 10621
rect 2369 10569 2421 10621
rect 2421 10569 2437 10621
rect 2437 10569 2489 10621
rect 2489 10569 2505 10621
rect 2505 10569 2557 10621
rect 2557 10569 2573 10621
rect 2573 10569 2625 10621
rect 2625 10569 2641 10621
rect 2641 10569 2663 10621
rect 2127 10557 2663 10569
rect 2127 10505 2149 10557
rect 2149 10505 2165 10557
rect 2165 10505 2217 10557
rect 2217 10505 2233 10557
rect 2233 10505 2285 10557
rect 2285 10505 2301 10557
rect 2301 10505 2353 10557
rect 2353 10505 2369 10557
rect 2369 10505 2421 10557
rect 2421 10505 2437 10557
rect 2437 10505 2489 10557
rect 2489 10505 2505 10557
rect 2505 10505 2557 10557
rect 2557 10505 2573 10557
rect 2573 10505 2625 10557
rect 2625 10505 2641 10557
rect 2641 10505 2663 10557
rect 2127 10493 2663 10505
rect 2127 10441 2149 10493
rect 2149 10441 2165 10493
rect 2165 10441 2217 10493
rect 2217 10441 2233 10493
rect 2233 10441 2285 10493
rect 2285 10441 2301 10493
rect 2301 10441 2353 10493
rect 2353 10441 2369 10493
rect 2369 10441 2421 10493
rect 2421 10441 2437 10493
rect 2437 10441 2489 10493
rect 2489 10441 2505 10493
rect 2505 10441 2557 10493
rect 2557 10441 2573 10493
rect 2573 10441 2625 10493
rect 2625 10441 2641 10493
rect 2641 10441 2663 10493
rect 2127 10429 2663 10441
rect 2127 10377 2149 10429
rect 2149 10377 2165 10429
rect 2165 10377 2217 10429
rect 2217 10377 2233 10429
rect 2233 10377 2285 10429
rect 2285 10377 2301 10429
rect 2301 10377 2353 10429
rect 2353 10377 2369 10429
rect 2369 10377 2421 10429
rect 2421 10377 2437 10429
rect 2437 10377 2489 10429
rect 2489 10377 2505 10429
rect 2505 10377 2557 10429
rect 2557 10377 2573 10429
rect 2573 10377 2625 10429
rect 2625 10377 2641 10429
rect 2641 10377 2663 10429
rect 2127 10365 2663 10377
rect 2127 10354 2149 10365
rect 2149 10354 2165 10365
rect 2165 10354 2217 10365
rect 2217 10354 2233 10365
rect 2233 10354 2285 10365
rect 2285 10354 2301 10365
rect 2301 10354 2353 10365
rect 2353 10354 2369 10365
rect 2369 10354 2421 10365
rect 2421 10354 2437 10365
rect 2437 10354 2489 10365
rect 2489 10354 2505 10365
rect 2505 10354 2557 10365
rect 2557 10354 2573 10365
rect 2573 10354 2625 10365
rect 2625 10354 2641 10365
rect 2641 10354 2663 10365
rect 2127 10313 2149 10329
rect 2149 10313 2165 10329
rect 2165 10313 2183 10329
rect 2207 10313 2217 10329
rect 2217 10313 2233 10329
rect 2233 10313 2263 10329
rect 2287 10313 2301 10329
rect 2301 10313 2343 10329
rect 2367 10313 2369 10329
rect 2369 10313 2421 10329
rect 2421 10313 2423 10329
rect 2447 10313 2489 10329
rect 2489 10313 2503 10329
rect 2527 10313 2557 10329
rect 2557 10313 2573 10329
rect 2573 10313 2583 10329
rect 2607 10313 2625 10329
rect 2625 10313 2641 10329
rect 2641 10313 2663 10329
rect 2127 10301 2183 10313
rect 2207 10301 2263 10313
rect 2287 10301 2343 10313
rect 2367 10301 2423 10313
rect 2447 10301 2503 10313
rect 2527 10301 2583 10313
rect 2607 10301 2663 10313
rect 2127 10273 2149 10301
rect 2149 10273 2165 10301
rect 2165 10273 2183 10301
rect 2207 10273 2217 10301
rect 2217 10273 2233 10301
rect 2233 10273 2263 10301
rect 2287 10273 2301 10301
rect 2301 10273 2343 10301
rect 2367 10273 2369 10301
rect 2369 10273 2421 10301
rect 2421 10273 2423 10301
rect 2447 10273 2489 10301
rect 2489 10273 2503 10301
rect 2527 10273 2557 10301
rect 2557 10273 2573 10301
rect 2573 10273 2583 10301
rect 2607 10273 2625 10301
rect 2625 10273 2641 10301
rect 2641 10273 2663 10301
rect 2127 10237 2183 10248
rect 2207 10237 2263 10248
rect 2287 10237 2343 10248
rect 2367 10237 2423 10248
rect 2447 10237 2503 10248
rect 2527 10237 2583 10248
rect 2607 10237 2663 10248
rect 2127 10192 2149 10237
rect 2149 10192 2165 10237
rect 2165 10192 2183 10237
rect 2207 10192 2217 10237
rect 2217 10192 2233 10237
rect 2233 10192 2263 10237
rect 2287 10192 2301 10237
rect 2301 10192 2343 10237
rect 2367 10192 2369 10237
rect 2369 10192 2421 10237
rect 2421 10192 2423 10237
rect 2447 10192 2489 10237
rect 2489 10192 2503 10237
rect 2527 10192 2557 10237
rect 2557 10192 2573 10237
rect 2573 10192 2583 10237
rect 2607 10192 2625 10237
rect 2625 10192 2641 10237
rect 2641 10192 2663 10237
rect 2127 10121 2149 10167
rect 2149 10121 2165 10167
rect 2165 10121 2183 10167
rect 2207 10121 2217 10167
rect 2217 10121 2233 10167
rect 2233 10121 2263 10167
rect 2287 10121 2301 10167
rect 2301 10121 2343 10167
rect 2367 10121 2369 10167
rect 2369 10121 2421 10167
rect 2421 10121 2423 10167
rect 2447 10121 2489 10167
rect 2489 10121 2503 10167
rect 2527 10121 2557 10167
rect 2557 10121 2573 10167
rect 2573 10121 2583 10167
rect 2607 10121 2625 10167
rect 2625 10121 2641 10167
rect 2641 10121 2663 10167
rect 2127 10111 2183 10121
rect 2207 10111 2263 10121
rect 2287 10111 2343 10121
rect 2367 10111 2423 10121
rect 2447 10111 2503 10121
rect 2527 10111 2583 10121
rect 2607 10111 2663 10121
rect 2127 10057 2149 10086
rect 2149 10057 2165 10086
rect 2165 10057 2183 10086
rect 2207 10057 2217 10086
rect 2217 10057 2233 10086
rect 2233 10057 2263 10086
rect 2287 10057 2301 10086
rect 2301 10057 2343 10086
rect 2367 10057 2369 10086
rect 2369 10057 2421 10086
rect 2421 10057 2423 10086
rect 2447 10057 2489 10086
rect 2489 10057 2503 10086
rect 2527 10057 2557 10086
rect 2557 10057 2573 10086
rect 2573 10057 2583 10086
rect 2607 10057 2625 10086
rect 2625 10057 2641 10086
rect 2641 10057 2663 10086
rect 2127 10045 2183 10057
rect 2207 10045 2263 10057
rect 2287 10045 2343 10057
rect 2367 10045 2423 10057
rect 2447 10045 2503 10057
rect 2527 10045 2583 10057
rect 2607 10045 2663 10057
rect 2127 10030 2149 10045
rect 2149 10030 2165 10045
rect 2165 10030 2183 10045
rect 2207 10030 2217 10045
rect 2217 10030 2233 10045
rect 2233 10030 2263 10045
rect 2287 10030 2301 10045
rect 2301 10030 2343 10045
rect 2367 10030 2369 10045
rect 2369 10030 2421 10045
rect 2421 10030 2423 10045
rect 2447 10030 2489 10045
rect 2489 10030 2503 10045
rect 2527 10030 2557 10045
rect 2557 10030 2573 10045
rect 2573 10030 2583 10045
rect 2607 10030 2625 10045
rect 2625 10030 2641 10045
rect 2641 10030 2663 10045
rect 2127 9993 2149 10005
rect 2149 9993 2165 10005
rect 2165 9993 2183 10005
rect 2207 9993 2217 10005
rect 2217 9993 2233 10005
rect 2233 9993 2263 10005
rect 2287 9993 2301 10005
rect 2301 9993 2343 10005
rect 2367 9993 2369 10005
rect 2369 9993 2421 10005
rect 2421 9993 2423 10005
rect 2447 9993 2489 10005
rect 2489 9993 2503 10005
rect 2527 9993 2557 10005
rect 2557 9993 2573 10005
rect 2573 9993 2583 10005
rect 2607 9993 2625 10005
rect 2625 9993 2641 10005
rect 2641 9993 2663 10005
rect 2127 9981 2183 9993
rect 2207 9981 2263 9993
rect 2287 9981 2343 9993
rect 2367 9981 2423 9993
rect 2447 9981 2503 9993
rect 2527 9981 2583 9993
rect 2607 9981 2663 9993
rect 2127 9949 2149 9981
rect 2149 9949 2165 9981
rect 2165 9949 2183 9981
rect 2207 9949 2217 9981
rect 2217 9949 2233 9981
rect 2233 9949 2263 9981
rect 2287 9949 2301 9981
rect 2301 9949 2343 9981
rect 2367 9949 2369 9981
rect 2369 9949 2421 9981
rect 2421 9949 2423 9981
rect 2447 9949 2489 9981
rect 2489 9949 2503 9981
rect 2527 9949 2557 9981
rect 2557 9949 2573 9981
rect 2573 9949 2583 9981
rect 2607 9949 2625 9981
rect 2625 9949 2641 9981
rect 2641 9949 2663 9981
rect 2127 9917 2183 9924
rect 2207 9917 2263 9924
rect 2287 9917 2343 9924
rect 2367 9917 2423 9924
rect 2447 9917 2503 9924
rect 2527 9917 2583 9924
rect 2607 9917 2663 9924
rect 2127 9868 2149 9917
rect 2149 9868 2165 9917
rect 2165 9868 2183 9917
rect 2207 9868 2217 9917
rect 2217 9868 2233 9917
rect 2233 9868 2263 9917
rect 2287 9868 2301 9917
rect 2301 9868 2343 9917
rect 2367 9868 2369 9917
rect 2369 9868 2421 9917
rect 2421 9868 2423 9917
rect 2447 9868 2489 9917
rect 2489 9868 2503 9917
rect 2527 9868 2557 9917
rect 2557 9868 2573 9917
rect 2573 9868 2583 9917
rect 2607 9868 2625 9917
rect 2625 9868 2641 9917
rect 2641 9868 2663 9917
rect 2127 8559 2149 8608
rect 2149 8559 2165 8608
rect 2165 8559 2217 8608
rect 2217 8559 2233 8608
rect 2233 8559 2285 8608
rect 2285 8559 2301 8608
rect 2301 8559 2353 8608
rect 2353 8559 2369 8608
rect 2369 8559 2421 8608
rect 2421 8559 2437 8608
rect 2437 8559 2489 8608
rect 2489 8559 2505 8608
rect 2505 8559 2557 8608
rect 2557 8559 2573 8608
rect 2573 8559 2625 8608
rect 2625 8559 2641 8608
rect 2641 8559 2663 8608
rect 2127 8547 2663 8559
rect 2127 8495 2149 8547
rect 2149 8495 2165 8547
rect 2165 8495 2217 8547
rect 2217 8495 2233 8547
rect 2233 8495 2285 8547
rect 2285 8495 2301 8547
rect 2301 8495 2353 8547
rect 2353 8495 2369 8547
rect 2369 8495 2421 8547
rect 2421 8495 2437 8547
rect 2437 8495 2489 8547
rect 2489 8495 2505 8547
rect 2505 8495 2557 8547
rect 2557 8495 2573 8547
rect 2573 8495 2625 8547
rect 2625 8495 2641 8547
rect 2641 8495 2663 8547
rect 2127 8483 2663 8495
rect 2127 8431 2149 8483
rect 2149 8431 2165 8483
rect 2165 8431 2217 8483
rect 2217 8431 2233 8483
rect 2233 8431 2285 8483
rect 2285 8431 2301 8483
rect 2301 8431 2353 8483
rect 2353 8431 2369 8483
rect 2369 8431 2421 8483
rect 2421 8431 2437 8483
rect 2437 8431 2489 8483
rect 2489 8431 2505 8483
rect 2505 8431 2557 8483
rect 2557 8431 2573 8483
rect 2573 8431 2625 8483
rect 2625 8431 2641 8483
rect 2641 8431 2663 8483
rect 2127 8419 2663 8431
rect 2127 8367 2149 8419
rect 2149 8367 2165 8419
rect 2165 8367 2217 8419
rect 2217 8367 2233 8419
rect 2233 8367 2285 8419
rect 2285 8367 2301 8419
rect 2301 8367 2353 8419
rect 2353 8367 2369 8419
rect 2369 8367 2421 8419
rect 2421 8367 2437 8419
rect 2437 8367 2489 8419
rect 2489 8367 2505 8419
rect 2505 8367 2557 8419
rect 2557 8367 2573 8419
rect 2573 8367 2625 8419
rect 2625 8367 2641 8419
rect 2641 8367 2663 8419
rect 2127 8355 2663 8367
rect 2127 8303 2149 8355
rect 2149 8303 2165 8355
rect 2165 8303 2217 8355
rect 2217 8303 2233 8355
rect 2233 8303 2285 8355
rect 2285 8303 2301 8355
rect 2301 8303 2353 8355
rect 2353 8303 2369 8355
rect 2369 8303 2421 8355
rect 2421 8303 2437 8355
rect 2437 8303 2489 8355
rect 2489 8303 2505 8355
rect 2505 8303 2557 8355
rect 2557 8303 2573 8355
rect 2573 8303 2625 8355
rect 2625 8303 2641 8355
rect 2641 8303 2663 8355
rect 2127 8291 2663 8303
rect 2127 8239 2149 8291
rect 2149 8239 2165 8291
rect 2165 8239 2217 8291
rect 2217 8239 2233 8291
rect 2233 8239 2285 8291
rect 2285 8239 2301 8291
rect 2301 8239 2353 8291
rect 2353 8239 2369 8291
rect 2369 8239 2421 8291
rect 2421 8239 2437 8291
rect 2437 8239 2489 8291
rect 2489 8239 2505 8291
rect 2505 8239 2557 8291
rect 2557 8239 2573 8291
rect 2573 8239 2625 8291
rect 2625 8239 2641 8291
rect 2641 8239 2663 8291
rect 2127 8227 2663 8239
rect 2127 8175 2149 8227
rect 2149 8175 2165 8227
rect 2165 8175 2217 8227
rect 2217 8175 2233 8227
rect 2233 8175 2285 8227
rect 2285 8175 2301 8227
rect 2301 8175 2353 8227
rect 2353 8175 2369 8227
rect 2369 8175 2421 8227
rect 2421 8175 2437 8227
rect 2437 8175 2489 8227
rect 2489 8175 2505 8227
rect 2505 8175 2557 8227
rect 2557 8175 2573 8227
rect 2573 8175 2625 8227
rect 2625 8175 2641 8227
rect 2641 8175 2663 8227
rect 2127 8163 2663 8175
rect 2127 8152 2149 8163
rect 2149 8152 2165 8163
rect 2165 8152 2217 8163
rect 2217 8152 2233 8163
rect 2233 8152 2285 8163
rect 2285 8152 2301 8163
rect 2301 8152 2353 8163
rect 2353 8152 2369 8163
rect 2369 8152 2421 8163
rect 2421 8152 2437 8163
rect 2437 8152 2489 8163
rect 2489 8152 2505 8163
rect 2505 8152 2557 8163
rect 2557 8152 2573 8163
rect 2573 8152 2625 8163
rect 2625 8152 2641 8163
rect 2641 8152 2663 8163
rect 2127 8111 2149 8127
rect 2149 8111 2165 8127
rect 2165 8111 2183 8127
rect 2207 8111 2217 8127
rect 2217 8111 2233 8127
rect 2233 8111 2263 8127
rect 2287 8111 2301 8127
rect 2301 8111 2343 8127
rect 2367 8111 2369 8127
rect 2369 8111 2421 8127
rect 2421 8111 2423 8127
rect 2447 8111 2489 8127
rect 2489 8111 2503 8127
rect 2527 8111 2557 8127
rect 2557 8111 2573 8127
rect 2573 8111 2583 8127
rect 2607 8111 2625 8127
rect 2625 8111 2641 8127
rect 2641 8111 2663 8127
rect 2127 8099 2183 8111
rect 2207 8099 2263 8111
rect 2287 8099 2343 8111
rect 2367 8099 2423 8111
rect 2447 8099 2503 8111
rect 2527 8099 2583 8111
rect 2607 8099 2663 8111
rect 2127 8071 2149 8099
rect 2149 8071 2165 8099
rect 2165 8071 2183 8099
rect 2207 8071 2217 8099
rect 2217 8071 2233 8099
rect 2233 8071 2263 8099
rect 2287 8071 2301 8099
rect 2301 8071 2343 8099
rect 2367 8071 2369 8099
rect 2369 8071 2421 8099
rect 2421 8071 2423 8099
rect 2447 8071 2489 8099
rect 2489 8071 2503 8099
rect 2527 8071 2557 8099
rect 2557 8071 2573 8099
rect 2573 8071 2583 8099
rect 2607 8071 2625 8099
rect 2625 8071 2641 8099
rect 2641 8071 2663 8099
rect 2127 8035 2183 8046
rect 2207 8035 2263 8046
rect 2287 8035 2343 8046
rect 2367 8035 2423 8046
rect 2447 8035 2503 8046
rect 2527 8035 2583 8046
rect 2607 8035 2663 8046
rect 2127 7990 2149 8035
rect 2149 7990 2165 8035
rect 2165 7990 2183 8035
rect 2207 7990 2217 8035
rect 2217 7990 2233 8035
rect 2233 7990 2263 8035
rect 2287 7990 2301 8035
rect 2301 7990 2343 8035
rect 2367 7990 2369 8035
rect 2369 7990 2421 8035
rect 2421 7990 2423 8035
rect 2447 7990 2489 8035
rect 2489 7990 2503 8035
rect 2527 7990 2557 8035
rect 2557 7990 2573 8035
rect 2573 7990 2583 8035
rect 2607 7990 2625 8035
rect 2625 7990 2641 8035
rect 2641 7990 2663 8035
rect 2127 7919 2149 7965
rect 2149 7919 2165 7965
rect 2165 7919 2183 7965
rect 2207 7919 2217 7965
rect 2217 7919 2233 7965
rect 2233 7919 2263 7965
rect 2287 7919 2301 7965
rect 2301 7919 2343 7965
rect 2367 7919 2369 7965
rect 2369 7919 2421 7965
rect 2421 7919 2423 7965
rect 2447 7919 2489 7965
rect 2489 7919 2503 7965
rect 2527 7919 2557 7965
rect 2557 7919 2573 7965
rect 2573 7919 2583 7965
rect 2607 7919 2625 7965
rect 2625 7919 2641 7965
rect 2641 7919 2663 7965
rect 2127 7909 2183 7919
rect 2207 7909 2263 7919
rect 2287 7909 2343 7919
rect 2367 7909 2423 7919
rect 2447 7909 2503 7919
rect 2527 7909 2583 7919
rect 2607 7909 2663 7919
rect 2127 7855 2149 7884
rect 2149 7855 2165 7884
rect 2165 7855 2183 7884
rect 2207 7855 2217 7884
rect 2217 7855 2233 7884
rect 2233 7855 2263 7884
rect 2287 7855 2301 7884
rect 2301 7855 2343 7884
rect 2367 7855 2369 7884
rect 2369 7855 2421 7884
rect 2421 7855 2423 7884
rect 2447 7855 2489 7884
rect 2489 7855 2503 7884
rect 2527 7855 2557 7884
rect 2557 7855 2573 7884
rect 2573 7855 2583 7884
rect 2607 7855 2625 7884
rect 2625 7855 2641 7884
rect 2641 7855 2663 7884
rect 2127 7843 2183 7855
rect 2207 7843 2263 7855
rect 2287 7843 2343 7855
rect 2367 7843 2423 7855
rect 2447 7843 2503 7855
rect 2527 7843 2583 7855
rect 2607 7843 2663 7855
rect 2127 7828 2149 7843
rect 2149 7828 2165 7843
rect 2165 7828 2183 7843
rect 2207 7828 2217 7843
rect 2217 7828 2233 7843
rect 2233 7828 2263 7843
rect 2287 7828 2301 7843
rect 2301 7828 2343 7843
rect 2367 7828 2369 7843
rect 2369 7828 2421 7843
rect 2421 7828 2423 7843
rect 2447 7828 2489 7843
rect 2489 7828 2503 7843
rect 2527 7828 2557 7843
rect 2557 7828 2573 7843
rect 2573 7828 2583 7843
rect 2607 7828 2625 7843
rect 2625 7828 2641 7843
rect 2641 7828 2663 7843
rect 2127 7791 2149 7803
rect 2149 7791 2165 7803
rect 2165 7791 2183 7803
rect 2207 7791 2217 7803
rect 2217 7791 2233 7803
rect 2233 7791 2263 7803
rect 2287 7791 2301 7803
rect 2301 7791 2343 7803
rect 2367 7791 2369 7803
rect 2369 7791 2421 7803
rect 2421 7791 2423 7803
rect 2447 7791 2489 7803
rect 2489 7791 2503 7803
rect 2527 7791 2557 7803
rect 2557 7791 2573 7803
rect 2573 7791 2583 7803
rect 2607 7791 2625 7803
rect 2625 7791 2641 7803
rect 2641 7791 2663 7803
rect 2127 7779 2183 7791
rect 2207 7779 2263 7791
rect 2287 7779 2343 7791
rect 2367 7779 2423 7791
rect 2447 7779 2503 7791
rect 2527 7779 2583 7791
rect 2607 7779 2663 7791
rect 2127 7747 2149 7779
rect 2149 7747 2165 7779
rect 2165 7747 2183 7779
rect 2207 7747 2217 7779
rect 2217 7747 2233 7779
rect 2233 7747 2263 7779
rect 2287 7747 2301 7779
rect 2301 7747 2343 7779
rect 2367 7747 2369 7779
rect 2369 7747 2421 7779
rect 2421 7747 2423 7779
rect 2447 7747 2489 7779
rect 2489 7747 2503 7779
rect 2527 7747 2557 7779
rect 2557 7747 2573 7779
rect 2573 7747 2583 7779
rect 2607 7747 2625 7779
rect 2625 7747 2641 7779
rect 2641 7747 2663 7779
rect 2127 7715 2183 7722
rect 2207 7715 2263 7722
rect 2287 7715 2343 7722
rect 2367 7715 2423 7722
rect 2447 7715 2503 7722
rect 2527 7715 2583 7722
rect 2607 7715 2663 7722
rect 2127 7666 2149 7715
rect 2149 7666 2165 7715
rect 2165 7666 2183 7715
rect 2207 7666 2217 7715
rect 2217 7666 2233 7715
rect 2233 7666 2263 7715
rect 2287 7666 2301 7715
rect 2301 7666 2343 7715
rect 2367 7666 2369 7715
rect 2369 7666 2421 7715
rect 2421 7666 2423 7715
rect 2447 7666 2489 7715
rect 2489 7666 2503 7715
rect 2527 7666 2557 7715
rect 2557 7666 2573 7715
rect 2573 7666 2583 7715
rect 2607 7666 2625 7715
rect 2625 7666 2641 7715
rect 2641 7666 2663 7715
rect 2127 6449 2149 6498
rect 2149 6449 2165 6498
rect 2165 6449 2217 6498
rect 2217 6449 2233 6498
rect 2233 6449 2285 6498
rect 2285 6449 2301 6498
rect 2301 6449 2353 6498
rect 2353 6449 2369 6498
rect 2369 6449 2421 6498
rect 2421 6449 2437 6498
rect 2437 6449 2489 6498
rect 2489 6449 2505 6498
rect 2505 6449 2557 6498
rect 2557 6449 2573 6498
rect 2573 6449 2625 6498
rect 2625 6449 2641 6498
rect 2641 6449 2663 6498
rect 2127 6437 2663 6449
rect 2127 6385 2149 6437
rect 2149 6385 2165 6437
rect 2165 6385 2217 6437
rect 2217 6385 2233 6437
rect 2233 6385 2285 6437
rect 2285 6385 2301 6437
rect 2301 6385 2353 6437
rect 2353 6385 2369 6437
rect 2369 6385 2421 6437
rect 2421 6385 2437 6437
rect 2437 6385 2489 6437
rect 2489 6385 2505 6437
rect 2505 6385 2557 6437
rect 2557 6385 2573 6437
rect 2573 6385 2625 6437
rect 2625 6385 2641 6437
rect 2641 6385 2663 6437
rect 2127 6373 2663 6385
rect 2127 6321 2149 6373
rect 2149 6321 2165 6373
rect 2165 6321 2217 6373
rect 2217 6321 2233 6373
rect 2233 6321 2285 6373
rect 2285 6321 2301 6373
rect 2301 6321 2353 6373
rect 2353 6321 2369 6373
rect 2369 6321 2421 6373
rect 2421 6321 2437 6373
rect 2437 6321 2489 6373
rect 2489 6321 2505 6373
rect 2505 6321 2557 6373
rect 2557 6321 2573 6373
rect 2573 6321 2625 6373
rect 2625 6321 2641 6373
rect 2641 6321 2663 6373
rect 2127 6309 2663 6321
rect 2127 6257 2149 6309
rect 2149 6257 2165 6309
rect 2165 6257 2217 6309
rect 2217 6257 2233 6309
rect 2233 6257 2285 6309
rect 2285 6257 2301 6309
rect 2301 6257 2353 6309
rect 2353 6257 2369 6309
rect 2369 6257 2421 6309
rect 2421 6257 2437 6309
rect 2437 6257 2489 6309
rect 2489 6257 2505 6309
rect 2505 6257 2557 6309
rect 2557 6257 2573 6309
rect 2573 6257 2625 6309
rect 2625 6257 2641 6309
rect 2641 6257 2663 6309
rect 2127 6245 2663 6257
rect 2127 6193 2149 6245
rect 2149 6193 2165 6245
rect 2165 6193 2217 6245
rect 2217 6193 2233 6245
rect 2233 6193 2285 6245
rect 2285 6193 2301 6245
rect 2301 6193 2353 6245
rect 2353 6193 2369 6245
rect 2369 6193 2421 6245
rect 2421 6193 2437 6245
rect 2437 6193 2489 6245
rect 2489 6193 2505 6245
rect 2505 6193 2557 6245
rect 2557 6193 2573 6245
rect 2573 6193 2625 6245
rect 2625 6193 2641 6245
rect 2641 6193 2663 6245
rect 2127 6181 2663 6193
rect 2127 6129 2149 6181
rect 2149 6129 2165 6181
rect 2165 6129 2217 6181
rect 2217 6129 2233 6181
rect 2233 6129 2285 6181
rect 2285 6129 2301 6181
rect 2301 6129 2353 6181
rect 2353 6129 2369 6181
rect 2369 6129 2421 6181
rect 2421 6129 2437 6181
rect 2437 6129 2489 6181
rect 2489 6129 2505 6181
rect 2505 6129 2557 6181
rect 2557 6129 2573 6181
rect 2573 6129 2625 6181
rect 2625 6129 2641 6181
rect 2641 6129 2663 6181
rect 2127 6117 2663 6129
rect 2127 6065 2149 6117
rect 2149 6065 2165 6117
rect 2165 6065 2217 6117
rect 2217 6065 2233 6117
rect 2233 6065 2285 6117
rect 2285 6065 2301 6117
rect 2301 6065 2353 6117
rect 2353 6065 2369 6117
rect 2369 6065 2421 6117
rect 2421 6065 2437 6117
rect 2437 6065 2489 6117
rect 2489 6065 2505 6117
rect 2505 6065 2557 6117
rect 2557 6065 2573 6117
rect 2573 6065 2625 6117
rect 2625 6065 2641 6117
rect 2641 6065 2663 6117
rect 2127 6053 2663 6065
rect 2127 6042 2149 6053
rect 2149 6042 2165 6053
rect 2165 6042 2217 6053
rect 2217 6042 2233 6053
rect 2233 6042 2285 6053
rect 2285 6042 2301 6053
rect 2301 6042 2353 6053
rect 2353 6042 2369 6053
rect 2369 6042 2421 6053
rect 2421 6042 2437 6053
rect 2437 6042 2489 6053
rect 2489 6042 2505 6053
rect 2505 6042 2557 6053
rect 2557 6042 2573 6053
rect 2573 6042 2625 6053
rect 2625 6042 2641 6053
rect 2641 6042 2663 6053
rect 2127 6001 2149 6017
rect 2149 6001 2165 6017
rect 2165 6001 2183 6017
rect 2207 6001 2217 6017
rect 2217 6001 2233 6017
rect 2233 6001 2263 6017
rect 2287 6001 2301 6017
rect 2301 6001 2343 6017
rect 2367 6001 2369 6017
rect 2369 6001 2421 6017
rect 2421 6001 2423 6017
rect 2447 6001 2489 6017
rect 2489 6001 2503 6017
rect 2527 6001 2557 6017
rect 2557 6001 2573 6017
rect 2573 6001 2583 6017
rect 2607 6001 2625 6017
rect 2625 6001 2641 6017
rect 2641 6001 2663 6017
rect 2127 5989 2183 6001
rect 2207 5989 2263 6001
rect 2287 5989 2343 6001
rect 2367 5989 2423 6001
rect 2447 5989 2503 6001
rect 2527 5989 2583 6001
rect 2607 5989 2663 6001
rect 2127 5961 2149 5989
rect 2149 5961 2165 5989
rect 2165 5961 2183 5989
rect 2207 5961 2217 5989
rect 2217 5961 2233 5989
rect 2233 5961 2263 5989
rect 2287 5961 2301 5989
rect 2301 5961 2343 5989
rect 2367 5961 2369 5989
rect 2369 5961 2421 5989
rect 2421 5961 2423 5989
rect 2447 5961 2489 5989
rect 2489 5961 2503 5989
rect 2527 5961 2557 5989
rect 2557 5961 2573 5989
rect 2573 5961 2583 5989
rect 2607 5961 2625 5989
rect 2625 5961 2641 5989
rect 2641 5961 2663 5989
rect 2127 5925 2183 5936
rect 2207 5925 2263 5936
rect 2287 5925 2343 5936
rect 2367 5925 2423 5936
rect 2447 5925 2503 5936
rect 2527 5925 2583 5936
rect 2607 5925 2663 5936
rect 2127 5880 2149 5925
rect 2149 5880 2165 5925
rect 2165 5880 2183 5925
rect 2207 5880 2217 5925
rect 2217 5880 2233 5925
rect 2233 5880 2263 5925
rect 2287 5880 2301 5925
rect 2301 5880 2343 5925
rect 2367 5880 2369 5925
rect 2369 5880 2421 5925
rect 2421 5880 2423 5925
rect 2447 5880 2489 5925
rect 2489 5880 2503 5925
rect 2527 5880 2557 5925
rect 2557 5880 2573 5925
rect 2573 5880 2583 5925
rect 2607 5880 2625 5925
rect 2625 5880 2641 5925
rect 2641 5880 2663 5925
rect 2127 5809 2149 5855
rect 2149 5809 2165 5855
rect 2165 5809 2183 5855
rect 2207 5809 2217 5855
rect 2217 5809 2233 5855
rect 2233 5809 2263 5855
rect 2287 5809 2301 5855
rect 2301 5809 2343 5855
rect 2367 5809 2369 5855
rect 2369 5809 2421 5855
rect 2421 5809 2423 5855
rect 2447 5809 2489 5855
rect 2489 5809 2503 5855
rect 2527 5809 2557 5855
rect 2557 5809 2573 5855
rect 2573 5809 2583 5855
rect 2607 5809 2625 5855
rect 2625 5809 2641 5855
rect 2641 5809 2663 5855
rect 2127 5799 2183 5809
rect 2207 5799 2263 5809
rect 2287 5799 2343 5809
rect 2367 5799 2423 5809
rect 2447 5799 2503 5809
rect 2527 5799 2583 5809
rect 2607 5799 2663 5809
rect 2127 5745 2149 5774
rect 2149 5745 2165 5774
rect 2165 5745 2183 5774
rect 2207 5745 2217 5774
rect 2217 5745 2233 5774
rect 2233 5745 2263 5774
rect 2287 5745 2301 5774
rect 2301 5745 2343 5774
rect 2367 5745 2369 5774
rect 2369 5745 2421 5774
rect 2421 5745 2423 5774
rect 2447 5745 2489 5774
rect 2489 5745 2503 5774
rect 2527 5745 2557 5774
rect 2557 5745 2573 5774
rect 2573 5745 2583 5774
rect 2607 5745 2625 5774
rect 2625 5745 2641 5774
rect 2641 5745 2663 5774
rect 2127 5733 2183 5745
rect 2207 5733 2263 5745
rect 2287 5733 2343 5745
rect 2367 5733 2423 5745
rect 2447 5733 2503 5745
rect 2527 5733 2583 5745
rect 2607 5733 2663 5745
rect 2127 5718 2149 5733
rect 2149 5718 2165 5733
rect 2165 5718 2183 5733
rect 2207 5718 2217 5733
rect 2217 5718 2233 5733
rect 2233 5718 2263 5733
rect 2287 5718 2301 5733
rect 2301 5718 2343 5733
rect 2367 5718 2369 5733
rect 2369 5718 2421 5733
rect 2421 5718 2423 5733
rect 2447 5718 2489 5733
rect 2489 5718 2503 5733
rect 2527 5718 2557 5733
rect 2557 5718 2573 5733
rect 2573 5718 2583 5733
rect 2607 5718 2625 5733
rect 2625 5718 2641 5733
rect 2641 5718 2663 5733
rect 2127 5681 2149 5693
rect 2149 5681 2165 5693
rect 2165 5681 2183 5693
rect 2207 5681 2217 5693
rect 2217 5681 2233 5693
rect 2233 5681 2263 5693
rect 2287 5681 2301 5693
rect 2301 5681 2343 5693
rect 2367 5681 2369 5693
rect 2369 5681 2421 5693
rect 2421 5681 2423 5693
rect 2447 5681 2489 5693
rect 2489 5681 2503 5693
rect 2527 5681 2557 5693
rect 2557 5681 2573 5693
rect 2573 5681 2583 5693
rect 2607 5681 2625 5693
rect 2625 5681 2641 5693
rect 2641 5681 2663 5693
rect 2127 5669 2183 5681
rect 2207 5669 2263 5681
rect 2287 5669 2343 5681
rect 2367 5669 2423 5681
rect 2447 5669 2503 5681
rect 2527 5669 2583 5681
rect 2607 5669 2663 5681
rect 2127 5637 2149 5669
rect 2149 5637 2165 5669
rect 2165 5637 2183 5669
rect 2207 5637 2217 5669
rect 2217 5637 2233 5669
rect 2233 5637 2263 5669
rect 2287 5637 2301 5669
rect 2301 5637 2343 5669
rect 2367 5637 2369 5669
rect 2369 5637 2421 5669
rect 2421 5637 2423 5669
rect 2447 5637 2489 5669
rect 2489 5637 2503 5669
rect 2527 5637 2557 5669
rect 2557 5637 2573 5669
rect 2573 5637 2583 5669
rect 2607 5637 2625 5669
rect 2625 5637 2641 5669
rect 2641 5637 2663 5669
rect 2127 5605 2183 5612
rect 2207 5605 2263 5612
rect 2287 5605 2343 5612
rect 2367 5605 2423 5612
rect 2447 5605 2503 5612
rect 2527 5605 2583 5612
rect 2607 5605 2663 5612
rect 2127 5556 2149 5605
rect 2149 5556 2165 5605
rect 2165 5556 2183 5605
rect 2207 5556 2217 5605
rect 2217 5556 2233 5605
rect 2233 5556 2263 5605
rect 2287 5556 2301 5605
rect 2301 5556 2343 5605
rect 2367 5556 2369 5605
rect 2369 5556 2421 5605
rect 2421 5556 2423 5605
rect 2447 5556 2489 5605
rect 2489 5556 2503 5605
rect 2527 5556 2557 5605
rect 2557 5556 2573 5605
rect 2573 5556 2583 5605
rect 2607 5556 2625 5605
rect 2625 5556 2641 5605
rect 2641 5556 2663 5605
rect 2127 4385 2149 4434
rect 2149 4385 2165 4434
rect 2165 4385 2217 4434
rect 2217 4385 2233 4434
rect 2233 4385 2285 4434
rect 2285 4385 2301 4434
rect 2301 4385 2353 4434
rect 2353 4385 2369 4434
rect 2369 4385 2421 4434
rect 2421 4385 2437 4434
rect 2437 4385 2489 4434
rect 2489 4385 2505 4434
rect 2505 4385 2557 4434
rect 2557 4385 2573 4434
rect 2573 4385 2625 4434
rect 2625 4385 2641 4434
rect 2641 4385 2663 4434
rect 2127 4373 2663 4385
rect 2127 4321 2149 4373
rect 2149 4321 2165 4373
rect 2165 4321 2217 4373
rect 2217 4321 2233 4373
rect 2233 4321 2285 4373
rect 2285 4321 2301 4373
rect 2301 4321 2353 4373
rect 2353 4321 2369 4373
rect 2369 4321 2421 4373
rect 2421 4321 2437 4373
rect 2437 4321 2489 4373
rect 2489 4321 2505 4373
rect 2505 4321 2557 4373
rect 2557 4321 2573 4373
rect 2573 4321 2625 4373
rect 2625 4321 2641 4373
rect 2641 4321 2663 4373
rect 2127 4309 2663 4321
rect 2127 4257 2149 4309
rect 2149 4257 2165 4309
rect 2165 4257 2217 4309
rect 2217 4257 2233 4309
rect 2233 4257 2285 4309
rect 2285 4257 2301 4309
rect 2301 4257 2353 4309
rect 2353 4257 2369 4309
rect 2369 4257 2421 4309
rect 2421 4257 2437 4309
rect 2437 4257 2489 4309
rect 2489 4257 2505 4309
rect 2505 4257 2557 4309
rect 2557 4257 2573 4309
rect 2573 4257 2625 4309
rect 2625 4257 2641 4309
rect 2641 4257 2663 4309
rect 2127 4245 2663 4257
rect 2127 4193 2149 4245
rect 2149 4193 2165 4245
rect 2165 4193 2217 4245
rect 2217 4193 2233 4245
rect 2233 4193 2285 4245
rect 2285 4193 2301 4245
rect 2301 4193 2353 4245
rect 2353 4193 2369 4245
rect 2369 4193 2421 4245
rect 2421 4193 2437 4245
rect 2437 4193 2489 4245
rect 2489 4193 2505 4245
rect 2505 4193 2557 4245
rect 2557 4193 2573 4245
rect 2573 4193 2625 4245
rect 2625 4193 2641 4245
rect 2641 4193 2663 4245
rect 2127 4181 2663 4193
rect 2127 4129 2149 4181
rect 2149 4129 2165 4181
rect 2165 4129 2217 4181
rect 2217 4129 2233 4181
rect 2233 4129 2285 4181
rect 2285 4129 2301 4181
rect 2301 4129 2353 4181
rect 2353 4129 2369 4181
rect 2369 4129 2421 4181
rect 2421 4129 2437 4181
rect 2437 4129 2489 4181
rect 2489 4129 2505 4181
rect 2505 4129 2557 4181
rect 2557 4129 2573 4181
rect 2573 4129 2625 4181
rect 2625 4129 2641 4181
rect 2641 4129 2663 4181
rect 2127 4117 2663 4129
rect 2127 4065 2149 4117
rect 2149 4065 2165 4117
rect 2165 4065 2217 4117
rect 2217 4065 2233 4117
rect 2233 4065 2285 4117
rect 2285 4065 2301 4117
rect 2301 4065 2353 4117
rect 2353 4065 2369 4117
rect 2369 4065 2421 4117
rect 2421 4065 2437 4117
rect 2437 4065 2489 4117
rect 2489 4065 2505 4117
rect 2505 4065 2557 4117
rect 2557 4065 2573 4117
rect 2573 4065 2625 4117
rect 2625 4065 2641 4117
rect 2641 4065 2663 4117
rect 2127 4053 2663 4065
rect 2127 4001 2149 4053
rect 2149 4001 2165 4053
rect 2165 4001 2217 4053
rect 2217 4001 2233 4053
rect 2233 4001 2285 4053
rect 2285 4001 2301 4053
rect 2301 4001 2353 4053
rect 2353 4001 2369 4053
rect 2369 4001 2421 4053
rect 2421 4001 2437 4053
rect 2437 4001 2489 4053
rect 2489 4001 2505 4053
rect 2505 4001 2557 4053
rect 2557 4001 2573 4053
rect 2573 4001 2625 4053
rect 2625 4001 2641 4053
rect 2641 4001 2663 4053
rect 2127 3989 2663 4001
rect 2127 3978 2149 3989
rect 2149 3978 2165 3989
rect 2165 3978 2217 3989
rect 2217 3978 2233 3989
rect 2233 3978 2285 3989
rect 2285 3978 2301 3989
rect 2301 3978 2353 3989
rect 2353 3978 2369 3989
rect 2369 3978 2421 3989
rect 2421 3978 2437 3989
rect 2437 3978 2489 3989
rect 2489 3978 2505 3989
rect 2505 3978 2557 3989
rect 2557 3978 2573 3989
rect 2573 3978 2625 3989
rect 2625 3978 2641 3989
rect 2641 3978 2663 3989
rect 2127 3937 2149 3953
rect 2149 3937 2165 3953
rect 2165 3937 2183 3953
rect 2207 3937 2217 3953
rect 2217 3937 2233 3953
rect 2233 3937 2263 3953
rect 2287 3937 2301 3953
rect 2301 3937 2343 3953
rect 2367 3937 2369 3953
rect 2369 3937 2421 3953
rect 2421 3937 2423 3953
rect 2447 3937 2489 3953
rect 2489 3937 2503 3953
rect 2527 3937 2557 3953
rect 2557 3937 2573 3953
rect 2573 3937 2583 3953
rect 2607 3937 2625 3953
rect 2625 3937 2641 3953
rect 2641 3937 2663 3953
rect 2127 3925 2183 3937
rect 2207 3925 2263 3937
rect 2287 3925 2343 3937
rect 2367 3925 2423 3937
rect 2447 3925 2503 3937
rect 2527 3925 2583 3937
rect 2607 3925 2663 3937
rect 2127 3897 2149 3925
rect 2149 3897 2165 3925
rect 2165 3897 2183 3925
rect 2207 3897 2217 3925
rect 2217 3897 2233 3925
rect 2233 3897 2263 3925
rect 2287 3897 2301 3925
rect 2301 3897 2343 3925
rect 2367 3897 2369 3925
rect 2369 3897 2421 3925
rect 2421 3897 2423 3925
rect 2447 3897 2489 3925
rect 2489 3897 2503 3925
rect 2527 3897 2557 3925
rect 2557 3897 2573 3925
rect 2573 3897 2583 3925
rect 2607 3897 2625 3925
rect 2625 3897 2641 3925
rect 2641 3897 2663 3925
rect 2127 3861 2183 3872
rect 2207 3861 2263 3872
rect 2287 3861 2343 3872
rect 2367 3861 2423 3872
rect 2447 3861 2503 3872
rect 2527 3861 2583 3872
rect 2607 3861 2663 3872
rect 2127 3816 2149 3861
rect 2149 3816 2165 3861
rect 2165 3816 2183 3861
rect 2207 3816 2217 3861
rect 2217 3816 2233 3861
rect 2233 3816 2263 3861
rect 2287 3816 2301 3861
rect 2301 3816 2343 3861
rect 2367 3816 2369 3861
rect 2369 3816 2421 3861
rect 2421 3816 2423 3861
rect 2447 3816 2489 3861
rect 2489 3816 2503 3861
rect 2527 3816 2557 3861
rect 2557 3816 2573 3861
rect 2573 3816 2583 3861
rect 2607 3816 2625 3861
rect 2625 3816 2641 3861
rect 2641 3816 2663 3861
rect 2127 3745 2149 3791
rect 2149 3745 2165 3791
rect 2165 3745 2183 3791
rect 2207 3745 2217 3791
rect 2217 3745 2233 3791
rect 2233 3745 2263 3791
rect 2287 3745 2301 3791
rect 2301 3745 2343 3791
rect 2367 3745 2369 3791
rect 2369 3745 2421 3791
rect 2421 3745 2423 3791
rect 2447 3745 2489 3791
rect 2489 3745 2503 3791
rect 2527 3745 2557 3791
rect 2557 3745 2573 3791
rect 2573 3745 2583 3791
rect 2607 3745 2625 3791
rect 2625 3745 2641 3791
rect 2641 3745 2663 3791
rect 2127 3735 2183 3745
rect 2207 3735 2263 3745
rect 2287 3735 2343 3745
rect 2367 3735 2423 3745
rect 2447 3735 2503 3745
rect 2527 3735 2583 3745
rect 2607 3735 2663 3745
rect 2127 3681 2149 3710
rect 2149 3681 2165 3710
rect 2165 3681 2183 3710
rect 2207 3681 2217 3710
rect 2217 3681 2233 3710
rect 2233 3681 2263 3710
rect 2287 3681 2301 3710
rect 2301 3681 2343 3710
rect 2367 3681 2369 3710
rect 2369 3681 2421 3710
rect 2421 3681 2423 3710
rect 2447 3681 2489 3710
rect 2489 3681 2503 3710
rect 2527 3681 2557 3710
rect 2557 3681 2573 3710
rect 2573 3681 2583 3710
rect 2607 3681 2625 3710
rect 2625 3681 2641 3710
rect 2641 3681 2663 3710
rect 2127 3669 2183 3681
rect 2207 3669 2263 3681
rect 2287 3669 2343 3681
rect 2367 3669 2423 3681
rect 2447 3669 2503 3681
rect 2527 3669 2583 3681
rect 2607 3669 2663 3681
rect 2127 3654 2149 3669
rect 2149 3654 2165 3669
rect 2165 3654 2183 3669
rect 2207 3654 2217 3669
rect 2217 3654 2233 3669
rect 2233 3654 2263 3669
rect 2287 3654 2301 3669
rect 2301 3654 2343 3669
rect 2367 3654 2369 3669
rect 2369 3654 2421 3669
rect 2421 3654 2423 3669
rect 2447 3654 2489 3669
rect 2489 3654 2503 3669
rect 2527 3654 2557 3669
rect 2557 3654 2573 3669
rect 2573 3654 2583 3669
rect 2607 3654 2625 3669
rect 2625 3654 2641 3669
rect 2641 3654 2663 3669
rect 2127 3617 2149 3629
rect 2149 3617 2165 3629
rect 2165 3617 2183 3629
rect 2207 3617 2217 3629
rect 2217 3617 2233 3629
rect 2233 3617 2263 3629
rect 2287 3617 2301 3629
rect 2301 3617 2343 3629
rect 2367 3617 2369 3629
rect 2369 3617 2421 3629
rect 2421 3617 2423 3629
rect 2447 3617 2489 3629
rect 2489 3617 2503 3629
rect 2527 3617 2557 3629
rect 2557 3617 2573 3629
rect 2573 3617 2583 3629
rect 2607 3617 2625 3629
rect 2625 3617 2641 3629
rect 2641 3617 2663 3629
rect 2127 3605 2183 3617
rect 2207 3605 2263 3617
rect 2287 3605 2343 3617
rect 2367 3605 2423 3617
rect 2447 3605 2503 3617
rect 2527 3605 2583 3617
rect 2607 3605 2663 3617
rect 2127 3573 2149 3605
rect 2149 3573 2165 3605
rect 2165 3573 2183 3605
rect 2207 3573 2217 3605
rect 2217 3573 2233 3605
rect 2233 3573 2263 3605
rect 2287 3573 2301 3605
rect 2301 3573 2343 3605
rect 2367 3573 2369 3605
rect 2369 3573 2421 3605
rect 2421 3573 2423 3605
rect 2447 3573 2489 3605
rect 2489 3573 2503 3605
rect 2527 3573 2557 3605
rect 2557 3573 2573 3605
rect 2573 3573 2583 3605
rect 2607 3573 2625 3605
rect 2625 3573 2641 3605
rect 2641 3573 2663 3605
rect 2127 3541 2183 3548
rect 2207 3541 2263 3548
rect 2287 3541 2343 3548
rect 2367 3541 2423 3548
rect 2447 3541 2503 3548
rect 2527 3541 2583 3548
rect 2607 3541 2663 3548
rect 2127 3492 2149 3541
rect 2149 3492 2165 3541
rect 2165 3492 2183 3541
rect 2207 3492 2217 3541
rect 2217 3492 2233 3541
rect 2233 3492 2263 3541
rect 2287 3492 2301 3541
rect 2301 3492 2343 3541
rect 2367 3492 2369 3541
rect 2369 3492 2421 3541
rect 2421 3492 2423 3541
rect 2447 3492 2489 3541
rect 2489 3492 2503 3541
rect 2527 3492 2557 3541
rect 2557 3492 2573 3541
rect 2573 3492 2583 3541
rect 2607 3492 2625 3541
rect 2625 3492 2641 3541
rect 2641 3492 2663 3541
rect 2127 2191 2149 2240
rect 2149 2191 2165 2240
rect 2165 2191 2217 2240
rect 2217 2191 2233 2240
rect 2233 2191 2285 2240
rect 2285 2191 2301 2240
rect 2301 2191 2353 2240
rect 2353 2191 2369 2240
rect 2369 2191 2421 2240
rect 2421 2191 2437 2240
rect 2437 2191 2489 2240
rect 2489 2191 2505 2240
rect 2505 2191 2557 2240
rect 2557 2191 2573 2240
rect 2573 2191 2625 2240
rect 2625 2191 2641 2240
rect 2641 2191 2663 2240
rect 2127 2179 2663 2191
rect 2127 2127 2149 2179
rect 2149 2127 2165 2179
rect 2165 2127 2217 2179
rect 2217 2127 2233 2179
rect 2233 2127 2285 2179
rect 2285 2127 2301 2179
rect 2301 2127 2353 2179
rect 2353 2127 2369 2179
rect 2369 2127 2421 2179
rect 2421 2127 2437 2179
rect 2437 2127 2489 2179
rect 2489 2127 2505 2179
rect 2505 2127 2557 2179
rect 2557 2127 2573 2179
rect 2573 2127 2625 2179
rect 2625 2127 2641 2179
rect 2641 2127 2663 2179
rect 2127 2115 2663 2127
rect 2127 2063 2149 2115
rect 2149 2063 2165 2115
rect 2165 2063 2217 2115
rect 2217 2063 2233 2115
rect 2233 2063 2285 2115
rect 2285 2063 2301 2115
rect 2301 2063 2353 2115
rect 2353 2063 2369 2115
rect 2369 2063 2421 2115
rect 2421 2063 2437 2115
rect 2437 2063 2489 2115
rect 2489 2063 2505 2115
rect 2505 2063 2557 2115
rect 2557 2063 2573 2115
rect 2573 2063 2625 2115
rect 2625 2063 2641 2115
rect 2641 2063 2663 2115
rect 2127 2051 2663 2063
rect 2127 1999 2149 2051
rect 2149 1999 2165 2051
rect 2165 1999 2217 2051
rect 2217 1999 2233 2051
rect 2233 1999 2285 2051
rect 2285 1999 2301 2051
rect 2301 1999 2353 2051
rect 2353 1999 2369 2051
rect 2369 1999 2421 2051
rect 2421 1999 2437 2051
rect 2437 1999 2489 2051
rect 2489 1999 2505 2051
rect 2505 1999 2557 2051
rect 2557 1999 2573 2051
rect 2573 1999 2625 2051
rect 2625 1999 2641 2051
rect 2641 1999 2663 2051
rect 2127 1987 2663 1999
rect 2127 1935 2149 1987
rect 2149 1935 2165 1987
rect 2165 1935 2217 1987
rect 2217 1935 2233 1987
rect 2233 1935 2285 1987
rect 2285 1935 2301 1987
rect 2301 1935 2353 1987
rect 2353 1935 2369 1987
rect 2369 1935 2421 1987
rect 2421 1935 2437 1987
rect 2437 1935 2489 1987
rect 2489 1935 2505 1987
rect 2505 1935 2557 1987
rect 2557 1935 2573 1987
rect 2573 1935 2625 1987
rect 2625 1935 2641 1987
rect 2641 1935 2663 1987
rect 2127 1923 2663 1935
rect 2127 1871 2149 1923
rect 2149 1871 2165 1923
rect 2165 1871 2217 1923
rect 2217 1871 2233 1923
rect 2233 1871 2285 1923
rect 2285 1871 2301 1923
rect 2301 1871 2353 1923
rect 2353 1871 2369 1923
rect 2369 1871 2421 1923
rect 2421 1871 2437 1923
rect 2437 1871 2489 1923
rect 2489 1871 2505 1923
rect 2505 1871 2557 1923
rect 2557 1871 2573 1923
rect 2573 1871 2625 1923
rect 2625 1871 2641 1923
rect 2641 1871 2663 1923
rect 2127 1859 2663 1871
rect 2127 1807 2149 1859
rect 2149 1807 2165 1859
rect 2165 1807 2217 1859
rect 2217 1807 2233 1859
rect 2233 1807 2285 1859
rect 2285 1807 2301 1859
rect 2301 1807 2353 1859
rect 2353 1807 2369 1859
rect 2369 1807 2421 1859
rect 2421 1807 2437 1859
rect 2437 1807 2489 1859
rect 2489 1807 2505 1859
rect 2505 1807 2557 1859
rect 2557 1807 2573 1859
rect 2573 1807 2625 1859
rect 2625 1807 2641 1859
rect 2641 1807 2663 1859
rect 2127 1795 2663 1807
rect 2127 1784 2149 1795
rect 2149 1784 2165 1795
rect 2165 1784 2217 1795
rect 2217 1784 2233 1795
rect 2233 1784 2285 1795
rect 2285 1784 2301 1795
rect 2301 1784 2353 1795
rect 2353 1784 2369 1795
rect 2369 1784 2421 1795
rect 2421 1784 2437 1795
rect 2437 1784 2489 1795
rect 2489 1784 2505 1795
rect 2505 1784 2557 1795
rect 2557 1784 2573 1795
rect 2573 1784 2625 1795
rect 2625 1784 2641 1795
rect 2641 1784 2663 1795
rect 2127 1743 2149 1759
rect 2149 1743 2165 1759
rect 2165 1743 2183 1759
rect 2207 1743 2217 1759
rect 2217 1743 2233 1759
rect 2233 1743 2263 1759
rect 2287 1743 2301 1759
rect 2301 1743 2343 1759
rect 2367 1743 2369 1759
rect 2369 1743 2421 1759
rect 2421 1743 2423 1759
rect 2447 1743 2489 1759
rect 2489 1743 2503 1759
rect 2527 1743 2557 1759
rect 2557 1743 2573 1759
rect 2573 1743 2583 1759
rect 2607 1743 2625 1759
rect 2625 1743 2641 1759
rect 2641 1743 2663 1759
rect 2127 1731 2183 1743
rect 2207 1731 2263 1743
rect 2287 1731 2343 1743
rect 2367 1731 2423 1743
rect 2447 1731 2503 1743
rect 2527 1731 2583 1743
rect 2607 1731 2663 1743
rect 2127 1703 2149 1731
rect 2149 1703 2165 1731
rect 2165 1703 2183 1731
rect 2207 1703 2217 1731
rect 2217 1703 2233 1731
rect 2233 1703 2263 1731
rect 2287 1703 2301 1731
rect 2301 1703 2343 1731
rect 2367 1703 2369 1731
rect 2369 1703 2421 1731
rect 2421 1703 2423 1731
rect 2447 1703 2489 1731
rect 2489 1703 2503 1731
rect 2527 1703 2557 1731
rect 2557 1703 2573 1731
rect 2573 1703 2583 1731
rect 2607 1703 2625 1731
rect 2625 1703 2641 1731
rect 2641 1703 2663 1731
rect 2127 1667 2183 1678
rect 2207 1667 2263 1678
rect 2287 1667 2343 1678
rect 2367 1667 2423 1678
rect 2447 1667 2503 1678
rect 2527 1667 2583 1678
rect 2607 1667 2663 1678
rect 2127 1622 2149 1667
rect 2149 1622 2165 1667
rect 2165 1622 2183 1667
rect 2207 1622 2217 1667
rect 2217 1622 2233 1667
rect 2233 1622 2263 1667
rect 2287 1622 2301 1667
rect 2301 1622 2343 1667
rect 2367 1622 2369 1667
rect 2369 1622 2421 1667
rect 2421 1622 2423 1667
rect 2447 1622 2489 1667
rect 2489 1622 2503 1667
rect 2527 1622 2557 1667
rect 2557 1622 2573 1667
rect 2573 1622 2583 1667
rect 2607 1622 2625 1667
rect 2625 1622 2641 1667
rect 2641 1622 2663 1667
rect 2127 1551 2149 1597
rect 2149 1551 2165 1597
rect 2165 1551 2183 1597
rect 2207 1551 2217 1597
rect 2217 1551 2233 1597
rect 2233 1551 2263 1597
rect 2287 1551 2301 1597
rect 2301 1551 2343 1597
rect 2367 1551 2369 1597
rect 2369 1551 2421 1597
rect 2421 1551 2423 1597
rect 2447 1551 2489 1597
rect 2489 1551 2503 1597
rect 2527 1551 2557 1597
rect 2557 1551 2573 1597
rect 2573 1551 2583 1597
rect 2607 1551 2625 1597
rect 2625 1551 2641 1597
rect 2641 1551 2663 1597
rect 2127 1541 2183 1551
rect 2207 1541 2263 1551
rect 2287 1541 2343 1551
rect 2367 1541 2423 1551
rect 2447 1541 2503 1551
rect 2527 1541 2583 1551
rect 2607 1541 2663 1551
rect 2127 1487 2149 1516
rect 2149 1487 2165 1516
rect 2165 1487 2183 1516
rect 2207 1487 2217 1516
rect 2217 1487 2233 1516
rect 2233 1487 2263 1516
rect 2287 1487 2301 1516
rect 2301 1487 2343 1516
rect 2367 1487 2369 1516
rect 2369 1487 2421 1516
rect 2421 1487 2423 1516
rect 2447 1487 2489 1516
rect 2489 1487 2503 1516
rect 2527 1487 2557 1516
rect 2557 1487 2573 1516
rect 2573 1487 2583 1516
rect 2607 1487 2625 1516
rect 2625 1487 2641 1516
rect 2641 1487 2663 1516
rect 2127 1475 2183 1487
rect 2207 1475 2263 1487
rect 2287 1475 2343 1487
rect 2367 1475 2423 1487
rect 2447 1475 2503 1487
rect 2527 1475 2583 1487
rect 2607 1475 2663 1487
rect 2127 1460 2149 1475
rect 2149 1460 2165 1475
rect 2165 1460 2183 1475
rect 2207 1460 2217 1475
rect 2217 1460 2233 1475
rect 2233 1460 2263 1475
rect 2287 1460 2301 1475
rect 2301 1460 2343 1475
rect 2367 1460 2369 1475
rect 2369 1460 2421 1475
rect 2421 1460 2423 1475
rect 2447 1460 2489 1475
rect 2489 1460 2503 1475
rect 2527 1460 2557 1475
rect 2557 1460 2573 1475
rect 2573 1460 2583 1475
rect 2607 1460 2625 1475
rect 2625 1460 2641 1475
rect 2641 1460 2663 1475
rect 2127 1423 2149 1435
rect 2149 1423 2165 1435
rect 2165 1423 2183 1435
rect 2207 1423 2217 1435
rect 2217 1423 2233 1435
rect 2233 1423 2263 1435
rect 2287 1423 2301 1435
rect 2301 1423 2343 1435
rect 2367 1423 2369 1435
rect 2369 1423 2421 1435
rect 2421 1423 2423 1435
rect 2447 1423 2489 1435
rect 2489 1423 2503 1435
rect 2527 1423 2557 1435
rect 2557 1423 2573 1435
rect 2573 1423 2583 1435
rect 2607 1423 2625 1435
rect 2625 1423 2641 1435
rect 2641 1423 2663 1435
rect 2127 1411 2183 1423
rect 2207 1411 2263 1423
rect 2287 1411 2343 1423
rect 2367 1411 2423 1423
rect 2447 1411 2503 1423
rect 2527 1411 2583 1423
rect 2607 1411 2663 1423
rect 2127 1379 2149 1411
rect 2149 1379 2165 1411
rect 2165 1379 2183 1411
rect 2207 1379 2217 1411
rect 2217 1379 2233 1411
rect 2233 1379 2263 1411
rect 2287 1379 2301 1411
rect 2301 1379 2343 1411
rect 2367 1379 2369 1411
rect 2369 1379 2421 1411
rect 2421 1379 2423 1411
rect 2447 1379 2489 1411
rect 2489 1379 2503 1411
rect 2527 1379 2557 1411
rect 2557 1379 2573 1411
rect 2573 1379 2583 1411
rect 2607 1379 2625 1411
rect 2625 1379 2641 1411
rect 2641 1379 2663 1411
rect 2127 1347 2183 1354
rect 2207 1347 2263 1354
rect 2287 1347 2343 1354
rect 2367 1347 2423 1354
rect 2447 1347 2503 1354
rect 2527 1347 2583 1354
rect 2607 1347 2663 1354
rect 2127 1298 2149 1347
rect 2149 1298 2165 1347
rect 2165 1298 2183 1347
rect 2207 1298 2217 1347
rect 2217 1298 2233 1347
rect 2233 1298 2263 1347
rect 2287 1298 2301 1347
rect 2301 1298 2343 1347
rect 2367 1298 2369 1347
rect 2369 1298 2421 1347
rect 2421 1298 2423 1347
rect 2447 1298 2489 1347
rect 2489 1298 2503 1347
rect 2527 1298 2557 1347
rect 2557 1298 2573 1347
rect 2573 1298 2583 1347
rect 2607 1298 2625 1347
rect 2625 1298 2641 1347
rect 2641 1298 2663 1347
rect 2104 85 2160 141
rect 2192 85 2248 141
rect 2280 85 2336 141
rect 2368 85 2424 141
rect 2456 85 2512 141
rect 2543 85 2599 141
rect 2630 85 2686 141
rect 2104 5 2160 61
rect 2192 5 2248 61
rect 2280 5 2336 61
rect 2368 5 2424 61
rect 2456 5 2512 61
rect 2543 5 2599 61
rect 2630 5 2686 61
<< metal3 >>
rect 286 38420 3170 39714
rect 286 37964 727 38420
rect 1263 37964 2127 38420
rect 2663 37964 3170 38420
rect 286 37939 3170 37964
rect 286 37883 727 37939
rect 783 37883 807 37939
rect 863 37883 887 37939
rect 943 37883 967 37939
rect 1023 37883 1047 37939
rect 1103 37883 1127 37939
rect 1183 37883 1207 37939
rect 1263 37883 2127 37939
rect 2183 37883 2207 37939
rect 2263 37883 2287 37939
rect 2343 37883 2367 37939
rect 2423 37883 2447 37939
rect 2503 37883 2527 37939
rect 2583 37883 2607 37939
rect 2663 37883 3170 37939
rect 286 37858 3170 37883
rect 286 37802 727 37858
rect 783 37802 807 37858
rect 863 37802 887 37858
rect 943 37802 967 37858
rect 1023 37802 1047 37858
rect 1103 37802 1127 37858
rect 1183 37802 1207 37858
rect 1263 37802 2127 37858
rect 2183 37802 2207 37858
rect 2263 37802 2287 37858
rect 2343 37802 2367 37858
rect 2423 37802 2447 37858
rect 2503 37802 2527 37858
rect 2583 37802 2607 37858
rect 2663 37802 3170 37858
rect 286 37777 3170 37802
rect 286 37721 727 37777
rect 783 37721 807 37777
rect 863 37721 887 37777
rect 943 37721 967 37777
rect 1023 37721 1047 37777
rect 1103 37721 1127 37777
rect 1183 37721 1207 37777
rect 1263 37721 2127 37777
rect 2183 37721 2207 37777
rect 2263 37721 2287 37777
rect 2343 37721 2367 37777
rect 2423 37721 2447 37777
rect 2503 37721 2527 37777
rect 2583 37721 2607 37777
rect 2663 37721 3170 37777
rect 286 37696 3170 37721
rect 286 37640 727 37696
rect 783 37640 807 37696
rect 863 37640 887 37696
rect 943 37640 967 37696
rect 1023 37640 1047 37696
rect 1103 37640 1127 37696
rect 1183 37640 1207 37696
rect 1263 37640 2127 37696
rect 2183 37640 2207 37696
rect 2263 37640 2287 37696
rect 2343 37640 2367 37696
rect 2423 37640 2447 37696
rect 2503 37640 2527 37696
rect 2583 37640 2607 37696
rect 2663 37640 3170 37696
rect 286 37615 3170 37640
rect 286 37559 727 37615
rect 783 37559 807 37615
rect 863 37559 887 37615
rect 943 37559 967 37615
rect 1023 37559 1047 37615
rect 1103 37559 1127 37615
rect 1183 37559 1207 37615
rect 1263 37559 2127 37615
rect 2183 37559 2207 37615
rect 2263 37559 2287 37615
rect 2343 37559 2367 37615
rect 2423 37559 2447 37615
rect 2503 37559 2527 37615
rect 2583 37559 2607 37615
rect 2663 37559 3170 37615
rect 286 37534 3170 37559
rect 286 37478 727 37534
rect 783 37478 807 37534
rect 863 37478 887 37534
rect 943 37478 967 37534
rect 1023 37478 1047 37534
rect 1103 37478 1127 37534
rect 1183 37478 1207 37534
rect 1263 37478 2127 37534
rect 2183 37478 2207 37534
rect 2263 37478 2287 37534
rect 2343 37478 2367 37534
rect 2423 37478 2447 37534
rect 2503 37478 2527 37534
rect 2583 37478 2607 37534
rect 2663 37478 3170 37534
rect 286 36366 3170 37478
rect 286 35910 727 36366
rect 1263 35910 2127 36366
rect 2663 35910 3170 36366
rect 286 35885 3170 35910
rect 286 35829 727 35885
rect 783 35829 807 35885
rect 863 35829 887 35885
rect 943 35829 967 35885
rect 1023 35829 1047 35885
rect 1103 35829 1127 35885
rect 1183 35829 1207 35885
rect 1263 35829 2127 35885
rect 2183 35829 2207 35885
rect 2263 35829 2287 35885
rect 2343 35829 2367 35885
rect 2423 35829 2447 35885
rect 2503 35829 2527 35885
rect 2583 35829 2607 35885
rect 2663 35829 3170 35885
rect 286 35804 3170 35829
rect 286 35748 727 35804
rect 783 35748 807 35804
rect 863 35748 887 35804
rect 943 35748 967 35804
rect 1023 35748 1047 35804
rect 1103 35748 1127 35804
rect 1183 35748 1207 35804
rect 1263 35748 2127 35804
rect 2183 35748 2207 35804
rect 2263 35748 2287 35804
rect 2343 35748 2367 35804
rect 2423 35748 2447 35804
rect 2503 35748 2527 35804
rect 2583 35748 2607 35804
rect 2663 35748 3170 35804
rect 286 35723 3170 35748
rect 286 35667 727 35723
rect 783 35667 807 35723
rect 863 35667 887 35723
rect 943 35667 967 35723
rect 1023 35667 1047 35723
rect 1103 35667 1127 35723
rect 1183 35667 1207 35723
rect 1263 35667 2127 35723
rect 2183 35667 2207 35723
rect 2263 35667 2287 35723
rect 2343 35667 2367 35723
rect 2423 35667 2447 35723
rect 2503 35667 2527 35723
rect 2583 35667 2607 35723
rect 2663 35667 3170 35723
rect 286 35642 3170 35667
rect 286 35586 727 35642
rect 783 35586 807 35642
rect 863 35586 887 35642
rect 943 35586 967 35642
rect 1023 35586 1047 35642
rect 1103 35586 1127 35642
rect 1183 35586 1207 35642
rect 1263 35586 2127 35642
rect 2183 35586 2207 35642
rect 2263 35586 2287 35642
rect 2343 35586 2367 35642
rect 2423 35586 2447 35642
rect 2503 35586 2527 35642
rect 2583 35586 2607 35642
rect 2663 35586 3170 35642
rect 286 35561 3170 35586
rect 286 35505 727 35561
rect 783 35505 807 35561
rect 863 35505 887 35561
rect 943 35505 967 35561
rect 1023 35505 1047 35561
rect 1103 35505 1127 35561
rect 1183 35505 1207 35561
rect 1263 35505 2127 35561
rect 2183 35505 2207 35561
rect 2263 35505 2287 35561
rect 2343 35505 2367 35561
rect 2423 35505 2447 35561
rect 2503 35505 2527 35561
rect 2583 35505 2607 35561
rect 2663 35505 3170 35561
rect 286 35480 3170 35505
rect 286 35424 727 35480
rect 783 35424 807 35480
rect 863 35424 887 35480
rect 943 35424 967 35480
rect 1023 35424 1047 35480
rect 1103 35424 1127 35480
rect 1183 35424 1207 35480
rect 1263 35424 2127 35480
rect 2183 35424 2207 35480
rect 2263 35424 2287 35480
rect 2343 35424 2367 35480
rect 2423 35424 2447 35480
rect 2503 35424 2527 35480
rect 2583 35424 2607 35480
rect 2663 35424 3170 35480
rect 286 34147 3170 35424
rect 286 33691 727 34147
rect 1263 33691 2127 34147
rect 2663 33691 3170 34147
rect 286 33666 3170 33691
rect 286 33610 727 33666
rect 783 33610 807 33666
rect 863 33610 887 33666
rect 943 33610 967 33666
rect 1023 33610 1047 33666
rect 1103 33610 1127 33666
rect 1183 33610 1207 33666
rect 1263 33610 2127 33666
rect 2183 33610 2207 33666
rect 2263 33610 2287 33666
rect 2343 33610 2367 33666
rect 2423 33610 2447 33666
rect 2503 33610 2527 33666
rect 2583 33610 2607 33666
rect 2663 33610 3170 33666
rect 286 33585 3170 33610
rect 286 33529 727 33585
rect 783 33529 807 33585
rect 863 33529 887 33585
rect 943 33529 967 33585
rect 1023 33529 1047 33585
rect 1103 33529 1127 33585
rect 1183 33529 1207 33585
rect 1263 33529 2127 33585
rect 2183 33529 2207 33585
rect 2263 33529 2287 33585
rect 2343 33529 2367 33585
rect 2423 33529 2447 33585
rect 2503 33529 2527 33585
rect 2583 33529 2607 33585
rect 2663 33529 3170 33585
rect 286 33504 3170 33529
rect 286 33448 727 33504
rect 783 33448 807 33504
rect 863 33448 887 33504
rect 943 33448 967 33504
rect 1023 33448 1047 33504
rect 1103 33448 1127 33504
rect 1183 33448 1207 33504
rect 1263 33448 2127 33504
rect 2183 33448 2207 33504
rect 2263 33448 2287 33504
rect 2343 33448 2367 33504
rect 2423 33448 2447 33504
rect 2503 33448 2527 33504
rect 2583 33448 2607 33504
rect 2663 33448 3170 33504
rect 286 33423 3170 33448
rect 286 33367 727 33423
rect 783 33367 807 33423
rect 863 33367 887 33423
rect 943 33367 967 33423
rect 1023 33367 1047 33423
rect 1103 33367 1127 33423
rect 1183 33367 1207 33423
rect 1263 33367 2127 33423
rect 2183 33367 2207 33423
rect 2263 33367 2287 33423
rect 2343 33367 2367 33423
rect 2423 33367 2447 33423
rect 2503 33367 2527 33423
rect 2583 33367 2607 33423
rect 2663 33367 3170 33423
rect 286 33342 3170 33367
rect 286 33286 727 33342
rect 783 33286 807 33342
rect 863 33286 887 33342
rect 943 33286 967 33342
rect 1023 33286 1047 33342
rect 1103 33286 1127 33342
rect 1183 33286 1207 33342
rect 1263 33286 2127 33342
rect 2183 33286 2207 33342
rect 2263 33286 2287 33342
rect 2343 33286 2367 33342
rect 2423 33286 2447 33342
rect 2503 33286 2527 33342
rect 2583 33286 2607 33342
rect 2663 33286 3170 33342
rect 286 33261 3170 33286
rect 286 33205 727 33261
rect 783 33205 807 33261
rect 863 33205 887 33261
rect 943 33205 967 33261
rect 1023 33205 1047 33261
rect 1103 33205 1127 33261
rect 1183 33205 1207 33261
rect 1263 33205 2127 33261
rect 2183 33205 2207 33261
rect 2263 33205 2287 33261
rect 2343 33205 2367 33261
rect 2423 33205 2447 33261
rect 2503 33205 2527 33261
rect 2583 33205 2607 33261
rect 2663 33205 3170 33261
rect 286 32018 3170 33205
rect 286 31562 727 32018
rect 1263 31562 2127 32018
rect 2663 31562 3170 32018
rect 286 31537 3170 31562
rect 286 31481 727 31537
rect 783 31481 807 31537
rect 863 31481 887 31537
rect 943 31481 967 31537
rect 1023 31481 1047 31537
rect 1103 31481 1127 31537
rect 1183 31481 1207 31537
rect 1263 31481 2127 31537
rect 2183 31481 2207 31537
rect 2263 31481 2287 31537
rect 2343 31481 2367 31537
rect 2423 31481 2447 31537
rect 2503 31481 2527 31537
rect 2583 31481 2607 31537
rect 2663 31481 3170 31537
rect 286 31456 3170 31481
rect 286 31400 727 31456
rect 783 31400 807 31456
rect 863 31400 887 31456
rect 943 31400 967 31456
rect 1023 31400 1047 31456
rect 1103 31400 1127 31456
rect 1183 31400 1207 31456
rect 1263 31400 2127 31456
rect 2183 31400 2207 31456
rect 2263 31400 2287 31456
rect 2343 31400 2367 31456
rect 2423 31400 2447 31456
rect 2503 31400 2527 31456
rect 2583 31400 2607 31456
rect 2663 31400 3170 31456
rect 286 31375 3170 31400
rect 286 31319 727 31375
rect 783 31319 807 31375
rect 863 31319 887 31375
rect 943 31319 967 31375
rect 1023 31319 1047 31375
rect 1103 31319 1127 31375
rect 1183 31319 1207 31375
rect 1263 31319 2127 31375
rect 2183 31319 2207 31375
rect 2263 31319 2287 31375
rect 2343 31319 2367 31375
rect 2423 31319 2447 31375
rect 2503 31319 2527 31375
rect 2583 31319 2607 31375
rect 2663 31319 3170 31375
rect 286 31294 3170 31319
rect 286 31238 727 31294
rect 783 31238 807 31294
rect 863 31238 887 31294
rect 943 31238 967 31294
rect 1023 31238 1047 31294
rect 1103 31238 1127 31294
rect 1183 31238 1207 31294
rect 1263 31238 2127 31294
rect 2183 31238 2207 31294
rect 2263 31238 2287 31294
rect 2343 31238 2367 31294
rect 2423 31238 2447 31294
rect 2503 31238 2527 31294
rect 2583 31238 2607 31294
rect 2663 31238 3170 31294
rect 286 31213 3170 31238
rect 286 31157 727 31213
rect 783 31157 807 31213
rect 863 31157 887 31213
rect 943 31157 967 31213
rect 1023 31157 1047 31213
rect 1103 31157 1127 31213
rect 1183 31157 1207 31213
rect 1263 31157 2127 31213
rect 2183 31157 2207 31213
rect 2263 31157 2287 31213
rect 2343 31157 2367 31213
rect 2423 31157 2447 31213
rect 2503 31157 2527 31213
rect 2583 31157 2607 31213
rect 2663 31157 3170 31213
rect 286 31132 3170 31157
rect 286 31076 727 31132
rect 783 31076 807 31132
rect 863 31076 887 31132
rect 943 31076 967 31132
rect 1023 31076 1047 31132
rect 1103 31076 1127 31132
rect 1183 31076 1207 31132
rect 1263 31076 2127 31132
rect 2183 31076 2207 31132
rect 2263 31076 2287 31132
rect 2343 31076 2367 31132
rect 2423 31076 2447 31132
rect 2503 31076 2527 31132
rect 2583 31076 2607 31132
rect 2663 31076 3170 31132
rect 286 29869 3170 31076
rect 286 29413 727 29869
rect 1263 29413 2127 29869
rect 2663 29413 3170 29869
rect 286 29388 3170 29413
rect 286 29332 727 29388
rect 783 29332 807 29388
rect 863 29332 887 29388
rect 943 29332 967 29388
rect 1023 29332 1047 29388
rect 1103 29332 1127 29388
rect 1183 29332 1207 29388
rect 1263 29332 2127 29388
rect 2183 29332 2207 29388
rect 2263 29332 2287 29388
rect 2343 29332 2367 29388
rect 2423 29332 2447 29388
rect 2503 29332 2527 29388
rect 2583 29332 2607 29388
rect 2663 29332 3170 29388
rect 286 29307 3170 29332
rect 286 29251 727 29307
rect 783 29251 807 29307
rect 863 29251 887 29307
rect 943 29251 967 29307
rect 1023 29251 1047 29307
rect 1103 29251 1127 29307
rect 1183 29251 1207 29307
rect 1263 29251 2127 29307
rect 2183 29251 2207 29307
rect 2263 29251 2287 29307
rect 2343 29251 2367 29307
rect 2423 29251 2447 29307
rect 2503 29251 2527 29307
rect 2583 29251 2607 29307
rect 2663 29251 3170 29307
rect 286 29226 3170 29251
rect 286 29170 727 29226
rect 783 29170 807 29226
rect 863 29170 887 29226
rect 943 29170 967 29226
rect 1023 29170 1047 29226
rect 1103 29170 1127 29226
rect 1183 29170 1207 29226
rect 1263 29170 2127 29226
rect 2183 29170 2207 29226
rect 2263 29170 2287 29226
rect 2343 29170 2367 29226
rect 2423 29170 2447 29226
rect 2503 29170 2527 29226
rect 2583 29170 2607 29226
rect 2663 29170 3170 29226
rect 286 29145 3170 29170
rect 286 29089 727 29145
rect 783 29089 807 29145
rect 863 29089 887 29145
rect 943 29089 967 29145
rect 1023 29089 1047 29145
rect 1103 29089 1127 29145
rect 1183 29089 1207 29145
rect 1263 29089 2127 29145
rect 2183 29089 2207 29145
rect 2263 29089 2287 29145
rect 2343 29089 2367 29145
rect 2423 29089 2447 29145
rect 2503 29089 2527 29145
rect 2583 29089 2607 29145
rect 2663 29089 3170 29145
rect 286 29064 3170 29089
rect 286 29008 727 29064
rect 783 29008 807 29064
rect 863 29008 887 29064
rect 943 29008 967 29064
rect 1023 29008 1047 29064
rect 1103 29008 1127 29064
rect 1183 29008 1207 29064
rect 1263 29008 2127 29064
rect 2183 29008 2207 29064
rect 2263 29008 2287 29064
rect 2343 29008 2367 29064
rect 2423 29008 2447 29064
rect 2503 29008 2527 29064
rect 2583 29008 2607 29064
rect 2663 29008 3170 29064
rect 286 28983 3170 29008
rect 286 28927 727 28983
rect 783 28927 807 28983
rect 863 28927 887 28983
rect 943 28927 967 28983
rect 1023 28927 1047 28983
rect 1103 28927 1127 28983
rect 1183 28927 1207 28983
rect 1263 28927 2127 28983
rect 2183 28927 2207 28983
rect 2263 28927 2287 28983
rect 2343 28927 2367 28983
rect 2423 28927 2447 28983
rect 2503 28927 2527 28983
rect 2583 28927 2607 28983
rect 2663 28927 3170 28983
rect 286 27862 3170 28927
rect 286 27406 727 27862
rect 1263 27406 2127 27862
rect 2663 27406 3170 27862
rect 286 27381 3170 27406
rect 286 27325 727 27381
rect 783 27325 807 27381
rect 863 27325 887 27381
rect 943 27325 967 27381
rect 1023 27325 1047 27381
rect 1103 27325 1127 27381
rect 1183 27325 1207 27381
rect 1263 27325 2127 27381
rect 2183 27325 2207 27381
rect 2263 27325 2287 27381
rect 2343 27325 2367 27381
rect 2423 27325 2447 27381
rect 2503 27325 2527 27381
rect 2583 27325 2607 27381
rect 2663 27325 3170 27381
rect 286 27300 3170 27325
rect 286 27244 727 27300
rect 783 27244 807 27300
rect 863 27244 887 27300
rect 943 27244 967 27300
rect 1023 27244 1047 27300
rect 1103 27244 1127 27300
rect 1183 27244 1207 27300
rect 1263 27244 2127 27300
rect 2183 27244 2207 27300
rect 2263 27244 2287 27300
rect 2343 27244 2367 27300
rect 2423 27244 2447 27300
rect 2503 27244 2527 27300
rect 2583 27244 2607 27300
rect 2663 27244 3170 27300
rect 286 27219 3170 27244
rect 286 27163 727 27219
rect 783 27163 807 27219
rect 863 27163 887 27219
rect 943 27163 967 27219
rect 1023 27163 1047 27219
rect 1103 27163 1127 27219
rect 1183 27163 1207 27219
rect 1263 27163 2127 27219
rect 2183 27163 2207 27219
rect 2263 27163 2287 27219
rect 2343 27163 2367 27219
rect 2423 27163 2447 27219
rect 2503 27163 2527 27219
rect 2583 27163 2607 27219
rect 2663 27163 3170 27219
rect 286 27138 3170 27163
rect 286 27082 727 27138
rect 783 27082 807 27138
rect 863 27082 887 27138
rect 943 27082 967 27138
rect 1023 27082 1047 27138
rect 1103 27082 1127 27138
rect 1183 27082 1207 27138
rect 1263 27082 2127 27138
rect 2183 27082 2207 27138
rect 2263 27082 2287 27138
rect 2343 27082 2367 27138
rect 2423 27082 2447 27138
rect 2503 27082 2527 27138
rect 2583 27082 2607 27138
rect 2663 27082 3170 27138
rect 286 27057 3170 27082
rect 286 27001 727 27057
rect 783 27001 807 27057
rect 863 27001 887 27057
rect 943 27001 967 27057
rect 1023 27001 1047 27057
rect 1103 27001 1127 27057
rect 1183 27001 1207 27057
rect 1263 27001 2127 27057
rect 2183 27001 2207 27057
rect 2263 27001 2287 27057
rect 2343 27001 2367 27057
rect 2423 27001 2447 27057
rect 2503 27001 2527 27057
rect 2583 27001 2607 27057
rect 2663 27001 3170 27057
rect 286 26976 3170 27001
rect 286 26920 727 26976
rect 783 26920 807 26976
rect 863 26920 887 26976
rect 943 26920 967 26976
rect 1023 26920 1047 26976
rect 1103 26920 1127 26976
rect 1183 26920 1207 26976
rect 1263 26920 2127 26976
rect 2183 26920 2207 26976
rect 2263 26920 2287 26976
rect 2343 26920 2367 26976
rect 2423 26920 2447 26976
rect 2503 26920 2527 26976
rect 2583 26920 2607 26976
rect 2663 26920 3170 26976
rect 286 25676 3170 26920
rect 286 25220 727 25676
rect 1263 25220 2127 25676
rect 2663 25220 3170 25676
rect 286 25195 3170 25220
rect 286 25139 727 25195
rect 783 25139 807 25195
rect 863 25139 887 25195
rect 943 25139 967 25195
rect 1023 25139 1047 25195
rect 1103 25139 1127 25195
rect 1183 25139 1207 25195
rect 1263 25139 2127 25195
rect 2183 25139 2207 25195
rect 2263 25139 2287 25195
rect 2343 25139 2367 25195
rect 2423 25139 2447 25195
rect 2503 25139 2527 25195
rect 2583 25139 2607 25195
rect 2663 25139 3170 25195
rect 286 25114 3170 25139
rect 286 25058 727 25114
rect 783 25058 807 25114
rect 863 25058 887 25114
rect 943 25058 967 25114
rect 1023 25058 1047 25114
rect 1103 25058 1127 25114
rect 1183 25058 1207 25114
rect 1263 25058 2127 25114
rect 2183 25058 2207 25114
rect 2263 25058 2287 25114
rect 2343 25058 2367 25114
rect 2423 25058 2447 25114
rect 2503 25058 2527 25114
rect 2583 25058 2607 25114
rect 2663 25058 3170 25114
rect 286 25033 3170 25058
rect 286 24977 727 25033
rect 783 24977 807 25033
rect 863 24977 887 25033
rect 943 24977 967 25033
rect 1023 24977 1047 25033
rect 1103 24977 1127 25033
rect 1183 24977 1207 25033
rect 1263 24977 2127 25033
rect 2183 24977 2207 25033
rect 2263 24977 2287 25033
rect 2343 24977 2367 25033
rect 2423 24977 2447 25033
rect 2503 24977 2527 25033
rect 2583 24977 2607 25033
rect 2663 24977 3170 25033
rect 286 24952 3170 24977
rect 286 24896 727 24952
rect 783 24896 807 24952
rect 863 24896 887 24952
rect 943 24896 967 24952
rect 1023 24896 1047 24952
rect 1103 24896 1127 24952
rect 1183 24896 1207 24952
rect 1263 24896 2127 24952
rect 2183 24896 2207 24952
rect 2263 24896 2287 24952
rect 2343 24896 2367 24952
rect 2423 24896 2447 24952
rect 2503 24896 2527 24952
rect 2583 24896 2607 24952
rect 2663 24896 3170 24952
rect 286 24871 3170 24896
rect 286 24815 727 24871
rect 783 24815 807 24871
rect 863 24815 887 24871
rect 943 24815 967 24871
rect 1023 24815 1047 24871
rect 1103 24815 1127 24871
rect 1183 24815 1207 24871
rect 1263 24815 2127 24871
rect 2183 24815 2207 24871
rect 2263 24815 2287 24871
rect 2343 24815 2367 24871
rect 2423 24815 2447 24871
rect 2503 24815 2527 24871
rect 2583 24815 2607 24871
rect 2663 24815 3170 24871
rect 286 24790 3170 24815
rect 286 24734 727 24790
rect 783 24734 807 24790
rect 863 24734 887 24790
rect 943 24734 967 24790
rect 1023 24734 1047 24790
rect 1103 24734 1127 24790
rect 1183 24734 1207 24790
rect 1263 24734 2127 24790
rect 2183 24734 2207 24790
rect 2263 24734 2287 24790
rect 2343 24734 2367 24790
rect 2423 24734 2447 24790
rect 2503 24734 2527 24790
rect 2583 24734 2607 24790
rect 2663 24734 3170 24790
rect 286 23528 3170 24734
rect 286 23072 727 23528
rect 1263 23072 2127 23528
rect 2663 23072 3170 23528
rect 286 23047 3170 23072
rect 286 22991 727 23047
rect 783 22991 807 23047
rect 863 22991 887 23047
rect 943 22991 967 23047
rect 1023 22991 1047 23047
rect 1103 22991 1127 23047
rect 1183 22991 1207 23047
rect 1263 22991 2127 23047
rect 2183 22991 2207 23047
rect 2263 22991 2287 23047
rect 2343 22991 2367 23047
rect 2423 22991 2447 23047
rect 2503 22991 2527 23047
rect 2583 22991 2607 23047
rect 2663 22991 3170 23047
rect 286 22966 3170 22991
rect 286 22910 727 22966
rect 783 22910 807 22966
rect 863 22910 887 22966
rect 943 22910 967 22966
rect 1023 22910 1047 22966
rect 1103 22910 1127 22966
rect 1183 22910 1207 22966
rect 1263 22910 2127 22966
rect 2183 22910 2207 22966
rect 2263 22910 2287 22966
rect 2343 22910 2367 22966
rect 2423 22910 2447 22966
rect 2503 22910 2527 22966
rect 2583 22910 2607 22966
rect 2663 22910 3170 22966
rect 286 22885 3170 22910
rect 286 22829 727 22885
rect 783 22829 807 22885
rect 863 22829 887 22885
rect 943 22829 967 22885
rect 1023 22829 1047 22885
rect 1103 22829 1127 22885
rect 1183 22829 1207 22885
rect 1263 22829 2127 22885
rect 2183 22829 2207 22885
rect 2263 22829 2287 22885
rect 2343 22829 2367 22885
rect 2423 22829 2447 22885
rect 2503 22829 2527 22885
rect 2583 22829 2607 22885
rect 2663 22829 3170 22885
rect 286 22804 3170 22829
rect 286 22748 727 22804
rect 783 22748 807 22804
rect 863 22748 887 22804
rect 943 22748 967 22804
rect 1023 22748 1047 22804
rect 1103 22748 1127 22804
rect 1183 22748 1207 22804
rect 1263 22748 2127 22804
rect 2183 22748 2207 22804
rect 2263 22748 2287 22804
rect 2343 22748 2367 22804
rect 2423 22748 2447 22804
rect 2503 22748 2527 22804
rect 2583 22748 2607 22804
rect 2663 22748 3170 22804
rect 286 22723 3170 22748
rect 286 22667 727 22723
rect 783 22667 807 22723
rect 863 22667 887 22723
rect 943 22667 967 22723
rect 1023 22667 1047 22723
rect 1103 22667 1127 22723
rect 1183 22667 1207 22723
rect 1263 22667 2127 22723
rect 2183 22667 2207 22723
rect 2263 22667 2287 22723
rect 2343 22667 2367 22723
rect 2423 22667 2447 22723
rect 2503 22667 2527 22723
rect 2583 22667 2607 22723
rect 2663 22667 3170 22723
rect 286 22642 3170 22667
rect 286 22586 727 22642
rect 783 22586 807 22642
rect 863 22586 887 22642
rect 943 22586 967 22642
rect 1023 22586 1047 22642
rect 1103 22586 1127 22642
rect 1183 22586 1207 22642
rect 1263 22586 2127 22642
rect 2183 22586 2207 22642
rect 2263 22586 2287 22642
rect 2343 22586 2367 22642
rect 2423 22586 2447 22642
rect 2503 22586 2527 22642
rect 2583 22586 2607 22642
rect 2663 22586 3170 22642
rect 286 21358 3170 22586
rect 286 20902 727 21358
rect 1263 20902 2127 21358
rect 2663 20902 3170 21358
rect 286 20877 3170 20902
rect 286 20821 727 20877
rect 783 20821 807 20877
rect 863 20821 887 20877
rect 943 20821 967 20877
rect 1023 20821 1047 20877
rect 1103 20821 1127 20877
rect 1183 20821 1207 20877
rect 1263 20821 2127 20877
rect 2183 20821 2207 20877
rect 2263 20821 2287 20877
rect 2343 20821 2367 20877
rect 2423 20821 2447 20877
rect 2503 20821 2527 20877
rect 2583 20821 2607 20877
rect 2663 20821 3170 20877
rect 286 20796 3170 20821
rect 286 20740 727 20796
rect 783 20740 807 20796
rect 863 20740 887 20796
rect 943 20740 967 20796
rect 1023 20740 1047 20796
rect 1103 20740 1127 20796
rect 1183 20740 1207 20796
rect 1263 20740 2127 20796
rect 2183 20740 2207 20796
rect 2263 20740 2287 20796
rect 2343 20740 2367 20796
rect 2423 20740 2447 20796
rect 2503 20740 2527 20796
rect 2583 20740 2607 20796
rect 2663 20740 3170 20796
rect 286 20715 3170 20740
rect 286 20659 727 20715
rect 783 20659 807 20715
rect 863 20659 887 20715
rect 943 20659 967 20715
rect 1023 20659 1047 20715
rect 1103 20659 1127 20715
rect 1183 20659 1207 20715
rect 1263 20659 2127 20715
rect 2183 20659 2207 20715
rect 2263 20659 2287 20715
rect 2343 20659 2367 20715
rect 2423 20659 2447 20715
rect 2503 20659 2527 20715
rect 2583 20659 2607 20715
rect 2663 20659 3170 20715
rect 286 20634 3170 20659
rect 286 20578 727 20634
rect 783 20578 807 20634
rect 863 20578 887 20634
rect 943 20578 967 20634
rect 1023 20578 1047 20634
rect 1103 20578 1127 20634
rect 1183 20578 1207 20634
rect 1263 20578 2127 20634
rect 2183 20578 2207 20634
rect 2263 20578 2287 20634
rect 2343 20578 2367 20634
rect 2423 20578 2447 20634
rect 2503 20578 2527 20634
rect 2583 20578 2607 20634
rect 2663 20578 3170 20634
rect 286 20553 3170 20578
rect 286 20497 727 20553
rect 783 20497 807 20553
rect 863 20497 887 20553
rect 943 20497 967 20553
rect 1023 20497 1047 20553
rect 1103 20497 1127 20553
rect 1183 20497 1207 20553
rect 1263 20497 2127 20553
rect 2183 20497 2207 20553
rect 2263 20497 2287 20553
rect 2343 20497 2367 20553
rect 2423 20497 2447 20553
rect 2503 20497 2527 20553
rect 2583 20497 2607 20553
rect 2663 20497 3170 20553
rect 286 20472 3170 20497
rect 286 20416 727 20472
rect 783 20416 807 20472
rect 863 20416 887 20472
rect 943 20416 967 20472
rect 1023 20416 1047 20472
rect 1103 20416 1127 20472
rect 1183 20416 1207 20472
rect 1263 20416 2127 20472
rect 2183 20416 2207 20472
rect 2263 20416 2287 20472
rect 2343 20416 2367 20472
rect 2423 20416 2447 20472
rect 2503 20416 2527 20472
rect 2583 20416 2607 20472
rect 2663 20416 3170 20472
rect 286 19254 3170 20416
rect 286 18798 727 19254
rect 1263 18798 2127 19254
rect 2663 18798 3170 19254
rect 286 18773 3170 18798
rect 286 18717 727 18773
rect 783 18717 807 18773
rect 863 18717 887 18773
rect 943 18717 967 18773
rect 1023 18717 1047 18773
rect 1103 18717 1127 18773
rect 1183 18717 1207 18773
rect 1263 18717 2127 18773
rect 2183 18717 2207 18773
rect 2263 18717 2287 18773
rect 2343 18717 2367 18773
rect 2423 18717 2447 18773
rect 2503 18717 2527 18773
rect 2583 18717 2607 18773
rect 2663 18717 3170 18773
rect 286 18692 3170 18717
rect 286 18636 727 18692
rect 783 18636 807 18692
rect 863 18636 887 18692
rect 943 18636 967 18692
rect 1023 18636 1047 18692
rect 1103 18636 1127 18692
rect 1183 18636 1207 18692
rect 1263 18636 2127 18692
rect 2183 18636 2207 18692
rect 2263 18636 2287 18692
rect 2343 18636 2367 18692
rect 2423 18636 2447 18692
rect 2503 18636 2527 18692
rect 2583 18636 2607 18692
rect 2663 18636 3170 18692
rect 286 18611 3170 18636
rect 286 18555 727 18611
rect 783 18555 807 18611
rect 863 18555 887 18611
rect 943 18555 967 18611
rect 1023 18555 1047 18611
rect 1103 18555 1127 18611
rect 1183 18555 1207 18611
rect 1263 18555 2127 18611
rect 2183 18555 2207 18611
rect 2263 18555 2287 18611
rect 2343 18555 2367 18611
rect 2423 18555 2447 18611
rect 2503 18555 2527 18611
rect 2583 18555 2607 18611
rect 2663 18555 3170 18611
rect 286 18530 3170 18555
rect 286 18474 727 18530
rect 783 18474 807 18530
rect 863 18474 887 18530
rect 943 18474 967 18530
rect 1023 18474 1047 18530
rect 1103 18474 1127 18530
rect 1183 18474 1207 18530
rect 1263 18474 2127 18530
rect 2183 18474 2207 18530
rect 2263 18474 2287 18530
rect 2343 18474 2367 18530
rect 2423 18474 2447 18530
rect 2503 18474 2527 18530
rect 2583 18474 2607 18530
rect 2663 18474 3170 18530
rect 286 18449 3170 18474
rect 286 18393 727 18449
rect 783 18393 807 18449
rect 863 18393 887 18449
rect 943 18393 967 18449
rect 1023 18393 1047 18449
rect 1103 18393 1127 18449
rect 1183 18393 1207 18449
rect 1263 18393 2127 18449
rect 2183 18393 2207 18449
rect 2263 18393 2287 18449
rect 2343 18393 2367 18449
rect 2423 18393 2447 18449
rect 2503 18393 2527 18449
rect 2583 18393 2607 18449
rect 2663 18393 3170 18449
rect 286 18368 3170 18393
rect 286 18312 727 18368
rect 783 18312 807 18368
rect 863 18312 887 18368
rect 943 18312 967 18368
rect 1023 18312 1047 18368
rect 1103 18312 1127 18368
rect 1183 18312 1207 18368
rect 1263 18312 2127 18368
rect 2183 18312 2207 18368
rect 2263 18312 2287 18368
rect 2343 18312 2367 18368
rect 2423 18312 2447 18368
rect 2503 18312 2527 18368
rect 2583 18312 2607 18368
rect 2663 18312 3170 18368
rect 286 17143 3170 18312
rect 286 16687 727 17143
rect 1263 16687 2127 17143
rect 2663 16687 3170 17143
rect 286 16662 3170 16687
rect 286 16606 727 16662
rect 783 16606 807 16662
rect 863 16606 887 16662
rect 943 16606 967 16662
rect 1023 16606 1047 16662
rect 1103 16606 1127 16662
rect 1183 16606 1207 16662
rect 1263 16606 2127 16662
rect 2183 16606 2207 16662
rect 2263 16606 2287 16662
rect 2343 16606 2367 16662
rect 2423 16606 2447 16662
rect 2503 16606 2527 16662
rect 2583 16606 2607 16662
rect 2663 16606 3170 16662
rect 286 16581 3170 16606
rect 286 16525 727 16581
rect 783 16525 807 16581
rect 863 16525 887 16581
rect 943 16525 967 16581
rect 1023 16525 1047 16581
rect 1103 16525 1127 16581
rect 1183 16525 1207 16581
rect 1263 16525 2127 16581
rect 2183 16525 2207 16581
rect 2263 16525 2287 16581
rect 2343 16525 2367 16581
rect 2423 16525 2447 16581
rect 2503 16525 2527 16581
rect 2583 16525 2607 16581
rect 2663 16525 3170 16581
rect 286 16500 3170 16525
rect 286 16444 727 16500
rect 783 16444 807 16500
rect 863 16444 887 16500
rect 943 16444 967 16500
rect 1023 16444 1047 16500
rect 1103 16444 1127 16500
rect 1183 16444 1207 16500
rect 1263 16444 2127 16500
rect 2183 16444 2207 16500
rect 2263 16444 2287 16500
rect 2343 16444 2367 16500
rect 2423 16444 2447 16500
rect 2503 16444 2527 16500
rect 2583 16444 2607 16500
rect 2663 16444 3170 16500
rect 286 16419 3170 16444
rect 286 16363 727 16419
rect 783 16363 807 16419
rect 863 16363 887 16419
rect 943 16363 967 16419
rect 1023 16363 1047 16419
rect 1103 16363 1127 16419
rect 1183 16363 1207 16419
rect 1263 16363 2127 16419
rect 2183 16363 2207 16419
rect 2263 16363 2287 16419
rect 2343 16363 2367 16419
rect 2423 16363 2447 16419
rect 2503 16363 2527 16419
rect 2583 16363 2607 16419
rect 2663 16363 3170 16419
rect 286 16338 3170 16363
rect 286 16282 727 16338
rect 783 16282 807 16338
rect 863 16282 887 16338
rect 943 16282 967 16338
rect 1023 16282 1047 16338
rect 1103 16282 1127 16338
rect 1183 16282 1207 16338
rect 1263 16282 2127 16338
rect 2183 16282 2207 16338
rect 2263 16282 2287 16338
rect 2343 16282 2367 16338
rect 2423 16282 2447 16338
rect 2503 16282 2527 16338
rect 2583 16282 2607 16338
rect 2663 16282 3170 16338
rect 286 16257 3170 16282
rect 286 16201 727 16257
rect 783 16201 807 16257
rect 863 16201 887 16257
rect 943 16201 967 16257
rect 1023 16201 1047 16257
rect 1103 16201 1127 16257
rect 1183 16201 1207 16257
rect 1263 16201 2127 16257
rect 2183 16201 2207 16257
rect 2263 16201 2287 16257
rect 2343 16201 2367 16257
rect 2423 16201 2447 16257
rect 2503 16201 2527 16257
rect 2583 16201 2607 16257
rect 2663 16201 3170 16257
rect 286 15006 3170 16201
rect 286 14550 727 15006
rect 1263 14550 2127 15006
rect 2663 14550 3170 15006
rect 286 14525 3170 14550
rect 286 14469 727 14525
rect 783 14469 807 14525
rect 863 14469 887 14525
rect 943 14469 967 14525
rect 1023 14469 1047 14525
rect 1103 14469 1127 14525
rect 1183 14469 1207 14525
rect 1263 14469 2127 14525
rect 2183 14469 2207 14525
rect 2263 14469 2287 14525
rect 2343 14469 2367 14525
rect 2423 14469 2447 14525
rect 2503 14469 2527 14525
rect 2583 14469 2607 14525
rect 2663 14469 3170 14525
rect 286 14444 3170 14469
rect 286 14388 727 14444
rect 783 14388 807 14444
rect 863 14388 887 14444
rect 943 14388 967 14444
rect 1023 14388 1047 14444
rect 1103 14388 1127 14444
rect 1183 14388 1207 14444
rect 1263 14388 2127 14444
rect 2183 14388 2207 14444
rect 2263 14388 2287 14444
rect 2343 14388 2367 14444
rect 2423 14388 2447 14444
rect 2503 14388 2527 14444
rect 2583 14388 2607 14444
rect 2663 14388 3170 14444
rect 286 14363 3170 14388
rect 286 14307 727 14363
rect 783 14307 807 14363
rect 863 14307 887 14363
rect 943 14307 967 14363
rect 1023 14307 1047 14363
rect 1103 14307 1127 14363
rect 1183 14307 1207 14363
rect 1263 14307 2127 14363
rect 2183 14307 2207 14363
rect 2263 14307 2287 14363
rect 2343 14307 2367 14363
rect 2423 14307 2447 14363
rect 2503 14307 2527 14363
rect 2583 14307 2607 14363
rect 2663 14307 3170 14363
rect 286 14282 3170 14307
rect 286 14226 727 14282
rect 783 14226 807 14282
rect 863 14226 887 14282
rect 943 14226 967 14282
rect 1023 14226 1047 14282
rect 1103 14226 1127 14282
rect 1183 14226 1207 14282
rect 1263 14226 2127 14282
rect 2183 14226 2207 14282
rect 2263 14226 2287 14282
rect 2343 14226 2367 14282
rect 2423 14226 2447 14282
rect 2503 14226 2527 14282
rect 2583 14226 2607 14282
rect 2663 14226 3170 14282
rect 286 14201 3170 14226
rect 286 14145 727 14201
rect 783 14145 807 14201
rect 863 14145 887 14201
rect 943 14145 967 14201
rect 1023 14145 1047 14201
rect 1103 14145 1127 14201
rect 1183 14145 1207 14201
rect 1263 14145 2127 14201
rect 2183 14145 2207 14201
rect 2263 14145 2287 14201
rect 2343 14145 2367 14201
rect 2423 14145 2447 14201
rect 2503 14145 2527 14201
rect 2583 14145 2607 14201
rect 2663 14145 3170 14201
rect 286 14120 3170 14145
rect 286 14064 727 14120
rect 783 14064 807 14120
rect 863 14064 887 14120
rect 943 14064 967 14120
rect 1023 14064 1047 14120
rect 1103 14064 1127 14120
rect 1183 14064 1207 14120
rect 1263 14064 2127 14120
rect 2183 14064 2207 14120
rect 2263 14064 2287 14120
rect 2343 14064 2367 14120
rect 2423 14064 2447 14120
rect 2503 14064 2527 14120
rect 2583 14064 2607 14120
rect 2663 14064 3170 14120
rect 110 13701 176 13707
rect 110 13637 111 13701
rect 175 13637 176 13701
rect 110 13620 176 13637
rect 110 13556 111 13620
rect 175 13556 176 13620
rect 110 13539 176 13556
rect 110 13475 111 13539
rect 175 13475 176 13539
rect 110 13458 176 13475
rect 110 13394 111 13458
rect 175 13394 176 13458
rect 110 13377 176 13394
rect 110 13313 111 13377
rect 175 13313 176 13377
rect 110 13296 176 13313
rect 110 13232 111 13296
rect 175 13232 176 13296
rect 110 13215 176 13232
rect 110 13151 111 13215
rect 175 13151 176 13215
rect 110 13133 176 13151
rect 110 13069 111 13133
rect 175 13069 176 13133
rect 110 13051 176 13069
rect 110 12987 111 13051
rect 175 12987 176 13051
rect 110 12969 176 12987
rect 110 12905 111 12969
rect 175 12905 176 12969
rect 110 12887 176 12905
rect 110 12823 111 12887
rect 175 12823 176 12887
rect 110 12817 176 12823
rect 286 12904 3170 14064
rect 286 12448 727 12904
rect 1263 12448 2127 12904
rect 2663 12448 3170 12904
rect 3280 13701 3346 13707
rect 3280 13637 3281 13701
rect 3345 13637 3346 13701
rect 3280 13620 3346 13637
rect 3280 13556 3281 13620
rect 3345 13556 3346 13620
rect 3280 13539 3346 13556
rect 3280 13475 3281 13539
rect 3345 13475 3346 13539
rect 3280 13458 3346 13475
rect 3280 13394 3281 13458
rect 3345 13394 3346 13458
rect 3280 13377 3346 13394
rect 3280 13313 3281 13377
rect 3345 13313 3346 13377
rect 3280 13296 3346 13313
rect 3280 13232 3281 13296
rect 3345 13232 3346 13296
rect 3280 13215 3346 13232
rect 3280 13151 3281 13215
rect 3345 13151 3346 13215
rect 3280 13133 3346 13151
rect 3280 13069 3281 13133
rect 3345 13069 3346 13133
rect 3280 13051 3346 13069
rect 3280 12987 3281 13051
rect 3345 12987 3346 13051
rect 3280 12969 3346 12987
rect 3280 12905 3281 12969
rect 3345 12905 3346 12969
rect 3280 12887 3346 12905
rect 3280 12823 3281 12887
rect 3345 12823 3346 12887
rect 3280 12817 3346 12823
rect 286 12423 3170 12448
rect 286 12367 727 12423
rect 783 12367 807 12423
rect 863 12367 887 12423
rect 943 12367 967 12423
rect 1023 12367 1047 12423
rect 1103 12367 1127 12423
rect 1183 12367 1207 12423
rect 1263 12367 2127 12423
rect 2183 12367 2207 12423
rect 2263 12367 2287 12423
rect 2343 12367 2367 12423
rect 2423 12367 2447 12423
rect 2503 12367 2527 12423
rect 2583 12367 2607 12423
rect 2663 12367 3170 12423
rect 286 12342 3170 12367
rect 286 12286 727 12342
rect 783 12286 807 12342
rect 863 12286 887 12342
rect 943 12286 967 12342
rect 1023 12286 1047 12342
rect 1103 12286 1127 12342
rect 1183 12286 1207 12342
rect 1263 12286 2127 12342
rect 2183 12286 2207 12342
rect 2263 12286 2287 12342
rect 2343 12286 2367 12342
rect 2423 12286 2447 12342
rect 2503 12286 2527 12342
rect 2583 12286 2607 12342
rect 2663 12286 3170 12342
rect 286 12261 3170 12286
rect 286 12205 727 12261
rect 783 12205 807 12261
rect 863 12205 887 12261
rect 943 12205 967 12261
rect 1023 12205 1047 12261
rect 1103 12205 1127 12261
rect 1183 12205 1207 12261
rect 1263 12205 2127 12261
rect 2183 12205 2207 12261
rect 2263 12205 2287 12261
rect 2343 12205 2367 12261
rect 2423 12205 2447 12261
rect 2503 12205 2527 12261
rect 2583 12205 2607 12261
rect 2663 12205 3170 12261
rect 286 12180 3170 12205
rect 286 12124 727 12180
rect 783 12124 807 12180
rect 863 12124 887 12180
rect 943 12124 967 12180
rect 1023 12124 1047 12180
rect 1103 12124 1127 12180
rect 1183 12124 1207 12180
rect 1263 12124 2127 12180
rect 2183 12124 2207 12180
rect 2263 12124 2287 12180
rect 2343 12124 2367 12180
rect 2423 12124 2447 12180
rect 2503 12124 2527 12180
rect 2583 12124 2607 12180
rect 2663 12124 3170 12180
rect 286 12099 3170 12124
rect 286 12043 727 12099
rect 783 12043 807 12099
rect 863 12043 887 12099
rect 943 12043 967 12099
rect 1023 12043 1047 12099
rect 1103 12043 1127 12099
rect 1183 12043 1207 12099
rect 1263 12043 2127 12099
rect 2183 12043 2207 12099
rect 2263 12043 2287 12099
rect 2343 12043 2367 12099
rect 2423 12043 2447 12099
rect 2503 12043 2527 12099
rect 2583 12043 2607 12099
rect 2663 12043 3170 12099
rect 286 12018 3170 12043
rect 286 11962 727 12018
rect 783 11962 807 12018
rect 863 11962 887 12018
rect 943 11962 967 12018
rect 1023 11962 1047 12018
rect 1103 11962 1127 12018
rect 1183 11962 1207 12018
rect 1263 11962 2127 12018
rect 2183 11962 2207 12018
rect 2263 11962 2287 12018
rect 2343 11962 2367 12018
rect 2423 11962 2447 12018
rect 2503 11962 2527 12018
rect 2583 11962 2607 12018
rect 2663 11962 3170 12018
rect 286 10810 3170 11962
rect 286 10354 727 10810
rect 1263 10354 2127 10810
rect 2663 10354 3170 10810
rect 286 10329 3170 10354
rect 286 10273 727 10329
rect 783 10273 807 10329
rect 863 10273 887 10329
rect 943 10273 967 10329
rect 1023 10273 1047 10329
rect 1103 10273 1127 10329
rect 1183 10273 1207 10329
rect 1263 10273 2127 10329
rect 2183 10273 2207 10329
rect 2263 10273 2287 10329
rect 2343 10273 2367 10329
rect 2423 10273 2447 10329
rect 2503 10273 2527 10329
rect 2583 10273 2607 10329
rect 2663 10273 3170 10329
rect 286 10248 3170 10273
rect 286 10192 727 10248
rect 783 10192 807 10248
rect 863 10192 887 10248
rect 943 10192 967 10248
rect 1023 10192 1047 10248
rect 1103 10192 1127 10248
rect 1183 10192 1207 10248
rect 1263 10192 2127 10248
rect 2183 10192 2207 10248
rect 2263 10192 2287 10248
rect 2343 10192 2367 10248
rect 2423 10192 2447 10248
rect 2503 10192 2527 10248
rect 2583 10192 2607 10248
rect 2663 10192 3170 10248
rect 286 10167 3170 10192
rect 286 10111 727 10167
rect 783 10111 807 10167
rect 863 10111 887 10167
rect 943 10111 967 10167
rect 1023 10111 1047 10167
rect 1103 10111 1127 10167
rect 1183 10111 1207 10167
rect 1263 10111 2127 10167
rect 2183 10111 2207 10167
rect 2263 10111 2287 10167
rect 2343 10111 2367 10167
rect 2423 10111 2447 10167
rect 2503 10111 2527 10167
rect 2583 10111 2607 10167
rect 2663 10111 3170 10167
rect 286 10086 3170 10111
rect 286 10030 727 10086
rect 783 10030 807 10086
rect 863 10030 887 10086
rect 943 10030 967 10086
rect 1023 10030 1047 10086
rect 1103 10030 1127 10086
rect 1183 10030 1207 10086
rect 1263 10030 2127 10086
rect 2183 10030 2207 10086
rect 2263 10030 2287 10086
rect 2343 10030 2367 10086
rect 2423 10030 2447 10086
rect 2503 10030 2527 10086
rect 2583 10030 2607 10086
rect 2663 10030 3170 10086
rect 286 10005 3170 10030
rect 286 9949 727 10005
rect 783 9949 807 10005
rect 863 9949 887 10005
rect 943 9949 967 10005
rect 1023 9949 1047 10005
rect 1103 9949 1127 10005
rect 1183 9949 1207 10005
rect 1263 9949 2127 10005
rect 2183 9949 2207 10005
rect 2263 9949 2287 10005
rect 2343 9949 2367 10005
rect 2423 9949 2447 10005
rect 2503 9949 2527 10005
rect 2583 9949 2607 10005
rect 2663 9949 3170 10005
rect 286 9924 3170 9949
rect 286 9868 727 9924
rect 783 9868 807 9924
rect 863 9868 887 9924
rect 943 9868 967 9924
rect 1023 9868 1047 9924
rect 1103 9868 1127 9924
rect 1183 9868 1207 9924
rect 1263 9868 2127 9924
rect 2183 9868 2207 9924
rect 2263 9868 2287 9924
rect 2343 9868 2367 9924
rect 2423 9868 2447 9924
rect 2503 9868 2527 9924
rect 2583 9868 2607 9924
rect 2663 9868 3170 9924
rect 286 8608 3170 9868
rect 286 8152 727 8608
rect 1263 8152 2127 8608
rect 2663 8152 3170 8608
rect 286 8127 3170 8152
rect 286 8071 727 8127
rect 783 8071 807 8127
rect 863 8071 887 8127
rect 943 8071 967 8127
rect 1023 8071 1047 8127
rect 1103 8071 1127 8127
rect 1183 8071 1207 8127
rect 1263 8071 2127 8127
rect 2183 8071 2207 8127
rect 2263 8071 2287 8127
rect 2343 8071 2367 8127
rect 2423 8071 2447 8127
rect 2503 8071 2527 8127
rect 2583 8071 2607 8127
rect 2663 8071 3170 8127
rect 286 8046 3170 8071
rect 286 7990 727 8046
rect 783 7990 807 8046
rect 863 7990 887 8046
rect 943 7990 967 8046
rect 1023 7990 1047 8046
rect 1103 7990 1127 8046
rect 1183 7990 1207 8046
rect 1263 7990 2127 8046
rect 2183 7990 2207 8046
rect 2263 7990 2287 8046
rect 2343 7990 2367 8046
rect 2423 7990 2447 8046
rect 2503 7990 2527 8046
rect 2583 7990 2607 8046
rect 2663 7990 3170 8046
rect 286 7965 3170 7990
rect 286 7909 727 7965
rect 783 7909 807 7965
rect 863 7909 887 7965
rect 943 7909 967 7965
rect 1023 7909 1047 7965
rect 1103 7909 1127 7965
rect 1183 7909 1207 7965
rect 1263 7909 2127 7965
rect 2183 7909 2207 7965
rect 2263 7909 2287 7965
rect 2343 7909 2367 7965
rect 2423 7909 2447 7965
rect 2503 7909 2527 7965
rect 2583 7909 2607 7965
rect 2663 7909 3170 7965
rect 286 7884 3170 7909
rect 286 7828 727 7884
rect 783 7828 807 7884
rect 863 7828 887 7884
rect 943 7828 967 7884
rect 1023 7828 1047 7884
rect 1103 7828 1127 7884
rect 1183 7828 1207 7884
rect 1263 7828 2127 7884
rect 2183 7828 2207 7884
rect 2263 7828 2287 7884
rect 2343 7828 2367 7884
rect 2423 7828 2447 7884
rect 2503 7828 2527 7884
rect 2583 7828 2607 7884
rect 2663 7828 3170 7884
rect 286 7803 3170 7828
rect 286 7747 727 7803
rect 783 7747 807 7803
rect 863 7747 887 7803
rect 943 7747 967 7803
rect 1023 7747 1047 7803
rect 1103 7747 1127 7803
rect 1183 7747 1207 7803
rect 1263 7747 2127 7803
rect 2183 7747 2207 7803
rect 2263 7747 2287 7803
rect 2343 7747 2367 7803
rect 2423 7747 2447 7803
rect 2503 7747 2527 7803
rect 2583 7747 2607 7803
rect 2663 7747 3170 7803
rect 286 7722 3170 7747
rect 286 7666 727 7722
rect 783 7666 807 7722
rect 863 7666 887 7722
rect 943 7666 967 7722
rect 1023 7666 1047 7722
rect 1103 7666 1127 7722
rect 1183 7666 1207 7722
rect 1263 7666 2127 7722
rect 2183 7666 2207 7722
rect 2263 7666 2287 7722
rect 2343 7666 2367 7722
rect 2423 7666 2447 7722
rect 2503 7666 2527 7722
rect 2583 7666 2607 7722
rect 2663 7666 3170 7722
rect 286 6498 3170 7666
rect 286 6042 727 6498
rect 1263 6042 2127 6498
rect 2663 6042 3170 6498
rect 286 6017 3170 6042
rect 286 5961 727 6017
rect 783 5961 807 6017
rect 863 5961 887 6017
rect 943 5961 967 6017
rect 1023 5961 1047 6017
rect 1103 5961 1127 6017
rect 1183 5961 1207 6017
rect 1263 5961 2127 6017
rect 2183 5961 2207 6017
rect 2263 5961 2287 6017
rect 2343 5961 2367 6017
rect 2423 5961 2447 6017
rect 2503 5961 2527 6017
rect 2583 5961 2607 6017
rect 2663 5961 3170 6017
rect 286 5936 3170 5961
rect 286 5880 727 5936
rect 783 5880 807 5936
rect 863 5880 887 5936
rect 943 5880 967 5936
rect 1023 5880 1047 5936
rect 1103 5880 1127 5936
rect 1183 5880 1207 5936
rect 1263 5880 2127 5936
rect 2183 5880 2207 5936
rect 2263 5880 2287 5936
rect 2343 5880 2367 5936
rect 2423 5880 2447 5936
rect 2503 5880 2527 5936
rect 2583 5880 2607 5936
rect 2663 5880 3170 5936
rect 286 5855 3170 5880
rect 286 5799 727 5855
rect 783 5799 807 5855
rect 863 5799 887 5855
rect 943 5799 967 5855
rect 1023 5799 1047 5855
rect 1103 5799 1127 5855
rect 1183 5799 1207 5855
rect 1263 5799 2127 5855
rect 2183 5799 2207 5855
rect 2263 5799 2287 5855
rect 2343 5799 2367 5855
rect 2423 5799 2447 5855
rect 2503 5799 2527 5855
rect 2583 5799 2607 5855
rect 2663 5799 3170 5855
rect 286 5774 3170 5799
rect 286 5718 727 5774
rect 783 5718 807 5774
rect 863 5718 887 5774
rect 943 5718 967 5774
rect 1023 5718 1047 5774
rect 1103 5718 1127 5774
rect 1183 5718 1207 5774
rect 1263 5718 2127 5774
rect 2183 5718 2207 5774
rect 2263 5718 2287 5774
rect 2343 5718 2367 5774
rect 2423 5718 2447 5774
rect 2503 5718 2527 5774
rect 2583 5718 2607 5774
rect 2663 5718 3170 5774
rect 286 5693 3170 5718
rect 286 5637 727 5693
rect 783 5637 807 5693
rect 863 5637 887 5693
rect 943 5637 967 5693
rect 1023 5637 1047 5693
rect 1103 5637 1127 5693
rect 1183 5637 1207 5693
rect 1263 5637 2127 5693
rect 2183 5637 2207 5693
rect 2263 5637 2287 5693
rect 2343 5637 2367 5693
rect 2423 5637 2447 5693
rect 2503 5637 2527 5693
rect 2583 5637 2607 5693
rect 2663 5637 3170 5693
rect 286 5612 3170 5637
rect 286 5556 727 5612
rect 783 5556 807 5612
rect 863 5556 887 5612
rect 943 5556 967 5612
rect 1023 5556 1047 5612
rect 1103 5556 1127 5612
rect 1183 5556 1207 5612
rect 1263 5556 2127 5612
rect 2183 5556 2207 5612
rect 2263 5556 2287 5612
rect 2343 5556 2367 5612
rect 2423 5556 2447 5612
rect 2503 5556 2527 5612
rect 2583 5556 2607 5612
rect 2663 5556 3170 5612
rect 286 4434 3170 5556
rect 286 3978 727 4434
rect 1263 3978 2127 4434
rect 2663 3978 3170 4434
rect 286 3953 3170 3978
rect 286 3897 727 3953
rect 783 3897 807 3953
rect 863 3897 887 3953
rect 943 3897 967 3953
rect 1023 3897 1047 3953
rect 1103 3897 1127 3953
rect 1183 3897 1207 3953
rect 1263 3897 2127 3953
rect 2183 3897 2207 3953
rect 2263 3897 2287 3953
rect 2343 3897 2367 3953
rect 2423 3897 2447 3953
rect 2503 3897 2527 3953
rect 2583 3897 2607 3953
rect 2663 3897 3170 3953
rect 286 3872 3170 3897
rect 286 3816 727 3872
rect 783 3816 807 3872
rect 863 3816 887 3872
rect 943 3816 967 3872
rect 1023 3816 1047 3872
rect 1103 3816 1127 3872
rect 1183 3816 1207 3872
rect 1263 3816 2127 3872
rect 2183 3816 2207 3872
rect 2263 3816 2287 3872
rect 2343 3816 2367 3872
rect 2423 3816 2447 3872
rect 2503 3816 2527 3872
rect 2583 3816 2607 3872
rect 2663 3816 3170 3872
rect 286 3791 3170 3816
rect 286 3735 727 3791
rect 783 3735 807 3791
rect 863 3735 887 3791
rect 943 3735 967 3791
rect 1023 3735 1047 3791
rect 1103 3735 1127 3791
rect 1183 3735 1207 3791
rect 1263 3735 2127 3791
rect 2183 3735 2207 3791
rect 2263 3735 2287 3791
rect 2343 3735 2367 3791
rect 2423 3735 2447 3791
rect 2503 3735 2527 3791
rect 2583 3735 2607 3791
rect 2663 3735 3170 3791
rect 286 3710 3170 3735
rect 286 3654 727 3710
rect 783 3654 807 3710
rect 863 3654 887 3710
rect 943 3654 967 3710
rect 1023 3654 1047 3710
rect 1103 3654 1127 3710
rect 1183 3654 1207 3710
rect 1263 3654 2127 3710
rect 2183 3654 2207 3710
rect 2263 3654 2287 3710
rect 2343 3654 2367 3710
rect 2423 3654 2447 3710
rect 2503 3654 2527 3710
rect 2583 3654 2607 3710
rect 2663 3654 3170 3710
rect 286 3629 3170 3654
rect 286 3573 727 3629
rect 783 3573 807 3629
rect 863 3573 887 3629
rect 943 3573 967 3629
rect 1023 3573 1047 3629
rect 1103 3573 1127 3629
rect 1183 3573 1207 3629
rect 1263 3573 2127 3629
rect 2183 3573 2207 3629
rect 2263 3573 2287 3629
rect 2343 3573 2367 3629
rect 2423 3573 2447 3629
rect 2503 3573 2527 3629
rect 2583 3573 2607 3629
rect 2663 3573 3170 3629
rect 286 3548 3170 3573
rect 286 3492 727 3548
rect 783 3492 807 3548
rect 863 3492 887 3548
rect 943 3492 967 3548
rect 1023 3492 1047 3548
rect 1103 3492 1127 3548
rect 1183 3492 1207 3548
rect 1263 3492 2127 3548
rect 2183 3492 2207 3548
rect 2263 3492 2287 3548
rect 2343 3492 2367 3548
rect 2423 3492 2447 3548
rect 2503 3492 2527 3548
rect 2583 3492 2607 3548
rect 2663 3492 3170 3548
rect 286 2240 3170 3492
rect 286 1784 727 2240
rect 1263 1784 2127 2240
rect 2663 1784 3170 2240
rect 286 1759 3170 1784
rect 286 1703 727 1759
rect 783 1703 807 1759
rect 863 1703 887 1759
rect 943 1703 967 1759
rect 1023 1703 1047 1759
rect 1103 1703 1127 1759
rect 1183 1703 1207 1759
rect 1263 1703 2127 1759
rect 2183 1703 2207 1759
rect 2263 1703 2287 1759
rect 2343 1703 2367 1759
rect 2423 1703 2447 1759
rect 2503 1703 2527 1759
rect 2583 1703 2607 1759
rect 2663 1703 3170 1759
rect 286 1678 3170 1703
rect 286 1622 727 1678
rect 783 1622 807 1678
rect 863 1622 887 1678
rect 943 1622 967 1678
rect 1023 1622 1047 1678
rect 1103 1622 1127 1678
rect 1183 1622 1207 1678
rect 1263 1622 2127 1678
rect 2183 1622 2207 1678
rect 2263 1622 2287 1678
rect 2343 1622 2367 1678
rect 2423 1622 2447 1678
rect 2503 1622 2527 1678
rect 2583 1622 2607 1678
rect 2663 1622 3170 1678
rect 286 1597 3170 1622
rect 286 1541 727 1597
rect 783 1541 807 1597
rect 863 1541 887 1597
rect 943 1541 967 1597
rect 1023 1541 1047 1597
rect 1103 1541 1127 1597
rect 1183 1541 1207 1597
rect 1263 1541 2127 1597
rect 2183 1541 2207 1597
rect 2263 1541 2287 1597
rect 2343 1541 2367 1597
rect 2423 1541 2447 1597
rect 2503 1541 2527 1597
rect 2583 1541 2607 1597
rect 2663 1541 3170 1597
rect 286 1516 3170 1541
rect 286 1460 727 1516
rect 783 1460 807 1516
rect 863 1460 887 1516
rect 943 1460 967 1516
rect 1023 1460 1047 1516
rect 1103 1460 1127 1516
rect 1183 1460 1207 1516
rect 1263 1460 2127 1516
rect 2183 1460 2207 1516
rect 2263 1460 2287 1516
rect 2343 1460 2367 1516
rect 2423 1460 2447 1516
rect 2503 1460 2527 1516
rect 2583 1460 2607 1516
rect 2663 1460 3170 1516
rect 286 1435 3170 1460
rect 286 1379 727 1435
rect 783 1379 807 1435
rect 863 1379 887 1435
rect 943 1379 967 1435
rect 1023 1379 1047 1435
rect 1103 1379 1127 1435
rect 1183 1379 1207 1435
rect 1263 1379 2127 1435
rect 2183 1379 2207 1435
rect 2263 1379 2287 1435
rect 2343 1379 2367 1435
rect 2423 1379 2447 1435
rect 2503 1379 2527 1435
rect 2583 1379 2607 1435
rect 2663 1379 3170 1435
rect 286 1354 3170 1379
rect 286 1298 727 1354
rect 783 1298 807 1354
rect 863 1298 887 1354
rect 943 1298 967 1354
rect 1023 1298 1047 1354
rect 1103 1298 1127 1354
rect 1183 1298 1207 1354
rect 1263 1298 2127 1354
rect 2183 1298 2207 1354
rect 2263 1298 2287 1354
rect 2343 1298 2367 1354
rect 2423 1298 2447 1354
rect 2503 1298 2527 1354
rect 2583 1298 2607 1354
rect 2663 1298 3170 1354
rect 286 286 3170 1298
rect 695 141 1295 166
rect 695 85 704 141
rect 760 85 792 141
rect 848 85 880 141
rect 936 85 968 141
rect 1024 85 1056 141
rect 1112 85 1143 141
rect 1199 85 1230 141
rect 1286 85 1295 141
rect 695 61 1295 85
rect 695 5 704 61
rect 760 5 792 61
rect 848 5 880 61
rect 936 5 968 61
rect 1024 5 1056 61
rect 1112 5 1143 61
rect 1199 5 1230 61
rect 1286 5 1295 61
rect 695 0 1295 5
rect 1495 141 1895 166
rect 1495 85 1504 141
rect 1560 85 1585 141
rect 1641 85 1666 141
rect 1722 85 1747 141
rect 1495 61 1747 85
rect 1495 5 1504 61
rect 1560 5 1585 61
rect 1641 5 1666 61
rect 1722 5 1747 61
rect 1883 5 1895 141
rect 1495 0 1895 5
rect 2095 141 2695 166
rect 2095 85 2104 141
rect 2160 85 2192 141
rect 2248 85 2280 141
rect 2336 85 2368 141
rect 2424 85 2456 141
rect 2512 85 2543 141
rect 2599 85 2630 141
rect 2686 85 2695 141
rect 2095 61 2695 85
rect 2095 5 2104 61
rect 2160 5 2192 61
rect 2248 5 2280 61
rect 2336 5 2368 61
rect 2424 5 2456 61
rect 2512 5 2543 61
rect 2599 5 2630 61
rect 2686 5 2695 61
rect 2095 0 2695 5
<< via3 >>
rect 111 13698 175 13701
rect 111 13642 115 13698
rect 115 13642 171 13698
rect 171 13642 175 13698
rect 111 13637 175 13642
rect 111 13617 175 13620
rect 111 13561 115 13617
rect 115 13561 171 13617
rect 171 13561 175 13617
rect 111 13556 175 13561
rect 111 13536 175 13539
rect 111 13480 115 13536
rect 115 13480 171 13536
rect 171 13480 175 13536
rect 111 13475 175 13480
rect 111 13455 175 13458
rect 111 13399 115 13455
rect 115 13399 171 13455
rect 171 13399 175 13455
rect 111 13394 175 13399
rect 111 13374 175 13377
rect 111 13318 115 13374
rect 115 13318 171 13374
rect 171 13318 175 13374
rect 111 13313 175 13318
rect 111 13292 175 13296
rect 111 13236 115 13292
rect 115 13236 171 13292
rect 171 13236 175 13292
rect 111 13232 175 13236
rect 111 13210 175 13215
rect 111 13154 115 13210
rect 115 13154 171 13210
rect 171 13154 175 13210
rect 111 13151 175 13154
rect 111 13128 175 13133
rect 111 13072 115 13128
rect 115 13072 171 13128
rect 171 13072 175 13128
rect 111 13069 175 13072
rect 111 13046 175 13051
rect 111 12990 115 13046
rect 115 12990 171 13046
rect 171 12990 175 13046
rect 111 12987 175 12990
rect 111 12964 175 12969
rect 111 12908 115 12964
rect 115 12908 171 12964
rect 171 12908 175 12964
rect 111 12905 175 12908
rect 111 12882 175 12887
rect 111 12826 115 12882
rect 115 12826 171 12882
rect 171 12826 175 12882
rect 111 12823 175 12826
rect 3281 13698 3345 13701
rect 3281 13642 3285 13698
rect 3285 13642 3341 13698
rect 3341 13642 3345 13698
rect 3281 13637 3345 13642
rect 3281 13617 3345 13620
rect 3281 13561 3285 13617
rect 3285 13561 3341 13617
rect 3341 13561 3345 13617
rect 3281 13556 3345 13561
rect 3281 13536 3345 13539
rect 3281 13480 3285 13536
rect 3285 13480 3341 13536
rect 3341 13480 3345 13536
rect 3281 13475 3345 13480
rect 3281 13455 3345 13458
rect 3281 13399 3285 13455
rect 3285 13399 3341 13455
rect 3341 13399 3345 13455
rect 3281 13394 3345 13399
rect 3281 13374 3345 13377
rect 3281 13318 3285 13374
rect 3285 13318 3341 13374
rect 3341 13318 3345 13374
rect 3281 13313 3345 13318
rect 3281 13292 3345 13296
rect 3281 13236 3285 13292
rect 3285 13236 3341 13292
rect 3341 13236 3345 13292
rect 3281 13232 3345 13236
rect 3281 13210 3345 13215
rect 3281 13154 3285 13210
rect 3285 13154 3341 13210
rect 3341 13154 3345 13210
rect 3281 13151 3345 13154
rect 3281 13128 3345 13133
rect 3281 13072 3285 13128
rect 3285 13072 3341 13128
rect 3341 13072 3345 13128
rect 3281 13069 3345 13072
rect 3281 13046 3345 13051
rect 3281 12990 3285 13046
rect 3285 12990 3341 13046
rect 3341 12990 3345 13046
rect 3281 12987 3345 12990
rect 3281 12964 3345 12969
rect 3281 12908 3285 12964
rect 3285 12908 3341 12964
rect 3341 12908 3345 12964
rect 3281 12905 3345 12908
rect 3281 12882 3345 12887
rect 3281 12826 3285 12882
rect 3285 12826 3341 12882
rect 3341 12826 3345 12882
rect 3281 12823 3345 12826
<< metal4 >>
rect 0 39964 3456 40000
rect 0 39728 215 39964
rect 451 39728 536 39964
rect 772 39728 856 39964
rect 1092 39728 1176 39964
rect 1412 39728 1496 39964
rect 1732 39728 1816 39964
rect 2052 39728 2136 39964
rect 2372 39728 2456 39964
rect 2692 39728 2776 39964
rect 3012 39728 3456 39964
rect 0 39640 3456 39728
rect 0 39404 215 39640
rect 451 39404 536 39640
rect 772 39404 856 39640
rect 1092 39404 1176 39640
rect 1412 39404 1496 39640
rect 1732 39404 1816 39640
rect 2052 39404 2136 39640
rect 2372 39404 2456 39640
rect 2692 39404 2776 39640
rect 3012 39404 3456 39640
rect 0 39316 3456 39404
rect 0 39080 215 39316
rect 451 39080 536 39316
rect 772 39080 856 39316
rect 1092 39080 1176 39316
rect 1412 39080 1496 39316
rect 1732 39080 1816 39316
rect 2052 39080 2136 39316
rect 2372 39080 2456 39316
rect 2692 39080 2776 39316
rect 3012 39080 3456 39316
rect 0 38992 3456 39080
rect 0 38756 215 38992
rect 451 38756 536 38992
rect 772 38756 856 38992
rect 1092 38756 1176 38992
rect 1412 38756 1496 38992
rect 1732 38756 1816 38992
rect 2052 38756 2136 38992
rect 2372 38756 2456 38992
rect 2692 38756 2776 38992
rect 3012 38756 3456 38992
rect 0 38668 3456 38756
rect 0 38432 215 38668
rect 451 38432 536 38668
rect 772 38432 856 38668
rect 1092 38432 1176 38668
rect 1412 38432 1496 38668
rect 1732 38432 1816 38668
rect 2052 38432 2136 38668
rect 2372 38432 2456 38668
rect 2692 38432 2776 38668
rect 3012 38432 3456 38668
rect 0 38344 3456 38432
rect 0 38108 215 38344
rect 451 38108 536 38344
rect 772 38108 856 38344
rect 1092 38108 1176 38344
rect 1412 38108 1496 38344
rect 1732 38108 1816 38344
rect 2052 38108 2136 38344
rect 2372 38108 2456 38344
rect 2692 38108 2776 38344
rect 3012 38108 3456 38344
rect 0 38020 3456 38108
rect 0 37784 215 38020
rect 451 37784 536 38020
rect 772 37784 856 38020
rect 1092 37784 1176 38020
rect 1412 37784 1496 38020
rect 1732 37784 1816 38020
rect 2052 37784 2136 38020
rect 2372 37784 2456 38020
rect 2692 37784 2776 38020
rect 3012 37784 3456 38020
rect 0 37696 3456 37784
rect 0 37460 215 37696
rect 451 37460 536 37696
rect 772 37460 856 37696
rect 1092 37460 1176 37696
rect 1412 37460 1496 37696
rect 1732 37460 1816 37696
rect 2052 37460 2136 37696
rect 2372 37460 2456 37696
rect 2692 37460 2776 37696
rect 3012 37460 3456 37696
rect 0 37372 3456 37460
rect 0 37136 215 37372
rect 451 37136 536 37372
rect 772 37136 856 37372
rect 1092 37136 1176 37372
rect 1412 37136 1496 37372
rect 1732 37136 1816 37372
rect 2052 37136 2136 37372
rect 2372 37136 2456 37372
rect 2692 37136 2776 37372
rect 3012 37136 3456 37372
rect 0 37048 3456 37136
rect 0 36812 215 37048
rect 451 36812 536 37048
rect 772 36812 856 37048
rect 1092 36812 1176 37048
rect 1412 36812 1496 37048
rect 1732 36812 1816 37048
rect 2052 36812 2136 37048
rect 2372 36812 2456 37048
rect 2692 36812 2776 37048
rect 3012 36812 3456 37048
rect 0 36724 3456 36812
rect 0 36488 215 36724
rect 451 36488 536 36724
rect 772 36488 856 36724
rect 1092 36488 1176 36724
rect 1412 36488 1496 36724
rect 1732 36488 1816 36724
rect 2052 36488 2136 36724
rect 2372 36488 2456 36724
rect 2692 36488 2776 36724
rect 3012 36488 3456 36724
rect 0 36400 3456 36488
rect 0 36164 215 36400
rect 451 36164 536 36400
rect 772 36164 856 36400
rect 1092 36164 1176 36400
rect 1412 36164 1496 36400
rect 1732 36164 1816 36400
rect 2052 36164 2136 36400
rect 2372 36164 2456 36400
rect 2692 36164 2776 36400
rect 3012 36164 3456 36400
rect 0 36076 3456 36164
rect 0 35840 215 36076
rect 451 35840 536 36076
rect 772 35840 856 36076
rect 1092 35840 1176 36076
rect 1412 35840 1496 36076
rect 1732 35840 1816 36076
rect 2052 35840 2136 36076
rect 2372 35840 2456 36076
rect 2692 35840 2776 36076
rect 3012 35840 3456 36076
rect 0 35752 3456 35840
rect 0 35516 215 35752
rect 451 35516 536 35752
rect 772 35516 856 35752
rect 1092 35516 1176 35752
rect 1412 35516 1496 35752
rect 1732 35516 1816 35752
rect 2052 35516 2136 35752
rect 2372 35516 2456 35752
rect 2692 35516 2776 35752
rect 3012 35516 3456 35752
rect 0 35428 3456 35516
rect 0 35192 215 35428
rect 451 35192 536 35428
rect 772 35192 856 35428
rect 1092 35192 1176 35428
rect 1412 35192 1496 35428
rect 1732 35192 1816 35428
rect 2052 35192 2136 35428
rect 2372 35192 2456 35428
rect 2692 35192 2776 35428
rect 3012 35192 3456 35428
rect 0 35157 3456 35192
rect 0 18972 3456 19000
rect 0 18736 215 18972
rect 451 18736 536 18972
rect 772 18736 856 18972
rect 1092 18736 1176 18972
rect 1412 18736 1496 18972
rect 1732 18736 1816 18972
rect 2052 18736 2136 18972
rect 2372 18736 2456 18972
rect 2692 18736 2776 18972
rect 3012 18736 3456 18972
rect 0 18636 3456 18736
rect 0 18400 215 18636
rect 451 18400 536 18636
rect 772 18400 856 18636
rect 1092 18400 1176 18636
rect 1412 18400 1496 18636
rect 1732 18400 1816 18636
rect 2052 18400 2136 18636
rect 2372 18400 2456 18636
rect 2692 18400 2776 18636
rect 3012 18400 3456 18636
rect 0 18300 3456 18400
rect 0 18064 215 18300
rect 451 18064 536 18300
rect 772 18064 856 18300
rect 1092 18064 1176 18300
rect 1412 18064 1496 18300
rect 1732 18064 1816 18300
rect 2052 18064 2136 18300
rect 2372 18064 2456 18300
rect 2692 18064 2776 18300
rect 3012 18064 3456 18300
rect 0 17964 3456 18064
rect 0 17728 215 17964
rect 451 17728 536 17964
rect 772 17728 856 17964
rect 1092 17728 1176 17964
rect 1412 17728 1496 17964
rect 1732 17728 1816 17964
rect 2052 17728 2136 17964
rect 2372 17728 2456 17964
rect 2692 17728 2776 17964
rect 3012 17728 3456 17964
rect 0 17628 3456 17728
rect 0 17392 215 17628
rect 451 17392 536 17628
rect 772 17392 856 17628
rect 1092 17392 1176 17628
rect 1412 17392 1496 17628
rect 1732 17392 1816 17628
rect 2052 17392 2136 17628
rect 2372 17392 2456 17628
rect 2692 17392 2776 17628
rect 3012 17392 3456 17628
rect 0 17292 3456 17392
rect 0 17056 215 17292
rect 451 17056 536 17292
rect 772 17056 856 17292
rect 1092 17056 1176 17292
rect 1412 17056 1496 17292
rect 1732 17056 1816 17292
rect 2052 17056 2136 17292
rect 2372 17056 2456 17292
rect 2692 17056 2776 17292
rect 3012 17056 3456 17292
rect 0 16956 3456 17056
rect 0 16720 215 16956
rect 451 16720 536 16956
rect 772 16720 856 16956
rect 1092 16720 1176 16956
rect 1412 16720 1496 16956
rect 1732 16720 1816 16956
rect 2052 16720 2136 16956
rect 2372 16720 2456 16956
rect 2692 16720 2776 16956
rect 3012 16720 3456 16956
rect 0 16620 3456 16720
rect 0 16384 215 16620
rect 451 16384 536 16620
rect 772 16384 856 16620
rect 1092 16384 1176 16620
rect 1412 16384 1496 16620
rect 1732 16384 1816 16620
rect 2052 16384 2136 16620
rect 2372 16384 2456 16620
rect 2692 16384 2776 16620
rect 3012 16384 3456 16620
rect 0 16284 3456 16384
rect 0 16048 215 16284
rect 451 16048 536 16284
rect 772 16048 856 16284
rect 1092 16048 1176 16284
rect 1412 16048 1496 16284
rect 1732 16048 1816 16284
rect 2052 16048 2136 16284
rect 2372 16048 2456 16284
rect 2692 16048 2776 16284
rect 3012 16048 3456 16284
rect 0 15948 3456 16048
rect 0 15712 215 15948
rect 451 15712 536 15948
rect 772 15712 856 15948
rect 1092 15712 1176 15948
rect 1412 15712 1496 15948
rect 1732 15712 1816 15948
rect 2052 15712 2136 15948
rect 2372 15712 2456 15948
rect 2692 15712 2776 15948
rect 3012 15712 3456 15948
rect 0 15612 3456 15712
rect 0 15376 215 15612
rect 451 15376 536 15612
rect 772 15376 856 15612
rect 1092 15376 1176 15612
rect 1412 15376 1496 15612
rect 1732 15376 1816 15612
rect 2052 15376 2136 15612
rect 2372 15376 2456 15612
rect 2692 15376 2776 15612
rect 3012 15376 3456 15612
rect 0 15276 3456 15376
rect 0 15040 215 15276
rect 451 15040 536 15276
rect 772 15040 856 15276
rect 1092 15040 1176 15276
rect 1412 15040 1496 15276
rect 1732 15040 1816 15276
rect 2052 15040 2136 15276
rect 2372 15040 2456 15276
rect 2692 15040 2776 15276
rect 3012 15040 3456 15276
rect 0 14940 3456 15040
rect 0 14704 215 14940
rect 451 14704 536 14940
rect 772 14704 856 14940
rect 1092 14704 1176 14940
rect 1412 14704 1496 14940
rect 1732 14704 1816 14940
rect 2052 14704 2136 14940
rect 2372 14704 2456 14940
rect 2692 14704 2776 14940
rect 3012 14704 3456 14940
rect 0 14604 3456 14704
rect 0 14368 215 14604
rect 451 14368 536 14604
rect 772 14368 856 14604
rect 1092 14368 1176 14604
rect 1412 14368 1496 14604
rect 1732 14368 1816 14604
rect 2052 14368 2136 14604
rect 2372 14368 2456 14604
rect 2692 14368 2776 14604
rect 3012 14368 3456 14604
rect 0 14268 3456 14368
rect 0 14032 215 14268
rect 451 14032 536 14268
rect 772 14032 856 14268
rect 1092 14032 1176 14268
rect 1412 14032 1496 14268
rect 1732 14032 1816 14268
rect 2052 14032 2136 14268
rect 2372 14032 2456 14268
rect 2692 14032 2776 14268
rect 3012 14032 3456 14268
rect 0 14007 3456 14032
rect 0 13701 3456 13707
rect 0 13637 111 13701
rect 175 13663 3281 13701
rect 175 13637 216 13663
rect 0 13620 216 13637
rect 0 13556 111 13620
rect 175 13556 216 13620
rect 0 13539 216 13556
rect 0 13475 111 13539
rect 175 13475 216 13539
rect 0 13458 216 13475
rect 0 13394 111 13458
rect 175 13427 216 13458
rect 452 13427 537 13663
rect 773 13427 857 13663
rect 1093 13427 1177 13663
rect 1413 13427 1497 13663
rect 1733 13427 1817 13663
rect 2053 13427 2137 13663
rect 2373 13427 2457 13663
rect 2693 13427 2777 13663
rect 3013 13637 3281 13663
rect 3345 13637 3456 13701
rect 3013 13620 3456 13637
rect 3013 13556 3281 13620
rect 3345 13556 3456 13620
rect 3013 13539 3456 13556
rect 3013 13475 3281 13539
rect 3345 13475 3456 13539
rect 3013 13458 3456 13475
rect 3013 13427 3281 13458
rect 175 13394 3281 13427
rect 3345 13394 3456 13458
rect 0 13377 3456 13394
rect 0 13313 111 13377
rect 175 13313 3281 13377
rect 3345 13313 3456 13377
rect 0 13296 3456 13313
rect 0 13232 111 13296
rect 175 13232 3281 13296
rect 3345 13232 3456 13296
rect 0 13215 3456 13232
rect 0 13151 111 13215
rect 175 13151 3281 13215
rect 3345 13151 3456 13215
rect 0 13133 3456 13151
rect 0 13069 111 13133
rect 175 13097 3281 13133
rect 175 13069 216 13097
rect 0 13051 216 13069
rect 0 12987 111 13051
rect 175 12987 216 13051
rect 0 12969 216 12987
rect 0 12905 111 12969
rect 175 12905 216 12969
rect 0 12887 216 12905
rect 0 12823 111 12887
rect 175 12861 216 12887
rect 452 12861 537 13097
rect 773 12861 857 13097
rect 1093 12861 1177 13097
rect 1413 12861 1497 13097
rect 1733 12861 1817 13097
rect 2053 12861 2137 13097
rect 2373 12861 2457 13097
rect 2693 12861 2777 13097
rect 3013 13069 3281 13097
rect 3345 13069 3456 13133
rect 3013 13051 3456 13069
rect 3013 12987 3281 13051
rect 3345 12987 3456 13051
rect 3013 12969 3456 12987
rect 3013 12905 3281 12969
rect 3345 12905 3456 12969
rect 3013 12887 3456 12905
rect 3013 12861 3281 12887
rect 175 12823 3281 12861
rect 3345 12823 3456 12887
rect 0 12817 3456 12823
rect 0 12493 3456 12537
rect 0 12257 215 12493
rect 451 12257 536 12493
rect 772 12257 856 12493
rect 1092 12257 1176 12493
rect 1412 12257 1496 12493
rect 1732 12257 1816 12493
rect 2052 12257 2136 12493
rect 2372 12257 2456 12493
rect 2692 12257 2776 12493
rect 3012 12257 3456 12493
rect 0 11927 3456 12257
rect 0 11691 215 11927
rect 451 11691 536 11927
rect 772 11691 856 11927
rect 1092 11691 1176 11927
rect 1412 11691 1496 11927
rect 1732 11691 1816 11927
rect 2052 11691 2136 11927
rect 2372 11691 2456 11927
rect 2692 11691 2776 11927
rect 3012 11691 3456 11927
rect 0 11647 3456 11691
rect 0 11281 3456 11347
rect 0 10625 3456 11221
rect 0 10329 215 10565
rect 451 10329 536 10565
rect 772 10329 856 10565
rect 1092 10329 1176 10565
rect 1412 10329 1496 10565
rect 1732 10329 1816 10565
rect 2052 10329 2136 10565
rect 2372 10329 2456 10565
rect 2692 10329 2776 10565
rect 3012 10329 3456 10565
rect 0 9673 3456 10269
rect 0 9547 3456 9613
rect 0 9203 3456 9247
rect 0 8967 216 9203
rect 452 8967 537 9203
rect 773 8967 857 9203
rect 1093 8967 1177 9203
rect 1413 8967 1497 9203
rect 1733 8967 1817 9203
rect 2053 8967 2137 9203
rect 2373 8967 2457 9203
rect 2693 8967 2777 9203
rect 3013 8967 3456 9203
rect 0 8597 3456 8967
rect 0 8361 216 8597
rect 452 8361 537 8597
rect 773 8361 857 8597
rect 1093 8361 1177 8597
rect 1413 8361 1497 8597
rect 1733 8361 1817 8597
rect 2053 8361 2137 8597
rect 2373 8361 2457 8597
rect 2693 8361 2777 8597
rect 3013 8361 3456 8597
rect 0 8317 3456 8361
rect 0 7993 3456 8037
rect 0 7757 215 7993
rect 451 7757 536 7993
rect 772 7757 856 7993
rect 1092 7757 1176 7993
rect 1412 7757 1496 7993
rect 1732 7757 1816 7993
rect 2052 7757 2136 7993
rect 2372 7757 2456 7993
rect 2692 7757 2776 7993
rect 3012 7757 3456 7993
rect 0 7627 3456 7757
rect 0 7391 215 7627
rect 451 7391 536 7627
rect 772 7391 856 7627
rect 1092 7391 1176 7627
rect 1412 7391 1496 7627
rect 1732 7391 1816 7627
rect 2052 7391 2136 7627
rect 2372 7391 2456 7627
rect 2692 7391 2776 7627
rect 3012 7391 3456 7627
rect 0 7347 3456 7391
rect 0 7023 3456 7067
rect 0 6787 215 7023
rect 451 6787 536 7023
rect 772 6787 856 7023
rect 1092 6787 1176 7023
rect 1412 6787 1496 7023
rect 1732 6787 1816 7023
rect 2052 6787 2136 7023
rect 2372 6787 2456 7023
rect 2692 6787 2776 7023
rect 3012 6787 3456 7023
rect 0 6657 3456 6787
rect 0 6421 215 6657
rect 451 6421 536 6657
rect 772 6421 856 6657
rect 1092 6421 1176 6657
rect 1412 6421 1496 6657
rect 1732 6421 1816 6657
rect 2052 6421 2136 6657
rect 2372 6421 2456 6657
rect 2692 6421 2776 6657
rect 3012 6421 3456 6657
rect 0 6377 3456 6421
rect 0 6053 3456 6097
rect 0 5817 215 6053
rect 451 5817 536 6053
rect 772 5817 856 6053
rect 1092 5817 1176 6053
rect 1412 5817 1496 6053
rect 1732 5817 1816 6053
rect 2052 5817 2136 6053
rect 2372 5817 2456 6053
rect 2692 5817 2776 6053
rect 3012 5817 3456 6053
rect 0 5447 3456 5817
rect 0 5211 215 5447
rect 451 5211 536 5447
rect 772 5211 856 5447
rect 1092 5211 1176 5447
rect 1412 5211 1496 5447
rect 1732 5211 1816 5447
rect 2052 5211 2136 5447
rect 2372 5211 2456 5447
rect 2692 5211 2776 5447
rect 3012 5211 3456 5447
rect 0 5167 3456 5211
rect 0 4843 3456 4887
rect 0 4607 215 4843
rect 451 4607 536 4843
rect 772 4607 856 4843
rect 1092 4607 1176 4843
rect 1412 4607 1496 4843
rect 1732 4607 1816 4843
rect 2052 4607 2136 4843
rect 2372 4607 2456 4843
rect 2692 4607 2776 4843
rect 3012 4607 3456 4843
rect 0 4237 3456 4607
rect 0 4001 215 4237
rect 451 4001 536 4237
rect 772 4001 856 4237
rect 1092 4001 1176 4237
rect 1412 4001 1496 4237
rect 1732 4001 1816 4237
rect 2052 4001 2136 4237
rect 2372 4001 2456 4237
rect 2692 4001 2776 4237
rect 3012 4001 3456 4237
rect 0 3957 3456 4001
rect 0 3633 3456 3677
rect 0 3397 215 3633
rect 451 3397 536 3633
rect 772 3397 856 3633
rect 1092 3397 1176 3633
rect 1412 3397 1496 3633
rect 1732 3397 1816 3633
rect 2052 3397 2136 3633
rect 2372 3397 2456 3633
rect 2692 3397 2776 3633
rect 3012 3397 3456 3633
rect 0 3267 3456 3397
rect 0 3031 215 3267
rect 451 3031 536 3267
rect 772 3031 856 3267
rect 1092 3031 1176 3267
rect 1412 3031 1496 3267
rect 1732 3031 1816 3267
rect 2052 3031 2136 3267
rect 2372 3031 2456 3267
rect 2692 3031 2776 3267
rect 3012 3031 3456 3267
rect 0 2987 3456 3031
rect 0 2663 3456 2707
rect 0 2427 215 2663
rect 451 2427 536 2663
rect 772 2427 856 2663
rect 1092 2427 1176 2663
rect 1412 2427 1496 2663
rect 1732 2427 1816 2663
rect 2052 2427 2136 2663
rect 2372 2427 2456 2663
rect 2692 2427 2776 2663
rect 3012 2427 3456 2663
rect 0 2057 3456 2427
rect 0 1821 215 2057
rect 451 1821 536 2057
rect 772 1821 856 2057
rect 1092 1821 1176 2057
rect 1412 1821 1496 2057
rect 1732 1821 1816 2057
rect 2052 1821 2136 2057
rect 2372 1821 2456 2057
rect 2692 1821 2776 2057
rect 3012 1821 3456 2057
rect 0 1777 3456 1821
rect 0 1452 3456 1497
rect 0 1216 215 1452
rect 451 1216 536 1452
rect 772 1216 856 1452
rect 1092 1216 1176 1452
rect 1412 1216 1496 1452
rect 1732 1216 1816 1452
rect 2052 1216 2136 1452
rect 2372 1216 2456 1452
rect 2692 1216 2776 1452
rect 3012 1216 3456 1452
rect 0 1070 3456 1216
rect 0 834 215 1070
rect 451 834 536 1070
rect 772 834 856 1070
rect 1092 834 1176 1070
rect 1412 834 1496 1070
rect 1732 834 1816 1070
rect 2052 834 2136 1070
rect 2372 834 2456 1070
rect 2692 834 2776 1070
rect 3012 834 3456 1070
rect 0 688 3456 834
rect 0 452 215 688
rect 451 452 536 688
rect 772 452 856 688
rect 1092 452 1176 688
rect 1412 452 1496 688
rect 1732 452 1816 688
rect 2052 452 2136 688
rect 2372 452 2456 688
rect 2692 452 2776 688
rect 3012 452 3456 688
rect 0 407 3456 452
<< via4 >>
rect 215 39728 451 39964
rect 536 39728 772 39964
rect 856 39728 1092 39964
rect 1176 39728 1412 39964
rect 1496 39728 1732 39964
rect 1816 39728 2052 39964
rect 2136 39728 2372 39964
rect 2456 39728 2692 39964
rect 2776 39728 3012 39964
rect 215 39404 451 39640
rect 536 39404 772 39640
rect 856 39404 1092 39640
rect 1176 39404 1412 39640
rect 1496 39404 1732 39640
rect 1816 39404 2052 39640
rect 2136 39404 2372 39640
rect 2456 39404 2692 39640
rect 2776 39404 3012 39640
rect 215 39080 451 39316
rect 536 39080 772 39316
rect 856 39080 1092 39316
rect 1176 39080 1412 39316
rect 1496 39080 1732 39316
rect 1816 39080 2052 39316
rect 2136 39080 2372 39316
rect 2456 39080 2692 39316
rect 2776 39080 3012 39316
rect 215 38756 451 38992
rect 536 38756 772 38992
rect 856 38756 1092 38992
rect 1176 38756 1412 38992
rect 1496 38756 1732 38992
rect 1816 38756 2052 38992
rect 2136 38756 2372 38992
rect 2456 38756 2692 38992
rect 2776 38756 3012 38992
rect 215 38432 451 38668
rect 536 38432 772 38668
rect 856 38432 1092 38668
rect 1176 38432 1412 38668
rect 1496 38432 1732 38668
rect 1816 38432 2052 38668
rect 2136 38432 2372 38668
rect 2456 38432 2692 38668
rect 2776 38432 3012 38668
rect 215 38108 451 38344
rect 536 38108 772 38344
rect 856 38108 1092 38344
rect 1176 38108 1412 38344
rect 1496 38108 1732 38344
rect 1816 38108 2052 38344
rect 2136 38108 2372 38344
rect 2456 38108 2692 38344
rect 2776 38108 3012 38344
rect 215 37784 451 38020
rect 536 37784 772 38020
rect 856 37784 1092 38020
rect 1176 37784 1412 38020
rect 1496 37784 1732 38020
rect 1816 37784 2052 38020
rect 2136 37784 2372 38020
rect 2456 37784 2692 38020
rect 2776 37784 3012 38020
rect 215 37460 451 37696
rect 536 37460 772 37696
rect 856 37460 1092 37696
rect 1176 37460 1412 37696
rect 1496 37460 1732 37696
rect 1816 37460 2052 37696
rect 2136 37460 2372 37696
rect 2456 37460 2692 37696
rect 2776 37460 3012 37696
rect 215 37136 451 37372
rect 536 37136 772 37372
rect 856 37136 1092 37372
rect 1176 37136 1412 37372
rect 1496 37136 1732 37372
rect 1816 37136 2052 37372
rect 2136 37136 2372 37372
rect 2456 37136 2692 37372
rect 2776 37136 3012 37372
rect 215 36812 451 37048
rect 536 36812 772 37048
rect 856 36812 1092 37048
rect 1176 36812 1412 37048
rect 1496 36812 1732 37048
rect 1816 36812 2052 37048
rect 2136 36812 2372 37048
rect 2456 36812 2692 37048
rect 2776 36812 3012 37048
rect 215 36488 451 36724
rect 536 36488 772 36724
rect 856 36488 1092 36724
rect 1176 36488 1412 36724
rect 1496 36488 1732 36724
rect 1816 36488 2052 36724
rect 2136 36488 2372 36724
rect 2456 36488 2692 36724
rect 2776 36488 3012 36724
rect 215 36164 451 36400
rect 536 36164 772 36400
rect 856 36164 1092 36400
rect 1176 36164 1412 36400
rect 1496 36164 1732 36400
rect 1816 36164 2052 36400
rect 2136 36164 2372 36400
rect 2456 36164 2692 36400
rect 2776 36164 3012 36400
rect 215 35840 451 36076
rect 536 35840 772 36076
rect 856 35840 1092 36076
rect 1176 35840 1412 36076
rect 1496 35840 1732 36076
rect 1816 35840 2052 36076
rect 2136 35840 2372 36076
rect 2456 35840 2692 36076
rect 2776 35840 3012 36076
rect 215 35516 451 35752
rect 536 35516 772 35752
rect 856 35516 1092 35752
rect 1176 35516 1412 35752
rect 1496 35516 1732 35752
rect 1816 35516 2052 35752
rect 2136 35516 2372 35752
rect 2456 35516 2692 35752
rect 2776 35516 3012 35752
rect 215 35192 451 35428
rect 536 35192 772 35428
rect 856 35192 1092 35428
rect 1176 35192 1412 35428
rect 1496 35192 1732 35428
rect 1816 35192 2052 35428
rect 2136 35192 2372 35428
rect 2456 35192 2692 35428
rect 2776 35192 3012 35428
rect 215 18736 451 18972
rect 536 18736 772 18972
rect 856 18736 1092 18972
rect 1176 18736 1412 18972
rect 1496 18736 1732 18972
rect 1816 18736 2052 18972
rect 2136 18736 2372 18972
rect 2456 18736 2692 18972
rect 2776 18736 3012 18972
rect 215 18400 451 18636
rect 536 18400 772 18636
rect 856 18400 1092 18636
rect 1176 18400 1412 18636
rect 1496 18400 1732 18636
rect 1816 18400 2052 18636
rect 2136 18400 2372 18636
rect 2456 18400 2692 18636
rect 2776 18400 3012 18636
rect 215 18064 451 18300
rect 536 18064 772 18300
rect 856 18064 1092 18300
rect 1176 18064 1412 18300
rect 1496 18064 1732 18300
rect 1816 18064 2052 18300
rect 2136 18064 2372 18300
rect 2456 18064 2692 18300
rect 2776 18064 3012 18300
rect 215 17728 451 17964
rect 536 17728 772 17964
rect 856 17728 1092 17964
rect 1176 17728 1412 17964
rect 1496 17728 1732 17964
rect 1816 17728 2052 17964
rect 2136 17728 2372 17964
rect 2456 17728 2692 17964
rect 2776 17728 3012 17964
rect 215 17392 451 17628
rect 536 17392 772 17628
rect 856 17392 1092 17628
rect 1176 17392 1412 17628
rect 1496 17392 1732 17628
rect 1816 17392 2052 17628
rect 2136 17392 2372 17628
rect 2456 17392 2692 17628
rect 2776 17392 3012 17628
rect 215 17056 451 17292
rect 536 17056 772 17292
rect 856 17056 1092 17292
rect 1176 17056 1412 17292
rect 1496 17056 1732 17292
rect 1816 17056 2052 17292
rect 2136 17056 2372 17292
rect 2456 17056 2692 17292
rect 2776 17056 3012 17292
rect 215 16720 451 16956
rect 536 16720 772 16956
rect 856 16720 1092 16956
rect 1176 16720 1412 16956
rect 1496 16720 1732 16956
rect 1816 16720 2052 16956
rect 2136 16720 2372 16956
rect 2456 16720 2692 16956
rect 2776 16720 3012 16956
rect 215 16384 451 16620
rect 536 16384 772 16620
rect 856 16384 1092 16620
rect 1176 16384 1412 16620
rect 1496 16384 1732 16620
rect 1816 16384 2052 16620
rect 2136 16384 2372 16620
rect 2456 16384 2692 16620
rect 2776 16384 3012 16620
rect 215 16048 451 16284
rect 536 16048 772 16284
rect 856 16048 1092 16284
rect 1176 16048 1412 16284
rect 1496 16048 1732 16284
rect 1816 16048 2052 16284
rect 2136 16048 2372 16284
rect 2456 16048 2692 16284
rect 2776 16048 3012 16284
rect 215 15712 451 15948
rect 536 15712 772 15948
rect 856 15712 1092 15948
rect 1176 15712 1412 15948
rect 1496 15712 1732 15948
rect 1816 15712 2052 15948
rect 2136 15712 2372 15948
rect 2456 15712 2692 15948
rect 2776 15712 3012 15948
rect 215 15376 451 15612
rect 536 15376 772 15612
rect 856 15376 1092 15612
rect 1176 15376 1412 15612
rect 1496 15376 1732 15612
rect 1816 15376 2052 15612
rect 2136 15376 2372 15612
rect 2456 15376 2692 15612
rect 2776 15376 3012 15612
rect 215 15040 451 15276
rect 536 15040 772 15276
rect 856 15040 1092 15276
rect 1176 15040 1412 15276
rect 1496 15040 1732 15276
rect 1816 15040 2052 15276
rect 2136 15040 2372 15276
rect 2456 15040 2692 15276
rect 2776 15040 3012 15276
rect 215 14704 451 14940
rect 536 14704 772 14940
rect 856 14704 1092 14940
rect 1176 14704 1412 14940
rect 1496 14704 1732 14940
rect 1816 14704 2052 14940
rect 2136 14704 2372 14940
rect 2456 14704 2692 14940
rect 2776 14704 3012 14940
rect 215 14368 451 14604
rect 536 14368 772 14604
rect 856 14368 1092 14604
rect 1176 14368 1412 14604
rect 1496 14368 1732 14604
rect 1816 14368 2052 14604
rect 2136 14368 2372 14604
rect 2456 14368 2692 14604
rect 2776 14368 3012 14604
rect 215 14032 451 14268
rect 536 14032 772 14268
rect 856 14032 1092 14268
rect 1176 14032 1412 14268
rect 1496 14032 1732 14268
rect 1816 14032 2052 14268
rect 2136 14032 2372 14268
rect 2456 14032 2692 14268
rect 2776 14032 3012 14268
rect 216 13427 452 13663
rect 537 13427 773 13663
rect 857 13427 1093 13663
rect 1177 13427 1413 13663
rect 1497 13427 1733 13663
rect 1817 13427 2053 13663
rect 2137 13427 2373 13663
rect 2457 13427 2693 13663
rect 2777 13427 3013 13663
rect 216 12861 452 13097
rect 537 12861 773 13097
rect 857 12861 1093 13097
rect 1177 12861 1413 13097
rect 1497 12861 1733 13097
rect 1817 12861 2053 13097
rect 2137 12861 2373 13097
rect 2457 12861 2693 13097
rect 2777 12861 3013 13097
rect 215 12257 451 12493
rect 536 12257 772 12493
rect 856 12257 1092 12493
rect 1176 12257 1412 12493
rect 1496 12257 1732 12493
rect 1816 12257 2052 12493
rect 2136 12257 2372 12493
rect 2456 12257 2692 12493
rect 2776 12257 3012 12493
rect 215 11691 451 11927
rect 536 11691 772 11927
rect 856 11691 1092 11927
rect 1176 11691 1412 11927
rect 1496 11691 1732 11927
rect 1816 11691 2052 11927
rect 2136 11691 2372 11927
rect 2456 11691 2692 11927
rect 2776 11691 3012 11927
rect 215 10329 451 10565
rect 536 10329 772 10565
rect 856 10329 1092 10565
rect 1176 10329 1412 10565
rect 1496 10329 1732 10565
rect 1816 10329 2052 10565
rect 2136 10329 2372 10565
rect 2456 10329 2692 10565
rect 2776 10329 3012 10565
rect 216 8967 452 9203
rect 537 8967 773 9203
rect 857 8967 1093 9203
rect 1177 8967 1413 9203
rect 1497 8967 1733 9203
rect 1817 8967 2053 9203
rect 2137 8967 2373 9203
rect 2457 8967 2693 9203
rect 2777 8967 3013 9203
rect 216 8361 452 8597
rect 537 8361 773 8597
rect 857 8361 1093 8597
rect 1177 8361 1413 8597
rect 1497 8361 1733 8597
rect 1817 8361 2053 8597
rect 2137 8361 2373 8597
rect 2457 8361 2693 8597
rect 2777 8361 3013 8597
rect 215 7757 451 7993
rect 536 7757 772 7993
rect 856 7757 1092 7993
rect 1176 7757 1412 7993
rect 1496 7757 1732 7993
rect 1816 7757 2052 7993
rect 2136 7757 2372 7993
rect 2456 7757 2692 7993
rect 2776 7757 3012 7993
rect 215 7391 451 7627
rect 536 7391 772 7627
rect 856 7391 1092 7627
rect 1176 7391 1412 7627
rect 1496 7391 1732 7627
rect 1816 7391 2052 7627
rect 2136 7391 2372 7627
rect 2456 7391 2692 7627
rect 2776 7391 3012 7627
rect 215 6787 451 7023
rect 536 6787 772 7023
rect 856 6787 1092 7023
rect 1176 6787 1412 7023
rect 1496 6787 1732 7023
rect 1816 6787 2052 7023
rect 2136 6787 2372 7023
rect 2456 6787 2692 7023
rect 2776 6787 3012 7023
rect 215 6421 451 6657
rect 536 6421 772 6657
rect 856 6421 1092 6657
rect 1176 6421 1412 6657
rect 1496 6421 1732 6657
rect 1816 6421 2052 6657
rect 2136 6421 2372 6657
rect 2456 6421 2692 6657
rect 2776 6421 3012 6657
rect 215 5817 451 6053
rect 536 5817 772 6053
rect 856 5817 1092 6053
rect 1176 5817 1412 6053
rect 1496 5817 1732 6053
rect 1816 5817 2052 6053
rect 2136 5817 2372 6053
rect 2456 5817 2692 6053
rect 2776 5817 3012 6053
rect 215 5211 451 5447
rect 536 5211 772 5447
rect 856 5211 1092 5447
rect 1176 5211 1412 5447
rect 1496 5211 1732 5447
rect 1816 5211 2052 5447
rect 2136 5211 2372 5447
rect 2456 5211 2692 5447
rect 2776 5211 3012 5447
rect 215 4607 451 4843
rect 536 4607 772 4843
rect 856 4607 1092 4843
rect 1176 4607 1412 4843
rect 1496 4607 1732 4843
rect 1816 4607 2052 4843
rect 2136 4607 2372 4843
rect 2456 4607 2692 4843
rect 2776 4607 3012 4843
rect 215 4001 451 4237
rect 536 4001 772 4237
rect 856 4001 1092 4237
rect 1176 4001 1412 4237
rect 1496 4001 1732 4237
rect 1816 4001 2052 4237
rect 2136 4001 2372 4237
rect 2456 4001 2692 4237
rect 2776 4001 3012 4237
rect 215 3397 451 3633
rect 536 3397 772 3633
rect 856 3397 1092 3633
rect 1176 3397 1412 3633
rect 1496 3397 1732 3633
rect 1816 3397 2052 3633
rect 2136 3397 2372 3633
rect 2456 3397 2692 3633
rect 2776 3397 3012 3633
rect 215 3031 451 3267
rect 536 3031 772 3267
rect 856 3031 1092 3267
rect 1176 3031 1412 3267
rect 1496 3031 1732 3267
rect 1816 3031 2052 3267
rect 2136 3031 2372 3267
rect 2456 3031 2692 3267
rect 2776 3031 3012 3267
rect 215 2427 451 2663
rect 536 2427 772 2663
rect 856 2427 1092 2663
rect 1176 2427 1412 2663
rect 1496 2427 1732 2663
rect 1816 2427 2052 2663
rect 2136 2427 2372 2663
rect 2456 2427 2692 2663
rect 2776 2427 3012 2663
rect 215 1821 451 2057
rect 536 1821 772 2057
rect 856 1821 1092 2057
rect 1176 1821 1412 2057
rect 1496 1821 1732 2057
rect 1816 1821 2052 2057
rect 2136 1821 2372 2057
rect 2456 1821 2692 2057
rect 2776 1821 3012 2057
rect 215 1216 451 1452
rect 536 1216 772 1452
rect 856 1216 1092 1452
rect 1176 1216 1412 1452
rect 1496 1216 1732 1452
rect 1816 1216 2052 1452
rect 2136 1216 2372 1452
rect 2456 1216 2692 1452
rect 2776 1216 3012 1452
rect 215 834 451 1070
rect 536 834 772 1070
rect 856 834 1092 1070
rect 1176 834 1412 1070
rect 1496 834 1732 1070
rect 1816 834 2052 1070
rect 2136 834 2372 1070
rect 2456 834 2692 1070
rect 2776 834 3012 1070
rect 215 452 451 688
rect 536 452 772 688
rect 856 452 1092 688
rect 1176 452 1412 688
rect 1496 452 1732 688
rect 1816 452 2052 688
rect 2136 452 2372 688
rect 2456 452 2692 688
rect 2776 452 3012 688
<< metal5 >>
rect 0 39964 3456 40000
rect 0 39728 215 39964
rect 451 39728 536 39964
rect 772 39728 856 39964
rect 1092 39728 1176 39964
rect 1412 39728 1496 39964
rect 1732 39728 1816 39964
rect 2052 39728 2136 39964
rect 2372 39728 2456 39964
rect 2692 39728 2776 39964
rect 3012 39728 3456 39964
rect 0 39640 3456 39728
rect 0 39404 215 39640
rect 451 39404 536 39640
rect 772 39404 856 39640
rect 1092 39404 1176 39640
rect 1412 39404 1496 39640
rect 1732 39404 1816 39640
rect 2052 39404 2136 39640
rect 2372 39404 2456 39640
rect 2692 39404 2776 39640
rect 3012 39404 3456 39640
rect 0 39316 3456 39404
rect 0 39080 215 39316
rect 451 39080 536 39316
rect 772 39080 856 39316
rect 1092 39080 1176 39316
rect 1412 39080 1496 39316
rect 1732 39080 1816 39316
rect 2052 39080 2136 39316
rect 2372 39080 2456 39316
rect 2692 39080 2776 39316
rect 3012 39080 3456 39316
rect 0 38992 3456 39080
rect 0 38756 215 38992
rect 451 38756 536 38992
rect 772 38756 856 38992
rect 1092 38756 1176 38992
rect 1412 38756 1496 38992
rect 1732 38756 1816 38992
rect 2052 38756 2136 38992
rect 2372 38756 2456 38992
rect 2692 38756 2776 38992
rect 3012 38756 3456 38992
rect 0 38668 3456 38756
rect 0 38432 215 38668
rect 451 38432 536 38668
rect 772 38432 856 38668
rect 1092 38432 1176 38668
rect 1412 38432 1496 38668
rect 1732 38432 1816 38668
rect 2052 38432 2136 38668
rect 2372 38432 2456 38668
rect 2692 38432 2776 38668
rect 3012 38432 3456 38668
rect 0 38344 3456 38432
rect 0 38108 215 38344
rect 451 38108 536 38344
rect 772 38108 856 38344
rect 1092 38108 1176 38344
rect 1412 38108 1496 38344
rect 1732 38108 1816 38344
rect 2052 38108 2136 38344
rect 2372 38108 2456 38344
rect 2692 38108 2776 38344
rect 3012 38108 3456 38344
rect 0 38020 3456 38108
rect 0 37784 215 38020
rect 451 37784 536 38020
rect 772 37784 856 38020
rect 1092 37784 1176 38020
rect 1412 37784 1496 38020
rect 1732 37784 1816 38020
rect 2052 37784 2136 38020
rect 2372 37784 2456 38020
rect 2692 37784 2776 38020
rect 3012 37784 3456 38020
rect 0 37696 3456 37784
rect 0 37460 215 37696
rect 451 37460 536 37696
rect 772 37460 856 37696
rect 1092 37460 1176 37696
rect 1412 37460 1496 37696
rect 1732 37460 1816 37696
rect 2052 37460 2136 37696
rect 2372 37460 2456 37696
rect 2692 37460 2776 37696
rect 3012 37460 3456 37696
rect 0 37372 3456 37460
rect 0 37136 215 37372
rect 451 37136 536 37372
rect 772 37136 856 37372
rect 1092 37136 1176 37372
rect 1412 37136 1496 37372
rect 1732 37136 1816 37372
rect 2052 37136 2136 37372
rect 2372 37136 2456 37372
rect 2692 37136 2776 37372
rect 3012 37136 3456 37372
rect 0 37048 3456 37136
rect 0 36812 215 37048
rect 451 36812 536 37048
rect 772 36812 856 37048
rect 1092 36812 1176 37048
rect 1412 36812 1496 37048
rect 1732 36812 1816 37048
rect 2052 36812 2136 37048
rect 2372 36812 2456 37048
rect 2692 36812 2776 37048
rect 3012 36812 3456 37048
rect 0 36724 3456 36812
rect 0 36488 215 36724
rect 451 36488 536 36724
rect 772 36488 856 36724
rect 1092 36488 1176 36724
rect 1412 36488 1496 36724
rect 1732 36488 1816 36724
rect 2052 36488 2136 36724
rect 2372 36488 2456 36724
rect 2692 36488 2776 36724
rect 3012 36488 3456 36724
rect 0 36400 3456 36488
rect 0 36164 215 36400
rect 451 36164 536 36400
rect 772 36164 856 36400
rect 1092 36164 1176 36400
rect 1412 36164 1496 36400
rect 1732 36164 1816 36400
rect 2052 36164 2136 36400
rect 2372 36164 2456 36400
rect 2692 36164 2776 36400
rect 3012 36164 3456 36400
rect 0 36076 3456 36164
rect 0 35840 215 36076
rect 451 35840 536 36076
rect 772 35840 856 36076
rect 1092 35840 1176 36076
rect 1412 35840 1496 36076
rect 1732 35840 1816 36076
rect 2052 35840 2136 36076
rect 2372 35840 2456 36076
rect 2692 35840 2776 36076
rect 3012 35840 3456 36076
rect 0 35752 3456 35840
rect 0 35516 215 35752
rect 451 35516 536 35752
rect 772 35516 856 35752
rect 1092 35516 1176 35752
rect 1412 35516 1496 35752
rect 1732 35516 1816 35752
rect 2052 35516 2136 35752
rect 2372 35516 2456 35752
rect 2692 35516 2776 35752
rect 3012 35516 3456 35752
rect 0 35428 3456 35516
rect 0 35192 215 35428
rect 451 35192 536 35428
rect 772 35192 856 35428
rect 1092 35192 1176 35428
rect 1412 35192 1496 35428
rect 1732 35192 1816 35428
rect 2052 35192 2136 35428
rect 2372 35192 2456 35428
rect 2692 35192 2776 35428
rect 3012 35192 3456 35428
rect 0 35157 3456 35192
rect 0 18972 3456 18997
rect 0 18736 215 18972
rect 451 18736 536 18972
rect 772 18736 856 18972
rect 1092 18736 1176 18972
rect 1412 18736 1496 18972
rect 1732 18736 1816 18972
rect 2052 18736 2136 18972
rect 2372 18736 2456 18972
rect 2692 18736 2776 18972
rect 3012 18736 3456 18972
rect 0 18636 3456 18736
rect 0 18400 215 18636
rect 451 18400 536 18636
rect 772 18400 856 18636
rect 1092 18400 1176 18636
rect 1412 18400 1496 18636
rect 1732 18400 1816 18636
rect 2052 18400 2136 18636
rect 2372 18400 2456 18636
rect 2692 18400 2776 18636
rect 3012 18400 3456 18636
rect 0 18300 3456 18400
rect 0 18064 215 18300
rect 451 18064 536 18300
rect 772 18064 856 18300
rect 1092 18064 1176 18300
rect 1412 18064 1496 18300
rect 1732 18064 1816 18300
rect 2052 18064 2136 18300
rect 2372 18064 2456 18300
rect 2692 18064 2776 18300
rect 3012 18064 3456 18300
rect 0 17964 3456 18064
rect 0 17728 215 17964
rect 451 17728 536 17964
rect 772 17728 856 17964
rect 1092 17728 1176 17964
rect 1412 17728 1496 17964
rect 1732 17728 1816 17964
rect 2052 17728 2136 17964
rect 2372 17728 2456 17964
rect 2692 17728 2776 17964
rect 3012 17728 3456 17964
rect 0 17628 3456 17728
rect 0 17392 215 17628
rect 451 17392 536 17628
rect 772 17392 856 17628
rect 1092 17392 1176 17628
rect 1412 17392 1496 17628
rect 1732 17392 1816 17628
rect 2052 17392 2136 17628
rect 2372 17392 2456 17628
rect 2692 17392 2776 17628
rect 3012 17392 3456 17628
rect 0 17292 3456 17392
rect 0 17056 215 17292
rect 451 17056 536 17292
rect 772 17056 856 17292
rect 1092 17056 1176 17292
rect 1412 17056 1496 17292
rect 1732 17056 1816 17292
rect 2052 17056 2136 17292
rect 2372 17056 2456 17292
rect 2692 17056 2776 17292
rect 3012 17056 3456 17292
rect 0 16956 3456 17056
rect 0 16720 215 16956
rect 451 16720 536 16956
rect 772 16720 856 16956
rect 1092 16720 1176 16956
rect 1412 16720 1496 16956
rect 1732 16720 1816 16956
rect 2052 16720 2136 16956
rect 2372 16720 2456 16956
rect 2692 16720 2776 16956
rect 3012 16720 3456 16956
rect 0 16620 3456 16720
rect 0 16384 215 16620
rect 451 16384 536 16620
rect 772 16384 856 16620
rect 1092 16384 1176 16620
rect 1412 16384 1496 16620
rect 1732 16384 1816 16620
rect 2052 16384 2136 16620
rect 2372 16384 2456 16620
rect 2692 16384 2776 16620
rect 3012 16384 3456 16620
rect 0 16284 3456 16384
rect 0 16048 215 16284
rect 451 16048 536 16284
rect 772 16048 856 16284
rect 1092 16048 1176 16284
rect 1412 16048 1496 16284
rect 1732 16048 1816 16284
rect 2052 16048 2136 16284
rect 2372 16048 2456 16284
rect 2692 16048 2776 16284
rect 3012 16048 3456 16284
rect 0 15948 3456 16048
rect 0 15712 215 15948
rect 451 15712 536 15948
rect 772 15712 856 15948
rect 1092 15712 1176 15948
rect 1412 15712 1496 15948
rect 1732 15712 1816 15948
rect 2052 15712 2136 15948
rect 2372 15712 2456 15948
rect 2692 15712 2776 15948
rect 3012 15712 3456 15948
rect 0 15612 3456 15712
rect 0 15376 215 15612
rect 451 15376 536 15612
rect 772 15376 856 15612
rect 1092 15376 1176 15612
rect 1412 15376 1496 15612
rect 1732 15376 1816 15612
rect 2052 15376 2136 15612
rect 2372 15376 2456 15612
rect 2692 15376 2776 15612
rect 3012 15376 3456 15612
rect 0 15276 3456 15376
rect 0 15040 215 15276
rect 451 15040 536 15276
rect 772 15040 856 15276
rect 1092 15040 1176 15276
rect 1412 15040 1496 15276
rect 1732 15040 1816 15276
rect 2052 15040 2136 15276
rect 2372 15040 2456 15276
rect 2692 15040 2776 15276
rect 3012 15040 3456 15276
rect 0 14940 3456 15040
rect 0 14704 215 14940
rect 451 14704 536 14940
rect 772 14704 856 14940
rect 1092 14704 1176 14940
rect 1412 14704 1496 14940
rect 1732 14704 1816 14940
rect 2052 14704 2136 14940
rect 2372 14704 2456 14940
rect 2692 14704 2776 14940
rect 3012 14704 3456 14940
rect 0 14604 3456 14704
rect 0 14368 215 14604
rect 451 14368 536 14604
rect 772 14368 856 14604
rect 1092 14368 1176 14604
rect 1412 14368 1496 14604
rect 1732 14368 1816 14604
rect 2052 14368 2136 14604
rect 2372 14368 2456 14604
rect 2692 14368 2776 14604
rect 3012 14368 3456 14604
rect 0 14268 3456 14368
rect 0 14032 215 14268
rect 451 14032 536 14268
rect 772 14032 856 14268
rect 1092 14032 1176 14268
rect 1412 14032 1496 14268
rect 1732 14032 1816 14268
rect 2052 14032 2136 14268
rect 2372 14032 2456 14268
rect 2692 14032 2776 14268
rect 3012 14032 3456 14268
rect 0 14007 3456 14032
rect 0 13663 3456 13687
rect 0 13427 216 13663
rect 452 13427 537 13663
rect 773 13427 857 13663
rect 1093 13427 1177 13663
rect 1413 13427 1497 13663
rect 1733 13427 1817 13663
rect 2053 13427 2137 13663
rect 2373 13427 2457 13663
rect 2693 13427 2777 13663
rect 3013 13427 3456 13663
rect 0 13097 3456 13427
rect 0 12861 216 13097
rect 452 12861 537 13097
rect 773 12861 857 13097
rect 1093 12861 1177 13097
rect 1413 12861 1497 13097
rect 1733 12861 1817 13097
rect 2053 12861 2137 13097
rect 2373 12861 2457 13097
rect 2693 12861 2777 13097
rect 3013 12861 3456 13097
rect 0 12837 3456 12861
rect 0 12493 3456 12517
rect 0 12257 215 12493
rect 451 12257 536 12493
rect 772 12257 856 12493
rect 1092 12257 1176 12493
rect 1412 12257 1496 12493
rect 1732 12257 1816 12493
rect 2052 12257 2136 12493
rect 2372 12257 2456 12493
rect 2692 12257 2776 12493
rect 3012 12257 3456 12493
rect 0 11927 3456 12257
rect 0 11691 215 11927
rect 451 11691 536 11927
rect 772 11691 856 11927
rect 1092 11691 1176 11927
rect 1412 11691 1496 11927
rect 1732 11691 1816 11927
rect 2052 11691 2136 11927
rect 2372 11691 2456 11927
rect 2692 11691 2776 11927
rect 3012 11691 3456 11927
rect 0 11667 3456 11691
rect 0 10565 3456 11347
rect 0 10329 215 10565
rect 451 10329 536 10565
rect 772 10329 856 10565
rect 1092 10329 1176 10565
rect 1412 10329 1496 10565
rect 1732 10329 1816 10565
rect 2052 10329 2136 10565
rect 2372 10329 2456 10565
rect 2692 10329 2776 10565
rect 3012 10329 3456 10565
rect 0 9547 3456 10329
rect 0 9203 3456 9227
rect 0 8967 216 9203
rect 452 8967 537 9203
rect 773 8967 857 9203
rect 1093 8967 1177 9203
rect 1413 8967 1497 9203
rect 1733 8967 1817 9203
rect 2053 8967 2137 9203
rect 2373 8967 2457 9203
rect 2693 8967 2777 9203
rect 3013 8967 3456 9203
rect 0 8597 3456 8967
rect 0 8361 216 8597
rect 452 8361 537 8597
rect 773 8361 857 8597
rect 1093 8361 1177 8597
rect 1413 8361 1497 8597
rect 1733 8361 1817 8597
rect 2053 8361 2137 8597
rect 2373 8361 2457 8597
rect 2693 8361 2777 8597
rect 3013 8361 3456 8597
rect 0 8337 3456 8361
rect 0 7993 3456 8017
rect 0 7757 215 7993
rect 451 7757 536 7993
rect 772 7757 856 7993
rect 1092 7757 1176 7993
rect 1412 7757 1496 7993
rect 1732 7757 1816 7993
rect 2052 7757 2136 7993
rect 2372 7757 2456 7993
rect 2692 7757 2776 7993
rect 3012 7757 3456 7993
rect 0 7627 3456 7757
rect 0 7391 215 7627
rect 451 7391 536 7627
rect 772 7391 856 7627
rect 1092 7391 1176 7627
rect 1412 7391 1496 7627
rect 1732 7391 1816 7627
rect 2052 7391 2136 7627
rect 2372 7391 2456 7627
rect 2692 7391 2776 7627
rect 3012 7391 3456 7627
rect 0 7367 3456 7391
rect 0 7023 3456 7047
rect 0 6787 215 7023
rect 451 6787 536 7023
rect 772 6787 856 7023
rect 1092 6787 1176 7023
rect 1412 6787 1496 7023
rect 1732 6787 1816 7023
rect 2052 6787 2136 7023
rect 2372 6787 2456 7023
rect 2692 6787 2776 7023
rect 3012 6787 3456 7023
rect 0 6657 3456 6787
rect 0 6421 215 6657
rect 451 6421 536 6657
rect 772 6421 856 6657
rect 1092 6421 1176 6657
rect 1412 6421 1496 6657
rect 1732 6421 1816 6657
rect 2052 6421 2136 6657
rect 2372 6421 2456 6657
rect 2692 6421 2776 6657
rect 3012 6421 3456 6657
rect 0 6397 3456 6421
rect 0 6053 3456 6077
rect 0 5817 215 6053
rect 451 5817 536 6053
rect 772 5817 856 6053
rect 1092 5817 1176 6053
rect 1412 5817 1496 6053
rect 1732 5817 1816 6053
rect 2052 5817 2136 6053
rect 2372 5817 2456 6053
rect 2692 5817 2776 6053
rect 3012 5817 3456 6053
rect 0 5447 3456 5817
rect 0 5211 215 5447
rect 451 5211 536 5447
rect 772 5211 856 5447
rect 1092 5211 1176 5447
rect 1412 5211 1496 5447
rect 1732 5211 1816 5447
rect 2052 5211 2136 5447
rect 2372 5211 2456 5447
rect 2692 5211 2776 5447
rect 3012 5211 3456 5447
rect 0 5187 3456 5211
rect 0 4843 3456 4867
rect 0 4607 215 4843
rect 451 4607 536 4843
rect 772 4607 856 4843
rect 1092 4607 1176 4843
rect 1412 4607 1496 4843
rect 1732 4607 1816 4843
rect 2052 4607 2136 4843
rect 2372 4607 2456 4843
rect 2692 4607 2776 4843
rect 3012 4607 3456 4843
rect 0 4237 3456 4607
rect 0 4001 215 4237
rect 451 4001 536 4237
rect 772 4001 856 4237
rect 1092 4001 1176 4237
rect 1412 4001 1496 4237
rect 1732 4001 1816 4237
rect 2052 4001 2136 4237
rect 2372 4001 2456 4237
rect 2692 4001 2776 4237
rect 3012 4001 3456 4237
rect 0 3977 3456 4001
rect 0 3633 3456 3657
rect 0 3397 215 3633
rect 451 3397 536 3633
rect 772 3397 856 3633
rect 1092 3397 1176 3633
rect 1412 3397 1496 3633
rect 1732 3397 1816 3633
rect 2052 3397 2136 3633
rect 2372 3397 2456 3633
rect 2692 3397 2776 3633
rect 3012 3397 3456 3633
rect 0 3267 3456 3397
rect 0 3031 215 3267
rect 451 3031 536 3267
rect 772 3031 856 3267
rect 1092 3031 1176 3267
rect 1412 3031 1496 3267
rect 1732 3031 1816 3267
rect 2052 3031 2136 3267
rect 2372 3031 2456 3267
rect 2692 3031 2776 3267
rect 3012 3031 3456 3267
rect 0 3007 3456 3031
rect 0 2663 3456 2687
rect 0 2427 215 2663
rect 451 2427 536 2663
rect 772 2427 856 2663
rect 1092 2427 1176 2663
rect 1412 2427 1496 2663
rect 1732 2427 1816 2663
rect 2052 2427 2136 2663
rect 2372 2427 2456 2663
rect 2692 2427 2776 2663
rect 3012 2427 3456 2663
rect 0 2057 3456 2427
rect 0 1821 215 2057
rect 451 1821 536 2057
rect 772 1821 856 2057
rect 1092 1821 1176 2057
rect 1412 1821 1496 2057
rect 1732 1821 1816 2057
rect 2052 1821 2136 2057
rect 2372 1821 2456 2057
rect 2692 1821 2776 2057
rect 3012 1821 3456 2057
rect 0 1797 3456 1821
rect 0 1452 3456 1477
rect 0 1216 215 1452
rect 451 1216 536 1452
rect 772 1216 856 1452
rect 1092 1216 1176 1452
rect 1412 1216 1496 1452
rect 1732 1216 1816 1452
rect 2052 1216 2136 1452
rect 2372 1216 2456 1452
rect 2692 1216 2776 1452
rect 3012 1216 3456 1452
rect 0 1070 3456 1216
rect 0 834 215 1070
rect 451 834 536 1070
rect 772 834 856 1070
rect 1092 834 1176 1070
rect 1412 834 1496 1070
rect 1732 834 1816 1070
rect 2052 834 2136 1070
rect 2372 834 2456 1070
rect 2692 834 2776 1070
rect 3012 834 3456 1070
rect 0 688 3456 834
rect 0 452 215 688
rect 451 452 536 688
rect 772 452 856 688
rect 1092 452 1176 688
rect 1412 452 1496 688
rect 1732 452 1816 688
rect 2052 452 2136 688
rect 2372 452 2456 688
rect 2692 452 2776 688
rect 3012 452 3456 688
rect 0 427 3456 452
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_0
timestamp 1707688321
transform -1 0 2880 0 -1 38972
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_1
timestamp 1707688321
transform -1 0 2880 0 -1 36842
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_2
timestamp 1707688321
transform -1 0 2880 0 -1 34712
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_3
timestamp 1707688321
transform -1 0 2880 0 1 30582
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_4
timestamp 1707688321
transform -1 0 2880 0 -1 30452
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_5
timestamp 1707688321
transform -1 0 2880 0 1 26322
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_6
timestamp 1707688321
transform -1 0 2880 0 -1 26192
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_7
timestamp 1707688321
transform -1 0 2880 0 1 22062
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_8
timestamp 1707688321
transform -1 0 2880 0 -1 21932
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_9
timestamp 1707688321
transform -1 0 2880 0 1 17802
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_10
timestamp 1707688321
transform -1 0 2880 0 -1 17672
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_11
timestamp 1707688321
transform -1 0 2880 0 1 13542
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_12
timestamp 1707688321
transform -1 0 2880 0 -1 13412
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_13
timestamp 1707688321
transform -1 0 2880 0 1 9282
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_14
timestamp 1707688321
transform -1 0 2880 0 -1 9152
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_15
timestamp 1707688321
transform -1 0 2880 0 1 5022
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_16
timestamp 1707688321
transform -1 0 2880 0 -1 4892
box -82 -32 2386 2032
use nfet_CDNS_55959141808712  nfet_CDNS_55959141808712_17
timestamp 1707688321
transform -1 0 2880 0 1 762
box -82 -32 2386 2032
<< labels >>
flabel metal3 s 1495 0 1895 166 3 FreeSans 520 0 0 0 cpos
port 1 nsew power bidirectional
flabel metal3 s 2095 0 2695 166 3 FreeSans 520 0 0 0 cneg
port 2 nsew ground bidirectional
flabel metal3 s 695 0 1295 166 3 FreeSans 520 0 0 0 cneg
port 2 nsew ground bidirectional
flabel metal5 s 3202 35157 3456 40000 3 FreeSans 520 180 0 0 vssio
port 3 nsew ground bidirectional
flabel metal5 s 3202 12837 3456 13687 3 FreeSans 520 180 0 0 vddio_q
port 4 nsew power bidirectional
flabel metal5 s 3202 14007 3456 18997 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 3202 11667 3456 12517 3 FreeSans 520 180 0 0 vssio_q
port 6 nsew ground bidirectional
flabel metal5 s 3202 1797 3456 2687 3 FreeSans 520 180 0 0 vccd
port 7 nsew power bidirectional
flabel metal5 s 3202 7367 3456 8017 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal5 s 3202 3977 3456 4867 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 3202 427 3456 1477 3 FreeSans 520 180 0 0 vcchib
port 9 nsew power bidirectional
flabel metal5 s 3202 6397 3456 7047 3 FreeSans 520 180 0 0 vswitch
port 10 nsew power bidirectional
flabel metal5 s 3202 5187 3456 6077 3 FreeSans 520 180 0 0 vssio
port 3 nsew ground bidirectional
flabel metal5 s 3263 3007 3456 3657 3 FreeSans 520 180 0 0 vdda
port 11 nsew power bidirectional
flabel metal5 s 3202 8337 3456 9227 3 FreeSans 520 180 0 0 vssd
port 12 nsew ground bidirectional
flabel metal5 s 3202 9547 3456 11347 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 vssd
port 12 nsew ground bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 vdda
port 11 nsew power bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 vssio_q
port 6 nsew ground bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 vssio
port 3 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 vswitch
port 10 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 vcchib
port 9 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 0 7367 254 8017 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 vccd
port 7 nsew power bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 vssio
port 3 nsew ground bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 vddio_q
port 4 nsew power bidirectional
flabel metal4 s 3202 14007 3456 19000 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 3202 35157 3456 39999 3 FreeSans 520 180 0 0 vssio
port 3 nsew ground bidirectional
flabel metal4 s 3202 9673 3456 10269 3 FreeSans 520 180 0 0 amuxbus_b
port 13 nsew signal bidirectional
flabel metal4 s 3202 1777 3456 2707 3 FreeSans 520 180 0 0 vccd
port 7 nsew power bidirectional
flabel metal4 s 3202 12817 3456 13707 3 FreeSans 520 180 0 0 vddio_q
port 4 nsew power bidirectional
flabel metal4 s 3202 7347 3456 8037 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 3202 3957 3456 4887 3 FreeSans 520 180 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 3202 407 3456 1497 3 FreeSans 520 180 0 0 vcchib
port 9 nsew power bidirectional
flabel metal4 s 3202 6377 3456 7067 3 FreeSans 520 180 0 0 vswitch
port 10 nsew power bidirectional
flabel metal4 s 3202 5167 3456 6097 3 FreeSans 520 180 0 0 vssio
port 3 nsew ground bidirectional
flabel metal4 s 3202 11647 3456 12537 3 FreeSans 520 180 0 0 vssio_q
port 6 nsew ground bidirectional
flabel metal4 s 3263 2987 3456 3677 3 FreeSans 520 180 0 0 vdda
port 11 nsew power bidirectional
flabel metal4 s 3202 8317 3456 9247 3 FreeSans 520 180 0 0 vssd
port 12 nsew ground bidirectional
flabel metal4 s 3202 10625 3456 11221 3 FreeSans 520 180 0 0 amuxbus_a
port 14 nsew signal bidirectional
flabel metal4 s 3202 9547 3456 9613 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 3202 10329 3456 10565 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 3202 11281 3456 11347 3 FreeSans 520 180 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 amuxbus_a
port 14 nsew signal bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 vssd
port 12 nsew ground bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 vdda
port 11 nsew power bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 vssio_q
port 6 nsew ground bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 vssio
port 3 nsew ground bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 vswitch
port 10 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 vcchib
port 9 nsew power bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 vssa
port 8 nsew ground bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 vccd
port 7 nsew power bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 amuxbus_b
port 13 nsew signal bidirectional
flabel metal4 s 0 35157 254 39999 3 FreeSans 520 0 0 0 vssio
port 3 nsew ground bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 vddio
port 5 nsew power bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 vddio_q
port 4 nsew power bidirectional
flabel metal2 s 2095 0 2695 242 3 FreeSans 520 0 0 0 cneg
port 2 nsew ground bidirectional
flabel metal2 s 695 0 1295 242 3 FreeSans 520 0 0 0 cneg
port 2 nsew ground bidirectional
flabel metal2 s 1495 0 1895 242 3 FreeSans 520 0 0 0 cpos
port 1 nsew power bidirectional
flabel comment s 2618 329 2618 329 0 FreeSans 400 0 0 0 condiode
rlabel metal3 s 2095 0 2695 166 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 0 1295 39165 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2095 0 2695 39165 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39333 1463 39341 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39319 1449 39333 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39305 1435 39319 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39291 1421 39305 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39277 1407 39291 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39263 1393 39277 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39249 1379 39263 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39235 1365 39249 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39221 1351 39235 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39207 1337 39221 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39193 1323 39207 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39179 1309 39193 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39165 1295 39179 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1927 39333 2695 39341 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1941 39319 2695 39333 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1955 39305 2695 39319 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1969 39291 2695 39305 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1983 39277 2695 39291 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1997 39263 2695 39277 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2011 39249 2695 39263 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2025 39235 2695 39249 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2039 39221 2695 39235 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2053 39207 2695 39221 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2067 39193 2695 39207 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2081 39179 2695 39193 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2095 39165 2695 39179 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 39341 2695 39782 1 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1495 0 1895 39063 1 cpos
port 1 nsew power bidirectional
rlabel metal4 s 0 8317 3456 9247 1 vssd
port 12 nsew ground bidirectional
rlabel metal4 s 0 2987 3456 3677 1 vdda
port 11 nsew power bidirectional
rlabel metal4 s 0 6377 3456 7067 1 vswitch
port 10 nsew power bidirectional
rlabel metal4 s 0 407 3456 1497 1 vcchib
port 9 nsew power bidirectional
rlabel metal5 s 0 9547 3456 11347 1 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 7347 3456 8037 1 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 9547 3456 9613 1 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 10329 3456 10565 1 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 11281 3456 11347 1 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 1777 3456 2707 1 vccd
port 7 nsew power bidirectional
rlabel metal4 s 0 11647 3456 12537 1 vssio_q
port 6 nsew ground bidirectional
rlabel metal5 s 0 14007 3456 18997 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 3957 3456 4887 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 14007 3456 19000 1 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 12817 3456 13707 1 vddio_q
port 4 nsew power bidirectional
rlabel metal5 s 0 35157 3456 40000 1 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 0 5167 3456 6097 1 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 0 35157 3456 40000 1 vssio
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 3456 40000
string GDS_END 9654072
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8300788
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
