magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 189 636
<< pmos >>
rect 0 0 100 600
<< pdiff >>
rect -50 0 0 600
rect 100 0 150 600
<< poly >>
rect 0 600 100 632
rect 0 -32 100 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 636
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_1
timestamp 1707688321
transform 1 0 100 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80642596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80641710
<< end >>
