magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 35 3488 61 4329
rect 1081 3565 1431 4292
rect 2533 3488 2559 4329
<< pwell >>
rect 790 4304 998 4390
rect 790 3467 998 3553
<< psubdiff >>
rect 816 4330 840 4364
rect 874 4330 914 4364
rect 948 4330 972 4364
rect 816 3493 840 3527
rect 874 3493 914 3527
rect 948 3493 972 3527
<< nsubdiff >>
rect 1330 4176 1364 4225
rect 1330 4108 1364 4142
rect 1330 4040 1364 4074
rect 1330 3972 1364 4006
rect 1330 3904 1364 3938
rect 1330 3836 1364 3870
rect 1330 3768 1364 3802
rect 1330 3700 1364 3734
rect 1330 3632 1364 3666
<< psubdiffcont >>
rect 840 4330 874 4364
rect 914 4330 948 4364
rect 840 3493 874 3527
rect 914 3493 948 3527
<< nsubdiffcont >>
rect 1330 4142 1364 4176
rect 1330 4074 1364 4108
rect 1330 4006 1364 4040
rect 1330 3938 1364 3972
rect 1330 3870 1364 3904
rect 1330 3802 1364 3836
rect 1330 3734 1364 3768
rect 1330 3666 1364 3700
<< poly >>
rect 869 4008 1003 4024
rect 869 3974 885 4008
rect 919 3974 953 4008
rect 987 3974 1003 4008
rect 869 3958 1003 3974
rect 1086 4008 1220 4024
rect 1086 3974 1102 4008
rect 1136 3974 1170 4008
rect 1204 3974 1220 4008
rect 1086 3958 1220 3974
rect 869 3883 1003 3899
rect 869 3849 885 3883
rect 919 3849 953 3883
rect 987 3849 1003 3883
rect 869 3833 1003 3849
rect 1086 3883 1220 3899
rect 1086 3849 1102 3883
rect 1136 3849 1170 3883
rect 1204 3849 1220 3883
rect 1086 3833 1220 3849
rect 428 3506 562 3522
rect 428 3472 444 3506
rect 478 3472 512 3506
rect 546 3472 562 3506
rect 2032 3506 2166 3522
rect 428 3456 562 3472
rect 2032 3472 2048 3506
rect 2082 3472 2116 3506
rect 2150 3472 2166 3506
rect 2032 3456 2166 3472
rect 971 1872 1105 1888
rect 971 1838 987 1872
rect 1021 1838 1055 1872
rect 1089 1838 1105 1872
rect 971 1822 1105 1838
rect 1489 1872 1623 1888
rect 1489 1838 1505 1872
rect 1539 1838 1573 1872
rect 1607 1838 1623 1872
rect 1489 1822 1623 1838
<< polycont >>
rect 885 3974 919 4008
rect 953 3974 987 4008
rect 1102 3974 1136 4008
rect 1170 3974 1204 4008
rect 885 3849 919 3883
rect 953 3849 987 3883
rect 1102 3849 1136 3883
rect 1170 3849 1204 3883
rect 444 3472 478 3506
rect 512 3472 546 3506
rect 2048 3472 2082 3506
rect 2116 3472 2150 3506
rect 987 1838 1021 1872
rect 1055 1838 1089 1872
rect 1505 1838 1539 1872
rect 1573 1838 1607 1872
<< locali >>
rect 816 4330 820 4364
rect 874 4330 892 4364
rect 948 4330 972 4364
rect 823 4199 857 4237
rect 823 4127 857 4165
rect 930 4121 964 4170
rect 397 4010 431 4058
rect 397 3928 431 3976
rect 397 3846 431 3894
rect 397 3764 431 3812
rect 397 3682 431 3730
rect 397 3600 431 3648
rect 1125 4132 1159 4170
rect 1231 4132 1265 4214
rect 1330 4176 1364 4214
rect 1330 4108 1364 4135
rect 573 4010 607 4058
rect 1330 4040 1364 4056
rect 573 3928 607 3976
rect 869 3974 885 4008
rect 940 3974 953 4008
rect 1086 3974 1102 4008
rect 1137 3974 1170 4008
rect 1209 3974 1220 4008
rect 573 3846 607 3894
rect 1330 3972 1364 3977
rect 1330 3931 1364 3938
rect 869 3849 885 3883
rect 940 3849 953 3883
rect 1097 3849 1102 3883
rect 1169 3849 1170 3883
rect 1204 3849 1220 3883
rect 1330 3851 1364 3870
rect 573 3764 607 3812
rect 573 3682 607 3730
rect 573 3600 607 3648
rect 823 3692 857 3730
rect 823 3620 857 3658
rect 930 3677 964 3715
rect 1125 3689 1159 3746
rect 1231 3721 1265 3759
rect 1330 3771 1364 3802
rect 1330 3700 1364 3734
rect 1125 3598 1159 3655
rect 1330 3611 1364 3657
rect 1987 4010 2021 4058
rect 1987 3928 2021 3976
rect 1987 3846 2021 3894
rect 1987 3764 2021 3812
rect 1987 3682 2021 3730
rect 1987 3600 2021 3648
rect 2163 4010 2197 4058
rect 2163 3928 2197 3976
rect 2163 3846 2197 3894
rect 2163 3764 2197 3812
rect 2163 3682 2197 3730
rect 2163 3600 2197 3648
rect 428 3472 437 3506
rect 478 3472 509 3506
rect 546 3472 562 3506
rect 816 3493 820 3527
rect 874 3493 892 3527
rect 948 3493 972 3527
rect 2032 3472 2048 3506
rect 2085 3472 2116 3506
rect 2157 3472 2166 3506
rect 971 1838 983 1872
rect 1021 1838 1055 1872
rect 1089 1838 1105 1872
rect 1489 1838 1505 1872
rect 1539 1838 1573 1872
rect 1611 1838 1623 1872
rect 926 1704 960 1742
rect 926 1632 960 1670
rect 1102 1704 1136 1742
rect 1102 1632 1136 1670
rect 1458 1704 1492 1742
rect 1458 1632 1492 1670
rect 1634 1704 1668 1742
rect 1634 1632 1668 1670
<< viali >>
rect 820 4330 840 4364
rect 840 4330 854 4364
rect 892 4330 914 4364
rect 914 4330 926 4364
rect 823 4237 857 4271
rect 1231 4214 1265 4248
rect 823 4165 857 4199
rect 823 4093 857 4127
rect 930 4170 964 4204
rect 397 4058 431 4092
rect 397 3976 431 4010
rect 397 3894 431 3928
rect 397 3812 431 3846
rect 397 3730 431 3764
rect 397 3648 431 3682
rect 397 3566 431 3600
rect 573 4058 607 4092
rect 930 4087 964 4121
rect 1125 4170 1159 4204
rect 1125 4098 1159 4132
rect 1231 4098 1265 4132
rect 1330 4214 1364 4248
rect 1330 4142 1364 4169
rect 1330 4135 1364 4142
rect 573 3976 607 4010
rect 1330 4074 1364 4090
rect 1330 4056 1364 4074
rect 906 3974 919 4008
rect 919 3974 940 4008
rect 978 3974 987 4008
rect 987 3974 1012 4008
rect 1103 3974 1136 4008
rect 1136 3974 1137 4008
rect 1175 3974 1204 4008
rect 1204 3974 1209 4008
rect 1330 4006 1364 4011
rect 1330 3977 1364 4006
rect 573 3894 607 3928
rect 1330 3904 1364 3931
rect 1330 3897 1364 3904
rect 906 3849 919 3883
rect 919 3849 940 3883
rect 978 3849 987 3883
rect 987 3849 1012 3883
rect 1063 3849 1097 3883
rect 1135 3849 1136 3883
rect 1136 3849 1169 3883
rect 573 3812 607 3846
rect 1330 3836 1364 3851
rect 1330 3817 1364 3836
rect 573 3730 607 3764
rect 573 3648 607 3682
rect 573 3566 607 3600
rect 823 3730 857 3764
rect 823 3658 857 3692
rect 930 3715 964 3749
rect 930 3643 964 3677
rect 1125 3746 1159 3780
rect 1125 3655 1159 3689
rect 1231 3759 1265 3793
rect 1231 3687 1265 3721
rect 1330 3768 1364 3771
rect 1330 3737 1364 3768
rect 823 3586 857 3620
rect 1125 3564 1159 3598
rect 1330 3666 1364 3691
rect 1330 3657 1364 3666
rect 1330 3577 1364 3611
rect 1987 4058 2021 4092
rect 1987 3976 2021 4010
rect 1987 3894 2021 3928
rect 1987 3812 2021 3846
rect 1987 3730 2021 3764
rect 1987 3648 2021 3682
rect 1987 3566 2021 3600
rect 2163 4058 2197 4092
rect 2163 3976 2197 4010
rect 2163 3894 2197 3928
rect 2163 3812 2197 3846
rect 2163 3730 2197 3764
rect 2163 3648 2197 3682
rect 2163 3566 2197 3600
rect 437 3472 444 3506
rect 444 3472 471 3506
rect 509 3472 512 3506
rect 512 3472 543 3506
rect 820 3493 840 3527
rect 840 3493 854 3527
rect 892 3493 914 3527
rect 914 3493 926 3527
rect 2051 3472 2082 3506
rect 2082 3472 2085 3506
rect 2123 3472 2150 3506
rect 2150 3472 2157 3506
rect 983 1838 987 1872
rect 987 1838 1017 1872
rect 1055 1838 1089 1872
rect 1505 1838 1539 1872
rect 1577 1838 1607 1872
rect 1607 1838 1611 1872
rect 926 1742 960 1776
rect 926 1670 960 1704
rect 926 1598 960 1632
rect 1102 1742 1136 1776
rect 1102 1670 1136 1704
rect 1102 1598 1136 1632
rect 1458 1742 1492 1776
rect 1458 1670 1492 1704
rect 1458 1598 1492 1632
rect 1634 1742 1668 1776
rect 1634 1670 1668 1704
rect 1634 1598 1668 1632
<< metal1 >>
rect 721 4364 938 4370
rect 721 4330 820 4364
rect 854 4330 892 4364
rect 926 4330 938 4364
rect 111 4222 681 4329
rect 721 4324 938 4330
rect 721 4271 863 4324
tri 863 4290 897 4324 nw
rect 721 4237 823 4271
rect 857 4237 863 4271
tri 357 4214 365 4222 ne
rect 365 4214 463 4222
tri 463 4214 471 4222 nw
tri 365 4204 375 4214 ne
rect 375 4204 453 4214
tri 453 4204 463 4214 nw
tri 375 4199 380 4204 ne
rect 380 4199 448 4204
tri 448 4199 453 4204 nw
rect 721 4199 863 4237
rect 1225 4248 1370 4260
tri 380 4188 391 4199 ne
rect 391 4092 437 4199
tri 437 4188 448 4199 nw
rect 721 4165 823 4199
rect 857 4165 863 4199
rect 721 4127 863 4165
rect 391 4058 397 4092
rect 431 4058 437 4092
rect 391 4010 437 4058
rect 391 3976 397 4010
rect 431 3976 437 4010
rect 391 3928 437 3976
rect 391 3894 397 3928
rect 431 3894 437 3928
rect 391 3846 437 3894
rect 391 3812 397 3846
rect 431 3812 437 3846
rect 391 3764 437 3812
rect 391 3730 397 3764
rect 431 3730 437 3764
tri 388 3715 391 3718 se
rect 391 3715 437 3730
tri 365 3692 388 3715 se
rect 388 3692 437 3715
tri 357 3684 365 3692 se
rect 365 3684 437 3692
rect 325 3682 437 3684
rect 325 3648 397 3682
rect 431 3648 437 3682
rect 325 3600 437 3648
rect 325 3566 397 3600
rect 431 3566 437 3600
rect 325 3554 437 3566
rect 564 4092 616 4104
rect 564 4058 573 4092
rect 607 4058 616 4092
rect 564 4010 616 4058
rect 564 3976 573 4010
rect 607 3976 616 4010
rect 564 3928 616 3976
rect 564 3894 573 3928
rect 607 3894 616 3928
rect 564 3846 616 3894
rect 564 3812 573 3846
rect 607 3812 616 3846
rect 564 3764 616 3812
rect 564 3755 573 3764
rect 607 3755 616 3764
rect 564 3691 616 3703
rect 564 3600 616 3639
rect 564 3566 573 3600
rect 607 3566 616 3600
rect 564 3554 616 3566
rect 721 4093 823 4127
rect 857 4093 863 4127
rect 721 4081 863 4093
rect 924 4204 1168 4216
rect 924 4170 930 4204
rect 964 4197 1125 4204
rect 1159 4197 1168 4204
rect 964 4170 1116 4197
rect 924 4145 1116 4170
rect 924 4133 1168 4145
rect 924 4121 1116 4133
rect 924 4087 930 4121
rect 964 4087 1116 4121
rect 924 4081 1116 4087
rect 1225 4214 1231 4248
rect 1265 4214 1330 4248
rect 1364 4214 1370 4248
rect 1980 4222 2537 4329
rect 1225 4169 1370 4214
tri 2123 4188 2157 4222 ne
rect 1225 4135 1330 4169
rect 1364 4135 1370 4169
rect 1225 4132 1370 4135
rect 1225 4098 1231 4132
rect 1265 4098 1370 4132
rect 1225 4090 1370 4098
rect 1225 4086 1330 4090
tri 1290 4081 1295 4086 ne
rect 1295 4081 1330 4086
rect 721 4075 845 4081
tri 845 4075 851 4081 nw
rect 924 4075 1168 4081
tri 1295 4075 1301 4081 ne
rect 1301 4075 1330 4081
rect 721 4056 826 4075
tri 826 4056 845 4075 nw
tri 1301 4056 1320 4075 ne
rect 1320 4056 1330 4075
rect 1364 4056 1370 4090
rect 721 4052 822 4056
tri 822 4052 826 4056 nw
tri 1320 4052 1324 4056 ne
rect 721 3793 817 4052
tri 817 4047 822 4052 nw
rect 845 3968 851 4020
rect 903 4008 915 4020
rect 967 4008 1097 4020
rect 903 3974 906 4008
rect 967 3974 978 4008
rect 1012 3974 1097 4008
rect 903 3968 915 3974
rect 967 3968 1097 3974
rect 1149 3968 1163 4020
rect 1215 3968 1274 4020
tri 1188 3934 1222 3968 ne
rect 894 3883 1057 3892
rect 894 3849 906 3883
rect 940 3849 978 3883
rect 1012 3849 1057 3883
rect 894 3840 1057 3849
rect 1109 3840 1123 3892
rect 1175 3840 1181 3892
tri 817 3793 834 3810 sw
rect 1222 3793 1274 3968
rect 721 3792 834 3793
tri 834 3792 835 3793 sw
rect 721 3780 835 3792
tri 835 3780 847 3792 sw
rect 1119 3780 1165 3792
rect 721 3776 847 3780
tri 847 3776 851 3780 sw
rect 721 3764 863 3776
rect 721 3730 823 3764
rect 857 3730 863 3764
rect 721 3692 863 3730
rect 721 3658 823 3692
rect 857 3658 863 3692
rect 721 3620 863 3658
rect 921 3753 973 3761
rect 921 3689 973 3701
rect 1119 3746 1125 3780
rect 1159 3746 1165 3780
rect 1119 3689 1165 3746
tri 1118 3655 1119 3656 se
rect 1119 3655 1125 3689
rect 1159 3655 1165 3689
rect 1222 3759 1231 3793
rect 1265 3759 1274 3793
rect 1222 3721 1274 3759
rect 1222 3687 1231 3721
rect 1265 3687 1274 3721
rect 1222 3675 1274 3687
rect 1324 4011 1370 4056
rect 1324 3977 1330 4011
rect 1364 3977 1370 4011
rect 1324 3931 1370 3977
rect 1324 3897 1330 3931
rect 1364 3897 1370 3931
rect 1324 3851 1370 3897
rect 1324 3817 1330 3851
rect 1364 3817 1370 3851
rect 1324 3771 1370 3817
rect 1324 3737 1330 3771
rect 1364 3737 1370 3771
rect 1324 3691 1370 3737
rect 1324 3657 1330 3691
rect 1364 3657 1370 3691
tri 1111 3648 1118 3655 se
rect 1118 3648 1165 3655
tri 1165 3648 1173 3656 sw
tri 1316 3648 1324 3656 se
rect 1324 3648 1370 3657
rect 921 3631 973 3637
tri 1094 3631 1111 3648 se
rect 1111 3631 1173 3648
tri 1173 3631 1190 3648 sw
tri 1299 3631 1316 3648 se
rect 1316 3631 1370 3648
tri 1085 3622 1094 3631 se
rect 1094 3622 1190 3631
tri 1190 3622 1199 3631 sw
tri 1290 3622 1299 3631 se
rect 1299 3622 1370 3631
rect 721 3586 823 3620
rect 857 3586 863 3620
rect 721 3564 863 3586
rect 1062 3616 1370 3622
tri 863 3564 866 3567 sw
rect 327 3527 334 3554
tri 334 3527 361 3554 nw
rect 721 3533 866 3564
tri 866 3533 897 3564 sw
rect 721 3527 938 3533
tri 327 3520 334 3527 nw
rect 408 3463 414 3515
rect 466 3506 478 3515
rect 530 3506 555 3515
rect 471 3472 478 3506
rect 543 3472 555 3506
rect 721 3493 820 3527
rect 854 3493 892 3527
rect 926 3493 938 3527
rect 1062 3500 1101 3616
rect 1217 3611 1370 3616
rect 1217 3577 1330 3611
rect 1364 3577 1370 3611
rect 1217 3500 1370 3577
rect 1978 4092 2030 4104
rect 1978 4058 1987 4092
rect 2021 4058 2030 4092
rect 1978 4010 2030 4058
rect 1978 3976 1987 4010
rect 2021 3976 2030 4010
rect 1978 3928 2030 3976
rect 1978 3894 1987 3928
rect 2021 3894 2030 3928
rect 1978 3846 2030 3894
rect 1978 3812 1987 3846
rect 2021 3812 2030 3846
rect 1978 3764 2030 3812
rect 1978 3730 1987 3764
rect 2021 3730 2030 3764
rect 1978 3690 2030 3730
rect 1978 3626 2030 3638
rect 1978 3566 1987 3574
rect 2021 3566 2030 3574
rect 1978 3554 2030 3566
rect 2157 4092 2203 4222
tri 2203 4188 2237 4222 nw
tri 2483 4188 2517 4222 nw
rect 2157 4058 2163 4092
rect 2197 4058 2203 4092
rect 2157 4010 2203 4058
rect 2157 3976 2163 4010
rect 2197 3976 2203 4010
rect 2157 3928 2203 3976
rect 2157 3894 2163 3928
rect 2197 3894 2203 3928
rect 2157 3846 2203 3894
rect 2157 3812 2163 3846
rect 2197 3812 2203 3846
rect 2157 3764 2203 3812
rect 2157 3730 2163 3764
rect 2197 3730 2203 3764
rect 2157 3684 2203 3730
tri 2203 3684 2237 3718 sw
rect 2157 3682 2269 3684
rect 2157 3648 2163 3682
rect 2197 3648 2269 3682
rect 2157 3600 2269 3648
rect 2157 3566 2163 3600
rect 2197 3566 2269 3600
rect 2157 3554 2269 3566
tri 2233 3520 2267 3554 ne
rect 1062 3494 1370 3500
rect 721 3487 938 3493
rect 466 3463 478 3472
rect 530 3463 555 3472
rect 1818 3463 1824 3515
rect 1876 3463 1888 3515
rect 1940 3506 2169 3515
rect 1940 3472 2051 3506
rect 2085 3472 2123 3506
rect 2157 3472 2169 3506
rect 1940 3463 2169 3472
rect 703 3169 1697 3369
rect 141 3070 935 3122
rect 987 3070 999 3122
rect 1051 3070 2447 3122
rect 849 2938 855 2990
rect 907 2938 919 2990
rect 971 2938 977 2990
rect 1542 2858 1548 2910
rect 1600 2858 1612 2910
rect 1664 2858 1670 2910
rect 1818 2858 1824 2910
rect 1876 2858 1888 2910
rect 1940 2858 1946 2910
rect 1057 2824 1602 2830
rect 1057 2772 1101 2824
rect 1153 2772 1165 2824
rect 1217 2772 1602 2824
rect 1057 2756 1602 2772
rect 354 2642 541 2741
rect 1057 2704 1101 2756
rect 1153 2704 1165 2756
rect 1217 2704 1602 2756
rect 1057 2688 1602 2704
rect 1057 2636 1101 2688
rect 1153 2636 1165 2688
rect 1217 2636 1602 2688
rect 1057 2630 1602 2636
rect 166 2547 257 2581
rect 1057 2538 1537 2590
rect 163 2464 227 2501
rect 1057 2458 1537 2510
rect 141 2374 494 2426
rect 546 2374 558 2426
rect 610 2374 1011 2426
rect 1063 2374 1075 2426
rect 1127 2374 1201 2426
rect 141 2290 1468 2342
rect 1520 2290 1532 2342
rect 1584 2290 1984 2342
rect 2036 2290 2048 2342
rect 2100 2290 2499 2342
rect 925 1829 931 1881
rect 983 1872 995 1881
rect 1047 1872 1101 1881
rect 1047 1838 1055 1872
rect 1089 1838 1101 1872
rect 983 1829 995 1838
rect 1047 1829 1101 1838
rect 1493 1872 1548 1881
rect 1600 1872 1612 1881
rect 1493 1838 1505 1872
rect 1539 1838 1548 1872
rect 1611 1838 1612 1872
rect 1493 1829 1548 1838
rect 1600 1829 1612 1838
rect 1664 1829 1670 1881
rect 920 1776 966 1788
tri 900 1742 920 1762 se
rect 920 1742 926 1776
rect 960 1742 966 1776
tri 886 1728 900 1742 se
rect 900 1728 966 1742
rect 845 1704 966 1728
rect 845 1670 926 1704
rect 960 1670 966 1704
rect 845 1632 966 1670
rect 845 1598 926 1632
rect 960 1598 966 1632
rect 845 1427 966 1598
rect 1081 1776 1142 1788
rect 1081 1742 1102 1776
rect 1136 1742 1142 1776
rect 1081 1716 1142 1742
rect 1133 1704 1142 1716
rect 1136 1670 1142 1704
rect 1133 1664 1142 1670
rect 1081 1652 1142 1664
rect 1133 1632 1142 1652
rect 1081 1598 1102 1600
rect 1136 1598 1142 1632
rect 1081 1586 1142 1598
rect 1452 1776 1514 1788
rect 1452 1742 1458 1776
rect 1492 1742 1514 1776
rect 1452 1716 1514 1742
rect 1452 1704 1462 1716
rect 1452 1670 1458 1704
rect 1452 1664 1462 1670
rect 1452 1652 1514 1664
rect 1452 1632 1462 1652
rect 1452 1598 1458 1632
rect 1492 1598 1514 1600
rect 1452 1586 1514 1598
rect 1628 1776 1674 1788
rect 1628 1742 1634 1776
rect 1668 1742 1674 1776
rect 1628 1728 1674 1742
tri 1674 1728 1708 1762 sw
rect 1628 1704 1749 1728
rect 1628 1670 1634 1704
rect 1668 1670 1749 1704
rect 1628 1632 1749 1670
rect 1628 1598 1634 1632
rect 1668 1598 1749 1632
tri 966 1433 1000 1467 sw
tri 1594 1433 1628 1467 se
rect 845 1375 867 1427
rect 919 1375 966 1427
rect 845 1346 966 1375
rect 845 1294 867 1346
rect 919 1294 966 1346
rect 845 1265 966 1294
rect 845 1213 867 1265
rect 919 1213 966 1265
rect 845 1207 966 1213
rect 1628 1207 1749 1598
rect 1329 606 1381 612
tri 1295 516 1329 550 se
rect 1329 542 1381 554
rect 926 490 1329 516
tri 1381 516 1415 550 sw
rect 1381 490 1700 516
rect 926 484 1700 490
rect 800 414 935 448
tri 935 414 969 448 sw
rect 800 402 969 414
tri 969 402 981 414 sw
tri 892 399 895 402 ne
rect 895 399 981 402
tri 981 399 984 402 sw
rect 1677 399 1683 451
rect 1735 399 1749 451
rect 1801 399 2004 451
tri 895 358 936 399 ne
rect 936 362 984 399
tri 984 362 1021 399 sw
rect 936 358 1021 362
tri 936 325 969 358 ne
rect 969 352 1021 358
rect 969 288 1021 300
rect 969 230 1021 236
rect 842 196 941 202
rect 507 67 840 155
rect 842 144 865 196
rect 917 144 941 196
rect 842 132 941 144
rect 842 80 865 132
rect 917 80 941 132
rect 842 74 941 80
<< via1 >>
rect 564 3730 573 3755
rect 573 3730 607 3755
rect 607 3730 616 3755
rect 564 3703 616 3730
rect 564 3682 616 3691
rect 564 3648 573 3682
rect 573 3648 607 3682
rect 607 3648 616 3682
rect 564 3639 616 3648
rect 1116 4170 1125 4197
rect 1125 4170 1159 4197
rect 1159 4170 1168 4197
rect 1116 4145 1168 4170
rect 1116 4132 1168 4133
rect 1116 4098 1125 4132
rect 1125 4098 1159 4132
rect 1159 4098 1168 4132
rect 1116 4081 1168 4098
rect 851 3968 903 4020
rect 915 4008 967 4020
rect 1097 4008 1149 4020
rect 915 3974 940 4008
rect 940 3974 967 4008
rect 1097 3974 1103 4008
rect 1103 3974 1137 4008
rect 1137 3974 1149 4008
rect 915 3968 967 3974
rect 1097 3968 1149 3974
rect 1163 4008 1215 4020
rect 1163 3974 1175 4008
rect 1175 3974 1209 4008
rect 1209 3974 1215 4008
rect 1163 3968 1215 3974
rect 1057 3883 1109 3892
rect 1057 3849 1063 3883
rect 1063 3849 1097 3883
rect 1097 3849 1109 3883
rect 1057 3840 1109 3849
rect 1123 3883 1175 3892
rect 1123 3849 1135 3883
rect 1135 3849 1169 3883
rect 1169 3849 1175 3883
rect 1123 3840 1175 3849
rect 921 3749 973 3753
rect 921 3715 930 3749
rect 930 3715 964 3749
rect 964 3715 973 3749
rect 921 3701 973 3715
rect 921 3677 973 3689
rect 921 3643 930 3677
rect 930 3643 964 3677
rect 964 3643 973 3677
rect 921 3637 973 3643
rect 414 3506 466 3515
rect 478 3506 530 3515
rect 414 3472 437 3506
rect 437 3472 466 3506
rect 478 3472 509 3506
rect 509 3472 530 3506
rect 1101 3598 1217 3616
rect 1101 3564 1125 3598
rect 1125 3564 1159 3598
rect 1159 3564 1217 3598
rect 1101 3500 1217 3564
rect 1978 3682 2030 3690
rect 1978 3648 1987 3682
rect 1987 3648 2021 3682
rect 2021 3648 2030 3682
rect 1978 3638 2030 3648
rect 1978 3600 2030 3626
rect 1978 3574 1987 3600
rect 1987 3574 2021 3600
rect 2021 3574 2030 3600
rect 414 3463 466 3472
rect 478 3463 530 3472
rect 1824 3463 1876 3515
rect 1888 3463 1940 3515
rect 935 3070 987 3122
rect 999 3070 1051 3122
rect 855 2938 907 2990
rect 919 2938 971 2990
rect 1548 2858 1600 2910
rect 1612 2858 1664 2910
rect 1824 2858 1876 2910
rect 1888 2858 1940 2910
rect 1101 2772 1153 2824
rect 1165 2772 1217 2824
rect 1101 2704 1153 2756
rect 1165 2704 1217 2756
rect 1101 2636 1153 2688
rect 1165 2636 1217 2688
rect 494 2374 546 2426
rect 558 2374 610 2426
rect 1011 2374 1063 2426
rect 1075 2374 1127 2426
rect 1468 2290 1520 2342
rect 1532 2290 1584 2342
rect 1984 2290 2036 2342
rect 2048 2290 2100 2342
rect 931 1829 983 1881
rect 995 1872 1047 1881
rect 995 1838 1017 1872
rect 1017 1838 1047 1872
rect 995 1829 1047 1838
rect 1548 1872 1600 1881
rect 1548 1838 1577 1872
rect 1577 1838 1600 1872
rect 1548 1829 1600 1838
rect 1612 1829 1664 1881
rect 1081 1704 1133 1716
rect 1081 1670 1102 1704
rect 1102 1670 1133 1704
rect 1081 1664 1133 1670
rect 1081 1632 1133 1652
rect 1081 1600 1102 1632
rect 1102 1600 1133 1632
rect 1462 1704 1514 1716
rect 1462 1670 1492 1704
rect 1492 1670 1514 1704
rect 1462 1664 1514 1670
rect 1462 1632 1514 1652
rect 1462 1600 1492 1632
rect 1492 1600 1514 1632
rect 867 1375 919 1427
rect 867 1294 919 1346
rect 867 1213 919 1265
rect 1329 554 1381 606
rect 1329 490 1381 542
rect 1683 399 1735 451
rect 1749 399 1801 451
rect 969 300 1021 352
rect 969 236 1021 288
rect 865 144 917 196
rect 865 80 917 132
<< metal2 >>
rect 1116 4197 1168 4203
rect 1116 4133 1168 4145
tri 1168 4127 1202 4161 sw
rect 1168 4081 1331 4127
rect 1116 4077 1331 4081
tri 1331 4077 1381 4127 sw
rect 1116 4075 1381 4077
tri 1295 4041 1329 4075 ne
rect 845 3968 851 4020
rect 903 3968 915 4020
rect 967 3968 973 4020
rect 1091 3968 1097 4020
rect 1149 3968 1163 4020
rect 1215 3970 1247 4020
tri 1247 3970 1297 4020 sw
rect 1215 3968 1297 3970
tri 887 3934 921 3968 ne
rect 564 3755 616 3761
rect 564 3691 616 3703
rect 408 3463 414 3515
rect 466 3463 478 3515
rect 530 3463 536 3515
tri 442 3429 476 3463 ne
tri 442 2990 476 3024 se
rect 476 2990 536 3463
rect 419 2938 536 2990
rect 438 2910 444 2938
tri 444 2910 472 2938 nw
tri 438 2904 444 2910 nw
tri 530 2426 564 2460 se
rect 564 2426 616 3639
rect 921 3753 973 3968
tri 1211 3934 1245 3968 ne
rect 921 3689 973 3701
rect 921 3631 973 3637
tri 971 3122 1005 3156 se
rect 1005 3122 1057 3892
rect 1109 3840 1123 3892
rect 1175 3840 1181 3892
tri 1057 3806 1091 3840 nw
rect 929 3070 935 3122
rect 987 3070 999 3122
rect 1051 3070 1057 3122
tri 971 3036 1005 3070 ne
rect 849 2938 855 2990
rect 907 2938 919 2990
rect 971 2938 977 2990
tri 891 2910 919 2938 ne
rect 919 2910 977 2938
tri 919 2904 925 2910 ne
rect 488 2374 494 2426
rect 546 2374 558 2426
rect 610 2374 616 2426
rect 925 1881 977 2910
rect 1005 2608 1057 3070
rect 1101 3616 1217 3622
rect 1101 2824 1217 3500
rect 1153 2772 1165 2824
rect 1101 2756 1217 2772
rect 1153 2704 1165 2756
rect 1101 2688 1217 2704
rect 1153 2636 1165 2688
rect 1101 2630 1217 2636
tri 1057 2608 1065 2616 sw
rect 1005 2594 1065 2608
tri 1005 2534 1065 2594 ne
tri 1065 2534 1139 2608 sw
tri 1065 2460 1139 2534 ne
tri 1139 2460 1213 2534 sw
tri 1139 2438 1161 2460 ne
rect 1005 2374 1011 2426
rect 1063 2374 1075 2426
rect 1127 2374 1133 2426
tri 1047 2342 1079 2374 ne
rect 1079 2342 1133 2374
tri 1079 2340 1081 2342 ne
tri 977 1881 1011 1915 sw
rect 925 1829 931 1881
rect 983 1829 995 1881
rect 1047 1829 1053 1881
rect 1081 1716 1133 2342
rect 1081 1652 1133 1664
rect 1081 1594 1133 1600
rect 842 1427 941 1433
rect 842 1375 867 1427
rect 919 1375 941 1427
rect 842 1346 941 1375
rect 842 1294 867 1346
rect 919 1294 941 1346
rect 842 1265 941 1294
rect 842 1213 867 1265
rect 919 1213 941 1265
rect 842 196 941 1213
rect 1161 399 1213 2460
rect 969 352 1021 358
rect 969 288 1021 300
tri 1021 282 1055 316 sw
tri 1211 282 1245 316 se
rect 1245 282 1297 3968
rect 1329 606 1381 4075
rect 1978 3690 2030 3696
rect 1978 3626 2030 3638
rect 1818 3463 1824 3515
rect 1876 3463 1888 3515
rect 1940 3463 1946 3515
tri 1860 3429 1894 3463 ne
tri 1860 2910 1894 2944 se
rect 1894 2910 1946 3463
rect 1542 2858 1548 2910
rect 1600 2858 1612 2910
rect 1664 2858 1670 2910
rect 1818 2858 1824 2910
rect 1876 2858 1888 2910
rect 1940 2858 1946 2910
tri 1584 2824 1618 2858 ne
rect 1462 2290 1468 2342
rect 1520 2290 1532 2342
rect 1584 2290 1590 2342
rect 1462 1716 1514 2290
tri 1514 2256 1548 2290 nw
tri 1584 1881 1618 1915 se
rect 1618 1881 1670 2858
rect 1978 2342 2030 3574
tri 2030 2342 2064 2376 sw
rect 1978 2290 1984 2342
rect 2036 2290 2048 2342
rect 2100 2290 2106 2342
rect 1542 1829 1548 1881
rect 1600 1829 1612 1881
rect 1664 1829 1670 1881
rect 1462 1652 1514 1664
rect 1462 1594 1514 1600
rect 1329 542 1381 554
rect 1329 484 1381 490
rect 1677 399 1683 451
rect 1735 399 1749 451
rect 1801 399 1807 451
tri 1721 365 1755 399 ne
tri 1297 282 1331 316 sw
rect 1021 270 1352 282
tri 1352 270 1364 282 sw
rect 1021 236 1364 270
rect 969 230 1364 236
tri 1364 230 1404 270 sw
tri 1330 196 1364 230 ne
rect 1364 196 1404 230
tri 1404 196 1438 230 sw
tri 1721 196 1755 230 se
rect 1755 196 1807 399
rect 842 144 865 196
rect 917 144 941 196
tri 1364 144 1416 196 ne
rect 1416 144 1807 196
rect 842 132 941 144
rect 842 80 865 132
rect 917 80 941 132
rect 842 74 941 80
use nfet_CDNS_5595914180817  nfet_CDNS_5595914180817_0
timestamp 1707688321
transform -1 0 1091 0 1 1590
box -79 -32 199 232
use nfet_CDNS_5595914180817  nfet_CDNS_5595914180817_1
timestamp 1707688321
transform 1 0 1503 0 1 1590
box -79 -32 199 232
use nfet_CDNS_5595914180825  nfet_CDNS_5595914180825_0
timestamp 1707688321
transform -1 0 919 0 1 3601
box -79 -32 129 232
use nfet_CDNS_5595914180825  nfet_CDNS_5595914180825_1
timestamp 1707688321
transform 1 0 869 0 -1 4256
box -79 -32 129 232
use pfet_CDNS_5595914180813  pfet_CDNS_5595914180813_0
timestamp 1707688321
transform -1 0 2152 0 1 3554
box -119 -66 239 666
use pfet_CDNS_5595914180813  pfet_CDNS_5595914180813_1
timestamp 1707688321
transform 1 0 442 0 1 3554
box -119 -66 239 666
use pfet_CDNS_5595914180824  pfet_CDNS_5595914180824_0
timestamp 1707688321
transform 1 0 1170 0 -1 4256
box -89 -36 139 236
use pfet_CDNS_5595914180824  pfet_CDNS_5595914180824_1
timestamp 1707688321
transform 1 0 1170 0 -1 3801
box -89 -36 139 236
use sky130_fd_io__amuxsplitv2_switch_levelshifter  sky130_fd_io__amuxsplitv2_switch_levelshifter_0
timestamp 1707688321
transform -1 0 2574 0 1 0
box -28 14 1320 4329
use sky130_fd_io__amuxsplitv2_switch_levelshifter  sky130_fd_io__amuxsplitv2_switch_levelshifter_1
timestamp 1707688321
transform 1 0 20 0 1 0
box -28 14 1320 4329
<< labels >>
flabel metal1 s 163 2464 227 2501 3 FreeSans 200 0 0 0 hold
port 2 nsew
flabel metal1 s 153 3078 231 3113 3 FreeSans 200 0 0 0 in_lv
port 3 nsew
flabel metal1 s 166 2547 257 2581 3 FreeSans 200 0 0 0 reset
port 4 nsew
flabel metal1 s 157 2296 247 2333 3 FreeSans 200 0 0 0 out_h
port 5 nsew
flabel metal1 s 162 2383 247 2418 3 FreeSans 200 0 0 0 out_h_n
port 6 nsew
flabel metal1 s 354 2642 541 2741 3 FreeSans 200 0 0 0 vccd
port 7 nsew
flabel metal1 s 283 4227 405 4264 3 FreeSans 200 0 0 0 vdda
port 8 nsew
flabel metal1 s 507 67 840 155 3 FreeSans 200 0 0 0 vssa
port 9 nsew
flabel metal1 s 2041 4234 2169 4256 3 FreeSans 200 0 0 0 vswitch
port 10 nsew
flabel metal1 s 737 4070 789 4211 3 FreeSans 400 0 0 0 vssd
port 11 nsew
<< properties >>
string GDS_END 729346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 699522
<< end >>
