magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 16604 -12035 22272 -8403
<< nwell >>
rect -401 6562 26385 6864
rect -401 4996 -167 6562
rect 1189 4996 1491 6562
rect -401 4694 1491 4996
rect -401 54 -99 4694
rect 301 3970 1825 4292
rect 301 264 6369 3970
rect 26083 -26 26385 6562
<< pwell >>
rect -73 6182 1129 6490
rect -73 5278 149 6182
rect 907 5278 1129 6182
rect -73 5056 1129 5278
rect 1551 5686 25964 6494
rect 1551 5516 6481 5686
rect 1551 4966 4049 5516
rect 1551 4634 1773 4966
rect 19 4412 1773 4634
rect 19 160 241 4412
rect 19 -62 6651 160
rect 25038 23 25964 5686
rect 25208 -62 25964 23
<< mvpsubdiff >>
rect -47 6430 -23 6464
rect 11 6430 49 6464
rect 83 6430 121 6464
rect 155 6430 193 6464
rect 227 6430 264 6464
rect 298 6430 335 6464
rect 369 6430 406 6464
rect 440 6430 477 6464
rect 511 6430 548 6464
rect 582 6430 619 6464
rect 653 6430 690 6464
rect 724 6430 761 6464
rect 795 6430 832 6464
rect 866 6430 903 6464
rect 937 6430 974 6464
rect 1008 6430 1045 6464
rect 1079 6430 1103 6464
rect -47 6378 1103 6430
rect -47 6344 57 6378
rect 91 6344 126 6378
rect 160 6344 195 6378
rect 229 6344 265 6378
rect 299 6344 335 6378
rect 369 6344 405 6378
rect 439 6344 475 6378
rect 509 6344 545 6378
rect 579 6344 615 6378
rect 649 6344 685 6378
rect 719 6344 755 6378
rect 789 6344 825 6378
rect 859 6344 895 6378
rect 929 6344 965 6378
rect 999 6344 1035 6378
rect 1069 6344 1103 6378
rect -13 6310 1103 6344
rect -47 6276 21 6310
rect 55 6276 91 6310
rect 125 6276 161 6310
rect 195 6276 231 6310
rect 265 6276 301 6310
rect 335 6276 371 6310
rect 405 6276 441 6310
rect 475 6276 511 6310
rect 545 6276 581 6310
rect 615 6276 651 6310
rect 685 6276 721 6310
rect 755 6276 791 6310
rect 825 6276 861 6310
rect 895 6276 931 6310
rect 965 6276 1001 6310
rect 1035 6276 1103 6310
rect -47 6273 1103 6276
rect -13 6272 1103 6273
rect -13 6242 1069 6272
rect -13 6239 89 6242
rect -47 6237 89 6239
rect -47 6203 21 6237
rect 55 6208 89 6237
rect 123 6208 159 6242
rect 193 6208 229 6242
rect 263 6208 299 6242
rect 333 6208 369 6242
rect 403 6208 439 6242
rect 473 6208 509 6242
rect 543 6208 579 6242
rect 613 6208 649 6242
rect 683 6208 720 6242
rect 754 6208 791 6242
rect 825 6208 862 6242
rect 896 6208 933 6242
rect 967 6240 1069 6242
rect 967 6208 1001 6240
rect 55 6203 123 6208
rect -47 6202 123 6203
rect -13 6168 123 6202
rect -47 6164 89 6168
rect -47 6132 21 6164
rect -13 6130 21 6132
rect 55 6134 89 6164
rect 55 6130 123 6134
rect -13 6098 123 6130
rect -47 6094 123 6098
rect -47 6091 89 6094
rect -47 6062 21 6091
rect -13 6057 21 6062
rect 55 6060 89 6091
rect 933 6206 1001 6208
rect 1035 6238 1069 6240
rect 1035 6206 1103 6238
rect 933 6202 1103 6206
rect 933 6172 1069 6202
rect 967 6170 1069 6172
rect 967 6138 1001 6170
rect 933 6136 1001 6138
rect 1035 6168 1069 6170
rect 1035 6136 1103 6168
rect 933 6132 1103 6136
rect 933 6102 1069 6132
rect 55 6057 123 6060
rect -13 6028 123 6057
rect -47 6020 123 6028
rect -47 6018 89 6020
rect -47 5992 21 6018
rect -13 5984 21 5992
rect 55 5986 89 6018
rect 55 5984 123 5986
rect -13 5958 123 5984
rect -47 5946 123 5958
rect -47 5945 89 5946
rect -47 5922 21 5945
rect -13 5911 21 5922
rect 55 5912 89 5945
rect 55 5911 123 5912
rect -13 5888 123 5911
rect -47 5873 123 5888
rect -47 5872 89 5873
rect -47 5852 21 5872
rect -13 5838 21 5852
rect 55 5839 89 5872
rect 55 5838 123 5839
rect -13 5818 123 5838
rect -47 5800 123 5818
rect -47 5799 89 5800
rect -47 5782 21 5799
rect -13 5765 21 5782
rect 55 5766 89 5799
rect 55 5765 123 5766
rect -13 5748 123 5765
rect -47 5727 123 5748
rect -47 5726 89 5727
rect -47 5712 21 5726
rect -13 5692 21 5712
rect 55 5693 89 5726
rect 55 5692 123 5693
rect -13 5678 123 5692
rect -47 5654 123 5678
rect -47 5653 89 5654
rect -47 5642 21 5653
rect -13 5619 21 5642
rect 55 5620 89 5653
rect 55 5619 123 5620
rect -13 5608 123 5619
rect -47 5581 123 5608
rect -47 5580 89 5581
rect -47 5572 21 5580
rect -13 5546 21 5572
rect 55 5547 89 5580
rect 55 5546 123 5547
rect -13 5538 123 5546
rect -47 5508 123 5538
rect -47 5507 89 5508
rect -47 5502 21 5507
rect -13 5473 21 5502
rect 55 5474 89 5507
rect 55 5473 123 5474
rect -13 5468 123 5473
rect -47 5435 123 5468
rect -47 5434 89 5435
rect -47 5432 21 5434
rect -13 5400 21 5432
rect 55 5401 89 5434
rect 55 5400 123 5401
rect -13 5398 123 5400
rect -47 5362 123 5398
rect 967 6100 1069 6102
rect 967 6068 1001 6100
rect 933 6066 1001 6068
rect 1035 6098 1069 6100
rect 1035 6066 1103 6098
rect 933 6062 1103 6066
rect 933 6032 1069 6062
rect 967 6030 1069 6032
rect 967 5998 1001 6030
rect 933 5996 1001 5998
rect 1035 6028 1069 6030
rect 1035 5996 1103 6028
rect 933 5992 1103 5996
rect 933 5962 1069 5992
rect 967 5960 1069 5962
rect 967 5928 1001 5960
rect 933 5926 1001 5928
rect 1035 5958 1069 5960
rect 1035 5926 1103 5958
rect 933 5922 1103 5926
rect 933 5891 1069 5922
rect 967 5890 1069 5891
rect 967 5857 1001 5890
rect 933 5856 1001 5857
rect 1035 5888 1069 5890
rect 1035 5856 1103 5888
rect 933 5852 1103 5856
rect 933 5820 1069 5852
rect 967 5786 1001 5820
rect 1035 5818 1069 5820
rect 1035 5786 1103 5818
rect 933 5782 1103 5786
rect 933 5750 1069 5782
rect 933 5749 1001 5750
rect 967 5716 1001 5749
rect 1035 5748 1069 5750
rect 1035 5716 1103 5748
rect 967 5715 1103 5716
rect 933 5712 1103 5715
rect 933 5680 1069 5712
rect 933 5678 1001 5680
rect 967 5646 1001 5678
rect 1035 5678 1069 5680
rect 1035 5646 1103 5678
rect 967 5644 1103 5646
rect 933 5642 1103 5644
rect 933 5610 1069 5642
rect 933 5607 1001 5610
rect 967 5576 1001 5607
rect 1035 5608 1069 5610
rect 1035 5576 1103 5608
rect 967 5573 1103 5576
rect 933 5572 1103 5573
rect 933 5539 1069 5572
rect 933 5536 1001 5539
rect 967 5505 1001 5536
rect 1035 5538 1069 5539
rect 1035 5505 1103 5538
rect 967 5502 1103 5505
rect 933 5468 1069 5502
rect 933 5465 1001 5468
rect 967 5434 1001 5465
rect 1035 5434 1103 5468
rect 967 5432 1103 5434
rect 967 5431 1069 5432
rect 933 5398 1069 5431
rect 933 5397 1103 5398
rect 933 5394 1001 5397
rect -13 5328 21 5362
rect 55 5328 89 5362
rect -47 5252 123 5328
rect 967 5363 1001 5394
rect 1035 5363 1103 5397
rect 967 5362 1103 5363
rect 967 5360 1069 5362
rect 933 5328 1069 5360
rect 933 5326 1103 5328
rect 933 5323 1001 5326
rect 967 5292 1001 5323
rect 1035 5292 1103 5326
rect 967 5289 1069 5292
rect 933 5258 1069 5289
rect 933 5255 1103 5258
rect 933 5252 1001 5255
rect -47 5218 -23 5252
rect 11 5218 46 5252
rect 80 5218 115 5252
rect 149 5218 184 5252
rect 218 5218 253 5252
rect -47 5184 253 5218
rect -47 5150 -23 5184
rect 11 5150 46 5184
rect 80 5150 115 5184
rect 149 5150 184 5184
rect 218 5150 253 5184
rect 967 5221 1001 5252
rect 1035 5221 1103 5255
rect 967 5187 1069 5221
rect 967 5184 1103 5187
rect 967 5150 1001 5184
rect 1035 5150 1103 5184
rect -47 5116 1069 5150
rect -47 5082 -23 5116
rect 11 5082 48 5116
rect 82 5082 119 5116
rect 153 5082 190 5116
rect 224 5082 261 5116
rect 295 5082 332 5116
rect 366 5082 403 5116
rect 437 5082 473 5116
rect 507 5082 543 5116
rect 577 5082 613 5116
rect 647 5082 683 5116
rect 717 5082 753 5116
rect 787 5082 823 5116
rect 857 5082 893 5116
rect 927 5082 963 5116
rect 997 5082 1103 5116
rect 1577 6460 25938 6468
rect 1577 6426 1601 6460
rect 1635 6426 1670 6460
rect 1704 6426 1739 6460
rect 1773 6426 1808 6460
rect 1842 6426 1877 6460
rect 1911 6426 1946 6460
rect 1980 6426 2015 6460
rect 2049 6426 2084 6460
rect 2118 6426 2153 6460
rect 2187 6426 2222 6460
rect 2256 6426 2291 6460
rect 2325 6426 2360 6460
rect 2394 6426 2429 6460
rect 2463 6426 2498 6460
rect 2532 6426 2567 6460
rect 2601 6426 2636 6460
rect 2670 6426 2705 6460
rect 2739 6426 2774 6460
rect 2808 6426 2843 6460
rect 2877 6426 2912 6460
rect 2946 6426 2981 6460
rect 3015 6426 3050 6460
rect 3084 6426 3119 6460
rect 3153 6426 3188 6460
rect 3222 6426 3257 6460
rect 3291 6426 3326 6460
rect 3360 6426 3395 6460
rect 3429 6426 3464 6460
rect 3498 6426 3533 6460
rect 3567 6426 3602 6460
rect 3636 6426 3671 6460
rect 3705 6426 3740 6460
rect 3774 6426 3809 6460
rect 3843 6426 3878 6460
rect 3912 6426 3947 6460
rect 3981 6426 4016 6460
rect 4050 6426 4085 6460
rect 4119 6426 4154 6460
rect 4188 6426 4223 6460
rect 4257 6426 4292 6460
rect 4326 6426 4361 6460
rect 4395 6426 4430 6460
rect 4464 6426 4499 6460
rect 4533 6426 4568 6460
rect 4602 6426 4637 6460
rect 4671 6426 4706 6460
rect 4740 6426 4775 6460
rect 4809 6426 4844 6460
rect 1577 6392 4844 6426
rect 1577 6358 1601 6392
rect 1635 6358 1670 6392
rect 1704 6358 1739 6392
rect 1773 6358 1808 6392
rect 1842 6358 1877 6392
rect 1911 6358 1946 6392
rect 1980 6358 2015 6392
rect 2049 6358 2084 6392
rect 2118 6358 2153 6392
rect 2187 6358 2222 6392
rect 2256 6358 2291 6392
rect 2325 6358 2360 6392
rect 2394 6358 2429 6392
rect 2463 6358 2498 6392
rect 2532 6358 2567 6392
rect 2601 6358 2636 6392
rect 2670 6358 2705 6392
rect 2739 6358 2774 6392
rect 2808 6358 2843 6392
rect 2877 6358 2912 6392
rect 2946 6358 2981 6392
rect 3015 6358 3050 6392
rect 3084 6358 3119 6392
rect 3153 6358 3188 6392
rect 3222 6358 3257 6392
rect 3291 6358 3326 6392
rect 3360 6358 3395 6392
rect 3429 6358 3464 6392
rect 3498 6358 3533 6392
rect 3567 6358 3602 6392
rect 3636 6358 3671 6392
rect 3705 6358 3740 6392
rect 3774 6358 3809 6392
rect 3843 6358 3878 6392
rect 3912 6358 3947 6392
rect 3981 6358 4016 6392
rect 4050 6358 4085 6392
rect 4119 6358 4154 6392
rect 4188 6358 4223 6392
rect 4257 6358 4292 6392
rect 4326 6358 4361 6392
rect 4395 6358 4430 6392
rect 4464 6358 4499 6392
rect 4533 6358 4568 6392
rect 4602 6358 4637 6392
rect 4671 6358 4706 6392
rect 4740 6358 4775 6392
rect 4809 6358 4844 6392
rect 1577 6324 4844 6358
rect 1577 6290 1601 6324
rect 1635 6290 1670 6324
rect 1704 6290 1739 6324
rect 1773 6290 1808 6324
rect 1842 6290 1877 6324
rect 1911 6290 1946 6324
rect 1980 6290 2015 6324
rect 2049 6290 2084 6324
rect 2118 6290 2153 6324
rect 2187 6290 2222 6324
rect 2256 6290 2291 6324
rect 2325 6290 2360 6324
rect 2394 6290 2429 6324
rect 2463 6290 2498 6324
rect 2532 6290 2567 6324
rect 2601 6290 2636 6324
rect 2670 6290 2705 6324
rect 2739 6290 2774 6324
rect 2808 6290 2843 6324
rect 2877 6290 2912 6324
rect 2946 6290 2981 6324
rect 3015 6290 3050 6324
rect 3084 6290 3119 6324
rect 3153 6290 3188 6324
rect 3222 6290 3257 6324
rect 3291 6290 3326 6324
rect 3360 6290 3395 6324
rect 3429 6290 3464 6324
rect 3498 6290 3533 6324
rect 3567 6290 3602 6324
rect 3636 6290 3671 6324
rect 3705 6290 3740 6324
rect 3774 6290 3809 6324
rect 3843 6290 3878 6324
rect 3912 6290 3947 6324
rect 3981 6290 4016 6324
rect 4050 6290 4085 6324
rect 4119 6290 4154 6324
rect 4188 6290 4223 6324
rect 4257 6290 4292 6324
rect 4326 6290 4361 6324
rect 4395 6290 4430 6324
rect 4464 6290 4499 6324
rect 4533 6290 4568 6324
rect 4602 6290 4637 6324
rect 4671 6290 4706 6324
rect 4740 6290 4775 6324
rect 4809 6290 4844 6324
rect 1577 6256 4844 6290
rect 1577 6222 1601 6256
rect 1635 6222 1670 6256
rect 1704 6222 1739 6256
rect 1773 6222 1808 6256
rect 1842 6222 1877 6256
rect 1911 6222 1946 6256
rect 1980 6222 2015 6256
rect 2049 6222 2084 6256
rect 2118 6222 2153 6256
rect 2187 6222 2222 6256
rect 2256 6222 2291 6256
rect 2325 6222 2360 6256
rect 2394 6222 2429 6256
rect 2463 6222 2498 6256
rect 2532 6222 2567 6256
rect 2601 6222 2636 6256
rect 2670 6222 2705 6256
rect 2739 6222 2774 6256
rect 2808 6222 2843 6256
rect 2877 6222 2912 6256
rect 2946 6222 2981 6256
rect 3015 6222 3050 6256
rect 3084 6222 3119 6256
rect 3153 6222 3188 6256
rect 3222 6222 3257 6256
rect 3291 6222 3326 6256
rect 3360 6222 3395 6256
rect 3429 6222 3464 6256
rect 3498 6222 3533 6256
rect 3567 6222 3602 6256
rect 3636 6222 3671 6256
rect 3705 6222 3740 6256
rect 3774 6222 3809 6256
rect 3843 6222 3878 6256
rect 3912 6222 3947 6256
rect 3981 6222 4016 6256
rect 4050 6222 4085 6256
rect 4119 6222 4154 6256
rect 4188 6222 4223 6256
rect 4257 6222 4292 6256
rect 4326 6222 4361 6256
rect 4395 6222 4430 6256
rect 4464 6222 4499 6256
rect 4533 6222 4568 6256
rect 4602 6222 4637 6256
rect 4671 6222 4706 6256
rect 4740 6222 4775 6256
rect 4809 6222 4844 6256
rect 1577 6188 4844 6222
rect 1577 6154 1601 6188
rect 1635 6154 1670 6188
rect 1704 6154 1739 6188
rect 1773 6154 1808 6188
rect 1842 6154 1877 6188
rect 1911 6154 1946 6188
rect 1980 6154 2015 6188
rect 2049 6154 2084 6188
rect 2118 6154 2153 6188
rect 2187 6154 2222 6188
rect 2256 6154 2291 6188
rect 2325 6154 2360 6188
rect 2394 6154 2429 6188
rect 2463 6154 2498 6188
rect 2532 6154 2567 6188
rect 2601 6154 2636 6188
rect 2670 6154 2705 6188
rect 2739 6154 2774 6188
rect 2808 6154 2843 6188
rect 2877 6154 2912 6188
rect 2946 6154 2981 6188
rect 3015 6154 3050 6188
rect 3084 6154 3119 6188
rect 3153 6154 3188 6188
rect 3222 6154 3257 6188
rect 3291 6154 3326 6188
rect 3360 6154 3395 6188
rect 3429 6154 3464 6188
rect 3498 6154 3533 6188
rect 3567 6154 3602 6188
rect 3636 6154 3671 6188
rect 3705 6154 3740 6188
rect 3774 6154 3809 6188
rect 3843 6154 3878 6188
rect 3912 6154 3947 6188
rect 3981 6154 4016 6188
rect 4050 6154 4085 6188
rect 4119 6154 4154 6188
rect 4188 6154 4223 6188
rect 4257 6154 4292 6188
rect 4326 6154 4361 6188
rect 4395 6154 4430 6188
rect 4464 6154 4499 6188
rect 4533 6154 4568 6188
rect 4602 6154 4637 6188
rect 4671 6154 4706 6188
rect 4740 6154 4775 6188
rect 4809 6154 4844 6188
rect 1577 6120 4844 6154
rect 1577 6086 1601 6120
rect 1635 6086 1670 6120
rect 1704 6086 1739 6120
rect 1773 6086 1808 6120
rect 1842 6086 1877 6120
rect 1911 6086 1946 6120
rect 1980 6086 2015 6120
rect 2049 6086 2084 6120
rect 2118 6086 2153 6120
rect 2187 6086 2222 6120
rect 2256 6086 2291 6120
rect 2325 6086 2360 6120
rect 2394 6086 2429 6120
rect 2463 6086 2498 6120
rect 2532 6086 2567 6120
rect 2601 6086 2636 6120
rect 2670 6086 2705 6120
rect 2739 6086 2774 6120
rect 2808 6086 2843 6120
rect 2877 6086 2912 6120
rect 2946 6086 2981 6120
rect 3015 6086 3050 6120
rect 3084 6086 3119 6120
rect 3153 6086 3188 6120
rect 3222 6086 3257 6120
rect 3291 6086 3326 6120
rect 3360 6086 3395 6120
rect 3429 6086 3464 6120
rect 3498 6086 3533 6120
rect 3567 6086 3602 6120
rect 3636 6086 3671 6120
rect 3705 6086 3740 6120
rect 3774 6086 3809 6120
rect 3843 6086 3878 6120
rect 3912 6086 3947 6120
rect 3981 6086 4016 6120
rect 4050 6086 4085 6120
rect 4119 6086 4154 6120
rect 4188 6086 4223 6120
rect 4257 6086 4292 6120
rect 4326 6086 4361 6120
rect 4395 6086 4430 6120
rect 4464 6086 4499 6120
rect 4533 6086 4568 6120
rect 4602 6086 4637 6120
rect 4671 6086 4706 6120
rect 4740 6086 4775 6120
rect 4809 6086 4844 6120
rect 1577 6052 4844 6086
rect 1577 6018 1601 6052
rect 1635 6018 1670 6052
rect 1704 6018 1739 6052
rect 1773 6018 1808 6052
rect 1842 6018 1877 6052
rect 1911 6018 1946 6052
rect 1980 6018 2015 6052
rect 2049 6018 2084 6052
rect 2118 6018 2153 6052
rect 2187 6018 2222 6052
rect 2256 6018 2291 6052
rect 2325 6018 2360 6052
rect 2394 6018 2429 6052
rect 2463 6018 2498 6052
rect 2532 6018 2567 6052
rect 2601 6018 2636 6052
rect 2670 6018 2705 6052
rect 2739 6018 2774 6052
rect 2808 6018 2843 6052
rect 2877 6018 2912 6052
rect 2946 6018 2981 6052
rect 3015 6018 3050 6052
rect 3084 6018 3119 6052
rect 3153 6018 3188 6052
rect 3222 6018 3257 6052
rect 3291 6018 3326 6052
rect 3360 6018 3395 6052
rect 3429 6018 3464 6052
rect 3498 6018 3533 6052
rect 3567 6018 3602 6052
rect 3636 6018 3671 6052
rect 3705 6018 3740 6052
rect 3774 6018 3809 6052
rect 3843 6018 3878 6052
rect 3912 6018 3947 6052
rect 3981 6018 4016 6052
rect 4050 6018 4085 6052
rect 4119 6018 4154 6052
rect 4188 6018 4223 6052
rect 4257 6018 4292 6052
rect 4326 6018 4361 6052
rect 4395 6018 4430 6052
rect 4464 6018 4499 6052
rect 4533 6018 4568 6052
rect 4602 6018 4637 6052
rect 4671 6018 4706 6052
rect 4740 6018 4775 6052
rect 4809 6018 4844 6052
rect 1577 5984 4844 6018
rect 1577 5950 1601 5984
rect 1635 5950 1670 5984
rect 1704 5950 1739 5984
rect 1773 5950 1808 5984
rect 1842 5950 1877 5984
rect 1911 5950 1946 5984
rect 1980 5950 2015 5984
rect 2049 5950 2084 5984
rect 2118 5950 2153 5984
rect 2187 5950 2222 5984
rect 2256 5950 2291 5984
rect 2325 5950 2360 5984
rect 2394 5950 2429 5984
rect 2463 5950 2498 5984
rect 2532 5950 2567 5984
rect 2601 5950 2636 5984
rect 2670 5950 2705 5984
rect 2739 5950 2774 5984
rect 2808 5950 2843 5984
rect 2877 5950 2912 5984
rect 2946 5950 2981 5984
rect 3015 5950 3050 5984
rect 3084 5950 3119 5984
rect 3153 5950 3188 5984
rect 3222 5950 3257 5984
rect 3291 5950 3326 5984
rect 3360 5950 3395 5984
rect 3429 5950 3464 5984
rect 3498 5950 3533 5984
rect 3567 5950 3602 5984
rect 3636 5950 3671 5984
rect 3705 5950 3740 5984
rect 3774 5950 3809 5984
rect 3843 5950 3878 5984
rect 3912 5950 3947 5984
rect 3981 5950 4016 5984
rect 4050 5950 4085 5984
rect 4119 5950 4154 5984
rect 4188 5950 4223 5984
rect 4257 5950 4292 5984
rect 4326 5950 4361 5984
rect 4395 5950 4430 5984
rect 4464 5950 4499 5984
rect 4533 5950 4568 5984
rect 4602 5950 4637 5984
rect 4671 5950 4706 5984
rect 4740 5950 4775 5984
rect 4809 5950 4844 5984
rect 1577 5916 4844 5950
rect 1577 5882 1601 5916
rect 1635 5882 1670 5916
rect 1704 5882 1739 5916
rect 1773 5882 1808 5916
rect 1842 5882 1877 5916
rect 1911 5882 1946 5916
rect 1980 5882 2015 5916
rect 2049 5882 2084 5916
rect 2118 5882 2153 5916
rect 2187 5882 2222 5916
rect 2256 5882 2291 5916
rect 2325 5882 2360 5916
rect 2394 5882 2429 5916
rect 2463 5882 2498 5916
rect 2532 5882 2567 5916
rect 2601 5882 2636 5916
rect 2670 5882 2705 5916
rect 2739 5882 2774 5916
rect 2808 5882 2843 5916
rect 2877 5882 2912 5916
rect 2946 5882 2981 5916
rect 3015 5882 3050 5916
rect 3084 5882 3119 5916
rect 3153 5882 3188 5916
rect 3222 5882 3257 5916
rect 3291 5882 3326 5916
rect 3360 5882 3395 5916
rect 3429 5882 3464 5916
rect 3498 5882 3533 5916
rect 3567 5882 3602 5916
rect 3636 5882 3671 5916
rect 3705 5882 3740 5916
rect 3774 5882 3809 5916
rect 3843 5882 3878 5916
rect 3912 5882 3947 5916
rect 3981 5882 4016 5916
rect 4050 5882 4085 5916
rect 4119 5882 4154 5916
rect 4188 5882 4223 5916
rect 4257 5882 4292 5916
rect 4326 5882 4361 5916
rect 4395 5882 4430 5916
rect 4464 5882 4499 5916
rect 4533 5882 4568 5916
rect 4602 5882 4637 5916
rect 4671 5882 4706 5916
rect 4740 5882 4775 5916
rect 4809 5882 4844 5916
rect 1577 5848 4844 5882
rect 1577 5814 1601 5848
rect 1635 5814 1670 5848
rect 1704 5814 1739 5848
rect 1773 5814 1808 5848
rect 1842 5814 1877 5848
rect 1911 5814 1946 5848
rect 1980 5814 2015 5848
rect 2049 5814 2084 5848
rect 2118 5814 2153 5848
rect 2187 5814 2222 5848
rect 2256 5814 2291 5848
rect 2325 5814 2360 5848
rect 2394 5814 2429 5848
rect 2463 5814 2498 5848
rect 2532 5814 2567 5848
rect 2601 5814 2636 5848
rect 2670 5814 2705 5848
rect 2739 5814 2774 5848
rect 2808 5814 2843 5848
rect 2877 5814 2912 5848
rect 2946 5814 2981 5848
rect 3015 5814 3050 5848
rect 3084 5814 3119 5848
rect 3153 5814 3188 5848
rect 3222 5814 3257 5848
rect 3291 5814 3326 5848
rect 3360 5814 3395 5848
rect 3429 5814 3464 5848
rect 3498 5814 3533 5848
rect 3567 5814 3602 5848
rect 3636 5814 3671 5848
rect 3705 5814 3740 5848
rect 3774 5814 3809 5848
rect 3843 5814 3878 5848
rect 3912 5814 3947 5848
rect 3981 5814 4016 5848
rect 4050 5814 4085 5848
rect 4119 5814 4154 5848
rect 4188 5814 4223 5848
rect 4257 5814 4292 5848
rect 4326 5814 4361 5848
rect 4395 5814 4430 5848
rect 4464 5814 4499 5848
rect 4533 5814 4568 5848
rect 4602 5814 4637 5848
rect 4671 5814 4706 5848
rect 4740 5814 4775 5848
rect 4809 5814 4844 5848
rect 1577 5780 4844 5814
rect 1577 5746 1601 5780
rect 1635 5746 1670 5780
rect 1704 5746 1739 5780
rect 1773 5746 1808 5780
rect 1842 5746 1877 5780
rect 1911 5746 1946 5780
rect 1980 5746 2015 5780
rect 2049 5746 2084 5780
rect 2118 5746 2153 5780
rect 2187 5746 2222 5780
rect 2256 5746 2291 5780
rect 2325 5746 2360 5780
rect 2394 5746 2429 5780
rect 2463 5746 2498 5780
rect 2532 5746 2567 5780
rect 2601 5746 2636 5780
rect 2670 5746 2705 5780
rect 2739 5746 2774 5780
rect 2808 5746 2843 5780
rect 2877 5746 2912 5780
rect 2946 5746 2981 5780
rect 3015 5746 3050 5780
rect 3084 5746 3119 5780
rect 3153 5746 3188 5780
rect 3222 5746 3257 5780
rect 3291 5746 3326 5780
rect 3360 5746 3395 5780
rect 3429 5746 3464 5780
rect 3498 5746 3533 5780
rect 3567 5746 3602 5780
rect 3636 5746 3671 5780
rect 3705 5746 3740 5780
rect 3774 5746 3809 5780
rect 3843 5746 3878 5780
rect 3912 5746 3947 5780
rect 3981 5746 4016 5780
rect 4050 5746 4085 5780
rect 4119 5746 4154 5780
rect 4188 5746 4223 5780
rect 4257 5746 4292 5780
rect 4326 5746 4361 5780
rect 4395 5746 4430 5780
rect 4464 5746 4499 5780
rect 4533 5746 4568 5780
rect 4602 5746 4637 5780
rect 4671 5746 4706 5780
rect 4740 5746 4775 5780
rect 4809 5746 4844 5780
rect 25210 6444 25938 6460
rect 25210 5746 25268 6444
rect 1577 5712 4844 5746
rect 6421 5712 25268 5746
rect 1577 5678 1611 5712
rect 1645 5678 1681 5712
rect 1715 5678 1751 5712
rect 1785 5678 1821 5712
rect 1855 5678 1891 5712
rect 1925 5678 1961 5712
rect 1995 5678 2030 5712
rect 2064 5678 2099 5712
rect 2133 5678 2168 5712
rect 2202 5678 2237 5712
rect 2271 5678 2306 5712
rect 2340 5678 2375 5712
rect 1577 5644 2375 5678
rect 1577 5610 1645 5644
rect 1679 5610 1718 5644
rect 1752 5610 1791 5644
rect 1825 5610 1864 5644
rect 1898 5610 1937 5644
rect 1971 5610 2010 5644
rect 2044 5610 2083 5644
rect 2117 5610 2156 5644
rect 2190 5610 2229 5644
rect 2263 5610 2302 5644
rect 2336 5610 2375 5644
rect 1577 5604 2375 5610
rect 1611 5576 2375 5604
rect 1611 5575 1713 5576
rect 1611 5570 1645 5575
rect 1577 5541 1645 5570
rect 1679 5542 1713 5575
rect 1747 5542 1787 5576
rect 1821 5542 1861 5576
rect 1895 5542 1935 5576
rect 1969 5542 2009 5576
rect 2043 5542 2083 5576
rect 2117 5542 2156 5576
rect 2190 5542 2229 5576
rect 2263 5542 2302 5576
rect 2336 5542 2375 5576
rect 6421 5542 6455 5712
rect 25064 5612 25149 5627
rect 1679 5541 4023 5542
rect 1577 5533 4023 5541
rect 1611 5506 4023 5533
rect 1611 5499 1645 5506
rect 1577 5472 1645 5499
rect 1679 5505 4023 5506
rect 1679 5472 1713 5505
rect 1577 5471 1713 5472
rect 1747 5471 1781 5505
rect 1815 5471 1850 5505
rect 1884 5471 1919 5505
rect 1953 5471 1988 5505
rect 2022 5471 2057 5505
rect 2091 5471 2126 5505
rect 2160 5471 2195 5505
rect 2229 5471 2264 5505
rect 2298 5471 2333 5505
rect 1577 5462 2333 5471
rect 1611 5437 2333 5462
rect 1611 5428 1645 5437
rect 1577 5403 1645 5428
rect 1679 5434 1781 5437
rect 1679 5403 1713 5434
rect 1577 5400 1713 5403
rect 1747 5403 1781 5434
rect 1815 5403 1850 5437
rect 1884 5403 1919 5437
rect 1953 5403 1988 5437
rect 2022 5403 2057 5437
rect 2091 5403 2126 5437
rect 2160 5403 2195 5437
rect 2229 5403 2264 5437
rect 2298 5403 2333 5437
rect 1747 5400 2333 5403
rect 1577 5391 2333 5400
rect 1611 5369 2333 5391
rect 1611 5368 1781 5369
rect 1611 5357 1645 5368
rect 1577 5334 1645 5357
rect 1679 5363 1781 5368
rect 1679 5334 1713 5363
rect 1577 5329 1713 5334
rect 1747 5335 1781 5363
rect 1815 5335 1850 5369
rect 1884 5335 1919 5369
rect 1953 5335 1988 5369
rect 2022 5335 2057 5369
rect 2091 5335 2126 5369
rect 2160 5335 2195 5369
rect 2229 5335 2264 5369
rect 2298 5335 2333 5369
rect 1747 5329 2333 5335
rect 1577 5320 2333 5329
rect 1611 5301 2333 5320
rect 1611 5299 1781 5301
rect 1611 5286 1645 5299
rect 1577 5265 1645 5286
rect 1679 5292 1781 5299
rect 1679 5265 1713 5292
rect 1577 5258 1713 5265
rect 1747 5267 1781 5292
rect 1815 5267 1850 5301
rect 1884 5267 1919 5301
rect 1953 5267 1988 5301
rect 2022 5267 2057 5301
rect 2091 5267 2126 5301
rect 2160 5267 2195 5301
rect 2229 5267 2264 5301
rect 2298 5267 2333 5301
rect 1747 5258 2333 5267
rect 1577 5249 2333 5258
rect 1611 5233 2333 5249
rect 1611 5230 1781 5233
rect 1611 5215 1645 5230
rect 1577 5196 1645 5215
rect 1679 5221 1781 5230
rect 1679 5196 1713 5221
rect 1577 5187 1713 5196
rect 1747 5199 1781 5221
rect 1815 5199 1850 5233
rect 1884 5199 1919 5233
rect 1953 5199 1988 5233
rect 2022 5199 2057 5233
rect 2091 5199 2126 5233
rect 2160 5199 2195 5233
rect 2229 5199 2264 5233
rect 2298 5199 2333 5233
rect 1747 5187 2333 5199
rect 1577 5178 2333 5187
rect 1611 5165 2333 5178
rect 1611 5161 1781 5165
rect 1611 5144 1645 5161
rect 1577 5127 1645 5144
rect 1679 5150 1781 5161
rect 1679 5127 1713 5150
rect 1577 5116 1713 5127
rect 1747 5131 1781 5150
rect 1815 5131 1850 5165
rect 1884 5131 1919 5165
rect 1953 5131 1988 5165
rect 2022 5131 2057 5165
rect 2091 5131 2126 5165
rect 2160 5131 2195 5165
rect 2229 5131 2264 5165
rect 2298 5131 2333 5165
rect 1747 5116 2333 5131
rect 1577 5107 2333 5116
rect 1611 5097 2333 5107
rect 1611 5092 1781 5097
rect 1611 5073 1645 5092
rect 1577 5058 1645 5073
rect 1679 5079 1781 5092
rect 1679 5058 1713 5079
rect 1577 5045 1713 5058
rect 1747 5063 1781 5079
rect 1815 5063 1850 5097
rect 1884 5063 1919 5097
rect 1953 5063 1988 5097
rect 2022 5063 2057 5097
rect 2091 5063 2126 5097
rect 2160 5063 2195 5097
rect 2229 5063 2264 5097
rect 2298 5063 2333 5097
rect 1747 5045 2333 5063
rect 1577 5036 2333 5045
rect 1611 5029 2333 5036
rect 1611 5023 1781 5029
rect 1611 5002 1645 5023
rect 1577 4989 1645 5002
rect 1679 5008 1781 5023
rect 1679 4989 1713 5008
rect 1577 4974 1713 4989
rect 1747 4995 1781 5008
rect 1815 4995 1850 5029
rect 1884 4995 1919 5029
rect 1953 4995 1988 5029
rect 2022 4995 2057 5029
rect 2091 4995 2126 5029
rect 2160 4995 2195 5029
rect 2229 4995 2264 5029
rect 2298 4995 2333 5029
rect 3999 4995 4023 5505
rect 1747 4992 4023 4995
rect 1577 4965 1747 4974
rect 1611 4954 1747 4965
rect 1611 4931 1645 4954
rect 1577 4920 1645 4931
rect 1679 4937 1747 4954
rect 1679 4920 1713 4937
rect 1577 4903 1713 4920
rect 1577 4894 1747 4903
rect 1611 4885 1747 4894
rect 1611 4860 1645 4885
rect 1577 4851 1645 4860
rect 1679 4866 1747 4885
rect 1679 4851 1713 4866
rect 1577 4832 1713 4851
rect 1577 4823 1747 4832
rect 1611 4816 1747 4823
rect 1611 4789 1645 4816
rect 1577 4782 1645 4789
rect 1679 4794 1747 4816
rect 1679 4782 1713 4794
rect 1577 4760 1713 4782
rect 1577 4752 1747 4760
rect 1611 4747 1747 4752
rect 1611 4718 1645 4747
rect 1577 4713 1645 4718
rect 1679 4722 1747 4747
rect 1679 4713 1713 4722
rect 1577 4688 1713 4713
rect 1577 4680 1747 4688
rect 1611 4678 1747 4680
rect 1611 4646 1645 4678
rect 1577 4644 1645 4646
rect 1679 4650 1747 4678
rect 1679 4644 1713 4650
rect 1577 4616 1713 4644
rect 1577 4609 1747 4616
rect 1577 4608 1645 4609
rect 45 4574 79 4608
rect 113 4574 150 4608
rect 184 4574 220 4608
rect 254 4574 290 4608
rect 324 4574 360 4608
rect 394 4574 430 4608
rect 464 4574 500 4608
rect 534 4574 570 4608
rect 604 4574 640 4608
rect 674 4574 710 4608
rect 744 4574 780 4608
rect 814 4574 850 4608
rect 884 4574 920 4608
rect 954 4574 990 4608
rect 1024 4574 1060 4608
rect 1094 4574 1130 4608
rect 1164 4574 1200 4608
rect 1234 4574 1282 4608
rect 1316 4574 1356 4608
rect 1390 4574 1430 4608
rect 1464 4574 1504 4608
rect 1538 4574 1577 4608
rect 1611 4575 1645 4608
rect 1679 4578 1747 4609
rect 1679 4575 1713 4578
rect 1611 4574 1713 4575
rect 45 4544 1713 4574
rect 45 4540 1747 4544
rect 45 4506 113 4540
rect 147 4506 186 4540
rect 220 4506 259 4540
rect 293 4506 332 4540
rect 366 4506 405 4540
rect 439 4506 478 4540
rect 512 4506 551 4540
rect 585 4506 624 4540
rect 658 4506 696 4540
rect 730 4506 768 4540
rect 802 4506 840 4540
rect 874 4506 912 4540
rect 946 4506 984 4540
rect 1018 4506 1056 4540
rect 1090 4506 1128 4540
rect 1162 4506 1200 4540
rect 1234 4506 1282 4540
rect 1316 4506 1355 4540
rect 1389 4506 1428 4540
rect 1462 4506 1501 4540
rect 1535 4506 1573 4540
rect 1607 4506 1645 4540
rect 1679 4506 1747 4540
rect 147 4472 1713 4506
rect 215 4438 254 4472
rect 288 4438 327 4472
rect 361 4438 400 4472
rect 434 4438 473 4472
rect 507 4438 546 4472
rect 580 4438 619 4472
rect 653 4438 692 4472
rect 726 4438 765 4472
rect 799 4438 838 4472
rect 872 4438 911 4472
rect 945 4438 984 4472
rect 1018 4438 1056 4472
rect 1090 4438 1128 4472
rect 1162 4438 1200 4472
rect 1234 4438 1282 4472
rect 1316 4438 1360 4472
rect 1394 4438 1438 4472
rect 1472 4438 1516 4472
rect 1550 4438 1593 4472
rect 1627 4438 1747 4472
rect 79 3860 215 3894
rect 45 3859 215 3860
rect 45 3826 113 3859
rect 79 3825 113 3826
rect 147 3825 181 3859
rect 79 3792 215 3825
rect 45 3790 215 3792
rect 45 3758 113 3790
rect 79 3756 113 3758
rect 147 3756 181 3790
rect 79 3724 215 3756
rect 45 3721 215 3724
rect 45 3690 113 3721
rect 79 3687 113 3690
rect 147 3687 181 3721
rect 79 3656 215 3687
rect 45 3652 215 3656
rect 45 3622 113 3652
rect 79 3618 113 3622
rect 147 3618 181 3652
rect 79 3588 215 3618
rect 45 3583 215 3588
rect 45 3554 113 3583
rect 79 3549 113 3554
rect 147 3549 181 3583
rect 79 3520 215 3549
rect 45 3514 215 3520
rect 45 3486 113 3514
rect 79 3480 113 3486
rect 147 3480 181 3514
rect 79 3452 215 3480
rect 45 3445 215 3452
rect 45 3418 113 3445
rect 79 3411 113 3418
rect 147 3411 181 3445
rect 79 3384 215 3411
rect 45 3376 215 3384
rect 45 3350 113 3376
rect 79 3342 113 3350
rect 147 3342 181 3376
rect 79 3316 215 3342
rect 45 3307 215 3316
rect 45 3282 113 3307
rect 79 3273 113 3282
rect 147 3273 181 3307
rect 79 3248 215 3273
rect 45 3238 215 3248
rect 45 3214 113 3238
rect 79 3204 113 3214
rect 147 3204 181 3238
rect 79 3180 215 3204
rect 45 3169 215 3180
rect 45 3146 113 3169
rect 79 3135 113 3146
rect 147 3135 181 3169
rect 79 3112 215 3135
rect 45 3100 215 3112
rect 45 3078 113 3100
rect 79 3066 113 3078
rect 147 3066 181 3100
rect 79 3044 215 3066
rect 45 3031 215 3044
rect 45 3010 113 3031
rect 79 2997 113 3010
rect 147 2997 181 3031
rect 79 2976 215 2997
rect 45 2962 215 2976
rect 45 2942 113 2962
rect 79 2928 113 2942
rect 147 2928 181 2962
rect 79 2908 215 2928
rect 45 2893 215 2908
rect 45 2874 113 2893
rect 79 2859 113 2874
rect 147 2859 181 2893
rect 79 2840 215 2859
rect 45 2824 215 2840
rect 45 2806 113 2824
rect 79 2790 113 2806
rect 147 2790 181 2824
rect 79 2772 215 2790
rect 45 2755 215 2772
rect 45 2738 113 2755
rect 79 2721 113 2738
rect 147 2721 181 2755
rect 79 2704 215 2721
rect 45 2686 215 2704
rect 45 2670 113 2686
rect 79 2652 113 2670
rect 147 2652 181 2686
rect 79 2636 215 2652
rect 45 2617 215 2636
rect 45 2602 113 2617
rect 79 2583 113 2602
rect 147 2583 181 2617
rect 79 2568 215 2583
rect 45 2548 215 2568
rect 45 2534 113 2548
rect 79 2514 113 2534
rect 147 2514 181 2548
rect 79 2500 215 2514
rect 45 2479 215 2500
rect 45 2466 113 2479
rect 79 2445 113 2466
rect 147 2445 181 2479
rect 79 2432 215 2445
rect 45 2410 215 2432
rect 45 2398 113 2410
rect 79 2376 113 2398
rect 147 2376 181 2410
rect 79 2364 215 2376
rect 45 2341 215 2364
rect 45 2330 113 2341
rect 79 2307 113 2330
rect 147 2307 181 2341
rect 79 2296 215 2307
rect 45 2272 215 2296
rect 45 2262 113 2272
rect 79 2238 113 2262
rect 147 2238 181 2272
rect 79 2228 215 2238
rect 45 2203 215 2228
rect 45 2194 113 2203
rect 79 2169 113 2194
rect 147 2169 181 2203
rect 79 2160 215 2169
rect 45 2134 215 2160
rect 45 2126 113 2134
rect 79 2100 113 2126
rect 147 2100 181 2134
rect 79 2092 215 2100
rect 45 2065 215 2092
rect 45 2058 113 2065
rect 79 2031 113 2058
rect 147 2031 181 2065
rect 79 2024 215 2031
rect 45 1996 215 2024
rect 45 1990 113 1996
rect 79 1962 113 1990
rect 147 1962 181 1996
rect 79 1956 215 1962
rect 45 1927 215 1956
rect 45 1922 113 1927
rect 79 1893 113 1922
rect 147 1893 181 1927
rect 79 1888 215 1893
rect 45 1858 215 1888
rect 45 1854 113 1858
rect 79 1824 113 1854
rect 147 1824 181 1858
rect 79 1820 215 1824
rect 45 1789 215 1820
rect 45 1786 113 1789
rect 79 1755 113 1786
rect 147 1755 181 1789
rect 79 1752 215 1755
rect 45 1720 215 1752
rect 45 1718 113 1720
rect 79 1686 113 1718
rect 147 1686 181 1720
rect 79 1684 215 1686
rect 45 1651 215 1684
rect 45 1650 113 1651
rect 79 1617 113 1650
rect 147 1617 181 1651
rect 79 1616 215 1617
rect 45 1582 215 1616
rect 79 1548 113 1582
rect 147 1548 181 1582
rect 45 1513 215 1548
rect 79 1479 113 1513
rect 147 1479 181 1513
rect 45 1444 215 1479
rect 79 1410 113 1444
rect 147 1410 181 1444
rect 45 1375 215 1410
rect 79 1341 113 1375
rect 147 1341 181 1375
rect 45 1306 215 1341
rect 79 1272 113 1306
rect 147 1272 181 1306
rect 45 1237 215 1272
rect 79 1203 113 1237
rect 147 1203 181 1237
rect 45 1168 215 1203
rect 79 1134 113 1168
rect 147 1134 181 1168
rect 45 1099 215 1134
rect 79 1065 113 1099
rect 147 1065 181 1099
rect 45 1030 215 1065
rect 79 996 113 1030
rect 147 996 181 1030
rect 45 961 215 996
rect 79 927 113 961
rect 147 927 181 961
rect 45 892 215 927
rect 79 858 113 892
rect 147 858 181 892
rect 45 823 215 858
rect 79 789 113 823
rect 147 789 181 823
rect 45 754 215 789
rect 79 720 113 754
rect 147 720 181 754
rect 45 685 215 720
rect 79 651 113 685
rect 147 651 181 685
rect 45 616 215 651
rect 79 582 113 616
rect 147 582 181 616
rect 45 547 215 582
rect 79 513 113 547
rect 147 513 181 547
rect 45 478 215 513
rect 79 444 113 478
rect 147 444 181 478
rect 45 409 215 444
rect 79 375 113 409
rect 147 375 181 409
rect 45 340 215 375
rect 79 306 113 340
rect 147 306 181 340
rect 45 271 215 306
rect 79 237 113 271
rect 147 237 181 271
rect 45 202 215 237
rect 79 168 113 202
rect 147 168 181 202
rect 45 134 215 168
rect 45 -36 6625 134
rect 25134 49 25149 5612
rect 25234 2058 25268 5712
rect 25914 2058 25938 6444
rect 25234 2023 25938 2058
rect 25234 1989 25268 2023
rect 25302 1989 25336 2023
rect 25370 1989 25404 2023
rect 25438 1989 25472 2023
rect 25506 1989 25540 2023
rect 25574 1989 25608 2023
rect 25642 1989 25676 2023
rect 25710 1989 25744 2023
rect 25778 1989 25812 2023
rect 25846 1989 25880 2023
rect 25914 1989 25938 2023
rect 25234 1954 25938 1989
rect 25234 1920 25268 1954
rect 25302 1920 25336 1954
rect 25370 1920 25404 1954
rect 25438 1920 25472 1954
rect 25506 1920 25540 1954
rect 25574 1920 25608 1954
rect 25642 1920 25676 1954
rect 25710 1920 25744 1954
rect 25778 1920 25812 1954
rect 25846 1920 25880 1954
rect 25914 1920 25938 1954
rect 25234 1885 25938 1920
rect 25234 1851 25268 1885
rect 25302 1851 25336 1885
rect 25370 1851 25404 1885
rect 25438 1851 25472 1885
rect 25506 1851 25540 1885
rect 25574 1851 25608 1885
rect 25642 1851 25676 1885
rect 25710 1851 25744 1885
rect 25778 1851 25812 1885
rect 25846 1851 25880 1885
rect 25914 1851 25938 1885
rect 25234 1816 25938 1851
rect 25234 1782 25268 1816
rect 25302 1782 25336 1816
rect 25370 1782 25404 1816
rect 25438 1782 25472 1816
rect 25506 1782 25540 1816
rect 25574 1782 25608 1816
rect 25642 1782 25676 1816
rect 25710 1782 25744 1816
rect 25778 1782 25812 1816
rect 25846 1782 25880 1816
rect 25914 1782 25938 1816
rect 25234 1747 25938 1782
rect 25234 1713 25268 1747
rect 25302 1713 25336 1747
rect 25370 1713 25404 1747
rect 25438 1713 25472 1747
rect 25506 1713 25540 1747
rect 25574 1713 25608 1747
rect 25642 1713 25676 1747
rect 25710 1713 25744 1747
rect 25778 1713 25812 1747
rect 25846 1713 25880 1747
rect 25914 1713 25938 1747
rect 25234 1678 25938 1713
rect 25234 1644 25268 1678
rect 25302 1644 25336 1678
rect 25370 1644 25404 1678
rect 25438 1644 25472 1678
rect 25506 1644 25540 1678
rect 25574 1644 25608 1678
rect 25642 1644 25676 1678
rect 25710 1644 25744 1678
rect 25778 1644 25812 1678
rect 25846 1644 25880 1678
rect 25914 1644 25938 1678
rect 25234 1609 25938 1644
rect 25234 1575 25268 1609
rect 25302 1575 25336 1609
rect 25370 1575 25404 1609
rect 25438 1575 25472 1609
rect 25506 1575 25540 1609
rect 25574 1575 25608 1609
rect 25642 1575 25676 1609
rect 25710 1575 25744 1609
rect 25778 1575 25812 1609
rect 25846 1575 25880 1609
rect 25914 1575 25938 1609
rect 25234 1540 25938 1575
rect 25234 1506 25268 1540
rect 25302 1506 25336 1540
rect 25370 1506 25404 1540
rect 25438 1506 25472 1540
rect 25506 1506 25540 1540
rect 25574 1506 25608 1540
rect 25642 1506 25676 1540
rect 25710 1506 25744 1540
rect 25778 1506 25812 1540
rect 25846 1506 25880 1540
rect 25914 1506 25938 1540
rect 25234 1471 25938 1506
rect 25234 1437 25268 1471
rect 25302 1437 25336 1471
rect 25370 1437 25404 1471
rect 25438 1437 25472 1471
rect 25506 1437 25540 1471
rect 25574 1437 25608 1471
rect 25642 1437 25676 1471
rect 25710 1437 25744 1471
rect 25778 1437 25812 1471
rect 25846 1437 25880 1471
rect 25914 1437 25938 1471
rect 25234 1402 25938 1437
rect 25234 1368 25268 1402
rect 25302 1368 25336 1402
rect 25370 1368 25404 1402
rect 25438 1368 25472 1402
rect 25506 1368 25540 1402
rect 25574 1368 25608 1402
rect 25642 1368 25676 1402
rect 25710 1368 25744 1402
rect 25778 1368 25812 1402
rect 25846 1368 25880 1402
rect 25914 1368 25938 1402
rect 25234 1333 25938 1368
rect 25234 1299 25268 1333
rect 25302 1299 25336 1333
rect 25370 1299 25404 1333
rect 25438 1299 25472 1333
rect 25506 1299 25540 1333
rect 25574 1299 25608 1333
rect 25642 1299 25676 1333
rect 25710 1299 25744 1333
rect 25778 1299 25812 1333
rect 25846 1299 25880 1333
rect 25914 1299 25938 1333
rect 25234 1264 25938 1299
rect 25234 1230 25268 1264
rect 25302 1230 25336 1264
rect 25370 1230 25404 1264
rect 25438 1230 25472 1264
rect 25506 1230 25540 1264
rect 25574 1230 25608 1264
rect 25642 1230 25676 1264
rect 25710 1230 25744 1264
rect 25778 1230 25812 1264
rect 25846 1230 25880 1264
rect 25914 1230 25938 1264
rect 25234 1195 25938 1230
rect 25234 1161 25268 1195
rect 25302 1161 25336 1195
rect 25370 1161 25404 1195
rect 25438 1161 25472 1195
rect 25506 1161 25540 1195
rect 25574 1161 25608 1195
rect 25642 1161 25676 1195
rect 25710 1161 25744 1195
rect 25778 1161 25812 1195
rect 25846 1161 25880 1195
rect 25914 1161 25938 1195
rect 25234 1126 25938 1161
rect 25234 1092 25268 1126
rect 25302 1092 25336 1126
rect 25370 1092 25404 1126
rect 25438 1092 25472 1126
rect 25506 1092 25540 1126
rect 25574 1092 25608 1126
rect 25642 1092 25676 1126
rect 25710 1092 25744 1126
rect 25778 1092 25812 1126
rect 25846 1092 25880 1126
rect 25914 1092 25938 1126
rect 25234 1057 25938 1092
rect 25234 1023 25268 1057
rect 25302 1023 25336 1057
rect 25370 1023 25404 1057
rect 25438 1023 25472 1057
rect 25506 1023 25540 1057
rect 25574 1023 25608 1057
rect 25642 1023 25676 1057
rect 25710 1023 25744 1057
rect 25778 1023 25812 1057
rect 25846 1023 25880 1057
rect 25914 1023 25938 1057
rect 25234 988 25938 1023
rect 25234 954 25268 988
rect 25302 954 25336 988
rect 25370 954 25404 988
rect 25438 954 25472 988
rect 25506 954 25540 988
rect 25574 954 25608 988
rect 25642 954 25676 988
rect 25710 954 25744 988
rect 25778 954 25812 988
rect 25846 954 25880 988
rect 25914 954 25938 988
rect 25234 919 25938 954
rect 25234 885 25268 919
rect 25302 885 25336 919
rect 25370 885 25404 919
rect 25438 885 25472 919
rect 25506 885 25540 919
rect 25574 885 25608 919
rect 25642 885 25676 919
rect 25710 885 25744 919
rect 25778 885 25812 919
rect 25846 885 25880 919
rect 25914 885 25938 919
rect 25234 850 25938 885
rect 25234 816 25268 850
rect 25302 816 25336 850
rect 25370 816 25404 850
rect 25438 816 25472 850
rect 25506 816 25540 850
rect 25574 816 25608 850
rect 25642 816 25676 850
rect 25710 816 25744 850
rect 25778 816 25812 850
rect 25846 816 25880 850
rect 25914 816 25938 850
rect 25234 781 25938 816
rect 25234 747 25268 781
rect 25302 747 25336 781
rect 25370 747 25404 781
rect 25438 747 25472 781
rect 25506 747 25540 781
rect 25574 747 25608 781
rect 25642 747 25676 781
rect 25710 747 25744 781
rect 25778 747 25812 781
rect 25846 747 25880 781
rect 25914 747 25938 781
rect 25234 712 25938 747
rect 25234 678 25268 712
rect 25302 678 25336 712
rect 25370 678 25404 712
rect 25438 678 25472 712
rect 25506 678 25540 712
rect 25574 678 25608 712
rect 25642 678 25676 712
rect 25710 678 25744 712
rect 25778 678 25812 712
rect 25846 678 25880 712
rect 25914 678 25938 712
rect 25234 643 25938 678
rect 25234 609 25268 643
rect 25302 609 25336 643
rect 25370 609 25404 643
rect 25438 609 25472 643
rect 25506 609 25540 643
rect 25574 609 25608 643
rect 25642 609 25676 643
rect 25710 609 25744 643
rect 25778 609 25812 643
rect 25846 609 25880 643
rect 25914 609 25938 643
rect 25234 574 25938 609
rect 25234 540 25268 574
rect 25302 540 25336 574
rect 25370 540 25404 574
rect 25438 540 25472 574
rect 25506 540 25540 574
rect 25574 540 25608 574
rect 25642 540 25676 574
rect 25710 540 25744 574
rect 25778 540 25812 574
rect 25846 540 25880 574
rect 25914 540 25938 574
rect 25234 505 25938 540
rect 25234 471 25268 505
rect 25302 471 25336 505
rect 25370 471 25404 505
rect 25438 471 25472 505
rect 25506 471 25540 505
rect 25574 471 25608 505
rect 25642 471 25676 505
rect 25710 471 25744 505
rect 25778 471 25812 505
rect 25846 471 25880 505
rect 25914 471 25938 505
rect 25234 436 25938 471
rect 25234 402 25268 436
rect 25302 402 25336 436
rect 25370 402 25404 436
rect 25438 402 25472 436
rect 25506 402 25540 436
rect 25574 402 25608 436
rect 25642 402 25676 436
rect 25710 402 25744 436
rect 25778 402 25812 436
rect 25846 402 25880 436
rect 25914 402 25938 436
rect 25234 367 25938 402
rect 25234 333 25268 367
rect 25302 333 25336 367
rect 25370 333 25404 367
rect 25438 333 25472 367
rect 25506 333 25540 367
rect 25574 333 25608 367
rect 25642 333 25676 367
rect 25710 333 25744 367
rect 25778 333 25812 367
rect 25846 333 25880 367
rect 25914 333 25938 367
rect 25234 298 25938 333
rect 25234 264 25268 298
rect 25302 264 25336 298
rect 25370 264 25404 298
rect 25438 264 25472 298
rect 25506 264 25540 298
rect 25574 264 25608 298
rect 25642 264 25676 298
rect 25710 264 25744 298
rect 25778 264 25812 298
rect 25846 264 25880 298
rect 25914 264 25938 298
rect 25234 229 25938 264
rect 25234 195 25268 229
rect 25302 195 25336 229
rect 25370 195 25404 229
rect 25438 195 25472 229
rect 25506 195 25540 229
rect 25574 195 25608 229
rect 25642 195 25676 229
rect 25710 195 25744 229
rect 25778 195 25812 229
rect 25846 195 25880 229
rect 25914 195 25938 229
rect 25234 160 25938 195
rect 25234 126 25268 160
rect 25302 126 25336 160
rect 25370 126 25404 160
rect 25438 126 25472 160
rect 25506 126 25540 160
rect 25574 126 25608 160
rect 25642 126 25676 160
rect 25710 126 25744 160
rect 25778 126 25812 160
rect 25846 126 25880 160
rect 25914 126 25938 160
rect 25234 91 25938 126
rect 25234 57 25268 91
rect 25302 57 25336 91
rect 25370 57 25404 91
rect 25438 57 25472 91
rect 25506 57 25540 91
rect 25574 57 25608 91
rect 25642 57 25676 91
rect 25710 57 25744 91
rect 25778 57 25812 91
rect 25846 57 25880 91
rect 25914 57 25938 91
rect 25234 22 25938 57
rect 25234 -12 25268 22
rect 25302 -12 25336 22
rect 25370 -12 25404 22
rect 25438 -12 25472 22
rect 25506 -12 25540 22
rect 25574 -12 25608 22
rect 25642 -12 25676 22
rect 25710 -12 25744 22
rect 25778 -12 25812 22
rect 25846 -12 25880 22
rect 25914 -12 25938 22
rect 25234 -36 25938 -12
<< mvnsubdiff >>
rect -335 6594 -311 6798
rect 1083 6764 1118 6798
rect 1152 6764 1187 6798
rect 1221 6764 1289 6798
rect 1323 6764 1358 6798
rect 1392 6764 1427 6798
rect 1461 6764 1496 6798
rect 1530 6764 1565 6798
rect 1599 6764 1634 6798
rect 1668 6764 1703 6798
rect 1737 6764 1772 6798
rect 1806 6764 1841 6798
rect 1875 6764 1910 6798
rect 1944 6764 1978 6798
rect 2012 6764 2046 6798
rect 1083 6730 2046 6764
rect 1083 6696 1118 6730
rect 1152 6696 1187 6730
rect 1221 6696 1323 6730
rect 1357 6696 1396 6730
rect 1430 6696 1469 6730
rect 1503 6696 1542 6730
rect 1576 6696 1614 6730
rect 1648 6696 1686 6730
rect 1720 6696 1758 6730
rect 1792 6696 1830 6730
rect 1864 6696 1902 6730
rect 1936 6696 1974 6730
rect 2008 6696 2046 6730
rect 1083 6692 2046 6696
rect 1083 6662 1255 6692
rect 1083 6628 1118 6662
rect 1152 6628 1187 6662
rect 1221 6658 1255 6662
rect 1289 6662 2046 6692
rect 1289 6661 1391 6662
rect 1289 6658 1323 6661
rect 1221 6628 1323 6658
rect -335 6525 -233 6560
rect -301 6491 -267 6525
rect -335 6456 -233 6491
rect 1255 6627 1323 6628
rect 1357 6628 1391 6661
rect 1425 6628 1464 6662
rect 1498 6628 1537 6662
rect 1571 6628 1610 6662
rect 1644 6628 1683 6662
rect 1717 6628 1756 6662
rect 1790 6628 1829 6662
rect 1863 6628 1902 6662
rect 1936 6628 1974 6662
rect 2008 6628 2046 6662
rect 2148 6764 2183 6798
rect 2217 6764 2252 6798
rect 2286 6764 2321 6798
rect 2355 6764 2390 6798
rect 2424 6764 2459 6798
rect 2493 6764 2528 6798
rect 2562 6764 2597 6798
rect 2631 6764 2666 6798
rect 2700 6764 2735 6798
rect 2769 6764 2804 6798
rect 2838 6764 2873 6798
rect 2907 6764 2942 6798
rect 2976 6764 3011 6798
rect 3045 6764 3080 6798
rect 3114 6764 3149 6798
rect 3183 6764 3218 6798
rect 3252 6764 3287 6798
rect 3321 6764 3356 6798
rect 3390 6764 3425 6798
rect 3459 6764 3494 6798
rect 3528 6764 3563 6798
rect 3597 6764 3632 6798
rect 3666 6764 3701 6798
rect 3735 6764 3770 6798
rect 3804 6764 3839 6798
rect 3873 6764 3908 6798
rect 3942 6764 3977 6798
rect 4011 6764 4046 6798
rect 4080 6764 4115 6798
rect 4149 6764 4184 6798
rect 4218 6764 4253 6798
rect 4287 6764 4322 6798
rect 4356 6764 4391 6798
rect 4425 6764 4460 6798
rect 4494 6764 4529 6798
rect 4563 6764 4598 6798
rect 4632 6764 4667 6798
rect 4701 6764 4736 6798
rect 4770 6764 4805 6798
rect 4839 6764 4874 6798
rect 4908 6764 4943 6798
rect 4977 6764 5012 6798
rect 5046 6764 5081 6798
rect 5115 6764 5150 6798
rect 5184 6764 5219 6798
rect 5253 6764 5288 6798
rect 5322 6764 5357 6798
rect 5391 6764 5426 6798
rect 5460 6764 5495 6798
rect 5529 6764 5564 6798
rect 5598 6764 5633 6798
rect 5667 6764 5702 6798
rect 5736 6764 5771 6798
rect 5805 6764 5840 6798
rect 5874 6764 5909 6798
rect 5943 6764 5978 6798
rect 6012 6764 6047 6798
rect 6081 6764 6116 6798
rect 6150 6764 6185 6798
rect 6219 6764 6254 6798
rect 6288 6764 6323 6798
rect 6357 6764 6392 6798
rect 6426 6764 6461 6798
rect 6495 6764 6530 6798
rect 6564 6764 6599 6798
rect 2148 6730 6599 6764
rect 26217 6764 26319 6798
rect 26217 6730 26285 6764
rect 2148 6696 2183 6730
rect 2217 6696 2252 6730
rect 2286 6696 2321 6730
rect 2355 6696 2390 6730
rect 2424 6696 2459 6730
rect 2493 6696 2528 6730
rect 2562 6696 2597 6730
rect 2631 6696 2666 6730
rect 2700 6696 2735 6730
rect 2769 6696 2804 6730
rect 2838 6696 2873 6730
rect 2907 6696 2942 6730
rect 2976 6696 3011 6730
rect 3045 6696 3080 6730
rect 3114 6696 3149 6730
rect 3183 6696 3218 6730
rect 3252 6696 3287 6730
rect 3321 6696 3356 6730
rect 3390 6696 3425 6730
rect 3459 6696 3494 6730
rect 3528 6696 3563 6730
rect 3597 6696 3632 6730
rect 3666 6696 3701 6730
rect 3735 6696 3770 6730
rect 3804 6696 3839 6730
rect 3873 6696 3908 6730
rect 3942 6696 3977 6730
rect 4011 6696 4046 6730
rect 4080 6696 4115 6730
rect 4149 6696 4184 6730
rect 4218 6696 4253 6730
rect 26251 6696 26319 6730
rect 2148 6662 4253 6696
rect 2148 6628 2183 6662
rect 2217 6628 2252 6662
rect 2286 6628 2321 6662
rect 2355 6628 2390 6662
rect 2424 6628 2459 6662
rect 2493 6628 2528 6662
rect 2562 6628 2597 6662
rect 2631 6628 2666 6662
rect 2700 6628 2735 6662
rect 2769 6628 2804 6662
rect 2838 6628 2873 6662
rect 2907 6628 2942 6662
rect 2976 6628 3011 6662
rect 3045 6628 3080 6662
rect 3114 6628 3149 6662
rect 3183 6628 3218 6662
rect 3252 6628 3287 6662
rect 3321 6628 3356 6662
rect 3390 6628 3425 6662
rect 3459 6628 3494 6662
rect 3528 6628 3563 6662
rect 3597 6628 3632 6662
rect 3666 6628 3701 6662
rect 3735 6628 3770 6662
rect 3804 6628 3839 6662
rect 3873 6628 3908 6662
rect 3942 6628 3977 6662
rect 4011 6628 4046 6662
rect 4080 6628 4115 6662
rect 4149 6628 4184 6662
rect 4218 6628 4253 6662
rect 26183 6695 26319 6696
rect 26183 6661 26285 6695
rect 26183 6628 26217 6661
rect 1357 6627 1425 6628
rect 1255 6622 1425 6627
rect 1289 6592 1425 6622
rect 1289 6588 1323 6592
rect 1255 6558 1323 6588
rect 1357 6558 1391 6592
rect 1255 6552 1425 6558
rect 1289 6523 1425 6552
rect 1289 6518 1323 6523
rect 1255 6489 1323 6518
rect 1357 6522 1425 6523
rect 1357 6489 1391 6522
rect 1255 6488 1391 6489
rect 1255 6482 1425 6488
rect -301 6422 -267 6456
rect -335 6387 -233 6422
rect -301 6353 -267 6387
rect -335 6318 -233 6353
rect -301 6284 -267 6318
rect -335 6249 -233 6284
rect -301 6215 -267 6249
rect -335 6180 -233 6215
rect -301 6146 -267 6180
rect -335 6111 -233 6146
rect -301 6077 -267 6111
rect -335 6042 -233 6077
rect -301 6008 -267 6042
rect -335 5973 -233 6008
rect -301 5939 -267 5973
rect -335 5904 -233 5939
rect -301 5870 -267 5904
rect -335 5835 -233 5870
rect -301 5801 -267 5835
rect -335 5766 -233 5801
rect -301 5732 -267 5766
rect -335 5697 -233 5732
rect -301 5663 -267 5697
rect -335 5628 -233 5663
rect -301 5594 -267 5628
rect -335 5558 -233 5594
rect -301 5524 -267 5558
rect -335 5488 -233 5524
rect -301 5454 -267 5488
rect -335 5418 -233 5454
rect -301 5384 -267 5418
rect -335 5348 -233 5384
rect -301 5314 -267 5348
rect -335 5278 -233 5314
rect -301 5244 -267 5278
rect -335 5208 -233 5244
rect -301 5174 -267 5208
rect -335 5138 -233 5174
rect -301 5104 -267 5138
rect -335 5068 -233 5104
rect 1289 6454 1425 6482
rect 26149 6627 26217 6628
rect 26251 6627 26319 6661
rect 26149 6626 26319 6627
rect 26149 6593 26285 6626
rect 26183 6592 26285 6593
rect 26183 6559 26217 6592
rect 26149 6558 26217 6559
rect 26251 6558 26319 6592
rect 26149 6524 26285 6558
rect 26183 6523 26319 6524
rect 26183 6490 26217 6523
rect 26149 6489 26217 6490
rect 26251 6490 26319 6523
rect 26251 6489 26285 6490
rect 1289 6448 1323 6454
rect 1255 6420 1323 6448
rect 1357 6452 1425 6454
rect 1357 6420 1391 6452
rect 1255 6418 1391 6420
rect 1255 6412 1425 6418
rect 1289 6385 1425 6412
rect 1289 6378 1323 6385
rect 1255 6351 1323 6378
rect 1357 6382 1425 6385
rect 1357 6351 1391 6382
rect 1255 6348 1391 6351
rect 1255 6342 1425 6348
rect 1289 6316 1425 6342
rect 1289 6308 1323 6316
rect 1255 6282 1323 6308
rect 1357 6312 1425 6316
rect 1357 6282 1391 6312
rect 1255 6278 1391 6282
rect 1255 6272 1425 6278
rect 1289 6247 1425 6272
rect 1289 6238 1323 6247
rect 1255 6213 1323 6238
rect 1357 6242 1425 6247
rect 1357 6213 1391 6242
rect 1255 6208 1391 6213
rect 1255 6202 1425 6208
rect 1289 6178 1425 6202
rect 1289 6168 1323 6178
rect 1255 6144 1323 6168
rect 1357 6172 1425 6178
rect 1357 6144 1391 6172
rect 1255 6138 1391 6144
rect 1255 6132 1425 6138
rect 1289 6109 1425 6132
rect 1289 6098 1323 6109
rect 1255 6075 1323 6098
rect 1357 6102 1425 6109
rect 1357 6075 1391 6102
rect 1255 6068 1391 6075
rect 1255 6062 1425 6068
rect 1289 6040 1425 6062
rect 1289 6028 1323 6040
rect 1255 6006 1323 6028
rect 1357 6032 1425 6040
rect 1357 6006 1391 6032
rect 1255 5998 1391 6006
rect 1255 5992 1425 5998
rect 1289 5971 1425 5992
rect 1289 5958 1323 5971
rect 1255 5937 1323 5958
rect 1357 5962 1425 5971
rect 1357 5937 1391 5962
rect 1255 5928 1391 5937
rect 1255 5922 1425 5928
rect 1289 5902 1425 5922
rect 1289 5888 1323 5902
rect 1255 5868 1323 5888
rect 1357 5892 1425 5902
rect 1357 5868 1391 5892
rect 1255 5858 1391 5868
rect 1255 5852 1425 5858
rect 1289 5833 1425 5852
rect 1289 5818 1323 5833
rect 1255 5799 1323 5818
rect 1357 5822 1425 5833
rect 1357 5799 1391 5822
rect 1255 5788 1391 5799
rect 1255 5782 1425 5788
rect 1289 5764 1425 5782
rect 1289 5748 1323 5764
rect 1255 5730 1323 5748
rect 1357 5751 1425 5764
rect 1357 5730 1391 5751
rect 1255 5717 1391 5730
rect 1255 5711 1425 5717
rect 1289 5695 1425 5711
rect 1289 5677 1323 5695
rect 1255 5661 1323 5677
rect 1357 5680 1425 5695
rect 1357 5661 1391 5680
rect 1255 5646 1391 5661
rect 1255 5640 1425 5646
rect 1289 5626 1425 5640
rect 1289 5606 1323 5626
rect 1255 5592 1323 5606
rect 1357 5609 1425 5626
rect 1357 5592 1391 5609
rect 1255 5575 1391 5592
rect 1255 5569 1425 5575
rect 1289 5557 1425 5569
rect 1289 5535 1323 5557
rect 1255 5523 1323 5535
rect 1357 5538 1425 5557
rect 1357 5523 1391 5538
rect 1255 5504 1391 5523
rect 1255 5498 1425 5504
rect 1289 5488 1425 5498
rect 1289 5464 1323 5488
rect 1255 5454 1323 5464
rect 1357 5467 1425 5488
rect 1357 5454 1391 5467
rect 1255 5433 1391 5454
rect 1255 5427 1425 5433
rect 1289 5419 1425 5427
rect 1289 5393 1323 5419
rect 1255 5385 1323 5393
rect 1357 5396 1425 5419
rect 1357 5385 1391 5396
rect 1255 5362 1391 5385
rect 1255 5356 1425 5362
rect 1289 5350 1425 5356
rect 1289 5322 1323 5350
rect 1255 5316 1323 5322
rect 1357 5325 1425 5350
rect 1357 5316 1391 5325
rect 1255 5291 1391 5316
rect 1255 5285 1425 5291
rect 1289 5281 1425 5285
rect 1289 5251 1323 5281
rect 1255 5247 1323 5251
rect 1357 5254 1425 5281
rect 1357 5247 1391 5254
rect 1255 5220 1391 5247
rect 1255 5214 1425 5220
rect 1289 5212 1425 5214
rect 1289 5180 1323 5212
rect 1255 5178 1323 5180
rect 1357 5183 1425 5212
rect 1357 5178 1391 5183
rect 1255 5149 1391 5178
rect 1255 5143 1425 5149
rect 1289 5142 1425 5143
rect 1289 5109 1323 5142
rect 1255 5108 1323 5109
rect 1357 5112 1425 5142
rect 1357 5108 1391 5112
rect -301 5034 -267 5068
rect -335 4998 -233 5034
rect -335 4896 -301 4964
rect 1255 5078 1391 5108
rect 1255 5072 1425 5078
rect 1289 5038 1323 5072
rect 1357 5041 1425 5072
rect 1357 5038 1391 5041
rect 1255 5007 1391 5038
rect 1255 5002 1425 5007
rect 1255 5001 1323 5002
rect 1289 4968 1323 5001
rect 1357 4970 1425 5002
rect 1357 4968 1391 4970
rect 1289 4967 1391 4968
rect 1255 4936 1391 4967
rect 1255 4932 1425 4936
rect 1255 4930 1323 4932
rect -199 4896 -165 4930
rect -131 4896 -97 4930
rect -63 4896 -29 4930
rect 5 4896 39 4930
rect 73 4896 107 4930
rect 141 4896 175 4930
rect 209 4896 243 4930
rect 277 4896 311 4930
rect 345 4896 379 4930
rect 413 4896 447 4930
rect 481 4896 515 4930
rect 549 4896 583 4930
rect 617 4896 651 4930
rect 685 4896 719 4930
rect 753 4896 787 4930
rect 821 4896 855 4930
rect 889 4896 923 4930
rect 957 4896 991 4930
rect 1025 4896 1059 4930
rect 1093 4896 1164 4930
rect 1198 4896 1255 4930
rect 1289 4898 1323 4930
rect 1357 4899 1425 4932
rect 1357 4898 1391 4899
rect 1289 4896 1391 4898
rect -335 4865 1391 4896
rect -335 4862 1425 4865
rect -335 4828 -267 4862
rect -233 4828 -197 4862
rect -163 4828 -127 4862
rect -93 4828 -57 4862
rect -23 4828 13 4862
rect 47 4828 83 4862
rect 117 4828 153 4862
rect 187 4828 223 4862
rect 257 4828 293 4862
rect 327 4828 363 4862
rect 397 4828 433 4862
rect 467 4828 503 4862
rect 537 4828 573 4862
rect 607 4828 643 4862
rect 677 4828 713 4862
rect 747 4828 783 4862
rect 817 4828 852 4862
rect 886 4828 921 4862
rect 955 4828 990 4862
rect 1024 4828 1059 4862
rect 1093 4828 1141 4862
rect 1175 4828 1232 4862
rect 1266 4828 1323 4862
rect 1357 4828 1425 4862
rect -233 4794 1391 4828
rect -165 4760 -129 4794
rect -95 4760 -59 4794
rect -25 4760 11 4794
rect 45 4760 81 4794
rect 115 4760 151 4794
rect 185 4760 221 4794
rect 255 4760 291 4794
rect 325 4760 361 4794
rect 395 4760 431 4794
rect 465 4760 501 4794
rect 535 4760 571 4794
rect 605 4760 641 4794
rect 675 4760 711 4794
rect 745 4760 781 4794
rect 815 4760 851 4794
rect 885 4760 921 4794
rect 955 4760 990 4794
rect 1024 4760 1059 4794
rect 1093 4760 1141 4794
rect 1175 4760 1212 4794
rect 1246 4760 1283 4794
rect 1317 4760 1425 4794
rect -301 4250 -165 4284
rect -335 4249 -165 4250
rect -335 4216 -267 4249
rect -301 4215 -267 4216
rect -233 4215 -199 4249
rect -301 4182 -165 4215
rect -335 4180 -165 4182
rect -335 4148 -267 4180
rect -301 4146 -267 4148
rect -233 4146 -199 4180
rect -301 4114 -165 4146
rect -335 4111 -165 4114
rect -335 4080 -267 4111
rect -301 4077 -267 4080
rect -233 4077 -199 4111
rect -301 4046 -165 4077
rect -335 4042 -165 4046
rect -335 4012 -267 4042
rect -301 4008 -267 4012
rect -233 4008 -199 4042
rect -301 3978 -165 4008
rect -335 3973 -165 3978
rect -335 3944 -267 3973
rect -301 3939 -267 3944
rect -233 3939 -199 3973
rect -301 3910 -165 3939
rect -335 3904 -165 3910
rect -335 3876 -267 3904
rect -301 3870 -267 3876
rect -233 3870 -199 3904
rect -301 3842 -165 3870
rect -335 3835 -165 3842
rect -335 3808 -267 3835
rect -301 3801 -267 3808
rect -233 3801 -199 3835
rect -301 3774 -165 3801
rect -335 3766 -165 3774
rect -335 3740 -267 3766
rect -301 3732 -267 3740
rect -233 3732 -199 3766
rect -301 3706 -165 3732
rect -335 3697 -165 3706
rect -335 3672 -267 3697
rect -301 3663 -267 3672
rect -233 3663 -199 3697
rect -301 3638 -165 3663
rect -335 3628 -165 3638
rect -335 3604 -267 3628
rect -301 3594 -267 3604
rect -233 3594 -199 3628
rect -301 3570 -165 3594
rect -335 3559 -165 3570
rect -335 3536 -267 3559
rect -301 3525 -267 3536
rect -233 3525 -199 3559
rect -301 3502 -165 3525
rect -335 3490 -165 3502
rect -335 3468 -267 3490
rect -301 3456 -267 3468
rect -233 3456 -199 3490
rect -301 3434 -165 3456
rect -335 3421 -165 3434
rect -335 3400 -267 3421
rect -301 3387 -267 3400
rect -233 3387 -199 3421
rect -301 3366 -165 3387
rect -335 3352 -165 3366
rect -335 3332 -267 3352
rect -301 3318 -267 3332
rect -233 3318 -199 3352
rect -301 3298 -165 3318
rect -335 3283 -165 3298
rect -335 3264 -267 3283
rect -301 3249 -267 3264
rect -233 3249 -199 3283
rect -301 3230 -165 3249
rect -335 3214 -165 3230
rect -335 3196 -267 3214
rect -301 3180 -267 3196
rect -233 3180 -199 3214
rect -301 3162 -165 3180
rect -335 3145 -165 3162
rect -335 3128 -267 3145
rect -301 3111 -267 3128
rect -233 3111 -199 3145
rect -301 3094 -165 3111
rect -335 3076 -165 3094
rect -335 3060 -267 3076
rect -301 3042 -267 3060
rect -233 3042 -199 3076
rect -301 3026 -165 3042
rect -335 3007 -165 3026
rect -335 2992 -267 3007
rect -301 2973 -267 2992
rect -233 2973 -199 3007
rect -301 2958 -165 2973
rect -335 2938 -165 2958
rect -335 2924 -267 2938
rect -301 2904 -267 2924
rect -233 2904 -199 2938
rect -301 2890 -165 2904
rect -335 2869 -165 2890
rect -335 2856 -267 2869
rect -301 2835 -267 2856
rect -233 2835 -199 2869
rect -301 2822 -165 2835
rect -335 2800 -165 2822
rect -335 2788 -267 2800
rect -301 2766 -267 2788
rect -233 2766 -199 2800
rect -301 2754 -165 2766
rect -335 2731 -165 2754
rect -335 2720 -267 2731
rect -301 2697 -267 2720
rect -233 2697 -199 2731
rect -301 2686 -165 2697
rect -335 2662 -165 2686
rect -335 2652 -267 2662
rect -301 2628 -267 2652
rect -233 2628 -199 2662
rect -301 2618 -165 2628
rect -335 2593 -165 2618
rect -335 2584 -267 2593
rect -301 2559 -267 2584
rect -233 2559 -199 2593
rect -301 2550 -165 2559
rect -335 2524 -165 2550
rect -335 2516 -267 2524
rect -301 2490 -267 2516
rect -233 2490 -199 2524
rect -301 2482 -165 2490
rect -335 2455 -165 2482
rect -335 2448 -267 2455
rect -301 2421 -267 2448
rect -233 2421 -199 2455
rect -301 2414 -165 2421
rect -335 2386 -165 2414
rect -335 2380 -267 2386
rect -301 2352 -267 2380
rect -233 2352 -199 2386
rect -301 2346 -165 2352
rect -335 2317 -165 2346
rect -335 2312 -267 2317
rect -301 2283 -267 2312
rect -233 2283 -199 2317
rect -301 2278 -165 2283
rect -335 2248 -165 2278
rect -335 2244 -267 2248
rect -301 2214 -267 2244
rect -233 2214 -199 2248
rect -301 2210 -165 2214
rect -335 2179 -165 2210
rect -335 2176 -267 2179
rect -301 2145 -267 2176
rect -233 2145 -199 2179
rect -301 2142 -165 2145
rect -335 2110 -165 2142
rect -335 2108 -267 2110
rect -301 2076 -267 2108
rect -233 2076 -199 2110
rect -301 2074 -165 2076
rect -335 2041 -165 2074
rect -335 2040 -267 2041
rect -301 2007 -267 2040
rect -233 2007 -199 2041
rect -301 2006 -165 2007
rect -335 1972 -165 2006
rect -301 1938 -267 1972
rect -233 1938 -199 1972
rect -335 1903 -165 1938
rect -301 1869 -267 1903
rect -233 1869 -199 1903
rect -335 1834 -165 1869
rect -301 1800 -267 1834
rect -233 1800 -199 1834
rect -335 1765 -165 1800
rect -301 1731 -267 1765
rect -233 1731 -199 1765
rect -335 1696 -165 1731
rect -301 1662 -267 1696
rect -233 1662 -199 1696
rect -335 1627 -165 1662
rect -301 1593 -267 1627
rect -233 1593 -199 1627
rect -335 1558 -165 1593
rect -301 1524 -267 1558
rect -233 1524 -199 1558
rect -335 1489 -165 1524
rect -301 1455 -267 1489
rect -233 1455 -199 1489
rect -335 1420 -165 1455
rect -301 1386 -267 1420
rect -233 1386 -199 1420
rect -335 1351 -165 1386
rect -301 1317 -267 1351
rect -233 1317 -199 1351
rect -335 1282 -165 1317
rect -301 1248 -267 1282
rect -233 1248 -199 1282
rect -335 1213 -165 1248
rect -301 1179 -267 1213
rect -233 1179 -199 1213
rect -335 1144 -165 1179
rect -301 1110 -267 1144
rect -233 1110 -199 1144
rect -335 1075 -165 1110
rect -301 1041 -267 1075
rect -233 1041 -199 1075
rect -335 1006 -165 1041
rect -301 972 -267 1006
rect -233 972 -199 1006
rect -335 937 -165 972
rect -301 903 -267 937
rect -233 903 -199 937
rect -335 868 -165 903
rect -301 834 -267 868
rect -233 834 -199 868
rect -335 799 -165 834
rect -301 765 -267 799
rect -233 765 -199 799
rect -335 730 -165 765
rect -301 696 -267 730
rect -233 696 -199 730
rect -335 661 -165 696
rect -301 627 -267 661
rect -233 627 -199 661
rect -335 592 -165 627
rect -301 558 -267 592
rect -233 558 -199 592
rect -335 523 -165 558
rect -301 489 -267 523
rect -233 489 -199 523
rect -335 454 -165 489
rect -301 420 -267 454
rect -233 420 -199 454
rect -335 385 -165 420
rect -301 351 -267 385
rect -233 351 -199 385
rect -335 316 -165 351
rect -301 282 -267 316
rect -233 282 -199 316
rect -335 247 -165 282
rect -301 213 -267 247
rect -233 213 -199 247
rect -335 178 -165 213
rect -301 144 -267 178
rect -233 144 -199 178
rect -335 120 -165 144
rect 367 4202 435 4226
rect 401 4192 435 4202
rect 469 4192 506 4226
rect 540 4192 577 4226
rect 611 4192 649 4226
rect 683 4192 721 4226
rect 755 4192 793 4226
rect 827 4192 865 4226
rect 899 4192 937 4226
rect 971 4192 1009 4226
rect 1043 4192 1081 4226
rect 1115 4192 1153 4226
rect 1187 4192 1225 4226
rect 1259 4192 1297 4226
rect 1331 4192 1369 4226
rect 1403 4192 1441 4226
rect 1475 4192 1513 4226
rect 1547 4192 1585 4226
rect 1619 4192 1657 4226
rect 1691 4202 1759 4226
rect 1691 4192 1725 4202
rect 367 4134 401 4168
rect 367 4066 401 4100
rect 1725 4125 1759 4168
rect 367 3998 401 4032
rect 367 3930 401 3964
rect 367 3862 401 3896
rect 367 3794 401 3828
rect 367 3726 401 3760
rect 367 3658 401 3692
rect 367 3590 401 3624
rect 367 3522 401 3556
rect 367 3454 401 3488
rect 367 3386 401 3420
rect 1725 4048 1759 4091
rect 1725 3972 1759 4014
rect 1725 3904 1759 3938
rect 1725 3870 1749 3904
rect 1783 3870 1817 3904
rect 1851 3870 1883 3904
rect 1987 3870 2021 3904
rect 2055 3870 2089 3904
rect 2123 3870 2157 3904
rect 2191 3870 2225 3904
rect 2259 3870 2293 3904
rect 2327 3870 2361 3904
rect 2395 3870 2429 3904
rect 2463 3870 2497 3904
rect 2531 3870 2565 3904
rect 2599 3870 2633 3904
rect 2667 3870 2701 3904
rect 2735 3870 2769 3904
rect 2803 3870 2837 3904
rect 2871 3870 2905 3904
rect 2939 3870 2973 3904
rect 3007 3870 3041 3904
rect 3075 3870 3109 3904
rect 3143 3870 3177 3904
rect 3211 3870 3245 3904
rect 3279 3870 3313 3904
rect 3347 3870 3381 3904
rect 3415 3870 3449 3904
rect 3483 3870 3517 3904
rect 3551 3870 3585 3904
rect 3619 3870 3653 3904
rect 3687 3870 3721 3904
rect 3755 3870 3789 3904
rect 3823 3870 3857 3904
rect 3891 3870 3925 3904
rect 3959 3870 3993 3904
rect 4027 3870 4062 3904
rect 4096 3870 4131 3904
rect 4165 3870 4200 3904
rect 4234 3870 4269 3904
rect 4303 3870 4338 3904
rect 4372 3870 4407 3904
rect 4441 3870 4476 3904
rect 4510 3870 4545 3904
rect 4579 3870 4614 3904
rect 4648 3870 4683 3904
rect 4717 3870 4752 3904
rect 4786 3870 4821 3904
rect 4855 3870 4890 3904
rect 4924 3870 4959 3904
rect 4993 3870 5028 3904
rect 5062 3870 5097 3904
rect 5131 3870 5166 3904
rect 5200 3870 5235 3904
rect 5269 3870 5304 3904
rect 5338 3870 5373 3904
rect 5407 3870 5442 3904
rect 5476 3870 5511 3904
rect 5545 3870 5580 3904
rect 5614 3870 5649 3904
rect 5683 3870 5718 3904
rect 5752 3870 5787 3904
rect 5821 3870 5856 3904
rect 5890 3870 5925 3904
rect 5959 3870 5994 3904
rect 6028 3870 6063 3904
rect 6097 3870 6132 3904
rect 6166 3870 6201 3904
rect 6235 3880 6303 3904
rect 6235 3870 6269 3880
rect 1725 3802 1883 3870
rect 1985 3802 2063 3870
rect 1725 3765 2063 3802
rect 1725 3731 1883 3765
rect 1917 3731 1951 3765
rect 1985 3731 2063 3765
rect 6269 3812 6303 3846
rect 6269 3744 6303 3778
rect 1725 3694 2063 3731
rect 1725 3660 1883 3694
rect 1917 3660 1951 3694
rect 1985 3660 2063 3694
rect 1725 3623 2063 3660
rect 1725 3589 1883 3623
rect 1917 3589 1951 3623
rect 1985 3589 2063 3623
rect 1725 3552 2063 3589
rect 1725 3518 1883 3552
rect 1917 3518 1951 3552
rect 1985 3518 2063 3552
rect 1725 3481 2063 3518
rect 1725 3447 1883 3481
rect 1917 3447 1951 3481
rect 1985 3447 2063 3481
rect 6269 3675 6303 3710
rect 6269 3606 6303 3641
rect 6269 3537 6303 3572
rect 1725 3410 2063 3447
rect 1725 3376 1883 3410
rect 1917 3376 1951 3410
rect 1985 3376 2063 3410
rect 367 3318 401 3352
rect 367 3250 401 3284
rect 1725 3339 2063 3376
rect 1725 3305 1883 3339
rect 1917 3305 1951 3339
rect 1985 3305 2063 3339
rect 6269 3468 6303 3503
rect 6269 3399 6303 3434
rect 6269 3330 6303 3365
rect 1725 3268 2063 3305
rect 1725 3234 1883 3268
rect 1917 3234 1951 3268
rect 1985 3234 2063 3268
rect 367 3182 401 3216
rect 1725 3227 2063 3234
rect 367 3114 401 3148
rect 1315 3197 2063 3227
rect 1315 3181 1883 3197
rect 1315 3147 1331 3181
rect 1365 3147 1399 3181
rect 1433 3147 1467 3181
rect 1501 3147 1535 3181
rect 1569 3147 1603 3181
rect 1637 3163 1883 3181
rect 1917 3163 1951 3197
rect 1985 3163 2063 3197
rect 1637 3147 2063 3163
rect 1315 3126 2063 3147
rect 1315 3110 1883 3126
rect 367 3046 401 3080
rect 1315 3076 1331 3110
rect 1365 3076 1399 3110
rect 1433 3076 1467 3110
rect 1501 3107 1883 3110
rect 1501 3076 1535 3107
rect 1315 3073 1535 3076
rect 1569 3073 1603 3107
rect 1637 3092 1883 3107
rect 1917 3092 1951 3126
rect 1985 3092 2063 3126
rect 1637 3073 2063 3092
rect 1315 3055 2063 3073
rect 367 2978 401 3012
rect 367 2910 401 2944
rect 367 2842 401 2876
rect 367 2774 401 2808
rect 1315 3039 1883 3055
rect 1315 3005 1331 3039
rect 1365 3005 1399 3039
rect 1433 3005 1467 3039
rect 1501 3033 1883 3039
rect 1501 3005 1535 3033
rect 1315 2999 1535 3005
rect 1569 2999 1603 3033
rect 1637 3021 1883 3033
rect 1917 3021 1951 3055
rect 1985 3021 2063 3055
rect 6269 3261 6303 3296
rect 6269 3192 6303 3227
rect 6269 3123 6303 3158
rect 6269 3054 6303 3089
rect 1637 2999 2063 3021
rect 1315 2984 2063 2999
rect 1315 2968 1883 2984
rect 1315 2934 1331 2968
rect 1365 2934 1399 2968
rect 1433 2934 1467 2968
rect 1501 2959 1883 2968
rect 1501 2934 1535 2959
rect 1315 2925 1535 2934
rect 1569 2925 1603 2959
rect 1637 2950 1883 2959
rect 1917 2950 1951 2984
rect 1985 2950 2063 2984
rect 1637 2925 2063 2950
rect 1315 2913 2063 2925
rect 1315 2897 1883 2913
rect 1315 2863 1331 2897
rect 1365 2863 1399 2897
rect 1433 2863 1467 2897
rect 1501 2885 1883 2897
rect 1501 2863 1535 2885
rect 1315 2851 1535 2863
rect 1569 2851 1603 2885
rect 1637 2879 1883 2885
rect 1917 2879 1951 2913
rect 1985 2879 2063 2913
rect 6269 2985 6303 3020
rect 6269 2916 6303 2951
rect 1637 2851 2063 2879
rect 1315 2842 2063 2851
rect 1315 2826 1883 2842
rect 1315 2792 1331 2826
rect 1365 2792 1399 2826
rect 1433 2792 1467 2826
rect 1501 2811 1883 2826
rect 1501 2792 1535 2811
rect 1315 2777 1535 2792
rect 1569 2777 1603 2811
rect 1637 2808 1883 2811
rect 1917 2808 1951 2842
rect 1985 2808 2063 2842
rect 1637 2777 2063 2808
rect 1315 2771 2063 2777
rect 1315 2755 1883 2771
rect 367 2706 401 2740
rect 367 2638 401 2672
rect 367 2570 401 2604
rect 367 2502 401 2536
rect 1315 2721 1331 2755
rect 1365 2721 1399 2755
rect 1433 2721 1467 2755
rect 1501 2737 1883 2755
rect 1917 2737 1951 2771
rect 1985 2737 2063 2771
rect 1501 2721 1535 2737
rect 1315 2703 1535 2721
rect 1569 2703 1603 2737
rect 1637 2703 2063 2737
rect 1315 2699 2063 2703
rect 1315 2684 1883 2699
rect 1315 2650 1331 2684
rect 1365 2650 1399 2684
rect 1433 2650 1467 2684
rect 1501 2665 1883 2684
rect 1917 2665 1951 2699
rect 1985 2665 2063 2699
rect 1501 2663 2063 2665
rect 1501 2650 1535 2663
rect 1315 2629 1535 2650
rect 1569 2629 1603 2663
rect 1637 2629 2063 2663
rect 6269 2847 6303 2882
rect 6269 2778 6303 2813
rect 6269 2709 6303 2744
rect 6269 2640 6303 2675
rect 1315 2627 2063 2629
rect 1315 2613 1883 2627
rect 1315 2579 1331 2613
rect 1365 2579 1399 2613
rect 1433 2579 1467 2613
rect 1501 2593 1883 2613
rect 1917 2593 1951 2627
rect 1985 2593 2063 2627
rect 1501 2589 2063 2593
rect 1501 2579 1535 2589
rect 1315 2555 1535 2579
rect 1569 2555 1603 2589
rect 1637 2555 2063 2589
rect 1315 2542 1883 2555
rect 1315 2508 1331 2542
rect 1365 2508 1399 2542
rect 1433 2508 1467 2542
rect 1501 2521 1883 2542
rect 1917 2521 1951 2555
rect 1985 2521 2063 2555
rect 1501 2515 2063 2521
rect 1501 2508 1535 2515
rect 367 2434 401 2468
rect 1315 2481 1535 2508
rect 1569 2481 1603 2515
rect 1637 2492 2063 2515
rect 6269 2571 6303 2606
rect 6269 2502 6303 2537
rect 1637 2483 2207 2492
rect 1637 2481 1883 2483
rect 1315 2471 1883 2481
rect 1315 2437 1331 2471
rect 1365 2437 1399 2471
rect 1433 2437 1467 2471
rect 1501 2449 1883 2471
rect 1917 2449 1951 2483
rect 1985 2458 2207 2483
rect 2241 2458 2275 2492
rect 2309 2458 2343 2492
rect 2377 2458 2411 2492
rect 2445 2458 2479 2492
rect 2513 2458 2547 2492
rect 2581 2458 2615 2492
rect 2649 2458 2683 2492
rect 2717 2458 2751 2492
rect 2785 2458 2820 2492
rect 2854 2458 2889 2492
rect 2923 2458 2958 2492
rect 2992 2458 3027 2492
rect 3061 2458 3096 2492
rect 3130 2458 3165 2492
rect 3199 2458 3234 2492
rect 3268 2458 3303 2492
rect 3337 2458 3372 2492
rect 3406 2458 3441 2492
rect 3475 2458 3510 2492
rect 3544 2458 3579 2492
rect 3613 2458 3648 2492
rect 3682 2458 3717 2492
rect 3751 2458 3786 2492
rect 3820 2458 3855 2492
rect 3889 2458 3924 2492
rect 3958 2458 3993 2492
rect 4027 2458 4062 2492
rect 4096 2458 4131 2492
rect 4165 2458 4200 2492
rect 4234 2458 4269 2492
rect 4303 2458 4338 2492
rect 4372 2458 4407 2492
rect 4441 2458 4476 2492
rect 4510 2458 4545 2492
rect 4579 2458 4614 2492
rect 4648 2458 4683 2492
rect 4717 2458 4752 2492
rect 4786 2458 4821 2492
rect 4855 2458 4890 2492
rect 4924 2458 4959 2492
rect 4993 2458 5028 2492
rect 5062 2458 5097 2492
rect 5131 2458 5166 2492
rect 5200 2458 5235 2492
rect 5269 2458 5304 2492
rect 5338 2458 5373 2492
rect 5407 2458 5442 2492
rect 5476 2458 5511 2492
rect 5545 2458 5580 2492
rect 5614 2458 5649 2492
rect 5683 2458 5718 2492
rect 5752 2458 5787 2492
rect 5821 2458 5856 2492
rect 5890 2458 5925 2492
rect 5959 2458 5994 2492
rect 6028 2458 6063 2492
rect 6097 2458 6132 2492
rect 6166 2458 6201 2492
rect 6235 2468 6269 2492
rect 6235 2458 6303 2468
rect 1985 2449 2063 2458
rect 1501 2442 2063 2449
rect 1501 2437 1535 2442
rect 367 2366 401 2400
rect 367 2298 401 2332
rect 367 2230 401 2264
rect 367 2162 401 2196
rect 367 2094 401 2128
rect 367 2026 401 2060
rect 367 1958 401 1992
rect 367 1890 401 1924
rect 1315 2408 1535 2437
rect 1569 2408 1603 2442
rect 1637 2411 2063 2442
rect 1637 2408 1883 2411
rect 1315 2400 1883 2408
rect 1315 2366 1331 2400
rect 1365 2366 1399 2400
rect 1433 2366 1467 2400
rect 1501 2377 1883 2400
rect 1917 2377 1951 2411
rect 1985 2377 2063 2411
rect 1501 2366 2063 2377
rect 1315 2328 2063 2366
rect 1315 2294 1331 2328
rect 1365 2294 1399 2328
rect 1433 2294 1467 2328
rect 1501 2294 2063 2328
rect 6269 2433 6303 2458
rect 6269 2364 6303 2399
rect 1315 2256 2063 2294
rect 1315 2222 1331 2256
rect 1365 2222 1399 2256
rect 1433 2222 1467 2256
rect 1501 2222 2063 2256
rect 1315 2184 2063 2222
rect 1315 2150 1331 2184
rect 1365 2150 1399 2184
rect 1433 2150 1467 2184
rect 1501 2150 2063 2184
rect 1315 2144 2063 2150
rect 1315 2112 1653 2144
rect 1315 2078 1331 2112
rect 1365 2078 1399 2112
rect 1433 2078 1467 2112
rect 1501 2078 1653 2112
rect 1315 2040 1653 2078
rect 1315 2006 1331 2040
rect 1365 2006 1399 2040
rect 1433 2006 1467 2040
rect 1501 2006 1653 2040
rect 1315 1968 1653 2006
rect 1315 1934 1331 1968
rect 1365 1934 1399 1968
rect 1433 1934 1467 1968
rect 1501 1934 1653 1968
rect 1315 1896 1653 1934
rect 1315 1862 1331 1896
rect 1365 1862 1399 1896
rect 1433 1862 1467 1896
rect 1501 1862 1653 1896
rect 367 1822 401 1856
rect 1315 1808 1653 1862
rect 367 1754 401 1788
rect 367 1686 401 1720
rect 367 1618 401 1652
rect 367 1550 401 1584
rect 367 1482 401 1516
rect 367 1414 401 1448
rect 367 1346 401 1380
rect 367 1278 401 1312
rect 367 1210 401 1244
rect 367 1142 401 1176
rect 367 1074 401 1108
rect 367 1006 401 1040
rect 367 938 401 972
rect 367 870 401 904
rect 367 802 401 836
rect 367 733 401 768
rect 367 664 401 699
rect 367 595 401 630
rect 367 526 401 561
rect 1607 1226 1653 1808
rect 2027 1226 2063 2144
rect 1607 1191 2063 1226
rect 1607 1157 1653 1191
rect 1687 1157 1721 1191
rect 1755 1157 1789 1191
rect 1823 1157 1857 1191
rect 1891 1157 1925 1191
rect 1959 1157 1993 1191
rect 2027 1157 2063 1191
rect 1607 1122 2063 1157
rect 1607 1088 1653 1122
rect 1687 1088 1721 1122
rect 1755 1088 1789 1122
rect 1823 1088 1857 1122
rect 1891 1088 1925 1122
rect 1959 1088 1993 1122
rect 2027 1088 2063 1122
rect 1607 1053 2063 1088
rect 1607 1019 1653 1053
rect 1687 1019 1721 1053
rect 1755 1019 1789 1053
rect 1823 1019 1857 1053
rect 1891 1019 1925 1053
rect 1959 1019 1993 1053
rect 2027 1019 2063 1053
rect 1607 984 2063 1019
rect 1607 950 1653 984
rect 1687 950 1721 984
rect 1755 950 1789 984
rect 1823 950 1857 984
rect 1891 950 1925 984
rect 1959 950 1993 984
rect 2027 950 2063 984
rect 1607 915 2063 950
rect 1607 881 1653 915
rect 1687 881 1721 915
rect 1755 881 1789 915
rect 1823 881 1857 915
rect 1891 881 1925 915
rect 1959 881 1993 915
rect 2027 881 2063 915
rect 1607 846 2063 881
rect 1607 812 1653 846
rect 1687 812 1721 846
rect 1755 812 1789 846
rect 1823 812 1857 846
rect 1891 812 1925 846
rect 1959 812 1993 846
rect 2027 812 2063 846
rect 1607 777 2063 812
rect 1607 743 1653 777
rect 1687 743 1721 777
rect 1755 743 1789 777
rect 1823 743 1857 777
rect 1891 743 1925 777
rect 1959 743 1993 777
rect 2027 743 2063 777
rect 1607 708 2063 743
rect 1607 674 1653 708
rect 1687 674 1721 708
rect 1755 674 1789 708
rect 1823 674 1857 708
rect 1891 674 1925 708
rect 1959 674 1993 708
rect 2027 674 2063 708
rect 1607 639 2063 674
rect 1607 605 1653 639
rect 1687 605 1721 639
rect 1755 605 1789 639
rect 1823 605 1857 639
rect 1891 605 1925 639
rect 1959 605 1993 639
rect 2027 605 2063 639
rect 1607 570 2063 605
rect 1607 536 1653 570
rect 1687 536 1721 570
rect 1755 536 1789 570
rect 1823 536 1857 570
rect 1891 536 1925 570
rect 1959 536 1993 570
rect 2027 536 2063 570
rect 367 457 401 492
rect 367 388 401 423
rect 1607 501 2063 536
rect 6269 2295 6303 2330
rect 6269 2226 6303 2261
rect 6269 2157 6303 2192
rect 6269 2088 6303 2123
rect 6269 2019 6303 2054
rect 6269 1950 6303 1985
rect 6269 1881 6303 1916
rect 6269 1812 6303 1847
rect 6269 1743 6303 1778
rect 6269 1674 6303 1709
rect 6269 1605 6303 1640
rect 6269 1536 6303 1571
rect 6269 1467 6303 1502
rect 6269 1398 6303 1433
rect 6269 1329 6303 1364
rect 6269 1260 6303 1295
rect 6269 1191 6303 1226
rect 6269 1122 6303 1157
rect 6269 1053 6303 1088
rect 6269 984 6303 1019
rect 6269 915 6303 950
rect 6269 846 6303 881
rect 6269 777 6303 812
rect 6269 708 6303 743
rect 6269 639 6303 674
rect 6269 570 6303 605
rect 1607 467 1653 501
rect 1687 467 1721 501
rect 1755 467 1789 501
rect 1823 467 1857 501
rect 1891 467 1925 501
rect 1959 467 1993 501
rect 2027 467 2063 501
rect 1607 432 2063 467
rect 1607 364 1653 432
rect 401 354 565 364
rect 367 330 565 354
rect 599 330 633 364
rect 667 330 701 364
rect 735 330 769 364
rect 803 330 837 364
rect 871 330 905 364
rect 939 330 973 364
rect 1007 330 1041 364
rect 1075 330 1109 364
rect 1143 330 1177 364
rect 1211 330 1245 364
rect 1279 330 1313 364
rect 1347 330 1381 364
rect 1415 330 1449 364
rect 1483 330 1517 364
rect 1551 330 1585 364
rect 1619 330 1653 364
rect 2027 364 2063 432
rect 6269 501 6303 536
rect 6269 432 6303 467
rect 6269 364 6303 398
rect 2027 330 2061 364
rect 2095 330 2129 364
rect 2163 330 2197 364
rect 2231 330 2265 364
rect 2299 330 2333 364
rect 2367 330 2401 364
rect 2435 330 2469 364
rect 2503 330 2537 364
rect 2571 330 2605 364
rect 2639 330 2673 364
rect 2707 330 2741 364
rect 2775 330 2809 364
rect 2843 330 2877 364
rect 2911 330 2945 364
rect 2979 330 3013 364
rect 3047 330 3081 364
rect 3115 330 3149 364
rect 3183 330 3217 364
rect 3251 330 3285 364
rect 3319 330 3353 364
rect 3387 330 3421 364
rect 3455 330 3489 364
rect 3523 330 3557 364
rect 3591 330 3625 364
rect 3659 330 3693 364
rect 3727 330 3761 364
rect 3795 330 3830 364
rect 3864 330 3899 364
rect 3933 330 3968 364
rect 4002 330 4037 364
rect 4071 330 4106 364
rect 4140 330 4175 364
rect 4209 330 4244 364
rect 4278 330 4313 364
rect 4347 330 4382 364
rect 4416 330 4451 364
rect 4485 330 4520 364
rect 4554 330 4589 364
rect 4623 330 4658 364
rect 4692 330 4727 364
rect 4761 330 4796 364
rect 4830 330 4865 364
rect 4899 330 4934 364
rect 4968 330 5003 364
rect 5037 330 5072 364
rect 5106 330 5141 364
rect 5175 330 5210 364
rect 5244 330 5279 364
rect 5313 330 5348 364
rect 5382 330 5417 364
rect 5451 330 5486 364
rect 5520 330 5555 364
rect 5589 330 5624 364
rect 5658 330 5693 364
rect 5727 330 5762 364
rect 5796 330 5831 364
rect 5865 330 5900 364
rect 5934 330 5969 364
rect 6003 330 6038 364
rect 6072 330 6107 364
rect 6141 330 6176 364
rect 6210 330 6245 364
rect 6279 330 6303 364
rect 26149 6456 26285 6489
rect 26149 6455 26319 6456
rect 26183 6454 26319 6455
rect 26183 6421 26217 6454
rect 26149 6420 26217 6421
rect 26251 6422 26319 6454
rect 26251 6420 26285 6422
rect 26149 6388 26285 6420
rect 26149 6386 26319 6388
rect 26183 6385 26319 6386
rect 26183 6352 26217 6385
rect 26149 6351 26217 6352
rect 26251 6354 26319 6385
rect 26251 6351 26285 6354
rect 26149 6320 26285 6351
rect 26149 6317 26319 6320
rect 26183 6316 26319 6317
rect 26183 6283 26217 6316
rect 26149 6282 26217 6283
rect 26251 6286 26319 6316
rect 26251 6282 26285 6286
rect 26149 6252 26285 6282
rect 26149 6248 26319 6252
rect 26183 6247 26319 6248
rect 26183 6214 26217 6247
rect 26149 6213 26217 6214
rect 26251 6218 26319 6247
rect 26251 6213 26285 6218
rect 26149 6184 26285 6213
rect 26149 6179 26319 6184
rect 26183 6178 26319 6179
rect 26183 6145 26217 6178
rect 26149 6144 26217 6145
rect 26251 6150 26319 6178
rect 26251 6144 26285 6150
rect 26149 6116 26285 6144
rect 26149 6110 26319 6116
rect 26183 6109 26319 6110
rect 26183 6076 26217 6109
rect 26149 6075 26217 6076
rect 26251 6082 26319 6109
rect 26251 6075 26285 6082
rect 26149 6048 26285 6075
rect 26149 6041 26319 6048
rect 26183 6040 26319 6041
rect 26183 6007 26217 6040
rect 26149 6006 26217 6007
rect 26251 6014 26319 6040
rect 26251 6006 26285 6014
rect 26149 5980 26285 6006
rect 26149 5972 26319 5980
rect 26183 5971 26319 5972
rect 26183 5938 26217 5971
rect 26149 5937 26217 5938
rect 26251 5946 26319 5971
rect 26251 5937 26285 5946
rect 26149 5912 26285 5937
rect 26149 5903 26319 5912
rect 26183 5902 26319 5903
rect 26183 5869 26217 5902
rect 26149 5868 26217 5869
rect 26251 5878 26319 5902
rect 26251 5868 26285 5878
rect 26149 5844 26285 5868
rect 26149 5834 26319 5844
rect 26183 5833 26319 5834
rect 26183 5800 26217 5833
rect 26149 5799 26217 5800
rect 26251 5810 26319 5833
rect 26251 5799 26285 5810
rect 26149 5776 26285 5799
rect 26149 5765 26319 5776
rect 26183 5764 26319 5765
rect 26183 5731 26217 5764
rect 26149 5730 26217 5731
rect 26251 5742 26319 5764
rect 26251 5730 26285 5742
rect 26149 5708 26285 5730
rect 26149 5696 26319 5708
rect 26183 5695 26319 5696
rect 26183 5662 26217 5695
rect 26149 5661 26217 5662
rect 26251 5674 26319 5695
rect 26251 5661 26285 5674
rect 26149 5640 26285 5661
rect 26149 5627 26319 5640
rect 26183 5626 26319 5627
rect 26183 5593 26217 5626
rect 26149 5592 26217 5593
rect 26251 5606 26319 5626
rect 26251 5592 26285 5606
rect 26149 5572 26285 5592
rect 26149 5558 26319 5572
rect 26183 5557 26319 5558
rect 26183 5524 26217 5557
rect 26149 5523 26217 5524
rect 26251 5538 26319 5557
rect 26251 5523 26285 5538
rect 26149 5504 26285 5523
rect 26149 5489 26319 5504
rect 26183 5488 26319 5489
rect 26183 5455 26217 5488
rect 26149 5454 26217 5455
rect 26251 5470 26319 5488
rect 26251 5454 26285 5470
rect 26149 5436 26285 5454
rect 26149 5420 26319 5436
rect 26183 5419 26319 5420
rect 26183 5386 26217 5419
rect 26149 5385 26217 5386
rect 26251 5402 26319 5419
rect 26251 5385 26285 5402
rect 26149 5368 26285 5385
rect 26149 5351 26319 5368
rect 26183 5350 26319 5351
rect 26183 5317 26217 5350
rect 26149 5316 26217 5317
rect 26251 5334 26319 5350
rect 26251 5316 26285 5334
rect 26149 5300 26285 5316
rect 26149 5282 26319 5300
rect 26183 5281 26319 5282
rect 26183 5248 26217 5281
rect 26149 5247 26217 5248
rect 26251 5266 26319 5281
rect 26251 5247 26285 5266
rect 26149 5232 26285 5247
rect 26149 5213 26319 5232
rect 26183 5212 26319 5213
rect 26183 5179 26217 5212
rect 26149 5178 26217 5179
rect 26251 5198 26319 5212
rect 26251 5178 26285 5198
rect 26149 5164 26285 5178
rect 26149 5144 26319 5164
rect 26183 5143 26319 5144
rect 26183 5110 26217 5143
rect 26149 5109 26217 5110
rect 26251 5130 26319 5143
rect 26251 5109 26285 5130
rect 26149 5096 26285 5109
rect 26149 5075 26319 5096
rect 26183 5074 26319 5075
rect 26183 5041 26217 5074
rect 26149 5040 26217 5041
rect 26251 5062 26319 5074
rect 26251 5040 26285 5062
rect 26149 5028 26285 5040
rect 26149 5006 26319 5028
rect 26183 5005 26319 5006
rect 26183 4972 26217 5005
rect 26149 4971 26217 4972
rect 26251 4994 26319 5005
rect 26251 4971 26285 4994
rect 26149 4960 26285 4971
rect 26149 4937 26319 4960
rect 26183 4936 26319 4937
rect 26183 4903 26217 4936
rect 26149 4902 26217 4903
rect 26251 4926 26319 4936
rect 26251 4902 26285 4926
rect 26149 4892 26285 4902
rect 26149 4868 26319 4892
rect 26183 4867 26319 4868
rect 26183 4834 26217 4867
rect 26149 4833 26217 4834
rect 26251 4858 26319 4867
rect 26251 4833 26285 4858
rect 26149 4824 26285 4833
rect 26149 4799 26319 4824
rect 26183 4798 26319 4799
rect 26183 4765 26217 4798
rect 26149 4764 26217 4765
rect 26251 4790 26319 4798
rect 26251 4764 26285 4790
rect 26149 4756 26285 4764
rect 26149 4730 26319 4756
rect 26183 4729 26319 4730
rect 26183 4696 26217 4729
rect 26149 4695 26217 4696
rect 26251 4722 26319 4729
rect 26251 4695 26285 4722
rect 26149 4688 26285 4695
rect 26149 4661 26319 4688
rect 26183 4660 26319 4661
rect 26183 4627 26217 4660
rect 26149 4626 26217 4627
rect 26251 4654 26319 4660
rect 26251 4626 26285 4654
rect 26149 4620 26285 4626
rect 26149 4592 26319 4620
rect 26183 4591 26319 4592
rect 26183 4558 26217 4591
rect 26149 4557 26217 4558
rect 26251 4586 26319 4591
rect 26251 4557 26285 4586
rect 26149 4552 26285 4557
rect 26149 4523 26319 4552
rect 26183 4522 26319 4523
rect 26183 4489 26217 4522
rect 26149 4488 26217 4489
rect 26251 4518 26319 4522
rect 26251 4488 26285 4518
rect 26149 4484 26285 4488
rect 26149 4454 26319 4484
rect 26183 4453 26319 4454
rect 26183 4420 26217 4453
rect 26149 4419 26217 4420
rect 26251 4450 26319 4453
rect 26251 4419 26285 4450
rect 26149 4416 26285 4419
rect 26149 4385 26319 4416
rect 26183 4384 26319 4385
rect 26183 4351 26217 4384
rect 26149 4350 26217 4351
rect 26251 4382 26319 4384
rect 26251 4350 26285 4382
rect 26149 4348 26285 4350
rect 26149 4316 26319 4348
rect 26183 4315 26319 4316
rect 26183 4282 26217 4315
rect 26149 4281 26217 4282
rect 26251 4314 26319 4315
rect 26251 4281 26285 4314
rect 26149 4280 26285 4281
rect 26149 4247 26319 4280
rect 26183 4246 26319 4247
rect 26183 4213 26217 4246
rect 26149 4178 26217 4213
rect 26149 40 26319 64
<< mvpsubdiffcont >>
rect -23 6430 11 6464
rect 49 6430 83 6464
rect 121 6430 155 6464
rect 193 6430 227 6464
rect 264 6430 298 6464
rect 335 6430 369 6464
rect 406 6430 440 6464
rect 477 6430 511 6464
rect 548 6430 582 6464
rect 619 6430 653 6464
rect 690 6430 724 6464
rect 761 6430 795 6464
rect 832 6430 866 6464
rect 903 6430 937 6464
rect 974 6430 1008 6464
rect 1045 6430 1079 6464
rect 57 6344 91 6378
rect 126 6344 160 6378
rect 195 6344 229 6378
rect 265 6344 299 6378
rect 335 6344 369 6378
rect 405 6344 439 6378
rect 475 6344 509 6378
rect 545 6344 579 6378
rect 615 6344 649 6378
rect 685 6344 719 6378
rect 755 6344 789 6378
rect 825 6344 859 6378
rect 895 6344 929 6378
rect 965 6344 999 6378
rect 1035 6344 1069 6378
rect -47 6310 -13 6344
rect 21 6276 55 6310
rect 91 6276 125 6310
rect 161 6276 195 6310
rect 231 6276 265 6310
rect 301 6276 335 6310
rect 371 6276 405 6310
rect 441 6276 475 6310
rect 511 6276 545 6310
rect 581 6276 615 6310
rect 651 6276 685 6310
rect 721 6276 755 6310
rect 791 6276 825 6310
rect 861 6276 895 6310
rect 931 6276 965 6310
rect 1001 6276 1035 6310
rect -47 6239 -13 6273
rect 21 6203 55 6237
rect 89 6208 123 6242
rect 159 6208 193 6242
rect 229 6208 263 6242
rect 299 6208 333 6242
rect 369 6208 403 6242
rect 439 6208 473 6242
rect 509 6208 543 6242
rect 579 6208 613 6242
rect 649 6208 683 6242
rect 720 6208 754 6242
rect 791 6208 825 6242
rect 862 6208 896 6242
rect 933 6208 967 6242
rect -47 6168 -13 6202
rect -47 6098 -13 6132
rect 21 6130 55 6164
rect 89 6134 123 6168
rect -47 6028 -13 6062
rect 21 6057 55 6091
rect 89 6060 123 6094
rect 1001 6206 1035 6240
rect 1069 6238 1103 6272
rect 933 6138 967 6172
rect 1001 6136 1035 6170
rect 1069 6168 1103 6202
rect -47 5958 -13 5992
rect 21 5984 55 6018
rect 89 5986 123 6020
rect -47 5888 -13 5922
rect 21 5911 55 5945
rect 89 5912 123 5946
rect -47 5818 -13 5852
rect 21 5838 55 5872
rect 89 5839 123 5873
rect -47 5748 -13 5782
rect 21 5765 55 5799
rect 89 5766 123 5800
rect -47 5678 -13 5712
rect 21 5692 55 5726
rect 89 5693 123 5727
rect -47 5608 -13 5642
rect 21 5619 55 5653
rect 89 5620 123 5654
rect -47 5538 -13 5572
rect 21 5546 55 5580
rect 89 5547 123 5581
rect -47 5468 -13 5502
rect 21 5473 55 5507
rect 89 5474 123 5508
rect -47 5398 -13 5432
rect 21 5400 55 5434
rect 89 5401 123 5435
rect 933 6068 967 6102
rect 1001 6066 1035 6100
rect 1069 6098 1103 6132
rect 933 5998 967 6032
rect 1001 5996 1035 6030
rect 1069 6028 1103 6062
rect 933 5928 967 5962
rect 1001 5926 1035 5960
rect 1069 5958 1103 5992
rect 933 5857 967 5891
rect 1001 5856 1035 5890
rect 1069 5888 1103 5922
rect 933 5786 967 5820
rect 1001 5786 1035 5820
rect 1069 5818 1103 5852
rect 933 5715 967 5749
rect 1001 5716 1035 5750
rect 1069 5748 1103 5782
rect 933 5644 967 5678
rect 1001 5646 1035 5680
rect 1069 5678 1103 5712
rect 933 5573 967 5607
rect 1001 5576 1035 5610
rect 1069 5608 1103 5642
rect 933 5502 967 5536
rect 1001 5505 1035 5539
rect 1069 5538 1103 5572
rect 1069 5468 1103 5502
rect 933 5431 967 5465
rect 1001 5434 1035 5468
rect 1069 5398 1103 5432
rect -47 5328 -13 5362
rect 21 5328 55 5362
rect 89 5328 123 5362
rect 933 5360 967 5394
rect 1001 5363 1035 5397
rect 1069 5328 1103 5362
rect 933 5289 967 5323
rect 1001 5292 1035 5326
rect 1069 5258 1103 5292
rect -23 5218 11 5252
rect 46 5218 80 5252
rect 115 5218 149 5252
rect 184 5218 218 5252
rect -23 5150 11 5184
rect 46 5150 80 5184
rect 115 5150 149 5184
rect 184 5150 218 5184
rect 253 5150 967 5252
rect 1001 5221 1035 5255
rect 1069 5187 1103 5221
rect 1001 5150 1035 5184
rect 1069 5116 1103 5150
rect -23 5082 11 5116
rect 48 5082 82 5116
rect 119 5082 153 5116
rect 190 5082 224 5116
rect 261 5082 295 5116
rect 332 5082 366 5116
rect 403 5082 437 5116
rect 473 5082 507 5116
rect 543 5082 577 5116
rect 613 5082 647 5116
rect 683 5082 717 5116
rect 753 5082 787 5116
rect 823 5082 857 5116
rect 893 5082 927 5116
rect 963 5082 997 5116
rect 1601 6426 1635 6460
rect 1670 6426 1704 6460
rect 1739 6426 1773 6460
rect 1808 6426 1842 6460
rect 1877 6426 1911 6460
rect 1946 6426 1980 6460
rect 2015 6426 2049 6460
rect 2084 6426 2118 6460
rect 2153 6426 2187 6460
rect 2222 6426 2256 6460
rect 2291 6426 2325 6460
rect 2360 6426 2394 6460
rect 2429 6426 2463 6460
rect 2498 6426 2532 6460
rect 2567 6426 2601 6460
rect 2636 6426 2670 6460
rect 2705 6426 2739 6460
rect 2774 6426 2808 6460
rect 2843 6426 2877 6460
rect 2912 6426 2946 6460
rect 2981 6426 3015 6460
rect 3050 6426 3084 6460
rect 3119 6426 3153 6460
rect 3188 6426 3222 6460
rect 3257 6426 3291 6460
rect 3326 6426 3360 6460
rect 3395 6426 3429 6460
rect 3464 6426 3498 6460
rect 3533 6426 3567 6460
rect 3602 6426 3636 6460
rect 3671 6426 3705 6460
rect 3740 6426 3774 6460
rect 3809 6426 3843 6460
rect 3878 6426 3912 6460
rect 3947 6426 3981 6460
rect 4016 6426 4050 6460
rect 4085 6426 4119 6460
rect 4154 6426 4188 6460
rect 4223 6426 4257 6460
rect 4292 6426 4326 6460
rect 4361 6426 4395 6460
rect 4430 6426 4464 6460
rect 4499 6426 4533 6460
rect 4568 6426 4602 6460
rect 4637 6426 4671 6460
rect 4706 6426 4740 6460
rect 4775 6426 4809 6460
rect 1601 6358 1635 6392
rect 1670 6358 1704 6392
rect 1739 6358 1773 6392
rect 1808 6358 1842 6392
rect 1877 6358 1911 6392
rect 1946 6358 1980 6392
rect 2015 6358 2049 6392
rect 2084 6358 2118 6392
rect 2153 6358 2187 6392
rect 2222 6358 2256 6392
rect 2291 6358 2325 6392
rect 2360 6358 2394 6392
rect 2429 6358 2463 6392
rect 2498 6358 2532 6392
rect 2567 6358 2601 6392
rect 2636 6358 2670 6392
rect 2705 6358 2739 6392
rect 2774 6358 2808 6392
rect 2843 6358 2877 6392
rect 2912 6358 2946 6392
rect 2981 6358 3015 6392
rect 3050 6358 3084 6392
rect 3119 6358 3153 6392
rect 3188 6358 3222 6392
rect 3257 6358 3291 6392
rect 3326 6358 3360 6392
rect 3395 6358 3429 6392
rect 3464 6358 3498 6392
rect 3533 6358 3567 6392
rect 3602 6358 3636 6392
rect 3671 6358 3705 6392
rect 3740 6358 3774 6392
rect 3809 6358 3843 6392
rect 3878 6358 3912 6392
rect 3947 6358 3981 6392
rect 4016 6358 4050 6392
rect 4085 6358 4119 6392
rect 4154 6358 4188 6392
rect 4223 6358 4257 6392
rect 4292 6358 4326 6392
rect 4361 6358 4395 6392
rect 4430 6358 4464 6392
rect 4499 6358 4533 6392
rect 4568 6358 4602 6392
rect 4637 6358 4671 6392
rect 4706 6358 4740 6392
rect 4775 6358 4809 6392
rect 1601 6290 1635 6324
rect 1670 6290 1704 6324
rect 1739 6290 1773 6324
rect 1808 6290 1842 6324
rect 1877 6290 1911 6324
rect 1946 6290 1980 6324
rect 2015 6290 2049 6324
rect 2084 6290 2118 6324
rect 2153 6290 2187 6324
rect 2222 6290 2256 6324
rect 2291 6290 2325 6324
rect 2360 6290 2394 6324
rect 2429 6290 2463 6324
rect 2498 6290 2532 6324
rect 2567 6290 2601 6324
rect 2636 6290 2670 6324
rect 2705 6290 2739 6324
rect 2774 6290 2808 6324
rect 2843 6290 2877 6324
rect 2912 6290 2946 6324
rect 2981 6290 3015 6324
rect 3050 6290 3084 6324
rect 3119 6290 3153 6324
rect 3188 6290 3222 6324
rect 3257 6290 3291 6324
rect 3326 6290 3360 6324
rect 3395 6290 3429 6324
rect 3464 6290 3498 6324
rect 3533 6290 3567 6324
rect 3602 6290 3636 6324
rect 3671 6290 3705 6324
rect 3740 6290 3774 6324
rect 3809 6290 3843 6324
rect 3878 6290 3912 6324
rect 3947 6290 3981 6324
rect 4016 6290 4050 6324
rect 4085 6290 4119 6324
rect 4154 6290 4188 6324
rect 4223 6290 4257 6324
rect 4292 6290 4326 6324
rect 4361 6290 4395 6324
rect 4430 6290 4464 6324
rect 4499 6290 4533 6324
rect 4568 6290 4602 6324
rect 4637 6290 4671 6324
rect 4706 6290 4740 6324
rect 4775 6290 4809 6324
rect 1601 6222 1635 6256
rect 1670 6222 1704 6256
rect 1739 6222 1773 6256
rect 1808 6222 1842 6256
rect 1877 6222 1911 6256
rect 1946 6222 1980 6256
rect 2015 6222 2049 6256
rect 2084 6222 2118 6256
rect 2153 6222 2187 6256
rect 2222 6222 2256 6256
rect 2291 6222 2325 6256
rect 2360 6222 2394 6256
rect 2429 6222 2463 6256
rect 2498 6222 2532 6256
rect 2567 6222 2601 6256
rect 2636 6222 2670 6256
rect 2705 6222 2739 6256
rect 2774 6222 2808 6256
rect 2843 6222 2877 6256
rect 2912 6222 2946 6256
rect 2981 6222 3015 6256
rect 3050 6222 3084 6256
rect 3119 6222 3153 6256
rect 3188 6222 3222 6256
rect 3257 6222 3291 6256
rect 3326 6222 3360 6256
rect 3395 6222 3429 6256
rect 3464 6222 3498 6256
rect 3533 6222 3567 6256
rect 3602 6222 3636 6256
rect 3671 6222 3705 6256
rect 3740 6222 3774 6256
rect 3809 6222 3843 6256
rect 3878 6222 3912 6256
rect 3947 6222 3981 6256
rect 4016 6222 4050 6256
rect 4085 6222 4119 6256
rect 4154 6222 4188 6256
rect 4223 6222 4257 6256
rect 4292 6222 4326 6256
rect 4361 6222 4395 6256
rect 4430 6222 4464 6256
rect 4499 6222 4533 6256
rect 4568 6222 4602 6256
rect 4637 6222 4671 6256
rect 4706 6222 4740 6256
rect 4775 6222 4809 6256
rect 1601 6154 1635 6188
rect 1670 6154 1704 6188
rect 1739 6154 1773 6188
rect 1808 6154 1842 6188
rect 1877 6154 1911 6188
rect 1946 6154 1980 6188
rect 2015 6154 2049 6188
rect 2084 6154 2118 6188
rect 2153 6154 2187 6188
rect 2222 6154 2256 6188
rect 2291 6154 2325 6188
rect 2360 6154 2394 6188
rect 2429 6154 2463 6188
rect 2498 6154 2532 6188
rect 2567 6154 2601 6188
rect 2636 6154 2670 6188
rect 2705 6154 2739 6188
rect 2774 6154 2808 6188
rect 2843 6154 2877 6188
rect 2912 6154 2946 6188
rect 2981 6154 3015 6188
rect 3050 6154 3084 6188
rect 3119 6154 3153 6188
rect 3188 6154 3222 6188
rect 3257 6154 3291 6188
rect 3326 6154 3360 6188
rect 3395 6154 3429 6188
rect 3464 6154 3498 6188
rect 3533 6154 3567 6188
rect 3602 6154 3636 6188
rect 3671 6154 3705 6188
rect 3740 6154 3774 6188
rect 3809 6154 3843 6188
rect 3878 6154 3912 6188
rect 3947 6154 3981 6188
rect 4016 6154 4050 6188
rect 4085 6154 4119 6188
rect 4154 6154 4188 6188
rect 4223 6154 4257 6188
rect 4292 6154 4326 6188
rect 4361 6154 4395 6188
rect 4430 6154 4464 6188
rect 4499 6154 4533 6188
rect 4568 6154 4602 6188
rect 4637 6154 4671 6188
rect 4706 6154 4740 6188
rect 4775 6154 4809 6188
rect 1601 6086 1635 6120
rect 1670 6086 1704 6120
rect 1739 6086 1773 6120
rect 1808 6086 1842 6120
rect 1877 6086 1911 6120
rect 1946 6086 1980 6120
rect 2015 6086 2049 6120
rect 2084 6086 2118 6120
rect 2153 6086 2187 6120
rect 2222 6086 2256 6120
rect 2291 6086 2325 6120
rect 2360 6086 2394 6120
rect 2429 6086 2463 6120
rect 2498 6086 2532 6120
rect 2567 6086 2601 6120
rect 2636 6086 2670 6120
rect 2705 6086 2739 6120
rect 2774 6086 2808 6120
rect 2843 6086 2877 6120
rect 2912 6086 2946 6120
rect 2981 6086 3015 6120
rect 3050 6086 3084 6120
rect 3119 6086 3153 6120
rect 3188 6086 3222 6120
rect 3257 6086 3291 6120
rect 3326 6086 3360 6120
rect 3395 6086 3429 6120
rect 3464 6086 3498 6120
rect 3533 6086 3567 6120
rect 3602 6086 3636 6120
rect 3671 6086 3705 6120
rect 3740 6086 3774 6120
rect 3809 6086 3843 6120
rect 3878 6086 3912 6120
rect 3947 6086 3981 6120
rect 4016 6086 4050 6120
rect 4085 6086 4119 6120
rect 4154 6086 4188 6120
rect 4223 6086 4257 6120
rect 4292 6086 4326 6120
rect 4361 6086 4395 6120
rect 4430 6086 4464 6120
rect 4499 6086 4533 6120
rect 4568 6086 4602 6120
rect 4637 6086 4671 6120
rect 4706 6086 4740 6120
rect 4775 6086 4809 6120
rect 1601 6018 1635 6052
rect 1670 6018 1704 6052
rect 1739 6018 1773 6052
rect 1808 6018 1842 6052
rect 1877 6018 1911 6052
rect 1946 6018 1980 6052
rect 2015 6018 2049 6052
rect 2084 6018 2118 6052
rect 2153 6018 2187 6052
rect 2222 6018 2256 6052
rect 2291 6018 2325 6052
rect 2360 6018 2394 6052
rect 2429 6018 2463 6052
rect 2498 6018 2532 6052
rect 2567 6018 2601 6052
rect 2636 6018 2670 6052
rect 2705 6018 2739 6052
rect 2774 6018 2808 6052
rect 2843 6018 2877 6052
rect 2912 6018 2946 6052
rect 2981 6018 3015 6052
rect 3050 6018 3084 6052
rect 3119 6018 3153 6052
rect 3188 6018 3222 6052
rect 3257 6018 3291 6052
rect 3326 6018 3360 6052
rect 3395 6018 3429 6052
rect 3464 6018 3498 6052
rect 3533 6018 3567 6052
rect 3602 6018 3636 6052
rect 3671 6018 3705 6052
rect 3740 6018 3774 6052
rect 3809 6018 3843 6052
rect 3878 6018 3912 6052
rect 3947 6018 3981 6052
rect 4016 6018 4050 6052
rect 4085 6018 4119 6052
rect 4154 6018 4188 6052
rect 4223 6018 4257 6052
rect 4292 6018 4326 6052
rect 4361 6018 4395 6052
rect 4430 6018 4464 6052
rect 4499 6018 4533 6052
rect 4568 6018 4602 6052
rect 4637 6018 4671 6052
rect 4706 6018 4740 6052
rect 4775 6018 4809 6052
rect 1601 5950 1635 5984
rect 1670 5950 1704 5984
rect 1739 5950 1773 5984
rect 1808 5950 1842 5984
rect 1877 5950 1911 5984
rect 1946 5950 1980 5984
rect 2015 5950 2049 5984
rect 2084 5950 2118 5984
rect 2153 5950 2187 5984
rect 2222 5950 2256 5984
rect 2291 5950 2325 5984
rect 2360 5950 2394 5984
rect 2429 5950 2463 5984
rect 2498 5950 2532 5984
rect 2567 5950 2601 5984
rect 2636 5950 2670 5984
rect 2705 5950 2739 5984
rect 2774 5950 2808 5984
rect 2843 5950 2877 5984
rect 2912 5950 2946 5984
rect 2981 5950 3015 5984
rect 3050 5950 3084 5984
rect 3119 5950 3153 5984
rect 3188 5950 3222 5984
rect 3257 5950 3291 5984
rect 3326 5950 3360 5984
rect 3395 5950 3429 5984
rect 3464 5950 3498 5984
rect 3533 5950 3567 5984
rect 3602 5950 3636 5984
rect 3671 5950 3705 5984
rect 3740 5950 3774 5984
rect 3809 5950 3843 5984
rect 3878 5950 3912 5984
rect 3947 5950 3981 5984
rect 4016 5950 4050 5984
rect 4085 5950 4119 5984
rect 4154 5950 4188 5984
rect 4223 5950 4257 5984
rect 4292 5950 4326 5984
rect 4361 5950 4395 5984
rect 4430 5950 4464 5984
rect 4499 5950 4533 5984
rect 4568 5950 4602 5984
rect 4637 5950 4671 5984
rect 4706 5950 4740 5984
rect 4775 5950 4809 5984
rect 1601 5882 1635 5916
rect 1670 5882 1704 5916
rect 1739 5882 1773 5916
rect 1808 5882 1842 5916
rect 1877 5882 1911 5916
rect 1946 5882 1980 5916
rect 2015 5882 2049 5916
rect 2084 5882 2118 5916
rect 2153 5882 2187 5916
rect 2222 5882 2256 5916
rect 2291 5882 2325 5916
rect 2360 5882 2394 5916
rect 2429 5882 2463 5916
rect 2498 5882 2532 5916
rect 2567 5882 2601 5916
rect 2636 5882 2670 5916
rect 2705 5882 2739 5916
rect 2774 5882 2808 5916
rect 2843 5882 2877 5916
rect 2912 5882 2946 5916
rect 2981 5882 3015 5916
rect 3050 5882 3084 5916
rect 3119 5882 3153 5916
rect 3188 5882 3222 5916
rect 3257 5882 3291 5916
rect 3326 5882 3360 5916
rect 3395 5882 3429 5916
rect 3464 5882 3498 5916
rect 3533 5882 3567 5916
rect 3602 5882 3636 5916
rect 3671 5882 3705 5916
rect 3740 5882 3774 5916
rect 3809 5882 3843 5916
rect 3878 5882 3912 5916
rect 3947 5882 3981 5916
rect 4016 5882 4050 5916
rect 4085 5882 4119 5916
rect 4154 5882 4188 5916
rect 4223 5882 4257 5916
rect 4292 5882 4326 5916
rect 4361 5882 4395 5916
rect 4430 5882 4464 5916
rect 4499 5882 4533 5916
rect 4568 5882 4602 5916
rect 4637 5882 4671 5916
rect 4706 5882 4740 5916
rect 4775 5882 4809 5916
rect 1601 5814 1635 5848
rect 1670 5814 1704 5848
rect 1739 5814 1773 5848
rect 1808 5814 1842 5848
rect 1877 5814 1911 5848
rect 1946 5814 1980 5848
rect 2015 5814 2049 5848
rect 2084 5814 2118 5848
rect 2153 5814 2187 5848
rect 2222 5814 2256 5848
rect 2291 5814 2325 5848
rect 2360 5814 2394 5848
rect 2429 5814 2463 5848
rect 2498 5814 2532 5848
rect 2567 5814 2601 5848
rect 2636 5814 2670 5848
rect 2705 5814 2739 5848
rect 2774 5814 2808 5848
rect 2843 5814 2877 5848
rect 2912 5814 2946 5848
rect 2981 5814 3015 5848
rect 3050 5814 3084 5848
rect 3119 5814 3153 5848
rect 3188 5814 3222 5848
rect 3257 5814 3291 5848
rect 3326 5814 3360 5848
rect 3395 5814 3429 5848
rect 3464 5814 3498 5848
rect 3533 5814 3567 5848
rect 3602 5814 3636 5848
rect 3671 5814 3705 5848
rect 3740 5814 3774 5848
rect 3809 5814 3843 5848
rect 3878 5814 3912 5848
rect 3947 5814 3981 5848
rect 4016 5814 4050 5848
rect 4085 5814 4119 5848
rect 4154 5814 4188 5848
rect 4223 5814 4257 5848
rect 4292 5814 4326 5848
rect 4361 5814 4395 5848
rect 4430 5814 4464 5848
rect 4499 5814 4533 5848
rect 4568 5814 4602 5848
rect 4637 5814 4671 5848
rect 4706 5814 4740 5848
rect 4775 5814 4809 5848
rect 1601 5746 1635 5780
rect 1670 5746 1704 5780
rect 1739 5746 1773 5780
rect 1808 5746 1842 5780
rect 1877 5746 1911 5780
rect 1946 5746 1980 5780
rect 2015 5746 2049 5780
rect 2084 5746 2118 5780
rect 2153 5746 2187 5780
rect 2222 5746 2256 5780
rect 2291 5746 2325 5780
rect 2360 5746 2394 5780
rect 2429 5746 2463 5780
rect 2498 5746 2532 5780
rect 2567 5746 2601 5780
rect 2636 5746 2670 5780
rect 2705 5746 2739 5780
rect 2774 5746 2808 5780
rect 2843 5746 2877 5780
rect 2912 5746 2946 5780
rect 2981 5746 3015 5780
rect 3050 5746 3084 5780
rect 3119 5746 3153 5780
rect 3188 5746 3222 5780
rect 3257 5746 3291 5780
rect 3326 5746 3360 5780
rect 3395 5746 3429 5780
rect 3464 5746 3498 5780
rect 3533 5746 3567 5780
rect 3602 5746 3636 5780
rect 3671 5746 3705 5780
rect 3740 5746 3774 5780
rect 3809 5746 3843 5780
rect 3878 5746 3912 5780
rect 3947 5746 3981 5780
rect 4016 5746 4050 5780
rect 4085 5746 4119 5780
rect 4154 5746 4188 5780
rect 4223 5746 4257 5780
rect 4292 5746 4326 5780
rect 4361 5746 4395 5780
rect 4430 5746 4464 5780
rect 4499 5746 4533 5780
rect 4568 5746 4602 5780
rect 4637 5746 4671 5780
rect 4706 5746 4740 5780
rect 4775 5746 4809 5780
rect 4844 5746 25210 6460
rect 4844 5712 6421 5746
rect 1611 5678 1645 5712
rect 1681 5678 1715 5712
rect 1751 5678 1785 5712
rect 1821 5678 1855 5712
rect 1891 5678 1925 5712
rect 1961 5678 1995 5712
rect 2030 5678 2064 5712
rect 2099 5678 2133 5712
rect 2168 5678 2202 5712
rect 2237 5678 2271 5712
rect 2306 5678 2340 5712
rect 1645 5610 1679 5644
rect 1718 5610 1752 5644
rect 1791 5610 1825 5644
rect 1864 5610 1898 5644
rect 1937 5610 1971 5644
rect 2010 5610 2044 5644
rect 2083 5610 2117 5644
rect 2156 5610 2190 5644
rect 2229 5610 2263 5644
rect 2302 5610 2336 5644
rect 1577 5570 1611 5604
rect 1645 5541 1679 5575
rect 1713 5542 1747 5576
rect 1787 5542 1821 5576
rect 1861 5542 1895 5576
rect 1935 5542 1969 5576
rect 2009 5542 2043 5576
rect 2083 5542 2117 5576
rect 2156 5542 2190 5576
rect 2229 5542 2263 5576
rect 2302 5542 2336 5576
rect 2375 5542 6421 5712
rect 1577 5499 1611 5533
rect 1645 5472 1679 5506
rect 1713 5471 1747 5505
rect 1781 5471 1815 5505
rect 1850 5471 1884 5505
rect 1919 5471 1953 5505
rect 1988 5471 2022 5505
rect 2057 5471 2091 5505
rect 2126 5471 2160 5505
rect 2195 5471 2229 5505
rect 2264 5471 2298 5505
rect 1577 5428 1611 5462
rect 1645 5403 1679 5437
rect 1713 5400 1747 5434
rect 1781 5403 1815 5437
rect 1850 5403 1884 5437
rect 1919 5403 1953 5437
rect 1988 5403 2022 5437
rect 2057 5403 2091 5437
rect 2126 5403 2160 5437
rect 2195 5403 2229 5437
rect 2264 5403 2298 5437
rect 1577 5357 1611 5391
rect 1645 5334 1679 5368
rect 1713 5329 1747 5363
rect 1781 5335 1815 5369
rect 1850 5335 1884 5369
rect 1919 5335 1953 5369
rect 1988 5335 2022 5369
rect 2057 5335 2091 5369
rect 2126 5335 2160 5369
rect 2195 5335 2229 5369
rect 2264 5335 2298 5369
rect 1577 5286 1611 5320
rect 1645 5265 1679 5299
rect 1713 5258 1747 5292
rect 1781 5267 1815 5301
rect 1850 5267 1884 5301
rect 1919 5267 1953 5301
rect 1988 5267 2022 5301
rect 2057 5267 2091 5301
rect 2126 5267 2160 5301
rect 2195 5267 2229 5301
rect 2264 5267 2298 5301
rect 1577 5215 1611 5249
rect 1645 5196 1679 5230
rect 1713 5187 1747 5221
rect 1781 5199 1815 5233
rect 1850 5199 1884 5233
rect 1919 5199 1953 5233
rect 1988 5199 2022 5233
rect 2057 5199 2091 5233
rect 2126 5199 2160 5233
rect 2195 5199 2229 5233
rect 2264 5199 2298 5233
rect 1577 5144 1611 5178
rect 1645 5127 1679 5161
rect 1713 5116 1747 5150
rect 1781 5131 1815 5165
rect 1850 5131 1884 5165
rect 1919 5131 1953 5165
rect 1988 5131 2022 5165
rect 2057 5131 2091 5165
rect 2126 5131 2160 5165
rect 2195 5131 2229 5165
rect 2264 5131 2298 5165
rect 1577 5073 1611 5107
rect 1645 5058 1679 5092
rect 1713 5045 1747 5079
rect 1781 5063 1815 5097
rect 1850 5063 1884 5097
rect 1919 5063 1953 5097
rect 1988 5063 2022 5097
rect 2057 5063 2091 5097
rect 2126 5063 2160 5097
rect 2195 5063 2229 5097
rect 2264 5063 2298 5097
rect 1577 5002 1611 5036
rect 1645 4989 1679 5023
rect 1713 4974 1747 5008
rect 1781 4995 1815 5029
rect 1850 4995 1884 5029
rect 1919 4995 1953 5029
rect 1988 4995 2022 5029
rect 2057 4995 2091 5029
rect 2126 4995 2160 5029
rect 2195 4995 2229 5029
rect 2264 4995 2298 5029
rect 2333 4995 3999 5505
rect 1577 4931 1611 4965
rect 1645 4920 1679 4954
rect 1713 4903 1747 4937
rect 1577 4860 1611 4894
rect 1645 4851 1679 4885
rect 1713 4832 1747 4866
rect 1577 4789 1611 4823
rect 1645 4782 1679 4816
rect 1713 4760 1747 4794
rect 1577 4718 1611 4752
rect 1645 4713 1679 4747
rect 1713 4688 1747 4722
rect 1577 4646 1611 4680
rect 1645 4644 1679 4678
rect 1713 4616 1747 4650
rect 79 4574 113 4608
rect 150 4574 184 4608
rect 220 4574 254 4608
rect 290 4574 324 4608
rect 360 4574 394 4608
rect 430 4574 464 4608
rect 500 4574 534 4608
rect 570 4574 604 4608
rect 640 4574 674 4608
rect 710 4574 744 4608
rect 780 4574 814 4608
rect 850 4574 884 4608
rect 920 4574 954 4608
rect 990 4574 1024 4608
rect 1060 4574 1094 4608
rect 1130 4574 1164 4608
rect 1200 4574 1234 4608
rect 1282 4574 1316 4608
rect 1356 4574 1390 4608
rect 1430 4574 1464 4608
rect 1504 4574 1538 4608
rect 1577 4574 1611 4608
rect 1645 4575 1679 4609
rect 1713 4544 1747 4578
rect 113 4506 147 4540
rect 186 4506 220 4540
rect 259 4506 293 4540
rect 332 4506 366 4540
rect 405 4506 439 4540
rect 478 4506 512 4540
rect 551 4506 585 4540
rect 624 4506 658 4540
rect 696 4506 730 4540
rect 768 4506 802 4540
rect 840 4506 874 4540
rect 912 4506 946 4540
rect 984 4506 1018 4540
rect 1056 4506 1090 4540
rect 1128 4506 1162 4540
rect 1200 4506 1234 4540
rect 1282 4506 1316 4540
rect 1355 4506 1389 4540
rect 1428 4506 1462 4540
rect 1501 4506 1535 4540
rect 1573 4506 1607 4540
rect 1645 4506 1679 4540
rect 45 4472 147 4506
rect 1713 4472 1747 4506
rect 45 3894 215 4472
rect 254 4438 288 4472
rect 327 4438 361 4472
rect 400 4438 434 4472
rect 473 4438 507 4472
rect 546 4438 580 4472
rect 619 4438 653 4472
rect 692 4438 726 4472
rect 765 4438 799 4472
rect 838 4438 872 4472
rect 911 4438 945 4472
rect 984 4438 1018 4472
rect 1056 4438 1090 4472
rect 1128 4438 1162 4472
rect 1200 4438 1234 4472
rect 1282 4438 1316 4472
rect 1360 4438 1394 4472
rect 1438 4438 1472 4472
rect 1516 4438 1550 4472
rect 1593 4438 1627 4472
rect 45 3860 79 3894
rect 45 3792 79 3826
rect 113 3825 147 3859
rect 181 3825 215 3859
rect 45 3724 79 3758
rect 113 3756 147 3790
rect 181 3756 215 3790
rect 45 3656 79 3690
rect 113 3687 147 3721
rect 181 3687 215 3721
rect 45 3588 79 3622
rect 113 3618 147 3652
rect 181 3618 215 3652
rect 45 3520 79 3554
rect 113 3549 147 3583
rect 181 3549 215 3583
rect 45 3452 79 3486
rect 113 3480 147 3514
rect 181 3480 215 3514
rect 45 3384 79 3418
rect 113 3411 147 3445
rect 181 3411 215 3445
rect 45 3316 79 3350
rect 113 3342 147 3376
rect 181 3342 215 3376
rect 45 3248 79 3282
rect 113 3273 147 3307
rect 181 3273 215 3307
rect 45 3180 79 3214
rect 113 3204 147 3238
rect 181 3204 215 3238
rect 45 3112 79 3146
rect 113 3135 147 3169
rect 181 3135 215 3169
rect 45 3044 79 3078
rect 113 3066 147 3100
rect 181 3066 215 3100
rect 45 2976 79 3010
rect 113 2997 147 3031
rect 181 2997 215 3031
rect 45 2908 79 2942
rect 113 2928 147 2962
rect 181 2928 215 2962
rect 45 2840 79 2874
rect 113 2859 147 2893
rect 181 2859 215 2893
rect 45 2772 79 2806
rect 113 2790 147 2824
rect 181 2790 215 2824
rect 45 2704 79 2738
rect 113 2721 147 2755
rect 181 2721 215 2755
rect 45 2636 79 2670
rect 113 2652 147 2686
rect 181 2652 215 2686
rect 45 2568 79 2602
rect 113 2583 147 2617
rect 181 2583 215 2617
rect 45 2500 79 2534
rect 113 2514 147 2548
rect 181 2514 215 2548
rect 45 2432 79 2466
rect 113 2445 147 2479
rect 181 2445 215 2479
rect 45 2364 79 2398
rect 113 2376 147 2410
rect 181 2376 215 2410
rect 45 2296 79 2330
rect 113 2307 147 2341
rect 181 2307 215 2341
rect 45 2228 79 2262
rect 113 2238 147 2272
rect 181 2238 215 2272
rect 45 2160 79 2194
rect 113 2169 147 2203
rect 181 2169 215 2203
rect 45 2092 79 2126
rect 113 2100 147 2134
rect 181 2100 215 2134
rect 45 2024 79 2058
rect 113 2031 147 2065
rect 181 2031 215 2065
rect 45 1956 79 1990
rect 113 1962 147 1996
rect 181 1962 215 1996
rect 45 1888 79 1922
rect 113 1893 147 1927
rect 181 1893 215 1927
rect 45 1820 79 1854
rect 113 1824 147 1858
rect 181 1824 215 1858
rect 45 1752 79 1786
rect 113 1755 147 1789
rect 181 1755 215 1789
rect 45 1684 79 1718
rect 113 1686 147 1720
rect 181 1686 215 1720
rect 45 1616 79 1650
rect 113 1617 147 1651
rect 181 1617 215 1651
rect 45 1548 79 1582
rect 113 1548 147 1582
rect 181 1548 215 1582
rect 45 1479 79 1513
rect 113 1479 147 1513
rect 181 1479 215 1513
rect 45 1410 79 1444
rect 113 1410 147 1444
rect 181 1410 215 1444
rect 45 1341 79 1375
rect 113 1341 147 1375
rect 181 1341 215 1375
rect 45 1272 79 1306
rect 113 1272 147 1306
rect 181 1272 215 1306
rect 45 1203 79 1237
rect 113 1203 147 1237
rect 181 1203 215 1237
rect 45 1134 79 1168
rect 113 1134 147 1168
rect 181 1134 215 1168
rect 45 1065 79 1099
rect 113 1065 147 1099
rect 181 1065 215 1099
rect 45 996 79 1030
rect 113 996 147 1030
rect 181 996 215 1030
rect 45 927 79 961
rect 113 927 147 961
rect 181 927 215 961
rect 45 858 79 892
rect 113 858 147 892
rect 181 858 215 892
rect 45 789 79 823
rect 113 789 147 823
rect 181 789 215 823
rect 45 720 79 754
rect 113 720 147 754
rect 181 720 215 754
rect 45 651 79 685
rect 113 651 147 685
rect 181 651 215 685
rect 45 582 79 616
rect 113 582 147 616
rect 181 582 215 616
rect 45 513 79 547
rect 113 513 147 547
rect 181 513 215 547
rect 45 444 79 478
rect 113 444 147 478
rect 181 444 215 478
rect 45 375 79 409
rect 113 375 147 409
rect 181 375 215 409
rect 45 306 79 340
rect 113 306 147 340
rect 181 306 215 340
rect 45 237 79 271
rect 113 237 147 271
rect 181 237 215 271
rect 45 168 79 202
rect 113 168 147 202
rect 181 168 215 202
rect 25268 2058 25914 6444
rect 25268 1989 25302 2023
rect 25336 1989 25370 2023
rect 25404 1989 25438 2023
rect 25472 1989 25506 2023
rect 25540 1989 25574 2023
rect 25608 1989 25642 2023
rect 25676 1989 25710 2023
rect 25744 1989 25778 2023
rect 25812 1989 25846 2023
rect 25880 1989 25914 2023
rect 25268 1920 25302 1954
rect 25336 1920 25370 1954
rect 25404 1920 25438 1954
rect 25472 1920 25506 1954
rect 25540 1920 25574 1954
rect 25608 1920 25642 1954
rect 25676 1920 25710 1954
rect 25744 1920 25778 1954
rect 25812 1920 25846 1954
rect 25880 1920 25914 1954
rect 25268 1851 25302 1885
rect 25336 1851 25370 1885
rect 25404 1851 25438 1885
rect 25472 1851 25506 1885
rect 25540 1851 25574 1885
rect 25608 1851 25642 1885
rect 25676 1851 25710 1885
rect 25744 1851 25778 1885
rect 25812 1851 25846 1885
rect 25880 1851 25914 1885
rect 25268 1782 25302 1816
rect 25336 1782 25370 1816
rect 25404 1782 25438 1816
rect 25472 1782 25506 1816
rect 25540 1782 25574 1816
rect 25608 1782 25642 1816
rect 25676 1782 25710 1816
rect 25744 1782 25778 1816
rect 25812 1782 25846 1816
rect 25880 1782 25914 1816
rect 25268 1713 25302 1747
rect 25336 1713 25370 1747
rect 25404 1713 25438 1747
rect 25472 1713 25506 1747
rect 25540 1713 25574 1747
rect 25608 1713 25642 1747
rect 25676 1713 25710 1747
rect 25744 1713 25778 1747
rect 25812 1713 25846 1747
rect 25880 1713 25914 1747
rect 25268 1644 25302 1678
rect 25336 1644 25370 1678
rect 25404 1644 25438 1678
rect 25472 1644 25506 1678
rect 25540 1644 25574 1678
rect 25608 1644 25642 1678
rect 25676 1644 25710 1678
rect 25744 1644 25778 1678
rect 25812 1644 25846 1678
rect 25880 1644 25914 1678
rect 25268 1575 25302 1609
rect 25336 1575 25370 1609
rect 25404 1575 25438 1609
rect 25472 1575 25506 1609
rect 25540 1575 25574 1609
rect 25608 1575 25642 1609
rect 25676 1575 25710 1609
rect 25744 1575 25778 1609
rect 25812 1575 25846 1609
rect 25880 1575 25914 1609
rect 25268 1506 25302 1540
rect 25336 1506 25370 1540
rect 25404 1506 25438 1540
rect 25472 1506 25506 1540
rect 25540 1506 25574 1540
rect 25608 1506 25642 1540
rect 25676 1506 25710 1540
rect 25744 1506 25778 1540
rect 25812 1506 25846 1540
rect 25880 1506 25914 1540
rect 25268 1437 25302 1471
rect 25336 1437 25370 1471
rect 25404 1437 25438 1471
rect 25472 1437 25506 1471
rect 25540 1437 25574 1471
rect 25608 1437 25642 1471
rect 25676 1437 25710 1471
rect 25744 1437 25778 1471
rect 25812 1437 25846 1471
rect 25880 1437 25914 1471
rect 25268 1368 25302 1402
rect 25336 1368 25370 1402
rect 25404 1368 25438 1402
rect 25472 1368 25506 1402
rect 25540 1368 25574 1402
rect 25608 1368 25642 1402
rect 25676 1368 25710 1402
rect 25744 1368 25778 1402
rect 25812 1368 25846 1402
rect 25880 1368 25914 1402
rect 25268 1299 25302 1333
rect 25336 1299 25370 1333
rect 25404 1299 25438 1333
rect 25472 1299 25506 1333
rect 25540 1299 25574 1333
rect 25608 1299 25642 1333
rect 25676 1299 25710 1333
rect 25744 1299 25778 1333
rect 25812 1299 25846 1333
rect 25880 1299 25914 1333
rect 25268 1230 25302 1264
rect 25336 1230 25370 1264
rect 25404 1230 25438 1264
rect 25472 1230 25506 1264
rect 25540 1230 25574 1264
rect 25608 1230 25642 1264
rect 25676 1230 25710 1264
rect 25744 1230 25778 1264
rect 25812 1230 25846 1264
rect 25880 1230 25914 1264
rect 25268 1161 25302 1195
rect 25336 1161 25370 1195
rect 25404 1161 25438 1195
rect 25472 1161 25506 1195
rect 25540 1161 25574 1195
rect 25608 1161 25642 1195
rect 25676 1161 25710 1195
rect 25744 1161 25778 1195
rect 25812 1161 25846 1195
rect 25880 1161 25914 1195
rect 25268 1092 25302 1126
rect 25336 1092 25370 1126
rect 25404 1092 25438 1126
rect 25472 1092 25506 1126
rect 25540 1092 25574 1126
rect 25608 1092 25642 1126
rect 25676 1092 25710 1126
rect 25744 1092 25778 1126
rect 25812 1092 25846 1126
rect 25880 1092 25914 1126
rect 25268 1023 25302 1057
rect 25336 1023 25370 1057
rect 25404 1023 25438 1057
rect 25472 1023 25506 1057
rect 25540 1023 25574 1057
rect 25608 1023 25642 1057
rect 25676 1023 25710 1057
rect 25744 1023 25778 1057
rect 25812 1023 25846 1057
rect 25880 1023 25914 1057
rect 25268 954 25302 988
rect 25336 954 25370 988
rect 25404 954 25438 988
rect 25472 954 25506 988
rect 25540 954 25574 988
rect 25608 954 25642 988
rect 25676 954 25710 988
rect 25744 954 25778 988
rect 25812 954 25846 988
rect 25880 954 25914 988
rect 25268 885 25302 919
rect 25336 885 25370 919
rect 25404 885 25438 919
rect 25472 885 25506 919
rect 25540 885 25574 919
rect 25608 885 25642 919
rect 25676 885 25710 919
rect 25744 885 25778 919
rect 25812 885 25846 919
rect 25880 885 25914 919
rect 25268 816 25302 850
rect 25336 816 25370 850
rect 25404 816 25438 850
rect 25472 816 25506 850
rect 25540 816 25574 850
rect 25608 816 25642 850
rect 25676 816 25710 850
rect 25744 816 25778 850
rect 25812 816 25846 850
rect 25880 816 25914 850
rect 25268 747 25302 781
rect 25336 747 25370 781
rect 25404 747 25438 781
rect 25472 747 25506 781
rect 25540 747 25574 781
rect 25608 747 25642 781
rect 25676 747 25710 781
rect 25744 747 25778 781
rect 25812 747 25846 781
rect 25880 747 25914 781
rect 25268 678 25302 712
rect 25336 678 25370 712
rect 25404 678 25438 712
rect 25472 678 25506 712
rect 25540 678 25574 712
rect 25608 678 25642 712
rect 25676 678 25710 712
rect 25744 678 25778 712
rect 25812 678 25846 712
rect 25880 678 25914 712
rect 25268 609 25302 643
rect 25336 609 25370 643
rect 25404 609 25438 643
rect 25472 609 25506 643
rect 25540 609 25574 643
rect 25608 609 25642 643
rect 25676 609 25710 643
rect 25744 609 25778 643
rect 25812 609 25846 643
rect 25880 609 25914 643
rect 25268 540 25302 574
rect 25336 540 25370 574
rect 25404 540 25438 574
rect 25472 540 25506 574
rect 25540 540 25574 574
rect 25608 540 25642 574
rect 25676 540 25710 574
rect 25744 540 25778 574
rect 25812 540 25846 574
rect 25880 540 25914 574
rect 25268 471 25302 505
rect 25336 471 25370 505
rect 25404 471 25438 505
rect 25472 471 25506 505
rect 25540 471 25574 505
rect 25608 471 25642 505
rect 25676 471 25710 505
rect 25744 471 25778 505
rect 25812 471 25846 505
rect 25880 471 25914 505
rect 25268 402 25302 436
rect 25336 402 25370 436
rect 25404 402 25438 436
rect 25472 402 25506 436
rect 25540 402 25574 436
rect 25608 402 25642 436
rect 25676 402 25710 436
rect 25744 402 25778 436
rect 25812 402 25846 436
rect 25880 402 25914 436
rect 25268 333 25302 367
rect 25336 333 25370 367
rect 25404 333 25438 367
rect 25472 333 25506 367
rect 25540 333 25574 367
rect 25608 333 25642 367
rect 25676 333 25710 367
rect 25744 333 25778 367
rect 25812 333 25846 367
rect 25880 333 25914 367
rect 25268 264 25302 298
rect 25336 264 25370 298
rect 25404 264 25438 298
rect 25472 264 25506 298
rect 25540 264 25574 298
rect 25608 264 25642 298
rect 25676 264 25710 298
rect 25744 264 25778 298
rect 25812 264 25846 298
rect 25880 264 25914 298
rect 25268 195 25302 229
rect 25336 195 25370 229
rect 25404 195 25438 229
rect 25472 195 25506 229
rect 25540 195 25574 229
rect 25608 195 25642 229
rect 25676 195 25710 229
rect 25744 195 25778 229
rect 25812 195 25846 229
rect 25880 195 25914 229
rect 25268 126 25302 160
rect 25336 126 25370 160
rect 25404 126 25438 160
rect 25472 126 25506 160
rect 25540 126 25574 160
rect 25608 126 25642 160
rect 25676 126 25710 160
rect 25744 126 25778 160
rect 25812 126 25846 160
rect 25880 126 25914 160
rect 25268 57 25302 91
rect 25336 57 25370 91
rect 25404 57 25438 91
rect 25472 57 25506 91
rect 25540 57 25574 91
rect 25608 57 25642 91
rect 25676 57 25710 91
rect 25744 57 25778 91
rect 25812 57 25846 91
rect 25880 57 25914 91
rect 25268 -12 25302 22
rect 25336 -12 25370 22
rect 25404 -12 25438 22
rect 25472 -12 25506 22
rect 25540 -12 25574 22
rect 25608 -12 25642 22
rect 25676 -12 25710 22
rect 25744 -12 25778 22
rect 25812 -12 25846 22
rect 25880 -12 25914 22
<< mvnsubdiffcont >>
rect -311 6628 1083 6798
rect 1118 6764 1152 6798
rect 1187 6764 1221 6798
rect 1289 6764 1323 6798
rect 1358 6764 1392 6798
rect 1427 6764 1461 6798
rect 1496 6764 1530 6798
rect 1565 6764 1599 6798
rect 1634 6764 1668 6798
rect 1703 6764 1737 6798
rect 1772 6764 1806 6798
rect 1841 6764 1875 6798
rect 1910 6764 1944 6798
rect 1978 6764 2012 6798
rect 1118 6696 1152 6730
rect 1187 6696 1221 6730
rect 1323 6696 1357 6730
rect 1396 6696 1430 6730
rect 1469 6696 1503 6730
rect 1542 6696 1576 6730
rect 1614 6696 1648 6730
rect 1686 6696 1720 6730
rect 1758 6696 1792 6730
rect 1830 6696 1864 6730
rect 1902 6696 1936 6730
rect 1974 6696 2008 6730
rect 1118 6628 1152 6662
rect 1187 6628 1221 6662
rect 1255 6658 1289 6692
rect -311 6594 -233 6628
rect -335 6560 -233 6594
rect -335 6491 -301 6525
rect -267 6491 -233 6525
rect 1323 6627 1357 6661
rect 1391 6628 1425 6662
rect 1464 6628 1498 6662
rect 1537 6628 1571 6662
rect 1610 6628 1644 6662
rect 1683 6628 1717 6662
rect 1756 6628 1790 6662
rect 1829 6628 1863 6662
rect 1902 6628 1936 6662
rect 1974 6628 2008 6662
rect 2046 6628 2148 6798
rect 2183 6764 2217 6798
rect 2252 6764 2286 6798
rect 2321 6764 2355 6798
rect 2390 6764 2424 6798
rect 2459 6764 2493 6798
rect 2528 6764 2562 6798
rect 2597 6764 2631 6798
rect 2666 6764 2700 6798
rect 2735 6764 2769 6798
rect 2804 6764 2838 6798
rect 2873 6764 2907 6798
rect 2942 6764 2976 6798
rect 3011 6764 3045 6798
rect 3080 6764 3114 6798
rect 3149 6764 3183 6798
rect 3218 6764 3252 6798
rect 3287 6764 3321 6798
rect 3356 6764 3390 6798
rect 3425 6764 3459 6798
rect 3494 6764 3528 6798
rect 3563 6764 3597 6798
rect 3632 6764 3666 6798
rect 3701 6764 3735 6798
rect 3770 6764 3804 6798
rect 3839 6764 3873 6798
rect 3908 6764 3942 6798
rect 3977 6764 4011 6798
rect 4046 6764 4080 6798
rect 4115 6764 4149 6798
rect 4184 6764 4218 6798
rect 4253 6764 4287 6798
rect 4322 6764 4356 6798
rect 4391 6764 4425 6798
rect 4460 6764 4494 6798
rect 4529 6764 4563 6798
rect 4598 6764 4632 6798
rect 4667 6764 4701 6798
rect 4736 6764 4770 6798
rect 4805 6764 4839 6798
rect 4874 6764 4908 6798
rect 4943 6764 4977 6798
rect 5012 6764 5046 6798
rect 5081 6764 5115 6798
rect 5150 6764 5184 6798
rect 5219 6764 5253 6798
rect 5288 6764 5322 6798
rect 5357 6764 5391 6798
rect 5426 6764 5460 6798
rect 5495 6764 5529 6798
rect 5564 6764 5598 6798
rect 5633 6764 5667 6798
rect 5702 6764 5736 6798
rect 5771 6764 5805 6798
rect 5840 6764 5874 6798
rect 5909 6764 5943 6798
rect 5978 6764 6012 6798
rect 6047 6764 6081 6798
rect 6116 6764 6150 6798
rect 6185 6764 6219 6798
rect 6254 6764 6288 6798
rect 6323 6764 6357 6798
rect 6392 6764 6426 6798
rect 6461 6764 6495 6798
rect 6530 6764 6564 6798
rect 6599 6730 26217 6798
rect 26285 6730 26319 6764
rect 2183 6696 2217 6730
rect 2252 6696 2286 6730
rect 2321 6696 2355 6730
rect 2390 6696 2424 6730
rect 2459 6696 2493 6730
rect 2528 6696 2562 6730
rect 2597 6696 2631 6730
rect 2666 6696 2700 6730
rect 2735 6696 2769 6730
rect 2804 6696 2838 6730
rect 2873 6696 2907 6730
rect 2942 6696 2976 6730
rect 3011 6696 3045 6730
rect 3080 6696 3114 6730
rect 3149 6696 3183 6730
rect 3218 6696 3252 6730
rect 3287 6696 3321 6730
rect 3356 6696 3390 6730
rect 3425 6696 3459 6730
rect 3494 6696 3528 6730
rect 3563 6696 3597 6730
rect 3632 6696 3666 6730
rect 3701 6696 3735 6730
rect 3770 6696 3804 6730
rect 3839 6696 3873 6730
rect 3908 6696 3942 6730
rect 3977 6696 4011 6730
rect 4046 6696 4080 6730
rect 4115 6696 4149 6730
rect 4184 6696 4218 6730
rect 4253 6696 26251 6730
rect 2183 6628 2217 6662
rect 2252 6628 2286 6662
rect 2321 6628 2355 6662
rect 2390 6628 2424 6662
rect 2459 6628 2493 6662
rect 2528 6628 2562 6662
rect 2597 6628 2631 6662
rect 2666 6628 2700 6662
rect 2735 6628 2769 6662
rect 2804 6628 2838 6662
rect 2873 6628 2907 6662
rect 2942 6628 2976 6662
rect 3011 6628 3045 6662
rect 3080 6628 3114 6662
rect 3149 6628 3183 6662
rect 3218 6628 3252 6662
rect 3287 6628 3321 6662
rect 3356 6628 3390 6662
rect 3425 6628 3459 6662
rect 3494 6628 3528 6662
rect 3563 6628 3597 6662
rect 3632 6628 3666 6662
rect 3701 6628 3735 6662
rect 3770 6628 3804 6662
rect 3839 6628 3873 6662
rect 3908 6628 3942 6662
rect 3977 6628 4011 6662
rect 4046 6628 4080 6662
rect 4115 6628 4149 6662
rect 4184 6628 4218 6662
rect 4253 6628 26183 6696
rect 26285 6661 26319 6695
rect 1255 6588 1289 6622
rect 1323 6558 1357 6592
rect 1391 6558 1425 6592
rect 1255 6518 1289 6552
rect 1323 6489 1357 6523
rect 1391 6488 1425 6522
rect -335 6422 -301 6456
rect -267 6422 -233 6456
rect -335 6353 -301 6387
rect -267 6353 -233 6387
rect -335 6284 -301 6318
rect -267 6284 -233 6318
rect -335 6215 -301 6249
rect -267 6215 -233 6249
rect -335 6146 -301 6180
rect -267 6146 -233 6180
rect -335 6077 -301 6111
rect -267 6077 -233 6111
rect -335 6008 -301 6042
rect -267 6008 -233 6042
rect -335 5939 -301 5973
rect -267 5939 -233 5973
rect -335 5870 -301 5904
rect -267 5870 -233 5904
rect -335 5801 -301 5835
rect -267 5801 -233 5835
rect -335 5732 -301 5766
rect -267 5732 -233 5766
rect -335 5663 -301 5697
rect -267 5663 -233 5697
rect -335 5594 -301 5628
rect -267 5594 -233 5628
rect -335 5524 -301 5558
rect -267 5524 -233 5558
rect -335 5454 -301 5488
rect -267 5454 -233 5488
rect -335 5384 -301 5418
rect -267 5384 -233 5418
rect -335 5314 -301 5348
rect -267 5314 -233 5348
rect -335 5244 -301 5278
rect -267 5244 -233 5278
rect -335 5174 -301 5208
rect -267 5174 -233 5208
rect -335 5104 -301 5138
rect -267 5104 -233 5138
rect 1255 6448 1289 6482
rect 26217 6627 26251 6661
rect 26149 6559 26183 6593
rect 26285 6592 26319 6626
rect 26217 6558 26251 6592
rect 26285 6524 26319 6558
rect 26149 6490 26183 6524
rect 26217 6489 26251 6523
rect 1323 6420 1357 6454
rect 1391 6418 1425 6452
rect 1255 6378 1289 6412
rect 1323 6351 1357 6385
rect 1391 6348 1425 6382
rect 1255 6308 1289 6342
rect 1323 6282 1357 6316
rect 1391 6278 1425 6312
rect 1255 6238 1289 6272
rect 1323 6213 1357 6247
rect 1391 6208 1425 6242
rect 1255 6168 1289 6202
rect 1323 6144 1357 6178
rect 1391 6138 1425 6172
rect 1255 6098 1289 6132
rect 1323 6075 1357 6109
rect 1391 6068 1425 6102
rect 1255 6028 1289 6062
rect 1323 6006 1357 6040
rect 1391 5998 1425 6032
rect 1255 5958 1289 5992
rect 1323 5937 1357 5971
rect 1391 5928 1425 5962
rect 1255 5888 1289 5922
rect 1323 5868 1357 5902
rect 1391 5858 1425 5892
rect 1255 5818 1289 5852
rect 1323 5799 1357 5833
rect 1391 5788 1425 5822
rect 1255 5748 1289 5782
rect 1323 5730 1357 5764
rect 1391 5717 1425 5751
rect 1255 5677 1289 5711
rect 1323 5661 1357 5695
rect 1391 5646 1425 5680
rect 1255 5606 1289 5640
rect 1323 5592 1357 5626
rect 1391 5575 1425 5609
rect 1255 5535 1289 5569
rect 1323 5523 1357 5557
rect 1391 5504 1425 5538
rect 1255 5464 1289 5498
rect 1323 5454 1357 5488
rect 1391 5433 1425 5467
rect 1255 5393 1289 5427
rect 1323 5385 1357 5419
rect 1391 5362 1425 5396
rect 1255 5322 1289 5356
rect 1323 5316 1357 5350
rect 1391 5291 1425 5325
rect 1255 5251 1289 5285
rect 1323 5247 1357 5281
rect 1391 5220 1425 5254
rect 1255 5180 1289 5214
rect 1323 5178 1357 5212
rect 1391 5149 1425 5183
rect 1255 5109 1289 5143
rect 1323 5108 1357 5142
rect -335 5034 -301 5068
rect -267 5034 -233 5068
rect -335 4964 -233 4998
rect -301 4930 -233 4964
rect 1391 5078 1425 5112
rect 1255 5038 1289 5072
rect 1323 5038 1357 5072
rect 1391 5007 1425 5041
rect 1255 4967 1289 5001
rect 1323 4968 1357 5002
rect 1391 4936 1425 4970
rect -301 4896 -199 4930
rect -165 4896 -131 4930
rect -97 4896 -63 4930
rect -29 4896 5 4930
rect 39 4896 73 4930
rect 107 4896 141 4930
rect 175 4896 209 4930
rect 243 4896 277 4930
rect 311 4896 345 4930
rect 379 4896 413 4930
rect 447 4896 481 4930
rect 515 4896 549 4930
rect 583 4896 617 4930
rect 651 4896 685 4930
rect 719 4896 753 4930
rect 787 4896 821 4930
rect 855 4896 889 4930
rect 923 4896 957 4930
rect 991 4896 1025 4930
rect 1059 4896 1093 4930
rect 1164 4896 1198 4930
rect 1255 4896 1289 4930
rect 1323 4898 1357 4932
rect 1391 4865 1425 4899
rect -267 4828 -233 4862
rect -197 4828 -163 4862
rect -127 4828 -93 4862
rect -57 4828 -23 4862
rect 13 4828 47 4862
rect 83 4828 117 4862
rect 153 4828 187 4862
rect 223 4828 257 4862
rect 293 4828 327 4862
rect 363 4828 397 4862
rect 433 4828 467 4862
rect 503 4828 537 4862
rect 573 4828 607 4862
rect 643 4828 677 4862
rect 713 4828 747 4862
rect 783 4828 817 4862
rect 852 4828 886 4862
rect 921 4828 955 4862
rect 990 4828 1024 4862
rect 1059 4828 1093 4862
rect 1141 4828 1175 4862
rect 1232 4828 1266 4862
rect 1323 4828 1357 4862
rect -335 4794 -233 4828
rect 1391 4794 1425 4828
rect -335 4284 -165 4794
rect -129 4760 -95 4794
rect -59 4760 -25 4794
rect 11 4760 45 4794
rect 81 4760 115 4794
rect 151 4760 185 4794
rect 221 4760 255 4794
rect 291 4760 325 4794
rect 361 4760 395 4794
rect 431 4760 465 4794
rect 501 4760 535 4794
rect 571 4760 605 4794
rect 641 4760 675 4794
rect 711 4760 745 4794
rect 781 4760 815 4794
rect 851 4760 885 4794
rect 921 4760 955 4794
rect 990 4760 1024 4794
rect 1059 4760 1093 4794
rect 1141 4760 1175 4794
rect 1212 4760 1246 4794
rect 1283 4760 1317 4794
rect -335 4250 -301 4284
rect -335 4182 -301 4216
rect -267 4215 -233 4249
rect -199 4215 -165 4249
rect -335 4114 -301 4148
rect -267 4146 -233 4180
rect -199 4146 -165 4180
rect -335 4046 -301 4080
rect -267 4077 -233 4111
rect -199 4077 -165 4111
rect -335 3978 -301 4012
rect -267 4008 -233 4042
rect -199 4008 -165 4042
rect -335 3910 -301 3944
rect -267 3939 -233 3973
rect -199 3939 -165 3973
rect -335 3842 -301 3876
rect -267 3870 -233 3904
rect -199 3870 -165 3904
rect -335 3774 -301 3808
rect -267 3801 -233 3835
rect -199 3801 -165 3835
rect -335 3706 -301 3740
rect -267 3732 -233 3766
rect -199 3732 -165 3766
rect -335 3638 -301 3672
rect -267 3663 -233 3697
rect -199 3663 -165 3697
rect -335 3570 -301 3604
rect -267 3594 -233 3628
rect -199 3594 -165 3628
rect -335 3502 -301 3536
rect -267 3525 -233 3559
rect -199 3525 -165 3559
rect -335 3434 -301 3468
rect -267 3456 -233 3490
rect -199 3456 -165 3490
rect -335 3366 -301 3400
rect -267 3387 -233 3421
rect -199 3387 -165 3421
rect -335 3298 -301 3332
rect -267 3318 -233 3352
rect -199 3318 -165 3352
rect -335 3230 -301 3264
rect -267 3249 -233 3283
rect -199 3249 -165 3283
rect -335 3162 -301 3196
rect -267 3180 -233 3214
rect -199 3180 -165 3214
rect -335 3094 -301 3128
rect -267 3111 -233 3145
rect -199 3111 -165 3145
rect -335 3026 -301 3060
rect -267 3042 -233 3076
rect -199 3042 -165 3076
rect -335 2958 -301 2992
rect -267 2973 -233 3007
rect -199 2973 -165 3007
rect -335 2890 -301 2924
rect -267 2904 -233 2938
rect -199 2904 -165 2938
rect -335 2822 -301 2856
rect -267 2835 -233 2869
rect -199 2835 -165 2869
rect -335 2754 -301 2788
rect -267 2766 -233 2800
rect -199 2766 -165 2800
rect -335 2686 -301 2720
rect -267 2697 -233 2731
rect -199 2697 -165 2731
rect -335 2618 -301 2652
rect -267 2628 -233 2662
rect -199 2628 -165 2662
rect -335 2550 -301 2584
rect -267 2559 -233 2593
rect -199 2559 -165 2593
rect -335 2482 -301 2516
rect -267 2490 -233 2524
rect -199 2490 -165 2524
rect -335 2414 -301 2448
rect -267 2421 -233 2455
rect -199 2421 -165 2455
rect -335 2346 -301 2380
rect -267 2352 -233 2386
rect -199 2352 -165 2386
rect -335 2278 -301 2312
rect -267 2283 -233 2317
rect -199 2283 -165 2317
rect -335 2210 -301 2244
rect -267 2214 -233 2248
rect -199 2214 -165 2248
rect -335 2142 -301 2176
rect -267 2145 -233 2179
rect -199 2145 -165 2179
rect -335 2074 -301 2108
rect -267 2076 -233 2110
rect -199 2076 -165 2110
rect -335 2006 -301 2040
rect -267 2007 -233 2041
rect -199 2007 -165 2041
rect -335 1938 -301 1972
rect -267 1938 -233 1972
rect -199 1938 -165 1972
rect -335 1869 -301 1903
rect -267 1869 -233 1903
rect -199 1869 -165 1903
rect -335 1800 -301 1834
rect -267 1800 -233 1834
rect -199 1800 -165 1834
rect -335 1731 -301 1765
rect -267 1731 -233 1765
rect -199 1731 -165 1765
rect -335 1662 -301 1696
rect -267 1662 -233 1696
rect -199 1662 -165 1696
rect -335 1593 -301 1627
rect -267 1593 -233 1627
rect -199 1593 -165 1627
rect -335 1524 -301 1558
rect -267 1524 -233 1558
rect -199 1524 -165 1558
rect -335 1455 -301 1489
rect -267 1455 -233 1489
rect -199 1455 -165 1489
rect -335 1386 -301 1420
rect -267 1386 -233 1420
rect -199 1386 -165 1420
rect -335 1317 -301 1351
rect -267 1317 -233 1351
rect -199 1317 -165 1351
rect -335 1248 -301 1282
rect -267 1248 -233 1282
rect -199 1248 -165 1282
rect -335 1179 -301 1213
rect -267 1179 -233 1213
rect -199 1179 -165 1213
rect -335 1110 -301 1144
rect -267 1110 -233 1144
rect -199 1110 -165 1144
rect -335 1041 -301 1075
rect -267 1041 -233 1075
rect -199 1041 -165 1075
rect -335 972 -301 1006
rect -267 972 -233 1006
rect -199 972 -165 1006
rect -335 903 -301 937
rect -267 903 -233 937
rect -199 903 -165 937
rect -335 834 -301 868
rect -267 834 -233 868
rect -199 834 -165 868
rect -335 765 -301 799
rect -267 765 -233 799
rect -199 765 -165 799
rect -335 696 -301 730
rect -267 696 -233 730
rect -199 696 -165 730
rect -335 627 -301 661
rect -267 627 -233 661
rect -199 627 -165 661
rect -335 558 -301 592
rect -267 558 -233 592
rect -199 558 -165 592
rect -335 489 -301 523
rect -267 489 -233 523
rect -199 489 -165 523
rect -335 420 -301 454
rect -267 420 -233 454
rect -199 420 -165 454
rect -335 351 -301 385
rect -267 351 -233 385
rect -199 351 -165 385
rect -335 282 -301 316
rect -267 282 -233 316
rect -199 282 -165 316
rect -335 213 -301 247
rect -267 213 -233 247
rect -199 213 -165 247
rect -335 144 -301 178
rect -267 144 -233 178
rect -199 144 -165 178
rect 367 4168 401 4202
rect 435 4192 469 4226
rect 506 4192 540 4226
rect 577 4192 611 4226
rect 649 4192 683 4226
rect 721 4192 755 4226
rect 793 4192 827 4226
rect 865 4192 899 4226
rect 937 4192 971 4226
rect 1009 4192 1043 4226
rect 1081 4192 1115 4226
rect 1153 4192 1187 4226
rect 1225 4192 1259 4226
rect 1297 4192 1331 4226
rect 1369 4192 1403 4226
rect 1441 4192 1475 4226
rect 1513 4192 1547 4226
rect 1585 4192 1619 4226
rect 1657 4192 1691 4226
rect 367 4100 401 4134
rect 367 4032 401 4066
rect 1725 4168 1759 4202
rect 1725 4091 1759 4125
rect 367 3964 401 3998
rect 367 3896 401 3930
rect 367 3828 401 3862
rect 367 3760 401 3794
rect 367 3692 401 3726
rect 367 3624 401 3658
rect 367 3556 401 3590
rect 367 3488 401 3522
rect 367 3420 401 3454
rect 367 3352 401 3386
rect 1725 4014 1759 4048
rect 1725 3938 1759 3972
rect 1749 3870 1783 3904
rect 1817 3870 1851 3904
rect 1883 3870 1987 3904
rect 2021 3870 2055 3904
rect 2089 3870 2123 3904
rect 2157 3870 2191 3904
rect 2225 3870 2259 3904
rect 2293 3870 2327 3904
rect 2361 3870 2395 3904
rect 2429 3870 2463 3904
rect 2497 3870 2531 3904
rect 2565 3870 2599 3904
rect 2633 3870 2667 3904
rect 2701 3870 2735 3904
rect 2769 3870 2803 3904
rect 2837 3870 2871 3904
rect 2905 3870 2939 3904
rect 2973 3870 3007 3904
rect 3041 3870 3075 3904
rect 3109 3870 3143 3904
rect 3177 3870 3211 3904
rect 3245 3870 3279 3904
rect 3313 3870 3347 3904
rect 3381 3870 3415 3904
rect 3449 3870 3483 3904
rect 3517 3870 3551 3904
rect 3585 3870 3619 3904
rect 3653 3870 3687 3904
rect 3721 3870 3755 3904
rect 3789 3870 3823 3904
rect 3857 3870 3891 3904
rect 3925 3870 3959 3904
rect 3993 3870 4027 3904
rect 4062 3870 4096 3904
rect 4131 3870 4165 3904
rect 4200 3870 4234 3904
rect 4269 3870 4303 3904
rect 4338 3870 4372 3904
rect 4407 3870 4441 3904
rect 4476 3870 4510 3904
rect 4545 3870 4579 3904
rect 4614 3870 4648 3904
rect 4683 3870 4717 3904
rect 4752 3870 4786 3904
rect 4821 3870 4855 3904
rect 4890 3870 4924 3904
rect 4959 3870 4993 3904
rect 5028 3870 5062 3904
rect 5097 3870 5131 3904
rect 5166 3870 5200 3904
rect 5235 3870 5269 3904
rect 5304 3870 5338 3904
rect 5373 3870 5407 3904
rect 5442 3870 5476 3904
rect 5511 3870 5545 3904
rect 5580 3870 5614 3904
rect 5649 3870 5683 3904
rect 5718 3870 5752 3904
rect 5787 3870 5821 3904
rect 5856 3870 5890 3904
rect 5925 3870 5959 3904
rect 5994 3870 6028 3904
rect 6063 3870 6097 3904
rect 6132 3870 6166 3904
rect 6201 3870 6235 3904
rect 1883 3802 1985 3870
rect 1883 3731 1917 3765
rect 1951 3731 1985 3765
rect 6269 3846 6303 3880
rect 6269 3778 6303 3812
rect 1883 3660 1917 3694
rect 1951 3660 1985 3694
rect 1883 3589 1917 3623
rect 1951 3589 1985 3623
rect 1883 3518 1917 3552
rect 1951 3518 1985 3552
rect 1883 3447 1917 3481
rect 1951 3447 1985 3481
rect 6269 3710 6303 3744
rect 6269 3641 6303 3675
rect 6269 3572 6303 3606
rect 6269 3503 6303 3537
rect 1883 3376 1917 3410
rect 1951 3376 1985 3410
rect 367 3284 401 3318
rect 367 3216 401 3250
rect 1883 3305 1917 3339
rect 1951 3305 1985 3339
rect 6269 3434 6303 3468
rect 6269 3365 6303 3399
rect 1883 3234 1917 3268
rect 1951 3234 1985 3268
rect 367 3148 401 3182
rect 367 3080 401 3114
rect 1331 3147 1365 3181
rect 1399 3147 1433 3181
rect 1467 3147 1501 3181
rect 1535 3147 1569 3181
rect 1603 3147 1637 3181
rect 1883 3163 1917 3197
rect 1951 3163 1985 3197
rect 1331 3076 1365 3110
rect 1399 3076 1433 3110
rect 1467 3076 1501 3110
rect 1535 3073 1569 3107
rect 1603 3073 1637 3107
rect 1883 3092 1917 3126
rect 1951 3092 1985 3126
rect 367 3012 401 3046
rect 367 2944 401 2978
rect 367 2876 401 2910
rect 367 2808 401 2842
rect 1331 3005 1365 3039
rect 1399 3005 1433 3039
rect 1467 3005 1501 3039
rect 1535 2999 1569 3033
rect 1603 2999 1637 3033
rect 1883 3021 1917 3055
rect 1951 3021 1985 3055
rect 6269 3296 6303 3330
rect 6269 3227 6303 3261
rect 6269 3158 6303 3192
rect 6269 3089 6303 3123
rect 1331 2934 1365 2968
rect 1399 2934 1433 2968
rect 1467 2934 1501 2968
rect 1535 2925 1569 2959
rect 1603 2925 1637 2959
rect 1883 2950 1917 2984
rect 1951 2950 1985 2984
rect 1331 2863 1365 2897
rect 1399 2863 1433 2897
rect 1467 2863 1501 2897
rect 1535 2851 1569 2885
rect 1603 2851 1637 2885
rect 1883 2879 1917 2913
rect 1951 2879 1985 2913
rect 6269 3020 6303 3054
rect 6269 2951 6303 2985
rect 367 2740 401 2774
rect 1331 2792 1365 2826
rect 1399 2792 1433 2826
rect 1467 2792 1501 2826
rect 1535 2777 1569 2811
rect 1603 2777 1637 2811
rect 1883 2808 1917 2842
rect 1951 2808 1985 2842
rect 367 2672 401 2706
rect 367 2604 401 2638
rect 367 2536 401 2570
rect 367 2468 401 2502
rect 1331 2721 1365 2755
rect 1399 2721 1433 2755
rect 1467 2721 1501 2755
rect 1883 2737 1917 2771
rect 1951 2737 1985 2771
rect 1535 2703 1569 2737
rect 1603 2703 1637 2737
rect 1331 2650 1365 2684
rect 1399 2650 1433 2684
rect 1467 2650 1501 2684
rect 1883 2665 1917 2699
rect 1951 2665 1985 2699
rect 1535 2629 1569 2663
rect 1603 2629 1637 2663
rect 6269 2882 6303 2916
rect 6269 2813 6303 2847
rect 6269 2744 6303 2778
rect 6269 2675 6303 2709
rect 1331 2579 1365 2613
rect 1399 2579 1433 2613
rect 1467 2579 1501 2613
rect 1883 2593 1917 2627
rect 1951 2593 1985 2627
rect 1535 2555 1569 2589
rect 1603 2555 1637 2589
rect 1331 2508 1365 2542
rect 1399 2508 1433 2542
rect 1467 2508 1501 2542
rect 1883 2521 1917 2555
rect 1951 2521 1985 2555
rect 367 2400 401 2434
rect 1535 2481 1569 2515
rect 1603 2481 1637 2515
rect 6269 2606 6303 2640
rect 6269 2537 6303 2571
rect 1331 2437 1365 2471
rect 1399 2437 1433 2471
rect 1467 2437 1501 2471
rect 1883 2449 1917 2483
rect 1951 2449 1985 2483
rect 2207 2458 2241 2492
rect 2275 2458 2309 2492
rect 2343 2458 2377 2492
rect 2411 2458 2445 2492
rect 2479 2458 2513 2492
rect 2547 2458 2581 2492
rect 2615 2458 2649 2492
rect 2683 2458 2717 2492
rect 2751 2458 2785 2492
rect 2820 2458 2854 2492
rect 2889 2458 2923 2492
rect 2958 2458 2992 2492
rect 3027 2458 3061 2492
rect 3096 2458 3130 2492
rect 3165 2458 3199 2492
rect 3234 2458 3268 2492
rect 3303 2458 3337 2492
rect 3372 2458 3406 2492
rect 3441 2458 3475 2492
rect 3510 2458 3544 2492
rect 3579 2458 3613 2492
rect 3648 2458 3682 2492
rect 3717 2458 3751 2492
rect 3786 2458 3820 2492
rect 3855 2458 3889 2492
rect 3924 2458 3958 2492
rect 3993 2458 4027 2492
rect 4062 2458 4096 2492
rect 4131 2458 4165 2492
rect 4200 2458 4234 2492
rect 4269 2458 4303 2492
rect 4338 2458 4372 2492
rect 4407 2458 4441 2492
rect 4476 2458 4510 2492
rect 4545 2458 4579 2492
rect 4614 2458 4648 2492
rect 4683 2458 4717 2492
rect 4752 2458 4786 2492
rect 4821 2458 4855 2492
rect 4890 2458 4924 2492
rect 4959 2458 4993 2492
rect 5028 2458 5062 2492
rect 5097 2458 5131 2492
rect 5166 2458 5200 2492
rect 5235 2458 5269 2492
rect 5304 2458 5338 2492
rect 5373 2458 5407 2492
rect 5442 2458 5476 2492
rect 5511 2458 5545 2492
rect 5580 2458 5614 2492
rect 5649 2458 5683 2492
rect 5718 2458 5752 2492
rect 5787 2458 5821 2492
rect 5856 2458 5890 2492
rect 5925 2458 5959 2492
rect 5994 2458 6028 2492
rect 6063 2458 6097 2492
rect 6132 2458 6166 2492
rect 6201 2458 6235 2492
rect 6269 2468 6303 2502
rect 367 2332 401 2366
rect 367 2264 401 2298
rect 367 2196 401 2230
rect 367 2128 401 2162
rect 367 2060 401 2094
rect 367 1992 401 2026
rect 367 1924 401 1958
rect 367 1856 401 1890
rect 1535 2408 1569 2442
rect 1603 2408 1637 2442
rect 1331 2366 1365 2400
rect 1399 2366 1433 2400
rect 1467 2366 1501 2400
rect 1883 2377 1917 2411
rect 1951 2377 1985 2411
rect 1331 2294 1365 2328
rect 1399 2294 1433 2328
rect 1467 2294 1501 2328
rect 6269 2399 6303 2433
rect 6269 2330 6303 2364
rect 1331 2222 1365 2256
rect 1399 2222 1433 2256
rect 1467 2222 1501 2256
rect 1331 2150 1365 2184
rect 1399 2150 1433 2184
rect 1467 2150 1501 2184
rect 1331 2078 1365 2112
rect 1399 2078 1433 2112
rect 1467 2078 1501 2112
rect 1331 2006 1365 2040
rect 1399 2006 1433 2040
rect 1467 2006 1501 2040
rect 1331 1934 1365 1968
rect 1399 1934 1433 1968
rect 1467 1934 1501 1968
rect 1331 1862 1365 1896
rect 1399 1862 1433 1896
rect 1467 1862 1501 1896
rect 367 1788 401 1822
rect 367 1720 401 1754
rect 367 1652 401 1686
rect 367 1584 401 1618
rect 367 1516 401 1550
rect 367 1448 401 1482
rect 367 1380 401 1414
rect 367 1312 401 1346
rect 367 1244 401 1278
rect 367 1176 401 1210
rect 367 1108 401 1142
rect 367 1040 401 1074
rect 367 972 401 1006
rect 367 904 401 938
rect 367 836 401 870
rect 367 768 401 802
rect 367 699 401 733
rect 367 630 401 664
rect 367 561 401 595
rect 367 492 401 526
rect 1653 1226 2027 2144
rect 1653 1157 1687 1191
rect 1721 1157 1755 1191
rect 1789 1157 1823 1191
rect 1857 1157 1891 1191
rect 1925 1157 1959 1191
rect 1993 1157 2027 1191
rect 1653 1088 1687 1122
rect 1721 1088 1755 1122
rect 1789 1088 1823 1122
rect 1857 1088 1891 1122
rect 1925 1088 1959 1122
rect 1993 1088 2027 1122
rect 1653 1019 1687 1053
rect 1721 1019 1755 1053
rect 1789 1019 1823 1053
rect 1857 1019 1891 1053
rect 1925 1019 1959 1053
rect 1993 1019 2027 1053
rect 1653 950 1687 984
rect 1721 950 1755 984
rect 1789 950 1823 984
rect 1857 950 1891 984
rect 1925 950 1959 984
rect 1993 950 2027 984
rect 1653 881 1687 915
rect 1721 881 1755 915
rect 1789 881 1823 915
rect 1857 881 1891 915
rect 1925 881 1959 915
rect 1993 881 2027 915
rect 1653 812 1687 846
rect 1721 812 1755 846
rect 1789 812 1823 846
rect 1857 812 1891 846
rect 1925 812 1959 846
rect 1993 812 2027 846
rect 1653 743 1687 777
rect 1721 743 1755 777
rect 1789 743 1823 777
rect 1857 743 1891 777
rect 1925 743 1959 777
rect 1993 743 2027 777
rect 1653 674 1687 708
rect 1721 674 1755 708
rect 1789 674 1823 708
rect 1857 674 1891 708
rect 1925 674 1959 708
rect 1993 674 2027 708
rect 1653 605 1687 639
rect 1721 605 1755 639
rect 1789 605 1823 639
rect 1857 605 1891 639
rect 1925 605 1959 639
rect 1993 605 2027 639
rect 1653 536 1687 570
rect 1721 536 1755 570
rect 1789 536 1823 570
rect 1857 536 1891 570
rect 1925 536 1959 570
rect 1993 536 2027 570
rect 367 423 401 457
rect 367 354 401 388
rect 6269 2261 6303 2295
rect 6269 2192 6303 2226
rect 6269 2123 6303 2157
rect 6269 2054 6303 2088
rect 6269 1985 6303 2019
rect 6269 1916 6303 1950
rect 6269 1847 6303 1881
rect 6269 1778 6303 1812
rect 6269 1709 6303 1743
rect 6269 1640 6303 1674
rect 6269 1571 6303 1605
rect 6269 1502 6303 1536
rect 6269 1433 6303 1467
rect 6269 1364 6303 1398
rect 6269 1295 6303 1329
rect 6269 1226 6303 1260
rect 6269 1157 6303 1191
rect 6269 1088 6303 1122
rect 6269 1019 6303 1053
rect 6269 950 6303 984
rect 6269 881 6303 915
rect 6269 812 6303 846
rect 6269 743 6303 777
rect 6269 674 6303 708
rect 6269 605 6303 639
rect 6269 536 6303 570
rect 1653 467 1687 501
rect 1721 467 1755 501
rect 1789 467 1823 501
rect 1857 467 1891 501
rect 1925 467 1959 501
rect 1993 467 2027 501
rect 565 330 599 364
rect 633 330 667 364
rect 701 330 735 364
rect 769 330 803 364
rect 837 330 871 364
rect 905 330 939 364
rect 973 330 1007 364
rect 1041 330 1075 364
rect 1109 330 1143 364
rect 1177 330 1211 364
rect 1245 330 1279 364
rect 1313 330 1347 364
rect 1381 330 1415 364
rect 1449 330 1483 364
rect 1517 330 1551 364
rect 1585 330 1619 364
rect 1653 330 2027 432
rect 6269 467 6303 501
rect 6269 398 6303 432
rect 2061 330 2095 364
rect 2129 330 2163 364
rect 2197 330 2231 364
rect 2265 330 2299 364
rect 2333 330 2367 364
rect 2401 330 2435 364
rect 2469 330 2503 364
rect 2537 330 2571 364
rect 2605 330 2639 364
rect 2673 330 2707 364
rect 2741 330 2775 364
rect 2809 330 2843 364
rect 2877 330 2911 364
rect 2945 330 2979 364
rect 3013 330 3047 364
rect 3081 330 3115 364
rect 3149 330 3183 364
rect 3217 330 3251 364
rect 3285 330 3319 364
rect 3353 330 3387 364
rect 3421 330 3455 364
rect 3489 330 3523 364
rect 3557 330 3591 364
rect 3625 330 3659 364
rect 3693 330 3727 364
rect 3761 330 3795 364
rect 3830 330 3864 364
rect 3899 330 3933 364
rect 3968 330 4002 364
rect 4037 330 4071 364
rect 4106 330 4140 364
rect 4175 330 4209 364
rect 4244 330 4278 364
rect 4313 330 4347 364
rect 4382 330 4416 364
rect 4451 330 4485 364
rect 4520 330 4554 364
rect 4589 330 4623 364
rect 4658 330 4692 364
rect 4727 330 4761 364
rect 4796 330 4830 364
rect 4865 330 4899 364
rect 4934 330 4968 364
rect 5003 330 5037 364
rect 5072 330 5106 364
rect 5141 330 5175 364
rect 5210 330 5244 364
rect 5279 330 5313 364
rect 5348 330 5382 364
rect 5417 330 5451 364
rect 5486 330 5520 364
rect 5555 330 5589 364
rect 5624 330 5658 364
rect 5693 330 5727 364
rect 5762 330 5796 364
rect 5831 330 5865 364
rect 5900 330 5934 364
rect 5969 330 6003 364
rect 6038 330 6072 364
rect 6107 330 6141 364
rect 6176 330 6210 364
rect 6245 330 6279 364
rect 26285 6456 26319 6490
rect 26149 6421 26183 6455
rect 26217 6420 26251 6454
rect 26285 6388 26319 6422
rect 26149 6352 26183 6386
rect 26217 6351 26251 6385
rect 26285 6320 26319 6354
rect 26149 6283 26183 6317
rect 26217 6282 26251 6316
rect 26285 6252 26319 6286
rect 26149 6214 26183 6248
rect 26217 6213 26251 6247
rect 26285 6184 26319 6218
rect 26149 6145 26183 6179
rect 26217 6144 26251 6178
rect 26285 6116 26319 6150
rect 26149 6076 26183 6110
rect 26217 6075 26251 6109
rect 26285 6048 26319 6082
rect 26149 6007 26183 6041
rect 26217 6006 26251 6040
rect 26285 5980 26319 6014
rect 26149 5938 26183 5972
rect 26217 5937 26251 5971
rect 26285 5912 26319 5946
rect 26149 5869 26183 5903
rect 26217 5868 26251 5902
rect 26285 5844 26319 5878
rect 26149 5800 26183 5834
rect 26217 5799 26251 5833
rect 26285 5776 26319 5810
rect 26149 5731 26183 5765
rect 26217 5730 26251 5764
rect 26285 5708 26319 5742
rect 26149 5662 26183 5696
rect 26217 5661 26251 5695
rect 26285 5640 26319 5674
rect 26149 5593 26183 5627
rect 26217 5592 26251 5626
rect 26285 5572 26319 5606
rect 26149 5524 26183 5558
rect 26217 5523 26251 5557
rect 26285 5504 26319 5538
rect 26149 5455 26183 5489
rect 26217 5454 26251 5488
rect 26285 5436 26319 5470
rect 26149 5386 26183 5420
rect 26217 5385 26251 5419
rect 26285 5368 26319 5402
rect 26149 5317 26183 5351
rect 26217 5316 26251 5350
rect 26285 5300 26319 5334
rect 26149 5248 26183 5282
rect 26217 5247 26251 5281
rect 26285 5232 26319 5266
rect 26149 5179 26183 5213
rect 26217 5178 26251 5212
rect 26285 5164 26319 5198
rect 26149 5110 26183 5144
rect 26217 5109 26251 5143
rect 26285 5096 26319 5130
rect 26149 5041 26183 5075
rect 26217 5040 26251 5074
rect 26285 5028 26319 5062
rect 26149 4972 26183 5006
rect 26217 4971 26251 5005
rect 26285 4960 26319 4994
rect 26149 4903 26183 4937
rect 26217 4902 26251 4936
rect 26285 4892 26319 4926
rect 26149 4834 26183 4868
rect 26217 4833 26251 4867
rect 26285 4824 26319 4858
rect 26149 4765 26183 4799
rect 26217 4764 26251 4798
rect 26285 4756 26319 4790
rect 26149 4696 26183 4730
rect 26217 4695 26251 4729
rect 26285 4688 26319 4722
rect 26149 4627 26183 4661
rect 26217 4626 26251 4660
rect 26285 4620 26319 4654
rect 26149 4558 26183 4592
rect 26217 4557 26251 4591
rect 26285 4552 26319 4586
rect 26149 4489 26183 4523
rect 26217 4488 26251 4522
rect 26285 4484 26319 4518
rect 26149 4420 26183 4454
rect 26217 4419 26251 4453
rect 26285 4416 26319 4450
rect 26149 4351 26183 4385
rect 26217 4350 26251 4384
rect 26285 4348 26319 4382
rect 26149 4282 26183 4316
rect 26217 4281 26251 4315
rect 26285 4280 26319 4314
rect 26149 4213 26183 4247
rect 26217 4178 26319 4246
rect 26149 64 26319 4178
<< poly >>
rect 155 6053 221 6069
rect 155 6019 171 6053
rect 205 6019 221 6053
rect 155 5985 221 6019
rect 155 5951 171 5985
rect 205 5951 221 5985
rect 155 5917 221 5951
rect 155 5883 171 5917
rect 205 5883 221 5917
rect 155 5849 221 5883
rect 155 5815 171 5849
rect 205 5815 221 5849
rect 155 5781 221 5815
rect 155 5747 171 5781
rect 205 5747 221 5781
rect 155 5713 221 5747
rect 155 5679 171 5713
rect 205 5679 221 5713
rect 155 5645 221 5679
rect 155 5611 171 5645
rect 205 5611 221 5645
rect 155 5577 221 5611
rect 155 5543 171 5577
rect 205 5543 221 5577
rect 155 5509 221 5543
rect 155 5475 171 5509
rect 205 5475 221 5509
rect 155 5441 221 5475
rect 155 5407 171 5441
rect 205 5407 221 5441
rect 155 5391 221 5407
rect 1513 4037 1585 4053
rect 1513 4003 1535 4037
rect 1569 4003 1585 4037
rect 1513 3969 1585 4003
rect 1513 3953 1535 3969
rect 1519 3935 1535 3953
rect 1569 3935 1585 3969
rect 1519 3901 1585 3935
rect 1519 3897 1535 3901
rect 1513 3867 1535 3897
rect 1569 3867 1585 3901
rect 1513 3833 1585 3867
rect 1513 3799 1535 3833
rect 1569 3799 1585 3833
rect 1513 3765 1585 3799
rect 1513 3731 1535 3765
rect 1569 3731 1585 3765
rect 1513 3697 1585 3731
rect 1513 3663 1535 3697
rect 1569 3663 1585 3697
rect 1513 3629 1585 3663
rect 1513 3595 1535 3629
rect 1569 3595 1585 3629
rect 1513 3561 1585 3595
rect 1513 3531 1535 3561
rect 1519 3527 1535 3531
rect 1569 3527 1585 3561
rect 1519 3493 1585 3527
rect 1519 3475 1535 3493
rect 1513 3459 1535 3475
rect 1569 3459 1585 3493
rect 1513 3425 1585 3459
rect 1513 3391 1535 3425
rect 1569 3391 1585 3425
rect 1513 3375 1585 3391
rect 2085 3715 2157 3731
rect 2085 3681 2101 3715
rect 2135 3681 2157 3715
rect 2085 3631 2157 3681
rect 2085 3620 2151 3631
rect 2085 3586 2101 3620
rect 2135 3586 2151 3620
rect 2085 3575 2151 3586
rect 2085 3525 2157 3575
rect 2085 3491 2101 3525
rect 2135 3491 2157 3525
rect 2085 3475 2157 3491
rect 1227 3213 1293 3229
rect 1227 3209 1243 3213
rect 1221 3179 1243 3209
rect 1277 3179 1293 3213
rect 1221 3145 1293 3179
rect 1221 3111 1243 3145
rect 1277 3111 1293 3145
rect 1221 3109 1293 3111
rect 1227 3095 1293 3109
rect 1221 3037 1293 3053
rect 1221 3003 1243 3037
rect 1277 3003 1293 3037
rect 1221 2953 1293 3003
rect 1227 2942 1293 2953
rect 1227 2908 1243 2942
rect 1277 2908 1293 2942
rect 1227 2897 1293 2908
rect 1221 2847 1293 2897
rect 1221 2813 1243 2847
rect 1277 2813 1293 2847
rect 1221 2797 1293 2813
rect 2085 3293 2157 3309
rect 2085 3259 2101 3293
rect 2135 3259 2157 3293
rect 2085 3209 2157 3259
rect 2085 3198 2151 3209
rect 2085 3164 2101 3198
rect 2135 3164 2151 3198
rect 2085 3153 2151 3164
rect 2085 3103 2157 3153
rect 2085 3069 2101 3103
rect 2135 3069 2157 3103
rect 2085 3053 2157 3069
rect 1221 2725 1293 2741
rect 1221 2691 1243 2725
rect 1277 2691 1293 2725
rect 1221 2641 1293 2691
rect 1227 2630 1293 2641
rect 1227 2596 1243 2630
rect 1277 2596 1293 2630
rect 1227 2585 1293 2596
rect 1221 2535 1293 2585
rect 1221 2501 1243 2535
rect 1277 2501 1293 2535
rect 1221 2485 1293 2501
rect 2085 2871 2157 2887
rect 2085 2837 2101 2871
rect 2135 2837 2157 2871
rect 2085 2787 2157 2837
rect 2085 2776 2151 2787
rect 2085 2742 2101 2776
rect 2135 2742 2151 2776
rect 2085 2731 2151 2742
rect 2085 2681 2157 2731
rect 2085 2647 2101 2681
rect 2135 2647 2157 2681
rect 2085 2631 2157 2647
rect 1221 2413 1293 2429
rect 1221 2379 1243 2413
rect 1277 2379 1293 2413
rect 1221 2341 1293 2379
rect 1221 2329 1243 2341
rect 1227 2307 1243 2329
rect 1277 2307 1293 2341
rect 1227 2273 1293 2307
rect 1221 2269 1293 2273
rect 1221 2235 1243 2269
rect 1277 2235 1293 2269
rect 1221 2197 1293 2235
rect 1221 2173 1243 2197
rect 1227 2163 1243 2173
rect 1277 2163 1293 2197
rect 1227 2125 1293 2163
rect 1227 2117 1243 2125
rect 1221 2091 1243 2117
rect 1277 2091 1293 2125
rect 1221 2053 1293 2091
rect 1221 2019 1243 2053
rect 1277 2019 1293 2053
rect 1221 2017 1293 2019
rect 1227 1982 1293 2017
rect 1227 1961 1243 1982
rect 1221 1948 1243 1961
rect 1277 1948 1293 1982
rect 1221 1911 1293 1948
rect 1221 1877 1243 1911
rect 1277 1877 1293 1911
rect 1221 1861 1293 1877
rect 1513 1679 1585 1695
rect 1513 1645 1535 1679
rect 1569 1645 1585 1679
rect 1513 1608 1585 1645
rect 1513 1595 1535 1608
rect 1519 1574 1535 1595
rect 1569 1574 1585 1608
rect 1519 1539 1585 1574
rect 1513 1537 1585 1539
rect 1513 1503 1535 1537
rect 1569 1503 1585 1537
rect 1513 1466 1585 1503
rect 1513 1439 1535 1466
rect 1519 1432 1535 1439
rect 1569 1432 1585 1466
rect 1519 1395 1585 1432
rect 1519 1383 1535 1395
rect 1513 1361 1535 1383
rect 1569 1361 1585 1395
rect 1513 1324 1585 1361
rect 1513 1290 1535 1324
rect 1569 1290 1585 1324
rect 1513 1283 1585 1290
rect 1519 1253 1585 1283
rect 1519 1227 1535 1253
rect 1513 1219 1535 1227
rect 1569 1219 1585 1253
rect 1513 1183 1585 1219
rect 1513 1149 1535 1183
rect 1569 1149 1585 1183
rect 1513 1127 1585 1149
rect 1519 1113 1585 1127
rect 1519 1079 1535 1113
rect 1569 1079 1585 1113
rect 1519 1071 1585 1079
rect 1513 1043 1585 1071
rect 1513 1009 1535 1043
rect 1569 1009 1585 1043
rect 1513 973 1585 1009
rect 1513 971 1535 973
rect 1519 939 1535 971
rect 1569 939 1585 973
rect 1519 915 1585 939
rect 1513 903 1585 915
rect 1513 869 1535 903
rect 1569 869 1585 903
rect 1513 833 1585 869
rect 1513 815 1535 833
rect 1519 799 1535 815
rect 1569 799 1585 833
rect 1519 763 1585 799
rect 1519 759 1535 763
rect 1513 729 1535 759
rect 1569 729 1585 763
rect 1513 693 1585 729
rect 1513 659 1535 693
rect 1569 659 1585 693
rect 1519 623 1585 659
rect 1519 603 1535 623
rect 1513 589 1535 603
rect 1569 589 1585 623
rect 1513 553 1585 589
rect 1513 519 1535 553
rect 1569 519 1585 553
rect 1513 503 1585 519
rect 2085 2303 2157 2319
rect 2085 2269 2101 2303
rect 2135 2269 2157 2303
rect 2085 2233 2157 2269
rect 2085 2199 2101 2233
rect 2135 2219 2157 2233
rect 2135 2199 2151 2219
rect 2085 2163 2151 2199
rect 2085 2129 2101 2163
rect 2135 2129 2157 2163
rect 2085 2093 2157 2129
rect 2085 2059 2101 2093
rect 2135 2063 2157 2093
rect 2135 2059 2151 2063
rect 2085 2023 2151 2059
rect 2085 1989 2101 2023
rect 2135 2007 2151 2023
rect 2135 1989 2157 2007
rect 2085 1953 2157 1989
rect 2085 1919 2101 1953
rect 2135 1919 2157 1953
rect 2085 1907 2157 1919
rect 2085 1883 2151 1907
rect 2085 1849 2101 1883
rect 2135 1851 2151 1883
rect 2135 1849 2157 1851
rect 2085 1813 2157 1849
rect 2085 1779 2101 1813
rect 2135 1779 2157 1813
rect 2085 1751 2157 1779
rect 2085 1743 2151 1751
rect 2085 1709 2101 1743
rect 2135 1709 2151 1743
rect 2085 1695 2151 1709
rect 2085 1673 2157 1695
rect 2085 1639 2101 1673
rect 2135 1639 2157 1673
rect 2085 1603 2157 1639
rect 2085 1569 2101 1603
rect 2135 1595 2157 1603
rect 2135 1569 2151 1595
rect 2085 1539 2151 1569
rect 2085 1533 2157 1539
rect 2085 1499 2101 1533
rect 2135 1499 2157 1533
rect 2085 1463 2157 1499
rect 2085 1429 2101 1463
rect 2135 1439 2157 1463
rect 2135 1429 2151 1439
rect 2085 1393 2151 1429
rect 2085 1359 2101 1393
rect 2135 1383 2151 1393
rect 2135 1359 2157 1383
rect 2085 1323 2157 1359
rect 2085 1289 2101 1323
rect 2135 1289 2157 1323
rect 2085 1283 2157 1289
rect 2085 1253 2151 1283
rect 2085 1219 2101 1253
rect 2135 1227 2151 1253
rect 2135 1219 2157 1227
rect 2085 1183 2157 1219
rect 2085 1149 2101 1183
rect 2135 1149 2157 1183
rect 2085 1127 2157 1149
rect 2085 1113 2151 1127
rect 2085 1079 2101 1113
rect 2135 1079 2151 1113
rect 2085 1071 2151 1079
rect 2085 1043 2157 1071
rect 2085 1009 2101 1043
rect 2135 1009 2157 1043
rect 2085 973 2157 1009
rect 2085 939 2101 973
rect 2135 971 2157 973
rect 2135 939 2151 971
rect 2085 915 2151 939
rect 2085 903 2157 915
rect 2085 869 2101 903
rect 2135 869 2157 903
rect 2085 833 2157 869
rect 2085 799 2101 833
rect 2135 815 2157 833
rect 2135 799 2151 815
rect 2085 763 2151 799
rect 2085 729 2101 763
rect 2135 759 2151 763
rect 2135 729 2157 759
rect 2085 693 2157 729
rect 2085 659 2101 693
rect 2135 659 2157 693
rect 2085 623 2151 659
rect 2085 589 2101 623
rect 2135 603 2151 623
rect 2135 589 2157 603
rect 2085 553 2157 589
rect 2085 519 2101 553
rect 2135 519 2157 553
rect 2085 503 2157 519
<< polycont >>
rect 171 6019 205 6053
rect 171 5951 205 5985
rect 171 5883 205 5917
rect 171 5815 205 5849
rect 171 5747 205 5781
rect 171 5679 205 5713
rect 171 5611 205 5645
rect 171 5543 205 5577
rect 171 5475 205 5509
rect 171 5407 205 5441
rect 1535 4003 1569 4037
rect 1535 3935 1569 3969
rect 1535 3867 1569 3901
rect 1535 3799 1569 3833
rect 1535 3731 1569 3765
rect 1535 3663 1569 3697
rect 1535 3595 1569 3629
rect 1535 3527 1569 3561
rect 1535 3459 1569 3493
rect 1535 3391 1569 3425
rect 2101 3681 2135 3715
rect 2101 3586 2135 3620
rect 2101 3491 2135 3525
rect 1243 3179 1277 3213
rect 1243 3111 1277 3145
rect 1243 3003 1277 3037
rect 1243 2908 1277 2942
rect 1243 2813 1277 2847
rect 2101 3259 2135 3293
rect 2101 3164 2135 3198
rect 2101 3069 2135 3103
rect 1243 2691 1277 2725
rect 1243 2596 1277 2630
rect 1243 2501 1277 2535
rect 2101 2837 2135 2871
rect 2101 2742 2135 2776
rect 2101 2647 2135 2681
rect 1243 2379 1277 2413
rect 1243 2307 1277 2341
rect 1243 2235 1277 2269
rect 1243 2163 1277 2197
rect 1243 2091 1277 2125
rect 1243 2019 1277 2053
rect 1243 1948 1277 1982
rect 1243 1877 1277 1911
rect 1535 1645 1569 1679
rect 1535 1574 1569 1608
rect 1535 1503 1569 1537
rect 1535 1432 1569 1466
rect 1535 1361 1569 1395
rect 1535 1290 1569 1324
rect 1535 1219 1569 1253
rect 1535 1149 1569 1183
rect 1535 1079 1569 1113
rect 1535 1009 1569 1043
rect 1535 939 1569 973
rect 1535 869 1569 903
rect 1535 799 1569 833
rect 1535 729 1569 763
rect 1535 659 1569 693
rect 1535 589 1569 623
rect 1535 519 1569 553
rect 2101 2269 2135 2303
rect 2101 2199 2135 2233
rect 2101 2129 2135 2163
rect 2101 2059 2135 2093
rect 2101 1989 2135 2023
rect 2101 1919 2135 1953
rect 2101 1849 2135 1883
rect 2101 1779 2135 1813
rect 2101 1709 2135 1743
rect 2101 1639 2135 1673
rect 2101 1569 2135 1603
rect 2101 1499 2135 1533
rect 2101 1429 2135 1463
rect 2101 1359 2135 1393
rect 2101 1289 2135 1323
rect 2101 1219 2135 1253
rect 2101 1149 2135 1183
rect 2101 1079 2135 1113
rect 2101 1009 2135 1043
rect 2101 939 2135 973
rect 2101 869 2135 903
rect 2101 799 2135 833
rect 2101 729 2135 763
rect 2101 659 2135 693
rect 2101 589 2135 623
rect 2101 519 2135 553
<< locali >>
rect -335 6594 -311 6798
rect 1083 6764 1118 6798
rect 1152 6766 1187 6798
rect 1221 6766 1289 6798
rect 1323 6766 1358 6798
rect 1392 6766 1427 6798
rect 1461 6766 1496 6798
rect 1530 6766 1565 6798
rect 1599 6766 1634 6798
rect 1668 6766 1703 6798
rect 1156 6764 1187 6766
rect 1083 6732 1122 6764
rect 1156 6732 1195 6764
rect 1229 6732 1268 6766
rect 1323 6764 1341 6766
rect 1392 6764 1413 6766
rect 1461 6764 1485 6766
rect 1530 6764 1557 6766
rect 1599 6764 1629 6766
rect 1668 6764 1701 6766
rect 1737 6764 1772 6798
rect 1806 6766 1841 6798
rect 1875 6766 1910 6798
rect 1944 6766 1978 6798
rect 2012 6766 2046 6798
rect 2148 6766 2183 6798
rect 2217 6766 2252 6798
rect 2286 6766 2321 6798
rect 2355 6766 2390 6798
rect 2424 6766 2459 6798
rect 1807 6764 1841 6766
rect 1879 6764 1910 6766
rect 1951 6764 1978 6766
rect 1302 6732 1341 6764
rect 1375 6732 1413 6764
rect 1447 6732 1485 6764
rect 1519 6732 1557 6764
rect 1591 6732 1629 6764
rect 1663 6732 1701 6764
rect 1735 6732 1773 6764
rect 1807 6732 1845 6764
rect 1879 6732 1917 6764
rect 1951 6732 1989 6764
rect 2023 6732 2046 6766
rect 2167 6764 2183 6766
rect 2239 6764 2252 6766
rect 2311 6764 2321 6766
rect 2383 6764 2390 6766
rect 2455 6764 2459 6766
rect 2493 6766 2528 6798
rect 2167 6732 2205 6764
rect 2239 6732 2277 6764
rect 2311 6732 2349 6764
rect 2383 6732 2421 6764
rect 2455 6732 2493 6764
rect 2527 6764 2528 6766
rect 2562 6766 2597 6798
rect 2631 6766 2666 6798
rect 2700 6766 2735 6798
rect 2769 6766 2804 6798
rect 2838 6766 2873 6798
rect 2907 6766 2942 6798
rect 2976 6766 3011 6798
rect 3045 6766 3080 6798
rect 3114 6766 3149 6798
rect 3183 6766 3218 6798
rect 3252 6766 3287 6798
rect 2562 6764 2565 6766
rect 2631 6764 2637 6766
rect 2700 6764 2709 6766
rect 2769 6764 2781 6766
rect 2838 6764 2853 6766
rect 2907 6764 2925 6766
rect 2976 6764 2997 6766
rect 3045 6764 3069 6766
rect 3114 6764 3141 6766
rect 3183 6764 3213 6766
rect 3252 6764 3285 6766
rect 3321 6764 3356 6798
rect 3390 6766 3425 6798
rect 3459 6766 3494 6798
rect 3528 6766 3563 6798
rect 3597 6766 3632 6798
rect 3666 6766 3701 6798
rect 3735 6766 3770 6798
rect 3804 6766 3839 6798
rect 3873 6766 3908 6798
rect 3942 6766 3977 6798
rect 4011 6766 4046 6798
rect 4080 6766 4115 6798
rect 3391 6764 3425 6766
rect 3463 6764 3494 6766
rect 3535 6764 3563 6766
rect 3607 6764 3632 6766
rect 3679 6764 3701 6766
rect 3751 6764 3770 6766
rect 3823 6764 3839 6766
rect 3895 6764 3908 6766
rect 3967 6764 3977 6766
rect 4039 6764 4046 6766
rect 4111 6764 4115 6766
rect 4149 6766 4184 6798
rect 4218 6766 4253 6798
rect 4287 6766 4322 6798
rect 4356 6766 4391 6798
rect 4425 6766 4460 6798
rect 4494 6766 4529 6798
rect 4563 6766 4598 6798
rect 4632 6766 4667 6798
rect 4701 6766 4736 6798
rect 4770 6766 4805 6798
rect 4839 6766 4874 6798
rect 4908 6766 4943 6798
rect 4977 6766 5012 6798
rect 5046 6766 5081 6798
rect 5115 6766 5150 6798
rect 5184 6766 5219 6798
rect 5253 6766 5288 6798
rect 5322 6766 5357 6798
rect 5391 6766 5426 6798
rect 5460 6766 5495 6798
rect 5529 6766 5564 6798
rect 5598 6766 5633 6798
rect 5667 6766 5702 6798
rect 5736 6766 5771 6798
rect 5805 6766 5840 6798
rect 5874 6766 5909 6798
rect 5943 6766 5978 6798
rect 6012 6766 6047 6798
rect 6081 6766 6116 6798
rect 6150 6766 6185 6798
rect 6219 6766 6254 6798
rect 6288 6766 6323 6798
rect 6357 6766 6392 6798
rect 6426 6766 6461 6798
rect 6495 6766 6530 6798
rect 6564 6766 6599 6798
rect 2527 6732 2565 6764
rect 2599 6732 2637 6764
rect 2671 6732 2709 6764
rect 2743 6732 2781 6764
rect 2815 6732 2853 6764
rect 2887 6732 2925 6764
rect 2959 6732 2997 6764
rect 3031 6732 3069 6764
rect 3103 6732 3141 6764
rect 3175 6732 3213 6764
rect 3247 6732 3285 6764
rect 3319 6732 3357 6764
rect 3391 6732 3429 6764
rect 3463 6732 3501 6764
rect 3535 6732 3573 6764
rect 3607 6732 3645 6764
rect 3679 6732 3717 6764
rect 3751 6732 3789 6764
rect 3823 6732 3861 6764
rect 3895 6732 3933 6764
rect 3967 6732 4005 6764
rect 4039 6732 4077 6764
rect 4111 6732 4149 6764
rect 1083 6730 2046 6732
rect 1083 6696 1118 6730
rect 1152 6696 1187 6730
rect 1221 6696 1323 6730
rect 1357 6696 1396 6730
rect 1430 6696 1469 6730
rect 1503 6696 1542 6730
rect 1576 6696 1614 6730
rect 1648 6696 1686 6730
rect 1720 6696 1758 6730
rect 1792 6696 1830 6730
rect 1864 6696 1902 6730
rect 1936 6696 1974 6730
rect 2008 6696 2046 6730
rect 1083 6694 2046 6696
rect 2148 6730 4149 6732
rect 26217 6764 26319 6798
rect 26217 6760 26285 6764
rect 2148 6696 2183 6730
rect 2217 6696 2252 6730
rect 2286 6696 2321 6730
rect 2355 6696 2390 6730
rect 2424 6696 2459 6730
rect 2493 6696 2528 6730
rect 2562 6696 2597 6730
rect 2631 6696 2666 6730
rect 2700 6696 2735 6730
rect 2769 6696 2804 6730
rect 2838 6696 2873 6730
rect 2907 6696 2942 6730
rect 2976 6696 3011 6730
rect 3045 6696 3080 6730
rect 3114 6696 3149 6730
rect 3183 6696 3218 6730
rect 3252 6696 3287 6730
rect 3321 6696 3356 6730
rect 3390 6696 3425 6730
rect 3459 6696 3494 6730
rect 3528 6696 3563 6730
rect 3597 6696 3632 6730
rect 3666 6696 3701 6730
rect 3735 6696 3770 6730
rect 3804 6696 3839 6730
rect 3873 6696 3908 6730
rect 3942 6696 3977 6730
rect 4011 6696 4046 6730
rect 4080 6696 4115 6730
rect 2148 6694 4149 6696
rect 1117 6662 1156 6694
rect 1190 6662 1229 6694
rect 1263 6692 1302 6694
rect 1117 6660 1118 6662
rect 1083 6628 1118 6660
rect 1152 6660 1156 6662
rect 1221 6660 1229 6662
rect 1289 6660 1302 6692
rect 1336 6661 1375 6694
rect 1409 6662 1448 6694
rect 1482 6662 1521 6694
rect 1555 6662 1594 6694
rect 1628 6662 1667 6694
rect 1701 6662 1740 6694
rect 1774 6662 1813 6694
rect 1847 6662 1886 6694
rect 1920 6662 1959 6694
rect 1993 6662 2032 6694
rect 1357 6660 1375 6661
rect 1425 6660 1448 6662
rect 1498 6660 1521 6662
rect 1571 6660 1594 6662
rect 1644 6660 1667 6662
rect 1717 6660 1740 6662
rect 1790 6660 1813 6662
rect 1863 6660 1886 6662
rect 1936 6660 1959 6662
rect 2008 6660 2032 6662
rect 2148 6660 2178 6694
rect 2212 6662 2251 6694
rect 2285 6662 2324 6694
rect 2358 6662 2397 6694
rect 2431 6662 2470 6694
rect 2504 6662 2543 6694
rect 2577 6662 2616 6694
rect 2650 6662 2689 6694
rect 2723 6662 2762 6694
rect 2796 6662 2835 6694
rect 2869 6662 2908 6694
rect 2217 6660 2251 6662
rect 1152 6628 1187 6660
rect 1221 6658 1255 6660
rect 1289 6658 1323 6660
rect 1221 6628 1323 6658
rect -335 6525 -303 6560
rect -335 6456 -303 6491
rect 1255 6627 1323 6628
rect 1357 6628 1391 6660
rect 1425 6628 1464 6660
rect 1498 6628 1537 6660
rect 1571 6628 1610 6660
rect 1644 6628 1683 6660
rect 1717 6628 1756 6660
rect 1790 6628 1829 6660
rect 1863 6628 1902 6660
rect 1936 6628 1974 6660
rect 2008 6628 2046 6660
rect 2148 6628 2183 6660
rect 2217 6628 2252 6660
rect 2286 6628 2321 6662
rect 2358 6660 2390 6662
rect 2431 6660 2459 6662
rect 2504 6660 2528 6662
rect 2577 6660 2597 6662
rect 2650 6660 2666 6662
rect 2723 6660 2735 6662
rect 2796 6660 2804 6662
rect 2869 6660 2873 6662
rect 2355 6628 2390 6660
rect 2424 6628 2459 6660
rect 2493 6628 2528 6660
rect 2562 6628 2597 6660
rect 2631 6628 2666 6660
rect 2700 6628 2735 6660
rect 2769 6628 2804 6660
rect 2838 6628 2873 6660
rect 2907 6660 2908 6662
rect 2942 6662 2981 6694
rect 3015 6662 3054 6694
rect 3088 6662 3127 6694
rect 3161 6662 3200 6694
rect 3234 6662 3273 6694
rect 3307 6662 3346 6694
rect 3380 6662 3419 6694
rect 3453 6662 3492 6694
rect 3526 6662 3565 6694
rect 3599 6662 3638 6694
rect 3672 6662 3711 6694
rect 3745 6662 3784 6694
rect 3818 6662 3857 6694
rect 3891 6662 3930 6694
rect 3964 6662 4003 6694
rect 4037 6662 4076 6694
rect 4110 6662 4149 6694
rect 2907 6628 2942 6660
rect 2976 6660 2981 6662
rect 3045 6660 3054 6662
rect 3114 6660 3127 6662
rect 3183 6660 3200 6662
rect 3252 6660 3273 6662
rect 3321 6660 3346 6662
rect 3390 6660 3419 6662
rect 3459 6660 3492 6662
rect 2976 6628 3011 6660
rect 3045 6628 3080 6660
rect 3114 6628 3149 6660
rect 3183 6628 3218 6660
rect 3252 6628 3287 6660
rect 3321 6628 3356 6660
rect 3390 6628 3425 6660
rect 3459 6628 3494 6660
rect 3528 6628 3563 6662
rect 3599 6660 3632 6662
rect 3672 6660 3701 6662
rect 3745 6660 3770 6662
rect 3818 6660 3839 6662
rect 3891 6660 3908 6662
rect 3964 6660 3977 6662
rect 4037 6660 4046 6662
rect 4110 6660 4115 6662
rect 3597 6628 3632 6660
rect 3666 6628 3701 6660
rect 3735 6628 3770 6660
rect 3804 6628 3839 6660
rect 3873 6628 3908 6660
rect 3942 6628 3977 6660
rect 4011 6628 4046 6660
rect 4080 6628 4115 6660
rect 26217 6730 26253 6760
rect 26251 6726 26253 6730
rect 26287 6726 26319 6730
rect 26251 6696 26319 6726
rect 26183 6695 26319 6696
rect 26183 6687 26285 6695
rect 4149 6628 4184 6660
rect 4218 6628 4253 6660
rect 26215 6661 26253 6687
rect 26215 6653 26217 6661
rect 26183 6628 26217 6653
rect 1357 6627 1425 6628
rect 1255 6622 1425 6627
rect 1393 6592 1425 6622
rect 1255 6552 1287 6588
rect 25 6464 66 6490
rect 100 6464 141 6490
rect 175 6464 216 6490
rect 250 6464 291 6490
rect 325 6464 365 6490
rect 399 6464 439 6490
rect 473 6464 513 6490
rect -335 6387 -303 6422
rect -335 6318 -303 6353
rect -335 6249 -303 6284
rect -335 6180 -303 6215
rect -335 6111 -303 6146
rect -335 6042 -303 6077
rect -335 5973 -303 6008
rect -335 5904 -303 5939
rect -335 5835 -303 5870
rect -335 5766 -303 5801
rect -335 5697 -303 5732
rect -335 5628 -303 5663
rect -335 5558 -303 5594
rect -335 5488 -303 5524
rect -335 5418 -303 5454
rect -335 5348 -303 5384
rect -335 5278 -303 5314
rect -335 5208 -303 5244
rect -335 5138 -303 5174
rect -335 5068 -303 5104
rect -47 6430 -23 6464
rect 25 6456 49 6464
rect 100 6456 121 6464
rect 175 6456 193 6464
rect 250 6456 264 6464
rect 325 6456 335 6464
rect 399 6456 406 6464
rect 473 6456 477 6464
rect 11 6430 49 6456
rect 83 6430 121 6456
rect 155 6430 193 6456
rect 227 6430 264 6456
rect 298 6430 335 6456
rect 369 6430 406 6456
rect 440 6430 477 6456
rect 511 6456 513 6464
rect 547 6464 587 6490
rect 621 6464 661 6490
rect 695 6464 735 6490
rect 769 6464 809 6490
rect 843 6464 883 6490
rect 917 6464 957 6490
rect 991 6464 1031 6490
rect 1255 6482 1287 6518
rect 1393 6522 1425 6558
rect 547 6456 548 6464
rect 511 6430 548 6456
rect 582 6456 587 6464
rect 653 6456 661 6464
rect 724 6456 735 6464
rect 795 6456 809 6464
rect 866 6456 883 6464
rect 937 6456 957 6464
rect 1008 6456 1031 6464
rect 582 6430 619 6456
rect 653 6430 690 6456
rect 724 6430 761 6456
rect 795 6430 832 6456
rect 866 6430 903 6456
rect 937 6430 974 6456
rect 1008 6430 1045 6456
rect 1079 6430 1103 6464
rect -47 6418 1103 6430
rect -47 6384 -9 6418
rect 25 6384 66 6418
rect 100 6384 141 6418
rect 175 6384 216 6418
rect 250 6384 291 6418
rect 325 6384 365 6418
rect 399 6384 439 6418
rect 473 6384 513 6418
rect 547 6384 587 6418
rect 621 6384 661 6418
rect 695 6384 735 6418
rect 769 6384 809 6418
rect 843 6384 883 6418
rect 917 6384 957 6418
rect 991 6384 1031 6418
rect 1065 6384 1103 6418
rect -47 6378 1103 6384
rect -47 6346 57 6378
rect -47 6344 23 6346
rect -13 6312 23 6344
rect 91 6346 126 6378
rect 160 6346 195 6378
rect 229 6346 265 6378
rect 299 6346 335 6378
rect 369 6346 405 6378
rect 439 6346 475 6378
rect 91 6344 98 6346
rect 160 6344 173 6346
rect 229 6344 248 6346
rect 299 6344 323 6346
rect 369 6344 398 6346
rect 439 6344 473 6346
rect 509 6344 545 6378
rect 579 6346 615 6378
rect 649 6346 685 6378
rect 719 6346 755 6378
rect 789 6346 825 6378
rect 859 6346 895 6378
rect 929 6346 965 6378
rect 582 6344 615 6346
rect 657 6344 685 6346
rect 732 6344 755 6346
rect 807 6344 825 6346
rect 882 6344 895 6346
rect 957 6344 965 6346
rect 999 6344 1035 6378
rect 1069 6344 1103 6378
rect 57 6312 98 6344
rect 132 6312 173 6344
rect 207 6312 248 6344
rect 282 6312 323 6344
rect 357 6312 398 6344
rect 432 6312 473 6344
rect 507 6312 548 6344
rect 582 6312 623 6344
rect 657 6312 698 6344
rect 732 6312 773 6344
rect 807 6312 848 6344
rect 882 6312 923 6344
rect 957 6312 1103 6344
rect -13 6310 1103 6312
rect -47 6276 21 6310
rect 55 6276 91 6310
rect 125 6276 161 6310
rect 195 6276 231 6310
rect 265 6276 301 6310
rect 335 6276 371 6310
rect 405 6276 441 6310
rect 475 6276 511 6310
rect 545 6276 581 6310
rect 615 6276 651 6310
rect 685 6276 721 6310
rect 755 6276 791 6310
rect 825 6276 861 6310
rect 895 6276 931 6310
rect 965 6276 1001 6310
rect 1035 6308 1103 6310
rect 1035 6276 1037 6308
rect -47 6274 1037 6276
rect 1071 6274 1103 6308
rect -47 6273 57 6274
rect -13 6240 57 6273
rect 91 6242 133 6274
rect 167 6242 209 6274
rect 243 6242 285 6274
rect 319 6242 361 6274
rect 395 6242 437 6274
rect 471 6242 513 6274
rect 547 6242 589 6274
rect 623 6242 665 6274
rect 699 6242 740 6274
rect 774 6242 815 6274
rect 849 6242 890 6274
rect 924 6242 965 6274
rect 999 6272 1103 6274
rect 123 6240 133 6242
rect 193 6240 209 6242
rect 263 6240 285 6242
rect 333 6240 361 6242
rect 403 6240 437 6242
rect -13 6239 89 6240
rect -47 6237 89 6239
rect -47 6234 21 6237
rect -47 6202 -15 6234
rect 19 6203 21 6234
rect 55 6208 89 6237
rect 123 6208 159 6240
rect 193 6208 229 6240
rect 263 6208 299 6240
rect 333 6208 369 6240
rect 403 6208 439 6240
rect 473 6208 509 6242
rect 547 6240 579 6242
rect 623 6240 649 6242
rect 699 6240 720 6242
rect 774 6240 791 6242
rect 849 6240 862 6242
rect 924 6240 933 6242
rect 999 6240 1069 6272
rect 543 6208 579 6240
rect 613 6208 649 6240
rect 683 6208 720 6240
rect 754 6208 791 6240
rect 825 6208 862 6240
rect 896 6208 933 6240
rect 967 6208 1001 6240
rect 55 6203 123 6208
rect 19 6200 123 6203
rect -13 6198 123 6200
rect -13 6168 57 6198
rect 91 6168 123 6198
rect -47 6164 57 6168
rect -47 6161 21 6164
rect -47 6132 -15 6161
rect 19 6130 21 6161
rect 55 6134 89 6164
rect 55 6130 123 6134
rect 19 6127 123 6130
rect -13 6122 123 6127
rect -13 6098 57 6122
rect -47 6091 57 6098
rect 91 6094 123 6122
rect 933 6206 1001 6208
rect 1035 6238 1069 6240
rect 1035 6233 1103 6238
rect 1035 6206 1037 6233
rect 933 6199 1037 6206
rect 1071 6202 1103 6233
rect 933 6198 1069 6199
rect 933 6172 965 6198
rect 999 6170 1069 6198
rect 999 6164 1001 6170
rect 967 6138 1001 6164
rect 933 6136 1001 6138
rect 1035 6168 1069 6170
rect 1035 6158 1103 6168
rect 1035 6136 1037 6158
rect 933 6124 1037 6136
rect 1071 6132 1103 6158
rect 933 6122 1069 6124
rect -47 6088 21 6091
rect -47 6062 -15 6088
rect 19 6057 21 6088
rect 55 6088 57 6091
rect 55 6060 89 6088
rect 390 6080 428 6114
rect 462 6080 500 6114
rect 534 6080 572 6114
rect 606 6080 644 6114
rect 678 6080 716 6114
rect 933 6102 965 6122
rect 999 6100 1069 6122
rect 999 6088 1001 6100
rect 55 6057 123 6060
rect 19 6054 123 6057
rect -13 6046 123 6054
rect -13 6028 57 6046
rect -47 6018 57 6028
rect 91 6020 123 6046
rect -47 6015 21 6018
rect -47 5992 -15 6015
rect 19 5984 21 6015
rect 55 6012 57 6018
rect 55 5986 89 6012
rect 55 5984 123 5986
rect 19 5981 123 5984
rect -13 5970 123 5981
rect -13 5958 57 5970
rect -47 5945 57 5958
rect 91 5946 123 5970
rect -47 5942 21 5945
rect -47 5922 -15 5942
rect 19 5911 21 5942
rect 55 5936 57 5945
rect 55 5912 89 5936
rect 55 5911 123 5912
rect 19 5908 123 5911
rect -13 5894 123 5908
rect -13 5888 57 5894
rect -47 5872 57 5888
rect 91 5873 123 5894
rect -47 5869 21 5872
rect -47 5852 -15 5869
rect 19 5838 21 5869
rect 55 5860 57 5872
rect 55 5839 89 5860
rect 55 5838 123 5839
rect 19 5835 123 5838
rect -13 5818 123 5835
rect -47 5799 57 5818
rect 91 5800 123 5818
rect -47 5795 21 5799
rect -47 5782 -15 5795
rect 19 5765 21 5795
rect 55 5784 57 5799
rect 55 5766 89 5784
rect 55 5765 123 5766
rect 19 5761 123 5765
rect -13 5748 123 5761
rect -47 5742 123 5748
rect -47 5726 57 5742
rect 91 5727 123 5742
rect -47 5721 21 5726
rect -47 5712 -15 5721
rect 19 5692 21 5721
rect 55 5708 57 5726
rect 55 5693 89 5708
rect 55 5692 123 5693
rect 19 5687 123 5692
rect -13 5678 123 5687
rect -47 5666 123 5678
rect -47 5653 57 5666
rect 91 5654 123 5666
rect -47 5647 21 5653
rect -47 5642 -15 5647
rect 19 5619 21 5647
rect 55 5632 57 5653
rect 55 5620 89 5632
rect 55 5619 123 5620
rect 19 5613 123 5619
rect -13 5608 123 5613
rect -47 5590 123 5608
rect -47 5580 57 5590
rect 91 5581 123 5590
rect -47 5573 21 5580
rect -47 5572 -15 5573
rect 19 5546 21 5573
rect 55 5556 57 5580
rect 55 5547 89 5556
rect 55 5546 123 5547
rect 19 5539 123 5546
rect -13 5538 123 5539
rect -47 5514 123 5538
rect -47 5507 57 5514
rect 91 5508 123 5514
rect -47 5502 21 5507
rect -13 5499 21 5502
rect 19 5473 21 5499
rect 55 5480 57 5507
rect 55 5474 89 5480
rect 55 5473 123 5474
rect -47 5465 -15 5468
rect 19 5465 123 5473
rect -47 5437 123 5465
rect -47 5434 57 5437
rect 91 5435 123 5437
rect -47 5432 21 5434
rect -13 5425 21 5432
rect 19 5400 21 5425
rect 55 5403 57 5434
rect 55 5401 89 5403
rect 55 5400 123 5401
rect -47 5391 -15 5398
rect 19 5391 123 5400
rect 171 6053 205 6069
rect 171 5985 205 6019
rect 967 6068 1001 6088
rect 933 6066 1001 6068
rect 1035 6098 1069 6100
rect 1035 6083 1103 6098
rect 1035 6066 1037 6083
rect 933 6049 1037 6066
rect 1071 6062 1103 6083
rect 933 6046 1069 6049
rect 933 6032 965 6046
rect 999 6030 1069 6046
rect 999 6012 1001 6030
rect 967 5998 1001 6012
rect 933 5996 1001 5998
rect 1035 6028 1069 6030
rect 1035 6008 1103 6028
rect 1035 5996 1037 6008
rect 933 5974 1037 5996
rect 1071 5992 1103 6008
rect 933 5970 1069 5974
rect 933 5962 965 5970
rect 171 5917 205 5951
rect 390 5924 428 5958
rect 462 5924 500 5958
rect 534 5924 572 5958
rect 606 5924 644 5958
rect 678 5924 716 5958
rect 999 5960 1069 5970
rect 999 5936 1001 5960
rect 967 5928 1001 5936
rect 933 5926 1001 5928
rect 1035 5958 1069 5960
rect 1035 5933 1103 5958
rect 1035 5926 1037 5933
rect 171 5849 205 5883
rect 171 5781 205 5815
rect 933 5899 1037 5926
rect 1071 5922 1103 5933
rect 933 5895 1069 5899
rect 933 5891 965 5895
rect 999 5890 1069 5895
rect 999 5861 1001 5890
rect 967 5857 1001 5861
rect 933 5856 1001 5857
rect 1035 5888 1069 5890
rect 1035 5858 1103 5888
rect 1035 5856 1037 5858
rect 933 5824 1037 5856
rect 1071 5852 1103 5858
rect 933 5820 1069 5824
rect 546 5768 584 5802
rect 618 5768 656 5802
rect 690 5768 728 5802
rect 999 5786 1001 5820
rect 1035 5818 1069 5820
rect 1035 5786 1103 5818
rect 933 5783 1103 5786
rect 171 5713 205 5747
rect 933 5750 1037 5783
rect 1071 5782 1103 5783
rect 933 5749 1001 5750
rect 967 5745 1001 5749
rect 999 5716 1001 5745
rect 1035 5749 1037 5750
rect 1035 5748 1069 5749
rect 1035 5716 1103 5748
rect 933 5711 965 5715
rect 999 5712 1103 5716
rect 999 5711 1069 5712
rect 933 5708 1069 5711
rect 171 5645 205 5679
rect 550 5658 588 5692
rect 622 5658 660 5692
rect 694 5658 732 5692
rect 933 5680 1037 5708
rect 933 5678 1001 5680
rect 967 5670 1001 5678
rect 171 5577 205 5611
rect 171 5509 205 5543
rect 999 5646 1001 5670
rect 1035 5674 1037 5680
rect 1071 5674 1103 5678
rect 1035 5646 1103 5674
rect 933 5636 965 5644
rect 999 5642 1103 5646
rect 999 5636 1069 5642
rect 933 5633 1069 5636
rect 933 5610 1037 5633
rect 933 5607 1001 5610
rect 967 5595 1001 5607
rect 999 5576 1001 5595
rect 1035 5599 1037 5610
rect 1071 5599 1103 5608
rect 1035 5576 1103 5599
rect 933 5561 965 5573
rect 999 5572 1103 5576
rect 999 5561 1069 5572
rect 933 5558 1069 5561
rect 933 5539 1037 5558
rect 933 5536 1001 5539
rect 550 5502 588 5536
rect 622 5502 660 5536
rect 694 5502 732 5536
rect 967 5520 1001 5536
rect 999 5505 1001 5520
rect 1035 5524 1037 5539
rect 1071 5524 1103 5538
rect 1035 5505 1103 5524
rect 999 5502 1103 5505
rect 171 5441 205 5475
rect 171 5391 205 5407
rect 933 5486 965 5502
rect 999 5486 1069 5502
rect 933 5484 1069 5486
rect 933 5468 1037 5484
rect 933 5465 1001 5468
rect 967 5445 1001 5465
rect 999 5434 1001 5445
rect 1035 5450 1037 5468
rect 1071 5450 1103 5468
rect 1035 5434 1103 5450
rect 999 5432 1103 5434
rect 933 5411 965 5431
rect 999 5411 1069 5432
rect 933 5410 1069 5411
rect 933 5397 1037 5410
rect 933 5394 1001 5397
rect -47 5362 123 5391
rect -13 5351 21 5362
rect 19 5328 21 5351
rect 55 5360 89 5362
rect 55 5328 57 5360
rect 630 5346 668 5380
rect 702 5346 740 5380
rect 967 5370 1001 5394
rect 999 5363 1001 5370
rect 1035 5376 1037 5397
rect 1071 5376 1103 5398
rect 1035 5363 1103 5376
rect 999 5362 1103 5363
rect -47 5317 -15 5328
rect 19 5326 57 5328
rect 91 5326 123 5328
rect 19 5317 123 5326
rect -47 5283 123 5317
rect -47 5277 57 5283
rect -47 5252 -15 5277
rect 19 5252 57 5277
rect 91 5252 123 5283
rect 933 5336 965 5360
rect 999 5336 1069 5362
rect 933 5326 1037 5336
rect 933 5323 1001 5326
rect 967 5295 1001 5323
rect 999 5292 1001 5295
rect 1035 5302 1037 5326
rect 1071 5302 1103 5328
rect 1035 5292 1103 5302
rect 933 5261 965 5289
rect 999 5262 1069 5292
rect 999 5261 1037 5262
rect 933 5255 1037 5261
rect 933 5252 1001 5255
rect -47 5218 -23 5252
rect 19 5243 46 5252
rect 91 5249 115 5252
rect 11 5218 46 5243
rect 80 5218 115 5249
rect 149 5218 184 5252
rect 218 5218 253 5252
rect 967 5221 1001 5252
rect 1035 5228 1037 5255
rect 1071 5228 1103 5258
rect 1035 5221 1103 5228
rect 967 5220 1069 5221
rect -47 5206 253 5218
rect -47 5203 57 5206
rect -47 5184 -15 5203
rect 19 5184 57 5203
rect 91 5184 253 5206
rect 999 5187 1069 5220
rect 999 5186 1103 5187
rect -47 5150 -23 5184
rect 19 5169 46 5184
rect 91 5172 115 5184
rect 11 5150 46 5169
rect 80 5150 115 5172
rect 149 5150 184 5184
rect 218 5150 253 5184
rect 967 5184 1103 5186
rect 967 5150 1001 5184
rect 1035 5150 1103 5184
rect -47 5148 1069 5150
rect -47 5129 715 5148
rect -47 5116 -15 5129
rect 19 5116 57 5129
rect 91 5116 715 5129
rect 749 5116 809 5148
rect 843 5116 904 5148
rect 938 5116 999 5148
rect -47 5082 -23 5116
rect 19 5095 48 5116
rect 91 5095 119 5116
rect 11 5082 48 5095
rect 82 5082 119 5095
rect 153 5082 190 5116
rect 224 5082 261 5116
rect 295 5082 332 5116
rect 366 5082 403 5116
rect 437 5082 473 5116
rect 507 5082 543 5116
rect 577 5082 613 5116
rect 647 5082 683 5116
rect 749 5114 753 5116
rect 717 5082 753 5114
rect 787 5114 809 5116
rect 787 5082 823 5114
rect 857 5082 893 5116
rect 938 5114 963 5116
rect 927 5082 963 5114
rect 997 5114 999 5116
rect 1033 5116 1069 5148
rect 1033 5114 1103 5116
rect 997 5082 1103 5114
rect 1255 6412 1287 6448
rect 1393 6452 1425 6488
rect 26149 6627 26217 6628
rect 26251 6653 26253 6661
rect 26287 6653 26319 6661
rect 26251 6627 26319 6653
rect 26149 6626 26319 6627
rect 26149 6614 26285 6626
rect 26149 6593 26181 6614
rect 26215 6592 26253 6614
rect 26215 6580 26217 6592
rect 26183 6559 26217 6580
rect 26149 6558 26217 6559
rect 26251 6580 26253 6592
rect 26287 6580 26319 6592
rect 26251 6558 26319 6580
rect 26149 6541 26285 6558
rect 26149 6524 26181 6541
rect 26215 6523 26253 6541
rect 26215 6507 26217 6523
rect 26183 6490 26217 6507
rect 26149 6489 26217 6490
rect 26251 6507 26253 6523
rect 26287 6507 26319 6524
rect 26251 6490 26319 6507
rect 26251 6489 26285 6490
rect 1255 6342 1287 6378
rect 1393 6382 1425 6418
rect 1255 6272 1287 6308
rect 1393 6312 1425 6348
rect 1255 6202 1287 6238
rect 1393 6242 1425 6278
rect 1255 6132 1287 6168
rect 1393 6172 1425 6208
rect 1255 6062 1287 6098
rect 1393 6102 1425 6138
rect 1255 5992 1287 6028
rect 1393 6032 1425 6068
rect 1255 5922 1287 5958
rect 1393 5962 1425 5998
rect 1255 5852 1287 5888
rect 1393 5892 1425 5928
rect 1255 5782 1287 5818
rect 1393 5822 1425 5858
rect 1255 5711 1287 5748
rect 1393 5751 1425 5788
rect 1255 5640 1287 5677
rect 1393 5680 1425 5717
rect 1255 5569 1287 5606
rect 1393 5609 1425 5646
rect 1255 5498 1287 5535
rect 1393 5538 1425 5575
rect 1255 5427 1287 5464
rect 1393 5467 1425 5504
rect 1255 5356 1287 5393
rect 1393 5396 1425 5433
rect 1255 5285 1287 5322
rect 1393 5325 1425 5362
rect 1255 5214 1287 5251
rect 1393 5254 1425 5291
rect 1255 5148 1287 5180
rect 1393 5183 1425 5220
rect 1393 5148 1425 5149
rect 1255 5143 1425 5148
rect 1289 5142 1425 5143
rect 1289 5109 1323 5142
rect -335 4998 -303 5034
rect -335 4828 -303 4964
rect 1255 5075 1287 5109
rect 1321 5108 1323 5109
rect 1357 5112 1425 5142
rect 1357 5109 1391 5112
rect 1357 5108 1359 5109
rect 1321 5075 1359 5108
rect 1393 5075 1425 5078
rect 1255 5072 1425 5075
rect 1289 5038 1323 5072
rect 1357 5041 1425 5072
rect 1357 5038 1391 5041
rect 1255 5036 1391 5038
rect 1255 5002 1287 5036
rect 1321 5002 1359 5036
rect 1393 5002 1425 5007
rect 1255 5001 1323 5002
rect 1289 4968 1323 5001
rect 1357 4970 1425 5002
rect 1357 4968 1391 4970
rect 1289 4967 1391 4968
rect 1255 4963 1391 4967
rect 1255 4930 1287 4963
rect 1321 4932 1359 4963
rect -197 4896 -165 4930
rect -131 4896 -97 4930
rect -63 4896 -29 4930
rect 5 4896 39 4930
rect 73 4896 107 4930
rect 141 4896 175 4930
rect 209 4896 243 4930
rect 277 4896 311 4930
rect 345 4896 379 4930
rect 413 4896 447 4930
rect 481 4896 515 4930
rect 549 4896 583 4930
rect 617 4896 651 4930
rect 685 4896 719 4930
rect 753 4896 787 4930
rect 821 4896 855 4930
rect 889 4896 923 4930
rect 957 4896 991 4930
rect 1025 4896 1059 4930
rect 1093 4896 1164 4930
rect 1198 4896 1255 4930
rect 1321 4929 1323 4932
rect 1289 4898 1323 4929
rect 1357 4929 1359 4932
rect 1393 4929 1425 4936
rect 1357 4899 1425 4929
rect 1357 4898 1391 4899
rect 1289 4896 1391 4898
rect -197 4890 1391 4896
rect -197 4862 1287 4890
rect -163 4828 -127 4862
rect -93 4828 -57 4862
rect -23 4828 13 4862
rect 47 4828 83 4862
rect 117 4828 153 4862
rect 187 4828 223 4862
rect 257 4828 293 4862
rect 327 4828 363 4862
rect 397 4828 433 4862
rect 467 4828 503 4862
rect 537 4828 573 4862
rect 607 4828 643 4862
rect 677 4828 713 4862
rect 747 4828 783 4862
rect 817 4828 852 4862
rect 886 4828 921 4862
rect 955 4828 990 4862
rect 1024 4828 1059 4862
rect 1093 4828 1141 4862
rect 1175 4828 1232 4862
rect 1266 4856 1287 4862
rect 1321 4862 1359 4890
rect 1321 4856 1323 4862
rect 1266 4828 1323 4856
rect 1357 4856 1359 4862
rect 1393 4856 1425 4865
rect 1357 4828 1425 4856
rect -197 4794 1391 4828
rect -165 4760 -129 4794
rect -95 4760 -59 4794
rect -25 4760 11 4794
rect 45 4760 81 4794
rect 115 4760 151 4794
rect 185 4760 221 4794
rect 255 4760 291 4794
rect 325 4760 361 4794
rect 395 4760 431 4794
rect 465 4760 501 4794
rect 535 4760 571 4794
rect 605 4760 641 4794
rect 675 4760 711 4794
rect 745 4760 781 4794
rect 815 4760 851 4794
rect 885 4760 921 4794
rect 955 4760 990 4794
rect 1024 4760 1059 4794
rect 1093 4760 1141 4794
rect 1175 4760 1212 4794
rect 1246 4760 1283 4794
rect 1317 4760 1425 4794
rect 1577 6460 1804 6468
rect 23006 6460 23045 6473
rect 23079 6460 23118 6473
rect 23152 6460 23191 6473
rect 23225 6460 23264 6473
rect 23298 6460 23337 6473
rect 23371 6460 23410 6473
rect 23444 6460 23483 6473
rect 23517 6460 23556 6473
rect 23590 6460 23629 6473
rect 23663 6460 23702 6473
rect 23736 6460 23775 6473
rect 23809 6460 23848 6473
rect 23882 6460 23921 6473
rect 23955 6460 23994 6473
rect 24028 6460 24067 6473
rect 24101 6460 24140 6473
rect 24174 6460 24213 6473
rect 24247 6460 24286 6473
rect 24320 6460 24359 6473
rect 24393 6460 24432 6473
rect 24466 6460 24505 6473
rect 24539 6460 24578 6473
rect 24612 6460 24651 6473
rect 24685 6460 24724 6473
rect 24758 6460 24797 6473
rect 24831 6460 24870 6473
rect 24904 6460 24943 6473
rect 24977 6460 25016 6473
rect 25050 6460 25089 6473
rect 25123 6460 25162 6473
rect 25196 6460 25235 6473
rect 1577 6426 1601 6460
rect 1635 6426 1670 6460
rect 1704 6426 1739 6460
rect 1773 6426 1804 6460
rect 1577 6392 1804 6426
rect 1577 6358 1601 6392
rect 1635 6358 1670 6392
rect 1704 6358 1739 6392
rect 1773 6367 1804 6392
rect 25210 6439 25235 6460
rect 25269 6444 25308 6473
rect 25342 6444 25381 6473
rect 25415 6444 25454 6473
rect 25488 6444 25527 6473
rect 25561 6444 25938 6473
rect 25210 6401 25268 6439
rect 25210 6367 25235 6401
rect 1773 6358 1808 6367
rect 1842 6358 1877 6367
rect 1911 6358 1946 6367
rect 1980 6358 2015 6367
rect 2049 6358 2084 6367
rect 2118 6358 2153 6367
rect 2187 6358 2222 6367
rect 2256 6358 2291 6367
rect 2325 6358 2360 6367
rect 2394 6358 2429 6367
rect 2463 6358 2498 6367
rect 2532 6358 2567 6367
rect 2601 6358 2636 6367
rect 2670 6358 2705 6367
rect 2739 6358 2774 6367
rect 2808 6358 2843 6367
rect 2877 6358 2912 6367
rect 2946 6358 2981 6367
rect 3015 6358 3050 6367
rect 3084 6358 3119 6367
rect 3153 6358 3188 6367
rect 3222 6358 3257 6367
rect 3291 6358 3326 6367
rect 3360 6358 3395 6367
rect 3429 6358 3464 6367
rect 3498 6358 3533 6367
rect 3567 6358 3602 6367
rect 3636 6358 3671 6367
rect 3705 6358 3740 6367
rect 3774 6358 3809 6367
rect 3843 6358 3878 6367
rect 3912 6358 3947 6367
rect 3981 6358 4016 6367
rect 4050 6358 4085 6367
rect 4119 6358 4154 6367
rect 4188 6358 4223 6367
rect 4257 6358 4292 6367
rect 4326 6358 4361 6367
rect 4395 6358 4430 6367
rect 4464 6358 4499 6367
rect 4533 6358 4568 6367
rect 4602 6358 4637 6367
rect 4671 6358 4706 6367
rect 4740 6358 4775 6367
rect 4809 6358 4844 6367
rect 1577 6324 4844 6358
rect 1577 6290 1601 6324
rect 1635 6294 1670 6324
rect 1704 6294 1739 6324
rect 1643 6290 1670 6294
rect 1715 6290 1739 6294
rect 1773 6290 1808 6324
rect 1842 6290 1877 6324
rect 1911 6290 1946 6324
rect 1980 6290 2015 6324
rect 2049 6290 2084 6324
rect 2118 6290 2153 6324
rect 2187 6290 2222 6324
rect 2256 6290 2291 6324
rect 2325 6290 2360 6324
rect 2394 6290 2429 6324
rect 2463 6290 2498 6324
rect 2532 6290 2567 6324
rect 2601 6290 2636 6324
rect 2670 6290 2705 6324
rect 2739 6290 2774 6324
rect 2808 6290 2843 6324
rect 2877 6290 2912 6324
rect 2946 6290 2981 6324
rect 3015 6290 3050 6324
rect 3084 6290 3119 6324
rect 3153 6290 3188 6324
rect 3222 6290 3257 6324
rect 3291 6290 3326 6324
rect 3360 6290 3395 6324
rect 3429 6290 3464 6324
rect 3498 6290 3533 6324
rect 3567 6290 3602 6324
rect 3636 6290 3671 6324
rect 3705 6290 3740 6324
rect 3774 6290 3809 6324
rect 3843 6290 3878 6324
rect 3912 6290 3947 6324
rect 3981 6290 4016 6324
rect 4050 6290 4085 6324
rect 4119 6290 4154 6324
rect 4188 6290 4223 6324
rect 4257 6290 4292 6324
rect 4326 6290 4361 6324
rect 4395 6290 4430 6324
rect 4464 6290 4499 6324
rect 4533 6290 4568 6324
rect 4602 6290 4637 6324
rect 4671 6290 4706 6324
rect 4740 6290 4775 6324
rect 4809 6290 4844 6324
rect 1577 6260 1609 6290
rect 1643 6260 1681 6290
rect 1715 6260 4844 6290
rect 1577 6256 4844 6260
rect 1577 6222 1601 6256
rect 1635 6222 1670 6256
rect 1704 6222 1739 6256
rect 1773 6222 1808 6256
rect 1842 6222 1877 6256
rect 1911 6222 1946 6256
rect 1980 6222 2015 6256
rect 2049 6222 2084 6256
rect 2118 6222 2153 6256
rect 2187 6222 2222 6256
rect 2256 6222 2291 6256
rect 2325 6222 2360 6256
rect 2394 6222 2429 6256
rect 2463 6222 2498 6256
rect 2532 6222 2567 6256
rect 2601 6222 2636 6256
rect 2670 6222 2705 6256
rect 2739 6222 2774 6256
rect 2808 6222 2843 6256
rect 2877 6222 2912 6256
rect 2946 6222 2981 6256
rect 3015 6222 3050 6256
rect 3084 6222 3119 6256
rect 3153 6222 3188 6256
rect 3222 6222 3257 6256
rect 3291 6222 3326 6256
rect 3360 6222 3395 6256
rect 3429 6222 3464 6256
rect 3498 6222 3533 6256
rect 3567 6222 3602 6256
rect 3636 6222 3671 6256
rect 3705 6222 3740 6256
rect 3774 6222 3809 6256
rect 3843 6222 3878 6256
rect 3912 6222 3947 6256
rect 3981 6222 4016 6256
rect 4050 6222 4085 6256
rect 4119 6222 4154 6256
rect 4188 6222 4223 6256
rect 4257 6222 4292 6256
rect 4326 6222 4361 6256
rect 4395 6222 4430 6256
rect 4464 6222 4499 6256
rect 4533 6222 4568 6256
rect 4602 6222 4637 6256
rect 4671 6222 4706 6256
rect 4740 6222 4775 6256
rect 4809 6222 4844 6256
rect 1577 6220 1681 6222
rect 1577 6188 1609 6220
rect 1643 6188 1681 6220
rect 1715 6188 4844 6222
rect 1577 6154 1601 6188
rect 1643 6186 1670 6188
rect 1635 6154 1670 6186
rect 1704 6154 1739 6188
rect 1773 6154 1808 6188
rect 1842 6154 1877 6188
rect 1911 6154 1946 6188
rect 1980 6154 2015 6188
rect 2049 6154 2084 6188
rect 2118 6154 2153 6188
rect 2187 6154 2222 6188
rect 2256 6154 2291 6188
rect 2325 6154 2360 6188
rect 2394 6154 2429 6188
rect 2463 6154 2498 6188
rect 2532 6154 2567 6188
rect 2601 6154 2636 6188
rect 2670 6154 2705 6188
rect 2739 6154 2774 6188
rect 2808 6154 2843 6188
rect 2877 6154 2912 6188
rect 2946 6154 2981 6188
rect 3015 6154 3050 6188
rect 3084 6154 3119 6188
rect 3153 6154 3188 6188
rect 3222 6154 3257 6188
rect 3291 6154 3326 6188
rect 3360 6154 3395 6188
rect 3429 6154 3464 6188
rect 3498 6154 3533 6188
rect 3567 6154 3602 6188
rect 3636 6154 3671 6188
rect 3705 6154 3740 6188
rect 3774 6154 3809 6188
rect 3843 6154 3878 6188
rect 3912 6154 3947 6188
rect 3981 6154 4016 6188
rect 4050 6154 4085 6188
rect 4119 6154 4154 6188
rect 4188 6154 4223 6188
rect 4257 6154 4292 6188
rect 4326 6154 4361 6188
rect 4395 6154 4430 6188
rect 4464 6154 4499 6188
rect 4533 6154 4568 6188
rect 4602 6154 4637 6188
rect 4671 6154 4706 6188
rect 4740 6154 4775 6188
rect 4809 6154 4844 6188
rect 1577 6149 4844 6154
rect 1577 6146 1681 6149
rect 1577 6120 1609 6146
rect 1643 6120 1681 6146
rect 1715 6120 4844 6149
rect 1577 6086 1601 6120
rect 1643 6112 1670 6120
rect 1715 6115 1739 6120
rect 1635 6086 1670 6112
rect 1704 6086 1739 6115
rect 1773 6086 1808 6120
rect 1842 6086 1877 6120
rect 1911 6086 1946 6120
rect 1980 6086 2015 6120
rect 2049 6086 2084 6120
rect 2118 6086 2153 6120
rect 2187 6086 2222 6120
rect 2256 6086 2291 6120
rect 2325 6086 2360 6120
rect 2394 6086 2429 6120
rect 2463 6086 2498 6120
rect 2532 6086 2567 6120
rect 2601 6086 2636 6120
rect 2670 6086 2705 6120
rect 2739 6086 2774 6120
rect 2808 6086 2843 6120
rect 2877 6086 2912 6120
rect 2946 6086 2981 6120
rect 3015 6086 3050 6120
rect 3084 6086 3119 6120
rect 3153 6086 3188 6120
rect 3222 6086 3257 6120
rect 3291 6086 3326 6120
rect 3360 6086 3395 6120
rect 3429 6086 3464 6120
rect 3498 6086 3533 6120
rect 3567 6086 3602 6120
rect 3636 6086 3671 6120
rect 3705 6086 3740 6120
rect 3774 6086 3809 6120
rect 3843 6086 3878 6120
rect 3912 6086 3947 6120
rect 3981 6086 4016 6120
rect 4050 6086 4085 6120
rect 4119 6086 4154 6120
rect 4188 6086 4223 6120
rect 4257 6086 4292 6120
rect 4326 6086 4361 6120
rect 4395 6086 4430 6120
rect 4464 6086 4499 6120
rect 4533 6086 4568 6120
rect 4602 6086 4637 6120
rect 4671 6086 4706 6120
rect 4740 6086 4775 6120
rect 4809 6086 4844 6120
rect 1577 6076 4844 6086
rect 1577 6072 1681 6076
rect 1577 6052 1609 6072
rect 1643 6052 1681 6072
rect 1715 6052 4844 6076
rect 1577 6018 1601 6052
rect 1643 6038 1670 6052
rect 1715 6042 1739 6052
rect 1635 6018 1670 6038
rect 1704 6018 1739 6042
rect 1773 6018 1808 6052
rect 1842 6018 1877 6052
rect 1911 6018 1946 6052
rect 1980 6018 2015 6052
rect 2049 6018 2084 6052
rect 2118 6018 2153 6052
rect 2187 6018 2222 6052
rect 2256 6018 2291 6052
rect 2325 6018 2360 6052
rect 2394 6018 2429 6052
rect 2463 6018 2498 6052
rect 2532 6018 2567 6052
rect 2601 6018 2636 6052
rect 2670 6018 2705 6052
rect 2739 6018 2774 6052
rect 2808 6018 2843 6052
rect 2877 6018 2912 6052
rect 2946 6018 2981 6052
rect 3015 6018 3050 6052
rect 3084 6018 3119 6052
rect 3153 6018 3188 6052
rect 3222 6018 3257 6052
rect 3291 6018 3326 6052
rect 3360 6018 3395 6052
rect 3429 6018 3464 6052
rect 3498 6018 3533 6052
rect 3567 6018 3602 6052
rect 3636 6018 3671 6052
rect 3705 6018 3740 6052
rect 3774 6018 3809 6052
rect 3843 6018 3878 6052
rect 3912 6018 3947 6052
rect 3981 6018 4016 6052
rect 4050 6018 4085 6052
rect 4119 6018 4154 6052
rect 4188 6018 4223 6052
rect 4257 6018 4292 6052
rect 4326 6018 4361 6052
rect 4395 6018 4430 6052
rect 4464 6018 4499 6052
rect 4533 6018 4568 6052
rect 4602 6018 4637 6052
rect 4671 6018 4706 6052
rect 4740 6018 4775 6052
rect 4809 6018 4844 6052
rect 1577 6003 4844 6018
rect 1577 5998 1681 6003
rect 1577 5984 1609 5998
rect 1643 5984 1681 5998
rect 1715 5984 4844 6003
rect 1577 5950 1601 5984
rect 1643 5964 1670 5984
rect 1715 5969 1739 5984
rect 1635 5950 1670 5964
rect 1704 5950 1739 5969
rect 1773 5950 1808 5984
rect 1842 5950 1877 5984
rect 1911 5950 1946 5984
rect 1980 5950 2015 5984
rect 2049 5950 2084 5984
rect 2118 5950 2153 5984
rect 2187 5950 2222 5984
rect 2256 5950 2291 5984
rect 2325 5950 2360 5984
rect 2394 5950 2429 5984
rect 2463 5950 2498 5984
rect 2532 5950 2567 5984
rect 2601 5950 2636 5984
rect 2670 5950 2705 5984
rect 2739 5950 2774 5984
rect 2808 5950 2843 5984
rect 2877 5950 2912 5984
rect 2946 5950 2981 5984
rect 3015 5950 3050 5984
rect 3084 5950 3119 5984
rect 3153 5950 3188 5984
rect 3222 5950 3257 5984
rect 3291 5950 3326 5984
rect 3360 5950 3395 5984
rect 3429 5950 3464 5984
rect 3498 5950 3533 5984
rect 3567 5950 3602 5984
rect 3636 5950 3671 5984
rect 3705 5950 3740 5984
rect 3774 5950 3809 5984
rect 3843 5950 3878 5984
rect 3912 5950 3947 5984
rect 3981 5950 4016 5984
rect 4050 5950 4085 5984
rect 4119 5950 4154 5984
rect 4188 5950 4223 5984
rect 4257 5950 4292 5984
rect 4326 5950 4361 5984
rect 4395 5950 4430 5984
rect 4464 5950 4499 5984
rect 4533 5950 4568 5984
rect 4602 5950 4637 5984
rect 4671 5950 4706 5984
rect 4740 5950 4775 5984
rect 4809 5950 4844 5984
rect 1577 5930 4844 5950
rect 1577 5924 1681 5930
rect 1577 5916 1609 5924
rect 1643 5916 1681 5924
rect 1715 5916 4844 5930
rect 1577 5882 1601 5916
rect 1643 5890 1670 5916
rect 1715 5896 1739 5916
rect 1635 5882 1670 5890
rect 1704 5882 1739 5896
rect 1773 5882 1808 5916
rect 1842 5882 1877 5916
rect 1911 5882 1946 5916
rect 1980 5882 2015 5916
rect 2049 5882 2084 5916
rect 2118 5882 2153 5916
rect 2187 5882 2222 5916
rect 2256 5882 2291 5916
rect 2325 5882 2360 5916
rect 2394 5882 2429 5916
rect 2463 5882 2498 5916
rect 2532 5882 2567 5916
rect 2601 5882 2636 5916
rect 2670 5882 2705 5916
rect 2739 5882 2774 5916
rect 2808 5882 2843 5916
rect 2877 5882 2912 5916
rect 2946 5882 2981 5916
rect 3015 5882 3050 5916
rect 3084 5882 3119 5916
rect 3153 5882 3188 5916
rect 3222 5882 3257 5916
rect 3291 5882 3326 5916
rect 3360 5882 3395 5916
rect 3429 5882 3464 5916
rect 3498 5882 3533 5916
rect 3567 5882 3602 5916
rect 3636 5882 3671 5916
rect 3705 5882 3740 5916
rect 3774 5882 3809 5916
rect 3843 5882 3878 5916
rect 3912 5882 3947 5916
rect 3981 5882 4016 5916
rect 4050 5882 4085 5916
rect 4119 5882 4154 5916
rect 4188 5882 4223 5916
rect 4257 5882 4292 5916
rect 4326 5882 4361 5916
rect 4395 5882 4430 5916
rect 4464 5882 4499 5916
rect 4533 5882 4568 5916
rect 4602 5882 4637 5916
rect 4671 5882 4706 5916
rect 4740 5882 4775 5916
rect 4809 5882 4844 5916
rect 1577 5857 4844 5882
rect 1577 5850 1681 5857
rect 1577 5848 1609 5850
rect 1643 5848 1681 5850
rect 1715 5848 4844 5857
rect 1577 5814 1601 5848
rect 1643 5816 1670 5848
rect 1715 5823 1739 5848
rect 1635 5814 1670 5816
rect 1704 5814 1739 5823
rect 1773 5814 1808 5848
rect 1842 5814 1877 5848
rect 1911 5814 1946 5848
rect 1980 5814 2015 5848
rect 2049 5814 2084 5848
rect 2118 5814 2153 5848
rect 2187 5814 2222 5848
rect 2256 5814 2291 5848
rect 2325 5814 2360 5848
rect 2394 5814 2429 5848
rect 2463 5814 2498 5848
rect 2532 5814 2567 5848
rect 2601 5814 2636 5848
rect 2670 5814 2705 5848
rect 2739 5814 2774 5848
rect 2808 5814 2843 5848
rect 2877 5814 2912 5848
rect 2946 5814 2981 5848
rect 3015 5814 3050 5848
rect 3084 5814 3119 5848
rect 3153 5814 3188 5848
rect 3222 5814 3257 5848
rect 3291 5814 3326 5848
rect 3360 5814 3395 5848
rect 3429 5814 3464 5848
rect 3498 5814 3533 5848
rect 3567 5814 3602 5848
rect 3636 5814 3671 5848
rect 3705 5814 3740 5848
rect 3774 5814 3809 5848
rect 3843 5814 3878 5848
rect 3912 5814 3947 5848
rect 3981 5814 4016 5848
rect 4050 5814 4085 5848
rect 4119 5814 4154 5848
rect 4188 5814 4223 5848
rect 4257 5814 4292 5848
rect 4326 5814 4361 5848
rect 4395 5814 4430 5848
rect 4464 5814 4499 5848
rect 4533 5814 4568 5848
rect 4602 5814 4637 5848
rect 4671 5814 4706 5848
rect 4740 5814 4775 5848
rect 4809 5814 4844 5848
rect 1577 5784 4844 5814
rect 1577 5780 1681 5784
rect 1715 5780 4844 5784
rect 1577 5746 1601 5780
rect 1635 5776 1670 5780
rect 1643 5746 1670 5776
rect 1715 5750 1739 5780
rect 1704 5746 1739 5750
rect 1773 5746 1808 5780
rect 1842 5746 1877 5780
rect 1911 5746 1946 5780
rect 1980 5746 2015 5780
rect 2049 5746 2084 5780
rect 2118 5746 2153 5780
rect 2187 5746 2222 5780
rect 2256 5746 2291 5780
rect 2325 5746 2360 5780
rect 2394 5746 2429 5780
rect 2463 5746 2498 5780
rect 2532 5746 2567 5780
rect 2601 5746 2636 5780
rect 2670 5746 2705 5780
rect 2739 5746 2774 5780
rect 2808 5746 2843 5780
rect 2877 5746 2912 5780
rect 2946 5746 2981 5780
rect 3015 5746 3050 5780
rect 3084 5746 3119 5780
rect 3153 5746 3188 5780
rect 3222 5746 3257 5780
rect 3291 5746 3326 5780
rect 3360 5746 3395 5780
rect 3429 5746 3464 5780
rect 3498 5746 3533 5780
rect 3567 5746 3602 5780
rect 3636 5746 3671 5780
rect 3705 5746 3740 5780
rect 3774 5746 3809 5780
rect 3843 5746 3878 5780
rect 3912 5746 3947 5780
rect 3981 5746 4016 5780
rect 4050 5746 4085 5780
rect 4119 5746 4154 5780
rect 4188 5746 4223 5780
rect 4257 5746 4292 5780
rect 4326 5746 4361 5780
rect 4395 5746 4430 5780
rect 4464 5746 4499 5780
rect 4533 5746 4568 5780
rect 4602 5746 4637 5780
rect 4671 5746 4706 5780
rect 4740 5746 4775 5780
rect 4809 5746 4844 5780
rect 25210 5746 25268 6367
rect 1577 5742 1609 5746
rect 1643 5742 4844 5746
rect 1577 5712 4844 5742
rect 6421 5712 25268 5746
rect 1577 5702 1611 5712
rect 1577 5668 1609 5702
rect 1645 5678 1681 5712
rect 1715 5678 1751 5712
rect 1785 5678 1821 5712
rect 1855 5678 1891 5712
rect 1925 5678 1961 5712
rect 1995 5678 2030 5712
rect 2064 5678 2099 5712
rect 2133 5678 2168 5712
rect 2202 5678 2237 5712
rect 2271 5678 2306 5712
rect 2340 5678 2375 5712
rect 1643 5677 1681 5678
rect 1715 5677 2375 5678
rect 1643 5668 2375 5677
rect 1577 5644 2375 5668
rect 6421 5654 6455 5712
rect 1577 5627 1645 5644
rect 1577 5604 1609 5627
rect 1643 5610 1645 5627
rect 1679 5638 1718 5644
rect 1679 5610 1681 5638
rect 1643 5604 1681 5610
rect 1715 5610 1718 5638
rect 1752 5610 1791 5644
rect 1825 5610 1864 5644
rect 1898 5610 1937 5644
rect 1971 5610 2010 5644
rect 2044 5610 2083 5644
rect 2117 5610 2156 5644
rect 2190 5610 2229 5644
rect 2263 5610 2302 5644
rect 2336 5610 2375 5644
rect 1715 5604 2375 5610
rect 1643 5593 2375 5604
rect 1611 5576 2375 5593
rect 1611 5575 1713 5576
rect 1611 5570 1645 5575
rect 1577 5552 1645 5570
rect 1577 5533 1609 5552
rect 1643 5541 1645 5552
rect 1679 5565 1713 5575
rect 1679 5541 1681 5565
rect 1747 5542 1787 5576
rect 1821 5542 1861 5576
rect 1895 5542 1935 5576
rect 1969 5542 2009 5576
rect 2043 5542 2083 5576
rect 2117 5542 2156 5576
rect 2190 5542 2229 5576
rect 2263 5542 2302 5576
rect 2336 5542 2375 5576
rect 6421 5542 6455 5548
rect 1643 5531 1681 5541
rect 1715 5531 4023 5542
rect 1643 5518 4023 5531
rect 1611 5506 4023 5518
rect 1611 5499 1645 5506
rect 1577 5477 1645 5499
rect 1577 5462 1609 5477
rect 1643 5472 1645 5477
rect 1679 5505 4023 5506
rect 1679 5492 1713 5505
rect 1679 5472 1681 5492
rect 1643 5458 1681 5472
rect 1747 5471 1781 5505
rect 1815 5471 1850 5505
rect 1884 5471 1919 5505
rect 1953 5471 1988 5505
rect 2022 5471 2057 5505
rect 2091 5471 2126 5505
rect 2160 5471 2195 5505
rect 2229 5471 2264 5505
rect 2298 5471 2333 5505
rect 1715 5458 2333 5471
rect 1643 5443 2333 5458
rect 1611 5437 2333 5443
rect 1611 5428 1645 5437
rect 1577 5403 1645 5428
rect 1679 5434 1781 5437
rect 1679 5419 1713 5434
rect 1679 5403 1681 5419
rect 1577 5402 1681 5403
rect 1577 5391 1609 5402
rect 1643 5385 1681 5402
rect 1747 5403 1781 5434
rect 1815 5403 1850 5437
rect 1884 5403 1919 5437
rect 1953 5403 1988 5437
rect 2022 5403 2057 5437
rect 2091 5403 2126 5437
rect 2160 5403 2195 5437
rect 2229 5403 2264 5437
rect 2298 5403 2333 5437
rect 1747 5400 2333 5403
rect 1715 5385 2333 5400
rect 1643 5369 2333 5385
rect 1643 5368 1781 5369
rect 1611 5357 1645 5368
rect 1577 5334 1645 5357
rect 1679 5363 1781 5368
rect 1679 5346 1713 5363
rect 1679 5334 1681 5346
rect 1577 5327 1681 5334
rect 1747 5335 1781 5363
rect 1815 5335 1850 5369
rect 1884 5335 1919 5369
rect 1953 5335 1988 5369
rect 2022 5335 2057 5369
rect 2091 5335 2126 5369
rect 2160 5335 2195 5369
rect 2229 5335 2264 5369
rect 2298 5335 2333 5369
rect 1747 5329 2333 5335
rect 1577 5320 1609 5327
rect 1643 5312 1681 5327
rect 1715 5312 2333 5329
rect 1643 5301 2333 5312
rect 1643 5299 1781 5301
rect 1643 5293 1645 5299
rect 1611 5286 1645 5293
rect 1577 5265 1645 5286
rect 1679 5292 1781 5299
rect 1679 5273 1713 5292
rect 1679 5265 1681 5273
rect 1577 5252 1681 5265
rect 1747 5267 1781 5292
rect 1815 5267 1850 5301
rect 1884 5267 1919 5301
rect 1953 5267 1988 5301
rect 2022 5267 2057 5301
rect 2091 5267 2126 5301
rect 2160 5267 2195 5301
rect 2229 5267 2264 5301
rect 2298 5267 2333 5301
rect 1747 5258 2333 5267
rect 1577 5249 1609 5252
rect 1643 5239 1681 5252
rect 1715 5239 2333 5258
rect 1643 5233 2333 5239
rect 1643 5230 1781 5233
rect 1643 5218 1645 5230
rect 1611 5215 1645 5218
rect 1577 5196 1645 5215
rect 1679 5221 1781 5230
rect 1679 5200 1713 5221
rect 1679 5196 1681 5200
rect 1577 5178 1681 5196
rect 1747 5199 1781 5221
rect 1815 5199 1850 5233
rect 1884 5199 1919 5233
rect 1953 5199 1988 5233
rect 2022 5199 2057 5233
rect 2091 5199 2126 5233
rect 2160 5199 2195 5233
rect 2229 5199 2264 5233
rect 2298 5199 2333 5233
rect 1747 5187 2333 5199
rect 1611 5177 1681 5178
rect 1643 5166 1681 5177
rect 1715 5166 2333 5187
rect 1643 5165 2333 5166
rect 1643 5161 1781 5165
rect 1577 5143 1609 5144
rect 1643 5143 1645 5161
rect 1577 5127 1645 5143
rect 1679 5150 1781 5161
rect 1679 5127 1713 5150
rect 1747 5131 1781 5150
rect 1815 5131 1850 5165
rect 1884 5131 1919 5165
rect 1953 5131 1988 5165
rect 2022 5131 2057 5165
rect 2091 5131 2126 5165
rect 2160 5131 2195 5165
rect 2229 5131 2264 5165
rect 2298 5131 2333 5165
rect 1577 5107 1681 5127
rect 1747 5116 2333 5131
rect 1611 5102 1681 5107
rect 1643 5093 1681 5102
rect 1715 5097 2333 5116
rect 1715 5093 1781 5097
rect 1643 5092 1781 5093
rect 1577 5068 1609 5073
rect 1643 5068 1645 5092
rect 1577 5058 1645 5068
rect 1679 5079 1781 5092
rect 1679 5058 1713 5079
rect 1577 5054 1713 5058
rect 1747 5063 1781 5079
rect 1815 5063 1850 5097
rect 1884 5063 1919 5097
rect 1953 5063 1988 5097
rect 2022 5063 2057 5097
rect 2091 5063 2126 5097
rect 2160 5063 2195 5097
rect 2229 5063 2264 5097
rect 2298 5063 2333 5097
rect 1577 5036 1681 5054
rect 1747 5045 2333 5063
rect 1611 5027 1681 5036
rect 1643 5023 1681 5027
rect 1577 4993 1609 5002
rect 1643 4993 1645 5023
rect 1577 4989 1645 4993
rect 1679 5020 1681 5023
rect 1715 5029 2333 5045
rect 1715 5020 1781 5029
rect 1679 5008 1781 5020
rect 1679 4989 1713 5008
rect 1577 4981 1713 4989
rect 1747 4995 1781 5008
rect 1815 4995 1850 5029
rect 1884 4995 1919 5029
rect 1953 4995 1988 5029
rect 2022 4995 2057 5029
rect 2091 4995 2126 5029
rect 2160 4995 2195 5029
rect 2229 4995 2264 5029
rect 2298 4995 2333 5029
rect 3999 4995 4023 5505
rect 4107 5428 4726 5508
rect 4107 5394 4181 5428
rect 1747 4992 4023 4995
rect 1577 4965 1681 4981
rect 1611 4954 1681 4965
rect 1611 4952 1645 4954
rect 1577 4918 1609 4931
rect 1643 4920 1645 4952
rect 1679 4947 1681 4954
rect 1715 4947 1747 4974
rect 1679 4937 1747 4947
rect 1679 4920 1713 4937
rect 1643 4918 1713 4920
rect 1577 4908 1713 4918
rect 1577 4894 1681 4908
rect 1611 4885 1681 4894
rect 1611 4877 1645 4885
rect 1577 4843 1609 4860
rect 1643 4851 1645 4877
rect 1679 4874 1681 4885
rect 1715 4874 1747 4903
rect 4107 4956 4181 4990
rect 4291 4956 4726 5428
rect 4107 4899 4726 4956
rect 5902 5428 6373 5508
rect 5902 4956 6189 5428
rect 6299 5394 6373 5428
rect 6299 4956 6373 4990
rect 5902 4899 6373 4956
rect 1679 4866 1747 4874
rect 1679 4851 1713 4866
rect 1643 4843 1713 4851
rect 1577 4835 1713 4843
rect 1577 4823 1681 4835
rect 1611 4816 1681 4823
rect 1611 4802 1645 4816
rect 1577 4768 1609 4789
rect 1643 4782 1645 4802
rect 1679 4801 1681 4816
rect 1715 4801 1747 4832
rect 1679 4794 1747 4801
rect 1679 4782 1713 4794
rect 1643 4768 1713 4782
rect 1577 4762 1713 4768
rect 1577 4752 1681 4762
rect 1611 4747 1681 4752
rect 1611 4727 1645 4747
rect 1577 4693 1609 4718
rect 1643 4713 1645 4727
rect 1679 4728 1681 4747
rect 1715 4728 1747 4760
rect 1679 4722 1747 4728
rect 1679 4713 1713 4722
rect 1643 4693 1713 4713
rect 1577 4689 1713 4693
rect 1577 4680 1681 4689
rect 1611 4678 1681 4680
rect 1611 4652 1645 4678
rect 1577 4618 1609 4646
rect 1643 4644 1645 4652
rect 1679 4655 1681 4678
rect 1715 4655 1747 4688
rect 1679 4650 1747 4655
rect 1679 4644 1713 4650
rect 1643 4618 1713 4644
rect 1577 4616 1713 4618
rect 1577 4609 1681 4616
rect 1577 4608 1645 4609
rect -335 4216 -303 4250
rect -197 4249 -165 4284
rect -335 4148 -303 4182
rect -197 4180 -165 4215
rect -335 4102 -303 4114
rect -197 4111 -165 4146
rect -335 4080 -267 4102
rect -301 4077 -267 4080
rect -233 4077 -231 4102
rect -301 4068 -231 4077
rect -197 4068 -165 4077
rect -301 4063 -165 4068
rect -335 4029 -303 4046
rect -269 4042 -165 4063
rect -269 4029 -267 4042
rect -335 4012 -267 4029
rect -301 4008 -267 4012
rect -233 4030 -199 4042
rect -233 4008 -231 4030
rect -301 3996 -231 4008
rect -197 3996 -165 4008
rect -301 3990 -165 3996
rect -335 3956 -303 3978
rect -269 3973 -165 3990
rect -269 3956 -267 3973
rect -335 3944 -267 3956
rect -301 3939 -267 3944
rect -233 3958 -199 3973
rect -233 3939 -231 3958
rect -301 3924 -231 3939
rect -197 3924 -165 3939
rect -301 3917 -165 3924
rect -335 3883 -303 3910
rect -269 3904 -165 3917
rect -269 3883 -267 3904
rect -335 3876 -267 3883
rect -301 3870 -267 3876
rect -233 3886 -199 3904
rect -233 3870 -231 3886
rect -301 3852 -231 3870
rect -197 3852 -165 3870
rect -301 3844 -165 3852
rect -335 3810 -303 3842
rect -269 3835 -165 3844
rect -269 3810 -267 3835
rect -335 3808 -267 3810
rect -301 3801 -267 3808
rect -233 3814 -199 3835
rect -233 3801 -231 3814
rect -301 3780 -231 3801
rect -197 3780 -165 3801
rect -301 3774 -165 3780
rect -335 3771 -165 3774
rect -335 3740 -303 3771
rect -269 3766 -165 3771
rect -269 3737 -267 3766
rect -301 3732 -267 3737
rect -233 3742 -199 3766
rect -233 3732 -231 3742
rect -301 3708 -231 3732
rect -197 3708 -165 3732
rect -301 3706 -165 3708
rect -335 3698 -165 3706
rect -335 3672 -303 3698
rect -269 3697 -165 3698
rect -269 3664 -267 3697
rect -301 3663 -267 3664
rect -233 3670 -199 3697
rect -233 3663 -231 3670
rect -301 3638 -231 3663
rect -335 3636 -231 3638
rect -197 3636 -165 3663
rect -335 3628 -165 3636
rect -335 3625 -267 3628
rect -335 3604 -303 3625
rect -269 3594 -267 3625
rect -233 3598 -199 3628
rect -233 3594 -231 3598
rect -269 3591 -231 3594
rect -301 3570 -231 3591
rect -335 3564 -231 3570
rect -197 3564 -165 3594
rect -335 3559 -165 3564
rect -335 3552 -267 3559
rect -335 3536 -303 3552
rect -269 3525 -267 3552
rect -233 3526 -199 3559
rect -233 3525 -231 3526
rect -269 3518 -231 3525
rect -301 3502 -231 3518
rect -335 3492 -231 3502
rect -197 3492 -165 3525
rect -335 3490 -165 3492
rect -335 3479 -267 3490
rect -335 3468 -303 3479
rect -269 3456 -267 3479
rect -233 3456 -199 3490
rect -269 3454 -165 3456
rect -269 3445 -231 3454
rect -301 3434 -231 3445
rect -335 3421 -231 3434
rect -197 3421 -165 3454
rect -335 3406 -267 3421
rect -335 3400 -303 3406
rect -269 3387 -267 3406
rect -233 3420 -231 3421
rect -233 3387 -199 3420
rect -269 3382 -165 3387
rect -269 3372 -231 3382
rect -301 3366 -231 3372
rect -335 3352 -231 3366
rect -197 3352 -165 3382
rect -335 3333 -267 3352
rect -335 3332 -303 3333
rect -269 3318 -267 3333
rect -233 3348 -231 3352
rect -233 3318 -199 3348
rect -269 3310 -165 3318
rect -269 3299 -231 3310
rect -301 3298 -231 3299
rect -335 3283 -231 3298
rect -197 3283 -165 3310
rect -335 3264 -267 3283
rect -301 3260 -267 3264
rect -269 3249 -267 3260
rect -233 3276 -231 3283
rect -233 3249 -199 3276
rect -269 3238 -165 3249
rect -335 3226 -303 3230
rect -269 3226 -231 3238
rect -335 3214 -231 3226
rect -197 3214 -165 3238
rect -335 3196 -267 3214
rect -301 3187 -267 3196
rect -269 3180 -267 3187
rect -233 3204 -231 3214
rect -233 3180 -199 3204
rect -269 3166 -165 3180
rect -335 3153 -303 3162
rect -269 3153 -231 3166
rect -335 3145 -231 3153
rect -197 3145 -165 3166
rect -335 3128 -267 3145
rect -301 3114 -267 3128
rect -269 3111 -267 3114
rect -233 3132 -231 3145
rect -233 3111 -199 3132
rect -269 3094 -165 3111
rect -335 3080 -303 3094
rect -269 3080 -231 3094
rect -335 3076 -231 3080
rect -197 3076 -165 3094
rect -335 3060 -267 3076
rect -301 3042 -267 3060
rect -233 3060 -231 3076
rect -233 3042 -199 3060
rect -301 3041 -165 3042
rect -335 3007 -303 3026
rect -269 3022 -165 3041
rect -269 3007 -231 3022
rect -197 3007 -165 3022
rect -335 2992 -267 3007
rect -301 2973 -267 2992
rect -233 2988 -231 3007
rect -233 2973 -199 2988
rect -301 2968 -165 2973
rect -335 2934 -303 2958
rect -269 2950 -165 2968
rect -269 2938 -231 2950
rect -197 2938 -165 2950
rect -269 2934 -267 2938
rect -335 2924 -267 2934
rect -301 2904 -267 2924
rect -233 2916 -231 2938
rect -233 2904 -199 2916
rect -301 2895 -165 2904
rect -335 2861 -303 2890
rect -269 2878 -165 2895
rect -269 2869 -231 2878
rect -197 2869 -165 2878
rect -269 2861 -267 2869
rect -335 2856 -267 2861
rect -301 2835 -267 2856
rect -233 2844 -231 2869
rect -233 2835 -199 2844
rect -301 2822 -165 2835
rect -335 2788 -303 2822
rect -269 2806 -165 2822
rect -269 2800 -231 2806
rect -197 2800 -165 2806
rect -269 2788 -267 2800
rect -301 2766 -267 2788
rect -233 2772 -231 2800
rect -233 2766 -199 2772
rect -301 2754 -165 2766
rect -335 2749 -165 2754
rect -335 2720 -303 2749
rect -269 2734 -165 2749
rect -269 2731 -231 2734
rect -197 2731 -165 2734
rect -269 2715 -267 2731
rect -301 2697 -267 2715
rect -233 2700 -231 2731
rect -233 2697 -199 2700
rect -301 2686 -165 2697
rect -335 2676 -165 2686
rect -335 2652 -303 2676
rect -269 2662 -165 2676
rect -269 2642 -267 2662
rect -301 2628 -267 2642
rect -233 2628 -231 2662
rect -301 2618 -165 2628
rect -335 2603 -165 2618
rect -335 2584 -303 2603
rect -269 2593 -165 2603
rect -269 2569 -267 2593
rect -301 2559 -267 2569
rect -233 2590 -199 2593
rect -233 2559 -231 2590
rect -301 2556 -231 2559
rect -197 2556 -165 2559
rect -301 2550 -165 2556
rect -335 2530 -165 2550
rect -335 2516 -303 2530
rect -269 2524 -165 2530
rect -269 2496 -267 2524
rect -301 2490 -267 2496
rect -233 2518 -199 2524
rect -233 2490 -231 2518
rect -301 2484 -231 2490
rect -197 2484 -165 2490
rect -301 2482 -165 2484
rect -335 2457 -165 2482
rect -335 2448 -303 2457
rect -269 2455 -165 2457
rect -269 2423 -267 2455
rect -301 2421 -267 2423
rect -233 2446 -199 2455
rect -233 2421 -231 2446
rect -301 2414 -231 2421
rect -335 2412 -231 2414
rect -197 2412 -165 2421
rect -335 2386 -165 2412
rect -335 2384 -267 2386
rect -335 2380 -303 2384
rect -269 2352 -267 2384
rect -233 2374 -199 2386
rect -233 2352 -231 2374
rect -269 2350 -231 2352
rect -301 2346 -231 2350
rect -335 2340 -231 2346
rect -197 2340 -165 2352
rect -335 2317 -165 2340
rect -335 2312 -267 2317
rect -301 2311 -267 2312
rect -269 2283 -267 2311
rect -233 2302 -199 2317
rect -233 2283 -231 2302
rect -335 2277 -303 2278
rect -269 2277 -231 2283
rect -335 2268 -231 2277
rect -197 2268 -165 2283
rect -335 2248 -165 2268
rect -335 2244 -267 2248
rect -301 2238 -267 2244
rect -269 2214 -267 2238
rect -233 2230 -199 2248
rect -233 2214 -231 2230
rect -335 2204 -303 2210
rect -269 2204 -231 2214
rect -335 2196 -231 2204
rect -197 2196 -165 2214
rect -335 2179 -165 2196
rect -335 2176 -267 2179
rect -301 2165 -267 2176
rect -269 2145 -267 2165
rect -233 2158 -199 2179
rect -233 2145 -231 2158
rect -335 2131 -303 2142
rect -269 2131 -231 2145
rect -335 2124 -231 2131
rect -197 2124 -165 2145
rect -335 2110 -165 2124
rect -335 2108 -267 2110
rect -301 2092 -267 2108
rect -269 2076 -267 2092
rect -233 2086 -199 2110
rect -233 2076 -231 2086
rect -335 2058 -303 2074
rect -269 2058 -231 2076
rect -335 2052 -231 2058
rect -197 2052 -165 2076
rect -335 2041 -165 2052
rect -335 2040 -267 2041
rect -301 2019 -267 2040
rect -269 2007 -267 2019
rect -233 2014 -199 2041
rect -233 2007 -231 2014
rect -335 1985 -303 2006
rect -269 1985 -231 2007
rect -335 1980 -231 1985
rect -197 1980 -165 2007
rect -335 1972 -165 1980
rect -301 1946 -267 1972
rect -269 1938 -267 1946
rect -233 1942 -199 1972
rect -233 1938 -231 1942
rect -335 1912 -303 1938
rect -269 1912 -231 1938
rect -335 1908 -231 1912
rect -197 1908 -165 1938
rect -335 1903 -165 1908
rect -301 1873 -267 1903
rect -269 1869 -267 1873
rect -233 1870 -199 1903
rect -233 1869 -231 1870
rect -335 1839 -303 1869
rect -269 1839 -231 1869
rect -335 1836 -231 1839
rect -197 1836 -165 1869
rect -335 1834 -165 1836
rect -301 1800 -267 1834
rect -233 1800 -199 1834
rect -335 1766 -303 1800
rect -269 1798 -165 1800
rect -269 1766 -231 1798
rect -335 1765 -231 1766
rect -197 1765 -165 1798
rect -301 1731 -267 1765
rect -233 1764 -231 1765
rect -233 1731 -199 1764
rect -335 1727 -165 1731
rect -335 1696 -303 1727
rect -269 1726 -165 1727
rect -269 1696 -231 1726
rect -197 1696 -165 1726
rect -269 1693 -267 1696
rect -301 1662 -267 1693
rect -233 1692 -231 1696
rect -233 1662 -199 1692
rect -335 1654 -165 1662
rect -335 1627 -303 1654
rect -269 1627 -231 1654
rect -197 1627 -165 1654
rect -269 1620 -267 1627
rect -301 1593 -267 1620
rect -233 1620 -231 1627
rect -233 1593 -199 1620
rect -335 1581 -165 1593
rect -335 1558 -303 1581
rect -269 1558 -231 1581
rect -197 1558 -165 1581
rect -269 1547 -267 1558
rect -301 1524 -267 1547
rect -233 1547 -231 1558
rect -233 1524 -199 1547
rect -335 1508 -165 1524
rect -335 1489 -303 1508
rect -269 1489 -231 1508
rect -197 1489 -165 1508
rect -269 1474 -267 1489
rect -301 1455 -267 1474
rect -233 1474 -231 1489
rect -233 1455 -199 1474
rect -335 1435 -165 1455
rect -335 1420 -303 1435
rect -269 1420 -231 1435
rect -197 1420 -165 1435
rect -269 1401 -267 1420
rect -301 1386 -267 1401
rect -233 1401 -231 1420
rect -233 1386 -199 1401
rect -335 1362 -165 1386
rect -335 1351 -303 1362
rect -269 1351 -231 1362
rect -197 1351 -165 1362
rect -269 1328 -267 1351
rect -301 1317 -267 1328
rect -233 1328 -231 1351
rect -233 1317 -199 1328
rect -335 1289 -165 1317
rect -335 1282 -303 1289
rect -269 1282 -231 1289
rect -197 1282 -165 1289
rect -269 1255 -267 1282
rect -301 1248 -267 1255
rect -233 1255 -231 1282
rect -233 1248 -199 1255
rect -335 1216 -165 1248
rect -335 1213 -303 1216
rect -269 1213 -231 1216
rect -197 1213 -165 1216
rect -269 1182 -267 1213
rect -301 1179 -267 1182
rect -233 1182 -231 1213
rect -233 1179 -199 1182
rect -335 1144 -165 1179
rect -301 1143 -267 1144
rect -269 1110 -267 1143
rect -233 1143 -199 1144
rect -233 1110 -231 1143
rect -335 1109 -303 1110
rect -269 1109 -231 1110
rect -197 1109 -165 1110
rect -335 1075 -165 1109
rect -301 1070 -267 1075
rect -269 1041 -267 1070
rect -233 1070 -199 1075
rect -233 1041 -231 1070
rect -335 1036 -303 1041
rect -269 1036 -231 1041
rect -197 1036 -165 1041
rect -335 1006 -165 1036
rect -301 997 -267 1006
rect -269 972 -267 997
rect -233 997 -199 1006
rect -233 972 -231 997
rect -335 963 -303 972
rect -269 963 -231 972
rect -197 963 -165 972
rect -335 937 -165 963
rect -301 924 -267 937
rect -269 903 -267 924
rect -233 924 -199 937
rect -233 903 -231 924
rect -335 890 -303 903
rect -269 890 -231 903
rect -197 890 -165 903
rect -335 868 -165 890
rect -301 851 -267 868
rect -269 834 -267 851
rect -233 851 -199 868
rect -233 834 -231 851
rect -335 817 -303 834
rect -269 817 -231 834
rect -197 817 -165 834
rect -335 799 -165 817
rect -301 778 -267 799
rect -269 765 -267 778
rect -233 778 -199 799
rect -233 765 -231 778
rect -335 744 -303 765
rect -269 744 -231 765
rect -197 744 -165 765
rect -335 730 -165 744
rect -301 705 -267 730
rect -269 696 -267 705
rect -233 705 -199 730
rect -233 696 -231 705
rect -335 671 -303 696
rect -269 671 -231 696
rect -197 671 -165 696
rect -335 661 -165 671
rect -301 632 -267 661
rect -269 627 -267 632
rect -233 632 -199 661
rect -233 627 -231 632
rect -335 598 -303 627
rect -269 598 -231 627
rect -197 598 -165 627
rect -335 592 -165 598
rect -301 559 -267 592
rect -269 558 -267 559
rect -233 559 -199 592
rect -233 558 -231 559
rect -335 525 -303 558
rect -269 525 -231 558
rect -197 525 -165 558
rect -335 523 -165 525
rect -301 489 -267 523
rect -233 489 -199 523
rect -335 486 -165 489
rect -335 454 -303 486
rect -269 454 -231 486
rect -197 454 -165 486
rect -269 452 -267 454
rect -301 420 -267 452
rect -233 452 -231 454
rect -233 420 -199 452
rect -335 413 -165 420
rect -335 385 -303 413
rect -269 385 -231 413
rect -197 385 -165 413
rect -269 379 -267 385
rect -301 351 -267 379
rect -233 379 -231 385
rect -233 351 -199 379
rect -335 340 -165 351
rect -335 316 -303 340
rect -269 316 -231 340
rect -197 316 -165 340
rect -269 306 -267 316
rect -301 282 -267 306
rect -233 306 -231 316
rect -233 282 -199 306
rect -335 267 -165 282
rect -335 247 -303 267
rect -269 247 -231 267
rect -197 247 -165 267
rect -269 233 -267 247
rect -301 213 -267 233
rect -233 233 -231 247
rect -233 213 -199 233
rect -335 194 -165 213
rect -335 178 -303 194
rect -269 178 -231 194
rect -197 178 -165 194
rect -269 160 -267 178
rect -301 144 -267 160
rect -233 160 -231 178
rect -233 144 -199 160
rect -335 120 -165 144
rect 45 4596 79 4608
rect 113 4596 150 4608
rect 45 4506 77 4596
rect 184 4574 220 4608
rect 254 4574 290 4608
rect 324 4574 360 4608
rect 394 4574 430 4608
rect 464 4574 500 4608
rect 534 4574 570 4608
rect 604 4574 640 4608
rect 674 4574 710 4608
rect 744 4577 780 4608
rect 814 4577 850 4608
rect 774 4574 780 4577
rect 847 4574 850 4577
rect 884 4577 920 4608
rect 884 4574 886 4577
rect 183 4543 740 4574
rect 774 4543 813 4574
rect 847 4543 886 4574
rect 954 4577 990 4608
rect 1024 4577 1060 4608
rect 1094 4577 1130 4608
rect 1164 4577 1200 4608
rect 1234 4577 1282 4608
rect 1316 4577 1356 4608
rect 954 4574 959 4577
rect 1024 4574 1032 4577
rect 1094 4574 1105 4577
rect 1164 4574 1177 4577
rect 1234 4574 1249 4577
rect 1316 4574 1321 4577
rect 920 4543 959 4574
rect 993 4543 1032 4574
rect 1066 4543 1105 4574
rect 1139 4543 1177 4574
rect 1211 4543 1249 4574
rect 1283 4543 1321 4574
rect 1355 4574 1356 4577
rect 1390 4577 1430 4608
rect 1390 4574 1393 4577
rect 1355 4543 1393 4574
rect 1427 4574 1430 4577
rect 1464 4577 1504 4608
rect 1538 4577 1577 4608
rect 1611 4577 1645 4608
rect 1464 4574 1465 4577
rect 1427 4543 1465 4574
rect 1499 4574 1504 4577
rect 1571 4574 1577 4577
rect 1643 4575 1645 4577
rect 1679 4582 1681 4609
rect 1715 4582 1747 4616
rect 1679 4578 1747 4582
rect 1679 4575 1713 4578
rect 1499 4543 1537 4574
rect 1571 4543 1609 4574
rect 1643 4544 1713 4575
rect 1643 4543 1747 4544
rect 183 4540 1681 4543
rect 183 4506 186 4540
rect 220 4506 259 4540
rect 293 4506 332 4540
rect 366 4506 405 4540
rect 439 4506 478 4540
rect 512 4506 551 4540
rect 585 4506 624 4540
rect 658 4506 696 4540
rect 730 4506 768 4540
rect 802 4506 840 4540
rect 874 4506 912 4540
rect 946 4506 984 4540
rect 1018 4506 1056 4540
rect 1090 4506 1128 4540
rect 1162 4506 1200 4540
rect 1234 4506 1282 4540
rect 1316 4506 1355 4540
rect 1389 4506 1428 4540
rect 1462 4506 1501 4540
rect 1535 4506 1573 4540
rect 1607 4506 1645 4540
rect 1679 4509 1681 4540
rect 1715 4509 1747 4543
rect 1877 4527 2358 4865
rect 2837 4527 4047 4865
rect 4199 4527 5244 4865
rect 5350 4526 6389 4865
rect 1679 4506 1747 4509
rect 183 4505 1713 4506
rect 183 4472 740 4505
rect 774 4472 815 4505
rect 849 4472 890 4505
rect 924 4472 965 4505
rect 999 4472 1040 4505
rect 1074 4472 1115 4505
rect 1149 4472 1190 4505
rect 1224 4472 1265 4505
rect 1299 4472 1340 4505
rect 1374 4472 1415 4505
rect 1449 4472 1490 4505
rect 1524 4472 1565 4505
rect 1599 4472 1713 4505
rect 215 4438 254 4472
rect 288 4438 327 4472
rect 361 4438 400 4472
rect 434 4438 473 4472
rect 507 4438 546 4472
rect 580 4438 619 4472
rect 653 4438 692 4472
rect 726 4471 740 4472
rect 799 4471 815 4472
rect 872 4471 890 4472
rect 945 4471 965 4472
rect 1018 4471 1040 4472
rect 1090 4471 1115 4472
rect 1162 4471 1190 4472
rect 1234 4471 1265 4472
rect 1316 4471 1340 4472
rect 1394 4471 1415 4472
rect 1472 4471 1490 4472
rect 1550 4471 1565 4472
rect 726 4438 765 4471
rect 799 4438 838 4471
rect 872 4438 911 4471
rect 945 4438 984 4471
rect 1018 4438 1056 4471
rect 1090 4438 1128 4471
rect 1162 4438 1200 4471
rect 1234 4438 1282 4471
rect 1316 4438 1360 4471
rect 1394 4438 1438 4471
rect 1472 4438 1516 4471
rect 1550 4438 1593 4471
rect 1627 4438 1747 4472
rect 1877 4319 2208 4369
rect 2351 4353 4075 4369
rect 1877 4281 2242 4319
rect 1877 4247 2208 4281
rect 45 3826 77 3860
rect 183 3859 215 3894
rect 45 3758 77 3792
rect 183 3790 215 3825
rect 45 3690 77 3724
rect 183 3721 215 3756
rect 45 3622 77 3656
rect 183 3652 215 3687
rect 45 3554 77 3588
rect 183 3583 215 3618
rect 45 3486 77 3520
rect 183 3514 215 3549
rect 45 3418 77 3452
rect 183 3445 215 3480
rect 45 3350 77 3384
rect 183 3376 215 3411
rect 45 3282 77 3316
rect 183 3307 215 3342
rect 45 3214 77 3248
rect 183 3238 215 3273
rect 45 3146 77 3180
rect 183 3169 215 3204
rect 45 3078 77 3112
rect 183 3100 215 3135
rect 45 3010 77 3044
rect 183 3031 215 3066
rect 45 2942 77 2976
rect 183 2962 215 2997
rect 45 2874 77 2908
rect 183 2893 215 2928
rect 45 2806 77 2840
rect 183 2824 215 2859
rect 45 2738 77 2772
rect 183 2755 215 2790
rect 45 2670 77 2704
rect 183 2686 215 2721
rect 45 2602 77 2636
rect 183 2617 215 2652
rect 45 2534 77 2568
rect 183 2548 215 2583
rect 45 2466 77 2500
rect 183 2479 215 2514
rect 45 2398 77 2432
rect 183 2410 215 2445
rect 45 2330 77 2364
rect 183 2341 215 2376
rect 79 2307 113 2330
rect 147 2307 181 2330
rect 79 2296 215 2307
rect 45 2291 215 2296
rect 45 2262 77 2291
rect 111 2272 149 2291
rect 183 2272 215 2291
rect 111 2257 113 2272
rect 79 2238 113 2257
rect 147 2257 149 2272
rect 147 2238 181 2257
rect 79 2228 215 2238
rect 45 2218 215 2228
rect 45 2194 77 2218
rect 111 2203 149 2218
rect 183 2203 215 2218
rect 111 2184 113 2203
rect 79 2169 113 2184
rect 147 2184 149 2203
rect 147 2169 181 2184
rect 79 2160 215 2169
rect 45 2145 215 2160
rect 45 2126 77 2145
rect 111 2134 149 2145
rect 183 2134 215 2145
rect 111 2111 113 2134
rect 79 2100 113 2111
rect 147 2111 149 2134
rect 147 2100 181 2111
rect 79 2092 215 2100
rect 45 2072 215 2092
rect 45 2058 77 2072
rect 111 2065 149 2072
rect 183 2065 215 2072
rect 111 2038 113 2065
rect 79 2031 113 2038
rect 147 2038 149 2065
rect 147 2031 181 2038
rect 79 2024 215 2031
rect 45 1999 215 2024
rect 45 1990 77 1999
rect 111 1996 149 1999
rect 183 1996 215 1999
rect 111 1965 113 1996
rect 79 1962 113 1965
rect 147 1965 149 1996
rect 147 1962 181 1965
rect 79 1956 215 1962
rect 45 1927 215 1956
rect 45 1926 113 1927
rect 45 1922 77 1926
rect 111 1893 113 1926
rect 147 1926 181 1927
rect 147 1893 149 1926
rect 111 1892 149 1893
rect 183 1892 215 1893
rect 79 1888 215 1892
rect 45 1858 215 1888
rect 45 1854 113 1858
rect 79 1853 113 1854
rect 111 1824 113 1853
rect 147 1853 181 1858
rect 147 1824 149 1853
rect 45 1819 77 1820
rect 111 1819 149 1824
rect 183 1819 215 1824
rect 45 1789 215 1819
rect 45 1786 113 1789
rect 79 1780 113 1786
rect 111 1755 113 1780
rect 147 1780 181 1789
rect 147 1755 149 1780
rect 45 1746 77 1752
rect 111 1746 149 1755
rect 183 1746 215 1755
rect 45 1720 215 1746
rect 45 1718 113 1720
rect 79 1707 113 1718
rect 111 1686 113 1707
rect 147 1707 181 1720
rect 147 1686 149 1707
rect 45 1673 77 1684
rect 111 1673 149 1686
rect 183 1673 215 1686
rect 45 1651 215 1673
rect 45 1650 113 1651
rect 79 1634 113 1650
rect 111 1617 113 1634
rect 147 1634 181 1651
rect 147 1617 149 1634
rect 45 1600 77 1616
rect 111 1600 149 1617
rect 183 1600 215 1617
rect 45 1582 215 1600
rect 79 1561 113 1582
rect 111 1548 113 1561
rect 147 1561 181 1582
rect 147 1548 149 1561
rect 45 1527 77 1548
rect 111 1527 149 1548
rect 183 1527 215 1548
rect 45 1513 215 1527
rect 79 1488 113 1513
rect 111 1479 113 1488
rect 147 1488 181 1513
rect 147 1479 149 1488
rect 45 1454 77 1479
rect 111 1454 149 1479
rect 183 1454 215 1479
rect 45 1444 215 1454
rect 79 1415 113 1444
rect 111 1410 113 1415
rect 147 1415 181 1444
rect 147 1410 149 1415
rect 45 1381 77 1410
rect 111 1381 149 1410
rect 183 1381 215 1410
rect 45 1375 215 1381
rect 79 1342 113 1375
rect 111 1341 113 1342
rect 147 1342 181 1375
rect 147 1341 149 1342
rect 45 1308 77 1341
rect 111 1308 149 1341
rect 183 1308 215 1341
rect 45 1306 215 1308
rect 79 1272 113 1306
rect 147 1272 181 1306
rect 45 1269 215 1272
rect 45 1237 77 1269
rect 111 1237 149 1269
rect 183 1237 215 1269
rect 111 1235 113 1237
rect 79 1203 113 1235
rect 147 1235 149 1237
rect 147 1203 181 1235
rect 45 1196 215 1203
rect 45 1168 77 1196
rect 111 1168 149 1196
rect 183 1168 215 1196
rect 111 1162 113 1168
rect 79 1134 113 1162
rect 147 1162 149 1168
rect 147 1134 181 1162
rect 45 1123 215 1134
rect 45 1099 77 1123
rect 111 1099 149 1123
rect 183 1099 215 1123
rect 111 1089 113 1099
rect 79 1065 113 1089
rect 147 1089 149 1099
rect 147 1065 181 1089
rect 45 1050 215 1065
rect 45 1030 77 1050
rect 111 1030 149 1050
rect 183 1030 215 1050
rect 111 1016 113 1030
rect 79 996 113 1016
rect 147 1016 149 1030
rect 147 996 181 1016
rect 45 977 215 996
rect 45 961 77 977
rect 111 961 149 977
rect 183 961 215 977
rect 111 943 113 961
rect 79 927 113 943
rect 147 943 149 961
rect 147 927 181 943
rect 45 904 215 927
rect 45 892 77 904
rect 111 892 149 904
rect 183 892 215 904
rect 111 870 113 892
rect 79 858 113 870
rect 147 870 149 892
rect 147 858 181 870
rect 45 831 215 858
rect 45 823 77 831
rect 111 823 149 831
rect 183 823 215 831
rect 111 797 113 823
rect 79 789 113 797
rect 147 797 149 823
rect 147 789 181 797
rect 45 758 215 789
rect 45 754 77 758
rect 111 754 149 758
rect 183 754 215 758
rect 111 724 113 754
rect 79 720 113 724
rect 147 724 149 754
rect 147 720 181 724
rect 45 685 215 720
rect 111 651 113 685
rect 147 651 149 685
rect 45 616 215 651
rect 79 612 113 616
rect 111 582 113 612
rect 147 612 181 616
rect 147 582 149 612
rect 45 578 77 582
rect 111 578 149 582
rect 183 578 215 582
rect 45 547 215 578
rect 79 539 113 547
rect 111 513 113 539
rect 147 539 181 547
rect 147 513 149 539
rect 45 505 77 513
rect 111 505 149 513
rect 183 505 215 513
rect 45 478 215 505
rect 79 466 113 478
rect 111 444 113 466
rect 147 466 181 478
rect 147 444 149 466
rect 45 432 77 444
rect 111 432 149 444
rect 183 432 215 444
rect 45 409 215 432
rect 79 393 113 409
rect 111 375 113 393
rect 147 393 181 409
rect 147 375 149 393
rect 45 359 77 375
rect 111 359 149 375
rect 183 359 215 375
rect 45 340 215 359
rect 79 320 113 340
rect 111 306 113 320
rect 147 320 181 340
rect 367 4202 435 4226
rect 401 4192 435 4202
rect 469 4192 506 4226
rect 540 4192 577 4226
rect 611 4192 649 4226
rect 683 4192 721 4226
rect 763 4192 793 4226
rect 837 4192 865 4226
rect 911 4192 937 4226
rect 985 4192 1009 4226
rect 1059 4192 1081 4226
rect 1133 4192 1153 4226
rect 1207 4192 1225 4226
rect 1281 4192 1297 4226
rect 1355 4192 1369 4226
rect 1429 4192 1441 4226
rect 1502 4192 1513 4226
rect 1575 4192 1585 4226
rect 1648 4192 1657 4226
rect 1721 4202 1759 4226
rect 1721 4192 1725 4202
rect 367 4134 401 4168
rect 1725 4125 1759 4168
rect 367 4066 401 4100
rect 367 3998 401 4032
rect 541 4020 1491 4119
rect 1535 4037 1569 4053
rect 367 3930 401 3964
rect 367 3862 401 3896
rect 541 3942 1491 3986
rect 541 3908 555 3942
rect 589 3908 627 3942
rect 661 3908 699 3942
rect 733 3908 771 3942
rect 805 3908 843 3942
rect 877 3908 915 3942
rect 949 3908 1075 3942
rect 1109 3908 1147 3942
rect 1181 3908 1219 3942
rect 1253 3908 1291 3942
rect 1325 3908 1363 3942
rect 1397 3908 1435 3942
rect 1469 3908 1491 3942
rect 541 3864 1491 3908
rect 1535 3969 1569 4003
rect 1535 3901 1569 3935
rect 1535 3833 1569 3867
rect 1725 4048 1759 4091
rect 1877 4209 2242 4247
rect 1877 4175 2208 4209
rect 1877 4137 2242 4175
rect 1877 4103 2208 4137
rect 1877 4065 2242 4103
rect 1877 4031 2208 4065
rect 2385 4319 4075 4353
rect 2351 4281 4075 4319
rect 2385 4247 4075 4281
rect 2351 4209 4075 4247
rect 2385 4175 4075 4209
rect 2351 4137 4075 4175
rect 2385 4103 4075 4137
rect 2351 4065 4075 4103
rect 2385 4031 4075 4065
rect 4179 4366 5312 4369
rect 4179 4332 5278 4366
rect 4179 4294 5312 4332
rect 4179 4260 5278 4294
rect 4179 4222 5312 4260
rect 4179 4188 5278 4222
rect 4179 4150 5312 4188
rect 4179 4116 5278 4150
rect 4179 4078 5312 4116
rect 4179 4044 5278 4078
rect 4179 4031 5312 4044
rect 5416 4366 6389 4369
rect 5450 4332 6389 4366
rect 5416 4294 6389 4332
rect 5450 4260 6389 4294
rect 5416 4222 6389 4260
rect 5450 4188 6389 4222
rect 5416 4150 6389 4188
rect 5450 4116 6389 4150
rect 5416 4078 6389 4116
rect 5450 4044 6389 4078
rect 5416 4031 6389 4044
rect 1725 3972 1759 4014
rect 1759 3938 4780 3942
rect 1725 3908 4780 3938
rect 4814 3908 5709 3942
rect 1725 3904 5709 3908
rect 5815 3904 6303 3942
rect 1725 3870 1749 3904
rect 1783 3870 1817 3904
rect 1851 3870 1883 3904
rect 1987 3870 2021 3904
rect 2055 3870 2089 3904
rect 2123 3870 2157 3904
rect 2191 3870 2225 3904
rect 2259 3870 2293 3904
rect 2327 3870 2361 3904
rect 2395 3870 2429 3904
rect 2463 3870 2497 3904
rect 2531 3870 2565 3904
rect 2599 3870 2633 3904
rect 2667 3870 2701 3904
rect 2735 3870 2769 3904
rect 2803 3870 2837 3904
rect 2871 3870 2905 3904
rect 2939 3870 2973 3904
rect 3007 3870 3041 3904
rect 3075 3870 3109 3904
rect 3143 3870 3177 3904
rect 3211 3870 3245 3904
rect 3279 3870 3313 3904
rect 3347 3870 3381 3904
rect 3415 3870 3449 3904
rect 3483 3870 3517 3904
rect 3551 3870 3585 3904
rect 3619 3870 3653 3904
rect 3687 3870 3721 3904
rect 3755 3870 3789 3904
rect 3823 3870 3857 3904
rect 3891 3870 3925 3904
rect 3959 3870 3993 3904
rect 4027 3870 4062 3904
rect 4096 3870 4131 3904
rect 4165 3870 4200 3904
rect 4234 3870 4269 3904
rect 4303 3870 4338 3904
rect 4372 3870 4407 3904
rect 4441 3870 4476 3904
rect 4510 3870 4545 3904
rect 4579 3870 4614 3904
rect 4648 3870 4683 3904
rect 4717 3870 4752 3904
rect 4786 3870 4821 3904
rect 4855 3870 4890 3904
rect 4924 3870 4959 3904
rect 4993 3870 5028 3904
rect 5062 3870 5097 3904
rect 5131 3870 5166 3904
rect 5200 3870 5235 3904
rect 5269 3870 5304 3904
rect 5338 3870 5373 3904
rect 5407 3870 5442 3904
rect 5476 3870 5511 3904
rect 5545 3870 5580 3904
rect 5614 3870 5649 3904
rect 5683 3870 5709 3904
rect 5821 3870 5856 3904
rect 5890 3870 5925 3904
rect 5959 3870 5994 3904
rect 6028 3870 6063 3904
rect 6097 3870 6132 3904
rect 6166 3870 6201 3904
rect 6235 3886 6303 3904
rect 6235 3870 6269 3886
rect 1725 3836 1883 3870
rect 367 3794 401 3828
rect 367 3726 401 3760
rect 541 3731 1491 3830
rect 1535 3765 1569 3799
rect 1985 3836 4780 3870
rect 4814 3836 5709 3870
rect 5815 3846 6269 3870
rect 5815 3836 6303 3846
rect 1985 3802 2048 3836
rect 6269 3814 6303 3836
rect 1535 3697 1569 3731
rect 367 3658 401 3692
rect 367 3590 401 3624
rect 541 3598 1491 3697
rect 1535 3629 1569 3663
rect 367 3522 401 3556
rect 367 3454 401 3488
rect 541 3520 1491 3564
rect 541 3486 555 3520
rect 589 3486 627 3520
rect 661 3486 699 3520
rect 733 3486 771 3520
rect 805 3486 843 3520
rect 877 3486 915 3520
rect 949 3486 1075 3520
rect 1109 3486 1147 3520
rect 1181 3486 1219 3520
rect 1253 3486 1291 3520
rect 1325 3486 1363 3520
rect 1397 3486 1435 3520
rect 1469 3486 1491 3520
rect 1535 3561 1569 3595
rect 1535 3493 1569 3527
rect 1535 3452 1569 3459
rect 367 3386 401 3420
rect 367 3320 401 3352
rect 367 3250 401 3284
rect 367 3182 401 3213
rect 367 3114 401 3140
rect 367 3046 401 3067
rect 458 3425 1569 3452
rect 458 3418 1535 3425
rect 458 3382 507 3418
rect 458 3348 463 3382
rect 497 3348 507 3382
rect 1535 3375 1569 3391
rect 1705 3746 1743 3780
rect 1777 3746 1815 3780
rect 458 3310 507 3348
rect 458 3276 463 3310
rect 497 3276 507 3310
rect 541 3309 1491 3364
rect 458 3238 507 3276
rect 458 3204 463 3238
rect 497 3204 507 3238
rect 458 3166 507 3204
rect 604 3226 1297 3275
rect 604 3192 757 3226
rect 791 3192 829 3226
rect 863 3192 901 3226
rect 935 3192 973 3226
rect 1007 3192 1045 3226
rect 1079 3192 1117 3226
rect 1151 3213 1297 3226
rect 1151 3192 1243 3213
rect 604 3176 1243 3192
rect 458 3132 463 3166
rect 497 3132 507 3166
rect 458 3094 507 3132
rect 1233 3148 1243 3176
rect 1277 3148 1297 3213
rect 1233 3145 1297 3148
rect 458 3060 463 3094
rect 497 3060 507 3094
rect 604 3098 1199 3119
rect 638 3064 676 3098
rect 710 3064 748 3098
rect 782 3064 820 3098
rect 854 3064 1199 3098
rect 604 3020 1199 3064
rect 1233 3111 1243 3145
rect 1277 3111 1297 3145
rect 1233 3110 1297 3111
rect 1233 3076 1243 3110
rect 1277 3076 1297 3110
rect 1233 3038 1297 3076
rect 367 2978 401 2994
rect 1233 3003 1243 3038
rect 1277 3003 1297 3038
rect 367 2910 401 2921
rect 657 2942 1199 2986
rect 657 2908 981 2942
rect 1015 2908 1053 2942
rect 1087 2908 1125 2942
rect 1159 2908 1199 2942
rect 657 2864 1199 2908
rect 1233 2942 1297 3003
rect 1233 2908 1243 2942
rect 1277 2908 1297 2942
rect 367 2842 401 2848
rect 1233 2847 1297 2908
rect 367 2774 401 2775
rect 367 2736 401 2740
rect 604 2786 1199 2830
rect 638 2752 676 2786
rect 710 2752 748 2786
rect 782 2752 820 2786
rect 854 2752 1199 2786
rect 604 2708 1199 2752
rect 1233 2813 1243 2847
rect 1277 2813 1297 2847
rect 1233 2725 1297 2813
rect 1233 2691 1243 2725
rect 1277 2691 1297 2725
rect 367 2663 401 2672
rect 367 2590 401 2604
rect 657 2630 1199 2674
rect 657 2596 894 2630
rect 928 2596 966 2630
rect 1000 2596 1038 2630
rect 1072 2596 1199 2630
rect 657 2552 1199 2596
rect 1233 2630 1297 2691
rect 1233 2596 1243 2630
rect 1277 2596 1297 2630
rect 367 2517 401 2536
rect 1233 2535 1297 2596
rect 367 2444 401 2468
rect 367 2371 401 2400
rect 604 2474 1199 2518
rect 638 2440 676 2474
rect 710 2440 748 2474
rect 782 2440 820 2474
rect 854 2440 1199 2474
rect 604 2396 1199 2440
rect 1233 2501 1243 2535
rect 1277 2501 1297 2535
rect 1233 2413 1297 2501
rect 1233 2379 1243 2413
rect 1277 2379 1297 2413
rect 367 2298 401 2332
rect 367 2230 401 2264
rect 657 2318 1199 2362
rect 657 2284 981 2318
rect 1015 2284 1053 2318
rect 1087 2284 1125 2318
rect 1159 2284 1199 2318
rect 657 2240 1199 2284
rect 1233 2341 1297 2379
rect 1233 2307 1243 2341
rect 1277 2307 1297 2341
rect 1233 2269 1297 2307
rect 1233 2227 1243 2269
rect 1277 2227 1297 2269
rect 367 2162 401 2191
rect 367 2094 401 2118
rect 604 2162 1199 2206
rect 638 2128 676 2162
rect 710 2128 748 2162
rect 782 2128 820 2162
rect 854 2128 1199 2162
rect 604 2084 1199 2128
rect 1233 2197 1297 2227
rect 1233 2155 1243 2197
rect 1277 2155 1297 2197
rect 1233 2125 1297 2155
rect 1233 2083 1243 2125
rect 1277 2083 1297 2125
rect 1233 2053 1297 2083
rect 367 2026 401 2045
rect 367 1958 401 1972
rect 657 2006 1199 2050
rect 657 1972 981 2006
rect 1015 1972 1053 2006
rect 1087 1972 1125 2006
rect 1159 1972 1199 2006
rect 657 1928 1199 1972
rect 1233 2011 1243 2053
rect 1277 2011 1297 2053
rect 1233 1982 1297 2011
rect 1233 1939 1243 1982
rect 1277 1939 1297 1982
rect 367 1890 401 1899
rect 1233 1911 1297 1939
rect 367 1822 401 1826
rect 604 1795 1199 1894
rect 1233 1867 1243 1911
rect 1277 1867 1297 1911
rect 1233 1861 1297 1867
rect 1331 3181 1637 3205
rect 1365 3147 1399 3181
rect 1433 3147 1467 3181
rect 1501 3147 1535 3181
rect 1569 3147 1603 3181
rect 1331 3110 1637 3147
rect 1365 3076 1399 3110
rect 1433 3076 1467 3110
rect 1501 3107 1637 3110
rect 1501 3076 1535 3107
rect 1331 3073 1535 3076
rect 1569 3073 1603 3107
rect 1331 3039 1637 3073
rect 1365 3005 1399 3039
rect 1433 3005 1467 3039
rect 1501 3033 1637 3039
rect 1501 3005 1535 3033
rect 1331 2999 1535 3005
rect 1569 2999 1603 3033
rect 1331 2968 1637 2999
rect 1365 2934 1399 2968
rect 1433 2934 1467 2968
rect 1501 2959 1637 2968
rect 1501 2934 1535 2959
rect 1331 2925 1535 2934
rect 1569 2925 1603 2959
rect 1331 2897 1637 2925
rect 1365 2863 1399 2897
rect 1433 2863 1467 2897
rect 1501 2885 1637 2897
rect 1501 2863 1535 2885
rect 1331 2851 1535 2863
rect 1569 2851 1603 2885
rect 1331 2826 1637 2851
rect 1365 2792 1399 2826
rect 1433 2792 1467 2826
rect 1501 2811 1637 2826
rect 1501 2792 1535 2811
rect 1331 2777 1535 2792
rect 1569 2777 1603 2811
rect 1331 2755 1637 2777
rect 1365 2721 1399 2755
rect 1433 2721 1467 2755
rect 1501 2737 1637 2755
rect 1501 2721 1535 2737
rect 1331 2703 1535 2721
rect 1569 2703 1603 2737
rect 1331 2684 1637 2703
rect 1365 2650 1399 2684
rect 1433 2650 1467 2684
rect 1501 2663 1637 2684
rect 1501 2650 1535 2663
rect 1331 2629 1535 2650
rect 1569 2629 1603 2663
rect 1331 2613 1637 2629
rect 1365 2579 1399 2613
rect 1433 2579 1467 2613
rect 1501 2589 1637 2613
rect 1501 2579 1535 2589
rect 1331 2555 1535 2579
rect 1569 2555 1603 2589
rect 1331 2542 1637 2555
rect 1365 2508 1399 2542
rect 1433 2508 1467 2542
rect 1501 2515 1637 2542
rect 1501 2508 1535 2515
rect 1331 2481 1535 2508
rect 1569 2481 1603 2515
rect 1331 2471 1637 2481
rect 1365 2437 1399 2471
rect 1433 2437 1467 2471
rect 1501 2442 1637 2471
rect 1501 2437 1535 2442
rect 1331 2408 1535 2437
rect 1569 2408 1603 2442
rect 1331 2400 1637 2408
rect 1365 2366 1399 2400
rect 1433 2366 1467 2400
rect 1501 2384 1637 2400
rect 1331 2328 1501 2366
rect 1365 2294 1399 2328
rect 1433 2294 1467 2328
rect 1671 2319 1849 3746
rect 1883 3765 2048 3802
rect 1917 3731 1951 3765
rect 1985 3731 2048 3765
rect 1883 3694 2048 3731
rect 2101 3727 2135 3731
rect 1917 3660 1951 3694
rect 1985 3660 2048 3694
rect 1883 3623 2048 3660
rect 1917 3589 1951 3623
rect 1985 3589 2048 3623
rect 1883 3552 2048 3589
rect 1917 3518 1951 3552
rect 1985 3518 2048 3552
rect 1883 3481 2048 3518
rect 1917 3447 1951 3481
rect 1985 3447 2048 3481
rect 1883 3410 2048 3447
rect 1917 3376 1951 3410
rect 1985 3376 2048 3410
rect 1883 3339 2048 3376
rect 1917 3305 1951 3339
rect 1985 3305 2048 3339
rect 1883 3268 2048 3305
rect 1917 3234 1951 3268
rect 1985 3234 2048 3268
rect 1883 3197 2048 3234
rect 1917 3163 1951 3197
rect 1985 3163 2048 3197
rect 1883 3126 2048 3163
rect 1917 3092 1951 3126
rect 1985 3092 2048 3126
rect 1883 3055 2048 3092
rect 1917 3021 1951 3055
rect 1985 3021 2048 3055
rect 1883 2984 2048 3021
rect 1917 2950 1951 2984
rect 1985 2950 2048 2984
rect 1883 2913 2048 2950
rect 1917 2879 1951 2913
rect 1985 2879 2048 2913
rect 1883 2842 2048 2879
rect 1917 2808 1951 2842
rect 1985 2808 2048 2842
rect 1883 2771 2048 2808
rect 1917 2737 1951 2771
rect 1985 2737 2048 2771
rect 1883 2699 2048 2737
rect 1917 2665 1951 2699
rect 1985 2665 2048 2699
rect 1883 2627 2048 2665
rect 2082 3715 2155 3727
rect 2082 3681 2101 3715
rect 2135 3681 2155 3715
rect 2245 3703 6187 3802
rect 6269 3744 6303 3778
rect 2082 3620 2155 3681
rect 6269 3675 6303 3708
rect 2082 3593 2101 3620
rect 2082 3559 2100 3593
rect 2135 3586 2155 3620
rect 2134 3559 2155 3586
rect 2082 3525 2155 3559
rect 2245 3620 6187 3669
rect 2245 3586 4893 3620
rect 4927 3586 4965 3620
rect 4999 3586 5504 3620
rect 5538 3586 5576 3620
rect 5610 3586 5648 3620
rect 5682 3586 5720 3620
rect 5754 3586 5792 3620
rect 5826 3586 6187 3620
rect 2245 3547 6187 3586
rect 6269 3606 6303 3636
rect 2082 3521 2101 3525
rect 2082 3487 2100 3521
rect 2135 3491 2155 3525
rect 6269 3537 6303 3564
rect 2134 3487 2155 3491
rect 2082 3293 2155 3487
rect 2245 3414 6187 3513
rect 6269 3468 6303 3492
rect 6269 3399 6303 3420
rect 2082 3259 2101 3293
rect 2135 3259 2155 3293
rect 2245 3276 6187 3375
rect 6269 3330 6303 3348
rect 2082 3198 2155 3259
rect 6269 3261 6303 3276
rect 2082 3164 2101 3198
rect 2135 3164 2155 3198
rect 2082 3103 2155 3164
rect 2245 3120 6187 3242
rect 6269 3192 6303 3204
rect 6269 3123 6303 3132
rect 2082 3069 2101 3103
rect 2135 3069 2155 3103
rect 2082 2871 2155 3069
rect 2245 2987 6187 3086
rect 6269 3054 6303 3059
rect 6269 2985 6303 2986
rect 2082 2837 2101 2871
rect 2135 2837 2155 2871
rect 2245 2854 6187 2953
rect 6269 2947 6303 2951
rect 6269 2874 6303 2882
rect 2082 2776 2155 2837
rect 2082 2742 2101 2776
rect 2135 2742 2155 2776
rect 2082 2681 2155 2742
rect 2242 2698 6187 2820
rect 6269 2801 6303 2813
rect 6269 2728 6303 2744
rect 2082 2647 2101 2681
rect 2135 2647 2155 2681
rect 2082 2631 2155 2647
rect 1917 2593 1951 2627
rect 1985 2593 2048 2627
rect 1883 2555 2048 2593
rect 2245 2565 6187 2664
rect 6269 2655 6303 2675
rect 6269 2582 6303 2606
rect 1917 2521 1951 2555
rect 1985 2531 2048 2555
rect 6269 2531 6303 2537
rect 1985 2521 6303 2531
rect 1883 2509 6303 2521
rect 1883 2492 6269 2509
rect 1883 2483 1906 2492
rect 1940 2483 2045 2492
rect 1940 2458 1951 2483
rect 1917 2449 1951 2458
rect 1985 2458 2045 2483
rect 2079 2458 2118 2492
rect 2152 2458 2191 2492
rect 2241 2458 2264 2492
rect 2309 2458 2337 2492
rect 2377 2458 2410 2492
rect 2445 2458 2479 2492
rect 2517 2458 2547 2492
rect 2590 2458 2615 2492
rect 2663 2458 2683 2492
rect 2736 2458 2751 2492
rect 2809 2458 2820 2492
rect 2882 2458 2889 2492
rect 2955 2458 2958 2492
rect 2992 2458 2994 2492
rect 3061 2458 3067 2492
rect 3130 2458 3140 2492
rect 3199 2458 3213 2492
rect 3268 2458 3286 2492
rect 3337 2458 3359 2492
rect 3406 2458 3432 2492
rect 3475 2458 3505 2492
rect 3544 2458 3578 2492
rect 3613 2458 3648 2492
rect 3685 2458 3717 2492
rect 3757 2458 3786 2492
rect 3829 2458 3855 2492
rect 3901 2458 3924 2492
rect 3973 2458 3993 2492
rect 4045 2458 4062 2492
rect 4117 2458 4131 2492
rect 4189 2458 4200 2492
rect 4261 2458 4269 2492
rect 4333 2458 4338 2492
rect 4405 2458 4407 2492
rect 4441 2458 4443 2492
rect 4510 2458 4515 2492
rect 4579 2458 4587 2492
rect 4648 2458 4659 2492
rect 4717 2458 4752 2492
rect 4786 2458 4821 2492
rect 4855 2458 4890 2492
rect 4924 2458 4959 2492
rect 4993 2458 5028 2492
rect 5062 2458 5097 2492
rect 5131 2458 5166 2492
rect 5200 2458 5235 2492
rect 5269 2458 5304 2492
rect 5338 2458 5373 2492
rect 5407 2458 5442 2492
rect 5476 2458 5511 2492
rect 5545 2458 5580 2492
rect 5614 2458 5649 2492
rect 5683 2458 5718 2492
rect 5752 2458 5787 2492
rect 5821 2458 5856 2492
rect 5890 2458 5925 2492
rect 5959 2458 5994 2492
rect 6028 2458 6063 2492
rect 6097 2458 6132 2492
rect 6166 2458 6201 2492
rect 6235 2468 6269 2492
rect 6235 2458 6303 2468
rect 1985 2449 6303 2458
rect 1883 2442 6303 2449
rect 1883 2420 2048 2442
rect 1883 2411 1906 2420
rect 1940 2411 2048 2420
rect 1940 2386 1951 2411
rect 1917 2377 1951 2386
rect 1985 2377 2048 2411
rect 6269 2436 6303 2442
rect 1883 2353 2048 2377
rect 2245 2364 6187 2408
rect 2245 2330 5504 2364
rect 5538 2330 5576 2364
rect 5610 2330 5648 2364
rect 5682 2330 5720 2364
rect 5754 2330 5792 2364
rect 5826 2330 6187 2364
rect 1331 2256 1501 2294
rect 1365 2222 1399 2256
rect 1433 2222 1467 2256
rect 1331 2184 1501 2222
rect 1365 2150 1399 2184
rect 1433 2150 1467 2184
rect 1331 2112 1501 2150
rect 1365 2078 1399 2112
rect 1433 2078 1467 2112
rect 1331 2040 1501 2078
rect 1365 2006 1399 2040
rect 1433 2006 1467 2040
rect 1331 1968 1501 2006
rect 1365 1934 1399 1968
rect 1433 1934 1467 1968
rect 1331 1896 1501 1934
rect 1365 1862 1399 1896
rect 1433 1862 1467 1896
rect 1331 1838 1501 1862
rect 1535 2303 2135 2319
rect 1535 2269 2101 2303
rect 2245 2286 6187 2330
rect 6269 2364 6303 2399
rect 6269 2295 6303 2329
rect 1535 2263 2135 2269
rect 367 1787 401 1788
rect 367 1714 401 1720
rect 541 1662 1491 1761
rect 1535 1679 1596 2263
rect 2084 2233 2135 2263
rect 2084 2199 2101 2233
rect 367 1641 401 1652
rect 1569 1645 1596 1679
rect 367 1567 401 1584
rect 367 1493 401 1516
rect 541 1584 1491 1628
rect 541 1550 1040 1584
rect 1074 1550 1112 1584
rect 1146 1550 1184 1584
rect 1218 1550 1256 1584
rect 1290 1550 1328 1584
rect 1362 1550 1400 1584
rect 1434 1550 1491 1584
rect 541 1506 1491 1550
rect 1535 1608 1596 1645
rect 1569 1574 1596 1608
rect 1535 1537 1596 1574
rect 1569 1503 1596 1537
rect 367 1419 401 1448
rect 367 1346 401 1380
rect 541 1428 1491 1472
rect 541 1394 604 1428
rect 638 1394 676 1428
rect 710 1394 748 1428
rect 782 1394 820 1428
rect 854 1394 1235 1428
rect 1269 1394 1307 1428
rect 1341 1394 1379 1428
rect 1413 1394 1451 1428
rect 1485 1394 1491 1428
rect 541 1350 1491 1394
rect 1535 1466 1596 1503
rect 1569 1432 1596 1466
rect 1535 1395 1596 1432
rect 1569 1361 1596 1395
rect 1535 1324 1596 1361
rect 367 1278 401 1311
rect 367 1210 401 1237
rect 541 1194 1491 1316
rect 1569 1290 1596 1324
rect 1535 1253 1596 1290
rect 1569 1219 1596 1253
rect 367 1142 401 1163
rect 1535 1183 1596 1219
rect 367 1074 401 1089
rect 541 1116 1491 1160
rect 541 1082 604 1116
rect 638 1082 676 1116
rect 710 1082 748 1116
rect 782 1082 820 1116
rect 854 1082 1235 1116
rect 1269 1082 1307 1116
rect 1341 1082 1379 1116
rect 1413 1082 1451 1116
rect 1485 1082 1491 1116
rect 541 1038 1491 1082
rect 1569 1149 1596 1183
rect 1535 1113 1596 1149
rect 1569 1079 1596 1113
rect 1535 1043 1596 1079
rect 367 1006 401 1015
rect 1569 1009 1596 1043
rect 367 938 401 941
rect 367 901 401 904
rect 541 882 1491 1004
rect 1535 973 1596 1009
rect 1569 939 1596 973
rect 1535 903 1596 939
rect 1569 869 1596 903
rect 367 827 401 836
rect 367 753 401 768
rect 541 726 1491 848
rect 1535 833 1596 869
rect 1569 799 1596 833
rect 1535 763 1596 799
rect 1569 729 1596 763
rect 367 679 401 699
rect 1535 693 1596 729
rect 367 605 401 630
rect 541 570 1491 692
rect 1569 659 1596 693
rect 1535 623 1596 659
rect 1569 589 1596 623
rect 367 531 401 561
rect 1535 553 1596 589
rect 367 457 401 492
rect 367 388 401 423
rect 367 330 401 349
rect 435 489 463 523
rect 497 489 507 523
rect 435 451 507 489
rect 435 417 463 451
rect 497 417 507 451
rect 147 306 149 320
rect 45 286 77 306
rect 111 286 149 306
rect 183 286 215 306
rect 45 271 215 286
rect 79 247 113 271
rect 111 237 113 247
rect 147 247 181 271
rect 147 237 149 247
rect 45 213 77 237
rect 111 213 149 237
rect 183 213 215 237
rect 45 202 215 213
rect 79 174 113 202
rect 111 168 113 174
rect 147 174 181 202
rect 147 168 149 174
rect 435 274 507 417
rect 541 414 1491 536
rect 1569 519 1596 553
rect 1535 503 1596 519
rect 1630 2144 2050 2168
rect 1630 1226 1653 2144
rect 2027 1226 2050 2144
rect 1630 1191 2050 1226
rect 1630 1157 1653 1191
rect 1687 1157 1721 1191
rect 1755 1157 1789 1191
rect 1823 1157 1857 1191
rect 1891 1157 1925 1191
rect 1959 1157 1993 1191
rect 2027 1157 2050 1191
rect 1630 1122 2050 1157
rect 1630 1088 1653 1122
rect 1687 1088 1721 1122
rect 1755 1088 1789 1122
rect 1823 1088 1857 1122
rect 1891 1088 1925 1122
rect 1959 1088 1993 1122
rect 2027 1088 2050 1122
rect 1630 1053 2050 1088
rect 1630 1019 1653 1053
rect 1687 1019 1721 1053
rect 1755 1019 1789 1053
rect 1823 1019 1857 1053
rect 1891 1019 1925 1053
rect 1959 1019 1993 1053
rect 2027 1019 2050 1053
rect 1630 984 2050 1019
rect 1630 950 1653 984
rect 1687 950 1721 984
rect 1755 950 1789 984
rect 1823 950 1857 984
rect 1891 950 1925 984
rect 1959 950 1993 984
rect 2027 950 2050 984
rect 1630 915 2050 950
rect 1630 881 1653 915
rect 1687 881 1721 915
rect 1755 881 1789 915
rect 1823 881 1857 915
rect 1891 881 1925 915
rect 1959 881 1993 915
rect 2027 881 2050 915
rect 1630 846 2050 881
rect 1630 812 1653 846
rect 1687 812 1721 846
rect 1755 812 1789 846
rect 1823 812 1857 846
rect 1891 812 1925 846
rect 1959 812 1993 846
rect 2027 812 2050 846
rect 1630 777 2050 812
rect 1630 743 1653 777
rect 1687 743 1721 777
rect 1755 743 1789 777
rect 1823 743 1857 777
rect 1891 743 1925 777
rect 1959 743 1993 777
rect 2027 743 2050 777
rect 1630 708 2050 743
rect 1630 674 1653 708
rect 1687 674 1721 708
rect 1755 674 1789 708
rect 1823 674 1857 708
rect 1891 674 1925 708
rect 1959 674 1993 708
rect 2027 674 2050 708
rect 1630 639 2050 674
rect 1630 605 1653 639
rect 1687 605 1721 639
rect 1755 605 1789 639
rect 1823 605 1857 639
rect 1891 605 1925 639
rect 1959 605 1993 639
rect 2027 605 2050 639
rect 1630 570 2050 605
rect 1630 536 1653 570
rect 1687 536 1721 570
rect 1755 536 1789 570
rect 1823 536 1857 570
rect 1891 536 1925 570
rect 1959 536 1993 570
rect 2027 536 2050 570
rect 1630 501 2050 536
rect 2084 2163 2135 2199
rect 2084 2129 2101 2163
rect 2245 2130 6187 2252
rect 6269 2226 6303 2256
rect 6269 2157 6303 2183
rect 2084 2093 2135 2129
rect 2084 2059 2101 2093
rect 2084 2023 2135 2059
rect 2084 1989 2101 2023
rect 2084 1953 2135 1989
rect 2245 2052 6187 2096
rect 2245 2018 5504 2052
rect 5538 2018 5576 2052
rect 5610 2018 5648 2052
rect 5682 2018 5720 2052
rect 5754 2018 5792 2052
rect 5826 2018 6187 2052
rect 2245 1974 6187 2018
rect 6269 2088 6303 2110
rect 6269 2019 6303 2037
rect 2084 1919 2101 1953
rect 6269 1950 6303 1964
rect 2084 1883 2135 1919
rect 2084 1849 2101 1883
rect 2084 1813 2135 1849
rect 2245 1818 6187 1940
rect 6269 1881 6303 1891
rect 2084 1779 2101 1813
rect 6269 1812 6303 1818
rect 2084 1743 2135 1779
rect 2084 1709 2101 1743
rect 2084 1673 2135 1709
rect 2084 1639 2101 1673
rect 2245 1740 6187 1784
rect 2245 1706 5504 1740
rect 5538 1706 5576 1740
rect 5610 1706 5648 1740
rect 5682 1706 5720 1740
rect 5754 1706 5792 1740
rect 5826 1706 6187 1740
rect 2245 1662 6187 1706
rect 6269 1743 6303 1745
rect 6269 1706 6303 1709
rect 2084 1603 2135 1639
rect 6269 1633 6303 1640
rect 2084 1569 2101 1603
rect 2084 1533 2135 1569
rect 2084 1499 2101 1533
rect 2245 1506 6187 1628
rect 6269 1560 6303 1571
rect 2084 1463 2135 1499
rect 6269 1487 6303 1502
rect 2084 1429 2101 1463
rect 2084 1393 2135 1429
rect 2084 1359 2101 1393
rect 2084 1323 2135 1359
rect 2245 1428 6187 1472
rect 2245 1394 5504 1428
rect 5538 1394 5576 1428
rect 5610 1394 5648 1428
rect 5682 1394 5720 1428
rect 5754 1394 5792 1428
rect 5826 1394 6187 1428
rect 2245 1350 6187 1394
rect 6269 1414 6303 1433
rect 2084 1289 2101 1323
rect 6269 1341 6303 1364
rect 2084 1253 2135 1289
rect 2084 1219 2101 1253
rect 2084 1183 2135 1219
rect 2245 1194 6187 1316
rect 6269 1268 6303 1295
rect 6269 1195 6303 1226
rect 2084 1149 2101 1183
rect 2084 1113 2135 1149
rect 2084 1079 2101 1113
rect 2084 1043 2135 1079
rect 2084 1009 2101 1043
rect 2245 1116 6187 1160
rect 2245 1082 5504 1116
rect 5538 1082 5576 1116
rect 5610 1082 5648 1116
rect 5682 1082 5720 1116
rect 5754 1082 5792 1116
rect 5826 1082 6187 1116
rect 2245 1038 6187 1082
rect 6269 1122 6303 1157
rect 6269 1053 6303 1088
rect 2084 973 2135 1009
rect 2084 939 2101 973
rect 2084 903 2135 939
rect 2084 869 2101 903
rect 2245 960 6187 1004
rect 2245 926 5134 960
rect 5168 926 5206 960
rect 5240 926 5278 960
rect 5312 926 5350 960
rect 5384 926 5422 960
rect 5456 926 6187 960
rect 2245 882 6187 926
rect 6269 984 6303 1015
rect 6521 3503 6559 3537
rect 6487 3462 6593 3503
rect 6521 3428 6559 3462
rect 6487 3387 6593 3428
rect 6521 3353 6559 3387
rect 6487 3312 6593 3353
rect 6521 3278 6559 3312
rect 6487 3238 6593 3278
rect 6521 3204 6559 3238
rect 6487 3164 6593 3204
rect 6521 3130 6559 3164
rect 6487 3090 6593 3130
rect 6521 3056 6559 3090
rect 6487 3016 6593 3056
rect 6521 2982 6559 3016
rect 6487 2942 6593 2982
rect 6521 2908 6559 2942
rect 6487 2868 6593 2908
rect 6521 2834 6559 2868
rect 6487 2794 6593 2834
rect 6521 2760 6559 2794
rect 6487 2720 6593 2760
rect 6521 2686 6559 2720
rect 6487 2646 6593 2686
rect 6521 2612 6559 2646
rect 6487 2572 6593 2612
rect 6521 2538 6559 2572
rect 6487 2498 6593 2538
rect 6521 2464 6559 2498
rect 6487 2424 6593 2464
rect 6521 2390 6559 2424
rect 6487 2350 6593 2390
rect 6521 2316 6559 2350
rect 6487 2276 6593 2316
rect 6521 2242 6559 2276
rect 6487 2202 6593 2242
rect 6521 2168 6559 2202
rect 6487 2128 6593 2168
rect 6521 2094 6559 2128
rect 6487 2054 6593 2094
rect 6521 2020 6559 2054
rect 25234 2058 25268 5712
rect 25914 2058 25938 6444
rect 6487 1980 6593 2020
rect 25234 2023 25792 2058
rect 25898 2023 25938 2058
rect 6521 1946 6559 1980
rect 25234 1989 25268 2023
rect 25302 1989 25336 2023
rect 25370 1989 25404 2023
rect 25438 1989 25472 2023
rect 25506 1989 25540 2023
rect 25574 1989 25608 2023
rect 25642 1989 25676 2023
rect 25710 1989 25744 2023
rect 25778 1989 25792 2023
rect 25914 1989 25938 2023
rect 6487 1906 6593 1946
rect 25234 1954 25792 1989
rect 25898 1954 25938 1989
rect 6521 1872 6559 1906
rect 25234 1920 25268 1954
rect 25302 1920 25336 1954
rect 25370 1920 25404 1954
rect 25438 1920 25472 1954
rect 25506 1920 25540 1954
rect 25574 1920 25608 1954
rect 25642 1920 25676 1954
rect 25710 1920 25744 1954
rect 25778 1920 25792 1954
rect 25914 1920 25938 1954
rect 6487 1832 6593 1872
rect 25234 1885 25792 1920
rect 25898 1885 25938 1920
rect 6521 1798 6559 1832
rect 25234 1851 25268 1885
rect 25302 1851 25336 1885
rect 25370 1851 25404 1885
rect 25438 1851 25472 1885
rect 25506 1851 25540 1885
rect 25574 1851 25608 1885
rect 25642 1851 25676 1885
rect 25710 1851 25744 1885
rect 25778 1851 25792 1885
rect 25914 1851 25938 1885
rect 6487 1758 6593 1798
rect 25234 1816 25792 1851
rect 25898 1816 25938 1851
rect 6521 1724 6559 1758
rect 25234 1782 25268 1816
rect 25302 1782 25336 1816
rect 25370 1782 25404 1816
rect 25438 1782 25472 1816
rect 25506 1782 25540 1816
rect 25574 1782 25608 1816
rect 25642 1782 25676 1816
rect 25710 1782 25744 1816
rect 25778 1782 25792 1816
rect 25914 1782 25938 1816
rect 25234 1747 25792 1782
rect 25898 1747 25938 1782
rect 6487 1684 6593 1724
rect 25234 1713 25268 1747
rect 25302 1713 25336 1747
rect 25370 1713 25404 1747
rect 25438 1713 25472 1747
rect 25506 1713 25540 1747
rect 25574 1713 25608 1747
rect 25642 1713 25676 1747
rect 25710 1713 25744 1747
rect 25778 1713 25792 1747
rect 25914 1713 25938 1747
rect 6521 1650 6559 1684
rect 25234 1678 25792 1713
rect 25898 1678 25938 1713
rect 6487 1610 6593 1650
rect 25234 1644 25268 1678
rect 25302 1644 25336 1678
rect 25370 1644 25404 1678
rect 25438 1644 25472 1678
rect 25506 1644 25540 1678
rect 25574 1644 25608 1678
rect 25642 1644 25676 1678
rect 25710 1644 25744 1678
rect 25778 1644 25792 1678
rect 25914 1644 25938 1678
rect 6521 1576 6559 1610
rect 25234 1609 25792 1644
rect 25898 1609 25938 1644
rect 6487 1536 6593 1576
rect 25234 1575 25268 1609
rect 25302 1575 25336 1609
rect 25370 1575 25404 1609
rect 25438 1575 25472 1609
rect 25506 1575 25540 1609
rect 25574 1575 25608 1609
rect 25642 1575 25676 1609
rect 25710 1575 25744 1609
rect 25778 1575 25792 1609
rect 25914 1575 25938 1609
rect 6521 1502 6559 1536
rect 25234 1540 25792 1575
rect 25898 1540 25938 1575
rect 6487 1462 6593 1502
rect 25234 1506 25268 1540
rect 25302 1506 25336 1540
rect 25370 1506 25404 1540
rect 25438 1506 25472 1540
rect 25506 1506 25540 1540
rect 25574 1506 25608 1540
rect 25642 1506 25676 1540
rect 25710 1506 25744 1540
rect 25778 1506 25792 1540
rect 25914 1506 25938 1540
rect 6521 1428 6559 1462
rect 25234 1471 25792 1506
rect 25898 1471 25938 1506
rect 6487 1388 6593 1428
rect 25234 1437 25268 1471
rect 25302 1437 25336 1471
rect 25370 1437 25404 1471
rect 25438 1437 25472 1471
rect 25506 1437 25540 1471
rect 25574 1437 25608 1471
rect 25642 1437 25676 1471
rect 25710 1437 25744 1471
rect 25778 1437 25792 1471
rect 25914 1437 25938 1471
rect 6521 1354 6559 1388
rect 25234 1402 25792 1437
rect 25898 1402 25938 1437
rect 6487 1314 6593 1354
rect 25234 1368 25268 1402
rect 25302 1368 25336 1402
rect 25370 1368 25404 1402
rect 25438 1368 25472 1402
rect 25506 1368 25540 1402
rect 25574 1368 25608 1402
rect 25642 1368 25676 1402
rect 25710 1368 25744 1402
rect 25778 1368 25792 1402
rect 25914 1368 25938 1402
rect 6521 1280 6559 1314
rect 25234 1333 25792 1368
rect 25898 1333 25938 1368
rect 6487 1240 6593 1280
rect 25234 1299 25268 1333
rect 25302 1299 25336 1333
rect 25370 1299 25404 1333
rect 25438 1299 25472 1333
rect 25506 1299 25540 1333
rect 25574 1299 25608 1333
rect 25642 1299 25676 1333
rect 25710 1299 25744 1333
rect 25778 1299 25792 1333
rect 25914 1299 25938 1333
rect 6521 1206 6559 1240
rect 25234 1264 25792 1299
rect 25898 1264 25938 1299
rect 6487 1166 6593 1206
rect 25234 1230 25268 1264
rect 25302 1230 25336 1264
rect 25370 1230 25404 1264
rect 25438 1230 25472 1264
rect 25506 1230 25540 1264
rect 25574 1230 25608 1264
rect 25642 1230 25676 1264
rect 25710 1230 25744 1264
rect 25778 1230 25792 1264
rect 25914 1230 25938 1264
rect 6521 1132 6559 1166
rect 25234 1195 25792 1230
rect 25898 1195 25938 1230
rect 25234 1161 25268 1195
rect 25302 1161 25336 1195
rect 25370 1161 25404 1195
rect 25438 1161 25472 1195
rect 25506 1161 25540 1195
rect 25574 1161 25608 1195
rect 25642 1161 25676 1195
rect 25710 1161 25744 1195
rect 25778 1161 25792 1195
rect 25914 1161 25938 1195
rect 6487 1092 6593 1132
rect 25234 1126 25792 1161
rect 25898 1126 25938 1161
rect 25234 1092 25268 1126
rect 25302 1092 25336 1126
rect 25370 1092 25404 1126
rect 25438 1092 25472 1126
rect 25506 1092 25540 1126
rect 25574 1092 25608 1126
rect 25642 1092 25676 1126
rect 25710 1092 25744 1126
rect 25778 1092 25792 1126
rect 25914 1092 25938 1126
rect 6521 1058 6559 1092
rect 6487 1018 6593 1058
rect 25234 1057 25792 1092
rect 25898 1057 25938 1092
rect 25234 1023 25268 1057
rect 25302 1023 25336 1057
rect 25370 1023 25404 1057
rect 25438 1023 25472 1057
rect 25506 1023 25540 1057
rect 25574 1023 25608 1057
rect 25642 1023 25676 1057
rect 25710 1023 25744 1057
rect 25778 1023 25792 1057
rect 25914 1023 25938 1057
rect 6521 984 6559 1018
rect 25234 988 25792 1023
rect 25898 988 25938 1023
rect 25234 954 25268 988
rect 25302 954 25336 988
rect 25370 954 25404 988
rect 25438 954 25472 988
rect 25506 954 25540 988
rect 25574 954 25608 988
rect 25642 954 25676 988
rect 25710 954 25744 988
rect 25778 954 25792 988
rect 25914 954 25938 988
rect 6269 915 6303 942
rect 25234 919 25792 954
rect 25898 919 25938 954
rect 2084 833 2135 869
rect 25234 885 25268 919
rect 25302 885 25336 919
rect 25370 885 25404 919
rect 25438 885 25472 919
rect 25506 885 25540 919
rect 25574 885 25608 919
rect 25642 885 25676 919
rect 25710 885 25744 919
rect 25778 915 25792 919
rect 25778 885 25812 915
rect 25846 885 25880 915
rect 25914 885 25938 919
rect 25234 876 25938 885
rect 2084 799 2101 833
rect 2084 763 2135 799
rect 2084 729 2101 763
rect 2084 693 2135 729
rect 2245 804 6187 848
rect 2245 770 5504 804
rect 5538 770 5576 804
rect 5610 770 5648 804
rect 5682 770 5720 804
rect 5754 770 5792 804
rect 5826 770 6187 804
rect 2245 726 6187 770
rect 6269 846 6303 869
rect 25234 850 25792 876
rect 25826 850 25864 876
rect 25898 850 25938 876
rect 25234 816 25268 850
rect 25302 816 25336 850
rect 25370 816 25404 850
rect 25438 816 25472 850
rect 25506 816 25540 850
rect 25574 816 25608 850
rect 25642 816 25676 850
rect 25710 816 25744 850
rect 25778 842 25792 850
rect 25846 842 25864 850
rect 25778 816 25812 842
rect 25846 816 25880 842
rect 25914 816 25938 850
rect 25234 803 25938 816
rect 6269 777 6303 796
rect 25234 781 25792 803
rect 25826 781 25864 803
rect 25898 781 25938 803
rect 2084 659 2101 693
rect 25234 747 25268 781
rect 25302 747 25336 781
rect 25370 747 25404 781
rect 25438 747 25472 781
rect 25506 747 25540 781
rect 25574 747 25608 781
rect 25642 747 25676 781
rect 25710 747 25744 781
rect 25778 769 25792 781
rect 25846 769 25864 781
rect 25778 747 25812 769
rect 25846 747 25880 769
rect 25914 747 25938 781
rect 25234 730 25938 747
rect 6269 708 6303 723
rect 2084 623 2135 659
rect 2084 589 2101 623
rect 2084 553 2135 589
rect 2245 648 6187 692
rect 2245 614 5134 648
rect 5168 614 5206 648
rect 5240 614 5278 648
rect 5312 614 5350 648
rect 5384 614 5422 648
rect 5456 614 6187 648
rect 2245 570 6187 614
rect 25234 712 25792 730
rect 25826 712 25864 730
rect 25898 712 25938 730
rect 25234 678 25268 712
rect 25302 678 25336 712
rect 25370 678 25404 712
rect 25438 678 25472 712
rect 25506 678 25540 712
rect 25574 678 25608 712
rect 25642 678 25676 712
rect 25710 678 25744 712
rect 25778 696 25792 712
rect 25846 696 25864 712
rect 25778 678 25812 696
rect 25846 678 25880 696
rect 25914 678 25938 712
rect 25234 657 25938 678
rect 6269 639 6303 650
rect 25234 643 25792 657
rect 25826 643 25864 657
rect 25898 643 25938 657
rect 25234 609 25268 643
rect 25302 609 25336 643
rect 25370 609 25404 643
rect 25438 609 25472 643
rect 25506 609 25540 643
rect 25574 609 25608 643
rect 25642 609 25676 643
rect 25710 609 25744 643
rect 25778 623 25792 643
rect 25846 623 25864 643
rect 25778 609 25812 623
rect 25846 609 25880 623
rect 25914 609 25938 643
rect 25234 584 25938 609
rect 6269 570 6303 577
rect 2084 519 2101 553
rect 25234 574 25792 584
rect 25826 574 25864 584
rect 25898 574 25938 584
rect 2084 503 2135 519
rect 1630 467 1653 501
rect 1687 467 1721 501
rect 1755 467 1789 501
rect 1823 467 1857 501
rect 1891 467 1925 501
rect 1959 467 1993 501
rect 2027 467 2050 501
rect 1630 432 2050 467
rect 1630 364 1653 432
rect 2027 364 2050 432
rect 2245 414 6187 536
rect 25234 540 25268 574
rect 25302 540 25336 574
rect 25370 540 25404 574
rect 25438 540 25472 574
rect 25506 540 25540 574
rect 25574 540 25608 574
rect 25642 540 25676 574
rect 25710 540 25744 574
rect 25778 550 25792 574
rect 25846 550 25864 574
rect 25778 540 25812 550
rect 25846 540 25880 550
rect 25914 540 25938 574
rect 25234 511 25938 540
rect 6269 501 6303 504
rect 25234 505 25792 511
rect 25826 505 25864 511
rect 25898 505 25938 511
rect 25234 471 25268 505
rect 25302 471 25336 505
rect 25370 471 25404 505
rect 25438 471 25472 505
rect 25506 471 25540 505
rect 25574 471 25608 505
rect 25642 471 25676 505
rect 25710 471 25744 505
rect 25778 477 25792 505
rect 25846 477 25864 505
rect 25778 471 25812 477
rect 25846 471 25880 477
rect 25914 471 25938 505
rect 6269 465 6303 467
rect 25234 438 25938 471
rect 25234 436 25792 438
rect 25826 436 25864 438
rect 25898 436 25938 438
rect 6269 364 6303 398
rect 25234 402 25268 436
rect 25302 402 25336 436
rect 25370 402 25404 436
rect 25438 402 25472 436
rect 25506 402 25540 436
rect 25574 402 25608 436
rect 25642 402 25676 436
rect 25710 402 25744 436
rect 25778 404 25792 436
rect 25846 404 25864 436
rect 25778 402 25812 404
rect 25846 402 25880 404
rect 25914 402 25938 436
rect 599 330 614 364
rect 667 330 687 364
rect 735 330 760 364
rect 803 330 833 364
rect 871 330 905 364
rect 940 330 973 364
rect 1013 330 1041 364
rect 1086 330 1109 364
rect 1159 330 1177 364
rect 1232 330 1245 364
rect 1305 330 1313 364
rect 1378 330 1381 364
rect 1415 330 1417 364
rect 1483 330 1490 364
rect 1551 330 1563 364
rect 1619 330 1636 364
rect 2034 330 2061 364
rect 2106 330 2129 364
rect 2178 330 2197 364
rect 2250 330 2265 364
rect 2322 330 2333 364
rect 2394 330 2401 364
rect 2466 330 2469 364
rect 2503 330 2504 364
rect 2571 330 2576 364
rect 2639 330 2648 364
rect 2707 330 2720 364
rect 2775 330 2792 364
rect 2843 330 2864 364
rect 2911 330 2936 364
rect 2979 330 3008 364
rect 3047 330 3080 364
rect 3115 330 3149 364
rect 3186 330 3217 364
rect 3258 330 3285 364
rect 3330 330 3353 364
rect 3402 330 3421 364
rect 3474 330 3489 364
rect 3546 330 3557 364
rect 3618 330 3625 364
rect 3690 330 3693 364
rect 3727 330 3728 364
rect 3795 330 3800 364
rect 3864 330 3872 364
rect 3933 330 3944 364
rect 4002 330 4016 364
rect 4071 330 4088 364
rect 4140 330 4160 364
rect 4209 330 4232 364
rect 4278 330 4304 364
rect 4347 330 4376 364
rect 4416 330 4448 364
rect 4485 330 4520 364
rect 4554 330 4589 364
rect 4626 330 4658 364
rect 4698 330 4727 364
rect 4761 330 4796 364
rect 4830 330 4865 364
rect 4899 330 4934 364
rect 4968 330 5003 364
rect 5037 330 5072 364
rect 5106 330 5141 364
rect 5175 330 5210 364
rect 5244 330 5279 364
rect 5313 330 5348 364
rect 5382 330 5417 364
rect 5451 330 5486 364
rect 5520 330 5555 364
rect 5589 330 5624 364
rect 5658 330 5693 364
rect 5727 330 5762 364
rect 5796 330 5831 364
rect 5865 330 5900 364
rect 5934 330 5969 364
rect 6003 330 6038 364
rect 6072 330 6107 364
rect 6141 330 6176 364
rect 6210 330 6245 364
rect 6279 330 6303 364
rect 25234 367 25938 402
rect 25234 333 25268 367
rect 25302 333 25336 367
rect 25370 333 25404 367
rect 25438 333 25472 367
rect 25506 333 25540 367
rect 25574 333 25608 367
rect 25642 333 25676 367
rect 25710 333 25744 367
rect 25778 365 25812 367
rect 25846 365 25880 367
rect 25778 333 25792 365
rect 25846 333 25864 365
rect 25914 333 25938 367
rect 25234 331 25792 333
rect 25826 331 25864 333
rect 25898 331 25938 333
rect 25234 298 25938 331
rect 435 168 677 274
rect 25234 264 25268 298
rect 25302 264 25336 298
rect 25370 264 25404 298
rect 25438 264 25472 298
rect 25506 264 25540 298
rect 25574 264 25608 298
rect 25642 264 25676 298
rect 25710 264 25744 298
rect 25778 292 25812 298
rect 25846 292 25880 298
rect 25778 264 25792 292
rect 25846 264 25864 292
rect 25914 264 25938 298
rect 25234 258 25792 264
rect 25826 258 25864 264
rect 25898 258 25938 264
rect 25234 229 25938 258
rect 25234 195 25268 229
rect 25302 195 25336 229
rect 25370 195 25404 229
rect 25438 195 25472 229
rect 25506 195 25540 229
rect 25574 195 25608 229
rect 25642 195 25676 229
rect 25710 195 25744 229
rect 25778 219 25812 229
rect 25846 219 25880 229
rect 25778 195 25792 219
rect 25846 195 25864 219
rect 25914 195 25938 229
rect 25234 185 25792 195
rect 25826 185 25864 195
rect 25898 185 25938 195
rect 45 140 77 168
rect 111 140 149 168
rect 183 140 215 168
rect 25234 160 25938 185
rect 45 134 215 140
rect 45 -36 6625 134
rect 25234 126 25268 160
rect 25302 126 25336 160
rect 25370 126 25404 160
rect 25438 126 25472 160
rect 25506 126 25540 160
rect 25574 126 25608 160
rect 25642 126 25676 160
rect 25710 126 25744 160
rect 25778 146 25812 160
rect 25846 146 25880 160
rect 25778 126 25792 146
rect 25846 126 25864 146
rect 25914 126 25938 160
rect 25234 112 25792 126
rect 25826 112 25864 126
rect 25898 112 25938 126
rect 25234 91 25938 112
rect 25234 57 25268 91
rect 25302 57 25336 91
rect 25370 57 25404 91
rect 25438 57 25472 91
rect 25506 57 25540 91
rect 25574 57 25608 91
rect 25642 57 25676 91
rect 25710 57 25744 91
rect 25778 73 25812 91
rect 25846 73 25880 91
rect 25778 57 25792 73
rect 25846 57 25864 73
rect 25914 57 25938 91
rect 25234 39 25792 57
rect 25826 39 25864 57
rect 25898 39 25938 57
rect 26149 6468 26285 6489
rect 26149 6455 26181 6468
rect 26215 6454 26253 6468
rect 26215 6434 26217 6454
rect 26183 6421 26217 6434
rect 26149 6420 26217 6421
rect 26251 6434 26253 6454
rect 26287 6434 26319 6456
rect 26251 6422 26319 6434
rect 26251 6420 26285 6422
rect 26149 6395 26285 6420
rect 26149 6386 26181 6395
rect 26215 6385 26253 6395
rect 26215 6361 26217 6385
rect 26183 6352 26217 6361
rect 26149 6351 26217 6352
rect 26251 6361 26253 6385
rect 26287 6361 26319 6388
rect 26251 6354 26319 6361
rect 26251 6351 26285 6354
rect 26149 6322 26285 6351
rect 26149 6317 26181 6322
rect 26215 6316 26253 6322
rect 26215 6288 26217 6316
rect 26183 6283 26217 6288
rect 26149 6282 26217 6283
rect 26251 6288 26253 6316
rect 26287 6288 26319 6320
rect 26251 6286 26319 6288
rect 26251 6282 26285 6286
rect 26149 6252 26285 6282
rect 26149 6249 26319 6252
rect 26149 6248 26181 6249
rect 26215 6247 26253 6249
rect 26215 6215 26217 6247
rect 26183 6214 26217 6215
rect 26149 6213 26217 6214
rect 26251 6215 26253 6247
rect 26287 6218 26319 6249
rect 26251 6213 26285 6215
rect 26149 6184 26285 6213
rect 26149 6179 26319 6184
rect 26183 6178 26319 6179
rect 26183 6176 26217 6178
rect 26149 6142 26181 6145
rect 26215 6144 26217 6176
rect 26251 6176 26319 6178
rect 26251 6144 26253 6176
rect 26287 6150 26319 6176
rect 26215 6142 26253 6144
rect 26149 6116 26285 6142
rect 26149 6110 26319 6116
rect 26183 6109 26319 6110
rect 26183 6103 26217 6109
rect 26149 6069 26181 6076
rect 26215 6075 26217 6103
rect 26251 6103 26319 6109
rect 26251 6075 26253 6103
rect 26287 6082 26319 6103
rect 26215 6069 26253 6075
rect 26149 6048 26285 6069
rect 26149 6041 26319 6048
rect 26183 6040 26319 6041
rect 26183 6030 26217 6040
rect 26149 5996 26181 6007
rect 26215 6006 26217 6030
rect 26251 6030 26319 6040
rect 26251 6006 26253 6030
rect 26287 6014 26319 6030
rect 26215 5996 26253 6006
rect 26149 5980 26285 5996
rect 26149 5972 26319 5980
rect 26183 5971 26319 5972
rect 26183 5957 26217 5971
rect 26149 5923 26181 5938
rect 26215 5937 26217 5957
rect 26251 5957 26319 5971
rect 26251 5937 26253 5957
rect 26287 5946 26319 5957
rect 26215 5923 26253 5937
rect 26149 5912 26285 5923
rect 26149 5903 26319 5912
rect 26183 5902 26319 5903
rect 26183 5884 26217 5902
rect 26149 5850 26181 5869
rect 26215 5868 26217 5884
rect 26251 5884 26319 5902
rect 26251 5868 26253 5884
rect 26287 5878 26319 5884
rect 26215 5850 26253 5868
rect 26149 5844 26285 5850
rect 26149 5834 26319 5844
rect 26183 5833 26319 5834
rect 26183 5811 26217 5833
rect 26149 5777 26181 5800
rect 26215 5799 26217 5811
rect 26251 5811 26319 5833
rect 26251 5799 26253 5811
rect 26287 5810 26319 5811
rect 26215 5777 26253 5799
rect 26149 5776 26285 5777
rect 26149 5765 26319 5776
rect 26183 5764 26319 5765
rect 26183 5738 26217 5764
rect 26149 5704 26181 5731
rect 26215 5730 26217 5738
rect 26251 5742 26319 5764
rect 26251 5738 26285 5742
rect 26251 5730 26253 5738
rect 26215 5704 26253 5730
rect 26287 5704 26319 5708
rect 26149 5696 26319 5704
rect 26183 5695 26319 5696
rect 26183 5665 26217 5695
rect 26149 5631 26181 5662
rect 26215 5661 26217 5665
rect 26251 5674 26319 5695
rect 26251 5665 26285 5674
rect 26251 5661 26253 5665
rect 26215 5631 26253 5661
rect 26287 5631 26319 5640
rect 26149 5627 26319 5631
rect 26183 5626 26319 5627
rect 26183 5593 26217 5626
rect 26149 5592 26217 5593
rect 26251 5606 26319 5626
rect 26251 5592 26285 5606
rect 26149 5558 26181 5592
rect 26215 5558 26253 5592
rect 26287 5558 26319 5572
rect 26183 5557 26319 5558
rect 26183 5524 26217 5557
rect 26149 5523 26217 5524
rect 26251 5538 26319 5557
rect 26251 5523 26285 5538
rect 26149 5519 26285 5523
rect 26149 5489 26181 5519
rect 26215 5488 26253 5519
rect 26215 5485 26217 5488
rect 26183 5455 26217 5485
rect 26149 5454 26217 5455
rect 26251 5485 26253 5488
rect 26287 5485 26319 5504
rect 26251 5470 26319 5485
rect 26251 5454 26285 5470
rect 26149 5446 26285 5454
rect 26149 5420 26181 5446
rect 26215 5419 26253 5446
rect 26215 5412 26217 5419
rect 26183 5386 26217 5412
rect 26149 5385 26217 5386
rect 26251 5412 26253 5419
rect 26287 5412 26319 5436
rect 26251 5402 26319 5412
rect 26251 5385 26285 5402
rect 26149 5373 26285 5385
rect 26149 5351 26181 5373
rect 26215 5350 26253 5373
rect 26215 5339 26217 5350
rect 26183 5317 26217 5339
rect 26149 5316 26217 5317
rect 26251 5339 26253 5350
rect 26287 5339 26319 5368
rect 26251 5334 26319 5339
rect 26251 5316 26285 5334
rect 26149 5300 26285 5316
rect 26149 5282 26181 5300
rect 26215 5281 26253 5300
rect 26215 5266 26217 5281
rect 26183 5248 26217 5266
rect 26149 5247 26217 5248
rect 26251 5266 26253 5281
rect 26287 5266 26319 5300
rect 26251 5247 26285 5266
rect 26149 5232 26285 5247
rect 26149 5227 26319 5232
rect 26149 5213 26181 5227
rect 26215 5212 26253 5227
rect 26215 5193 26217 5212
rect 26183 5179 26217 5193
rect 26149 5178 26217 5179
rect 26251 5193 26253 5212
rect 26287 5198 26319 5227
rect 26251 5178 26285 5193
rect 26149 5164 26285 5178
rect 26149 5154 26319 5164
rect 26149 5144 26181 5154
rect 26215 5143 26253 5154
rect 26215 5120 26217 5143
rect 26183 5110 26217 5120
rect 26149 5109 26217 5110
rect 26251 5120 26253 5143
rect 26287 5130 26319 5154
rect 26251 5109 26285 5120
rect 26149 5096 26285 5109
rect 26149 5081 26319 5096
rect 26149 5075 26181 5081
rect 26215 5074 26253 5081
rect 26215 5047 26217 5074
rect 26183 5041 26217 5047
rect 26149 5040 26217 5041
rect 26251 5047 26253 5074
rect 26287 5062 26319 5081
rect 26251 5040 26285 5047
rect 26149 5028 26285 5040
rect 26149 5008 26319 5028
rect 26149 5006 26181 5008
rect 26215 5005 26253 5008
rect 26215 4974 26217 5005
rect 26183 4972 26217 4974
rect 26149 4971 26217 4972
rect 26251 4974 26253 5005
rect 26287 4994 26319 5008
rect 26251 4971 26285 4974
rect 26149 4960 26285 4971
rect 26149 4937 26319 4960
rect 26183 4936 26319 4937
rect 26183 4935 26217 4936
rect 26149 4901 26181 4903
rect 26215 4902 26217 4935
rect 26251 4935 26319 4936
rect 26251 4902 26253 4935
rect 26287 4926 26319 4935
rect 26215 4901 26253 4902
rect 26149 4892 26285 4901
rect 26149 4868 26319 4892
rect 26183 4867 26319 4868
rect 26183 4862 26217 4867
rect 26149 4828 26181 4834
rect 26215 4833 26217 4862
rect 26251 4862 26319 4867
rect 26251 4833 26253 4862
rect 26287 4858 26319 4862
rect 26215 4828 26253 4833
rect 26149 4824 26285 4828
rect 26149 4799 26319 4824
rect 26183 4798 26319 4799
rect 26183 4789 26217 4798
rect 26149 4755 26181 4765
rect 26215 4764 26217 4789
rect 26251 4790 26319 4798
rect 26251 4789 26285 4790
rect 26251 4764 26253 4789
rect 26215 4755 26253 4764
rect 26287 4755 26319 4756
rect 26149 4730 26319 4755
rect 26183 4729 26319 4730
rect 26183 4716 26217 4729
rect 26149 4682 26181 4696
rect 26215 4695 26217 4716
rect 26251 4722 26319 4729
rect 26251 4716 26285 4722
rect 26251 4695 26253 4716
rect 26215 4682 26253 4695
rect 26287 4682 26319 4688
rect 26149 4661 26319 4682
rect 26183 4660 26319 4661
rect 26183 4643 26217 4660
rect 26149 4609 26181 4627
rect 26215 4626 26217 4643
rect 26251 4654 26319 4660
rect 26251 4643 26285 4654
rect 26251 4626 26253 4643
rect 26215 4609 26253 4626
rect 26287 4609 26319 4620
rect 26149 4592 26319 4609
rect 26183 4591 26319 4592
rect 26183 4570 26217 4591
rect 26149 4536 26181 4558
rect 26215 4557 26217 4570
rect 26251 4586 26319 4591
rect 26251 4570 26285 4586
rect 26251 4557 26253 4570
rect 26215 4536 26253 4557
rect 26287 4536 26319 4552
rect 26149 4523 26319 4536
rect 26183 4522 26319 4523
rect 26183 4497 26217 4522
rect 26149 4463 26181 4489
rect 26215 4488 26217 4497
rect 26251 4518 26319 4522
rect 26251 4497 26285 4518
rect 26251 4488 26253 4497
rect 26215 4463 26253 4488
rect 26287 4463 26319 4484
rect 26149 4454 26319 4463
rect 26183 4453 26319 4454
rect 26183 4424 26217 4453
rect 26149 4390 26181 4420
rect 26215 4419 26217 4424
rect 26251 4450 26319 4453
rect 26251 4424 26285 4450
rect 26251 4419 26253 4424
rect 26215 4390 26253 4419
rect 26287 4390 26319 4416
rect 26149 4385 26319 4390
rect 26183 4384 26319 4385
rect 26183 4351 26217 4384
rect 26251 4382 26319 4384
rect 26251 4351 26285 4382
rect 26149 4316 26181 4351
rect 26149 4247 26181 4282
rect 26287 4314 26319 4348
rect 26287 4246 26319 4280
rect 26149 4178 26181 4213
rect 26149 40 26181 64
rect 25234 22 25938 39
rect 25234 -12 25268 22
rect 25302 -12 25336 22
rect 25370 -12 25404 22
rect 25438 -12 25472 22
rect 25506 -12 25540 22
rect 25574 -12 25608 22
rect 25642 -12 25676 22
rect 25710 -12 25744 22
rect 25778 -12 25812 22
rect 25846 -12 25880 22
rect 25914 -12 25938 22
rect 25234 -36 25938 -12
rect 26287 40 26319 64
<< viali >>
rect -265 6732 -231 6766
rect -192 6732 -158 6766
rect -119 6732 -85 6766
rect -46 6732 -12 6766
rect 27 6732 61 6766
rect 100 6732 134 6766
rect 173 6732 207 6766
rect 246 6732 280 6766
rect 319 6732 353 6766
rect 392 6732 426 6766
rect 465 6732 499 6766
rect 538 6732 572 6766
rect 611 6732 645 6766
rect 684 6732 718 6766
rect 757 6732 791 6766
rect 830 6732 864 6766
rect 903 6732 937 6766
rect 976 6732 1010 6766
rect 1049 6732 1083 6766
rect 1122 6764 1152 6766
rect 1152 6764 1156 6766
rect 1195 6764 1221 6766
rect 1221 6764 1229 6766
rect 1122 6732 1156 6764
rect 1195 6732 1229 6764
rect 1268 6764 1289 6766
rect 1289 6764 1302 6766
rect 1341 6764 1358 6766
rect 1358 6764 1375 6766
rect 1413 6764 1427 6766
rect 1427 6764 1447 6766
rect 1485 6764 1496 6766
rect 1496 6764 1519 6766
rect 1557 6764 1565 6766
rect 1565 6764 1591 6766
rect 1629 6764 1634 6766
rect 1634 6764 1663 6766
rect 1701 6764 1703 6766
rect 1703 6764 1735 6766
rect 1773 6764 1806 6766
rect 1806 6764 1807 6766
rect 1845 6764 1875 6766
rect 1875 6764 1879 6766
rect 1917 6764 1944 6766
rect 1944 6764 1951 6766
rect 1989 6764 2012 6766
rect 2012 6764 2023 6766
rect 1268 6732 1302 6764
rect 1341 6732 1375 6764
rect 1413 6732 1447 6764
rect 1485 6732 1519 6764
rect 1557 6732 1591 6764
rect 1629 6732 1663 6764
rect 1701 6732 1735 6764
rect 1773 6732 1807 6764
rect 1845 6732 1879 6764
rect 1917 6732 1951 6764
rect 1989 6732 2023 6764
rect 2061 6732 2095 6766
rect 2133 6732 2148 6766
rect 2148 6732 2167 6766
rect 2205 6764 2217 6766
rect 2217 6764 2239 6766
rect 2277 6764 2286 6766
rect 2286 6764 2311 6766
rect 2349 6764 2355 6766
rect 2355 6764 2383 6766
rect 2421 6764 2424 6766
rect 2424 6764 2455 6766
rect 2205 6732 2239 6764
rect 2277 6732 2311 6764
rect 2349 6732 2383 6764
rect 2421 6732 2455 6764
rect 2493 6732 2527 6766
rect 2565 6764 2597 6766
rect 2597 6764 2599 6766
rect 2637 6764 2666 6766
rect 2666 6764 2671 6766
rect 2709 6764 2735 6766
rect 2735 6764 2743 6766
rect 2781 6764 2804 6766
rect 2804 6764 2815 6766
rect 2853 6764 2873 6766
rect 2873 6764 2887 6766
rect 2925 6764 2942 6766
rect 2942 6764 2959 6766
rect 2997 6764 3011 6766
rect 3011 6764 3031 6766
rect 3069 6764 3080 6766
rect 3080 6764 3103 6766
rect 3141 6764 3149 6766
rect 3149 6764 3175 6766
rect 3213 6764 3218 6766
rect 3218 6764 3247 6766
rect 3285 6764 3287 6766
rect 3287 6764 3319 6766
rect 3357 6764 3390 6766
rect 3390 6764 3391 6766
rect 3429 6764 3459 6766
rect 3459 6764 3463 6766
rect 3501 6764 3528 6766
rect 3528 6764 3535 6766
rect 3573 6764 3597 6766
rect 3597 6764 3607 6766
rect 3645 6764 3666 6766
rect 3666 6764 3679 6766
rect 3717 6764 3735 6766
rect 3735 6764 3751 6766
rect 3789 6764 3804 6766
rect 3804 6764 3823 6766
rect 3861 6764 3873 6766
rect 3873 6764 3895 6766
rect 3933 6764 3942 6766
rect 3942 6764 3967 6766
rect 4005 6764 4011 6766
rect 4011 6764 4039 6766
rect 4077 6764 4080 6766
rect 4080 6764 4111 6766
rect 4149 6764 4184 6766
rect 4184 6764 4218 6766
rect 4218 6764 4253 6766
rect 4253 6764 4287 6766
rect 4287 6764 4322 6766
rect 4322 6764 4356 6766
rect 4356 6764 4391 6766
rect 4391 6764 4425 6766
rect 4425 6764 4460 6766
rect 4460 6764 4494 6766
rect 4494 6764 4529 6766
rect 4529 6764 4563 6766
rect 4563 6764 4598 6766
rect 4598 6764 4632 6766
rect 4632 6764 4667 6766
rect 4667 6764 4701 6766
rect 4701 6764 4736 6766
rect 4736 6764 4770 6766
rect 4770 6764 4805 6766
rect 4805 6764 4839 6766
rect 4839 6764 4874 6766
rect 4874 6764 4908 6766
rect 4908 6764 4943 6766
rect 4943 6764 4977 6766
rect 4977 6764 5012 6766
rect 5012 6764 5046 6766
rect 5046 6764 5081 6766
rect 5081 6764 5115 6766
rect 5115 6764 5150 6766
rect 5150 6764 5184 6766
rect 5184 6764 5219 6766
rect 5219 6764 5253 6766
rect 5253 6764 5288 6766
rect 5288 6764 5322 6766
rect 5322 6764 5357 6766
rect 5357 6764 5391 6766
rect 5391 6764 5426 6766
rect 5426 6764 5460 6766
rect 5460 6764 5495 6766
rect 5495 6764 5529 6766
rect 5529 6764 5564 6766
rect 5564 6764 5598 6766
rect 5598 6764 5633 6766
rect 5633 6764 5667 6766
rect 5667 6764 5702 6766
rect 5702 6764 5736 6766
rect 5736 6764 5771 6766
rect 5771 6764 5805 6766
rect 5805 6764 5840 6766
rect 5840 6764 5874 6766
rect 5874 6764 5909 6766
rect 5909 6764 5943 6766
rect 5943 6764 5978 6766
rect 5978 6764 6012 6766
rect 6012 6764 6047 6766
rect 6047 6764 6081 6766
rect 6081 6764 6116 6766
rect 6116 6764 6150 6766
rect 6150 6764 6185 6766
rect 6185 6764 6219 6766
rect 6219 6764 6254 6766
rect 6254 6764 6288 6766
rect 6288 6764 6323 6766
rect 6323 6764 6357 6766
rect 6357 6764 6392 6766
rect 6392 6764 6426 6766
rect 6426 6764 6461 6766
rect 6461 6764 6495 6766
rect 6495 6764 6530 6766
rect 6530 6764 6564 6766
rect 6564 6764 6599 6766
rect 2565 6732 2599 6764
rect 2637 6732 2671 6764
rect 2709 6732 2743 6764
rect 2781 6732 2815 6764
rect 2853 6732 2887 6764
rect 2925 6732 2959 6764
rect 2997 6732 3031 6764
rect 3069 6732 3103 6764
rect 3141 6732 3175 6764
rect 3213 6732 3247 6764
rect 3285 6732 3319 6764
rect 3357 6732 3391 6764
rect 3429 6732 3463 6764
rect 3501 6732 3535 6764
rect 3573 6732 3607 6764
rect 3645 6732 3679 6764
rect 3717 6732 3751 6764
rect 3789 6732 3823 6764
rect 3861 6732 3895 6764
rect 3933 6732 3967 6764
rect 4005 6732 4039 6764
rect 4077 6732 4111 6764
rect 4149 6730 6599 6764
rect 6599 6730 26143 6766
rect 4149 6696 4184 6730
rect 4184 6696 4218 6730
rect 4218 6696 4253 6730
rect -231 6660 -197 6694
rect -158 6660 -124 6694
rect -85 6660 -51 6694
rect -12 6660 22 6694
rect 61 6660 95 6694
rect 134 6660 168 6694
rect 207 6660 241 6694
rect 280 6660 314 6694
rect 353 6660 387 6694
rect 426 6660 460 6694
rect 499 6660 533 6694
rect 572 6660 606 6694
rect 645 6660 679 6694
rect 718 6660 752 6694
rect 791 6660 825 6694
rect 864 6660 898 6694
rect 937 6660 971 6694
rect 1010 6660 1044 6694
rect 1083 6660 1117 6694
rect 1156 6662 1190 6694
rect 1229 6692 1263 6694
rect -303 6628 -197 6656
rect 1156 6660 1187 6662
rect 1187 6660 1190 6662
rect 1229 6660 1255 6692
rect 1255 6660 1263 6692
rect 1302 6661 1336 6694
rect 1375 6662 1409 6694
rect 1448 6662 1482 6694
rect 1521 6662 1555 6694
rect 1594 6662 1628 6694
rect 1667 6662 1701 6694
rect 1740 6662 1774 6694
rect 1813 6662 1847 6694
rect 1886 6662 1920 6694
rect 1959 6662 1993 6694
rect 1302 6660 1323 6661
rect 1323 6660 1336 6661
rect 1375 6660 1391 6662
rect 1391 6660 1409 6662
rect 1448 6660 1464 6662
rect 1464 6660 1482 6662
rect 1521 6660 1537 6662
rect 1537 6660 1555 6662
rect 1594 6660 1610 6662
rect 1610 6660 1628 6662
rect 1667 6660 1683 6662
rect 1683 6660 1701 6662
rect 1740 6660 1756 6662
rect 1756 6660 1774 6662
rect 1813 6660 1829 6662
rect 1829 6660 1847 6662
rect 1886 6660 1902 6662
rect 1902 6660 1920 6662
rect 1959 6660 1974 6662
rect 1974 6660 1993 6662
rect 2032 6660 2046 6694
rect 2046 6660 2066 6694
rect 2105 6660 2139 6694
rect 2178 6662 2212 6694
rect 2251 6662 2285 6694
rect 2324 6662 2358 6694
rect 2397 6662 2431 6694
rect 2470 6662 2504 6694
rect 2543 6662 2577 6694
rect 2616 6662 2650 6694
rect 2689 6662 2723 6694
rect 2762 6662 2796 6694
rect 2835 6662 2869 6694
rect 2178 6660 2183 6662
rect 2183 6660 2212 6662
rect 2251 6660 2252 6662
rect 2252 6660 2285 6662
rect -303 6560 -233 6628
rect -233 6560 -197 6628
rect -303 6525 -197 6560
rect -303 6491 -301 6525
rect -301 6491 -267 6525
rect -267 6491 -233 6525
rect -233 6491 -197 6525
rect -303 6456 -197 6491
rect 2324 6660 2355 6662
rect 2355 6660 2358 6662
rect 2397 6660 2424 6662
rect 2424 6660 2431 6662
rect 2470 6660 2493 6662
rect 2493 6660 2504 6662
rect 2543 6660 2562 6662
rect 2562 6660 2577 6662
rect 2616 6660 2631 6662
rect 2631 6660 2650 6662
rect 2689 6660 2700 6662
rect 2700 6660 2723 6662
rect 2762 6660 2769 6662
rect 2769 6660 2796 6662
rect 2835 6660 2838 6662
rect 2838 6660 2869 6662
rect 2908 6660 2942 6694
rect 2981 6662 3015 6694
rect 3054 6662 3088 6694
rect 3127 6662 3161 6694
rect 3200 6662 3234 6694
rect 3273 6662 3307 6694
rect 3346 6662 3380 6694
rect 3419 6662 3453 6694
rect 3492 6662 3526 6694
rect 3565 6662 3599 6694
rect 3638 6662 3672 6694
rect 3711 6662 3745 6694
rect 3784 6662 3818 6694
rect 3857 6662 3891 6694
rect 3930 6662 3964 6694
rect 4003 6662 4037 6694
rect 4076 6662 4110 6694
rect 4149 6662 4253 6696
rect 2981 6660 3011 6662
rect 3011 6660 3015 6662
rect 3054 6660 3080 6662
rect 3080 6660 3088 6662
rect 3127 6660 3149 6662
rect 3149 6660 3161 6662
rect 3200 6660 3218 6662
rect 3218 6660 3234 6662
rect 3273 6660 3287 6662
rect 3287 6660 3307 6662
rect 3346 6660 3356 6662
rect 3356 6660 3380 6662
rect 3419 6660 3425 6662
rect 3425 6660 3453 6662
rect 3492 6660 3494 6662
rect 3494 6660 3526 6662
rect 3565 6660 3597 6662
rect 3597 6660 3599 6662
rect 3638 6660 3666 6662
rect 3666 6660 3672 6662
rect 3711 6660 3735 6662
rect 3735 6660 3745 6662
rect 3784 6660 3804 6662
rect 3804 6660 3818 6662
rect 3857 6660 3873 6662
rect 3873 6660 3891 6662
rect 3930 6660 3942 6662
rect 3942 6660 3964 6662
rect 4003 6660 4011 6662
rect 4011 6660 4037 6662
rect 4076 6660 4080 6662
rect 4080 6660 4110 6662
rect 4149 6660 4184 6662
rect 4184 6660 4218 6662
rect 4218 6660 4253 6662
rect 4253 6660 26143 6730
rect 26181 6726 26215 6760
rect 26253 6730 26285 6760
rect 26285 6730 26287 6760
rect 26253 6726 26287 6730
rect 26181 6653 26183 6687
rect 26183 6653 26215 6687
rect 26253 6661 26285 6687
rect 26285 6661 26287 6687
rect 1287 6588 1289 6622
rect 1289 6592 1393 6622
rect 1289 6588 1323 6592
rect 1287 6558 1323 6588
rect 1323 6558 1357 6592
rect 1357 6558 1391 6592
rect 1391 6558 1393 6592
rect 1287 6552 1393 6558
rect 1287 6518 1289 6552
rect 1289 6523 1393 6552
rect 1289 6518 1323 6523
rect -9 6464 25 6490
rect 66 6464 100 6490
rect 141 6464 175 6490
rect 216 6464 250 6490
rect 291 6464 325 6490
rect 365 6464 399 6490
rect 439 6464 473 6490
rect -303 6422 -301 6456
rect -301 6422 -267 6456
rect -267 6422 -233 6456
rect -233 6422 -197 6456
rect -303 6387 -197 6422
rect -303 6353 -301 6387
rect -301 6353 -267 6387
rect -267 6353 -233 6387
rect -233 6353 -197 6387
rect -303 6318 -197 6353
rect -303 6284 -301 6318
rect -301 6284 -267 6318
rect -267 6284 -233 6318
rect -233 6284 -197 6318
rect -303 6249 -197 6284
rect -303 6215 -301 6249
rect -301 6215 -267 6249
rect -267 6215 -233 6249
rect -233 6215 -197 6249
rect -303 6180 -197 6215
rect -303 6146 -301 6180
rect -301 6146 -267 6180
rect -267 6146 -233 6180
rect -233 6146 -197 6180
rect -303 6111 -197 6146
rect -303 6077 -301 6111
rect -301 6077 -267 6111
rect -267 6077 -233 6111
rect -233 6077 -197 6111
rect -303 6042 -197 6077
rect -303 6008 -301 6042
rect -301 6008 -267 6042
rect -267 6008 -233 6042
rect -233 6008 -197 6042
rect -303 5973 -197 6008
rect -303 5939 -301 5973
rect -301 5939 -267 5973
rect -267 5939 -233 5973
rect -233 5939 -197 5973
rect -303 5904 -197 5939
rect -303 5870 -301 5904
rect -301 5870 -267 5904
rect -267 5870 -233 5904
rect -233 5870 -197 5904
rect -303 5835 -197 5870
rect -303 5801 -301 5835
rect -301 5801 -267 5835
rect -267 5801 -233 5835
rect -233 5801 -197 5835
rect -303 5766 -197 5801
rect -303 5732 -301 5766
rect -301 5732 -267 5766
rect -267 5732 -233 5766
rect -233 5732 -197 5766
rect -303 5697 -197 5732
rect -303 5663 -301 5697
rect -301 5663 -267 5697
rect -267 5663 -233 5697
rect -233 5663 -197 5697
rect -303 5628 -197 5663
rect -303 5594 -301 5628
rect -301 5594 -267 5628
rect -267 5594 -233 5628
rect -233 5594 -197 5628
rect -303 5558 -197 5594
rect -303 5524 -301 5558
rect -301 5524 -267 5558
rect -267 5524 -233 5558
rect -233 5524 -197 5558
rect -303 5488 -197 5524
rect -303 5454 -301 5488
rect -301 5454 -267 5488
rect -267 5454 -233 5488
rect -233 5454 -197 5488
rect -303 5418 -197 5454
rect -303 5384 -301 5418
rect -301 5384 -267 5418
rect -267 5384 -233 5418
rect -233 5384 -197 5418
rect -303 5348 -197 5384
rect -303 5314 -301 5348
rect -301 5314 -267 5348
rect -267 5314 -233 5348
rect -233 5314 -197 5348
rect -303 5278 -197 5314
rect -303 5244 -301 5278
rect -301 5244 -267 5278
rect -267 5244 -233 5278
rect -233 5244 -197 5278
rect -303 5208 -197 5244
rect -303 5174 -301 5208
rect -301 5174 -267 5208
rect -267 5174 -233 5208
rect -233 5174 -197 5208
rect -303 5138 -197 5174
rect -303 5104 -301 5138
rect -301 5104 -267 5138
rect -267 5104 -233 5138
rect -233 5104 -197 5138
rect -303 5068 -197 5104
rect -9 6456 11 6464
rect 11 6456 25 6464
rect 66 6456 83 6464
rect 83 6456 100 6464
rect 141 6456 155 6464
rect 155 6456 175 6464
rect 216 6456 227 6464
rect 227 6456 250 6464
rect 291 6456 298 6464
rect 298 6456 325 6464
rect 365 6456 369 6464
rect 369 6456 399 6464
rect 439 6456 440 6464
rect 440 6456 473 6464
rect 513 6456 547 6490
rect 587 6464 621 6490
rect 661 6464 695 6490
rect 735 6464 769 6490
rect 809 6464 843 6490
rect 883 6464 917 6490
rect 957 6464 991 6490
rect 1031 6464 1065 6490
rect 1287 6489 1323 6518
rect 1323 6489 1357 6523
rect 1357 6522 1393 6523
rect 1357 6489 1391 6522
rect 1287 6488 1391 6489
rect 1391 6488 1393 6522
rect 1287 6482 1393 6488
rect 587 6456 619 6464
rect 619 6456 621 6464
rect 661 6456 690 6464
rect 690 6456 695 6464
rect 735 6456 761 6464
rect 761 6456 769 6464
rect 809 6456 832 6464
rect 832 6456 843 6464
rect 883 6456 903 6464
rect 903 6456 917 6464
rect 957 6456 974 6464
rect 974 6456 991 6464
rect 1031 6456 1045 6464
rect 1045 6456 1065 6464
rect -9 6384 25 6418
rect 66 6384 100 6418
rect 141 6384 175 6418
rect 216 6384 250 6418
rect 291 6384 325 6418
rect 365 6384 399 6418
rect 439 6384 473 6418
rect 513 6384 547 6418
rect 587 6384 621 6418
rect 661 6384 695 6418
rect 735 6384 769 6418
rect 809 6384 843 6418
rect 883 6384 917 6418
rect 957 6384 991 6418
rect 1031 6384 1065 6418
rect 23 6312 57 6346
rect 98 6344 126 6346
rect 126 6344 132 6346
rect 173 6344 195 6346
rect 195 6344 207 6346
rect 248 6344 265 6346
rect 265 6344 282 6346
rect 323 6344 335 6346
rect 335 6344 357 6346
rect 398 6344 405 6346
rect 405 6344 432 6346
rect 473 6344 475 6346
rect 475 6344 507 6346
rect 548 6344 579 6346
rect 579 6344 582 6346
rect 623 6344 649 6346
rect 649 6344 657 6346
rect 698 6344 719 6346
rect 719 6344 732 6346
rect 773 6344 789 6346
rect 789 6344 807 6346
rect 848 6344 859 6346
rect 859 6344 882 6346
rect 923 6344 929 6346
rect 929 6344 957 6346
rect 98 6312 132 6344
rect 173 6312 207 6344
rect 248 6312 282 6344
rect 323 6312 357 6344
rect 398 6312 432 6344
rect 473 6312 507 6344
rect 548 6312 582 6344
rect 623 6312 657 6344
rect 698 6312 732 6344
rect 773 6312 807 6344
rect 848 6312 882 6344
rect 923 6312 957 6344
rect 1037 6274 1071 6308
rect 57 6242 91 6274
rect 133 6242 167 6274
rect 209 6242 243 6274
rect 285 6242 319 6274
rect 361 6242 395 6274
rect 437 6242 471 6274
rect 513 6242 547 6274
rect 589 6242 623 6274
rect 665 6242 699 6274
rect 740 6242 774 6274
rect 815 6242 849 6274
rect 890 6242 924 6274
rect 965 6242 999 6274
rect 57 6240 89 6242
rect 89 6240 91 6242
rect 133 6240 159 6242
rect 159 6240 167 6242
rect 209 6240 229 6242
rect 229 6240 243 6242
rect 285 6240 299 6242
rect 299 6240 319 6242
rect 361 6240 369 6242
rect 369 6240 395 6242
rect 437 6240 439 6242
rect 439 6240 471 6242
rect -15 6202 19 6234
rect 513 6240 543 6242
rect 543 6240 547 6242
rect 589 6240 613 6242
rect 613 6240 623 6242
rect 665 6240 683 6242
rect 683 6240 699 6242
rect 740 6240 754 6242
rect 754 6240 774 6242
rect 815 6240 825 6242
rect 825 6240 849 6242
rect 890 6240 896 6242
rect 896 6240 924 6242
rect 965 6240 967 6242
rect 967 6240 999 6242
rect -15 6200 -13 6202
rect -13 6200 19 6202
rect 57 6168 91 6198
rect 57 6164 89 6168
rect 89 6164 91 6168
rect -15 6132 19 6161
rect -15 6127 -13 6132
rect -13 6127 19 6132
rect 57 6094 91 6122
rect 1037 6202 1071 6233
rect 1037 6199 1069 6202
rect 1069 6199 1071 6202
rect 965 6172 999 6198
rect 965 6164 967 6172
rect 967 6164 999 6172
rect 1037 6132 1071 6158
rect 1037 6124 1069 6132
rect 1069 6124 1071 6132
rect -15 6062 19 6088
rect -15 6054 -13 6062
rect -13 6054 19 6062
rect 57 6088 89 6094
rect 89 6088 91 6094
rect 356 6080 390 6114
rect 428 6080 462 6114
rect 500 6080 534 6114
rect 572 6080 606 6114
rect 644 6080 678 6114
rect 716 6080 750 6114
rect 965 6102 999 6122
rect 965 6088 967 6102
rect 967 6088 999 6102
rect 57 6020 91 6046
rect -15 5992 19 6015
rect -15 5981 -13 5992
rect -13 5981 19 5992
rect 57 6012 89 6020
rect 89 6012 91 6020
rect 57 5946 91 5970
rect -15 5922 19 5942
rect -15 5908 -13 5922
rect -13 5908 19 5922
rect 57 5936 89 5946
rect 89 5936 91 5946
rect 57 5873 91 5894
rect -15 5852 19 5869
rect -15 5835 -13 5852
rect -13 5835 19 5852
rect 57 5860 89 5873
rect 89 5860 91 5873
rect 57 5800 91 5818
rect -15 5782 19 5795
rect -15 5761 -13 5782
rect -13 5761 19 5782
rect 57 5784 89 5800
rect 89 5784 91 5800
rect 57 5727 91 5742
rect -15 5712 19 5721
rect -15 5687 -13 5712
rect -13 5687 19 5712
rect 57 5708 89 5727
rect 89 5708 91 5727
rect 57 5654 91 5666
rect -15 5642 19 5647
rect -15 5613 -13 5642
rect -13 5613 19 5642
rect 57 5632 89 5654
rect 89 5632 91 5654
rect 57 5581 91 5590
rect -15 5572 19 5573
rect -15 5539 -13 5572
rect -13 5539 19 5572
rect 57 5556 89 5581
rect 89 5556 91 5581
rect 57 5508 91 5514
rect -15 5468 -13 5499
rect -13 5468 19 5499
rect 57 5480 89 5508
rect 89 5480 91 5508
rect -15 5465 19 5468
rect 57 5435 91 5437
rect -15 5398 -13 5425
rect -13 5398 19 5425
rect 57 5403 89 5435
rect 89 5403 91 5435
rect -15 5391 19 5398
rect 1037 6062 1071 6083
rect 1037 6049 1069 6062
rect 1069 6049 1071 6062
rect 965 6032 999 6046
rect 965 6012 967 6032
rect 967 6012 999 6032
rect 1037 5992 1071 6008
rect 1037 5974 1069 5992
rect 1069 5974 1071 5992
rect 965 5962 999 5970
rect 356 5924 390 5958
rect 428 5924 462 5958
rect 500 5924 534 5958
rect 572 5924 606 5958
rect 644 5924 678 5958
rect 716 5924 750 5958
rect 965 5936 967 5962
rect 967 5936 999 5962
rect 1037 5922 1071 5933
rect 1037 5899 1069 5922
rect 1069 5899 1071 5922
rect 965 5891 999 5895
rect 965 5861 967 5891
rect 967 5861 999 5891
rect 1037 5852 1071 5858
rect 1037 5824 1069 5852
rect 1069 5824 1071 5852
rect 512 5768 546 5802
rect 584 5768 618 5802
rect 656 5768 690 5802
rect 728 5768 762 5802
rect 965 5786 967 5820
rect 967 5786 999 5820
rect 1037 5782 1071 5783
rect 965 5715 967 5745
rect 967 5715 999 5745
rect 1037 5749 1069 5782
rect 1069 5749 1071 5782
rect 965 5711 999 5715
rect 516 5658 550 5692
rect 588 5658 622 5692
rect 660 5658 694 5692
rect 732 5658 766 5692
rect 965 5644 967 5670
rect 967 5644 999 5670
rect 1037 5678 1069 5708
rect 1069 5678 1071 5708
rect 1037 5674 1071 5678
rect 965 5636 999 5644
rect 965 5573 967 5595
rect 967 5573 999 5595
rect 1037 5608 1069 5633
rect 1069 5608 1071 5633
rect 1037 5599 1071 5608
rect 965 5561 999 5573
rect 516 5502 550 5536
rect 588 5502 622 5536
rect 660 5502 694 5536
rect 732 5502 766 5536
rect 965 5502 967 5520
rect 967 5502 999 5520
rect 1037 5538 1069 5558
rect 1069 5538 1071 5558
rect 1037 5524 1071 5538
rect 965 5486 999 5502
rect 1037 5468 1069 5484
rect 1069 5468 1071 5484
rect 965 5431 967 5445
rect 967 5431 999 5445
rect 1037 5450 1071 5468
rect 965 5411 999 5431
rect 1037 5398 1069 5410
rect 1069 5398 1071 5410
rect -15 5328 -13 5351
rect -13 5328 19 5351
rect 57 5328 89 5360
rect 89 5328 91 5360
rect 596 5346 630 5380
rect 668 5346 702 5380
rect 740 5346 774 5380
rect 965 5360 967 5370
rect 967 5360 999 5370
rect 1037 5376 1071 5398
rect -15 5317 19 5328
rect 57 5326 91 5328
rect -15 5252 19 5277
rect 57 5252 91 5283
rect 965 5336 999 5360
rect 1037 5328 1069 5336
rect 1069 5328 1071 5336
rect 965 5289 967 5295
rect 967 5289 999 5295
rect 1037 5302 1071 5328
rect 965 5261 999 5289
rect 1037 5258 1069 5262
rect 1069 5258 1071 5262
rect -15 5243 11 5252
rect 11 5243 19 5252
rect 57 5249 80 5252
rect 80 5249 91 5252
rect 1037 5228 1071 5258
rect -15 5184 19 5203
rect 57 5184 91 5206
rect 715 5186 749 5220
rect 798 5186 832 5220
rect 881 5186 915 5220
rect 965 5186 967 5220
rect 967 5186 999 5220
rect -15 5169 11 5184
rect 11 5169 19 5184
rect 57 5172 80 5184
rect 80 5172 91 5184
rect -15 5116 19 5129
rect 57 5116 91 5129
rect 715 5116 749 5148
rect 809 5116 843 5148
rect 904 5116 938 5148
rect -15 5095 11 5116
rect 11 5095 19 5116
rect 57 5095 82 5116
rect 82 5095 91 5116
rect 715 5114 717 5116
rect 717 5114 749 5116
rect 809 5114 823 5116
rect 823 5114 843 5116
rect 904 5114 927 5116
rect 927 5114 938 5116
rect 999 5114 1033 5148
rect 1287 6448 1289 6482
rect 1289 6454 1393 6482
rect 1289 6448 1323 6454
rect 1287 6420 1323 6448
rect 1323 6420 1357 6454
rect 1357 6452 1393 6454
rect 26253 6653 26287 6661
rect 26181 6593 26215 6614
rect 26181 6580 26183 6593
rect 26183 6580 26215 6593
rect 26253 6592 26285 6614
rect 26285 6592 26287 6614
rect 26253 6580 26287 6592
rect 26181 6524 26215 6541
rect 26181 6507 26183 6524
rect 26183 6507 26215 6524
rect 26253 6524 26285 6541
rect 26285 6524 26287 6541
rect 26253 6507 26287 6524
rect 1357 6420 1391 6452
rect 1287 6418 1391 6420
rect 1391 6418 1393 6452
rect 1287 6412 1393 6418
rect 1287 6378 1289 6412
rect 1289 6385 1393 6412
rect 1289 6378 1323 6385
rect 1287 6351 1323 6378
rect 1323 6351 1357 6385
rect 1357 6382 1393 6385
rect 1357 6351 1391 6382
rect 1287 6348 1391 6351
rect 1391 6348 1393 6382
rect 1287 6342 1393 6348
rect 1287 6308 1289 6342
rect 1289 6316 1393 6342
rect 1289 6308 1323 6316
rect 1287 6282 1323 6308
rect 1323 6282 1357 6316
rect 1357 6312 1393 6316
rect 1357 6282 1391 6312
rect 1287 6278 1391 6282
rect 1391 6278 1393 6312
rect 1287 6272 1393 6278
rect 1287 6238 1289 6272
rect 1289 6247 1393 6272
rect 1289 6238 1323 6247
rect 1287 6213 1323 6238
rect 1323 6213 1357 6247
rect 1357 6242 1393 6247
rect 1357 6213 1391 6242
rect 1287 6208 1391 6213
rect 1391 6208 1393 6242
rect 1287 6202 1393 6208
rect 1287 6168 1289 6202
rect 1289 6178 1393 6202
rect 1289 6168 1323 6178
rect 1287 6144 1323 6168
rect 1323 6144 1357 6178
rect 1357 6172 1393 6178
rect 1357 6144 1391 6172
rect 1287 6138 1391 6144
rect 1391 6138 1393 6172
rect 1287 6132 1393 6138
rect 1287 6098 1289 6132
rect 1289 6109 1393 6132
rect 1289 6098 1323 6109
rect 1287 6075 1323 6098
rect 1323 6075 1357 6109
rect 1357 6102 1393 6109
rect 1357 6075 1391 6102
rect 1287 6068 1391 6075
rect 1391 6068 1393 6102
rect 1287 6062 1393 6068
rect 1287 6028 1289 6062
rect 1289 6040 1393 6062
rect 1289 6028 1323 6040
rect 1287 6006 1323 6028
rect 1323 6006 1357 6040
rect 1357 6032 1393 6040
rect 1357 6006 1391 6032
rect 1287 5998 1391 6006
rect 1391 5998 1393 6032
rect 1287 5992 1393 5998
rect 1287 5958 1289 5992
rect 1289 5971 1393 5992
rect 1289 5958 1323 5971
rect 1287 5937 1323 5958
rect 1323 5937 1357 5971
rect 1357 5962 1393 5971
rect 1357 5937 1391 5962
rect 1287 5928 1391 5937
rect 1391 5928 1393 5962
rect 1287 5922 1393 5928
rect 1287 5888 1289 5922
rect 1289 5902 1393 5922
rect 1289 5888 1323 5902
rect 1287 5868 1323 5888
rect 1323 5868 1357 5902
rect 1357 5892 1393 5902
rect 1357 5868 1391 5892
rect 1287 5858 1391 5868
rect 1391 5858 1393 5892
rect 1287 5852 1393 5858
rect 1287 5818 1289 5852
rect 1289 5833 1393 5852
rect 1289 5818 1323 5833
rect 1287 5799 1323 5818
rect 1323 5799 1357 5833
rect 1357 5822 1393 5833
rect 1357 5799 1391 5822
rect 1287 5788 1391 5799
rect 1391 5788 1393 5822
rect 1287 5782 1393 5788
rect 1287 5748 1289 5782
rect 1289 5764 1393 5782
rect 1289 5748 1323 5764
rect 1287 5730 1323 5748
rect 1323 5730 1357 5764
rect 1357 5751 1393 5764
rect 1357 5730 1391 5751
rect 1287 5717 1391 5730
rect 1391 5717 1393 5751
rect 1287 5711 1393 5717
rect 1287 5677 1289 5711
rect 1289 5695 1393 5711
rect 1289 5677 1323 5695
rect 1287 5661 1323 5677
rect 1323 5661 1357 5695
rect 1357 5680 1393 5695
rect 1357 5661 1391 5680
rect 1287 5646 1391 5661
rect 1391 5646 1393 5680
rect 1287 5640 1393 5646
rect 1287 5606 1289 5640
rect 1289 5626 1393 5640
rect 1289 5606 1323 5626
rect 1287 5592 1323 5606
rect 1323 5592 1357 5626
rect 1357 5609 1393 5626
rect 1357 5592 1391 5609
rect 1287 5575 1391 5592
rect 1391 5575 1393 5609
rect 1287 5569 1393 5575
rect 1287 5535 1289 5569
rect 1289 5557 1393 5569
rect 1289 5535 1323 5557
rect 1287 5523 1323 5535
rect 1323 5523 1357 5557
rect 1357 5538 1393 5557
rect 1357 5523 1391 5538
rect 1287 5504 1391 5523
rect 1391 5504 1393 5538
rect 1287 5498 1393 5504
rect 1287 5464 1289 5498
rect 1289 5488 1393 5498
rect 1289 5464 1323 5488
rect 1287 5454 1323 5464
rect 1323 5454 1357 5488
rect 1357 5467 1393 5488
rect 1357 5454 1391 5467
rect 1287 5433 1391 5454
rect 1391 5433 1393 5467
rect 1287 5427 1393 5433
rect 1287 5393 1289 5427
rect 1289 5419 1393 5427
rect 1289 5393 1323 5419
rect 1287 5385 1323 5393
rect 1323 5385 1357 5419
rect 1357 5396 1393 5419
rect 1357 5385 1391 5396
rect 1287 5362 1391 5385
rect 1391 5362 1393 5396
rect 1287 5356 1393 5362
rect 1287 5322 1289 5356
rect 1289 5350 1393 5356
rect 1289 5322 1323 5350
rect 1287 5316 1323 5322
rect 1323 5316 1357 5350
rect 1357 5325 1393 5350
rect 1357 5316 1391 5325
rect 1287 5291 1391 5316
rect 1391 5291 1393 5325
rect 1287 5285 1393 5291
rect 1287 5251 1289 5285
rect 1289 5281 1393 5285
rect 1289 5251 1323 5281
rect 1287 5247 1323 5251
rect 1323 5247 1357 5281
rect 1357 5254 1393 5281
rect 1357 5247 1391 5254
rect 1287 5220 1391 5247
rect 1391 5220 1393 5254
rect 1287 5214 1393 5220
rect 1287 5180 1289 5214
rect 1289 5212 1393 5214
rect 1289 5180 1323 5212
rect 1287 5178 1323 5180
rect 1323 5178 1357 5212
rect 1357 5183 1393 5212
rect 1357 5178 1391 5183
rect 1287 5149 1391 5178
rect 1391 5149 1393 5183
rect 1287 5148 1393 5149
rect -303 5034 -301 5068
rect -301 5034 -267 5068
rect -267 5034 -233 5068
rect -233 5034 -197 5068
rect -303 4998 -197 5034
rect -303 4964 -233 4998
rect -303 4896 -301 4964
rect -301 4930 -233 4964
rect -233 4930 -197 4998
rect 1287 5075 1321 5109
rect 1359 5078 1391 5109
rect 1391 5078 1393 5109
rect 1359 5075 1393 5078
rect 1287 5002 1321 5036
rect 1359 5007 1391 5036
rect 1391 5007 1393 5036
rect 1359 5002 1393 5007
rect 1287 4930 1321 4963
rect 1359 4936 1391 4963
rect 1391 4936 1393 4963
rect -301 4896 -199 4930
rect -199 4896 -197 4930
rect 1287 4929 1289 4930
rect 1289 4929 1321 4930
rect 1359 4929 1393 4936
rect -303 4862 -197 4896
rect -303 4828 -267 4862
rect -267 4828 -233 4862
rect -303 4794 -233 4828
rect -233 4794 -197 4862
rect 1287 4856 1321 4890
rect 1359 4865 1391 4890
rect 1391 4865 1393 4890
rect 1359 4856 1393 4865
rect -303 4284 -197 4794
rect 1804 6460 23006 6473
rect 23045 6460 23079 6473
rect 23118 6460 23152 6473
rect 23191 6460 23225 6473
rect 23264 6460 23298 6473
rect 23337 6460 23371 6473
rect 23410 6460 23444 6473
rect 23483 6460 23517 6473
rect 23556 6460 23590 6473
rect 23629 6460 23663 6473
rect 23702 6460 23736 6473
rect 23775 6460 23809 6473
rect 23848 6460 23882 6473
rect 23921 6460 23955 6473
rect 23994 6460 24028 6473
rect 24067 6460 24101 6473
rect 24140 6460 24174 6473
rect 24213 6460 24247 6473
rect 24286 6460 24320 6473
rect 24359 6460 24393 6473
rect 24432 6460 24466 6473
rect 24505 6460 24539 6473
rect 24578 6460 24612 6473
rect 24651 6460 24685 6473
rect 24724 6460 24758 6473
rect 24797 6460 24831 6473
rect 24870 6460 24904 6473
rect 24943 6460 24977 6473
rect 25016 6460 25050 6473
rect 25089 6460 25123 6473
rect 25162 6460 25196 6473
rect 1804 6426 1808 6460
rect 1808 6426 1842 6460
rect 1842 6426 1877 6460
rect 1877 6426 1911 6460
rect 1911 6426 1946 6460
rect 1946 6426 1980 6460
rect 1980 6426 2015 6460
rect 2015 6426 2049 6460
rect 2049 6426 2084 6460
rect 2084 6426 2118 6460
rect 2118 6426 2153 6460
rect 2153 6426 2187 6460
rect 2187 6426 2222 6460
rect 2222 6426 2256 6460
rect 2256 6426 2291 6460
rect 2291 6426 2325 6460
rect 2325 6426 2360 6460
rect 2360 6426 2394 6460
rect 2394 6426 2429 6460
rect 2429 6426 2463 6460
rect 2463 6426 2498 6460
rect 2498 6426 2532 6460
rect 2532 6426 2567 6460
rect 2567 6426 2601 6460
rect 2601 6426 2636 6460
rect 2636 6426 2670 6460
rect 2670 6426 2705 6460
rect 2705 6426 2739 6460
rect 2739 6426 2774 6460
rect 2774 6426 2808 6460
rect 2808 6426 2843 6460
rect 2843 6426 2877 6460
rect 2877 6426 2912 6460
rect 2912 6426 2946 6460
rect 2946 6426 2981 6460
rect 2981 6426 3015 6460
rect 3015 6426 3050 6460
rect 3050 6426 3084 6460
rect 3084 6426 3119 6460
rect 3119 6426 3153 6460
rect 3153 6426 3188 6460
rect 3188 6426 3222 6460
rect 3222 6426 3257 6460
rect 3257 6426 3291 6460
rect 3291 6426 3326 6460
rect 3326 6426 3360 6460
rect 3360 6426 3395 6460
rect 3395 6426 3429 6460
rect 3429 6426 3464 6460
rect 3464 6426 3498 6460
rect 3498 6426 3533 6460
rect 3533 6426 3567 6460
rect 3567 6426 3602 6460
rect 3602 6426 3636 6460
rect 3636 6426 3671 6460
rect 3671 6426 3705 6460
rect 3705 6426 3740 6460
rect 3740 6426 3774 6460
rect 3774 6426 3809 6460
rect 3809 6426 3843 6460
rect 3843 6426 3878 6460
rect 3878 6426 3912 6460
rect 3912 6426 3947 6460
rect 3947 6426 3981 6460
rect 3981 6426 4016 6460
rect 4016 6426 4050 6460
rect 4050 6426 4085 6460
rect 4085 6426 4119 6460
rect 4119 6426 4154 6460
rect 4154 6426 4188 6460
rect 4188 6426 4223 6460
rect 4223 6426 4257 6460
rect 4257 6426 4292 6460
rect 4292 6426 4326 6460
rect 4326 6426 4361 6460
rect 4361 6426 4395 6460
rect 4395 6426 4430 6460
rect 4430 6426 4464 6460
rect 4464 6426 4499 6460
rect 4499 6426 4533 6460
rect 4533 6426 4568 6460
rect 4568 6426 4602 6460
rect 4602 6426 4637 6460
rect 4637 6426 4671 6460
rect 4671 6426 4706 6460
rect 4706 6426 4740 6460
rect 4740 6426 4775 6460
rect 4775 6426 4809 6460
rect 4809 6426 4844 6460
rect 1804 6392 4844 6426
rect 1804 6367 1808 6392
rect 1808 6367 1842 6392
rect 1842 6367 1877 6392
rect 1877 6367 1911 6392
rect 1911 6367 1946 6392
rect 1946 6367 1980 6392
rect 1980 6367 2015 6392
rect 2015 6367 2049 6392
rect 2049 6367 2084 6392
rect 2084 6367 2118 6392
rect 2118 6367 2153 6392
rect 2153 6367 2187 6392
rect 2187 6367 2222 6392
rect 2222 6367 2256 6392
rect 2256 6367 2291 6392
rect 2291 6367 2325 6392
rect 2325 6367 2360 6392
rect 2360 6367 2394 6392
rect 2394 6367 2429 6392
rect 2429 6367 2463 6392
rect 2463 6367 2498 6392
rect 2498 6367 2532 6392
rect 2532 6367 2567 6392
rect 2567 6367 2601 6392
rect 2601 6367 2636 6392
rect 2636 6367 2670 6392
rect 2670 6367 2705 6392
rect 2705 6367 2739 6392
rect 2739 6367 2774 6392
rect 2774 6367 2808 6392
rect 2808 6367 2843 6392
rect 2843 6367 2877 6392
rect 2877 6367 2912 6392
rect 2912 6367 2946 6392
rect 2946 6367 2981 6392
rect 2981 6367 3015 6392
rect 3015 6367 3050 6392
rect 3050 6367 3084 6392
rect 3084 6367 3119 6392
rect 3119 6367 3153 6392
rect 3153 6367 3188 6392
rect 3188 6367 3222 6392
rect 3222 6367 3257 6392
rect 3257 6367 3291 6392
rect 3291 6367 3326 6392
rect 3326 6367 3360 6392
rect 3360 6367 3395 6392
rect 3395 6367 3429 6392
rect 3429 6367 3464 6392
rect 3464 6367 3498 6392
rect 3498 6367 3533 6392
rect 3533 6367 3567 6392
rect 3567 6367 3602 6392
rect 3602 6367 3636 6392
rect 3636 6367 3671 6392
rect 3671 6367 3705 6392
rect 3705 6367 3740 6392
rect 3740 6367 3774 6392
rect 3774 6367 3809 6392
rect 3809 6367 3843 6392
rect 3843 6367 3878 6392
rect 3878 6367 3912 6392
rect 3912 6367 3947 6392
rect 3947 6367 3981 6392
rect 3981 6367 4016 6392
rect 4016 6367 4050 6392
rect 4050 6367 4085 6392
rect 4085 6367 4119 6392
rect 4119 6367 4154 6392
rect 4154 6367 4188 6392
rect 4188 6367 4223 6392
rect 4223 6367 4257 6392
rect 4257 6367 4292 6392
rect 4292 6367 4326 6392
rect 4326 6367 4361 6392
rect 4361 6367 4395 6392
rect 4395 6367 4430 6392
rect 4430 6367 4464 6392
rect 4464 6367 4499 6392
rect 4499 6367 4533 6392
rect 4533 6367 4568 6392
rect 4568 6367 4602 6392
rect 4602 6367 4637 6392
rect 4637 6367 4671 6392
rect 4671 6367 4706 6392
rect 4706 6367 4740 6392
rect 4740 6367 4775 6392
rect 4775 6367 4809 6392
rect 4809 6367 4844 6392
rect 4844 6367 23006 6460
rect 23045 6439 23079 6460
rect 23118 6439 23152 6460
rect 23191 6439 23225 6460
rect 23264 6439 23298 6460
rect 23337 6439 23371 6460
rect 23410 6439 23444 6460
rect 23483 6439 23517 6460
rect 23556 6439 23590 6460
rect 23629 6439 23663 6460
rect 23702 6439 23736 6460
rect 23775 6439 23809 6460
rect 23848 6439 23882 6460
rect 23921 6439 23955 6460
rect 23994 6439 24028 6460
rect 24067 6439 24101 6460
rect 24140 6439 24174 6460
rect 24213 6439 24247 6460
rect 24286 6439 24320 6460
rect 24359 6439 24393 6460
rect 24432 6439 24466 6460
rect 24505 6439 24539 6460
rect 24578 6439 24612 6460
rect 24651 6439 24685 6460
rect 24724 6439 24758 6460
rect 24797 6439 24831 6460
rect 24870 6439 24904 6460
rect 24943 6439 24977 6460
rect 25016 6439 25050 6460
rect 25089 6439 25123 6460
rect 25162 6439 25196 6460
rect 25235 6444 25269 6473
rect 25308 6444 25342 6473
rect 25381 6444 25415 6473
rect 25454 6444 25488 6473
rect 25527 6444 25561 6473
rect 25235 6439 25268 6444
rect 25268 6439 25269 6444
rect 25308 6439 25342 6444
rect 25381 6439 25415 6444
rect 25454 6439 25488 6444
rect 25527 6439 25561 6444
rect 23045 6367 23079 6401
rect 23118 6367 23152 6401
rect 23191 6367 23225 6401
rect 23264 6367 23298 6401
rect 23337 6367 23371 6401
rect 23410 6367 23444 6401
rect 23483 6367 23517 6401
rect 23556 6367 23590 6401
rect 23629 6367 23663 6401
rect 23702 6367 23736 6401
rect 23775 6367 23809 6401
rect 23848 6367 23882 6401
rect 23921 6367 23955 6401
rect 23994 6367 24028 6401
rect 24067 6367 24101 6401
rect 24140 6367 24174 6401
rect 24213 6367 24247 6401
rect 24286 6367 24320 6401
rect 24359 6367 24393 6401
rect 24432 6367 24466 6401
rect 24505 6367 24539 6401
rect 24578 6367 24612 6401
rect 24651 6367 24685 6401
rect 24724 6367 24758 6401
rect 24797 6367 24831 6401
rect 24870 6367 24904 6401
rect 24943 6367 24977 6401
rect 25016 6367 25050 6401
rect 25089 6367 25123 6401
rect 25162 6367 25196 6401
rect 25235 6367 25268 6401
rect 25268 6367 25269 6401
rect 25308 6367 25342 6401
rect 25381 6367 25415 6401
rect 25454 6367 25488 6401
rect 25527 6367 25561 6401
rect 1609 6290 1635 6294
rect 1635 6290 1643 6294
rect 1681 6290 1704 6294
rect 1704 6290 1715 6294
rect 1609 6260 1643 6290
rect 1681 6260 1715 6290
rect 1609 6188 1643 6220
rect 1681 6188 1715 6222
rect 1609 6186 1635 6188
rect 1635 6186 1643 6188
rect 1609 6120 1643 6146
rect 1681 6120 1715 6149
rect 1609 6112 1635 6120
rect 1635 6112 1643 6120
rect 1681 6115 1704 6120
rect 1704 6115 1715 6120
rect 1609 6052 1643 6072
rect 1681 6052 1715 6076
rect 1609 6038 1635 6052
rect 1635 6038 1643 6052
rect 1681 6042 1704 6052
rect 1704 6042 1715 6052
rect 1609 5984 1643 5998
rect 1681 5984 1715 6003
rect 1609 5964 1635 5984
rect 1635 5964 1643 5984
rect 1681 5969 1704 5984
rect 1704 5969 1715 5984
rect 1609 5916 1643 5924
rect 1681 5916 1715 5930
rect 1609 5890 1635 5916
rect 1635 5890 1643 5916
rect 1681 5896 1704 5916
rect 1704 5896 1715 5916
rect 1609 5848 1643 5850
rect 1681 5848 1715 5857
rect 1609 5816 1635 5848
rect 1635 5816 1643 5848
rect 1681 5823 1704 5848
rect 1704 5823 1715 5848
rect 1681 5780 1715 5784
rect 1609 5746 1635 5776
rect 1635 5746 1643 5776
rect 1681 5750 1704 5780
rect 1704 5750 1715 5780
rect 1609 5742 1643 5746
rect 1609 5678 1611 5702
rect 1611 5678 1643 5702
rect 1681 5678 1715 5711
rect 1609 5668 1643 5678
rect 1681 5677 1715 5678
rect 1609 5604 1643 5627
rect 1681 5604 1715 5638
rect 1609 5593 1611 5604
rect 1611 5593 1643 5604
rect 1609 5533 1643 5552
rect 1681 5542 1713 5565
rect 1713 5542 1715 5565
rect 4723 5548 6421 5654
rect 6421 5548 22973 5654
rect 23350 5620 23384 5654
rect 23423 5620 23457 5654
rect 23496 5620 23530 5654
rect 23569 5620 23603 5654
rect 23642 5620 23676 5654
rect 23715 5620 23749 5654
rect 23788 5620 23822 5654
rect 23861 5620 23895 5654
rect 23934 5620 23968 5654
rect 24007 5620 24041 5654
rect 24080 5620 24114 5654
rect 24153 5620 24187 5654
rect 24226 5620 24260 5654
rect 24299 5620 24333 5654
rect 24372 5620 24406 5654
rect 24445 5620 24479 5654
rect 24518 5620 24552 5654
rect 24591 5620 24625 5654
rect 24664 5620 24698 5654
rect 24737 5620 24771 5654
rect 24810 5620 24844 5654
rect 24883 5620 24917 5654
rect 24956 5620 24990 5654
rect 23350 5548 23384 5582
rect 23424 5548 23458 5582
rect 23498 5548 23532 5582
rect 23572 5548 23606 5582
rect 23646 5548 23680 5582
rect 23720 5548 23754 5582
rect 23795 5548 23829 5582
rect 23870 5548 23904 5582
rect 23945 5548 23979 5582
rect 24020 5548 24054 5582
rect 24095 5548 24129 5582
rect 24170 5548 24204 5582
rect 24245 5548 24279 5582
rect 24320 5548 24354 5582
rect 24395 5548 24429 5582
rect 24470 5548 24504 5582
rect 24545 5548 24579 5582
rect 24620 5548 24654 5582
rect 24695 5548 24729 5582
rect 24770 5548 24804 5582
rect 24845 5548 24879 5582
rect 24920 5548 24954 5582
rect 24995 5548 25029 5582
rect 25070 5548 25104 5582
rect 1609 5518 1611 5533
rect 1611 5518 1643 5533
rect 1681 5531 1715 5542
rect 1609 5462 1643 5477
rect 1609 5443 1611 5462
rect 1611 5443 1643 5462
rect 1681 5471 1713 5492
rect 1713 5471 1715 5492
rect 1681 5458 1715 5471
rect 1609 5391 1643 5402
rect 1609 5368 1611 5391
rect 1611 5368 1643 5391
rect 1681 5400 1713 5419
rect 1713 5400 1715 5419
rect 1681 5385 1715 5400
rect 1681 5329 1713 5346
rect 1713 5329 1715 5346
rect 1609 5320 1643 5327
rect 1609 5293 1611 5320
rect 1611 5293 1643 5320
rect 1681 5312 1715 5329
rect 1681 5258 1713 5273
rect 1713 5258 1715 5273
rect 1609 5249 1643 5252
rect 1609 5218 1611 5249
rect 1611 5218 1643 5249
rect 1681 5239 1715 5258
rect 1681 5187 1713 5200
rect 1713 5187 1715 5200
rect 1609 5144 1611 5177
rect 1611 5144 1643 5177
rect 1681 5166 1715 5187
rect 1609 5143 1643 5144
rect 1681 5116 1713 5127
rect 1713 5116 1715 5127
rect 1609 5073 1611 5102
rect 1611 5073 1643 5102
rect 1681 5093 1715 5116
rect 1609 5068 1643 5073
rect 1681 5045 1713 5054
rect 1713 5045 1715 5054
rect 1609 5002 1611 5027
rect 1611 5002 1643 5027
rect 1609 4993 1643 5002
rect 1681 5020 1715 5045
rect 1681 4974 1713 4981
rect 1713 4974 1715 4981
rect 1609 4931 1611 4952
rect 1611 4931 1643 4952
rect 1609 4918 1643 4931
rect 1681 4947 1715 4974
rect 1681 4903 1713 4908
rect 1713 4903 1715 4908
rect 1609 4860 1611 4877
rect 1611 4860 1643 4877
rect 1609 4843 1643 4860
rect 1681 4874 1715 4903
rect 25070 5476 25104 5510
rect 1681 4832 1713 4835
rect 1713 4832 1715 4835
rect 1609 4789 1611 4802
rect 1611 4789 1643 4802
rect 1609 4768 1643 4789
rect 1681 4801 1715 4832
rect 1681 4760 1713 4762
rect 1713 4760 1715 4762
rect 1609 4718 1611 4727
rect 1611 4718 1643 4727
rect 1609 4693 1643 4718
rect 1681 4728 1715 4760
rect 1681 4688 1713 4689
rect 1713 4688 1715 4689
rect 1609 4646 1611 4652
rect 1611 4646 1643 4652
rect 1609 4618 1643 4646
rect 1681 4655 1715 4688
rect -303 4250 -301 4284
rect -301 4250 -197 4284
rect -303 4249 -197 4250
rect -303 4216 -267 4249
rect -303 4182 -301 4216
rect -301 4215 -267 4216
rect -267 4215 -233 4249
rect -233 4215 -199 4249
rect -199 4215 -197 4249
rect -301 4182 -197 4215
rect -303 4180 -197 4182
rect -303 4148 -267 4180
rect -303 4114 -301 4148
rect -301 4146 -267 4148
rect -267 4146 -233 4180
rect -233 4146 -199 4180
rect -199 4146 -197 4180
rect -301 4114 -197 4146
rect -303 4111 -197 4114
rect -303 4102 -267 4111
rect -267 4102 -233 4111
rect -233 4102 -199 4111
rect -231 4077 -199 4102
rect -199 4077 -197 4111
rect -231 4068 -197 4077
rect -303 4046 -301 4063
rect -301 4046 -269 4063
rect -303 4029 -269 4046
rect -231 4008 -199 4030
rect -199 4008 -197 4030
rect -231 3996 -197 4008
rect -303 3978 -301 3990
rect -301 3978 -269 3990
rect -303 3956 -269 3978
rect -231 3939 -199 3958
rect -199 3939 -197 3958
rect -231 3924 -197 3939
rect -303 3910 -301 3917
rect -301 3910 -269 3917
rect -303 3883 -269 3910
rect -231 3870 -199 3886
rect -199 3870 -197 3886
rect -231 3852 -197 3870
rect -303 3842 -301 3844
rect -301 3842 -269 3844
rect -303 3810 -269 3842
rect -231 3801 -199 3814
rect -199 3801 -197 3814
rect -231 3780 -197 3801
rect -303 3740 -269 3771
rect -303 3737 -301 3740
rect -301 3737 -269 3740
rect -231 3732 -199 3742
rect -199 3732 -197 3742
rect -231 3708 -197 3732
rect -303 3672 -269 3698
rect -303 3664 -301 3672
rect -301 3664 -269 3672
rect -231 3663 -199 3670
rect -199 3663 -197 3670
rect -231 3636 -197 3663
rect -303 3604 -269 3625
rect -303 3591 -301 3604
rect -301 3591 -269 3604
rect -231 3594 -199 3598
rect -199 3594 -197 3598
rect -231 3564 -197 3594
rect -303 3536 -269 3552
rect -303 3518 -301 3536
rect -301 3518 -269 3536
rect -231 3525 -199 3526
rect -199 3525 -197 3526
rect -231 3492 -197 3525
rect -303 3468 -269 3479
rect -303 3445 -301 3468
rect -301 3445 -269 3468
rect -231 3421 -197 3454
rect -303 3400 -269 3406
rect -303 3372 -301 3400
rect -301 3372 -269 3400
rect -231 3420 -199 3421
rect -199 3420 -197 3421
rect -231 3352 -197 3382
rect -303 3332 -269 3333
rect -303 3299 -301 3332
rect -301 3299 -269 3332
rect -231 3348 -199 3352
rect -199 3348 -197 3352
rect -231 3283 -197 3310
rect -303 3230 -301 3260
rect -301 3230 -269 3260
rect -231 3276 -199 3283
rect -199 3276 -197 3283
rect -303 3226 -269 3230
rect -231 3214 -197 3238
rect -303 3162 -301 3187
rect -301 3162 -269 3187
rect -231 3204 -199 3214
rect -199 3204 -197 3214
rect -303 3153 -269 3162
rect -231 3145 -197 3166
rect -303 3094 -301 3114
rect -301 3094 -269 3114
rect -231 3132 -199 3145
rect -199 3132 -197 3145
rect -303 3080 -269 3094
rect -231 3076 -197 3094
rect -231 3060 -199 3076
rect -199 3060 -197 3076
rect -303 3026 -301 3041
rect -301 3026 -269 3041
rect -303 3007 -269 3026
rect -231 3007 -197 3022
rect -231 2988 -199 3007
rect -199 2988 -197 3007
rect -303 2958 -301 2968
rect -301 2958 -269 2968
rect -303 2934 -269 2958
rect -231 2938 -197 2950
rect -231 2916 -199 2938
rect -199 2916 -197 2938
rect -303 2890 -301 2895
rect -301 2890 -269 2895
rect -303 2861 -269 2890
rect -231 2869 -197 2878
rect -231 2844 -199 2869
rect -199 2844 -197 2869
rect -303 2788 -269 2822
rect -231 2800 -197 2806
rect -231 2772 -199 2800
rect -199 2772 -197 2800
rect -303 2720 -269 2749
rect -231 2731 -197 2734
rect -303 2715 -301 2720
rect -301 2715 -269 2720
rect -231 2700 -199 2731
rect -199 2700 -197 2731
rect -303 2652 -269 2676
rect -303 2642 -301 2652
rect -301 2642 -269 2652
rect -231 2628 -199 2662
rect -199 2628 -197 2662
rect -303 2584 -269 2603
rect -303 2569 -301 2584
rect -301 2569 -269 2584
rect -231 2559 -199 2590
rect -199 2559 -197 2590
rect -231 2556 -197 2559
rect -303 2516 -269 2530
rect -303 2496 -301 2516
rect -301 2496 -269 2516
rect -231 2490 -199 2518
rect -199 2490 -197 2518
rect -231 2484 -197 2490
rect -303 2448 -269 2457
rect -303 2423 -301 2448
rect -301 2423 -269 2448
rect -231 2421 -199 2446
rect -199 2421 -197 2446
rect -231 2412 -197 2421
rect -303 2380 -269 2384
rect -303 2350 -301 2380
rect -301 2350 -269 2380
rect -231 2352 -199 2374
rect -199 2352 -197 2374
rect -231 2340 -197 2352
rect -303 2278 -301 2311
rect -301 2278 -269 2311
rect -231 2283 -199 2302
rect -199 2283 -197 2302
rect -303 2277 -269 2278
rect -231 2268 -197 2283
rect -303 2210 -301 2238
rect -301 2210 -269 2238
rect -231 2214 -199 2230
rect -199 2214 -197 2230
rect -303 2204 -269 2210
rect -231 2196 -197 2214
rect -303 2142 -301 2165
rect -301 2142 -269 2165
rect -231 2145 -199 2158
rect -199 2145 -197 2158
rect -303 2131 -269 2142
rect -231 2124 -197 2145
rect -303 2074 -301 2092
rect -301 2074 -269 2092
rect -231 2076 -199 2086
rect -199 2076 -197 2086
rect -303 2058 -269 2074
rect -231 2052 -197 2076
rect -303 2006 -301 2019
rect -301 2006 -269 2019
rect -231 2007 -199 2014
rect -199 2007 -197 2014
rect -303 1985 -269 2006
rect -231 1980 -197 2007
rect -303 1938 -301 1946
rect -301 1938 -269 1946
rect -231 1938 -199 1942
rect -199 1938 -197 1942
rect -303 1912 -269 1938
rect -231 1908 -197 1938
rect -303 1869 -301 1873
rect -301 1869 -269 1873
rect -231 1869 -199 1870
rect -199 1869 -197 1870
rect -303 1839 -269 1869
rect -231 1836 -197 1869
rect -303 1766 -269 1800
rect -231 1765 -197 1798
rect -231 1764 -199 1765
rect -199 1764 -197 1765
rect -303 1696 -269 1727
rect -231 1696 -197 1726
rect -303 1693 -301 1696
rect -301 1693 -269 1696
rect -231 1692 -199 1696
rect -199 1692 -197 1696
rect -303 1627 -269 1654
rect -231 1627 -197 1654
rect -303 1620 -301 1627
rect -301 1620 -269 1627
rect -231 1620 -199 1627
rect -199 1620 -197 1627
rect -303 1558 -269 1581
rect -231 1558 -197 1581
rect -303 1547 -301 1558
rect -301 1547 -269 1558
rect -231 1547 -199 1558
rect -199 1547 -197 1558
rect -303 1489 -269 1508
rect -231 1489 -197 1508
rect -303 1474 -301 1489
rect -301 1474 -269 1489
rect -231 1474 -199 1489
rect -199 1474 -197 1489
rect -303 1420 -269 1435
rect -231 1420 -197 1435
rect -303 1401 -301 1420
rect -301 1401 -269 1420
rect -231 1401 -199 1420
rect -199 1401 -197 1420
rect -303 1351 -269 1362
rect -231 1351 -197 1362
rect -303 1328 -301 1351
rect -301 1328 -269 1351
rect -231 1328 -199 1351
rect -199 1328 -197 1351
rect -303 1282 -269 1289
rect -231 1282 -197 1289
rect -303 1255 -301 1282
rect -301 1255 -269 1282
rect -231 1255 -199 1282
rect -199 1255 -197 1282
rect -303 1213 -269 1216
rect -231 1213 -197 1216
rect -303 1182 -301 1213
rect -301 1182 -269 1213
rect -231 1182 -199 1213
rect -199 1182 -197 1213
rect -303 1110 -301 1143
rect -301 1110 -269 1143
rect -231 1110 -199 1143
rect -199 1110 -197 1143
rect -303 1109 -269 1110
rect -231 1109 -197 1110
rect -303 1041 -301 1070
rect -301 1041 -269 1070
rect -231 1041 -199 1070
rect -199 1041 -197 1070
rect -303 1036 -269 1041
rect -231 1036 -197 1041
rect -303 972 -301 997
rect -301 972 -269 997
rect -231 972 -199 997
rect -199 972 -197 997
rect -303 963 -269 972
rect -231 963 -197 972
rect -303 903 -301 924
rect -301 903 -269 924
rect -231 903 -199 924
rect -199 903 -197 924
rect -303 890 -269 903
rect -231 890 -197 903
rect -303 834 -301 851
rect -301 834 -269 851
rect -231 834 -199 851
rect -199 834 -197 851
rect -303 817 -269 834
rect -231 817 -197 834
rect -303 765 -301 778
rect -301 765 -269 778
rect -231 765 -199 778
rect -199 765 -197 778
rect -303 744 -269 765
rect -231 744 -197 765
rect -303 696 -301 705
rect -301 696 -269 705
rect -231 696 -199 705
rect -199 696 -197 705
rect -303 671 -269 696
rect -231 671 -197 696
rect -303 627 -301 632
rect -301 627 -269 632
rect -231 627 -199 632
rect -199 627 -197 632
rect -303 598 -269 627
rect -231 598 -197 627
rect -303 558 -301 559
rect -301 558 -269 559
rect -231 558 -199 559
rect -199 558 -197 559
rect -303 525 -269 558
rect -231 525 -197 558
rect -303 454 -269 486
rect -231 454 -197 486
rect -303 452 -301 454
rect -301 452 -269 454
rect -231 452 -199 454
rect -199 452 -197 454
rect -303 385 -269 413
rect -231 385 -197 413
rect -303 379 -301 385
rect -301 379 -269 385
rect -231 379 -199 385
rect -199 379 -197 385
rect -303 316 -269 340
rect -231 316 -197 340
rect -303 306 -301 316
rect -301 306 -269 316
rect -231 306 -199 316
rect -199 306 -197 316
rect -303 247 -269 267
rect -231 247 -197 267
rect -303 233 -301 247
rect -301 233 -269 247
rect -231 233 -199 247
rect -199 233 -197 247
rect -303 178 -269 194
rect -231 178 -197 194
rect -303 160 -301 178
rect -301 160 -269 178
rect -231 160 -199 178
rect -199 160 -197 178
rect 77 4574 79 4596
rect 79 4574 113 4596
rect 113 4574 150 4596
rect 150 4574 183 4596
rect 740 4574 744 4577
rect 744 4574 774 4577
rect 813 4574 814 4577
rect 814 4574 847 4577
rect 77 4540 183 4574
rect 740 4543 774 4574
rect 813 4543 847 4574
rect 886 4543 920 4577
rect 959 4574 990 4577
rect 990 4574 993 4577
rect 1032 4574 1060 4577
rect 1060 4574 1066 4577
rect 1105 4574 1130 4577
rect 1130 4574 1139 4577
rect 1177 4574 1200 4577
rect 1200 4574 1211 4577
rect 1249 4574 1282 4577
rect 1282 4574 1283 4577
rect 959 4543 993 4574
rect 1032 4543 1066 4574
rect 1105 4543 1139 4574
rect 1177 4543 1211 4574
rect 1249 4543 1283 4574
rect 1321 4543 1355 4577
rect 1393 4543 1427 4577
rect 1465 4543 1499 4577
rect 1537 4574 1538 4577
rect 1538 4574 1571 4577
rect 1609 4574 1611 4577
rect 1611 4574 1643 4577
rect 1681 4582 1715 4616
rect 1537 4543 1571 4574
rect 1609 4543 1643 4574
rect 77 4506 113 4540
rect 113 4506 147 4540
rect 77 4472 147 4506
rect 147 4472 183 4540
rect 1681 4509 1715 4543
rect 740 4472 774 4505
rect 815 4472 849 4505
rect 890 4472 924 4505
rect 965 4472 999 4505
rect 1040 4472 1074 4505
rect 1115 4472 1149 4505
rect 1190 4472 1224 4505
rect 1265 4472 1299 4505
rect 1340 4472 1374 4505
rect 1415 4472 1449 4505
rect 1490 4472 1524 4505
rect 1565 4472 1599 4505
rect 77 3894 183 4472
rect 740 4471 765 4472
rect 765 4471 774 4472
rect 815 4471 838 4472
rect 838 4471 849 4472
rect 890 4471 911 4472
rect 911 4471 924 4472
rect 965 4471 984 4472
rect 984 4471 999 4472
rect 1040 4471 1056 4472
rect 1056 4471 1074 4472
rect 1115 4471 1128 4472
rect 1128 4471 1149 4472
rect 1190 4471 1200 4472
rect 1200 4471 1224 4472
rect 1265 4471 1282 4472
rect 1282 4471 1299 4472
rect 1340 4471 1360 4472
rect 1360 4471 1374 4472
rect 1415 4471 1438 4472
rect 1438 4471 1449 4472
rect 1490 4471 1516 4472
rect 1516 4471 1524 4472
rect 1565 4471 1593 4472
rect 1593 4471 1599 4472
rect 2208 4319 2242 4353
rect 2208 4247 2242 4281
rect 77 3860 79 3894
rect 79 3860 183 3894
rect 77 3859 183 3860
rect 77 3826 113 3859
rect 77 3792 79 3826
rect 79 3825 113 3826
rect 113 3825 147 3859
rect 147 3825 181 3859
rect 181 3825 183 3859
rect 79 3792 183 3825
rect 77 3790 183 3792
rect 77 3758 113 3790
rect 77 3724 79 3758
rect 79 3756 113 3758
rect 113 3756 147 3790
rect 147 3756 181 3790
rect 181 3756 183 3790
rect 79 3724 183 3756
rect 77 3721 183 3724
rect 77 3690 113 3721
rect 77 3656 79 3690
rect 79 3687 113 3690
rect 113 3687 147 3721
rect 147 3687 181 3721
rect 181 3687 183 3721
rect 79 3656 183 3687
rect 77 3652 183 3656
rect 77 3622 113 3652
rect 77 3588 79 3622
rect 79 3618 113 3622
rect 113 3618 147 3652
rect 147 3618 181 3652
rect 181 3618 183 3652
rect 79 3588 183 3618
rect 77 3583 183 3588
rect 77 3554 113 3583
rect 77 3520 79 3554
rect 79 3549 113 3554
rect 113 3549 147 3583
rect 147 3549 181 3583
rect 181 3549 183 3583
rect 79 3520 183 3549
rect 77 3514 183 3520
rect 77 3486 113 3514
rect 77 3452 79 3486
rect 79 3480 113 3486
rect 113 3480 147 3514
rect 147 3480 181 3514
rect 181 3480 183 3514
rect 79 3452 183 3480
rect 77 3445 183 3452
rect 77 3418 113 3445
rect 77 3384 79 3418
rect 79 3411 113 3418
rect 113 3411 147 3445
rect 147 3411 181 3445
rect 181 3411 183 3445
rect 79 3384 183 3411
rect 77 3376 183 3384
rect 77 3350 113 3376
rect 77 3316 79 3350
rect 79 3342 113 3350
rect 113 3342 147 3376
rect 147 3342 181 3376
rect 181 3342 183 3376
rect 79 3316 183 3342
rect 77 3307 183 3316
rect 77 3282 113 3307
rect 77 3248 79 3282
rect 79 3273 113 3282
rect 113 3273 147 3307
rect 147 3273 181 3307
rect 181 3273 183 3307
rect 79 3248 183 3273
rect 77 3238 183 3248
rect 77 3214 113 3238
rect 77 3180 79 3214
rect 79 3204 113 3214
rect 113 3204 147 3238
rect 147 3204 181 3238
rect 181 3204 183 3238
rect 79 3180 183 3204
rect 77 3169 183 3180
rect 77 3146 113 3169
rect 77 3112 79 3146
rect 79 3135 113 3146
rect 113 3135 147 3169
rect 147 3135 181 3169
rect 181 3135 183 3169
rect 79 3112 183 3135
rect 77 3100 183 3112
rect 77 3078 113 3100
rect 77 3044 79 3078
rect 79 3066 113 3078
rect 113 3066 147 3100
rect 147 3066 181 3100
rect 181 3066 183 3100
rect 79 3044 183 3066
rect 77 3031 183 3044
rect 77 3010 113 3031
rect 77 2976 79 3010
rect 79 2997 113 3010
rect 113 2997 147 3031
rect 147 2997 181 3031
rect 181 2997 183 3031
rect 79 2976 183 2997
rect 77 2962 183 2976
rect 77 2942 113 2962
rect 77 2908 79 2942
rect 79 2928 113 2942
rect 113 2928 147 2962
rect 147 2928 181 2962
rect 181 2928 183 2962
rect 79 2908 183 2928
rect 77 2893 183 2908
rect 77 2874 113 2893
rect 77 2840 79 2874
rect 79 2859 113 2874
rect 113 2859 147 2893
rect 147 2859 181 2893
rect 181 2859 183 2893
rect 79 2840 183 2859
rect 77 2824 183 2840
rect 77 2806 113 2824
rect 77 2772 79 2806
rect 79 2790 113 2806
rect 113 2790 147 2824
rect 147 2790 181 2824
rect 181 2790 183 2824
rect 79 2772 183 2790
rect 77 2755 183 2772
rect 77 2738 113 2755
rect 77 2704 79 2738
rect 79 2721 113 2738
rect 113 2721 147 2755
rect 147 2721 181 2755
rect 181 2721 183 2755
rect 79 2704 183 2721
rect 77 2686 183 2704
rect 77 2670 113 2686
rect 77 2636 79 2670
rect 79 2652 113 2670
rect 113 2652 147 2686
rect 147 2652 181 2686
rect 181 2652 183 2686
rect 79 2636 183 2652
rect 77 2617 183 2636
rect 77 2602 113 2617
rect 77 2568 79 2602
rect 79 2583 113 2602
rect 113 2583 147 2617
rect 147 2583 181 2617
rect 181 2583 183 2617
rect 79 2568 183 2583
rect 77 2548 183 2568
rect 77 2534 113 2548
rect 77 2500 79 2534
rect 79 2514 113 2534
rect 113 2514 147 2548
rect 147 2514 181 2548
rect 181 2514 183 2548
rect 79 2500 183 2514
rect 77 2479 183 2500
rect 77 2466 113 2479
rect 77 2432 79 2466
rect 79 2445 113 2466
rect 113 2445 147 2479
rect 147 2445 181 2479
rect 181 2445 183 2479
rect 79 2432 183 2445
rect 77 2410 183 2432
rect 77 2398 113 2410
rect 77 2364 79 2398
rect 79 2376 113 2398
rect 113 2376 147 2410
rect 147 2376 181 2410
rect 181 2376 183 2410
rect 79 2364 183 2376
rect 77 2341 183 2364
rect 77 2330 113 2341
rect 113 2330 147 2341
rect 147 2330 181 2341
rect 181 2330 183 2341
rect 77 2262 111 2291
rect 149 2272 183 2291
rect 77 2257 79 2262
rect 79 2257 111 2262
rect 149 2257 181 2272
rect 181 2257 183 2272
rect 77 2194 111 2218
rect 149 2203 183 2218
rect 77 2184 79 2194
rect 79 2184 111 2194
rect 149 2184 181 2203
rect 181 2184 183 2203
rect 77 2126 111 2145
rect 149 2134 183 2145
rect 77 2111 79 2126
rect 79 2111 111 2126
rect 149 2111 181 2134
rect 181 2111 183 2134
rect 77 2058 111 2072
rect 149 2065 183 2072
rect 77 2038 79 2058
rect 79 2038 111 2058
rect 149 2038 181 2065
rect 181 2038 183 2065
rect 77 1990 111 1999
rect 149 1996 183 1999
rect 77 1965 79 1990
rect 79 1965 111 1990
rect 149 1965 181 1996
rect 181 1965 183 1996
rect 77 1922 111 1926
rect 77 1892 79 1922
rect 79 1892 111 1922
rect 149 1893 181 1926
rect 181 1893 183 1926
rect 149 1892 183 1893
rect 77 1820 79 1853
rect 79 1820 111 1853
rect 149 1824 181 1853
rect 181 1824 183 1853
rect 77 1819 111 1820
rect 149 1819 183 1824
rect 77 1752 79 1780
rect 79 1752 111 1780
rect 149 1755 181 1780
rect 181 1755 183 1780
rect 77 1746 111 1752
rect 149 1746 183 1755
rect 77 1684 79 1707
rect 79 1684 111 1707
rect 149 1686 181 1707
rect 181 1686 183 1707
rect 77 1673 111 1684
rect 149 1673 183 1686
rect 77 1616 79 1634
rect 79 1616 111 1634
rect 149 1617 181 1634
rect 181 1617 183 1634
rect 77 1600 111 1616
rect 149 1600 183 1617
rect 77 1548 79 1561
rect 79 1548 111 1561
rect 149 1548 181 1561
rect 181 1548 183 1561
rect 77 1527 111 1548
rect 149 1527 183 1548
rect 77 1479 79 1488
rect 79 1479 111 1488
rect 149 1479 181 1488
rect 181 1479 183 1488
rect 77 1454 111 1479
rect 149 1454 183 1479
rect 77 1410 79 1415
rect 79 1410 111 1415
rect 149 1410 181 1415
rect 181 1410 183 1415
rect 77 1381 111 1410
rect 149 1381 183 1410
rect 77 1341 79 1342
rect 79 1341 111 1342
rect 149 1341 181 1342
rect 181 1341 183 1342
rect 77 1308 111 1341
rect 149 1308 183 1341
rect 77 1237 111 1269
rect 149 1237 183 1269
rect 77 1235 79 1237
rect 79 1235 111 1237
rect 149 1235 181 1237
rect 181 1235 183 1237
rect 77 1168 111 1196
rect 149 1168 183 1196
rect 77 1162 79 1168
rect 79 1162 111 1168
rect 149 1162 181 1168
rect 181 1162 183 1168
rect 77 1099 111 1123
rect 149 1099 183 1123
rect 77 1089 79 1099
rect 79 1089 111 1099
rect 149 1089 181 1099
rect 181 1089 183 1099
rect 77 1030 111 1050
rect 149 1030 183 1050
rect 77 1016 79 1030
rect 79 1016 111 1030
rect 149 1016 181 1030
rect 181 1016 183 1030
rect 77 961 111 977
rect 149 961 183 977
rect 77 943 79 961
rect 79 943 111 961
rect 149 943 181 961
rect 181 943 183 961
rect 77 892 111 904
rect 149 892 183 904
rect 77 870 79 892
rect 79 870 111 892
rect 149 870 181 892
rect 181 870 183 892
rect 77 823 111 831
rect 149 823 183 831
rect 77 797 79 823
rect 79 797 111 823
rect 149 797 181 823
rect 181 797 183 823
rect 77 754 111 758
rect 149 754 183 758
rect 77 724 79 754
rect 79 724 111 754
rect 149 724 181 754
rect 181 724 183 754
rect 77 651 79 685
rect 79 651 111 685
rect 149 651 181 685
rect 181 651 183 685
rect 77 582 79 612
rect 79 582 111 612
rect 149 582 181 612
rect 181 582 183 612
rect 77 578 111 582
rect 149 578 183 582
rect 77 513 79 539
rect 79 513 111 539
rect 149 513 181 539
rect 181 513 183 539
rect 77 505 111 513
rect 149 505 183 513
rect 77 444 79 466
rect 79 444 111 466
rect 149 444 181 466
rect 181 444 183 466
rect 77 432 111 444
rect 149 432 183 444
rect 77 375 79 393
rect 79 375 111 393
rect 149 375 181 393
rect 181 375 183 393
rect 77 359 111 375
rect 149 359 183 375
rect 77 306 79 320
rect 79 306 111 320
rect 729 4192 755 4226
rect 755 4192 763 4226
rect 803 4192 827 4226
rect 827 4192 837 4226
rect 877 4192 899 4226
rect 899 4192 911 4226
rect 951 4192 971 4226
rect 971 4192 985 4226
rect 1025 4192 1043 4226
rect 1043 4192 1059 4226
rect 1099 4192 1115 4226
rect 1115 4192 1133 4226
rect 1173 4192 1187 4226
rect 1187 4192 1207 4226
rect 1247 4192 1259 4226
rect 1259 4192 1281 4226
rect 1321 4192 1331 4226
rect 1331 4192 1355 4226
rect 1395 4192 1403 4226
rect 1403 4192 1429 4226
rect 1468 4192 1475 4226
rect 1475 4192 1502 4226
rect 1541 4192 1547 4226
rect 1547 4192 1575 4226
rect 1614 4192 1619 4226
rect 1619 4192 1648 4226
rect 1687 4192 1691 4226
rect 1691 4192 1721 4226
rect 555 3908 589 3942
rect 627 3908 661 3942
rect 699 3908 733 3942
rect 771 3908 805 3942
rect 843 3908 877 3942
rect 915 3908 949 3942
rect 1075 3908 1109 3942
rect 1147 3908 1181 3942
rect 1219 3908 1253 3942
rect 1291 3908 1325 3942
rect 1363 3908 1397 3942
rect 1435 3908 1469 3942
rect 2208 4175 2242 4209
rect 2208 4103 2242 4137
rect 2208 4031 2242 4065
rect 2351 4319 2385 4353
rect 2351 4247 2385 4281
rect 2351 4175 2385 4209
rect 2351 4103 2385 4137
rect 2351 4031 2385 4065
rect 5278 4332 5312 4366
rect 5278 4260 5312 4294
rect 5278 4188 5312 4222
rect 5278 4116 5312 4150
rect 5278 4044 5312 4078
rect 5416 4332 5450 4366
rect 5416 4260 5450 4294
rect 5416 4188 5450 4222
rect 5416 4116 5450 4150
rect 5416 4044 5450 4078
rect 4780 3908 4814 3942
rect 5709 3904 5815 3942
rect 5709 3870 5718 3904
rect 5718 3870 5752 3904
rect 5752 3870 5787 3904
rect 5787 3870 5815 3904
rect 6269 3880 6303 3886
rect 4780 3836 4814 3870
rect 5709 3836 5815 3870
rect 6269 3852 6303 3880
rect 6269 3812 6303 3814
rect 555 3486 589 3520
rect 627 3486 661 3520
rect 699 3486 733 3520
rect 771 3486 805 3520
rect 843 3486 877 3520
rect 915 3486 949 3520
rect 1075 3486 1109 3520
rect 1147 3486 1181 3520
rect 1219 3486 1253 3520
rect 1291 3486 1325 3520
rect 1363 3486 1397 3520
rect 1435 3486 1469 3520
rect 367 3318 401 3320
rect 367 3286 401 3318
rect 367 3216 401 3247
rect 367 3213 401 3216
rect 367 3148 401 3174
rect 367 3140 401 3148
rect 367 3080 401 3101
rect 367 3067 401 3080
rect 463 3348 497 3382
rect 1671 3746 1705 3780
rect 1743 3746 1777 3780
rect 1815 3746 1849 3780
rect 463 3276 497 3310
rect 463 3204 497 3238
rect 757 3192 791 3226
rect 829 3192 863 3226
rect 901 3192 935 3226
rect 973 3192 1007 3226
rect 1045 3192 1079 3226
rect 1117 3192 1151 3226
rect 1243 3179 1277 3182
rect 463 3132 497 3166
rect 1243 3148 1277 3179
rect 463 3060 497 3094
rect 604 3064 638 3098
rect 676 3064 710 3098
rect 748 3064 782 3098
rect 820 3064 854 3098
rect 367 3012 401 3028
rect 1243 3076 1277 3110
rect 367 2994 401 3012
rect 1243 3037 1277 3038
rect 1243 3004 1277 3037
rect 367 2944 401 2955
rect 367 2921 401 2944
rect 367 2876 401 2882
rect 367 2848 401 2876
rect 981 2908 1015 2942
rect 1053 2908 1087 2942
rect 1125 2908 1159 2942
rect 367 2808 401 2809
rect 367 2775 401 2808
rect 367 2706 401 2736
rect 604 2752 638 2786
rect 676 2752 710 2786
rect 748 2752 782 2786
rect 820 2752 854 2786
rect 367 2702 401 2706
rect 367 2638 401 2663
rect 367 2629 401 2638
rect 367 2570 401 2590
rect 367 2556 401 2570
rect 894 2596 928 2630
rect 966 2596 1000 2630
rect 1038 2596 1072 2630
rect 367 2502 401 2517
rect 367 2483 401 2502
rect 367 2434 401 2444
rect 367 2410 401 2434
rect 604 2440 638 2474
rect 676 2440 710 2474
rect 748 2440 782 2474
rect 820 2440 854 2474
rect 367 2366 401 2371
rect 367 2337 401 2366
rect 367 2264 401 2298
rect 981 2284 1015 2318
rect 1053 2284 1087 2318
rect 1125 2284 1159 2318
rect 367 2196 401 2225
rect 1243 2235 1277 2261
rect 1243 2227 1277 2235
rect 367 2191 401 2196
rect 367 2128 401 2152
rect 367 2118 401 2128
rect 604 2128 638 2162
rect 676 2128 710 2162
rect 748 2128 782 2162
rect 820 2128 854 2162
rect 1243 2163 1277 2189
rect 1243 2155 1277 2163
rect 367 2060 401 2079
rect 367 2045 401 2060
rect 1243 2091 1277 2117
rect 1243 2083 1277 2091
rect 367 1992 401 2006
rect 367 1972 401 1992
rect 367 1924 401 1933
rect 981 1972 1015 2006
rect 1053 1972 1087 2006
rect 1125 1972 1159 2006
rect 1243 2019 1277 2045
rect 1243 2011 1277 2019
rect 1243 1948 1277 1973
rect 1243 1939 1277 1948
rect 367 1899 401 1924
rect 367 1856 401 1860
rect 367 1826 401 1856
rect 1243 1877 1277 1901
rect 1243 1867 1277 1877
rect 6269 3780 6303 3812
rect 6269 3710 6303 3742
rect 6269 3708 6303 3710
rect 2100 3586 2101 3593
rect 2101 3586 2134 3593
rect 2100 3559 2134 3586
rect 4893 3586 4927 3620
rect 4965 3586 4999 3620
rect 5504 3586 5538 3620
rect 5576 3586 5610 3620
rect 5648 3586 5682 3620
rect 5720 3586 5754 3620
rect 5792 3586 5826 3620
rect 6269 3641 6303 3670
rect 6269 3636 6303 3641
rect 6269 3572 6303 3598
rect 6269 3564 6303 3572
rect 2100 3491 2101 3521
rect 2101 3491 2134 3521
rect 2100 3487 2134 3491
rect 6269 3503 6303 3526
rect 6269 3492 6303 3503
rect 6269 3434 6303 3454
rect 6269 3420 6303 3434
rect 6269 3365 6303 3382
rect 6269 3348 6303 3365
rect 6269 3296 6303 3310
rect 6269 3276 6303 3296
rect 6269 3227 6303 3238
rect 6269 3204 6303 3227
rect 6269 3158 6303 3166
rect 6269 3132 6303 3158
rect 6269 3089 6303 3093
rect 6269 3059 6303 3089
rect 6269 2986 6303 3020
rect 6269 2916 6303 2947
rect 6269 2913 6303 2916
rect 6269 2847 6303 2874
rect 6269 2840 6303 2847
rect 6269 2778 6303 2801
rect 6269 2767 6303 2778
rect 6269 2709 6303 2728
rect 6269 2694 6303 2709
rect 6269 2640 6303 2655
rect 6269 2621 6303 2640
rect 6269 2571 6303 2582
rect 6269 2548 6303 2571
rect 6269 2502 6303 2509
rect 1906 2483 1940 2492
rect 1906 2458 1917 2483
rect 1917 2458 1940 2483
rect 2045 2458 2079 2492
rect 2118 2458 2152 2492
rect 2191 2458 2207 2492
rect 2207 2458 2225 2492
rect 2264 2458 2275 2492
rect 2275 2458 2298 2492
rect 2337 2458 2343 2492
rect 2343 2458 2371 2492
rect 2410 2458 2411 2492
rect 2411 2458 2444 2492
rect 2483 2458 2513 2492
rect 2513 2458 2517 2492
rect 2556 2458 2581 2492
rect 2581 2458 2590 2492
rect 2629 2458 2649 2492
rect 2649 2458 2663 2492
rect 2702 2458 2717 2492
rect 2717 2458 2736 2492
rect 2775 2458 2785 2492
rect 2785 2458 2809 2492
rect 2848 2458 2854 2492
rect 2854 2458 2882 2492
rect 2921 2458 2923 2492
rect 2923 2458 2955 2492
rect 2994 2458 3027 2492
rect 3027 2458 3028 2492
rect 3067 2458 3096 2492
rect 3096 2458 3101 2492
rect 3140 2458 3165 2492
rect 3165 2458 3174 2492
rect 3213 2458 3234 2492
rect 3234 2458 3247 2492
rect 3286 2458 3303 2492
rect 3303 2458 3320 2492
rect 3359 2458 3372 2492
rect 3372 2458 3393 2492
rect 3432 2458 3441 2492
rect 3441 2458 3466 2492
rect 3505 2458 3510 2492
rect 3510 2458 3539 2492
rect 3578 2458 3579 2492
rect 3579 2458 3612 2492
rect 3651 2458 3682 2492
rect 3682 2458 3685 2492
rect 3723 2458 3751 2492
rect 3751 2458 3757 2492
rect 3795 2458 3820 2492
rect 3820 2458 3829 2492
rect 3867 2458 3889 2492
rect 3889 2458 3901 2492
rect 3939 2458 3958 2492
rect 3958 2458 3973 2492
rect 4011 2458 4027 2492
rect 4027 2458 4045 2492
rect 4083 2458 4096 2492
rect 4096 2458 4117 2492
rect 4155 2458 4165 2492
rect 4165 2458 4189 2492
rect 4227 2458 4234 2492
rect 4234 2458 4261 2492
rect 4299 2458 4303 2492
rect 4303 2458 4333 2492
rect 4371 2458 4372 2492
rect 4372 2458 4405 2492
rect 4443 2458 4476 2492
rect 4476 2458 4477 2492
rect 4515 2458 4545 2492
rect 4545 2458 4549 2492
rect 4587 2458 4614 2492
rect 4614 2458 4621 2492
rect 4659 2458 4683 2492
rect 4683 2458 4693 2492
rect 6269 2475 6303 2502
rect 1906 2411 1940 2420
rect 1906 2386 1917 2411
rect 1917 2386 1940 2411
rect 6269 2433 6303 2436
rect 5504 2330 5538 2364
rect 5576 2330 5610 2364
rect 5648 2330 5682 2364
rect 5720 2330 5754 2364
rect 5792 2330 5826 2364
rect 6269 2402 6303 2433
rect 6269 2330 6303 2363
rect 6269 2329 6303 2330
rect 367 1754 401 1787
rect 367 1753 401 1754
rect 367 1686 401 1714
rect 367 1680 401 1686
rect 6269 2261 6303 2290
rect 6269 2256 6303 2261
rect 367 1618 401 1641
rect 367 1607 401 1618
rect 367 1550 401 1567
rect 367 1533 401 1550
rect 1040 1550 1074 1584
rect 1112 1550 1146 1584
rect 1184 1550 1218 1584
rect 1256 1550 1290 1584
rect 1328 1550 1362 1584
rect 1400 1550 1434 1584
rect 367 1482 401 1493
rect 367 1459 401 1482
rect 367 1414 401 1419
rect 367 1385 401 1414
rect 604 1394 638 1428
rect 676 1394 710 1428
rect 748 1394 782 1428
rect 820 1394 854 1428
rect 1235 1394 1269 1428
rect 1307 1394 1341 1428
rect 1379 1394 1413 1428
rect 1451 1394 1485 1428
rect 367 1312 401 1345
rect 367 1311 401 1312
rect 367 1244 401 1271
rect 367 1237 401 1244
rect 367 1176 401 1197
rect 367 1163 401 1176
rect 367 1108 401 1123
rect 367 1089 401 1108
rect 367 1040 401 1049
rect 367 1015 401 1040
rect 604 1082 638 1116
rect 676 1082 710 1116
rect 748 1082 782 1116
rect 820 1082 854 1116
rect 1235 1082 1269 1116
rect 1307 1082 1341 1116
rect 1379 1082 1413 1116
rect 1451 1082 1485 1116
rect 367 972 401 975
rect 367 941 401 972
rect 367 870 401 901
rect 367 867 401 870
rect 367 802 401 827
rect 367 793 401 802
rect 367 733 401 753
rect 367 719 401 733
rect 367 664 401 679
rect 367 645 401 664
rect 367 595 401 605
rect 367 571 401 595
rect 367 526 401 531
rect 367 497 401 526
rect 367 423 401 457
rect 367 354 401 383
rect 367 349 401 354
rect 463 489 497 523
rect 463 417 497 451
rect 149 306 181 320
rect 181 306 183 320
rect 77 286 111 306
rect 149 286 183 306
rect 77 237 79 247
rect 79 237 111 247
rect 149 237 181 247
rect 181 237 183 247
rect 77 213 111 237
rect 149 213 183 237
rect 77 168 79 174
rect 79 168 111 174
rect 149 168 181 174
rect 181 168 183 174
rect 6269 2192 6303 2217
rect 6269 2183 6303 2192
rect 6269 2123 6303 2144
rect 6269 2110 6303 2123
rect 5504 2018 5538 2052
rect 5576 2018 5610 2052
rect 5648 2018 5682 2052
rect 5720 2018 5754 2052
rect 5792 2018 5826 2052
rect 6269 2054 6303 2071
rect 6269 2037 6303 2054
rect 6269 1985 6303 1998
rect 6269 1964 6303 1985
rect 6269 1916 6303 1925
rect 6269 1891 6303 1916
rect 6269 1847 6303 1852
rect 6269 1818 6303 1847
rect 5504 1706 5538 1740
rect 5576 1706 5610 1740
rect 5648 1706 5682 1740
rect 5720 1706 5754 1740
rect 5792 1706 5826 1740
rect 6269 1778 6303 1779
rect 6269 1745 6303 1778
rect 6269 1674 6303 1706
rect 6269 1672 6303 1674
rect 6269 1605 6303 1633
rect 6269 1599 6303 1605
rect 6269 1536 6303 1560
rect 6269 1526 6303 1536
rect 5504 1394 5538 1428
rect 5576 1394 5610 1428
rect 5648 1394 5682 1428
rect 5720 1394 5754 1428
rect 5792 1394 5826 1428
rect 6269 1467 6303 1487
rect 6269 1453 6303 1467
rect 6269 1398 6303 1414
rect 6269 1380 6303 1398
rect 6269 1329 6303 1341
rect 6269 1307 6303 1329
rect 6269 1260 6303 1268
rect 6269 1234 6303 1260
rect 6269 1191 6303 1195
rect 6269 1161 6303 1191
rect 5504 1082 5538 1116
rect 5576 1082 5610 1116
rect 5648 1082 5682 1116
rect 5720 1082 5754 1116
rect 5792 1082 5826 1116
rect 6269 1088 6303 1122
rect 6269 1019 6303 1049
rect 6269 1015 6303 1019
rect 5134 926 5168 960
rect 5206 926 5240 960
rect 5278 926 5312 960
rect 5350 926 5384 960
rect 5422 926 5456 960
rect 6487 3503 6521 3537
rect 6559 3503 6593 3537
rect 6487 3428 6521 3462
rect 6559 3428 6593 3462
rect 6487 3353 6521 3387
rect 6559 3353 6593 3387
rect 25070 3316 25176 5472
rect 6487 3278 6521 3312
rect 6559 3278 6593 3312
rect 25142 3278 25176 3312
rect 25070 3243 25104 3277
rect 6487 3204 6521 3238
rect 6559 3204 6593 3238
rect 25142 3206 25176 3240
rect 25070 3170 25104 3204
rect 6487 3130 6521 3164
rect 6559 3130 6593 3164
rect 25142 3134 25176 3168
rect 25070 3097 25104 3131
rect 6487 3056 6521 3090
rect 6559 3056 6593 3090
rect 25142 3062 25176 3096
rect 25070 3024 25104 3058
rect 6487 2982 6521 3016
rect 6559 2982 6593 3016
rect 25142 2990 25176 3024
rect 25070 2951 25104 2985
rect 6487 2908 6521 2942
rect 6559 2908 6593 2942
rect 25142 2917 25176 2951
rect 25070 2878 25104 2912
rect 6487 2834 6521 2868
rect 6559 2834 6593 2868
rect 25142 2844 25176 2878
rect 25070 2805 25104 2839
rect 6487 2760 6521 2794
rect 6559 2760 6593 2794
rect 25142 2771 25176 2805
rect 25070 2732 25104 2766
rect 6487 2686 6521 2720
rect 6559 2686 6593 2720
rect 25142 2698 25176 2732
rect 25070 2659 25104 2693
rect 6487 2612 6521 2646
rect 6559 2612 6593 2646
rect 25142 2625 25176 2659
rect 25070 2586 25104 2620
rect 6487 2538 6521 2572
rect 6559 2538 6593 2572
rect 25142 2552 25176 2586
rect 25070 2513 25104 2547
rect 6487 2464 6521 2498
rect 6559 2464 6593 2498
rect 25142 2479 25176 2513
rect 25070 2440 25104 2474
rect 6487 2390 6521 2424
rect 6559 2390 6593 2424
rect 25142 2406 25176 2440
rect 25070 2367 25104 2401
rect 6487 2316 6521 2350
rect 6559 2316 6593 2350
rect 25142 2333 25176 2367
rect 25070 2294 25104 2328
rect 6487 2242 6521 2276
rect 6559 2242 6593 2276
rect 25142 2260 25176 2294
rect 25070 2221 25104 2255
rect 6487 2168 6521 2202
rect 6559 2168 6593 2202
rect 25142 2187 25176 2221
rect 25070 2148 25104 2182
rect 6487 2094 6521 2128
rect 6559 2094 6593 2128
rect 25142 2114 25176 2148
rect 25070 2075 25104 2109
rect 6487 2020 6521 2054
rect 6559 2020 6593 2054
rect 25142 2041 25176 2075
rect 25792 2058 25898 6133
rect 25070 2002 25104 2036
rect 25792 2023 25898 2058
rect 6487 1946 6521 1980
rect 6559 1946 6593 1980
rect 25142 1968 25176 2002
rect 25792 1989 25812 2023
rect 25812 1989 25846 2023
rect 25846 1989 25880 2023
rect 25880 1989 25898 2023
rect 25070 1929 25104 1963
rect 25792 1954 25898 1989
rect 6487 1872 6521 1906
rect 6559 1872 6593 1906
rect 25142 1895 25176 1929
rect 25792 1920 25812 1954
rect 25812 1920 25846 1954
rect 25846 1920 25880 1954
rect 25880 1920 25898 1954
rect 25070 1856 25104 1890
rect 25792 1885 25898 1920
rect 6487 1798 6521 1832
rect 6559 1798 6593 1832
rect 25142 1822 25176 1856
rect 25792 1851 25812 1885
rect 25812 1851 25846 1885
rect 25846 1851 25880 1885
rect 25880 1851 25898 1885
rect 25070 1783 25104 1817
rect 25792 1816 25898 1851
rect 6487 1724 6521 1758
rect 6559 1724 6593 1758
rect 25142 1749 25176 1783
rect 25792 1782 25812 1816
rect 25812 1782 25846 1816
rect 25846 1782 25880 1816
rect 25880 1782 25898 1816
rect 25792 1747 25898 1782
rect 25070 1710 25104 1744
rect 25792 1713 25812 1747
rect 25812 1713 25846 1747
rect 25846 1713 25880 1747
rect 25880 1713 25898 1747
rect 6487 1650 6521 1684
rect 6559 1650 6593 1684
rect 25142 1676 25176 1710
rect 25792 1678 25898 1713
rect 25070 1637 25104 1671
rect 25792 1644 25812 1678
rect 25812 1644 25846 1678
rect 25846 1644 25880 1678
rect 25880 1644 25898 1678
rect 6487 1576 6521 1610
rect 6559 1576 6593 1610
rect 25142 1603 25176 1637
rect 25792 1609 25898 1644
rect 25070 1564 25104 1598
rect 25792 1575 25812 1609
rect 25812 1575 25846 1609
rect 25846 1575 25880 1609
rect 25880 1575 25898 1609
rect 6487 1502 6521 1536
rect 6559 1502 6593 1536
rect 25142 1530 25176 1564
rect 25792 1540 25898 1575
rect 25070 1491 25104 1525
rect 25792 1506 25812 1540
rect 25812 1506 25846 1540
rect 25846 1506 25880 1540
rect 25880 1506 25898 1540
rect 6487 1428 6521 1462
rect 6559 1428 6593 1462
rect 25142 1457 25176 1491
rect 25792 1471 25898 1506
rect 25070 1418 25104 1452
rect 25792 1437 25812 1471
rect 25812 1437 25846 1471
rect 25846 1437 25880 1471
rect 25880 1437 25898 1471
rect 6487 1354 6521 1388
rect 6559 1354 6593 1388
rect 25142 1384 25176 1418
rect 25792 1402 25898 1437
rect 25070 1345 25104 1379
rect 25792 1368 25812 1402
rect 25812 1368 25846 1402
rect 25846 1368 25880 1402
rect 25880 1368 25898 1402
rect 6487 1280 6521 1314
rect 6559 1280 6593 1314
rect 25142 1311 25176 1345
rect 25792 1333 25898 1368
rect 25070 1272 25104 1306
rect 25792 1299 25812 1333
rect 25812 1299 25846 1333
rect 25846 1299 25880 1333
rect 25880 1299 25898 1333
rect 6487 1206 6521 1240
rect 6559 1206 6593 1240
rect 25142 1238 25176 1272
rect 25792 1264 25898 1299
rect 25070 1199 25104 1233
rect 25792 1230 25812 1264
rect 25812 1230 25846 1264
rect 25846 1230 25880 1264
rect 25880 1230 25898 1264
rect 6487 1132 6521 1166
rect 6559 1132 6593 1166
rect 25142 1165 25176 1199
rect 25792 1195 25898 1230
rect 25792 1161 25812 1195
rect 25812 1161 25846 1195
rect 25846 1161 25880 1195
rect 25880 1161 25898 1195
rect 25070 1126 25104 1160
rect 25792 1126 25898 1161
rect 25142 1092 25176 1126
rect 25792 1092 25812 1126
rect 25812 1092 25846 1126
rect 25846 1092 25880 1126
rect 25880 1092 25898 1126
rect 6487 1058 6521 1092
rect 6559 1058 6593 1092
rect 25070 1053 25104 1087
rect 25792 1057 25898 1092
rect 25142 1019 25176 1053
rect 25792 1023 25812 1057
rect 25812 1023 25846 1057
rect 25846 1023 25880 1057
rect 25880 1023 25898 1057
rect 6487 984 6521 1018
rect 6559 984 6593 1018
rect 25070 980 25104 1014
rect 25792 988 25898 1023
rect 6269 950 6303 976
rect 6269 942 6303 950
rect 25142 946 25176 980
rect 25792 954 25812 988
rect 25812 954 25846 988
rect 25846 954 25880 988
rect 25880 954 25898 988
rect 25070 907 25104 941
rect 25792 919 25898 954
rect 6269 881 6303 903
rect 6269 869 6303 881
rect 25142 873 25176 907
rect 25792 915 25812 919
rect 25812 915 25846 919
rect 25846 915 25880 919
rect 25880 915 25898 919
rect 5504 770 5538 804
rect 5576 770 5610 804
rect 5648 770 5682 804
rect 5720 770 5754 804
rect 5792 770 5826 804
rect 25070 834 25104 868
rect 25792 850 25826 876
rect 25864 850 25898 876
rect 6269 812 6303 830
rect 6269 796 6303 812
rect 25142 800 25176 834
rect 25792 842 25812 850
rect 25812 842 25826 850
rect 25864 842 25880 850
rect 25880 842 25898 850
rect 25070 761 25104 795
rect 25792 781 25826 803
rect 25864 781 25898 803
rect 6269 743 6303 757
rect 6269 723 6303 743
rect 25142 727 25176 761
rect 25792 769 25812 781
rect 25812 769 25826 781
rect 25864 769 25880 781
rect 25880 769 25898 781
rect 5134 614 5168 648
rect 5206 614 5240 648
rect 5278 614 5312 648
rect 5350 614 5384 648
rect 5422 614 5456 648
rect 25070 688 25104 722
rect 25792 712 25826 730
rect 25864 712 25898 730
rect 6269 674 6303 684
rect 6269 650 6303 674
rect 25142 654 25176 688
rect 25792 696 25812 712
rect 25812 696 25826 712
rect 25864 696 25880 712
rect 25880 696 25898 712
rect 25070 615 25104 649
rect 25792 643 25826 657
rect 25864 643 25898 657
rect 6269 605 6303 611
rect 6269 577 6303 605
rect 25142 581 25176 615
rect 25792 623 25812 643
rect 25812 623 25826 643
rect 25864 623 25880 643
rect 25880 623 25898 643
rect 25070 542 25104 576
rect 25792 574 25826 584
rect 25864 574 25898 584
rect 6269 536 6303 538
rect 6269 504 6303 536
rect 25142 508 25176 542
rect 25792 550 25812 574
rect 25812 550 25826 574
rect 25864 550 25880 574
rect 25880 550 25898 574
rect 25792 505 25826 511
rect 25864 505 25898 511
rect 25070 469 25104 503
rect 25792 477 25812 505
rect 25812 477 25826 505
rect 25864 477 25880 505
rect 25880 477 25898 505
rect 6269 432 6303 465
rect 25142 435 25176 469
rect 25792 436 25826 438
rect 25864 436 25898 438
rect 6269 431 6303 432
rect 25070 396 25104 430
rect 25792 404 25812 436
rect 25812 404 25826 436
rect 25864 404 25880 436
rect 25880 404 25898 436
rect 541 330 565 364
rect 565 330 575 364
rect 614 330 633 364
rect 633 330 648 364
rect 687 330 701 364
rect 701 330 721 364
rect 760 330 769 364
rect 769 330 794 364
rect 833 330 837 364
rect 837 330 867 364
rect 906 330 939 364
rect 939 330 940 364
rect 979 330 1007 364
rect 1007 330 1013 364
rect 1052 330 1075 364
rect 1075 330 1086 364
rect 1125 330 1143 364
rect 1143 330 1159 364
rect 1198 330 1211 364
rect 1211 330 1232 364
rect 1271 330 1279 364
rect 1279 330 1305 364
rect 1344 330 1347 364
rect 1347 330 1378 364
rect 1417 330 1449 364
rect 1449 330 1451 364
rect 1490 330 1517 364
rect 1517 330 1524 364
rect 1563 330 1585 364
rect 1585 330 1597 364
rect 1636 330 1653 364
rect 1653 330 1670 364
rect 1709 330 1743 364
rect 1782 330 1816 364
rect 1855 330 1889 364
rect 1928 330 1962 364
rect 2000 330 2027 364
rect 2027 330 2034 364
rect 2072 330 2095 364
rect 2095 330 2106 364
rect 2144 330 2163 364
rect 2163 330 2178 364
rect 2216 330 2231 364
rect 2231 330 2250 364
rect 2288 330 2299 364
rect 2299 330 2322 364
rect 2360 330 2367 364
rect 2367 330 2394 364
rect 2432 330 2435 364
rect 2435 330 2466 364
rect 2504 330 2537 364
rect 2537 330 2538 364
rect 2576 330 2605 364
rect 2605 330 2610 364
rect 2648 330 2673 364
rect 2673 330 2682 364
rect 2720 330 2741 364
rect 2741 330 2754 364
rect 2792 330 2809 364
rect 2809 330 2826 364
rect 2864 330 2877 364
rect 2877 330 2898 364
rect 2936 330 2945 364
rect 2945 330 2970 364
rect 3008 330 3013 364
rect 3013 330 3042 364
rect 3080 330 3081 364
rect 3081 330 3114 364
rect 3152 330 3183 364
rect 3183 330 3186 364
rect 3224 330 3251 364
rect 3251 330 3258 364
rect 3296 330 3319 364
rect 3319 330 3330 364
rect 3368 330 3387 364
rect 3387 330 3402 364
rect 3440 330 3455 364
rect 3455 330 3474 364
rect 3512 330 3523 364
rect 3523 330 3546 364
rect 3584 330 3591 364
rect 3591 330 3618 364
rect 3656 330 3659 364
rect 3659 330 3690 364
rect 3728 330 3761 364
rect 3761 330 3762 364
rect 3800 330 3830 364
rect 3830 330 3834 364
rect 3872 330 3899 364
rect 3899 330 3906 364
rect 3944 330 3968 364
rect 3968 330 3978 364
rect 4016 330 4037 364
rect 4037 330 4050 364
rect 4088 330 4106 364
rect 4106 330 4122 364
rect 4160 330 4175 364
rect 4175 330 4194 364
rect 4232 330 4244 364
rect 4244 330 4266 364
rect 4304 330 4313 364
rect 4313 330 4338 364
rect 4376 330 4382 364
rect 4382 330 4410 364
rect 4448 330 4451 364
rect 4451 330 4482 364
rect 4520 330 4554 364
rect 4592 330 4623 364
rect 4623 330 4626 364
rect 4664 330 4692 364
rect 4692 330 4698 364
rect 25142 362 25176 396
rect 25070 323 25104 357
rect 25792 333 25812 365
rect 25812 333 25826 365
rect 25864 333 25880 365
rect 25880 333 25898 365
rect 25792 331 25826 333
rect 25864 331 25898 333
rect 25142 289 25176 323
rect 677 168 783 274
rect 25070 250 25104 284
rect 25792 264 25812 292
rect 25812 264 25826 292
rect 25864 264 25880 292
rect 25880 264 25898 292
rect 25792 258 25826 264
rect 25864 258 25898 264
rect 25142 216 25176 250
rect 25070 177 25104 211
rect 25792 195 25812 219
rect 25812 195 25826 219
rect 25864 195 25880 219
rect 25880 195 25898 219
rect 25792 185 25826 195
rect 25864 185 25898 195
rect 77 140 111 168
rect 149 140 183 168
rect 25142 143 25176 177
rect 24413 104 24447 138
rect 24486 104 24520 138
rect 24559 104 24593 138
rect 24632 104 24666 138
rect 24705 104 24739 138
rect 24778 104 24812 138
rect 24851 104 24885 138
rect 24924 104 24958 138
rect 24997 104 25031 138
rect 25070 104 25104 138
rect 25792 126 25812 146
rect 25812 126 25826 146
rect 25864 126 25880 146
rect 25880 126 25898 146
rect 25792 112 25826 126
rect 25864 112 25898 126
rect 25142 70 25176 104
rect 24456 32 24490 66
rect 24528 32 24562 66
rect 24600 32 24634 66
rect 24672 32 24706 66
rect 24744 32 24778 66
rect 24816 32 24850 66
rect 24888 32 24922 66
rect 24960 32 24994 66
rect 25032 32 25066 66
rect 25792 57 25812 73
rect 25812 57 25826 73
rect 25864 57 25880 73
rect 25880 57 25898 73
rect 25792 39 25826 57
rect 25864 39 25898 57
rect 26181 6455 26215 6468
rect 26181 6434 26183 6455
rect 26183 6434 26215 6455
rect 26253 6456 26285 6468
rect 26285 6456 26287 6468
rect 26253 6434 26287 6456
rect 26181 6386 26215 6395
rect 26181 6361 26183 6386
rect 26183 6361 26215 6386
rect 26253 6388 26285 6395
rect 26285 6388 26287 6395
rect 26253 6361 26287 6388
rect 26181 6317 26215 6322
rect 26181 6288 26183 6317
rect 26183 6288 26215 6317
rect 26253 6320 26285 6322
rect 26285 6320 26287 6322
rect 26253 6288 26287 6320
rect 26181 6248 26215 6249
rect 26181 6215 26183 6248
rect 26183 6215 26215 6248
rect 26253 6218 26287 6249
rect 26253 6215 26285 6218
rect 26285 6215 26287 6218
rect 26181 6145 26183 6176
rect 26183 6145 26215 6176
rect 26181 6142 26215 6145
rect 26253 6150 26287 6176
rect 26253 6142 26285 6150
rect 26285 6142 26287 6150
rect 26181 6076 26183 6103
rect 26183 6076 26215 6103
rect 26181 6069 26215 6076
rect 26253 6082 26287 6103
rect 26253 6069 26285 6082
rect 26285 6069 26287 6082
rect 26181 6007 26183 6030
rect 26183 6007 26215 6030
rect 26181 5996 26215 6007
rect 26253 6014 26287 6030
rect 26253 5996 26285 6014
rect 26285 5996 26287 6014
rect 26181 5938 26183 5957
rect 26183 5938 26215 5957
rect 26181 5923 26215 5938
rect 26253 5946 26287 5957
rect 26253 5923 26285 5946
rect 26285 5923 26287 5946
rect 26181 5869 26183 5884
rect 26183 5869 26215 5884
rect 26181 5850 26215 5869
rect 26253 5878 26287 5884
rect 26253 5850 26285 5878
rect 26285 5850 26287 5878
rect 26181 5800 26183 5811
rect 26183 5800 26215 5811
rect 26181 5777 26215 5800
rect 26253 5810 26287 5811
rect 26253 5777 26285 5810
rect 26285 5777 26287 5810
rect 26181 5731 26183 5738
rect 26183 5731 26215 5738
rect 26181 5704 26215 5731
rect 26253 5708 26285 5738
rect 26285 5708 26287 5738
rect 26253 5704 26287 5708
rect 26181 5662 26183 5665
rect 26183 5662 26215 5665
rect 26181 5631 26215 5662
rect 26253 5640 26285 5665
rect 26285 5640 26287 5665
rect 26253 5631 26287 5640
rect 26181 5558 26215 5592
rect 26253 5572 26285 5592
rect 26285 5572 26287 5592
rect 26253 5558 26287 5572
rect 26181 5489 26215 5519
rect 26181 5485 26183 5489
rect 26183 5485 26215 5489
rect 26253 5504 26285 5519
rect 26285 5504 26287 5519
rect 26253 5485 26287 5504
rect 26181 5420 26215 5446
rect 26181 5412 26183 5420
rect 26183 5412 26215 5420
rect 26253 5436 26285 5446
rect 26285 5436 26287 5446
rect 26253 5412 26287 5436
rect 26181 5351 26215 5373
rect 26181 5339 26183 5351
rect 26183 5339 26215 5351
rect 26253 5368 26285 5373
rect 26285 5368 26287 5373
rect 26253 5339 26287 5368
rect 26181 5282 26215 5300
rect 26181 5266 26183 5282
rect 26183 5266 26215 5282
rect 26253 5266 26287 5300
rect 26181 5213 26215 5227
rect 26181 5193 26183 5213
rect 26183 5193 26215 5213
rect 26253 5198 26287 5227
rect 26253 5193 26285 5198
rect 26285 5193 26287 5198
rect 26181 5144 26215 5154
rect 26181 5120 26183 5144
rect 26183 5120 26215 5144
rect 26253 5130 26287 5154
rect 26253 5120 26285 5130
rect 26285 5120 26287 5130
rect 26181 5075 26215 5081
rect 26181 5047 26183 5075
rect 26183 5047 26215 5075
rect 26253 5062 26287 5081
rect 26253 5047 26285 5062
rect 26285 5047 26287 5062
rect 26181 5006 26215 5008
rect 26181 4974 26183 5006
rect 26183 4974 26215 5006
rect 26253 4994 26287 5008
rect 26253 4974 26285 4994
rect 26285 4974 26287 4994
rect 26181 4903 26183 4935
rect 26183 4903 26215 4935
rect 26181 4901 26215 4903
rect 26253 4926 26287 4935
rect 26253 4901 26285 4926
rect 26285 4901 26287 4926
rect 26181 4834 26183 4862
rect 26183 4834 26215 4862
rect 26181 4828 26215 4834
rect 26253 4858 26287 4862
rect 26253 4828 26285 4858
rect 26285 4828 26287 4858
rect 26181 4765 26183 4789
rect 26183 4765 26215 4789
rect 26181 4755 26215 4765
rect 26253 4756 26285 4789
rect 26285 4756 26287 4789
rect 26253 4755 26287 4756
rect 26181 4696 26183 4716
rect 26183 4696 26215 4716
rect 26181 4682 26215 4696
rect 26253 4688 26285 4716
rect 26285 4688 26287 4716
rect 26253 4682 26287 4688
rect 26181 4627 26183 4643
rect 26183 4627 26215 4643
rect 26181 4609 26215 4627
rect 26253 4620 26285 4643
rect 26285 4620 26287 4643
rect 26253 4609 26287 4620
rect 26181 4558 26183 4570
rect 26183 4558 26215 4570
rect 26181 4536 26215 4558
rect 26253 4552 26285 4570
rect 26285 4552 26287 4570
rect 26253 4536 26287 4552
rect 26181 4489 26183 4497
rect 26183 4489 26215 4497
rect 26181 4463 26215 4489
rect 26253 4484 26285 4497
rect 26285 4484 26287 4497
rect 26253 4463 26287 4484
rect 26181 4420 26183 4424
rect 26183 4420 26215 4424
rect 26181 4390 26215 4420
rect 26253 4416 26285 4424
rect 26285 4416 26287 4424
rect 26253 4390 26287 4416
rect 26181 4350 26217 4351
rect 26217 4350 26251 4351
rect 26251 4350 26285 4351
rect 26181 4348 26285 4350
rect 26285 4348 26287 4351
rect 26181 4316 26287 4348
rect 26181 4282 26183 4316
rect 26183 4315 26287 4316
rect 26183 4282 26217 4315
rect 26181 4281 26217 4282
rect 26217 4281 26251 4315
rect 26251 4314 26287 4315
rect 26251 4281 26285 4314
rect 26181 4280 26285 4281
rect 26285 4280 26287 4314
rect 26181 4247 26287 4280
rect 26181 4213 26183 4247
rect 26183 4246 26287 4247
rect 26183 4213 26217 4246
rect 26181 4178 26217 4213
rect 26217 4178 26287 4246
rect 26181 64 26287 4178
rect 26181 -147 26287 64
<< metal1 >>
rect -309 6766 26293 6772
rect -309 6732 -265 6766
rect -231 6732 -192 6766
rect -158 6732 -119 6766
rect -85 6732 -46 6766
rect -12 6732 27 6766
rect 61 6732 100 6766
rect 134 6732 173 6766
rect 207 6732 246 6766
rect 280 6732 319 6766
rect 353 6732 392 6766
rect 426 6732 465 6766
rect 499 6732 538 6766
rect 572 6732 611 6766
rect 645 6732 684 6766
rect 718 6732 757 6766
rect 791 6732 830 6766
rect 864 6732 903 6766
rect 937 6732 976 6766
rect 1010 6732 1049 6766
rect 1083 6732 1122 6766
rect 1156 6732 1195 6766
rect 1229 6732 1268 6766
rect 1302 6732 1341 6766
rect 1375 6732 1413 6766
rect 1447 6732 1485 6766
rect 1519 6732 1557 6766
rect 1591 6732 1629 6766
rect 1663 6732 1701 6766
rect 1735 6732 1773 6766
rect 1807 6732 1845 6766
rect 1879 6732 1917 6766
rect 1951 6732 1989 6766
rect 2023 6732 2061 6766
rect 2095 6732 2133 6766
rect 2167 6732 2205 6766
rect 2239 6732 2277 6766
rect 2311 6732 2349 6766
rect 2383 6732 2421 6766
rect 2455 6732 2493 6766
rect 2527 6732 2565 6766
rect 2599 6732 2637 6766
rect 2671 6732 2709 6766
rect 2743 6732 2781 6766
rect 2815 6732 2853 6766
rect 2887 6732 2925 6766
rect 2959 6732 2997 6766
rect 3031 6732 3069 6766
rect 3103 6732 3141 6766
rect 3175 6732 3213 6766
rect 3247 6732 3285 6766
rect 3319 6732 3357 6766
rect 3391 6732 3429 6766
rect 3463 6732 3501 6766
rect 3535 6732 3573 6766
rect 3607 6732 3645 6766
rect 3679 6732 3717 6766
rect 3751 6732 3789 6766
rect 3823 6732 3861 6766
rect 3895 6732 3933 6766
rect 3967 6732 4005 6766
rect 4039 6732 4077 6766
rect 4111 6732 4149 6766
rect -309 6694 4149 6732
rect -309 6660 -231 6694
rect -197 6660 -158 6694
rect -124 6660 -85 6694
rect -51 6660 -12 6694
rect 22 6660 61 6694
rect 95 6660 134 6694
rect 168 6660 207 6694
rect 241 6660 280 6694
rect 314 6660 353 6694
rect 387 6660 426 6694
rect 460 6660 499 6694
rect 533 6660 572 6694
rect 606 6660 645 6694
rect 679 6660 718 6694
rect 752 6660 791 6694
rect 825 6660 864 6694
rect 898 6660 937 6694
rect 971 6660 1010 6694
rect 1044 6660 1083 6694
rect 1117 6660 1156 6694
rect 1190 6660 1229 6694
rect 1263 6660 1302 6694
rect 1336 6660 1375 6694
rect 1409 6660 1448 6694
rect 1482 6660 1521 6694
rect 1555 6660 1594 6694
rect 1628 6660 1667 6694
rect 1701 6660 1740 6694
rect 1774 6660 1813 6694
rect 1847 6660 1886 6694
rect 1920 6660 1959 6694
rect 1993 6660 2032 6694
rect 2066 6660 2105 6694
rect 2139 6660 2178 6694
rect 2212 6660 2251 6694
rect 2285 6660 2324 6694
rect 2358 6660 2397 6694
rect 2431 6660 2470 6694
rect 2504 6660 2543 6694
rect 2577 6660 2616 6694
rect 2650 6660 2689 6694
rect 2723 6660 2762 6694
rect 2796 6660 2835 6694
rect 2869 6660 2908 6694
rect 2942 6660 2981 6694
rect 3015 6660 3054 6694
rect 3088 6660 3127 6694
rect 3161 6660 3200 6694
rect 3234 6660 3273 6694
rect 3307 6660 3346 6694
rect 3380 6660 3419 6694
rect 3453 6660 3492 6694
rect 3526 6660 3565 6694
rect 3599 6660 3638 6694
rect 3672 6660 3711 6694
rect 3745 6660 3784 6694
rect 3818 6660 3857 6694
rect 3891 6660 3930 6694
rect 3964 6660 4003 6694
rect 4037 6660 4076 6694
rect 4110 6660 4149 6694
rect 26143 6760 26293 6766
rect 26143 6726 26181 6760
rect 26215 6726 26253 6760
rect 26287 6726 26293 6760
rect 26143 6687 26293 6726
rect 26143 6660 26181 6687
rect -309 6656 26181 6660
rect -309 4102 -303 6656
rect -197 6654 26181 6656
rect -197 6653 -127 6654
tri -127 6653 -126 6654 nw
tri 1216 6653 1217 6654 ne
rect 1217 6653 1463 6654
tri 1463 6653 1464 6654 nw
tri 26124 6653 26125 6654 ne
rect 26125 6653 26181 6654
rect 26215 6653 26253 6687
rect 26287 6653 26293 6687
rect -197 6634 -146 6653
tri -146 6634 -127 6653 nw
tri 1217 6634 1236 6653 ne
rect 1236 6634 1444 6653
tri 1444 6634 1463 6653 nw
tri 26125 6634 26144 6653 ne
rect 26144 6634 26293 6653
rect -197 6622 -158 6634
tri -158 6622 -146 6634 nw
tri 1236 6622 1248 6634 ne
rect 1248 6622 1424 6634
rect -309 4068 -231 4102
rect -197 4068 -191 6622
tri -191 6589 -158 6622 nw
tri 1248 6589 1281 6622 ne
rect -21 6490 1077 6496
rect -21 6456 -9 6490
rect 25 6456 66 6490
rect 100 6456 141 6490
rect 175 6456 216 6490
rect 250 6456 291 6490
rect 325 6456 365 6490
rect 399 6456 439 6490
rect 473 6456 513 6490
rect 547 6456 587 6490
rect 621 6456 661 6490
rect 695 6456 735 6490
rect 769 6456 809 6490
rect 843 6456 883 6490
rect 917 6456 957 6490
rect 991 6456 1031 6490
rect 1065 6456 1077 6490
rect -21 6418 1077 6456
rect -21 6384 -9 6418
rect 25 6384 66 6418
rect 100 6384 141 6418
rect 175 6384 216 6418
rect 250 6384 291 6418
rect 325 6384 365 6418
rect 399 6384 439 6418
rect 473 6384 513 6418
rect 547 6384 587 6418
rect 621 6384 661 6418
rect 695 6384 735 6418
rect 769 6384 809 6418
rect 843 6384 883 6418
rect 917 6384 957 6418
rect 991 6384 1031 6418
rect 1065 6384 1077 6418
rect -21 6346 1077 6384
rect -21 6312 23 6346
rect 57 6312 98 6346
rect 132 6312 173 6346
rect 207 6312 248 6346
rect 282 6312 323 6346
rect 357 6312 398 6346
rect 432 6312 473 6346
rect 507 6312 548 6346
rect 582 6312 623 6346
rect 657 6312 698 6346
rect 732 6312 773 6346
rect 807 6312 848 6346
rect 882 6312 923 6346
rect 957 6312 1077 6346
rect -21 6308 1077 6312
rect -21 6274 1037 6308
rect 1071 6274 1077 6308
rect -21 6240 57 6274
rect 91 6240 133 6274
rect 167 6240 209 6274
rect 243 6240 285 6274
rect 319 6240 361 6274
rect 395 6240 437 6274
rect 471 6240 513 6274
rect 547 6240 589 6274
rect 623 6240 665 6274
rect 699 6240 740 6274
rect 774 6240 815 6274
rect 849 6240 890 6274
rect 924 6240 965 6274
rect 999 6240 1077 6274
rect -21 6234 1077 6240
rect -21 6200 -15 6234
rect 19 6233 161 6234
tri 161 6233 162 6234 nw
tri 894 6233 895 6234 ne
rect 895 6233 1077 6234
rect 19 6200 127 6233
rect -21 6199 127 6200
tri 127 6199 161 6233 nw
tri 895 6199 929 6233 ne
rect 929 6199 1037 6233
rect 1071 6199 1077 6233
rect -21 6198 126 6199
tri 126 6198 127 6199 nw
tri 929 6198 930 6199 ne
rect 930 6198 1077 6199
rect -21 6164 57 6198
rect 91 6164 97 6198
tri 97 6169 126 6198 nw
tri 930 6169 959 6198 ne
rect -21 6161 97 6164
rect -21 6127 -15 6161
rect 19 6127 97 6161
rect -21 6122 97 6127
rect -21 6088 57 6122
rect 91 6088 97 6122
rect 959 6164 965 6198
rect 999 6164 1077 6198
rect 959 6158 1077 6164
rect 959 6124 1037 6158
rect 1071 6124 1077 6158
rect 959 6122 1077 6124
rect 344 6114 826 6120
rect -21 6054 -15 6088
rect 19 6054 97 6088
rect -21 6046 97 6054
rect -21 6015 57 6046
rect -21 5981 -15 6015
rect 19 6012 57 6015
rect 91 6012 97 6046
rect 19 5981 97 6012
rect -21 5970 97 5981
rect -21 5942 57 5970
rect -21 5908 -15 5942
rect 19 5936 57 5942
rect 91 5936 97 5970
rect 19 5908 97 5936
rect -21 5894 97 5908
rect -21 5869 57 5894
rect -21 5835 -15 5869
rect 19 5860 57 5869
rect 91 5860 97 5894
rect 19 5835 97 5860
rect -21 5818 97 5835
rect -21 5795 57 5818
rect -21 5761 -15 5795
rect 19 5784 57 5795
rect 91 5784 97 5818
rect 19 5761 97 5784
rect -21 5742 97 5761
rect -21 5721 57 5742
rect -21 5687 -15 5721
rect 19 5708 57 5721
rect 91 5708 97 5742
rect 19 5687 97 5708
rect -21 5666 97 5687
rect -21 5647 57 5666
rect -21 5613 -15 5647
rect 19 5632 57 5647
rect 91 5632 97 5666
rect 19 5613 97 5632
rect -21 5590 97 5613
rect -21 5573 57 5590
rect -21 5539 -15 5573
rect 19 5556 57 5573
rect 91 5556 97 5590
rect 19 5539 97 5556
rect -21 5514 97 5539
rect -21 5499 57 5514
rect -21 5465 -15 5499
rect 19 5480 57 5499
rect 91 5480 97 5514
rect 19 5465 97 5480
rect -21 5437 97 5465
rect -21 5425 57 5437
rect -21 5391 -15 5425
rect 19 5403 57 5425
rect 91 5403 97 5437
rect 19 5391 97 5403
rect 211 5391 316 6097
rect 344 6080 356 6114
rect 390 6080 428 6114
rect 462 6080 500 6114
rect 534 6080 572 6114
rect 606 6080 644 6114
rect 678 6080 716 6114
rect 750 6088 826 6114
tri 826 6088 858 6120 sw
rect 959 6088 965 6122
rect 999 6088 1077 6122
rect 750 6083 858 6088
tri 858 6083 863 6088 sw
rect 959 6083 1077 6088
rect 750 6080 863 6083
rect 344 6074 863 6080
tri 863 6074 872 6083 sw
tri 806 6066 814 6074 ne
rect 814 6066 872 6074
tri 872 6066 880 6074 sw
tri 814 6054 826 6066 ne
rect 826 6054 880 6066
tri 826 6049 831 6054 ne
rect 831 6049 880 6054
tri 831 6046 834 6049 ne
rect -21 5360 97 5391
tri 239 5380 250 5391 ne
rect 250 5380 316 5391
tri 250 5366 264 5380 ne
rect -21 5351 57 5360
rect -21 5317 -15 5351
rect 19 5326 57 5351
rect 91 5326 97 5360
rect 19 5317 97 5326
rect -21 5283 97 5317
rect -21 5277 57 5283
rect -21 5243 -15 5277
rect 19 5249 57 5277
rect 91 5249 97 5283
rect 19 5243 97 5249
rect -21 5206 97 5243
rect -21 5203 57 5206
rect -21 5169 -15 5203
rect 19 5172 57 5203
rect 91 5172 97 5206
rect 19 5169 97 5172
rect -21 5129 97 5169
rect -21 5095 -15 5129
rect 19 5095 57 5129
rect 91 5095 97 5129
rect -21 4963 97 5095
tri 97 4963 100 4966 sw
rect -21 4929 100 4963
tri 100 4929 134 4963 sw
rect -21 4918 134 4929
tri 134 4918 145 4929 sw
tri -21 4908 -11 4918 ne
rect -11 4908 145 4918
tri 145 4908 155 4918 sw
tri -11 4890 7 4908 ne
rect 7 4890 155 4908
tri 155 4890 173 4908 sw
tri 7 4874 23 4890 ne
rect 23 4874 173 4890
tri 173 4874 189 4890 sw
tri 23 4856 41 4874 ne
rect 41 4856 189 4874
tri 41 4843 54 4856 ne
rect 54 4843 189 4856
tri 54 4835 62 4843 ne
rect 62 4835 189 4843
tri 62 4826 71 4835 ne
rect -309 4063 -191 4068
rect -309 4029 -303 4063
rect -269 4030 -191 4063
rect -269 4029 -231 4030
rect -309 3996 -231 4029
rect -197 3996 -191 4030
rect -309 3990 -191 3996
rect -309 3956 -303 3990
rect -269 3958 -191 3990
rect -269 3956 -231 3958
rect -309 3924 -231 3956
rect -197 3924 -191 3958
rect -309 3917 -191 3924
rect -309 3883 -303 3917
rect -269 3886 -191 3917
rect -269 3883 -231 3886
rect -309 3852 -231 3883
rect -197 3852 -191 3886
rect -309 3844 -191 3852
rect -309 3810 -303 3844
rect -269 3814 -191 3844
rect -269 3810 -231 3814
rect -309 3780 -231 3810
rect -197 3780 -191 3814
rect -309 3771 -191 3780
rect -309 3737 -303 3771
rect -269 3742 -191 3771
rect -269 3737 -231 3742
rect -309 3708 -231 3737
rect -197 3708 -191 3742
rect -309 3698 -191 3708
rect -309 3664 -303 3698
rect -269 3670 -191 3698
rect -269 3664 -231 3670
rect -309 3636 -231 3664
rect -197 3636 -191 3670
rect -309 3625 -191 3636
rect -309 3591 -303 3625
rect -269 3598 -191 3625
rect -269 3591 -231 3598
rect -309 3564 -231 3591
rect -197 3564 -191 3598
rect -309 3552 -191 3564
rect -309 3518 -303 3552
rect -269 3526 -191 3552
rect -269 3518 -231 3526
rect -309 3492 -231 3518
rect -197 3492 -191 3526
rect -309 3479 -191 3492
rect -309 3445 -303 3479
rect -269 3454 -191 3479
rect -269 3445 -231 3454
rect -309 3420 -231 3445
rect -197 3420 -191 3454
rect -309 3406 -191 3420
rect -309 3372 -303 3406
rect -269 3382 -191 3406
rect -269 3372 -231 3382
rect -309 3348 -231 3372
rect -197 3348 -191 3382
rect -309 3333 -191 3348
rect -309 3299 -303 3333
rect -269 3310 -191 3333
rect -269 3299 -231 3310
rect -309 3276 -231 3299
rect -197 3276 -191 3310
rect -309 3260 -191 3276
rect -309 3226 -303 3260
rect -269 3238 -191 3260
rect -269 3226 -231 3238
rect -309 3204 -231 3226
rect -197 3204 -191 3238
rect -309 3187 -191 3204
rect -309 3153 -303 3187
rect -269 3166 -191 3187
rect -269 3153 -231 3166
rect -309 3132 -231 3153
rect -197 3132 -191 3166
rect -309 3114 -191 3132
rect -309 3080 -303 3114
rect -269 3094 -191 3114
rect -269 3080 -231 3094
rect -309 3060 -231 3080
rect -197 3060 -191 3094
rect -309 3041 -191 3060
rect -309 3007 -303 3041
rect -269 3022 -191 3041
rect -269 3007 -231 3022
rect -309 2988 -231 3007
rect -197 2988 -191 3022
rect -309 2968 -191 2988
rect -309 2934 -303 2968
rect -269 2950 -191 2968
rect -269 2934 -231 2950
rect -309 2916 -231 2934
rect -197 2916 -191 2950
rect -309 2895 -191 2916
rect -309 2861 -303 2895
rect -269 2878 -191 2895
rect -269 2861 -231 2878
rect -309 2844 -231 2861
rect -197 2844 -191 2878
rect -309 2822 -191 2844
rect -309 2788 -303 2822
rect -269 2806 -191 2822
rect -269 2788 -231 2806
rect -309 2772 -231 2788
rect -197 2772 -191 2806
rect -309 2749 -191 2772
rect -309 2715 -303 2749
rect -269 2734 -191 2749
rect -269 2715 -231 2734
rect -309 2700 -231 2715
rect -197 2700 -191 2734
rect -309 2676 -191 2700
rect -309 2642 -303 2676
rect -269 2662 -191 2676
rect -269 2642 -231 2662
rect -309 2628 -231 2642
rect -197 2628 -191 2662
rect -309 2603 -191 2628
rect -309 2569 -303 2603
rect -269 2590 -191 2603
rect -269 2569 -231 2590
rect -309 2556 -231 2569
rect -197 2556 -191 2590
rect -309 2530 -191 2556
rect -309 2496 -303 2530
rect -269 2518 -191 2530
rect -269 2496 -231 2518
rect -309 2484 -231 2496
rect -197 2484 -191 2518
rect -309 2457 -191 2484
rect -309 2423 -303 2457
rect -269 2446 -191 2457
rect -269 2423 -231 2446
rect -309 2412 -231 2423
rect -197 2412 -191 2446
rect -309 2384 -191 2412
rect -309 2350 -303 2384
rect -269 2374 -191 2384
rect -269 2350 -231 2374
rect -309 2340 -231 2350
rect -197 2340 -191 2374
rect -309 2311 -191 2340
rect -309 2277 -303 2311
rect -269 2302 -191 2311
rect -269 2277 -231 2302
rect -309 2268 -231 2277
rect -197 2268 -191 2302
rect -309 2238 -191 2268
rect -309 2204 -303 2238
rect -269 2230 -191 2238
rect -269 2204 -231 2230
rect -309 2196 -231 2204
rect -197 2196 -191 2230
rect -309 2165 -191 2196
rect -309 2131 -303 2165
rect -269 2158 -191 2165
rect -269 2131 -231 2158
rect -309 2124 -231 2131
rect -197 2124 -191 2158
rect -309 2092 -191 2124
rect -309 2058 -303 2092
rect -269 2086 -191 2092
rect -269 2058 -231 2086
rect -309 2052 -231 2058
rect -197 2052 -191 2086
rect -309 2019 -191 2052
rect -309 1985 -303 2019
rect -269 2014 -191 2019
rect -269 1985 -231 2014
rect -309 1980 -231 1985
rect -197 1980 -191 2014
rect -309 1946 -191 1980
rect -309 1912 -303 1946
rect -269 1942 -191 1946
rect -269 1912 -231 1942
rect -309 1908 -231 1912
rect -197 1908 -191 1942
rect -309 1873 -191 1908
rect -309 1839 -303 1873
rect -269 1870 -191 1873
rect -269 1839 -231 1870
rect -309 1836 -231 1839
rect -197 1836 -191 1870
rect -309 1800 -191 1836
rect -309 1766 -303 1800
rect -269 1798 -191 1800
rect -269 1766 -231 1798
rect -309 1764 -231 1766
rect -197 1764 -191 1798
rect -309 1727 -191 1764
rect -309 1693 -303 1727
rect -269 1726 -191 1727
rect -269 1693 -231 1726
rect -309 1692 -231 1693
rect -197 1692 -191 1726
rect -309 1654 -191 1692
rect -309 1620 -303 1654
rect -269 1620 -231 1654
rect -197 1620 -191 1654
rect -309 1581 -191 1620
rect -309 1547 -303 1581
rect -269 1547 -231 1581
rect -197 1547 -191 1581
rect -309 1508 -191 1547
rect -309 1474 -303 1508
rect -269 1474 -231 1508
rect -197 1474 -191 1508
rect -309 1435 -191 1474
rect -309 1401 -303 1435
rect -269 1401 -231 1435
rect -197 1401 -191 1435
rect -309 1362 -191 1401
rect -309 1328 -303 1362
rect -269 1328 -231 1362
rect -197 1328 -191 1362
rect -309 1289 -191 1328
rect -309 1255 -303 1289
rect -269 1255 -231 1289
rect -197 1255 -191 1289
rect -309 1216 -191 1255
rect -309 1182 -303 1216
rect -269 1182 -231 1216
rect -197 1182 -191 1216
rect -309 1143 -191 1182
rect -309 1109 -303 1143
rect -269 1109 -231 1143
rect -197 1109 -191 1143
rect -309 1070 -191 1109
rect -309 1036 -303 1070
rect -269 1036 -231 1070
rect -197 1036 -191 1070
rect -309 997 -191 1036
rect -309 963 -303 997
rect -269 963 -231 997
rect -197 963 -191 997
rect -309 924 -191 963
rect -309 890 -303 924
rect -269 890 -231 924
rect -197 890 -191 924
rect -309 851 -191 890
rect -309 817 -303 851
rect -269 817 -231 851
rect -197 817 -191 851
rect -309 778 -191 817
rect -309 744 -303 778
rect -269 744 -231 778
rect -197 744 -191 778
rect -309 705 -191 744
rect -309 671 -303 705
rect -269 671 -231 705
rect -197 671 -191 705
rect -309 632 -191 671
rect -309 598 -303 632
rect -269 598 -231 632
rect -197 598 -191 632
rect -309 559 -191 598
rect -309 525 -303 559
rect -269 525 -231 559
rect -197 525 -191 559
rect -309 486 -191 525
rect -309 452 -303 486
rect -269 452 -231 486
rect -197 452 -191 486
rect -309 413 -191 452
rect -309 379 -303 413
rect -269 379 -231 413
rect -197 379 -191 413
rect -309 340 -191 379
rect -309 306 -303 340
rect -269 306 -231 340
rect -197 306 -191 340
rect -309 267 -191 306
rect -309 233 -303 267
rect -269 233 -231 267
rect -197 233 -191 267
rect -309 194 -191 233
rect -309 160 -303 194
rect -269 160 -231 194
rect -197 160 -191 194
rect -309 134 -191 160
rect 71 4596 189 4835
rect 71 2330 77 4596
rect 183 2330 189 4596
rect 71 2291 189 2330
rect 71 2257 77 2291
rect 111 2257 149 2291
rect 183 2257 189 2291
rect 71 2218 189 2257
rect 71 2184 77 2218
rect 111 2184 149 2218
rect 183 2184 189 2218
rect 71 2145 189 2184
rect 71 2111 77 2145
rect 111 2111 149 2145
rect 183 2111 189 2145
rect 71 2072 189 2111
rect 71 2038 77 2072
rect 111 2038 149 2072
rect 183 2038 189 2072
rect 71 1999 189 2038
rect 71 1965 77 1999
rect 111 1965 149 1999
rect 183 1965 189 1999
rect 71 1926 189 1965
rect 71 1892 77 1926
rect 111 1892 149 1926
rect 183 1892 189 1926
rect 71 1853 189 1892
rect 71 1819 77 1853
rect 111 1819 149 1853
rect 183 1819 189 1853
rect 71 1780 189 1819
rect 71 1746 77 1780
rect 111 1746 149 1780
rect 183 1746 189 1780
rect 71 1707 189 1746
rect 71 1673 77 1707
rect 111 1673 149 1707
rect 183 1673 189 1707
rect 71 1634 189 1673
rect 71 1600 77 1634
rect 111 1600 149 1634
rect 183 1600 189 1634
rect 71 1561 189 1600
rect 71 1527 77 1561
rect 111 1527 149 1561
rect 183 1527 189 1561
rect 71 1488 189 1527
rect 71 1454 77 1488
rect 111 1454 149 1488
rect 183 1454 189 1488
rect 71 1415 189 1454
rect 71 1381 77 1415
rect 111 1381 149 1415
rect 183 1381 189 1415
rect 71 1342 189 1381
rect 71 1308 77 1342
rect 111 1308 149 1342
rect 183 1308 189 1342
rect 71 1269 189 1308
rect 71 1235 77 1269
rect 111 1235 149 1269
rect 183 1235 189 1269
rect 71 1196 189 1235
rect 71 1162 77 1196
rect 111 1162 149 1196
rect 183 1162 189 1196
rect 71 1123 189 1162
rect 71 1089 77 1123
rect 111 1089 149 1123
rect 183 1089 189 1123
rect 71 1050 189 1089
rect 71 1016 77 1050
rect 111 1016 149 1050
rect 183 1016 189 1050
rect 71 977 189 1016
rect 71 943 77 977
rect 111 943 149 977
rect 183 943 189 977
rect 71 904 189 943
rect 71 870 77 904
rect 111 870 149 904
rect 183 870 189 904
rect 71 831 189 870
rect 71 797 77 831
rect 111 797 149 831
rect 183 797 189 831
rect 71 758 189 797
rect 71 724 77 758
rect 111 724 149 758
rect 183 724 189 758
rect 71 685 189 724
rect 71 651 77 685
rect 111 651 149 685
rect 183 651 189 685
rect 71 612 189 651
rect 71 578 77 612
rect 111 578 149 612
rect 183 578 189 612
rect 71 539 189 578
rect 71 505 77 539
rect 111 505 149 539
rect 183 505 189 539
rect 71 466 189 505
rect 71 432 77 466
rect 111 432 149 466
rect 183 432 189 466
rect 71 393 189 432
rect 71 359 77 393
rect 111 359 149 393
rect 183 359 189 393
rect 71 320 189 359
rect 71 286 77 320
rect 111 286 149 320
rect 183 286 189 320
rect 71 247 189 286
rect 71 213 77 247
rect 111 213 149 247
rect 183 213 189 247
rect 264 289 316 5380
rect 344 5958 762 5964
rect 344 5924 356 5958
rect 390 5924 428 5958
rect 462 5924 500 5958
rect 534 5924 572 5958
rect 606 5924 644 5958
rect 678 5924 716 5958
rect 750 5924 762 5958
rect 344 5918 762 5924
rect 344 5899 402 5918
tri 402 5899 421 5918 nw
rect 344 5895 398 5899
tri 398 5895 402 5899 nw
rect 344 3537 396 5895
tri 396 5893 398 5895 nw
tri 822 5824 834 5836 se
rect 834 5824 880 6049
tri 818 5820 822 5824 se
rect 822 5820 880 5824
tri 814 5816 818 5820 se
rect 818 5816 880 5820
tri 806 5808 814 5816 se
rect 814 5808 872 5816
tri 872 5808 880 5816 nw
rect 959 6049 1037 6083
rect 1071 6049 1077 6083
rect 959 6046 1077 6049
rect 959 6012 965 6046
rect 999 6012 1077 6046
rect 959 6008 1077 6012
rect 959 5974 1037 6008
rect 1071 5974 1077 6008
rect 959 5970 1077 5974
rect 959 5936 965 5970
rect 999 5936 1077 5970
rect 959 5933 1077 5936
rect 959 5899 1037 5933
rect 1071 5899 1077 5933
rect 959 5895 1077 5899
rect 959 5861 965 5895
rect 999 5861 1077 5895
rect 959 5858 1077 5861
rect 959 5824 1037 5858
rect 1071 5824 1077 5858
rect 959 5820 1077 5824
tri 493 5802 499 5808 se
rect 499 5802 850 5808
tri 459 5768 493 5802 se
rect 493 5768 512 5802
rect 546 5768 584 5802
rect 618 5768 656 5802
rect 690 5768 728 5802
rect 762 5786 850 5802
tri 850 5786 872 5808 nw
rect 959 5786 965 5820
rect 999 5786 1077 5820
rect 762 5783 847 5786
tri 847 5783 850 5786 nw
rect 959 5783 1077 5786
rect 762 5768 826 5783
tri 453 5762 459 5768 se
rect 459 5762 826 5768
tri 826 5762 847 5783 nw
tri 440 5749 453 5762 se
rect 453 5749 514 5762
tri 514 5749 527 5762 nw
rect 959 5749 1037 5783
rect 1071 5749 1077 5783
tri 436 5745 440 5749 se
rect 440 5745 510 5749
tri 510 5745 514 5749 nw
rect 959 5745 1077 5749
tri 424 5733 436 5745 se
rect 436 5733 476 5745
rect 424 3708 476 5733
tri 476 5711 510 5745 nw
rect 959 5711 965 5745
rect 999 5711 1077 5745
rect 959 5708 1077 5711
rect 504 5692 821 5698
rect 504 5658 516 5692
rect 550 5658 588 5692
rect 622 5658 660 5692
rect 694 5658 732 5692
rect 766 5674 821 5692
tri 821 5674 845 5698 sw
rect 959 5674 1037 5708
rect 1071 5674 1077 5708
rect 766 5670 845 5674
tri 845 5670 849 5674 sw
rect 959 5670 1077 5674
rect 766 5658 849 5670
rect 504 5655 849 5658
tri 849 5655 864 5670 sw
rect 504 5652 864 5655
tri 793 5636 809 5652 ne
rect 809 5636 864 5652
tri 809 5633 812 5636 ne
rect 812 5633 864 5636
tri 812 5627 818 5633 ne
rect 504 5536 778 5542
rect 504 5502 516 5536
rect 550 5502 588 5536
rect 622 5502 660 5536
rect 694 5502 732 5536
rect 766 5502 778 5536
rect 504 5496 778 5502
rect 504 5486 571 5496
tri 571 5486 581 5496 nw
rect 504 5484 569 5486
tri 569 5484 571 5486 nw
rect 504 3954 556 5484
tri 556 5471 569 5484 nw
tri 817 5410 818 5411 se
rect 818 5410 864 5633
tri 793 5386 817 5410 se
rect 817 5386 864 5410
rect 584 5383 864 5386
rect 584 5380 857 5383
rect 584 5346 596 5380
rect 630 5346 668 5380
rect 702 5346 740 5380
rect 774 5376 857 5380
tri 857 5376 864 5383 nw
rect 959 5636 965 5670
rect 999 5636 1077 5670
rect 959 5633 1077 5636
rect 959 5599 1037 5633
rect 1071 5599 1077 5633
rect 959 5595 1077 5599
rect 959 5561 965 5595
rect 999 5561 1077 5595
rect 959 5558 1077 5561
rect 959 5524 1037 5558
rect 1071 5524 1077 5558
rect 959 5520 1077 5524
rect 959 5486 965 5520
rect 999 5486 1077 5520
rect 959 5484 1077 5486
rect 959 5450 1037 5484
rect 1071 5450 1077 5484
rect 959 5445 1077 5450
rect 959 5411 965 5445
rect 999 5411 1077 5445
rect 959 5410 1077 5411
rect 959 5376 1037 5410
rect 1071 5376 1077 5410
rect 774 5370 851 5376
tri 851 5370 857 5376 nw
rect 959 5370 1077 5376
rect 774 5346 821 5370
rect 584 5340 821 5346
tri 821 5340 851 5370 nw
rect 584 5336 657 5340
tri 657 5336 661 5340 nw
rect 959 5336 965 5370
rect 999 5336 1077 5370
rect 584 4110 636 5336
tri 636 5315 657 5336 nw
rect 959 5302 1037 5336
rect 1071 5302 1077 5336
rect 959 5295 1077 5302
tri 929 5261 959 5291 se
rect 959 5261 965 5295
rect 999 5262 1077 5295
rect 999 5261 1037 5262
tri 896 5228 929 5261 se
rect 929 5228 1037 5261
rect 1071 5228 1077 5262
tri 894 5226 896 5228 se
rect 896 5226 1077 5228
rect 703 5220 1077 5226
rect 703 5186 715 5220
rect 749 5186 798 5220
rect 832 5186 881 5220
rect 915 5186 965 5220
rect 999 5186 1077 5220
rect 703 5148 1077 5186
rect 703 5114 715 5148
rect 749 5114 809 5148
rect 843 5114 904 5148
rect 938 5114 999 5148
rect 1033 5114 1077 5148
rect 703 4618 1077 5114
rect 1281 5148 1287 6622
rect 1393 6614 1424 6622
tri 1424 6614 1444 6634 nw
tri 26144 6614 26164 6634 ne
rect 26164 6614 26293 6634
rect 1393 6603 1413 6614
tri 1413 6603 1424 6614 nw
tri 26164 6603 26175 6614 ne
rect 1393 5148 1399 6603
tri 1399 6589 1413 6603 nw
rect 26175 6580 26181 6614
rect 26215 6580 26253 6614
rect 26287 6580 26293 6614
rect 26175 6541 26293 6580
rect 26175 6507 26181 6541
rect 26215 6507 26253 6541
rect 26287 6507 26293 6541
tri 1709 6473 1715 6479 se
rect 1715 6473 25586 6479
rect 1281 5109 1399 5148
rect 1281 5075 1287 5109
rect 1321 5075 1359 5109
rect 1393 5075 1399 5109
rect 1281 5036 1399 5075
rect 1281 5002 1287 5036
rect 1321 5002 1359 5036
rect 1393 5002 1399 5036
rect 1281 4963 1399 5002
rect 1281 4929 1287 4963
rect 1321 4929 1359 4963
rect 1393 4929 1399 4963
rect 1281 4890 1399 4929
rect 1281 4856 1287 4890
rect 1321 4856 1359 4890
rect 1393 4856 1399 4890
rect 1281 4844 1399 4856
tri 1603 6367 1709 6473 se
rect 1709 6367 1804 6473
rect 23006 6439 23045 6473
rect 23079 6439 23118 6473
rect 23152 6439 23191 6473
rect 23225 6439 23264 6473
rect 23298 6439 23337 6473
rect 23371 6439 23410 6473
rect 23444 6439 23483 6473
rect 23517 6439 23556 6473
rect 23590 6439 23629 6473
rect 23663 6439 23702 6473
rect 23736 6439 23775 6473
rect 23809 6439 23848 6473
rect 23882 6439 23921 6473
rect 23955 6439 23994 6473
rect 24028 6439 24067 6473
rect 24101 6439 24140 6473
rect 24174 6439 24213 6473
rect 24247 6439 24286 6473
rect 24320 6439 24359 6473
rect 24393 6439 24432 6473
rect 24466 6439 24505 6473
rect 24539 6439 24578 6473
rect 24612 6439 24651 6473
rect 24685 6439 24724 6473
rect 24758 6439 24797 6473
rect 24831 6439 24870 6473
rect 24904 6439 24943 6473
rect 24977 6439 25016 6473
rect 25050 6439 25089 6473
rect 25123 6439 25162 6473
rect 25196 6439 25235 6473
rect 25269 6439 25308 6473
rect 25342 6439 25381 6473
rect 25415 6439 25454 6473
rect 25488 6439 25527 6473
rect 25561 6468 25586 6473
tri 25586 6468 25597 6479 sw
rect 26175 6468 26293 6507
rect 25561 6439 25597 6468
rect 23006 6434 25597 6439
tri 25597 6434 25631 6468 sw
rect 26175 6434 26181 6468
rect 26215 6434 26253 6468
rect 26287 6434 26293 6468
rect 23006 6401 25631 6434
rect 23006 6367 23045 6401
rect 23079 6367 23118 6401
rect 23152 6367 23191 6401
rect 23225 6367 23264 6401
rect 23298 6367 23337 6401
rect 23371 6367 23410 6401
rect 23444 6367 23483 6401
rect 23517 6367 23556 6401
rect 23590 6367 23629 6401
rect 23663 6367 23702 6401
rect 23736 6367 23775 6401
rect 23809 6367 23848 6401
rect 23882 6367 23921 6401
rect 23955 6367 23994 6401
rect 24028 6367 24067 6401
rect 24101 6367 24140 6401
rect 24174 6367 24213 6401
rect 24247 6367 24286 6401
rect 24320 6367 24359 6401
rect 24393 6367 24432 6401
rect 24466 6367 24505 6401
rect 24539 6367 24578 6401
rect 24612 6367 24651 6401
rect 24685 6367 24724 6401
rect 24758 6367 24797 6401
rect 24831 6367 24870 6401
rect 24904 6367 24943 6401
rect 24977 6367 25016 6401
rect 25050 6367 25089 6401
rect 25123 6367 25162 6401
rect 25196 6367 25235 6401
rect 25269 6367 25308 6401
rect 25342 6367 25381 6401
rect 25415 6367 25454 6401
rect 25488 6367 25527 6401
rect 25561 6395 25631 6401
tri 25631 6395 25670 6434 sw
rect 26175 6395 26293 6434
rect 25561 6367 25670 6395
rect 1603 6361 25670 6367
tri 25670 6361 25704 6395 sw
rect 26175 6361 26181 6395
rect 26215 6361 26253 6395
rect 26287 6361 26293 6395
rect 1603 6352 1887 6361
tri 1887 6352 1896 6361 nw
tri 25538 6352 25547 6361 ne
rect 25547 6352 25704 6361
rect 1603 6333 1868 6352
tri 1868 6333 1887 6352 nw
tri 25547 6333 25566 6352 ne
rect 25566 6333 25704 6352
rect 1603 6322 1857 6333
tri 1857 6322 1868 6333 nw
tri 2096 6322 2107 6333 se
rect 2107 6322 25420 6333
tri 25420 6322 25431 6333 sw
tri 25566 6322 25577 6333 ne
rect 25577 6322 25704 6333
tri 25704 6322 25743 6361 sw
rect 26175 6322 26293 6361
rect 1603 6315 1850 6322
tri 1850 6315 1857 6322 nw
tri 2089 6315 2096 6322 se
rect 2096 6315 25431 6322
tri 25431 6315 25438 6322 sw
tri 25577 6315 25584 6322 ne
rect 25584 6315 25743 6322
rect 1603 6306 1841 6315
tri 1841 6306 1850 6315 nw
tri 2080 6306 2089 6315 se
rect 2089 6306 25438 6315
tri 25438 6306 25447 6315 sw
tri 25584 6306 25593 6315 ne
rect 25593 6306 25743 6315
rect 1603 6294 1823 6306
rect 1603 6260 1609 6294
rect 1643 6260 1681 6294
rect 1715 6288 1823 6294
tri 1823 6288 1841 6306 nw
tri 2062 6288 2080 6306 se
rect 2080 6288 25447 6306
tri 25447 6288 25465 6306 sw
tri 25593 6288 25611 6306 ne
rect 25611 6288 25743 6306
tri 25743 6288 25777 6322 sw
rect 26175 6288 26181 6322
rect 26215 6288 26253 6322
rect 26287 6288 26293 6322
rect 1715 6260 1794 6288
rect 1603 6259 1794 6260
tri 1794 6259 1823 6288 nw
tri 2033 6259 2062 6288 se
rect 2062 6281 25465 6288
rect 2062 6259 2107 6281
tri 2107 6259 2129 6281 nw
tri 25398 6259 25420 6281 ne
rect 25420 6259 25465 6281
rect 1603 6249 1784 6259
tri 1784 6249 1794 6259 nw
tri 2023 6249 2033 6259 se
rect 2033 6253 2101 6259
tri 2101 6253 2107 6259 nw
tri 25420 6253 25426 6259 ne
rect 25426 6253 25465 6259
rect 2033 6249 2097 6253
tri 2097 6249 2101 6253 nw
tri 2137 6249 2141 6253 se
rect 2141 6249 25386 6253
tri 25386 6249 25390 6253 sw
tri 25426 6249 25430 6253 ne
rect 25430 6249 25465 6253
tri 25465 6249 25504 6288 sw
tri 25611 6249 25650 6288 ne
rect 25650 6279 25777 6288
tri 25777 6279 25786 6288 sw
rect 25650 6249 25786 6279
tri 25786 6249 25816 6279 sw
rect 26175 6249 26293 6288
rect 1603 6241 1776 6249
tri 1776 6241 1784 6249 nw
tri 2015 6241 2023 6249 se
rect 2023 6241 2089 6249
tri 2089 6241 2097 6249 nw
tri 2129 6241 2137 6249 se
rect 2137 6247 25390 6249
tri 25390 6247 25392 6249 sw
tri 25430 6247 25432 6249 ne
rect 25432 6247 25504 6249
rect 2137 6241 25392 6247
tri 25392 6241 25398 6247 sw
tri 25432 6241 25438 6247 ne
rect 25438 6241 25504 6247
tri 25504 6241 25512 6249 sw
tri 25650 6241 25658 6249 ne
rect 25658 6241 25816 6249
rect 1603 6240 1775 6241
tri 1775 6240 1776 6241 nw
tri 2014 6240 2015 6241 se
rect 2015 6240 2067 6241
rect 1603 6222 1750 6240
rect 1603 6220 1681 6222
rect 1603 6186 1609 6220
rect 1643 6188 1681 6220
rect 1715 6215 1750 6222
tri 1750 6215 1775 6240 nw
tri 1989 6215 2014 6240 se
rect 2014 6219 2067 6240
tri 2067 6219 2089 6241 nw
tri 2107 6219 2129 6241 se
rect 2129 6219 25398 6241
rect 2014 6215 2063 6219
tri 2063 6215 2067 6219 nw
tri 2103 6215 2107 6219 se
rect 2107 6215 25398 6219
tri 25398 6215 25424 6241 sw
tri 25438 6215 25464 6241 ne
rect 25464 6215 25512 6241
tri 25512 6215 25538 6241 sw
tri 25658 6215 25684 6241 ne
rect 25684 6215 25816 6241
tri 25816 6215 25850 6249 sw
rect 26175 6215 26181 6249
rect 26215 6215 26253 6249
rect 26287 6215 26293 6249
rect 1715 6188 1721 6215
rect 1643 6186 1721 6188
tri 1721 6186 1750 6215 nw
tri 1960 6186 1989 6215 se
rect 1989 6186 2033 6215
rect 1603 6149 1721 6186
tri 1959 6185 1960 6186 se
rect 1960 6185 2033 6186
tri 2033 6185 2063 6215 nw
tri 2095 6207 2103 6215 se
rect 2103 6207 25424 6215
tri 25424 6207 25432 6215 sw
tri 25464 6207 25472 6215 ne
rect 25472 6207 25538 6215
tri 2073 6185 2095 6207 se
rect 2095 6201 25432 6207
rect 2095 6185 2141 6201
tri 1956 6182 1959 6185 se
rect 1959 6182 2027 6185
tri 1950 6176 1956 6182 se
rect 1956 6179 2027 6182
tri 2027 6179 2033 6185 nw
tri 2067 6179 2073 6185 se
rect 2073 6179 2141 6185
tri 2141 6179 2163 6201 nw
tri 25364 6179 25386 6201 ne
rect 25386 6185 25432 6201
tri 25432 6185 25454 6207 sw
tri 25472 6185 25494 6207 ne
rect 25494 6195 25538 6207
tri 25538 6195 25558 6215 sw
tri 25684 6195 25704 6215 ne
rect 25704 6195 25850 6215
tri 25850 6195 25870 6215 sw
rect 25494 6185 25558 6195
rect 25386 6179 25454 6185
rect 1956 6176 2024 6179
tri 2024 6176 2027 6179 nw
tri 2064 6176 2067 6179 se
rect 2067 6176 2138 6179
tri 2138 6176 2141 6179 nw
tri 25386 6176 25389 6179 ne
rect 25389 6176 25454 6179
tri 25454 6176 25463 6185 sw
tri 25494 6176 25503 6185 ne
rect 25503 6176 25558 6185
tri 25558 6176 25577 6195 sw
tri 25704 6176 25723 6195 ne
rect 25723 6176 25870 6195
tri 25870 6176 25889 6195 sw
rect 26175 6176 26293 6215
tri 1941 6167 1950 6176 se
rect 1950 6167 2015 6176
tri 2015 6167 2024 6176 nw
tri 2055 6167 2064 6176 se
rect 2064 6173 2135 6176
tri 2135 6173 2138 6176 nw
tri 25389 6173 25392 6176 ne
rect 25392 6173 25463 6176
tri 25463 6173 25466 6176 sw
tri 25503 6173 25506 6176 ne
rect 25506 6173 25577 6176
rect 2064 6167 2104 6173
rect 1603 6146 1681 6149
rect 1603 6112 1609 6146
rect 1643 6115 1681 6146
rect 1715 6115 1721 6149
tri 1916 6142 1941 6167 se
rect 1941 6145 1993 6167
tri 1993 6145 2015 6167 nw
tri 2033 6145 2055 6167 se
rect 2055 6145 2104 6167
rect 1941 6142 1990 6145
tri 1990 6142 1993 6145 nw
tri 2030 6142 2033 6145 se
rect 2033 6142 2104 6145
tri 2104 6142 2135 6173 nw
tri 2144 6142 2175 6173 se
rect 2175 6142 25352 6173
tri 25352 6142 25383 6173 sw
tri 25392 6142 25423 6173 ne
rect 25423 6167 25466 6173
tri 25466 6167 25472 6173 sw
tri 25506 6167 25512 6173 ne
rect 25512 6167 25577 6173
tri 25577 6167 25586 6176 sw
tri 25723 6167 25732 6176 ne
rect 25732 6167 25889 6176
rect 25423 6142 25472 6167
tri 25472 6142 25497 6167 sw
tri 25512 6142 25537 6167 ne
rect 25537 6142 25586 6167
tri 25586 6142 25611 6167 sw
tri 25732 6145 25754 6167 ne
rect 25754 6161 25889 6167
tri 25889 6161 25904 6176 sw
rect 25754 6145 25904 6161
tri 25754 6142 25757 6145 ne
rect 25757 6142 25904 6145
tri 1907 6133 1916 6142 se
rect 1916 6133 1981 6142
tri 1981 6133 1990 6142 nw
tri 2021 6133 2030 6142 se
rect 2030 6139 2101 6142
tri 2101 6139 2104 6142 nw
tri 2141 6139 2144 6142 se
rect 2144 6139 25383 6142
tri 25383 6139 25386 6142 sw
tri 25423 6139 25426 6142 ne
rect 25426 6139 25497 6142
rect 2030 6133 2095 6139
tri 2095 6133 2101 6139 nw
tri 2135 6133 2141 6139 se
rect 2141 6133 25386 6139
tri 25386 6133 25392 6139 sw
tri 25426 6133 25432 6139 ne
rect 25432 6133 25497 6139
tri 25497 6133 25506 6142 sw
tri 25537 6133 25546 6142 ne
rect 25546 6133 25611 6142
tri 25611 6133 25620 6142 sw
tri 25757 6133 25766 6142 ne
rect 25766 6133 25904 6142
rect 1643 6112 1721 6115
rect 1603 6076 1721 6112
tri 1885 6111 1907 6133 se
rect 1907 6111 1959 6133
tri 1959 6111 1981 6133 nw
tri 1999 6111 2021 6133 se
rect 2021 6111 2067 6133
tri 1867 6093 1885 6111 se
rect 1885 6105 1953 6111
tri 1953 6105 1959 6111 nw
tri 1993 6105 1999 6111 se
rect 1999 6105 2067 6111
tri 2067 6105 2095 6133 nw
tri 2107 6105 2135 6133 se
rect 2135 6121 25392 6133
rect 2135 6105 2175 6121
rect 1885 6093 1941 6105
tri 1941 6093 1953 6105 nw
tri 1981 6093 1993 6105 se
rect 1993 6099 2061 6105
tri 2061 6099 2067 6105 nw
tri 2101 6099 2107 6105 se
rect 2107 6099 2175 6105
tri 2175 6099 2197 6121 nw
tri 25330 6099 25352 6121 ne
rect 25352 6105 25392 6121
tri 25392 6105 25420 6133 sw
tri 25432 6105 25460 6133 ne
rect 25460 6111 25506 6133
tri 25506 6111 25528 6133 sw
tri 25546 6111 25568 6133 ne
rect 25568 6111 25620 6133
rect 25460 6105 25528 6111
rect 25352 6099 25420 6105
tri 25420 6099 25426 6105 sw
tri 25460 6099 25466 6105 ne
rect 25466 6099 25528 6105
tri 25528 6099 25540 6111 sw
tri 25568 6099 25580 6111 ne
rect 25580 6099 25620 6111
rect 1993 6093 2027 6099
rect 1603 6072 1681 6076
rect 1603 6038 1609 6072
rect 1643 6042 1681 6072
rect 1715 6042 1721 6076
rect 1643 6038 1721 6042
rect 1603 6003 1721 6038
rect 1603 5998 1681 6003
rect 1603 5964 1609 5998
rect 1643 5969 1681 5998
rect 1715 5969 1721 6003
rect 1643 5964 1721 5969
rect 1603 5930 1721 5964
rect 1603 5924 1681 5930
rect 1603 5890 1609 5924
rect 1643 5896 1681 5924
rect 1715 5896 1721 5930
rect 1643 5890 1721 5896
rect 1603 5857 1721 5890
rect 1603 5850 1681 5857
rect 1603 5816 1609 5850
rect 1643 5823 1681 5850
rect 1715 5823 1721 5857
rect 1643 5816 1721 5823
rect 1603 5784 1721 5816
rect 1603 5776 1681 5784
rect 1603 5742 1609 5776
rect 1643 5750 1681 5776
rect 1715 5750 1721 5784
rect 1643 5742 1721 5750
rect 1603 5711 1721 5742
rect 1603 5702 1681 5711
rect 1603 5668 1609 5702
rect 1643 5677 1681 5702
rect 1715 5677 1721 5711
rect 1643 5668 1721 5677
rect 1603 5638 1721 5668
rect 1603 5627 1681 5638
rect 1603 5593 1609 5627
rect 1643 5604 1681 5627
rect 1715 5604 1721 5638
rect 1643 5593 1721 5604
rect 1603 5565 1721 5593
rect 1603 5552 1681 5565
rect 1603 5518 1609 5552
rect 1643 5531 1681 5552
rect 1715 5531 1721 5565
rect 1643 5518 1721 5531
rect 1603 5492 1721 5518
rect 1603 5477 1681 5492
rect 1603 5443 1609 5477
rect 1643 5458 1681 5477
rect 1715 5458 1721 5492
rect 1643 5443 1721 5458
rect 1603 5419 1721 5443
rect 1603 5402 1681 5419
rect 1603 5368 1609 5402
rect 1643 5385 1681 5402
rect 1715 5385 1721 5419
rect 1643 5368 1721 5385
rect 1603 5346 1721 5368
rect 1603 5327 1681 5346
rect 1603 5293 1609 5327
rect 1643 5312 1681 5327
rect 1715 5312 1721 5346
rect 1643 5293 1721 5312
rect 1603 5273 1721 5293
rect 1603 5252 1681 5273
rect 1603 5218 1609 5252
rect 1643 5239 1681 5252
rect 1715 5239 1721 5273
rect 1643 5218 1721 5239
rect 1603 5200 1721 5218
rect 1603 5177 1681 5200
rect 1603 5143 1609 5177
rect 1643 5166 1681 5177
rect 1715 5166 1721 5200
rect 1643 5143 1721 5166
rect 1603 5127 1721 5143
rect 1603 5102 1681 5127
rect 1603 5068 1609 5102
rect 1643 5093 1681 5102
rect 1715 5093 1721 5127
rect 1643 5068 1721 5093
rect 1603 5054 1721 5068
rect 1603 5027 1681 5054
rect 1603 4993 1609 5027
rect 1643 5020 1681 5027
rect 1715 5020 1721 5054
rect 1643 4993 1721 5020
rect 1603 4981 1721 4993
rect 1603 4952 1681 4981
rect 1603 4918 1609 4952
rect 1643 4947 1681 4952
rect 1715 4947 1721 4981
rect 1643 4918 1721 4947
rect 1603 4908 1721 4918
rect 1603 4877 1681 4908
rect 1603 4843 1609 4877
rect 1643 4874 1681 4877
rect 1715 4874 1721 4908
rect 1643 4843 1721 4874
rect 1603 4835 1721 4843
rect 1603 4802 1681 4835
rect 1603 4768 1609 4802
rect 1643 4801 1681 4802
rect 1715 4801 1721 4835
rect 1643 4768 1721 4801
rect 1603 4762 1721 4768
rect 1603 4728 1681 4762
rect 1715 4728 1721 4762
rect 1603 4727 1721 4728
rect 1603 4693 1609 4727
rect 1643 4693 1721 4727
rect 1603 4689 1721 4693
rect 1603 4655 1681 4689
rect 1715 4655 1721 4689
rect 1603 4652 1721 4655
tri 1077 4618 1107 4648 sw
tri 1573 4618 1603 4648 se
rect 1603 4618 1609 4652
rect 1643 4618 1721 4652
rect 703 4616 1107 4618
tri 1107 4616 1109 4618 sw
tri 1571 4616 1573 4618 se
rect 1573 4616 1721 4618
rect 703 4583 1109 4616
tri 1109 4583 1142 4616 sw
tri 1538 4583 1571 4616 se
rect 1571 4583 1681 4616
rect 703 4582 1681 4583
rect 1715 4582 1721 4616
rect 703 4577 1721 4582
rect 703 4543 740 4577
rect 774 4543 813 4577
rect 847 4543 886 4577
rect 920 4543 959 4577
rect 993 4543 1032 4577
rect 1066 4543 1105 4577
rect 1139 4543 1177 4577
rect 1211 4543 1249 4577
rect 1283 4543 1321 4577
rect 1355 4543 1393 4577
rect 1427 4543 1465 4577
rect 1499 4543 1537 4577
rect 1571 4543 1609 4577
rect 1643 4543 1721 4577
rect 703 4509 1681 4543
rect 1715 4509 1721 4543
rect 703 4505 1721 4509
rect 703 4471 740 4505
rect 774 4471 815 4505
rect 849 4471 890 4505
rect 924 4471 965 4505
rect 999 4471 1040 4505
rect 1074 4471 1115 4505
rect 1149 4471 1190 4505
rect 1224 4471 1265 4505
rect 1299 4471 1340 4505
rect 1374 4471 1415 4505
rect 1449 4471 1490 4505
rect 1524 4471 1565 4505
rect 1599 4471 1721 4505
rect 703 4465 1721 4471
tri 1815 6041 1867 6093 se
rect 1867 6071 1919 6093
tri 1919 6071 1941 6093 nw
tri 1959 6071 1981 6093 se
rect 1981 6071 2027 6093
rect 1867 6041 1889 6071
tri 1889 6041 1919 6071 nw
tri 1947 6059 1959 6071 se
rect 1959 6065 2027 6071
tri 2027 6065 2061 6099 nw
tri 2067 6065 2101 6099 se
rect 2101 6093 2169 6099
tri 2169 6093 2175 6099 nw
tri 25352 6093 25358 6099 ne
rect 25358 6093 25426 6099
rect 2101 6065 2129 6093
rect 1959 6059 2021 6065
tri 2021 6059 2027 6065 nw
tri 2061 6059 2067 6065 se
rect 2067 6059 2129 6065
tri 1929 6041 1947 6059 se
rect 1947 6041 1993 6059
rect 717 4226 1733 4232
rect 717 4192 729 4226
rect 763 4192 803 4226
rect 837 4192 877 4226
rect 911 4192 951 4226
rect 985 4192 1025 4226
rect 1059 4192 1099 4226
rect 1133 4192 1173 4226
rect 1207 4192 1247 4226
rect 1281 4192 1321 4226
rect 1355 4192 1395 4226
rect 1429 4192 1468 4226
rect 1502 4192 1541 4226
rect 1575 4192 1614 4226
rect 1648 4192 1687 4226
rect 1721 4192 1733 4226
rect 717 4186 1733 4192
tri 636 4110 661 4135 sw
tri 1790 4110 1815 4135 se
rect 1815 4110 1867 6041
tri 1867 6019 1889 6041 nw
tri 1919 6031 1929 6041 se
rect 1929 6031 1993 6041
tri 1993 6031 2021 6059 nw
tri 2033 6031 2061 6059 se
rect 2061 6053 2129 6059
tri 2129 6053 2169 6093 nw
tri 2181 6065 2209 6093 se
rect 2209 6065 25318 6093
tri 25318 6065 25346 6093 sw
tri 25358 6065 25386 6093 ne
rect 25386 6065 25426 6093
tri 25426 6065 25460 6099 sw
tri 25466 6065 25500 6099 ne
rect 25500 6093 25540 6099
tri 25540 6093 25546 6099 sw
tri 25580 6093 25586 6099 ne
rect 25586 6093 25620 6099
tri 25620 6093 25660 6133 sw
tri 25766 6113 25786 6133 ne
rect 25500 6065 25546 6093
tri 2169 6053 2181 6065 se
rect 2181 6053 25346 6065
rect 2061 6035 2111 6053
tri 2111 6035 2129 6053 nw
tri 2151 6035 2169 6053 se
rect 2169 6041 25346 6053
rect 2169 6035 2209 6041
rect 2061 6031 2101 6035
tri 1907 6019 1919 6031 se
rect 1919 6019 1969 6031
rect 584 4103 1860 4110
tri 1860 4103 1867 4110 nw
tri 1895 6007 1907 6019 se
rect 1907 6007 1969 6019
tri 1969 6007 1993 6031 nw
tri 2027 6025 2033 6031 se
rect 2033 6025 2101 6031
tri 2101 6025 2111 6035 nw
tri 2141 6025 2151 6035 se
rect 2151 6025 2209 6035
tri 2009 6007 2027 6025 se
rect 2027 6007 2082 6025
rect 584 4078 1835 4103
tri 1835 4078 1860 4103 nw
rect 584 4071 1828 4078
tri 1828 4071 1835 4078 nw
rect 584 4065 1822 4071
tri 1822 4065 1828 4071 nw
tri 1889 4065 1895 4071 se
rect 1895 4065 1947 6007
tri 1947 5985 1969 6007 nw
tri 2008 6006 2009 6007 se
rect 2009 6006 2082 6007
tri 2082 6006 2101 6025 nw
tri 2122 6006 2141 6025 se
rect 2141 6006 2209 6025
rect 2008 5985 2061 6006
tri 2061 5985 2082 6006 nw
tri 2111 5995 2122 6006 se
rect 2122 5995 2209 6006
tri 2209 5995 2255 6041 nw
tri 25296 6013 25324 6041 ne
rect 25324 6031 25346 6041
tri 25346 6031 25380 6065 sw
tri 25386 6031 25420 6065 ne
rect 25420 6059 25460 6065
tri 25460 6059 25466 6065 sw
tri 25500 6059 25506 6065 ne
rect 25506 6059 25546 6065
tri 25546 6059 25580 6093 sw
tri 25586 6059 25620 6093 ne
rect 25620 6059 25660 6093
rect 25420 6031 25466 6059
tri 25466 6031 25494 6059 sw
tri 25506 6031 25534 6059 ne
rect 25534 6041 25580 6059
tri 25580 6041 25598 6059 sw
tri 25620 6041 25638 6059 ne
rect 25638 6041 25660 6059
rect 25534 6031 25598 6041
rect 25324 6025 25380 6031
tri 25380 6025 25386 6031 sw
tri 25420 6025 25426 6031 ne
rect 25426 6025 25494 6031
tri 25494 6025 25500 6031 sw
tri 25534 6025 25540 6031 ne
rect 25540 6025 25598 6031
tri 25598 6025 25614 6041 sw
tri 25638 6025 25654 6041 ne
rect 25654 6025 25660 6041
rect 25324 6013 25386 6025
tri 25386 6013 25398 6025 sw
tri 25426 6013 25438 6025 ne
rect 25438 6013 25500 6025
tri 4283 5995 4301 6013 se
rect 4301 5995 25283 6013
tri 25283 5995 25301 6013 sw
tri 25324 5995 25342 6013 ne
rect 25342 6006 25398 6013
tri 25398 6006 25405 6013 sw
tri 25438 6006 25445 6013 ne
rect 25445 6007 25500 6013
tri 25500 6007 25518 6025 sw
tri 25540 6007 25558 6025 ne
rect 25558 6019 25614 6025
tri 25614 6019 25620 6025 sw
tri 25654 6019 25660 6025 ne
tri 25660 6019 25734 6093 sw
rect 25558 6007 25620 6019
rect 25445 6006 25518 6007
rect 25342 5997 25405 6006
tri 25405 5997 25414 6006 sw
tri 25445 5997 25454 6006 ne
rect 25454 5997 25518 6006
rect 25342 5995 25414 5997
tri 2107 5991 2111 5995 se
rect 2111 5991 2205 5995
tri 2205 5991 2209 5995 nw
tri 4279 5991 4283 5995 se
rect 4283 5991 25301 5995
tri 25301 5991 25305 5995 sw
tri 25342 5991 25346 5995 ne
rect 25346 5991 25414 5995
tri 25414 5991 25420 5997 sw
tri 25454 5991 25460 5997 ne
rect 25460 5991 25518 5997
tri 25518 5991 25534 6007 sw
tri 25558 5991 25574 6007 ne
rect 25574 5997 25620 6007
tri 25620 5997 25642 6019 sw
tri 25660 5997 25682 6019 ne
rect 25574 5991 25642 5997
tri 2101 5985 2107 5991 se
rect 2107 5985 2199 5991
tri 2199 5985 2205 5991 nw
tri 4273 5985 4279 5991 se
rect 4279 5985 25305 5991
rect 584 4064 1821 4065
tri 1821 4064 1822 4065 nw
tri 1888 4064 1889 4065 se
rect 1889 4064 1947 4065
rect 584 4052 1809 4064
tri 1809 4052 1821 4064 nw
tri 1876 4052 1888 4064 se
rect 1888 4052 1947 4064
tri 958 4031 979 4052 ne
rect 979 4031 1045 4052
tri 1045 4031 1066 4052 nw
tri 1855 4031 1876 4052 se
rect 1876 4049 1947 4052
rect 1876 4031 1929 4049
tri 1929 4031 1947 4049 nw
tri 979 4027 983 4031 ne
tri 556 3954 581 3979 sw
rect 504 3942 955 3954
rect 504 3908 555 3942
rect 589 3908 627 3942
rect 661 3908 699 3942
rect 733 3908 771 3942
rect 805 3908 843 3942
rect 877 3908 915 3942
rect 949 3908 955 3942
rect 504 3896 955 3908
tri 974 3814 983 3823 se
rect 983 3814 1041 4031
tri 1041 4027 1045 4031 nw
tri 1851 4027 1855 4031 se
rect 1855 4027 1917 4031
tri 1843 4019 1851 4027 se
rect 1851 4019 1917 4027
tri 1917 4019 1929 4031 nw
tri 1840 4016 1843 4019 se
rect 1843 4016 1914 4019
tri 1914 4016 1917 4019 nw
tri 1821 3997 1840 4016 se
rect 1840 3997 1895 4016
tri 1895 3997 1914 4016 nw
tri 1778 3954 1821 3997 se
rect 1821 3954 1852 3997
tri 1852 3954 1895 3997 nw
rect 1069 3948 1846 3954
tri 1846 3948 1852 3954 nw
rect 1069 3942 1840 3948
tri 1840 3942 1846 3948 nw
rect 1069 3908 1075 3942
rect 1109 3908 1147 3942
rect 1181 3908 1219 3942
rect 1253 3908 1291 3942
rect 1325 3908 1363 3942
rect 1397 3908 1435 3942
rect 1469 3908 1806 3942
tri 1806 3908 1840 3942 nw
rect 1069 3896 1794 3908
tri 1794 3896 1806 3908 nw
tri 1041 3814 1050 3823 sw
tri 958 3798 974 3814 se
rect 974 3798 1050 3814
tri 1050 3798 1066 3814 sw
rect 932 3780 1861 3798
rect 932 3746 1671 3780
rect 1705 3746 1743 3780
rect 1777 3746 1815 3780
rect 1849 3746 1861 3780
rect 932 3740 1861 3746
tri 476 3708 481 3713 sw
rect 424 3698 481 3708
tri 481 3698 491 3708 sw
rect 424 3688 491 3698
tri 491 3688 501 3698 sw
tri 1998 3688 2008 3698 se
rect 2008 3688 2060 5985
tri 2060 5984 2061 5985 nw
tri 2100 5984 2101 5985 se
rect 2101 5984 2196 5985
rect 424 3676 1092 3688
tri 424 3670 430 3676 ne
rect 430 3670 1092 3676
tri 1980 3670 1998 3688 se
rect 1998 3676 2060 3688
rect 1998 3670 2054 3676
tri 2054 3670 2060 3676 nw
tri 2088 5972 2100 5984 se
rect 2100 5982 2196 5984
tri 2196 5982 2199 5985 nw
tri 2315 5982 2318 5985 se
rect 2318 5982 3814 5985
rect 2100 5972 2186 5982
tri 2186 5972 2196 5982 nw
tri 2305 5972 2315 5982 se
rect 2315 5972 3814 5982
tri 4260 5972 4273 5985 se
rect 4273 5972 25305 5985
tri 25305 5972 25324 5991 sw
tri 25346 5972 25365 5991 ne
rect 25365 5985 25420 5991
tri 25420 5985 25426 5991 sw
tri 25460 5985 25466 5991 ne
rect 25466 5985 25534 5991
tri 25534 5985 25540 5991 sw
tri 25574 5985 25580 5991 ne
rect 25580 5985 25642 5991
tri 25642 5985 25654 5997 sw
rect 25365 5984 25426 5985
tri 25426 5984 25427 5985 sw
tri 25466 5984 25467 5985 ne
rect 25467 5984 25540 5985
rect 25365 5972 25427 5984
tri 430 3636 464 3670 ne
rect 464 3636 1092 3670
tri 1946 3636 1980 3670 se
rect 1980 3636 2020 3670
tri 2020 3636 2054 3670 nw
tri 464 3632 468 3636 ne
rect 468 3632 1092 3636
tri 1942 3632 1946 3636 se
rect 1946 3632 2016 3636
tri 2016 3632 2020 3636 nw
tri 468 3630 470 3632 ne
rect 470 3630 1092 3632
tri 1940 3630 1942 3632 se
rect 1942 3630 2014 3632
tri 2014 3630 2016 3632 nw
tri 958 3620 968 3630 ne
rect 968 3626 1062 3630
tri 1062 3626 1066 3630 nw
tri 1936 3626 1940 3630 se
rect 1940 3626 2010 3630
tri 2010 3626 2014 3630 nw
tri 2084 3626 2088 3630 se
rect 2088 3626 2140 5972
tri 2140 5926 2186 5972 nw
tri 2259 5926 2305 5972 se
rect 2305 5926 3814 5972
tri 4214 5926 4260 5972 se
rect 4260 5931 25324 5972
tri 25324 5931 25365 5972 sw
tri 25365 5931 25406 5972 ne
rect 25406 5957 25427 5972
tri 25427 5957 25454 5984 sw
tri 25467 5957 25494 5984 ne
rect 25494 5963 25540 5984
tri 25540 5963 25562 5985 sw
tri 25580 5963 25602 5985 ne
rect 25494 5957 25562 5963
rect 25406 5951 25454 5957
tri 25454 5951 25460 5957 sw
tri 25494 5951 25500 5957 ne
rect 25500 5951 25562 5957
tri 25562 5951 25574 5963 sw
rect 25406 5931 25460 5951
rect 4260 5926 25365 5931
tri 25365 5926 25370 5931 sw
tri 25406 5926 25411 5931 ne
rect 25411 5929 25460 5931
tri 25460 5929 25482 5951 sw
tri 25500 5929 25522 5951 ne
rect 25411 5926 25482 5929
tri 2215 5882 2259 5926 se
rect 2259 5882 3814 5926
tri 4170 5882 4214 5926 se
rect 4214 5923 25370 5926
tri 25370 5923 25373 5926 sw
tri 25411 5923 25414 5926 ne
rect 25414 5923 25482 5926
rect 4214 5917 25373 5923
tri 25373 5917 25379 5923 sw
tri 25414 5917 25420 5923 ne
rect 25420 5917 25482 5923
tri 25482 5917 25494 5929 sw
rect 4214 5895 25379 5917
tri 25379 5895 25401 5917 sw
tri 25420 5895 25442 5917 ne
rect 4214 5882 25401 5895
tri 25401 5882 25414 5895 sw
tri 2196 5863 2215 5882 se
rect 2215 5863 3814 5882
rect 2196 5023 3814 5863
tri 4031 5743 4170 5882 se
rect 4170 5864 25414 5882
rect 4170 5836 4394 5864
tri 4394 5836 4422 5864 nw
tri 23280 5836 23308 5864 ne
rect 23308 5836 25414 5864
rect 4170 5796 4354 5836
tri 4354 5796 4394 5836 nw
tri 4394 5796 4434 5836 se
rect 4434 5796 23125 5836
rect 4170 5783 4341 5796
tri 4341 5783 4354 5796 nw
tri 4381 5783 4394 5796 se
rect 4394 5783 23125 5796
rect 4170 5743 4301 5783
tri 4301 5743 4341 5783 nw
tri 4341 5743 4381 5783 se
rect 4381 5743 23125 5783
tri 23125 5743 23218 5836 sw
tri 23308 5743 23401 5836 ne
rect 23401 5743 25414 5836
tri 3942 5654 4031 5743 se
rect 4031 5729 4287 5743
tri 4287 5729 4301 5743 nw
tri 4327 5729 4341 5743 se
rect 4341 5729 23218 5743
rect 4031 5689 4247 5729
tri 4247 5689 4287 5729 nw
tri 4309 5711 4327 5729 se
rect 4327 5711 23218 5729
tri 23218 5711 23250 5743 sw
tri 4287 5689 4309 5711 se
rect 4309 5689 23250 5711
tri 23401 5689 23455 5743 ne
rect 23455 5689 25414 5743
rect 4031 5654 4212 5689
tri 4212 5654 4247 5689 nw
rect 4287 5688 23250 5689
rect 4287 5660 4448 5688
tri 4448 5660 4476 5688 nw
tri 22997 5660 23025 5688 ne
rect 23025 5660 23250 5688
tri 25063 5660 25092 5689 ne
rect 25092 5660 25414 5689
rect 4287 5654 4442 5660
tri 4442 5654 4448 5660 nw
rect 4711 5654 22985 5660
tri 23025 5654 23031 5660 ne
rect 23031 5654 23250 5660
tri 3887 5599 3942 5654 se
rect 3942 5599 4157 5654
tri 4157 5599 4212 5654 nw
rect 3887 5548 4106 5599
tri 4106 5548 4157 5599 nw
rect 2168 4630 2797 4861
rect 2799 4860 2835 4861
tri 2168 4515 2283 4630 ne
rect 2283 4515 2797 4630
rect 2798 4516 2836 4860
rect 2799 4515 2835 4516
rect 2837 4515 2889 4861
rect 3887 4527 4077 5548
tri 4077 5519 4106 5548 nw
tri 2283 4371 2427 4515 ne
rect 2427 4424 2708 4515
tri 2708 4424 2799 4515 nw
rect 2427 4378 2662 4424
tri 2662 4378 2708 4424 nw
tri 4241 4378 4287 4424 se
rect 4287 4378 4387 5654
tri 4387 5599 4442 5654 nw
rect 4711 5548 4723 5654
rect 22973 5548 22985 5654
tri 23031 5643 23042 5654 ne
rect 4711 5542 22985 5548
tri 4501 5510 4505 5514 se
rect 4505 5510 6617 5514
tri 6617 5510 6621 5514 sw
tri 4467 5476 4501 5510 se
rect 4501 5476 6621 5510
tri 6621 5476 6655 5510 sw
tri 4463 5472 4467 5476 se
rect 4467 5472 6655 5476
tri 6655 5472 6659 5476 sw
rect 2427 4371 2655 4378
tri 2655 4371 2662 4378 nw
tri 4234 4371 4241 4378 se
rect 4241 4371 4387 4378
tri 2427 4366 2432 4371 ne
rect 2432 4366 2655 4371
tri 4229 4366 4234 4371 se
rect 4234 4366 4387 4371
tri 2432 4365 2433 4366 ne
rect 2433 4365 2655 4366
tri 4228 4365 4229 4366 se
rect 4229 4365 4387 4366
rect 2168 4353 2301 4365
rect 2303 4364 2339 4365
rect 2168 4319 2208 4353
rect 2242 4319 2301 4353
rect 2168 4281 2301 4319
rect 2168 4247 2208 4281
rect 2242 4247 2301 4281
rect 2168 4209 2301 4247
rect 2168 4175 2208 4209
rect 2242 4175 2301 4209
rect 2168 4137 2301 4175
rect 2168 4103 2208 4137
rect 2242 4103 2301 4137
rect 2168 4065 2301 4103
rect 2168 4031 2208 4065
rect 2242 4031 2301 4065
rect 2168 4019 2301 4031
rect 2302 4020 2340 4364
rect 2341 4353 2393 4365
rect 2341 4319 2351 4353
rect 2385 4319 2393 4353
tri 2433 4333 2465 4365 ne
rect 2341 4281 2393 4319
rect 2341 4247 2351 4281
rect 2385 4247 2393 4281
rect 2341 4209 2393 4247
rect 2341 4175 2351 4209
rect 2385 4175 2393 4209
rect 2341 4137 2393 4175
rect 2341 4103 2351 4137
rect 2385 4103 2393 4137
rect 2341 4065 2393 4103
rect 2341 4031 2351 4065
rect 2385 4031 2393 4065
rect 2303 4019 2339 4020
rect 2341 4019 2393 4031
rect 2465 4019 2655 4365
tri 2655 4019 2665 4029 sw
rect 4081 4019 4387 4365
tri 4415 5424 4463 5472 se
rect 4463 5424 6659 5472
rect 4415 5421 6659 5424
rect 4415 5414 5858 5421
tri 5858 5414 5865 5421 nw
tri 6446 5414 6453 5421 ne
rect 6453 5414 6659 5421
rect 2168 3942 2276 4019
tri 2276 3994 2301 4019 nw
rect 2465 4007 2665 4019
tri 2665 4007 2677 4019 sw
rect 2465 3982 2677 4007
tri 2677 3982 2702 4007 sw
tri 4390 3982 4415 4007 se
rect 4415 3982 4513 5414
tri 4513 5388 4539 5414 nw
tri 4735 5389 4760 5414 ne
tri 2276 3942 2294 3960 sw
rect 2465 3942 2702 3982
tri 2702 3942 2742 3982 sw
rect 2168 3935 2294 3942
tri 2294 3935 2301 3942 sw
rect 2465 3936 2742 3942
tri 2742 3936 2748 3942 sw
rect 2799 3936 4513 3982
tri 4542 5369 4546 5373 se
rect 4546 5369 4732 5373
rect 2168 3908 2395 3935
tri 2395 3908 2422 3935 sw
rect 2465 3908 2748 3936
tri 2748 3908 2776 3936 sw
rect 2168 3870 2422 3908
tri 2422 3870 2460 3908 sw
rect 2465 3905 4513 3908
tri 2465 3870 2500 3905 ne
rect 2500 3870 4513 3905
rect 2168 3865 2460 3870
tri 2460 3865 2465 3870 sw
tri 2500 3865 2505 3870 ne
rect 2505 3865 4513 3870
rect 2168 3836 2465 3865
tri 2465 3836 2494 3865 sw
tri 2505 3836 2534 3865 ne
rect 2534 3836 4513 3865
rect 2168 3829 2494 3836
tri 2494 3829 2501 3836 sw
tri 2534 3829 2541 3836 ne
rect 2541 3829 4513 3836
rect 2168 3814 2501 3829
tri 2501 3814 2516 3829 sw
tri 2541 3814 2556 3829 ne
rect 2556 3814 4513 3829
rect 2168 3789 2516 3814
tri 2516 3789 2541 3814 sw
tri 2556 3789 2581 3814 ne
rect 2581 3789 4513 3814
rect 2168 3780 2541 3789
tri 2541 3780 2550 3789 sw
tri 2581 3780 2590 3789 ne
rect 2590 3780 4513 3789
rect 2168 3777 2550 3780
tri 2550 3777 2553 3780 sw
tri 2590 3777 2593 3780 ne
rect 2593 3777 4513 3780
rect 2168 3752 2553 3777
tri 2553 3752 2578 3777 sw
tri 4390 3752 4415 3777 ne
rect 2168 3749 2578 3752
tri 2578 3749 2581 3752 sw
rect 2168 3742 4378 3749
tri 4378 3742 4385 3749 sw
rect 2168 3740 4385 3742
tri 4385 3740 4387 3742 sw
rect 2168 3667 4387 3740
tri 4311 3642 4336 3667 ne
rect 968 3624 1060 3626
tri 1060 3624 1062 3626 nw
tri 1934 3624 1936 3626 se
rect 1936 3624 2008 3626
tri 2008 3624 2010 3626 nw
tri 2082 3624 2084 3626 se
rect 2084 3624 2140 3626
rect 968 3620 1056 3624
tri 1056 3620 1060 3624 nw
tri 1930 3620 1934 3624 se
rect 1934 3620 2004 3624
tri 2004 3620 2008 3624 nw
tri 2078 3620 2082 3624 se
rect 2082 3620 2140 3624
tri 968 3605 983 3620 ne
tri 396 3537 416 3557 sw
rect 344 3532 416 3537
tri 416 3532 421 3537 sw
rect 344 3520 955 3532
tri 344 3486 378 3520 ne
rect 378 3486 555 3520
rect 589 3486 627 3520
rect 661 3486 699 3520
rect 733 3486 771 3520
rect 805 3486 843 3520
rect 877 3486 915 3520
rect 949 3486 955 3520
tri 378 3474 390 3486 ne
rect 390 3474 955 3486
tri 982 3420 983 3421 se
rect 983 3420 1041 3620
tri 1041 3605 1056 3620 nw
tri 1915 3605 1930 3620 se
rect 1930 3605 1989 3620
tri 1989 3605 2004 3620 nw
tri 2063 3605 2078 3620 se
rect 2078 3605 2140 3620
tri 1903 3593 1915 3605 se
rect 1915 3593 1977 3605
tri 1977 3593 1989 3605 nw
tri 2051 3593 2063 3605 se
rect 2063 3593 2140 3605
tri 1890 3580 1903 3593 se
rect 1903 3580 1943 3593
tri 1869 3559 1890 3580 se
rect 1890 3559 1943 3580
tri 1943 3559 1977 3593 nw
tri 2017 3559 2051 3593 se
rect 2051 3559 2100 3593
rect 2134 3559 2140 3593
tri 1860 3550 1869 3559 se
rect 1869 3550 1934 3559
tri 1934 3550 1943 3559 nw
tri 2008 3550 2017 3559 se
rect 2017 3550 2140 3559
tri 1847 3537 1860 3550 se
rect 1860 3537 1921 3550
tri 1921 3537 1934 3550 nw
tri 1995 3537 2008 3550 se
rect 2008 3537 2140 3550
tri 1842 3532 1847 3537 se
rect 1847 3532 1916 3537
tri 1916 3532 1921 3537 nw
tri 1990 3532 1995 3537 se
rect 1995 3532 2140 3537
rect 1069 3526 1910 3532
tri 1910 3526 1916 3532 nw
tri 1984 3526 1990 3532 se
rect 1990 3526 2140 3532
rect 1069 3521 1905 3526
tri 1905 3521 1910 3526 nw
tri 1979 3521 1984 3526 se
rect 1984 3521 2140 3526
rect 1069 3520 1890 3521
rect 1069 3486 1075 3520
rect 1109 3486 1147 3520
rect 1181 3486 1219 3520
rect 1253 3486 1291 3520
rect 1325 3486 1363 3520
rect 1397 3486 1435 3520
rect 1469 3506 1890 3520
tri 1890 3506 1905 3521 nw
tri 1964 3506 1979 3521 se
rect 1979 3506 2100 3521
rect 1469 3487 1871 3506
tri 1871 3487 1890 3506 nw
tri 1945 3487 1964 3506 se
rect 1964 3487 2100 3506
rect 2134 3487 2140 3521
rect 1469 3486 1859 3487
rect 1069 3475 1859 3486
tri 1859 3475 1871 3487 nw
tri 1933 3475 1945 3487 se
rect 1945 3475 2140 3487
rect 1069 3474 1858 3475
tri 1858 3474 1859 3475 nw
tri 1932 3474 1933 3475 se
rect 1933 3474 2140 3475
tri 1920 3462 1932 3474 se
rect 1932 3471 2140 3474
rect 1932 3462 2131 3471
tri 2131 3462 2140 3471 nw
rect 2185 3636 4299 3639
tri 4299 3636 4302 3639 sw
rect 2185 3630 4302 3636
tri 4302 3630 4308 3636 sw
rect 2185 3550 4308 3630
rect 2185 3541 4299 3550
tri 4299 3541 4308 3550 nw
rect 2185 3537 2252 3541
tri 2252 3537 2256 3541 nw
tri 4335 3537 4336 3538 se
rect 4336 3537 4387 3667
rect 2185 3526 2241 3537
tri 2241 3526 2252 3537 nw
tri 4324 3526 4335 3537 se
rect 4335 3526 4387 3537
tri 1912 3454 1920 3462 se
rect 1920 3454 2123 3462
tri 2123 3454 2131 3462 nw
tri 1890 3432 1912 3454 se
rect 1912 3447 2116 3454
tri 2116 3447 2123 3454 nw
rect 1912 3432 2101 3447
tri 2101 3432 2116 3447 nw
tri 2170 3432 2185 3447 se
rect 2185 3432 2231 3526
tri 2231 3516 2241 3526 nw
tri 4314 3516 4324 3526 se
rect 4324 3516 4387 3526
tri 4311 3513 4314 3516 se
rect 4314 3513 4387 3516
tri 1879 3421 1890 3432 se
rect 1890 3421 2032 3432
tri 1041 3420 1042 3421 sw
tri 1878 3420 1879 3421 se
rect 1879 3420 2032 3421
tri 2032 3420 2044 3432 nw
tri 2165 3427 2170 3432 se
rect 2170 3427 2231 3432
tri 2158 3420 2165 3427 se
rect 2165 3420 2224 3427
tri 2224 3420 2231 3427 nw
tri 2259 3503 2269 3513 se
rect 2269 3503 4387 3513
tri 958 3396 982 3420 se
rect 982 3396 1042 3420
tri 1042 3396 1066 3420 sw
tri 1854 3396 1878 3420 se
rect 1878 3396 2008 3420
tri 2008 3396 2032 3420 nw
tri 2136 3398 2158 3420 se
rect 2158 3398 2202 3420
tri 2202 3398 2224 3420 nw
rect 2259 3418 4387 3503
tri 2134 3396 2136 3398 se
rect 2136 3396 2200 3398
tri 2200 3396 2202 3398 nw
rect 932 3394 2006 3396
tri 2006 3394 2008 3396 nw
tri 2132 3394 2134 3396 se
rect 2134 3394 2198 3396
tri 2198 3394 2200 3396 nw
rect 457 3382 503 3394
rect 457 3348 463 3382
rect 497 3348 503 3382
rect 361 3320 407 3332
rect 361 3286 367 3320
rect 401 3286 407 3320
rect 361 3247 407 3286
rect 361 3213 367 3247
rect 401 3213 407 3247
rect 361 3174 407 3213
rect 361 3140 367 3174
rect 401 3140 407 3174
rect 361 3101 407 3140
rect 361 3067 367 3101
rect 401 3067 407 3101
rect 361 3028 407 3067
rect 361 2994 367 3028
rect 401 2994 407 3028
rect 361 2955 407 2994
rect 361 2921 367 2955
rect 401 2921 407 2955
rect 361 2882 407 2921
rect 361 2848 367 2882
rect 401 2848 407 2882
rect 361 2809 407 2848
rect 361 2775 367 2809
rect 401 2775 407 2809
rect 361 2736 407 2775
rect 361 2702 367 2736
rect 401 2702 407 2736
rect 361 2663 407 2702
rect 361 2629 367 2663
rect 401 2629 407 2663
rect 361 2590 407 2629
rect 361 2556 367 2590
rect 401 2556 407 2590
rect 361 2517 407 2556
rect 361 2483 367 2517
rect 401 2483 407 2517
rect 361 2444 407 2483
rect 361 2410 367 2444
rect 401 2410 407 2444
rect 361 2371 407 2410
rect 361 2337 367 2371
rect 401 2337 407 2371
rect 361 2298 407 2337
rect 361 2264 367 2298
rect 401 2264 407 2298
rect 361 2225 407 2264
rect 361 2191 367 2225
rect 401 2191 407 2225
rect 361 2152 407 2191
rect 361 2118 367 2152
rect 401 2118 407 2152
rect 361 2079 407 2118
rect 361 2045 367 2079
rect 401 2045 407 2079
rect 361 2006 407 2045
rect 361 1972 367 2006
rect 401 1972 407 2006
rect 361 1933 407 1972
rect 361 1899 367 1933
rect 401 1899 407 1933
rect 361 1860 407 1899
rect 361 1826 367 1860
rect 401 1826 407 1860
rect 361 1787 407 1826
rect 361 1753 367 1787
rect 401 1753 407 1787
rect 361 1714 407 1753
rect 361 1680 367 1714
rect 401 1680 407 1714
rect 361 1641 407 1680
rect 361 1607 367 1641
rect 401 1607 407 1641
rect 361 1567 407 1607
rect 361 1533 367 1567
rect 401 1533 407 1567
rect 361 1493 407 1533
rect 361 1459 367 1493
rect 401 1459 407 1493
rect 361 1419 407 1459
rect 361 1385 367 1419
rect 401 1385 407 1419
rect 361 1345 407 1385
rect 361 1311 367 1345
rect 401 1311 407 1345
rect 361 1271 407 1311
rect 361 1237 367 1271
rect 401 1237 407 1271
rect 361 1197 407 1237
rect 361 1163 367 1197
rect 401 1163 407 1197
rect 361 1123 407 1163
rect 361 1089 367 1123
rect 401 1089 407 1123
rect 361 1049 407 1089
rect 361 1015 367 1049
rect 401 1015 407 1049
rect 361 975 407 1015
rect 361 941 367 975
rect 401 941 407 975
rect 361 901 407 941
rect 361 867 367 901
rect 401 867 407 901
rect 361 827 407 867
rect 361 793 367 827
rect 401 793 407 827
rect 361 753 407 793
rect 361 719 367 753
rect 401 719 407 753
rect 361 679 407 719
rect 361 645 367 679
rect 401 645 407 679
rect 361 605 407 645
rect 361 571 367 605
rect 401 571 407 605
rect 361 531 407 571
rect 361 497 367 531
rect 401 497 407 531
rect 361 457 407 497
rect 361 423 367 457
rect 401 423 407 457
rect 361 383 407 423
rect 457 3310 503 3348
rect 932 3387 1999 3394
tri 1999 3387 2006 3394 nw
tri 2125 3387 2132 3394 se
rect 2132 3387 2191 3394
tri 2191 3387 2198 3394 nw
tri 4410 3387 4415 3392 se
rect 4415 3387 4513 3777
rect 932 3382 1994 3387
tri 1994 3382 1999 3387 nw
tri 2120 3382 2125 3387 se
rect 2125 3382 2186 3387
tri 2186 3382 2191 3387 nw
tri 4405 3382 4410 3387 se
rect 4410 3382 4513 3387
rect 932 3348 1960 3382
tri 1960 3348 1994 3382 nw
tri 2086 3348 2120 3382 se
rect 2120 3348 2152 3382
tri 2152 3348 2186 3382 nw
tri 4390 3367 4405 3382 se
rect 4405 3367 4513 3382
rect 932 3338 1950 3348
tri 1950 3338 1960 3348 nw
tri 2076 3338 2086 3348 se
rect 2086 3338 2142 3348
tri 2142 3338 2152 3348 nw
tri 2070 3332 2076 3338 se
rect 2076 3332 2136 3338
tri 2136 3332 2142 3338 nw
tri 2054 3316 2070 3332 se
rect 2070 3316 2120 3332
tri 2120 3316 2136 3332 nw
tri 2050 3312 2054 3316 se
rect 2054 3312 2116 3316
tri 2116 3312 2120 3316 nw
tri 2048 3310 2050 3312 se
rect 2050 3310 2114 3312
tri 2114 3310 2116 3312 nw
rect 457 3276 463 3310
rect 497 3276 503 3310
rect 457 3238 503 3276
rect 457 3204 463 3238
rect 497 3204 503 3238
rect 457 3166 503 3204
rect 457 3132 463 3166
rect 497 3132 503 3166
rect 457 3094 503 3132
rect 457 3060 463 3094
rect 497 3060 503 3094
rect 457 523 503 3060
rect 457 489 463 523
rect 497 489 503 523
rect 457 451 503 489
rect 569 3276 2080 3310
tri 2080 3276 2114 3310 nw
rect 569 3266 2070 3276
tri 2070 3266 2080 3276 nw
rect 2246 3270 4513 3367
tri 4390 3266 4394 3270 ne
rect 4394 3266 4513 3270
rect 569 3243 716 3266
tri 716 3243 739 3266 nw
tri 4394 3245 4415 3266 ne
rect 569 3132 714 3243
tri 714 3241 716 3243 nw
tri 2142 3241 2143 3242 se
rect 2143 3241 4366 3242
tri 2141 3240 2142 3241 se
rect 2142 3240 4366 3241
tri 2139 3238 2141 3240 se
rect 2141 3238 4366 3240
tri 742 3229 751 3238 se
rect 751 3229 4366 3238
rect 742 3226 4366 3229
rect 742 3192 757 3226
rect 791 3192 829 3226
rect 863 3192 901 3226
rect 935 3192 973 3226
rect 1007 3192 1045 3226
rect 1079 3192 1117 3226
rect 1151 3192 4366 3226
rect 742 3182 4366 3192
rect 742 3152 1243 3182
tri 888 3148 892 3152 ne
rect 892 3148 1243 3152
rect 1277 3148 4366 3182
tri 892 3135 905 3148 ne
rect 905 3135 4366 3148
tri 714 3132 717 3135 sw
tri 905 3132 908 3135 ne
rect 908 3132 4366 3135
rect 569 3130 717 3132
tri 717 3130 719 3132 sw
tri 908 3130 910 3132 ne
rect 910 3130 4366 3132
rect 569 3110 719 3130
tri 719 3110 739 3130 sw
tri 910 3110 930 3130 ne
rect 930 3117 4366 3130
rect 930 3114 2209 3117
tri 2209 3114 2212 3117 nw
rect 930 3110 2192 3114
rect 569 3098 860 3110
rect 569 3064 604 3098
rect 638 3064 676 3098
rect 710 3064 748 3098
rect 782 3064 820 3098
rect 854 3064 860 3098
tri 930 3076 964 3110 ne
rect 964 3076 1243 3110
rect 1277 3097 2192 3110
tri 2192 3097 2209 3114 nw
tri 4398 3097 4415 3114 se
rect 4415 3097 4513 3266
rect 1277 3096 2191 3097
tri 2191 3096 2192 3097 nw
tri 4397 3096 4398 3097 se
rect 4398 3096 4513 3097
rect 1277 3093 2188 3096
tri 2188 3093 2191 3096 nw
tri 4394 3093 4397 3096 se
rect 4397 3093 4513 3096
rect 1277 3089 2184 3093
tri 2184 3089 2188 3093 nw
tri 4390 3089 4394 3093 se
rect 4394 3089 4513 3093
rect 1277 3076 2154 3089
rect 569 2786 860 3064
tri 964 3059 981 3076 ne
rect 981 3059 2154 3076
tri 2154 3059 2184 3089 nw
tri 981 3056 984 3059 ne
rect 984 3056 2151 3059
tri 2151 3056 2154 3059 nw
tri 984 3038 1002 3056 ne
rect 1002 3038 2119 3056
tri 1002 3004 1036 3038 ne
rect 1036 3004 1243 3038
rect 1277 3024 2119 3038
tri 2119 3024 2151 3056 nw
rect 1277 3020 2115 3024
tri 2115 3020 2119 3024 nw
rect 1277 3004 2093 3020
tri 1036 2998 1042 3004 ne
rect 1042 2998 2093 3004
tri 2093 2998 2115 3020 nw
rect 2246 2997 4513 3089
tri 4538 2982 4542 2986 se
rect 4542 2982 4732 5369
tri 4510 2954 4538 2982 se
rect 4538 2954 4732 2982
rect 569 2752 604 2786
rect 638 2752 676 2786
rect 710 2752 748 2786
rect 782 2752 820 2786
rect 854 2752 860 2786
rect 569 2474 860 2752
rect 569 2440 604 2474
rect 638 2440 676 2474
rect 710 2440 748 2474
rect 782 2440 820 2474
rect 854 2440 860 2474
rect 569 2162 860 2440
rect 888 2953 2060 2954
tri 2060 2953 2061 2954 sw
tri 4509 2953 4510 2954 se
rect 4510 2953 4732 2954
rect 888 2951 2061 2953
tri 2061 2951 2063 2953 sw
rect 888 2947 2063 2951
tri 2063 2947 2067 2951 sw
rect 888 2942 2067 2947
rect 888 2908 981 2942
rect 1015 2908 1053 2942
rect 1087 2908 1125 2942
rect 1159 2913 2067 2942
tri 2067 2913 2101 2947 sw
rect 1159 2908 2101 2913
tri 2101 2908 2106 2913 sw
rect 888 2896 2106 2908
tri 2106 2896 2118 2908 sw
rect 888 2878 2118 2896
tri 2118 2878 2136 2896 sw
rect 888 2874 2136 2878
tri 2136 2874 2140 2878 sw
rect 888 2854 2140 2874
tri 2140 2854 2160 2874 sw
rect 2249 2854 4732 2953
rect 888 2840 2160 2854
tri 2160 2840 2174 2854 sw
tri 4445 2840 4459 2854 ne
rect 4459 2840 4732 2854
rect 888 2834 2174 2840
tri 2174 2834 2180 2840 sw
tri 4459 2834 4465 2840 ne
rect 4465 2834 4732 2840
rect 888 2829 2180 2834
tri 2180 2829 2185 2834 sw
tri 4465 2829 4470 2834 ne
rect 888 2826 2185 2829
tri 2185 2826 2188 2829 sw
rect 888 2817 4433 2826
tri 4433 2817 4442 2826 sw
rect 888 2696 4442 2817
rect 888 2694 4440 2696
tri 4440 2694 4442 2696 nw
rect 888 2687 4433 2694
tri 4433 2687 4440 2694 nw
rect 888 2686 2195 2687
tri 2195 2686 2196 2687 nw
rect 888 2684 2193 2686
tri 2193 2684 2195 2686 nw
rect 888 2672 2168 2684
tri 1104 2671 1105 2672 ne
rect 1105 2671 2168 2672
rect 888 2670 1103 2671
tri 1103 2670 1104 2671 sw
tri 1105 2670 1106 2671 ne
rect 1106 2670 2168 2671
rect 888 2668 1104 2670
tri 1104 2668 1106 2670 sw
tri 1106 2668 1108 2670 ne
rect 1108 2668 2168 2670
rect 888 2666 1106 2668
tri 1106 2666 1108 2668 sw
tri 1108 2666 1110 2668 ne
rect 1110 2666 2168 2668
rect 888 2664 1108 2666
tri 1108 2664 1110 2666 sw
tri 1110 2664 1112 2666 ne
rect 1112 2664 2168 2666
rect 888 2662 1110 2664
tri 1110 2662 1112 2664 sw
tri 1112 2662 1114 2664 ne
rect 1114 2662 2168 2664
rect 888 2660 1112 2662
tri 1112 2660 1114 2662 sw
tri 1114 2660 1116 2662 ne
rect 1116 2660 2168 2662
rect 888 2659 1114 2660
tri 1114 2659 1115 2660 sw
tri 1116 2659 1117 2660 ne
rect 1117 2659 2168 2660
tri 2168 2659 2193 2684 nw
tri 4445 2659 4470 2684 se
rect 4470 2659 4732 2834
rect 888 2658 1115 2659
tri 1115 2658 1116 2659 sw
tri 1117 2658 1118 2659 ne
rect 888 2643 1116 2658
rect 888 2630 1078 2642
rect 1080 2641 1116 2643
rect 1118 2655 2164 2659
tri 2164 2655 2168 2659 nw
rect 1118 2642 2151 2655
tri 2151 2642 2164 2655 nw
rect 888 2596 894 2630
rect 928 2596 966 2630
rect 1000 2596 1038 2630
rect 1072 2596 1078 2630
rect 888 2584 1078 2596
rect 1079 2585 1117 2641
rect 1118 2621 2130 2642
tri 2130 2621 2151 2642 nw
rect 2249 2637 4732 2659
rect 2249 2625 4720 2637
tri 4720 2625 4732 2637 nw
rect 4760 5171 5840 5414
tri 5840 5396 5858 5414 nw
tri 6453 5396 6471 5414 ne
rect 6471 5396 6659 5414
tri 6471 5394 6473 5396 ne
rect 4760 5069 4864 5171
tri 4864 5069 4966 5171 nw
tri 5560 5069 5662 5171 ne
rect 5662 5069 5840 5171
rect 4760 5065 4860 5069
tri 4860 5065 4864 5069 nw
tri 5022 5067 5024 5069 se
rect 5024 5067 5488 5069
tri 5488 5067 5490 5069 sw
tri 5662 5067 5664 5069 ne
rect 5664 5067 5840 5069
tri 5020 5065 5022 5067 se
rect 5022 5065 5490 5067
rect 4760 3942 4832 5065
tri 4832 5037 4860 5065 nw
tri 4992 5037 5020 5065 se
rect 5020 5060 5490 5065
tri 5490 5060 5497 5067 sw
tri 5664 5060 5671 5067 ne
rect 5020 5037 5497 5060
tri 5497 5037 5520 5060 sw
tri 4896 4941 4992 5037 se
rect 4992 4941 5520 5037
rect 4760 3908 4780 3942
rect 4814 3908 4832 3942
rect 4760 3870 4832 3908
rect 4760 3836 4780 3870
rect 4814 3836 4832 3870
rect 2249 2621 4716 2625
tri 4716 2621 4720 2625 nw
tri 4756 2621 4760 2625 se
rect 4760 2621 4832 3836
rect 1118 2612 2121 2621
tri 2121 2612 2130 2621 nw
rect 2249 2612 4707 2621
tri 4707 2612 4716 2621 nw
tri 4747 2612 4756 2621 se
rect 4756 2612 4832 2621
rect 1118 2586 2095 2612
tri 2095 2586 2121 2612 nw
rect 2249 2597 4692 2612
tri 4692 2597 4707 2612 nw
tri 4732 2597 4747 2612 se
rect 4747 2597 4832 2612
rect 2249 2586 4681 2597
tri 4681 2586 4692 2597 nw
tri 4721 2586 4732 2597 se
rect 4732 2586 4832 2597
rect 1080 2583 1116 2585
rect 888 2568 1116 2583
rect 1118 2584 2093 2586
tri 2093 2584 2095 2586 nw
rect 2249 2584 4679 2586
tri 4679 2584 4681 2586 nw
tri 4719 2584 4721 2586 se
rect 4721 2584 4832 2586
rect 1118 2582 2091 2584
tri 2091 2582 2093 2584 nw
rect 2249 2582 4677 2584
tri 4677 2582 4679 2584 nw
tri 4717 2582 4719 2584 se
rect 4719 2582 4832 2584
rect 888 2566 1114 2568
tri 1114 2566 1116 2568 nw
tri 1116 2566 1118 2568 se
rect 1118 2566 2074 2582
rect 888 2565 1113 2566
tri 1113 2565 1114 2566 nw
tri 1115 2565 1116 2566 se
rect 1116 2565 2074 2566
tri 2074 2565 2091 2582 nw
rect 2249 2565 4660 2582
tri 4660 2565 4677 2582 nw
tri 4700 2565 4717 2582 se
rect 4717 2565 4832 2582
rect 888 2564 1112 2565
tri 1112 2564 1113 2565 nw
tri 1114 2564 1115 2565 se
rect 1115 2564 1335 2565
rect 888 2562 1110 2564
tri 1110 2562 1112 2564 nw
tri 1112 2562 1114 2564 se
rect 1114 2562 1335 2564
rect 888 2560 1108 2562
tri 1108 2560 1110 2562 nw
tri 1110 2560 1112 2562 se
rect 1112 2560 1335 2562
rect 888 2558 1106 2560
tri 1106 2558 1108 2560 nw
tri 1108 2558 1110 2560 se
rect 1110 2558 1335 2560
rect 888 2556 1104 2558
tri 1104 2556 1106 2558 nw
tri 1106 2556 1108 2558 se
rect 1108 2556 1335 2558
rect 888 2555 1103 2556
tri 1103 2555 1104 2556 nw
tri 1105 2555 1106 2556 se
rect 1106 2555 1335 2556
tri 1104 2554 1105 2555 se
rect 1105 2554 1335 2555
rect 888 2548 1335 2554
tri 1335 2548 1352 2565 nw
tri 4683 2548 4700 2565 se
rect 4700 2548 4832 2565
rect 888 2538 1325 2548
tri 1325 2538 1335 2548 nw
tri 4673 2538 4683 2548 se
rect 4683 2538 4832 2548
rect 888 2513 1300 2538
tri 1300 2513 1325 2538 nw
tri 4648 2513 4673 2538 se
rect 4673 2531 4832 2538
rect 4673 2513 4814 2531
tri 4814 2513 4832 2531 nw
tri 4860 4905 4896 4941 se
rect 4896 4914 5051 4941
tri 5051 4914 5078 4941 nw
tri 5438 4914 5465 4941 ne
rect 5465 4914 5520 4941
tri 5520 4914 5643 5037 sw
rect 4896 4905 5026 4914
rect 4860 3620 5026 4905
tri 5026 4889 5051 4914 nw
tri 5465 4889 5490 4914 ne
rect 4860 3586 4893 3620
rect 4927 3586 4965 3620
rect 4999 3586 5026 3620
rect 888 2509 1296 2513
tri 1296 2509 1300 2513 nw
tri 4644 2509 4648 2513 se
rect 4648 2509 4810 2513
tri 4810 2509 4814 2513 nw
rect 888 2498 1285 2509
tri 1285 2498 1296 2509 nw
tri 1388 2498 1399 2509 se
rect 1399 2498 4799 2509
tri 4799 2498 4810 2509 nw
rect 888 2492 1279 2498
tri 1279 2492 1285 2498 nw
tri 1382 2492 1388 2498 se
rect 1388 2492 4776 2498
rect 888 2486 1273 2492
tri 1273 2486 1279 2492 nw
tri 1376 2486 1382 2492 se
rect 1382 2486 1906 2492
rect 888 2470 1257 2486
tri 1257 2470 1273 2486 nw
tri 1360 2470 1376 2486 se
rect 1376 2470 1906 2486
rect 888 2462 1249 2470
tri 1249 2462 1257 2470 nw
tri 1352 2462 1360 2470 se
rect 1360 2462 1906 2470
rect 888 2458 1245 2462
tri 1245 2458 1249 2462 nw
tri 1350 2460 1352 2462 se
rect 1352 2460 1906 2462
rect 1350 2458 1906 2460
rect 1940 2458 2045 2492
rect 2079 2458 2118 2492
rect 2152 2458 2191 2492
rect 2225 2458 2264 2492
rect 2298 2458 2337 2492
rect 2371 2458 2410 2492
rect 2444 2458 2483 2492
rect 2517 2458 2556 2492
rect 2590 2458 2629 2492
rect 2663 2458 2702 2492
rect 2736 2458 2775 2492
rect 2809 2458 2848 2492
rect 2882 2458 2921 2492
rect 2955 2458 2994 2492
rect 3028 2458 3067 2492
rect 3101 2458 3140 2492
rect 3174 2458 3213 2492
rect 3247 2458 3286 2492
rect 3320 2458 3359 2492
rect 3393 2458 3432 2492
rect 3466 2458 3505 2492
rect 3539 2458 3578 2492
rect 3612 2458 3651 2492
rect 3685 2458 3723 2492
rect 3757 2458 3795 2492
rect 3829 2458 3867 2492
rect 3901 2458 3939 2492
rect 3973 2458 4011 2492
rect 4045 2458 4083 2492
rect 4117 2458 4155 2492
rect 4189 2458 4227 2492
rect 4261 2458 4299 2492
rect 4333 2458 4371 2492
rect 4405 2458 4443 2492
rect 4477 2458 4515 2492
rect 4549 2458 4587 2492
rect 4621 2458 4659 2492
rect 4693 2475 4776 2492
tri 4776 2475 4799 2498 nw
tri 4856 2475 4860 2479 se
rect 4860 2475 5026 3586
rect 4693 2464 4765 2475
tri 4765 2464 4776 2475 nw
tri 4845 2464 4856 2475 se
rect 4856 2464 5026 2475
rect 4693 2458 4750 2464
rect 888 2440 1227 2458
tri 1227 2440 1245 2458 nw
rect 1350 2449 4750 2458
tri 4750 2449 4765 2464 nw
tri 4830 2449 4845 2464 se
rect 4845 2449 5026 2464
rect 1350 2440 2229 2449
tri 2229 2440 2238 2449 nw
tri 4821 2440 4830 2449 se
rect 4830 2440 5026 2449
rect 888 2436 1223 2440
tri 1223 2436 1227 2440 nw
rect 1350 2436 2225 2440
tri 2225 2436 2229 2440 nw
tri 4817 2436 4821 2440 se
rect 4821 2436 5026 2440
rect 888 2420 1207 2436
tri 1207 2420 1223 2436 nw
rect 1350 2421 2210 2436
tri 2210 2421 2225 2436 nw
tri 4802 2421 4817 2436 se
rect 4817 2421 5026 2436
rect 1350 2420 2191 2421
rect 888 2418 1205 2420
tri 1205 2418 1207 2420 nw
rect 1203 2417 1204 2418
tri 1204 2417 1205 2418 nw
rect 889 2416 1202 2417
tri 1203 2416 1204 2417 nw
rect 1350 2386 1906 2420
rect 1940 2402 2191 2420
tri 2191 2402 2210 2421 nw
tri 2271 2402 2290 2421 se
rect 2290 2402 5026 2421
rect 1940 2390 2179 2402
tri 2179 2390 2191 2402 nw
tri 2259 2390 2271 2402 se
rect 2271 2390 5026 2402
rect 1940 2386 2169 2390
rect 1350 2380 2169 2386
tri 2169 2380 2179 2390 nw
tri 2249 2380 2259 2390 se
rect 2259 2380 5026 2390
rect 569 2128 604 2162
rect 638 2128 676 2162
rect 710 2128 748 2162
rect 782 2128 820 2162
rect 854 2128 860 2162
rect 569 2018 860 2128
rect 889 2379 1202 2380
rect 888 2318 1203 2378
rect 888 2284 981 2318
rect 1015 2284 1053 2318
rect 1087 2284 1125 2318
rect 1159 2284 1203 2318
rect 888 2047 1203 2284
rect 1350 2376 2165 2380
tri 2165 2376 2169 2380 nw
tri 2245 2376 2249 2380 se
rect 2249 2376 5026 2380
rect 1350 2367 2156 2376
tri 2156 2367 2165 2376 nw
tri 2236 2367 2245 2376 se
rect 2245 2367 5026 2376
rect 1350 2364 2153 2367
tri 2153 2364 2156 2367 nw
tri 2233 2364 2236 2367 se
rect 2236 2364 5026 2367
rect 1350 2331 2120 2364
tri 2120 2331 2153 2364 nw
tri 2200 2331 2233 2364 se
rect 2233 2331 5026 2364
rect 1350 2330 2119 2331
tri 2119 2330 2120 2331 nw
tri 2199 2330 2200 2331 se
rect 2200 2330 5026 2331
rect 1350 2329 2118 2330
tri 2118 2329 2119 2330 nw
tri 2198 2329 2199 2330 se
rect 2199 2329 5026 2330
rect 1350 2326 2115 2329
tri 2115 2326 2118 2329 nw
tri 2195 2326 2198 2329 se
rect 2198 2326 5026 2329
rect 1350 2318 2107 2326
tri 2107 2318 2115 2326 nw
tri 2187 2318 2195 2326 se
rect 2195 2318 5026 2326
rect 1350 2316 2105 2318
tri 2105 2316 2107 2318 nw
tri 2185 2316 2187 2318 se
rect 2187 2316 5026 2318
rect 1350 2294 2083 2316
tri 2083 2294 2105 2316 nw
tri 2163 2294 2185 2316 se
rect 2185 2294 5026 2316
rect 1350 2290 2079 2294
tri 2079 2290 2083 2294 nw
tri 2159 2290 2163 2294 se
rect 2163 2290 5026 2294
tri 888 2045 890 2047 ne
rect 890 2045 1203 2047
tri 890 2031 904 2045 ne
rect 904 2031 1203 2045
tri 860 2018 873 2031 sw
tri 904 2018 917 2031 ne
rect 917 2018 1203 2031
rect 569 2011 873 2018
tri 873 2011 880 2018 sw
tri 917 2011 924 2018 ne
rect 924 2011 1203 2018
rect 569 2006 880 2011
tri 880 2006 885 2011 sw
tri 924 2006 929 2011 ne
rect 929 2006 1203 2011
rect 569 2003 885 2006
tri 885 2003 888 2006 sw
tri 929 2003 932 2006 ne
rect 932 2003 981 2006
rect 569 1972 888 2003
tri 888 1972 919 2003 sw
tri 932 1972 963 2003 ne
rect 963 1972 981 2003
rect 1015 1972 1053 2006
rect 1087 1972 1125 2006
rect 1159 1972 1203 2006
rect 569 1960 919 1972
tri 919 1960 931 1972 sw
tri 963 1960 975 1972 ne
rect 975 1960 1203 1972
rect 1231 2261 1289 2267
rect 1231 2227 1243 2261
rect 1277 2227 1289 2261
rect 1231 2189 1289 2227
rect 1231 2155 1243 2189
rect 1277 2155 1289 2189
rect 1231 2117 1289 2155
rect 1231 2083 1243 2117
rect 1277 2083 1289 2117
rect 1231 2045 1289 2083
rect 1231 2011 1243 2045
rect 1277 2011 1289 2045
rect 1231 1973 1289 2011
rect 569 1939 931 1960
tri 931 1939 952 1960 sw
rect 1231 1939 1243 1973
rect 1277 1939 1289 1973
rect 569 1929 952 1939
tri 952 1929 962 1939 sw
rect 569 1925 962 1929
tri 962 1925 966 1929 sw
rect 569 1901 966 1925
tri 966 1901 990 1925 sw
rect 1231 1901 1289 1939
rect 569 1886 990 1901
tri 990 1886 1005 1901 sw
rect 569 1867 1159 1886
tri 1159 1867 1178 1886 sw
rect 1231 1867 1243 1901
rect 1277 1867 1289 1901
rect 569 1861 1178 1867
tri 1178 1861 1184 1867 sw
rect 1231 1861 1289 1867
rect 569 1856 1184 1861
tri 1184 1856 1189 1861 sw
rect 569 1852 1189 1856
tri 1189 1852 1193 1856 sw
rect 569 1838 1193 1852
tri 1193 1838 1207 1852 sw
rect 1350 1838 2064 2290
tri 2064 2275 2079 2290 nw
tri 2144 2275 2159 2290 se
rect 2159 2275 5026 2290
tri 2126 2257 2144 2275 se
rect 2144 2257 5026 2275
tri 2125 2256 2126 2257 se
rect 2126 2256 5025 2257
tri 5025 2256 5026 2257 nw
rect 5054 4515 5296 4877
rect 5298 4876 5334 4877
rect 5297 4516 5335 4876
rect 5298 4515 5334 4516
rect 5336 4515 5462 4877
tri 2120 2251 2125 2256 se
rect 2125 2251 5017 2256
rect 2120 2248 5017 2251
tri 5017 2248 5025 2256 nw
rect 2120 2242 2231 2248
tri 2231 2242 2237 2248 nw
tri 5051 2242 5054 2245 se
rect 5054 2242 5244 4515
tri 5244 4463 5296 4515 nw
rect 2120 2148 2212 2242
tri 2212 2223 2231 2242 nw
tri 5032 2223 5051 2242 se
rect 5051 2223 5244 2242
tri 5030 2221 5032 2223 se
rect 5032 2221 5244 2223
tri 5029 2220 5030 2221 se
rect 5030 2220 5244 2221
rect 2249 2162 5244 2220
tri 5029 2159 5032 2162 ne
rect 5032 2159 5244 2162
tri 2212 2148 2223 2159 sw
tri 5032 2148 5043 2159 ne
rect 5043 2148 5244 2159
rect 2120 2144 2223 2148
tri 2223 2144 2227 2148 sw
tri 5043 2144 5047 2148 ne
rect 5047 2144 5244 2148
rect 2120 2134 2227 2144
tri 2227 2134 2237 2144 sw
tri 5047 2137 5054 2144 ne
rect 2120 1936 4989 2134
rect 2120 1929 2230 1936
tri 2230 1929 2237 1936 nw
tri 5050 1929 5054 1933 se
rect 5054 1929 5244 2144
rect 2120 1925 2226 1929
tri 2226 1925 2230 1929 nw
tri 5046 1925 5050 1929 se
rect 5050 1925 5244 1929
rect 569 1819 1207 1838
tri 1207 1819 1226 1838 sw
rect 569 1818 1226 1819
tri 1226 1818 1227 1819 sw
rect 2120 1818 2212 1925
tri 2212 1911 2226 1925 nw
tri 5032 1911 5046 1925 se
rect 5046 1911 5244 1925
tri 5029 1908 5032 1911 se
rect 5032 1908 5244 1911
rect 2249 1850 5244 1908
tri 5029 1825 5054 1850 ne
tri 2212 1818 2213 1819 sw
rect 569 1814 1227 1818
tri 1227 1814 1231 1818 sw
rect 569 1798 1231 1814
tri 1231 1798 1247 1814 sw
tri 2104 1798 2120 1814 se
rect 2120 1798 2213 1818
tri 2213 1798 2233 1818 sw
rect 569 1794 1247 1798
tri 1247 1794 1251 1798 sw
tri 2100 1794 2104 1798 se
rect 2104 1794 2233 1798
tri 2233 1794 2237 1798 sw
rect 569 1783 1251 1794
tri 1251 1783 1262 1794 sw
tri 2089 1783 2100 1794 se
rect 2100 1783 4989 1794
rect 569 1782 1262 1783
tri 1262 1782 1263 1783 sw
tri 2088 1782 2089 1783 se
rect 2089 1782 4989 1783
rect 569 1654 4989 1782
rect 569 1650 1003 1654
tri 1003 1650 1007 1654 nw
tri 1462 1650 1466 1654 ne
rect 1466 1650 4989 1654
rect 569 1637 990 1650
tri 990 1637 1003 1650 nw
tri 1466 1637 1479 1650 ne
rect 1479 1637 4989 1650
rect 569 1633 986 1637
tri 986 1633 990 1637 nw
tri 1479 1633 1483 1637 ne
rect 1483 1633 4989 1637
rect 569 1599 952 1633
tri 952 1599 986 1633 nw
tri 1483 1620 1496 1633 ne
rect 1496 1624 4989 1633
rect 1496 1620 2205 1624
tri 2205 1620 2209 1624 nw
tri 5053 1620 5054 1621 se
rect 5054 1620 5244 1850
rect 569 1596 949 1599
tri 949 1596 952 1599 nw
rect 569 1584 937 1596
tri 937 1584 949 1596 nw
tri 977 1584 989 1596 se
rect 989 1584 1440 1596
rect 569 1556 909 1584
tri 909 1556 937 1584 nw
tri 949 1556 977 1584 se
rect 977 1556 1040 1584
rect 569 1550 903 1556
tri 903 1550 909 1556 nw
tri 943 1550 949 1556 se
rect 949 1550 1040 1556
rect 1074 1550 1112 1584
rect 1146 1550 1184 1584
rect 1218 1550 1256 1584
rect 1290 1550 1328 1584
rect 1362 1550 1400 1584
rect 1434 1550 1440 1584
rect 569 1538 891 1550
tri 891 1538 903 1550 nw
tri 931 1538 943 1550 se
rect 943 1538 1440 1550
rect 569 1537 890 1538
tri 890 1537 891 1538 nw
tri 930 1537 931 1538 se
rect 931 1537 1440 1538
rect 569 1526 879 1537
tri 879 1526 890 1537 nw
tri 919 1526 930 1537 se
rect 930 1526 1440 1537
rect 569 1428 862 1526
tri 862 1509 879 1526 nw
tri 902 1509 919 1526 se
rect 919 1509 1440 1526
tri 899 1506 902 1509 se
rect 902 1506 1440 1509
rect 1496 1509 2184 1620
tri 2184 1599 2205 1620 nw
tri 5032 1599 5053 1620 se
rect 5053 1599 5244 1620
tri 5029 1596 5032 1599 se
rect 5032 1596 5244 1599
rect 2242 1538 5244 1596
tri 5029 1526 5041 1538 ne
rect 5041 1526 5244 1538
tri 5041 1514 5053 1526 ne
rect 5053 1514 5244 1526
tri 2184 1509 2189 1514 sw
tri 5053 1513 5054 1514 ne
tri 895 1502 899 1506 se
rect 899 1502 1222 1506
tri 1222 1502 1226 1506 nw
rect 1496 1502 2189 1509
tri 2189 1502 2196 1509 sw
rect 569 1394 604 1428
rect 638 1394 676 1428
rect 710 1394 748 1428
rect 782 1394 820 1428
rect 854 1394 862 1428
rect 569 1116 862 1394
rect 569 1082 604 1116
rect 638 1082 676 1116
rect 710 1082 748 1116
rect 782 1082 820 1116
rect 854 1082 862 1116
rect 569 869 862 1082
tri 890 1497 895 1502 se
rect 895 1497 1211 1502
rect 890 1491 1211 1497
tri 1211 1491 1222 1502 nw
rect 1496 1491 2196 1502
tri 2196 1491 2207 1502 sw
rect 890 1487 1207 1491
tri 1207 1487 1211 1491 nw
rect 1496 1487 2207 1491
tri 2207 1487 2211 1491 sw
rect 890 1482 1202 1487
tri 1202 1482 1207 1487 nw
rect 1496 1482 2211 1487
tri 2211 1482 2216 1487 sw
rect 890 1338 1201 1482
tri 1201 1481 1202 1482 nw
tri 1495 1481 1496 1482 se
rect 1496 1481 4989 1482
tri 1471 1457 1495 1481 se
rect 1495 1457 4989 1481
tri 1242 1453 1246 1457 se
rect 1246 1453 4989 1457
tri 1229 1440 1242 1453 se
rect 1242 1440 4989 1453
rect 1229 1428 4989 1440
rect 1229 1394 1235 1428
rect 1269 1394 1307 1428
rect 1341 1394 1379 1428
rect 1413 1394 1451 1428
rect 1485 1394 4989 1428
rect 1229 1380 4989 1394
tri 1229 1363 1246 1380 ne
rect 1246 1363 4989 1380
tri 1471 1354 1480 1363 ne
rect 1480 1354 4989 1363
tri 1480 1345 1489 1354 ne
rect 1489 1345 4989 1354
tri 1489 1341 1493 1345 ne
rect 1493 1341 4989 1345
tri 1201 1338 1204 1341 sw
tri 1493 1338 1496 1341 ne
rect 1496 1340 4989 1341
rect 1496 1338 2214 1340
tri 2214 1338 2216 1340 nw
rect 890 1316 1204 1338
tri 1204 1316 1226 1338 sw
rect 890 1194 1440 1316
rect 1496 1206 2184 1338
tri 2184 1308 2214 1338 nw
tri 5053 1308 5054 1309 se
rect 5054 1308 5244 1514
tri 5052 1307 5053 1308 se
rect 5053 1307 5244 1308
tri 5029 1284 5052 1307 se
rect 5052 1284 5244 1307
rect 2242 1226 5244 1284
rect 5272 4366 5370 4378
rect 5372 4377 5408 4378
rect 5272 4332 5278 4366
rect 5312 4332 5370 4366
rect 5272 4294 5370 4332
rect 5272 4260 5278 4294
rect 5312 4260 5370 4294
rect 5272 4222 5370 4260
rect 5272 4188 5278 4222
rect 5312 4188 5370 4222
rect 5272 4150 5370 4188
rect 5272 4116 5278 4150
rect 5312 4116 5370 4150
rect 5272 4078 5370 4116
rect 5272 4044 5278 4078
rect 5312 4044 5370 4078
rect 5272 4016 5370 4044
rect 5371 4017 5409 4377
rect 5410 4366 5462 4378
rect 5410 4332 5416 4366
rect 5450 4332 5462 4366
rect 5410 4294 5462 4332
rect 5410 4260 5416 4294
rect 5450 4260 5462 4294
rect 5410 4222 5462 4260
rect 5410 4188 5416 4222
rect 5450 4188 5462 4222
rect 5410 4150 5462 4188
rect 5410 4116 5416 4150
rect 5450 4116 5462 4150
rect 5410 4078 5462 4116
rect 5410 4044 5416 4078
rect 5450 4044 5462 4078
rect 5372 4016 5408 4017
rect 5410 4016 5462 4044
rect 5272 3942 5344 4016
tri 5344 3990 5370 4016 nw
tri 5344 3942 5353 3951 sw
rect 5272 3836 5353 3942
tri 5353 3836 5459 3942 sw
rect 5272 3833 5459 3836
tri 5459 3833 5462 3836 sw
tri 2184 1206 2201 1223 sw
rect 1496 1199 2201 1206
tri 2201 1199 2208 1206 sw
rect 1496 1198 2208 1199
tri 2208 1198 2209 1199 sw
rect 890 1175 1207 1194
tri 1207 1175 1226 1194 nw
rect 890 1042 1201 1175
tri 1201 1169 1207 1175 nw
tri 1490 1169 1496 1175 se
rect 1496 1169 5134 1198
tri 1482 1161 1490 1169 se
rect 1490 1161 5134 1169
tri 1471 1150 1482 1161 se
rect 1482 1150 5134 1161
tri 1233 1132 1251 1150 se
rect 1251 1132 5134 1150
tri 5268 1132 5272 1136 se
rect 5272 1132 5462 3833
tri 1229 1128 1233 1132 se
rect 1233 1128 5134 1132
rect 1229 1116 5134 1128
tri 5262 1126 5268 1132 se
rect 5268 1126 5462 1132
tri 5258 1122 5262 1126 se
rect 5262 1122 5462 1126
tri 5252 1116 5258 1122 se
rect 5258 1116 5462 1122
rect 1229 1082 1235 1116
rect 1269 1082 1307 1116
rect 1341 1082 1379 1116
rect 1413 1082 1451 1116
rect 1485 1082 5134 1116
tri 5218 1082 5252 1116 se
rect 5252 1082 5462 1116
rect 1229 1070 5134 1082
tri 1229 1058 1241 1070 ne
rect 1241 1058 1484 1070
tri 1484 1058 1496 1070 nw
tri 2157 1058 2169 1070 ne
rect 2169 1058 5134 1070
tri 5194 1058 5218 1082 se
rect 5218 1058 5462 1082
tri 1241 1053 1246 1058 ne
rect 1246 1053 1479 1058
tri 1479 1053 1484 1058 nw
tri 2169 1053 2174 1058 ne
rect 2174 1053 5134 1058
tri 5189 1053 5194 1058 se
rect 5194 1053 5462 1058
tri 1246 1049 1250 1053 ne
rect 1250 1049 1475 1053
tri 1475 1049 1479 1053 nw
tri 2174 1049 2178 1053 ne
rect 2178 1049 5134 1053
tri 5185 1049 5189 1053 se
rect 5189 1049 5462 1053
tri 1250 1043 1256 1049 ne
rect 1256 1043 1468 1049
tri 1201 1042 1202 1043 sw
tri 1256 1042 1257 1043 ne
rect 1257 1042 1468 1043
tri 1468 1042 1475 1049 nw
tri 2178 1042 2185 1049 ne
rect 2185 1042 5134 1049
tri 5178 1042 5185 1049 se
rect 5185 1042 5462 1049
rect 890 1015 1202 1042
tri 1202 1015 1229 1042 sw
tri 5151 1015 5178 1042 se
rect 5178 1015 5462 1042
rect 890 1014 1229 1015
tri 1229 1014 1230 1015 sw
tri 5150 1014 5151 1015 se
rect 5151 1014 5462 1015
rect 890 960 5462 1014
rect 890 926 5134 960
rect 5168 926 5206 960
rect 5240 926 5278 960
rect 5312 926 5350 960
rect 5384 926 5422 960
rect 5456 926 5462 960
rect 890 893 5462 926
tri 890 882 901 893 ne
rect 901 882 5462 893
tri 5095 879 5098 882 ne
rect 5098 879 5462 882
tri 862 869 872 879 sw
tri 5098 869 5108 879 ne
rect 5108 869 5462 879
rect 569 868 872 869
tri 872 868 873 869 sw
tri 5108 868 5109 869 ne
rect 5109 868 5462 869
rect 569 854 873 868
tri 873 854 887 868 sw
tri 5109 857 5120 868 ne
rect 569 720 5025 854
rect 569 577 862 720
tri 862 695 887 720 nw
tri 5098 695 5120 717 se
rect 5120 695 5462 868
tri 5095 692 5098 695 se
rect 5098 692 5462 695
tri 895 688 899 692 se
rect 899 688 5462 692
tri 891 684 895 688 se
rect 895 684 5462 688
tri 890 683 891 684 se
rect 891 683 5462 684
rect 890 648 5462 683
rect 890 614 5134 648
rect 5168 614 5206 648
rect 5240 614 5278 648
rect 5312 614 5350 648
rect 5384 614 5422 648
rect 5456 614 5462 648
rect 890 602 5462 614
rect 5490 3788 5643 4914
rect 5671 3942 5840 5067
rect 5671 3836 5709 3942
rect 5815 3836 5840 3942
rect 5671 3830 5840 3836
rect 5878 3906 6125 5393
rect 6473 5209 6659 5396
tri 6659 5209 6922 5472 sw
rect 6473 5198 6922 5209
rect 6473 5171 6975 5198
tri 6975 5171 7002 5198 nw
tri 6470 4942 6473 4945 se
rect 6473 4942 6922 5171
tri 6922 5118 6975 5171 nw
tri 6448 4920 6470 4942 se
rect 6470 4920 6922 4942
tri 6225 4913 6232 4920 se
rect 6232 4913 6922 4920
tri 23013 4913 23042 4942 se
rect 23042 4913 23250 5654
rect 23338 5654 25041 5660
rect 23338 5620 23350 5654
rect 23384 5620 23423 5654
rect 23457 5620 23496 5654
rect 23530 5620 23569 5654
rect 23603 5620 23642 5654
rect 23676 5620 23715 5654
rect 23749 5620 23788 5654
rect 23822 5620 23861 5654
rect 23895 5620 23934 5654
rect 23968 5620 24007 5654
rect 24041 5620 24080 5654
rect 24114 5620 24153 5654
rect 24187 5620 24226 5654
rect 24260 5620 24299 5654
rect 24333 5620 24372 5654
rect 24406 5620 24445 5654
rect 24479 5620 24518 5654
rect 24552 5620 24591 5654
rect 24625 5620 24664 5654
rect 24698 5620 24737 5654
rect 24771 5620 24810 5654
rect 24844 5620 24883 5654
rect 24917 5620 24956 5654
rect 24990 5620 25041 5654
rect 23338 5609 25041 5620
tri 25041 5609 25092 5660 sw
tri 25092 5609 25143 5660 ne
rect 25143 5609 25414 5660
rect 23338 5599 25092 5609
tri 25092 5599 25102 5609 sw
tri 25143 5599 25153 5609 ne
rect 25153 5599 25414 5609
rect 23338 5582 25102 5599
tri 25102 5582 25119 5599 sw
tri 25153 5582 25170 5599 ne
rect 25170 5582 25414 5599
rect 23338 5548 23350 5582
rect 23384 5548 23424 5582
rect 23458 5548 23498 5582
rect 23532 5548 23572 5582
rect 23606 5548 23646 5582
rect 23680 5548 23720 5582
rect 23754 5548 23795 5582
rect 23829 5548 23870 5582
rect 23904 5548 23945 5582
rect 23979 5548 24020 5582
rect 24054 5548 24095 5582
rect 24129 5548 24170 5582
rect 24204 5548 24245 5582
rect 24279 5548 24320 5582
rect 24354 5548 24395 5582
rect 24429 5548 24470 5582
rect 24504 5548 24545 5582
rect 24579 5548 24620 5582
rect 24654 5548 24695 5582
rect 24729 5548 24770 5582
rect 24804 5548 24845 5582
rect 24879 5548 24920 5582
rect 24954 5548 24995 5582
rect 25029 5548 25070 5582
rect 25104 5570 25119 5582
tri 25119 5570 25131 5582 sw
tri 25170 5570 25182 5582 ne
rect 25182 5570 25414 5582
rect 25104 5548 25131 5570
rect 23338 5542 25131 5548
tri 25131 5542 25159 5570 sw
tri 25182 5542 25210 5570 ne
tri 24913 5519 24936 5542 ne
rect 24936 5519 25159 5542
tri 25159 5519 25182 5542 sw
tri 24936 5510 24945 5519 ne
rect 24945 5510 25182 5519
tri 24945 5476 24979 5510 ne
rect 24979 5476 25070 5510
rect 25104 5476 25182 5510
tri 24979 5472 24983 5476 ne
rect 24983 5472 25182 5476
tri 24983 5414 25041 5472 ne
rect 25041 5414 25070 5472
tri 25041 5391 25064 5414 ne
tri 6200 4888 6225 4913 se
rect 6225 4888 6922 4913
tri 7245 4888 7270 4913 nw
tri 22988 4888 23013 4913 se
rect 23013 4888 23250 4913
tri 6189 4877 6200 4888 se
rect 6200 4877 6922 4888
tri 22977 4877 22988 4888 se
rect 22988 4877 23250 4888
tri 23250 4877 23331 4958 sw
tri 6153 4841 6189 4877 se
rect 6189 4866 6922 4877
tri 22966 4866 22977 4877 se
rect 22977 4875 23331 4877
tri 23331 4875 23333 4877 sw
rect 22977 4866 23333 4875
rect 6189 4841 6825 4866
rect 6153 4830 6825 4841
rect 6153 3951 6243 4830
tri 6243 4805 6268 4830 nw
tri 6739 4805 6764 4830 ne
rect 6764 4805 6825 4830
tri 6764 4793 6776 4805 ne
rect 6776 4793 6825 4805
tri 22893 4793 22966 4866 se
rect 22966 4810 23333 4866
tri 23333 4810 23398 4875 sw
tri 24332 4810 24397 4875 ne
rect 22966 4793 23398 4810
tri 23398 4793 23415 4810 sw
tri 6776 4765 6804 4793 ne
rect 6804 4776 6825 4793
rect 23042 4746 23250 4793
tri 6243 3951 6263 3971 sw
rect 6153 3948 6263 3951
tri 6263 3948 6266 3951 sw
rect 6153 3935 6266 3948
tri 6266 3935 6279 3948 sw
tri 6153 3923 6165 3935 ne
rect 6165 3923 6279 3935
tri 6125 3906 6142 3923 sw
tri 6165 3906 6182 3923 ne
rect 6182 3906 6279 3923
rect 5878 3886 6142 3906
tri 6142 3886 6162 3906 sw
tri 6182 3886 6202 3906 ne
rect 6202 3898 6279 3906
tri 6279 3898 6316 3935 sw
rect 6202 3886 6316 3898
rect 5878 3866 6162 3886
tri 6162 3866 6182 3886 sw
tri 6202 3866 6222 3886 ne
rect 6222 3866 6269 3886
tri 5643 3788 5668 3813 sw
rect 5490 3620 5850 3788
rect 5490 3586 5504 3620
rect 5538 3586 5576 3620
rect 5610 3586 5648 3620
rect 5682 3586 5720 3620
rect 5754 3586 5792 3620
rect 5826 3586 5850 3620
rect 5490 2364 5850 3586
rect 5490 2330 5504 2364
rect 5538 2330 5576 2364
rect 5610 2330 5648 2364
rect 5682 2330 5720 2364
rect 5754 2330 5792 2364
rect 5826 2330 5850 2364
rect 5490 2052 5850 2330
rect 5490 2018 5504 2052
rect 5538 2018 5576 2052
rect 5610 2018 5648 2052
rect 5682 2018 5720 2052
rect 5754 2018 5792 2052
rect 5826 2018 5850 2052
rect 5490 1740 5850 2018
rect 5490 1706 5504 1740
rect 5538 1706 5576 1740
rect 5610 1706 5648 1740
rect 5682 1706 5720 1740
rect 5754 1706 5792 1740
rect 5826 1706 5850 1740
rect 5490 1428 5850 1706
rect 5490 1394 5504 1428
rect 5538 1394 5576 1428
rect 5610 1394 5648 1428
rect 5682 1394 5720 1428
rect 5754 1394 5792 1428
rect 5826 1394 5850 1428
rect 5490 1116 5850 1394
rect 5490 1082 5504 1116
rect 5538 1082 5576 1116
rect 5610 1082 5648 1116
rect 5682 1082 5720 1116
rect 5754 1082 5792 1116
rect 5826 1082 5850 1116
rect 5490 804 5850 1082
rect 5490 770 5504 804
rect 5538 770 5576 804
rect 5610 770 5648 804
rect 5682 770 5720 804
rect 5754 770 5792 804
rect 5826 770 5850 804
tri 862 577 875 590 sw
tri 5477 577 5490 590 se
rect 5490 577 5850 770
rect 569 576 875 577
tri 875 576 876 577 sw
tri 5476 576 5477 577 se
rect 5477 576 5850 577
rect 569 565 876 576
tri 876 565 887 576 sw
tri 5465 565 5476 576 se
rect 5476 565 5850 576
rect 569 466 5850 565
tri 569 465 570 466 ne
rect 570 465 5850 466
rect 457 417 463 451
rect 497 417 503 451
tri 570 431 604 465 ne
rect 604 431 5850 465
tri 604 430 605 431 ne
rect 605 430 5850 431
rect 457 405 503 417
tri 605 405 630 430 ne
rect 630 405 5850 430
tri 630 398 637 405 ne
rect 637 398 5850 405
tri 4805 396 4807 398 ne
rect 4807 396 5850 398
tri 4807 395 4808 396 ne
rect 4808 395 5850 396
rect 361 349 367 383
rect 401 370 407 383
tri 407 370 432 395 sw
tri 4808 370 4833 395 ne
rect 4833 394 5850 395
rect 4833 370 5026 394
rect 401 364 4711 370
tri 4833 369 4834 370 ne
rect 401 349 541 364
rect 361 330 541 349
rect 575 330 614 364
rect 648 330 687 364
rect 721 330 760 364
rect 794 330 833 364
rect 867 330 906 364
rect 940 330 979 364
rect 1013 330 1052 364
rect 1086 330 1125 364
rect 1159 330 1198 364
rect 1232 330 1271 364
rect 1305 330 1344 364
rect 1378 330 1417 364
rect 1451 330 1490 364
rect 1524 330 1563 364
rect 1597 330 1636 364
rect 1670 330 1709 364
rect 1743 330 1782 364
rect 1816 330 1855 364
rect 1889 330 1928 364
rect 1962 330 2000 364
rect 2034 330 2072 364
rect 2106 330 2144 364
rect 2178 330 2216 364
rect 2250 330 2288 364
rect 2322 330 2360 364
rect 2394 330 2432 364
rect 2466 330 2504 364
rect 2538 330 2576 364
rect 2610 330 2648 364
rect 2682 330 2720 364
rect 2754 330 2792 364
rect 2826 330 2864 364
rect 2898 330 2936 364
rect 2970 330 3008 364
rect 3042 330 3080 364
rect 3114 330 3152 364
rect 3186 330 3224 364
rect 3258 330 3296 364
rect 3330 330 3368 364
rect 3402 330 3440 364
rect 3474 330 3512 364
rect 3546 330 3584 364
rect 3618 330 3656 364
rect 3690 330 3728 364
rect 3762 330 3800 364
rect 3834 330 3872 364
rect 3906 330 3944 364
rect 3978 330 4016 364
rect 4050 330 4088 364
rect 4122 330 4160 364
rect 4194 330 4232 364
rect 4266 330 4304 364
rect 4338 330 4376 364
rect 4410 330 4448 364
rect 4482 330 4520 364
rect 4554 330 4592 364
rect 4626 330 4664 364
rect 4698 330 4711 364
rect 361 314 4711 330
rect 4834 322 5026 370
tri 5026 369 5051 394 nw
tri 5633 369 5658 394 ne
rect 5658 322 5850 394
rect 5878 577 6182 3866
tri 6222 3852 6236 3866 ne
rect 6236 3852 6269 3866
rect 6303 3852 6316 3886
tri 6236 3830 6258 3852 ne
rect 6258 3830 6316 3852
tri 6258 3825 6263 3830 ne
rect 6263 3825 6316 3830
tri 6316 3825 6389 3898 sw
rect 5879 575 6181 576
rect 5878 539 6182 575
rect 5879 538 6181 539
rect 5878 430 6182 537
rect 6263 3814 6389 3825
rect 6263 3780 6269 3814
rect 6303 3780 6389 3814
rect 6263 3744 6389 3780
tri 6389 3744 6470 3825 sw
rect 6263 3742 6924 3744
rect 6263 3708 6269 3742
rect 6303 3708 6924 3742
rect 6263 3670 6924 3708
rect 6263 3636 6269 3670
rect 6303 3654 6924 3670
rect 6303 3636 6349 3654
rect 6263 3632 6349 3636
tri 6349 3632 6371 3654 nw
tri 6735 3632 6757 3654 ne
rect 6757 3632 6924 3654
rect 6263 3598 6309 3632
rect 6263 3564 6269 3598
rect 6303 3564 6309 3598
tri 6309 3592 6349 3632 nw
tri 6757 3592 6797 3632 ne
rect 6797 3592 6924 3632
tri 6797 3583 6806 3592 ne
rect 6263 3526 6309 3564
rect 6263 3492 6269 3526
rect 6303 3492 6309 3526
rect 6263 3454 6309 3492
rect 6263 3420 6269 3454
rect 6303 3420 6309 3454
rect 6263 3382 6309 3420
rect 6263 3348 6269 3382
rect 6303 3348 6309 3382
rect 6263 3310 6309 3348
rect 6263 3276 6269 3310
rect 6303 3276 6309 3310
rect 6263 3238 6309 3276
rect 6263 3204 6269 3238
rect 6303 3204 6309 3238
rect 6263 3166 6309 3204
rect 6263 3132 6269 3166
rect 6303 3132 6309 3166
rect 6263 3093 6309 3132
rect 6263 3059 6269 3093
rect 6303 3059 6309 3093
rect 6263 3020 6309 3059
rect 6263 2986 6269 3020
rect 6303 2986 6309 3020
rect 6263 2947 6309 2986
rect 6263 2913 6269 2947
rect 6303 2913 6309 2947
rect 6263 2874 6309 2913
rect 6263 2840 6269 2874
rect 6303 2840 6309 2874
rect 6263 2801 6309 2840
rect 6263 2767 6269 2801
rect 6303 2767 6309 2801
rect 6263 2728 6309 2767
rect 6263 2694 6269 2728
rect 6303 2694 6309 2728
rect 6263 2655 6309 2694
rect 6263 2621 6269 2655
rect 6303 2621 6309 2655
rect 6263 2582 6309 2621
rect 6263 2548 6269 2582
rect 6303 2548 6309 2582
rect 6263 2509 6309 2548
rect 6263 2475 6269 2509
rect 6303 2475 6309 2509
rect 6263 2436 6309 2475
rect 6263 2402 6269 2436
rect 6303 2402 6309 2436
rect 6263 2363 6309 2402
rect 6263 2329 6269 2363
rect 6303 2329 6309 2363
rect 6263 2290 6309 2329
rect 6263 2256 6269 2290
rect 6303 2256 6309 2290
rect 6263 2217 6309 2256
rect 6263 2183 6269 2217
rect 6303 2183 6309 2217
rect 6263 2144 6309 2183
rect 6263 2110 6269 2144
rect 6303 2110 6309 2144
rect 6263 2071 6309 2110
rect 6263 2037 6269 2071
rect 6303 2037 6309 2071
rect 6263 1998 6309 2037
rect 6263 1964 6269 1998
rect 6303 1964 6309 1998
rect 6263 1925 6309 1964
rect 6263 1891 6269 1925
rect 6303 1891 6309 1925
rect 6263 1852 6309 1891
rect 6263 1818 6269 1852
rect 6303 1818 6309 1852
rect 6263 1779 6309 1818
rect 6263 1745 6269 1779
rect 6303 1745 6309 1779
rect 6263 1706 6309 1745
rect 6263 1672 6269 1706
rect 6303 1672 6309 1706
rect 6263 1633 6309 1672
rect 6263 1599 6269 1633
rect 6303 1599 6309 1633
rect 6263 1560 6309 1599
rect 6263 1526 6269 1560
rect 6303 1526 6309 1560
rect 6263 1487 6309 1526
rect 6263 1453 6269 1487
rect 6303 1453 6309 1487
rect 6263 1414 6309 1453
rect 6263 1380 6269 1414
rect 6303 1380 6309 1414
rect 6263 1341 6309 1380
rect 6263 1307 6269 1341
rect 6303 1307 6309 1341
rect 6263 1268 6309 1307
rect 6263 1234 6269 1268
rect 6303 1234 6309 1268
rect 6263 1195 6309 1234
rect 6263 1161 6269 1195
rect 6303 1161 6309 1195
rect 6263 1122 6309 1161
rect 6263 1088 6269 1122
rect 6303 1088 6309 1122
rect 6263 1049 6309 1088
rect 6263 1015 6269 1049
rect 6303 1019 6309 1049
rect 6481 3537 6599 3549
rect 6481 3503 6487 3537
rect 6521 3503 6559 3537
rect 6593 3503 6599 3537
rect 6481 3462 6599 3503
rect 6481 3428 6487 3462
rect 6521 3428 6559 3462
rect 6593 3428 6599 3462
rect 6481 3387 6599 3428
rect 6481 3353 6487 3387
rect 6521 3353 6559 3387
rect 6593 3353 6599 3387
rect 6481 3312 6599 3353
rect 6481 3278 6487 3312
rect 6521 3278 6559 3312
rect 6593 3278 6599 3312
rect 6481 3238 6599 3278
rect 6481 3204 6487 3238
rect 6521 3204 6559 3238
rect 6593 3204 6599 3238
rect 6481 3164 6599 3204
rect 6481 3130 6487 3164
rect 6521 3130 6559 3164
rect 6593 3130 6599 3164
rect 6481 3090 6599 3130
rect 6481 3056 6487 3090
rect 6521 3056 6559 3090
rect 6593 3056 6599 3090
rect 6481 3016 6599 3056
rect 6481 2982 6487 3016
rect 6521 2982 6559 3016
rect 6593 2982 6599 3016
rect 6481 2942 6599 2982
rect 6481 2908 6487 2942
rect 6521 2908 6559 2942
rect 6593 2908 6599 2942
rect 6481 2868 6599 2908
rect 6481 2834 6487 2868
rect 6521 2834 6559 2868
rect 6593 2834 6599 2868
rect 6481 2794 6599 2834
rect 6481 2760 6487 2794
rect 6521 2760 6559 2794
rect 6593 2760 6599 2794
rect 6481 2720 6599 2760
rect 6481 2686 6487 2720
rect 6521 2686 6559 2720
rect 6593 2686 6599 2720
rect 6481 2646 6599 2686
rect 6481 2612 6487 2646
rect 6521 2612 6559 2646
rect 6593 2612 6599 2646
rect 6481 2572 6599 2612
rect 6481 2538 6487 2572
rect 6521 2538 6559 2572
rect 6593 2538 6599 2572
rect 6481 2498 6599 2538
rect 6481 2464 6487 2498
rect 6521 2464 6559 2498
rect 6593 2464 6599 2498
rect 6481 2424 6599 2464
rect 6481 2390 6487 2424
rect 6521 2390 6559 2424
rect 6593 2390 6599 2424
rect 6481 2350 6599 2390
rect 6481 2316 6487 2350
rect 6521 2316 6559 2350
rect 6593 2316 6599 2350
rect 6481 2276 6599 2316
rect 6481 2242 6487 2276
rect 6521 2242 6559 2276
rect 6593 2242 6599 2276
rect 6481 2202 6599 2242
rect 6481 2168 6487 2202
rect 6521 2168 6559 2202
rect 6593 2168 6599 2202
rect 6481 2128 6599 2168
rect 6481 2094 6487 2128
rect 6521 2094 6559 2128
rect 6593 2094 6599 2128
rect 6481 2054 6599 2094
rect 6481 2020 6487 2054
rect 6521 2020 6559 2054
rect 6593 2020 6599 2054
rect 6481 1980 6599 2020
rect 6481 1946 6487 1980
rect 6521 1946 6559 1980
rect 6593 1946 6599 1980
rect 6481 1906 6599 1946
rect 6481 1872 6487 1906
rect 6521 1872 6559 1906
rect 6593 1872 6599 1906
rect 6481 1832 6599 1872
rect 6481 1798 6487 1832
rect 6521 1798 6559 1832
rect 6593 1798 6599 1832
rect 6481 1758 6599 1798
rect 6481 1724 6487 1758
rect 6521 1724 6559 1758
rect 6593 1724 6599 1758
rect 6481 1684 6599 1724
rect 6481 1650 6487 1684
rect 6521 1650 6559 1684
rect 6593 1650 6599 1684
rect 6481 1610 6599 1650
rect 6481 1576 6487 1610
rect 6521 1576 6559 1610
rect 6593 1576 6599 1610
rect 6481 1536 6599 1576
rect 6481 1502 6487 1536
rect 6521 1502 6559 1536
rect 6593 1502 6599 1536
rect 6481 1462 6599 1502
rect 6481 1428 6487 1462
rect 6521 1428 6559 1462
rect 6593 1428 6599 1462
rect 6481 1388 6599 1428
rect 6481 1354 6487 1388
rect 6521 1354 6559 1388
rect 6593 1354 6599 1388
rect 6481 1314 6599 1354
rect 6481 1280 6487 1314
rect 6521 1280 6559 1314
rect 6593 1280 6599 1314
rect 6481 1240 6599 1280
rect 6481 1206 6487 1240
rect 6521 1206 6559 1240
rect 6593 1206 6599 1240
rect 6481 1166 6599 1206
rect 6481 1132 6487 1166
rect 6521 1132 6559 1166
rect 6593 1132 6599 1166
rect 6481 1092 6599 1132
rect 6481 1058 6487 1092
rect 6521 1058 6559 1092
rect 6593 1058 6599 1092
tri 6309 1019 6317 1027 sw
rect 6303 1018 6317 1019
tri 6317 1018 6318 1019 sw
rect 6481 1018 6599 1058
tri 6798 1019 6806 1027 se
rect 6806 1019 6924 3592
rect 6303 1015 6318 1018
rect 6263 984 6318 1015
tri 6318 984 6352 1018 sw
rect 6481 984 6487 1018
rect 6521 984 6559 1018
rect 6593 984 6599 1018
tri 6793 1014 6798 1019 se
rect 6798 1014 6924 1019
rect 6263 980 6352 984
tri 6352 980 6356 984 sw
rect 6263 976 6356 980
rect 6263 942 6269 976
rect 6303 972 6356 976
tri 6356 972 6364 980 sw
rect 6481 972 6599 984
tri 6759 980 6793 1014 se
rect 6793 980 6924 1014
tri 6751 972 6759 980 se
rect 6759 972 6924 980
rect 6303 946 6364 972
tri 6364 946 6390 972 sw
tri 6725 946 6751 972 se
rect 6751 946 6924 972
rect 6303 942 6390 946
rect 6263 941 6390 942
tri 6390 941 6395 946 sw
tri 6720 941 6725 946 se
rect 6725 941 6924 946
rect 6263 914 6395 941
tri 6395 914 6422 941 sw
tri 6693 914 6720 941 se
rect 6720 914 6924 941
rect 6263 907 6422 914
tri 6422 907 6429 914 sw
tri 6686 907 6693 914 se
rect 6693 907 6924 914
rect 6263 903 6429 907
rect 6263 869 6269 903
rect 6303 902 6429 903
tri 6429 902 6434 907 sw
tri 6681 902 6686 907 se
rect 6686 902 6924 907
rect 6303 869 6924 902
rect 6263 830 6924 869
rect 6263 796 6269 830
rect 6303 796 6924 830
rect 6263 757 6924 796
rect 6263 723 6269 757
rect 6303 723 6924 757
rect 6263 684 6924 723
rect 6263 650 6269 684
rect 6303 650 6924 684
rect 6263 611 6924 650
rect 6263 577 6269 611
rect 6303 577 6924 611
rect 6263 538 6924 577
rect 6263 504 6269 538
rect 6303 504 6924 538
rect 6263 465 6924 504
rect 6263 431 6269 465
rect 6303 431 6924 465
tri 6182 430 6183 431 sw
rect 5878 405 6183 430
tri 6183 405 6208 430 sw
rect 5878 396 6208 405
tri 6208 396 6217 405 sw
rect 5878 367 6217 396
tri 6217 367 6246 396 sw
rect 6263 390 6924 431
tri 6263 375 6278 390 ne
rect 6278 375 6924 390
rect 25064 3316 25070 5414
rect 25176 3316 25182 5472
rect 25064 3312 25182 3316
rect 25064 3278 25142 3312
rect 25176 3278 25182 3312
rect 25064 3277 25182 3278
rect 25064 3243 25070 3277
rect 25104 3243 25182 3277
rect 25064 3240 25182 3243
rect 25064 3206 25142 3240
rect 25176 3206 25182 3240
rect 25064 3204 25182 3206
rect 25064 3170 25070 3204
rect 25104 3170 25182 3204
rect 25064 3168 25182 3170
rect 25064 3134 25142 3168
rect 25176 3134 25182 3168
rect 25064 3131 25182 3134
rect 25064 3097 25070 3131
rect 25104 3097 25182 3131
rect 25064 3096 25182 3097
rect 25064 3062 25142 3096
rect 25176 3062 25182 3096
rect 25064 3058 25182 3062
rect 25064 3024 25070 3058
rect 25104 3024 25182 3058
rect 25064 2990 25142 3024
rect 25176 2990 25182 3024
rect 25064 2985 25182 2990
rect 25064 2951 25070 2985
rect 25104 2951 25182 2985
rect 25064 2917 25142 2951
rect 25176 2917 25182 2951
rect 25064 2912 25182 2917
rect 25064 2878 25070 2912
rect 25104 2878 25182 2912
rect 25064 2844 25142 2878
rect 25176 2844 25182 2878
rect 25064 2839 25182 2844
rect 25064 2805 25070 2839
rect 25104 2805 25182 2839
rect 25064 2771 25142 2805
rect 25176 2771 25182 2805
rect 25064 2766 25182 2771
rect 25064 2732 25070 2766
rect 25104 2732 25182 2766
rect 25064 2698 25142 2732
rect 25176 2698 25182 2732
rect 25064 2693 25182 2698
rect 25064 2659 25070 2693
rect 25104 2659 25182 2693
rect 25064 2625 25142 2659
rect 25176 2625 25182 2659
rect 25064 2620 25182 2625
rect 25064 2586 25070 2620
rect 25104 2586 25182 2620
rect 25064 2552 25142 2586
rect 25176 2552 25182 2586
rect 25064 2547 25182 2552
rect 25064 2513 25070 2547
rect 25104 2513 25182 2547
rect 25064 2479 25142 2513
rect 25176 2479 25182 2513
rect 25064 2474 25182 2479
rect 25064 2440 25070 2474
rect 25104 2440 25182 2474
rect 25064 2406 25142 2440
rect 25176 2406 25182 2440
rect 25064 2401 25182 2406
rect 25064 2367 25070 2401
rect 25104 2367 25182 2401
rect 25064 2333 25142 2367
rect 25176 2333 25182 2367
rect 25064 2328 25182 2333
rect 25064 2294 25070 2328
rect 25104 2294 25182 2328
rect 25064 2260 25142 2294
rect 25176 2260 25182 2294
rect 25064 2255 25182 2260
rect 25064 2221 25070 2255
rect 25104 2221 25182 2255
rect 25064 2187 25142 2221
rect 25176 2187 25182 2221
rect 25064 2182 25182 2187
rect 25064 2148 25070 2182
rect 25104 2148 25182 2182
rect 25064 2114 25142 2148
rect 25176 2114 25182 2148
rect 25064 2109 25182 2114
rect 25064 2075 25070 2109
rect 25104 2075 25182 2109
rect 25064 2041 25142 2075
rect 25176 2041 25182 2075
rect 25064 2036 25182 2041
rect 25064 2002 25070 2036
rect 25104 2002 25182 2036
rect 25064 1968 25142 2002
rect 25176 1968 25182 2002
rect 25064 1963 25182 1968
rect 25064 1929 25070 1963
rect 25104 1929 25182 1963
rect 25064 1895 25142 1929
rect 25176 1895 25182 1929
rect 25064 1890 25182 1895
rect 25064 1856 25070 1890
rect 25104 1856 25182 1890
rect 25064 1822 25142 1856
rect 25176 1822 25182 1856
rect 25064 1817 25182 1822
rect 25064 1783 25070 1817
rect 25104 1783 25182 1817
rect 25064 1749 25142 1783
rect 25176 1749 25182 1783
rect 25064 1744 25182 1749
rect 25064 1710 25070 1744
rect 25104 1710 25182 1744
rect 25064 1676 25142 1710
rect 25176 1676 25182 1710
rect 25064 1671 25182 1676
rect 25064 1637 25070 1671
rect 25104 1637 25182 1671
rect 25064 1603 25142 1637
rect 25176 1603 25182 1637
rect 25064 1598 25182 1603
rect 25064 1564 25070 1598
rect 25104 1564 25182 1598
rect 25064 1530 25142 1564
rect 25176 1530 25182 1564
rect 25064 1525 25182 1530
rect 25064 1491 25070 1525
rect 25104 1491 25182 1525
rect 25064 1457 25142 1491
rect 25176 1457 25182 1491
rect 25064 1452 25182 1457
rect 25064 1418 25070 1452
rect 25104 1418 25182 1452
rect 25064 1384 25142 1418
rect 25176 1384 25182 1418
rect 25064 1379 25182 1384
rect 25064 1345 25070 1379
rect 25104 1345 25182 1379
rect 25064 1311 25142 1345
rect 25176 1311 25182 1345
rect 25064 1306 25182 1311
rect 25064 1272 25070 1306
rect 25104 1272 25182 1306
rect 25064 1238 25142 1272
rect 25176 1238 25182 1272
rect 25064 1233 25182 1238
rect 25064 1199 25070 1233
rect 25104 1199 25182 1233
rect 25064 1165 25142 1199
rect 25176 1165 25182 1199
rect 25064 1160 25182 1165
rect 25064 1126 25070 1160
rect 25104 1126 25182 1160
rect 25064 1092 25142 1126
rect 25176 1092 25182 1126
rect 25064 1087 25182 1092
rect 25064 1053 25070 1087
rect 25104 1053 25182 1087
rect 25064 1019 25142 1053
rect 25176 1019 25182 1053
rect 25064 1014 25182 1019
rect 25064 980 25070 1014
rect 25104 980 25182 1014
rect 25064 946 25142 980
rect 25176 946 25182 980
rect 25064 941 25182 946
rect 25064 907 25070 941
rect 25104 907 25182 941
rect 25064 873 25142 907
rect 25176 873 25182 907
rect 25064 868 25182 873
rect 25064 834 25070 868
rect 25104 834 25182 868
rect 25064 800 25142 834
rect 25176 800 25182 834
rect 25064 795 25182 800
rect 25064 761 25070 795
rect 25104 761 25182 795
rect 25064 727 25142 761
rect 25176 727 25182 761
rect 25064 722 25182 727
rect 25064 688 25070 722
rect 25104 688 25182 722
rect 25064 654 25142 688
rect 25176 654 25182 688
rect 25064 649 25182 654
rect 25064 615 25070 649
rect 25104 615 25182 649
rect 25064 581 25142 615
rect 25176 581 25182 615
rect 25064 576 25182 581
rect 25064 542 25070 576
rect 25104 542 25182 576
rect 25064 508 25142 542
rect 25176 508 25182 542
rect 25064 503 25182 508
rect 25064 482 25070 503
rect 25104 482 25182 503
tri 3137 298 3153 314 ne
rect 3153 298 3181 314
tri 316 289 325 298 sw
tri 3153 289 3162 298 ne
rect 3162 289 3181 298
rect 264 284 325 289
tri 325 284 330 289 sw
tri 3162 284 3167 289 ne
rect 3167 284 3181 289
rect 264 280 330 284
tri 330 280 334 284 sw
tri 3167 280 3171 284 ne
rect 3171 280 3181 284
rect 264 274 334 280
tri 334 274 340 280 sw
rect 665 274 795 280
rect 264 267 340 274
tri 340 267 347 274 sw
rect 264 232 519 267
tri 264 223 273 232 ne
rect 273 223 519 232
tri 519 223 563 267 sw
rect 71 174 189 213
rect 71 140 77 174
rect 111 140 149 174
rect 183 140 189 174
tri 273 171 325 223 ne
rect 325 171 563 223
tri 541 168 544 171 ne
rect 544 168 563 171
tri 563 168 618 223 sw
rect 665 168 677 274
rect 783 168 795 274
tri 3171 270 3181 280 ne
rect 3949 289 3968 314
tri 3968 289 3993 314 nw
tri 4302 289 4327 314 ne
rect 4327 289 4357 314
tri 4357 289 4382 314 nw
rect 3949 284 3963 289
tri 3963 284 3968 289 nw
rect 3949 280 3959 284
tri 3959 280 3963 284 nw
tri 3949 270 3959 280 nw
tri 544 149 563 168 ne
rect 563 162 618 168
tri 618 162 624 168 sw
rect 665 162 795 168
rect 563 149 624 162
tri 624 149 637 162 sw
tri 563 143 569 149 ne
rect 569 143 637 149
tri 569 142 570 143 ne
rect 570 142 637 143
rect 71 114 189 140
tri 570 138 574 142 ne
rect 574 138 637 142
tri 574 128 584 138 ne
rect 584 128 637 138
tri 584 127 585 128 ne
rect 585 114 637 128
rect 665 143 723 162
tri 723 143 742 162 nw
rect 665 142 722 143
tri 722 142 723 143 nw
rect 5878 142 6246 367
tri 6431 362 6444 375 ne
rect 6444 362 6712 375
tri 6712 362 6725 375 nw
rect 25180 366 25182 482
rect 25064 362 25142 366
rect 25176 362 25182 366
tri 6444 357 6449 362 ne
rect 6449 357 6707 362
tri 6707 357 6712 362 nw
rect 25064 357 25182 362
tri 6449 324 6482 357 ne
rect 6482 322 6674 357
tri 6674 324 6707 357 nw
rect 25064 323 25070 357
rect 25104 323 25182 357
rect 25064 289 25142 323
rect 25176 289 25182 323
rect 25064 284 25182 289
rect 25064 250 25070 284
rect 25104 250 25182 284
rect 6815 142 7562 196
rect 8053 170 8799 224
rect 10938 170 11684 224
rect 12176 170 12922 224
rect 16298 170 17044 224
rect 25064 216 25142 250
rect 25176 216 25182 250
rect 25064 211 25182 216
rect 25064 177 25070 211
rect 25104 177 25182 211
tri 25039 144 25064 169 se
rect 25064 144 25142 177
rect 24401 143 25142 144
rect 25176 143 25182 177
rect 665 138 718 142
tri 718 138 722 142 nw
rect 24401 138 25182 143
rect 665 114 717 138
tri 717 137 718 138 nw
rect 24401 104 24413 138
rect 24447 104 24486 138
rect 24520 104 24559 138
rect 24593 104 24632 138
rect 24666 104 24705 138
rect 24739 104 24778 138
rect 24812 104 24851 138
rect 24885 104 24924 138
rect 24958 104 24997 138
rect 25031 104 25070 138
rect 25104 104 25182 138
rect 24401 70 25142 104
rect 25176 70 25182 104
rect 24401 66 25182 70
rect 24401 32 24456 66
rect 24490 32 24528 66
rect 24562 32 24600 66
rect 24634 32 24672 66
rect 24706 32 24744 66
rect 24778 32 24816 66
rect 24850 32 24888 66
rect 24922 32 24960 66
rect 24994 32 25032 66
rect 25066 32 25182 66
rect 24401 26 25182 32
rect 25210 461 25414 5570
rect 25211 459 25413 460
rect 25210 423 25414 459
rect 25211 422 25413 423
rect 25210 119 25414 421
rect 25442 214 25494 5917
rect 25522 214 25574 5951
rect 25602 214 25654 5985
rect 25682 214 25734 6019
rect 25786 915 25792 6133
rect 25898 915 25904 6133
rect 25786 876 25904 915
rect 25786 842 25792 876
rect 25826 842 25864 876
rect 25898 842 25904 876
rect 25786 803 25904 842
rect 25786 769 25792 803
rect 25826 769 25864 803
rect 25898 769 25904 803
rect 25786 730 25904 769
rect 25786 696 25792 730
rect 25826 696 25864 730
rect 25898 696 25904 730
rect 25786 657 25904 696
rect 25786 623 25792 657
rect 25826 623 25864 657
rect 25898 623 25904 657
rect 25786 584 25904 623
rect 25786 550 25792 584
rect 25826 550 25864 584
rect 25898 550 25904 584
rect 25786 511 25904 550
rect 25786 482 25792 511
rect 25826 482 25864 511
rect 25898 482 25904 511
rect 25786 366 25787 482
rect 25903 366 25904 482
rect 25786 365 25904 366
rect 25786 331 25792 365
rect 25826 331 25864 365
rect 25898 331 25904 365
rect 25786 292 25904 331
rect 25786 258 25792 292
rect 25826 258 25864 292
rect 25898 258 25904 292
rect 25786 219 25904 258
rect 25210 3 25222 119
rect 25402 9 25414 119
rect 25786 185 25792 219
rect 25826 185 25864 219
rect 25898 185 25904 219
rect 25786 146 25904 185
rect 25786 112 25792 146
rect 25826 112 25864 146
rect 25898 112 25904 146
rect 25786 73 25904 112
rect 25786 39 25792 73
rect 25826 39 25864 73
rect 25898 39 25904 73
rect 25786 27 25904 39
rect 26175 6142 26181 6176
rect 26215 6142 26253 6176
rect 26287 6142 26293 6176
rect 26175 6103 26293 6142
rect 26175 6069 26181 6103
rect 26215 6069 26253 6103
rect 26287 6069 26293 6103
rect 26175 6030 26293 6069
rect 26175 5996 26181 6030
rect 26215 5996 26253 6030
rect 26287 5996 26293 6030
rect 26175 5957 26293 5996
rect 26175 5923 26181 5957
rect 26215 5923 26253 5957
rect 26287 5923 26293 5957
rect 26175 5884 26293 5923
rect 26175 5850 26181 5884
rect 26215 5850 26253 5884
rect 26287 5850 26293 5884
rect 26175 5811 26293 5850
rect 26175 5777 26181 5811
rect 26215 5777 26253 5811
rect 26287 5777 26293 5811
rect 26175 5738 26293 5777
rect 26175 5704 26181 5738
rect 26215 5704 26253 5738
rect 26287 5704 26293 5738
rect 26175 5665 26293 5704
rect 26175 5631 26181 5665
rect 26215 5631 26253 5665
rect 26287 5631 26293 5665
rect 26175 5592 26293 5631
rect 26175 5558 26181 5592
rect 26215 5558 26253 5592
rect 26287 5558 26293 5592
rect 26175 5519 26293 5558
rect 26175 5485 26181 5519
rect 26215 5485 26253 5519
rect 26287 5485 26293 5519
rect 26175 5446 26293 5485
rect 26175 5412 26181 5446
rect 26215 5412 26253 5446
rect 26287 5412 26293 5446
rect 26175 5373 26293 5412
rect 26175 5339 26181 5373
rect 26215 5339 26253 5373
rect 26287 5339 26293 5373
rect 26175 5300 26293 5339
rect 26175 5266 26181 5300
rect 26215 5266 26253 5300
rect 26287 5266 26293 5300
rect 26175 5227 26293 5266
rect 26175 5193 26181 5227
rect 26215 5193 26253 5227
rect 26287 5193 26293 5227
rect 26175 5154 26293 5193
rect 26175 5120 26181 5154
rect 26215 5120 26253 5154
rect 26287 5120 26293 5154
rect 26175 5081 26293 5120
rect 26175 5047 26181 5081
rect 26215 5047 26253 5081
rect 26287 5047 26293 5081
rect 26175 5008 26293 5047
rect 26175 4974 26181 5008
rect 26215 4974 26253 5008
rect 26287 4974 26293 5008
rect 26175 4935 26293 4974
rect 26175 4901 26181 4935
rect 26215 4901 26253 4935
rect 26287 4901 26293 4935
rect 26175 4862 26293 4901
rect 26175 4828 26181 4862
rect 26215 4828 26253 4862
rect 26287 4828 26293 4862
rect 26175 4789 26293 4828
rect 26175 4755 26181 4789
rect 26215 4755 26253 4789
rect 26287 4755 26293 4789
rect 26175 4716 26293 4755
rect 26175 4682 26181 4716
rect 26215 4682 26253 4716
rect 26287 4682 26293 4716
rect 26175 4643 26293 4682
rect 26175 4609 26181 4643
rect 26215 4609 26253 4643
rect 26287 4609 26293 4643
rect 26175 4570 26293 4609
rect 26175 4536 26181 4570
rect 26215 4536 26253 4570
rect 26287 4536 26293 4570
rect 26175 4497 26293 4536
rect 26175 4463 26181 4497
rect 26215 4463 26253 4497
rect 26287 4463 26293 4497
rect 26175 4424 26293 4463
rect 26175 4390 26181 4424
rect 26215 4390 26253 4424
rect 26287 4390 26293 4424
rect 26175 4351 26293 4390
rect 25402 3 25408 9
tri 25408 3 25414 9 nw
rect 26175 -147 26181 4351
rect 26287 -147 26293 4351
rect 26175 -159 26293 -147
tri 24059 -4169 24175 -4053 se
rect 24175 -4169 24181 -4053
rect 24297 -4169 24321 -4053
tri 24028 -4200 24059 -4169 se
rect 24059 -4200 24290 -4169
tri 24290 -4200 24321 -4169 nw
rect 22237 -4316 22243 -4200
rect 22359 -4316 24174 -4200
tri 24174 -4316 24290 -4200 nw
rect 23459 -4514 23517 -4450
rect 16643 -8556 16771 -8437
rect 16995 -8910 17113 -8838
<< rmetal1 >>
rect 2797 4860 2799 4861
rect 2835 4860 2837 4861
rect 2797 4516 2798 4860
rect 2836 4516 2837 4860
rect 2797 4515 2799 4516
rect 2835 4515 2837 4516
rect 2301 4364 2303 4365
rect 2339 4364 2341 4365
rect 2301 4020 2302 4364
rect 2340 4020 2341 4364
rect 2301 4019 2303 4020
rect 2339 4019 2341 4020
rect 888 2671 1104 2672
tri 1104 2671 1105 2672 sw
tri 1103 2670 1104 2671 ne
rect 1104 2670 1105 2671
tri 1105 2670 1106 2671 sw
tri 1104 2668 1106 2670 ne
tri 1106 2668 1108 2670 sw
tri 1106 2666 1108 2668 ne
tri 1108 2666 1110 2668 sw
tri 1108 2664 1110 2666 ne
tri 1110 2664 1112 2666 sw
tri 1110 2662 1112 2664 ne
tri 1112 2662 1114 2664 sw
tri 1112 2660 1114 2662 ne
tri 1114 2660 1116 2662 sw
tri 1114 2659 1115 2660 ne
rect 1115 2659 1116 2660
tri 1116 2659 1117 2660 sw
tri 1115 2658 1116 2659 ne
rect 1116 2658 1117 2659
tri 1117 2658 1118 2659 sw
rect 888 2642 1080 2643
rect 1078 2641 1080 2642
rect 1116 2641 1118 2658
rect 1078 2585 1079 2641
rect 1117 2585 1118 2641
rect 1078 2584 1080 2585
rect 888 2583 1080 2584
rect 1116 2568 1118 2585
tri 1114 2566 1116 2568 se
tri 1116 2566 1118 2568 nw
tri 1113 2565 1114 2566 se
rect 1114 2565 1115 2566
tri 1115 2565 1116 2566 nw
tri 1112 2564 1113 2565 se
rect 1113 2564 1114 2565
tri 1114 2564 1115 2565 nw
tri 1110 2562 1112 2564 se
tri 1112 2562 1114 2564 nw
tri 1108 2560 1110 2562 se
tri 1110 2560 1112 2562 nw
tri 1106 2558 1108 2560 se
tri 1108 2558 1110 2560 nw
tri 1104 2556 1106 2558 se
tri 1106 2556 1108 2558 nw
tri 1103 2555 1104 2556 se
rect 1104 2555 1105 2556
tri 1105 2555 1106 2556 nw
rect 888 2554 1104 2555
tri 1104 2554 1105 2555 nw
rect 888 2417 1203 2418
rect 888 2416 889 2417
rect 1202 2416 1203 2417
rect 888 2379 889 2380
rect 1202 2379 1203 2380
rect 888 2378 1203 2379
rect 5296 4876 5298 4877
rect 5334 4876 5336 4877
rect 5296 4516 5297 4876
rect 5335 4516 5336 4876
rect 5296 4515 5298 4516
rect 5334 4515 5336 4516
rect 5370 4377 5372 4378
rect 5408 4377 5410 4378
rect 5370 4017 5371 4377
rect 5409 4017 5410 4377
rect 5370 4016 5372 4017
rect 5408 4016 5410 4017
rect 5878 576 6182 577
rect 5878 575 5879 576
rect 6181 575 6182 576
rect 5878 538 5879 539
rect 6181 538 6182 539
rect 5878 537 6182 538
rect 25210 460 25414 461
rect 25210 459 25211 460
rect 25413 459 25414 460
rect 25210 422 25211 423
rect 25413 422 25414 423
rect 25210 421 25414 422
<< via1 >>
rect 25064 469 25070 482
rect 25070 469 25104 482
rect 25104 469 25180 482
rect 25064 435 25142 469
rect 25142 435 25176 469
rect 25176 435 25180 469
rect 25064 430 25180 435
rect 25064 396 25070 430
rect 25070 396 25104 430
rect 25104 396 25180 430
rect 25064 366 25142 396
rect 25142 366 25176 396
rect 25176 366 25180 396
rect 25787 477 25792 482
rect 25792 477 25826 482
rect 25826 477 25864 482
rect 25864 477 25898 482
rect 25898 477 25903 482
rect 25787 438 25903 477
rect 25787 404 25792 438
rect 25792 404 25826 438
rect 25826 404 25864 438
rect 25864 404 25898 438
rect 25898 404 25903 438
rect 25787 366 25903 404
rect 25222 3 25402 119
rect 24181 -4169 24297 -4053
rect 22243 -4316 22359 -4200
<< metal2 >>
rect 25064 482 25903 490
rect 25180 366 25787 482
rect 25064 350 25903 366
rect 3181 -544 3949 322
rect 25210 3 25222 119
rect 25402 3 25414 119
tri 24903 -4053 25210 -3746 se
rect 25210 -3963 25414 3
rect 25210 -4053 25324 -3963
tri 25324 -4053 25414 -3963 nw
rect 24175 -4169 24181 -4053
rect 24297 -4169 25208 -4053
tri 25208 -4169 25324 -4053 nw
rect 22237 -4316 22243 -4200
rect 22359 -4316 22365 -4200
tri 22055 -7795 22237 -7613 se
rect 22237 -7667 22365 -4316
tri 22237 -7795 22365 -7667 nw
tri 21873 -7977 22055 -7795 se
tri 22055 -7977 22237 -7795 nw
tri 21691 -8159 21873 -7977 se
tri 21873 -8159 22055 -7977 nw
tri 21509 -8341 21691 -8159 se
tri 21691 -8341 21873 -8159 nw
tri 21472 -8378 21509 -8341 se
rect 21509 -8378 21654 -8341
tri 21654 -8378 21691 -8341 nw
rect 21472 -8685 21600 -8378
tri 21600 -8432 21654 -8378 nw
rect 21328 -8771 21444 -8685
<< metal3 >>
rect 17294 -11416 21619 -10860
<< metal4 >>
rect 12937 -10864 13477 -10631
tri 13477 -10864 13710 -10631 sw
rect 12937 -11416 17920 -10864
rect 12937 -11649 13477 -11416
tri 13477 -11649 13710 -11416 nw
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 1 0 4780 0 1 3836
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 1 0 1906 0 1 2386
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 2134 1 0 3487
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 497 1 0 417
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 1 0 4893 0 1 3586
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1707688321
transform 1 0 677 0 1 168
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_1
timestamp 1707688321
transform 1 0 5709 0 1 3836
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 1 0 1671 0 1 3746
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 1 0 596 0 1 5346
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform 0 1 894 1 0 2596
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1707688321
transform 0 1 981 1 0 2908
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1707688321
transform 0 1 981 1 0 1972
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1707688321
transform 0 1 981 1 0 2284
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1707688321
transform 1 0 1243 0 1 3004
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 0 1 463 1 0 3060
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1707688321
transform 0 1 2208 1 0 4031
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_2
timestamp 1707688321
transform 0 1 5278 1 0 4044
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_3
timestamp 1707688321
transform 0 1 2351 1 0 4031
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_4
timestamp 1707688321
transform 0 1 5416 1 0 4044
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 1 0 512 0 -1 5802
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1707688321
transform 1 0 516 0 1 5658
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1707688321
transform 1 0 516 0 1 5502
box 0 0 1 1
use L1M1_CDNS_52468879185301  L1M1_CDNS_52468879185301_0
timestamp 1707688321
transform 1 0 1363 0 1 1844
box -12 -6 118 616
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_0
timestamp 1707688321
transform 0 1 1075 -1 0 3520
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_1
timestamp 1707688321
transform 0 1 1075 -1 0 3942
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_2
timestamp 1707688321
transform 0 1 555 -1 0 3520
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_3
timestamp 1707688321
transform 0 1 555 -1 0 3942
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_4
timestamp 1707688321
transform 0 1 757 -1 0 3226
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_5
timestamp 1707688321
transform 0 -1 1434 1 0 1550
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_6
timestamp 1707688321
transform 1 0 1243 0 1 1867
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 1 0 356 0 -1 6114
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1707688321
transform 1 0 356 0 -1 5958
box 0 0 1 1
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1707688321
transform 0 -1 205 1 0 5403
box -12 -6 694 40
use L1M1_CDNS_52468879185948  L1M1_CDNS_52468879185948_0
timestamp 1707688321
transform 1 0 2811 0 1 3942
box -12 -6 1702 40
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_0
timestamp 1707688321
transform 0 1 560 -1 0 3384
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_1
timestamp 1707688321
transform 0 1 560 -1 0 3676
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_2
timestamp 1707688321
transform 0 1 560 -1 0 3786
box -12 -6 46 904
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_0
timestamp 1707688321
transform 0 -1 1464 -1 0 4098
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_1
timestamp 1707688321
transform 0 1 604 1 0 770
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_2
timestamp 1707688321
transform 0 1 604 1 0 458
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_3
timestamp 1707688321
transform 0 1 604 1 0 1706
box -12 -6 46 832
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1707688321
transform 0 1 604 -1 0 3098
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_1
timestamp 1707688321
transform 0 1 604 -1 0 2162
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_2
timestamp 1707688321
transform 0 1 604 -1 0 2786
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_3
timestamp 1707688321
transform 0 1 604 -1 0 2474
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_4
timestamp 1707688321
transform 0 1 604 1 0 1082
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_5
timestamp 1707688321
transform 0 1 604 1 0 1394
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_6
timestamp 1707688321
transform 0 1 1235 1 0 1082
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_7
timestamp 1707688321
transform 0 1 1235 1 0 1394
box 0 0 1 1
use L1M1_CDNS_524688791851067  L1M1_CDNS_524688791851067_0
timestamp 1707688321
transform 0 1 2250 1 0 3586
box -12 -6 46 2056
use L1M1_CDNS_524688791851067  L1M1_CDNS_524688791851067_1
timestamp 1707688321
transform 0 1 2310 1 0 3165
box -12 -6 46 2056
use L1M1_CDNS_524688791851067  L1M1_CDNS_524688791851067_2
timestamp 1707688321
transform 0 1 2265 1 0 3430
box -12 -6 46 2056
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_0
timestamp 1707688321
transform 0 1 5504 1 0 770
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_1
timestamp 1707688321
transform 0 1 5504 1 0 1082
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_2
timestamp 1707688321
transform 0 1 5504 1 0 2018
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_3
timestamp 1707688321
transform 0 1 5504 1 0 1706
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_4
timestamp 1707688321
transform 0 1 5504 1 0 1394
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_5
timestamp 1707688321
transform 0 1 5504 1 0 2330
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_6
timestamp 1707688321
transform 0 1 5504 1 0 3586
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_7
timestamp 1707688321
transform 0 -1 5456 1 0 926
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_8
timestamp 1707688321
transform 0 -1 5456 1 0 614
box 0 0 1 1
use L1M1_CDNS_524688791851562  L1M1_CDNS_524688791851562_0
timestamp 1707688321
transform 0 -1 6383 1 0 4530
box -12 -6 262 112
use L1M1_CDNS_524688791851563  L1M1_CDNS_524688791851563_0
timestamp 1707688321
transform 0 -1 4071 -1 0 4861
box -12 -6 334 184
use L1M1_CDNS_524688791851563  L1M1_CDNS_524688791851563_1
timestamp 1707688321
transform 0 1 3897 1 0 4031
box -12 -6 334 184
use L1M1_CDNS_524688791851563  L1M1_CDNS_524688791851563_2
timestamp 1707688321
transform 0 1 2174 1 0 4527
box -12 -6 334 184
use L1M1_CDNS_524688791851563  L1M1_CDNS_524688791851563_3
timestamp 1707688321
transform 0 1 2837 1 0 4527
box -12 -6 334 184
use L1M1_CDNS_524688791851563  L1M1_CDNS_524688791851563_4
timestamp 1707688321
transform 0 -1 5238 1 0 4527
box -12 -6 334 184
use L1M1_CDNS_524688791851564  L1M1_CDNS_524688791851564_0
timestamp 1707688321
transform 0 1 604 -1 0 1850
box -12 -6 46 544
use L1M1_CDNS_524688791851564  L1M1_CDNS_524688791851564_1
timestamp 1707688321
transform 0 1 896 1 0 926
box -12 -6 46 544
use L1M1_CDNS_524688791851564  L1M1_CDNS_524688791851564_2
timestamp 1707688321
transform 0 1 896 1 0 614
box -12 -6 46 544
use L1M1_CDNS_524688791851564  L1M1_CDNS_524688791851564_3
timestamp 1707688321
transform 0 1 896 1 0 1238
box -12 -6 46 544
use L1M1_CDNS_524688791851565  L1M1_CDNS_524688791851565_0
timestamp 1707688321
transform 0 1 2251 1 0 770
box -12 -6 46 2704
use L1M1_CDNS_524688791851565  L1M1_CDNS_524688791851565_1
timestamp 1707688321
transform 0 1 2285 1 0 1394
box -12 -6 46 2704
use L1M1_CDNS_524688791851565  L1M1_CDNS_524688791851565_2
timestamp 1707688321
transform 0 1 2285 1 0 2018
box -12 -6 46 2704
use L1M1_CDNS_524688791851565  L1M1_CDNS_524688791851565_3
timestamp 1707688321
transform 0 1 2285 1 0 2330
box -12 -6 46 2704
use L1M1_CDNS_524688791851565  L1M1_CDNS_524688791851565_4
timestamp 1707688321
transform 0 1 2285 1 0 1706
box -12 -6 46 2704
use L1M1_CDNS_524688791851566  L1M1_CDNS_524688791851566_0
timestamp 1707688321
transform 0 1 2286 1 0 458
box -12 -6 46 3496
use L1M1_CDNS_524688791851567  L1M1_CDNS_524688791851567_0
timestamp 1707688321
transform 0 1 2246 1 0 614
box -12 -6 46 2488
use L1M1_CDNS_524688791851567  L1M1_CDNS_524688791851567_1
timestamp 1707688321
transform 0 1 2246 1 0 926
box -12 -6 46 2488
use L1M1_CDNS_524688791851568  L1M1_CDNS_524688791851568_0
timestamp 1707688321
transform 1 0 1644 0 1 1846
box -12 -6 406 328
use L1M1_CDNS_524688791851569  L1M1_CDNS_524688791851569_0
timestamp 1707688321
transform 1 0 2250 0 1 5066
box -12 -6 1198 760
use L1M1_CDNS_524688791851570  L1M1_CDNS_524688791851570_0
timestamp 1707688321
transform 0 1 5350 1 0 4527
box -12 -6 334 112
use L1M1_CDNS_524688791851570  L1M1_CDNS_524688791851570_1
timestamp 1707688321
transform 0 -1 6383 1 0 4035
box -12 -6 334 112
use L1M1_CDNS_524688791851571  L1M1_CDNS_524688791851571_0
timestamp 1707688321
transform 0 1 2246 1 0 1238
box -12 -6 46 2992
use L1M1_CDNS_524688791851571  L1M1_CDNS_524688791851571_1
timestamp 1707688321
transform 0 1 2246 1 0 1550
box -12 -6 46 2992
use L1M1_CDNS_524688791851572  L1M1_CDNS_524688791851572_0
timestamp 1707688321
transform 0 1 2286 1 0 1082
box -12 -6 46 2848
use L1M1_CDNS_524688791851573  L1M1_CDNS_524688791851573_0
timestamp 1707688321
transform 1 0 2328 0 1 5858
box -12 -6 1486 112
use L1M1_CDNS_524688791851574  L1M1_CDNS_524688791851574_0
timestamp 1707688321
transform 1 0 3474 0 1 5066
box -12 -6 334 760
use L1M1_CDNS_524688791851575  L1M1_CDNS_524688791851575_0
timestamp 1707688321
transform 0 1 2256 1 0 3009
box -12 -6 46 2200
use L1M1_CDNS_524688791851575  L1M1_CDNS_524688791851575_1
timestamp 1707688321
transform 0 1 2256 1 0 3321
box -12 -6 46 2200
use L1M1_CDNS_524688791851575  L1M1_CDNS_524688791851575_2
timestamp 1707688321
transform 0 1 2242 1 0 2742
box -12 -6 46 2200
use L1M1_CDNS_524688791851576  L1M1_CDNS_524688791851576_0
timestamp 1707688321
transform 0 1 2255 1 0 2898
box -12 -6 46 2416
use L1M1_CDNS_524688791851577  L1M1_CDNS_524688791851577_0
timestamp 1707688321
transform 0 1 2255 1 0 2586
box -12 -6 46 2344
use L1M1_CDNS_524688791851578  L1M1_CDNS_524688791851578_0
timestamp 1707688321
transform 0 1 2250 1 0 3703
box -12 -6 46 2128
use L1M1_CDNS_524688791851579  L1M1_CDNS_524688791851579_0
timestamp 1707688321
transform 0 1 5902 1 0 4899
box -12 -6 478 184
use L1M1_CDNS_524688791851579  L1M1_CDNS_524688791851579_1
timestamp 1707688321
transform 0 -1 4726 1 0 4899
box -12 -6 478 184
use L1M1_CDNS_524688791851580  L1M1_CDNS_524688791851580_0
timestamp 1707688321
transform 0 -1 5238 1 0 1862
box -12 -6 46 2920
use L1M1_CDNS_524688791851580  L1M1_CDNS_524688791851580_1
timestamp 1707688321
transform 0 -1 5238 1 0 2174
box -12 -6 46 2920
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 1 0 25216 0 1 3
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 25787 1 0 360
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform 0 1 25064 1 0 360
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 1 0 22237 0 -1 -4200
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 24175 0 1 -4169
box 0 0 1 1
use M1M2_CDNS_524688791851187  M1M2_CDNS_524688791851187_0
timestamp 1707688321
transform 1 0 3181 0 1 -544
box 0 0 768 180
use M1M2_CDNS_524688791851498  M1M2_CDNS_524688791851498_0
timestamp 1707688321
transform 1 0 3181 0 1 270
box 0 0 768 52
use M3M4_CDNS_524688791851561  M3M4_CDNS_524688791851561_0
timestamp 1707688321
transform 1 0 17295 0 1 -11416
box -1 0 625 556
use nfet_CDNS_524688791851604  nfet_CDNS_524688791851604_0
timestamp 1707688321
transform 0 1 247 -1 0 6069
box -79 -26 335 626
use nfet_CDNS_524688791851604  nfet_CDNS_524688791851604_1
timestamp 1707688321
transform 0 1 247 -1 0 5647
box -79 -26 335 626
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_0
timestamp 1707688321
transform 0 -1 6183 -1 0 2319
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_1
timestamp 1707688321
transform 0 -1 6183 -1 0 2887
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_2
timestamp 1707688321
transform 0 -1 6183 -1 0 3731
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_3
timestamp 1707688321
transform 0 -1 6183 -1 0 3309
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_4
timestamp 1707688321
transform 0 -1 6183 -1 0 2007
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_5
timestamp 1707688321
transform 0 -1 6183 -1 0 1695
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_6
timestamp 1707688321
transform 0 -1 6183 -1 0 1383
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_7
timestamp 1707688321
transform 0 -1 6183 -1 0 1071
box -119 -66 375 4066
use pfet_CDNS_524688791851598  pfet_CDNS_524688791851598_8
timestamp 1707688321
transform 0 -1 6183 -1 0 759
box -119 -66 375 4066
use pfet_CDNS_524688791851601  pfet_CDNS_524688791851601_0
timestamp 1707688321
transform 0 -1 1487 -1 0 1695
box -119 -66 1311 1066
use pfet_CDNS_524688791851602  pfet_CDNS_524688791851602_0
timestamp 1707688321
transform 0 -1 1195 -1 0 3209
box -119 -66 1467 666
use pfet_CDNS_524688791851603  pfet_CDNS_524688791851603_0
timestamp 1707688321
transform 0 -1 1487 -1 0 4053
box -119 -66 375 1066
use pfet_CDNS_524688791851603  pfet_CDNS_524688791851603_1
timestamp 1707688321
transform 0 -1 1487 -1 0 3631
box -119 -66 375 1066
use PYres_CDNS_524688791851597  PYres_CDNS_524688791851597_0
timestamp 1707688321
transform -1 0 3993 0 1 4000
box -50 0 2132 400
use PYres_CDNS_524688791851597  PYres_CDNS_524688791851597_1
timestamp 1707688321
transform -1 0 6311 0 1 4000
box -50 0 2132 400
use PYres_CDNS_524688791851597  PYres_CDNS_524688791851597_2
timestamp 1707688321
transform 1 0 4233 0 1 4496
box -50 0 2132 400
use PYres_CDNS_524688791851597  PYres_CDNS_524688791851597_3
timestamp 1707688321
transform 1 0 1911 0 1 4496
box -50 0 2132 400
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1707688321
transform -1 0 6375 0 1 4990
box 0 0 2270 404
use sky130_fd_io__sio_pudrvr_reg_pu_natives  sky130_fd_io__sio_pudrvr_reg_pu_natives_0
timestamp 1707688321
transform 1 0 6455 0 1 -12115
box -184 0 18805 17853
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1707688321
transform 1 0 1026 0 1 2584
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851581  sky130_fd_io__tk_em1o_CDNS_524688791851581_0
timestamp 1707688321
transform 0 1 888 -1 0 2470
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851582  sky130_fd_io__tk_em1s_CDNS_524688791851582_0
timestamp 1707688321
transform 0 -1 6182 1 0 485
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851583  sky130_fd_io__tk_em1s_CDNS_524688791851583_0
timestamp 1707688321
transform 0 -1 25414 1 0 369
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851584  sky130_fd_io__tk_em1s_CDNS_524688791851584_0
timestamp 1707688321
transform -1 0 2889 0 1 4515
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851584  sky130_fd_io__tk_em1s_CDNS_524688791851584_1
timestamp 1707688321
transform -1 0 2393 0 1 4019
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851585  sky130_fd_io__tk_em1s_CDNS_524688791851585_0
timestamp 1707688321
transform -1 0 5462 0 1 4016
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851585  sky130_fd_io__tk_em1s_CDNS_524688791851585_1
timestamp 1707688321
transform -1 0 5388 0 1 4515
box 0 0 1 1
<< labels >>
flabel comment s 7700 4757 7700 4757 0 FreeSans 1000 0 0 0 condiode
flabel comment s 17539 -8656 17539 -8656 0 FreeSans 1000 0 0 0 condiode
flabel comment s 3747 5044 3747 5044 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 6536 5559 6536 5559 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 6541 3512 6541 3512 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 25475 686 25475 686 0 FreeSans 300 90 0 0 pug<0>
flabel comment s 13116 6967 13116 6967 0 FreeSans 1600 0 0 0 top cell boundary
flabel comment s 5151 4708 5151 4708 0 FreeSans 1000 0 0 0 I80
flabel comment s 25557 635 25557 635 0 FreeSans 300 90 0 0 pu_h_n<0>
flabel comment s 25637 641 25637 641 0 FreeSans 300 90 0 0 pu_h_n<1>
flabel comment s 2342 4611 2342 4611 0 FreeSans 1000 0 0 0 I79
flabel comment s 1026 1651 1026 1651 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 1492 1026 1492 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 1332 1026 1332 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 1180 1026 1180 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 555 1026 555 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 707 1026 707 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 866 1026 866 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 1026 1028 1026 1028 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 4769 1028 4769 1028 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 4769 865 4769 865 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 4769 715 4769 715 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 4769 560 4769 560 0 FreeSans 200 0 0 0 pdrvr0
flabel comment s 2142 4107 2142 4107 0 FreeSans 1000 0 0 0 I81
flabel comment s 5136 5094 5136 5094 0 FreeSans 1000 0 0 0 resd
flabel comment s 5172 4198 5172 4198 0 FreeSans 1000 0 0 0 I78
flabel comment s 611 132 611 132 0 FreeSans 200 90 0 0 nghs_h
flabel comment s 25039 6324 25039 6324 0 FreeSans 300 0 0 0 pug<1>
flabel comment s 25034 6074 25034 6074 0 FreeSans 300 0 0 0 pug<0>
flabel comment s 24989 6236 24989 6236 0 FreeSans 300 0 0 0 pu_h_n<1>
flabel comment s 24983 6156 24983 6156 0 FreeSans 300 0 0 0 pu_h_n<0>
flabel comment s 692 131 692 131 0 FreeSans 200 90 0 0 pghs_h
flabel comment s 2034 5394 2034 5394 0 FreeSans 300 90 0 0 pu_h_n<0>
flabel comment s 1921 5400 1921 5400 0 FreeSans 300 90 0 0 pu_h_n<1>
flabel comment s 2110 5445 2110 5445 0 FreeSans 300 90 0 0 pug<0>
flabel comment s 1833 5450 1833 5450 0 FreeSans 300 90 0 0 pug<1>
flabel comment s 25725 691 25725 691 0 FreeSans 300 90 0 0 pug<1>
flabel metal1 s 16995 -8910 17113 -8838 3 FreeSans 200 90 0 0 vgnd_io
port 2 nsew
flabel metal1 s 16298 170 17044 224 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal1 s 10938 170 11684 224 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal1 s 12176 170 12922 224 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal1 s 16643 -8556 16771 -8437 3 FreeSans 200 90 0 0 vcc_io
port 4 nsew
flabel metal1 s 6482 322 6674 355 3 FreeSans 200 180 0 0 vpb_drvr
port 5 nsew
flabel metal1 s 5878 142 6246 238 0 FreeSans 200 0 0 0 pad
port 3 nsew
flabel metal1 s 8053 170 8799 224 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal1 s 6815 142 7562 196 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal1 s 71 114 189 193 3 FreeSans 200 90 0 0 vnb
port 6 nsew
flabel metal1 s -309 134 -191 146 3 FreeSans 200 90 0 0 vcc_io
port 4 nsew
flabel metal1 s 5658 366 5850 378 3 FreeSans 200 90 0 0 vcc_io
port 4 nsew
flabel metal1 s 665 114 717 149 0 FreeSans 200 90 0 0 pghs_h
port 7 nsew
flabel metal1 s 585 114 637 149 0 FreeSans 200 90 0 0 nghs_h
port 8 nsew
flabel metal4 s 12970 -11617 13469 -10669 3 FreeSans 200 90 0 0 pad
port 3 nsew
flabel metal2 s 3181 -544 3949 -364 3 FreeSans 200 90 0 0 vpb_drvr
port 5 nsew
flabel metal2 s 21328 -8771 21444 -8685 7 FreeSans 200 90 0 0 vref_nng
port 9 nsew
<< properties >>
string GDS_END 96445916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95663210
string path 9.600 7.600 9.600 106.300 
<< end >>
