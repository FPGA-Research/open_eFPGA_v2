magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< locali >>
rect 5664 50491 5680 50525
rect 5714 50491 5730 50525
rect 7031 50425 7484 50459
rect 5554 50379 5570 50413
rect 5604 50379 5620 50413
rect 5664 50289 5680 50323
rect 5714 50289 5730 50323
rect 5664 50065 5680 50099
rect 5714 50065 5730 50099
rect 5554 49975 5570 50009
rect 5604 49975 5620 50009
rect 7031 49929 7484 49963
rect 5664 49863 5680 49897
rect 5714 49863 5730 49897
rect 5664 49701 5680 49735
rect 5714 49701 5730 49735
rect 7031 49635 7484 49669
rect 5554 49589 5570 49623
rect 5604 49589 5620 49623
rect 5664 49499 5680 49533
rect 5714 49499 5730 49533
rect 5664 49275 5680 49309
rect 5714 49275 5730 49309
rect 5554 49185 5570 49219
rect 5604 49185 5620 49219
rect 7031 49139 7484 49173
rect 5664 49073 5680 49107
rect 5714 49073 5730 49107
rect 5664 48911 5680 48945
rect 5714 48911 5730 48945
rect 7031 48845 7484 48879
rect 5554 48799 5570 48833
rect 5604 48799 5620 48833
rect 5664 48709 5680 48743
rect 5714 48709 5730 48743
rect 5664 48485 5680 48519
rect 5714 48485 5730 48519
rect 5554 48395 5570 48429
rect 5604 48395 5620 48429
rect 7031 48349 7484 48383
rect 5664 48283 5680 48317
rect 5714 48283 5730 48317
rect 5664 48121 5680 48155
rect 5714 48121 5730 48155
rect 7031 48055 7484 48089
rect 5554 48009 5570 48043
rect 5604 48009 5620 48043
rect 5664 47919 5680 47953
rect 5714 47919 5730 47953
rect 5664 47695 5680 47729
rect 5714 47695 5730 47729
rect 5554 47605 5570 47639
rect 5604 47605 5620 47639
rect 7031 47559 7484 47593
rect 5664 47493 5680 47527
rect 5714 47493 5730 47527
rect 5664 47331 5680 47365
rect 5714 47331 5730 47365
rect 7031 47265 7484 47299
rect 5554 47219 5570 47253
rect 5604 47219 5620 47253
rect 5664 47129 5680 47163
rect 5714 47129 5730 47163
rect 5664 46905 5680 46939
rect 5714 46905 5730 46939
rect 5554 46815 5570 46849
rect 5604 46815 5620 46849
rect 7031 46769 7484 46803
rect 5664 46703 5680 46737
rect 5714 46703 5730 46737
rect 5664 46541 5680 46575
rect 5714 46541 5730 46575
rect 7031 46475 7484 46509
rect 5554 46429 5570 46463
rect 5604 46429 5620 46463
rect 5664 46339 5680 46373
rect 5714 46339 5730 46373
rect 5664 46115 5680 46149
rect 5714 46115 5730 46149
rect 5554 46025 5570 46059
rect 5604 46025 5620 46059
rect 7031 45979 7484 46013
rect 5664 45913 5680 45947
rect 5714 45913 5730 45947
rect 5664 45751 5680 45785
rect 5714 45751 5730 45785
rect 7031 45685 7484 45719
rect 5554 45639 5570 45673
rect 5604 45639 5620 45673
rect 5664 45549 5680 45583
rect 5714 45549 5730 45583
rect 5664 45325 5680 45359
rect 5714 45325 5730 45359
rect 5554 45235 5570 45269
rect 5604 45235 5620 45269
rect 7031 45189 7484 45223
rect 5664 45123 5680 45157
rect 5714 45123 5730 45157
rect 5664 44961 5680 44995
rect 5714 44961 5730 44995
rect 7031 44895 7484 44929
rect 5554 44849 5570 44883
rect 5604 44849 5620 44883
rect 5664 44759 5680 44793
rect 5714 44759 5730 44793
rect 5664 44535 5680 44569
rect 5714 44535 5730 44569
rect 5554 44445 5570 44479
rect 5604 44445 5620 44479
rect 7031 44399 7484 44433
rect 5664 44333 5680 44367
rect 5714 44333 5730 44367
rect 5664 44171 5680 44205
rect 5714 44171 5730 44205
rect 7031 44105 7484 44139
rect 5554 44059 5570 44093
rect 5604 44059 5620 44093
rect 5664 43969 5680 44003
rect 5714 43969 5730 44003
rect 5664 43745 5680 43779
rect 5714 43745 5730 43779
rect 5554 43655 5570 43689
rect 5604 43655 5620 43689
rect 7031 43609 7484 43643
rect 5664 43543 5680 43577
rect 5714 43543 5730 43577
rect 5664 43381 5680 43415
rect 5714 43381 5730 43415
rect 7031 43315 7484 43349
rect 5554 43269 5570 43303
rect 5604 43269 5620 43303
rect 5664 43179 5680 43213
rect 5714 43179 5730 43213
rect 5664 42955 5680 42989
rect 5714 42955 5730 42989
rect 5554 42865 5570 42899
rect 5604 42865 5620 42899
rect 7031 42819 7484 42853
rect 5664 42753 5680 42787
rect 5714 42753 5730 42787
rect 5664 42591 5680 42625
rect 5714 42591 5730 42625
rect 7031 42525 7484 42559
rect 5554 42479 5570 42513
rect 5604 42479 5620 42513
rect 5664 42389 5680 42423
rect 5714 42389 5730 42423
rect 5664 42165 5680 42199
rect 5714 42165 5730 42199
rect 5554 42075 5570 42109
rect 5604 42075 5620 42109
rect 7031 42029 7484 42063
rect 5664 41963 5680 41997
rect 5714 41963 5730 41997
rect 5664 41801 5680 41835
rect 5714 41801 5730 41835
rect 7031 41735 7484 41769
rect 5554 41689 5570 41723
rect 5604 41689 5620 41723
rect 5664 41599 5680 41633
rect 5714 41599 5730 41633
rect 5664 41375 5680 41409
rect 5714 41375 5730 41409
rect 5554 41285 5570 41319
rect 5604 41285 5620 41319
rect 7031 41239 7484 41273
rect 5664 41173 5680 41207
rect 5714 41173 5730 41207
rect 5664 41011 5680 41045
rect 5714 41011 5730 41045
rect 7031 40945 7484 40979
rect 5554 40899 5570 40933
rect 5604 40899 5620 40933
rect 5664 40809 5680 40843
rect 5714 40809 5730 40843
rect 5664 40585 5680 40619
rect 5714 40585 5730 40619
rect 5554 40495 5570 40529
rect 5604 40495 5620 40529
rect 7031 40449 7484 40483
rect 5664 40383 5680 40417
rect 5714 40383 5730 40417
rect 5664 40221 5680 40255
rect 5714 40221 5730 40255
rect 7031 40155 7484 40189
rect 5554 40109 5570 40143
rect 5604 40109 5620 40143
rect 5664 40019 5680 40053
rect 5714 40019 5730 40053
rect 5664 39795 5680 39829
rect 5714 39795 5730 39829
rect 5554 39705 5570 39739
rect 5604 39705 5620 39739
rect 7031 39659 7484 39693
rect 5664 39593 5680 39627
rect 5714 39593 5730 39627
rect 5664 39431 5680 39465
rect 5714 39431 5730 39465
rect 7031 39365 7484 39399
rect 5554 39319 5570 39353
rect 5604 39319 5620 39353
rect 5664 39229 5680 39263
rect 5714 39229 5730 39263
rect 5664 39005 5680 39039
rect 5714 39005 5730 39039
rect 5554 38915 5570 38949
rect 5604 38915 5620 38949
rect 7031 38869 7484 38903
rect 5664 38803 5680 38837
rect 5714 38803 5730 38837
rect 5664 38641 5680 38675
rect 5714 38641 5730 38675
rect 7031 38575 7484 38609
rect 5554 38529 5570 38563
rect 5604 38529 5620 38563
rect 5664 38439 5680 38473
rect 5714 38439 5730 38473
rect 5664 38215 5680 38249
rect 5714 38215 5730 38249
rect 5554 38125 5570 38159
rect 5604 38125 5620 38159
rect 7031 38079 7484 38113
rect 5664 38013 5680 38047
rect 5714 38013 5730 38047
rect 5664 37851 5680 37885
rect 5714 37851 5730 37885
rect 7031 37785 7484 37819
rect 5554 37739 5570 37773
rect 5604 37739 5620 37773
rect 5664 37649 5680 37683
rect 5714 37649 5730 37683
rect 5664 37425 5680 37459
rect 5714 37425 5730 37459
rect 5554 37335 5570 37369
rect 5604 37335 5620 37369
rect 7031 37289 7484 37323
rect 5664 37223 5680 37257
rect 5714 37223 5730 37257
rect 5664 37061 5680 37095
rect 5714 37061 5730 37095
rect 7031 36995 7484 37029
rect 5554 36949 5570 36983
rect 5604 36949 5620 36983
rect 5664 36859 5680 36893
rect 5714 36859 5730 36893
rect 5664 36635 5680 36669
rect 5714 36635 5730 36669
rect 5554 36545 5570 36579
rect 5604 36545 5620 36579
rect 7031 36499 7484 36533
rect 5664 36433 5680 36467
rect 5714 36433 5730 36467
rect 5664 36271 5680 36305
rect 5714 36271 5730 36305
rect 7031 36205 7484 36239
rect 5554 36159 5570 36193
rect 5604 36159 5620 36193
rect 5664 36069 5680 36103
rect 5714 36069 5730 36103
rect 5664 35845 5680 35879
rect 5714 35845 5730 35879
rect 5554 35755 5570 35789
rect 5604 35755 5620 35789
rect 7031 35709 7484 35743
rect 5664 35643 5680 35677
rect 5714 35643 5730 35677
rect 5664 35481 5680 35515
rect 5714 35481 5730 35515
rect 7031 35415 7484 35449
rect 5554 35369 5570 35403
rect 5604 35369 5620 35403
rect 5664 35279 5680 35313
rect 5714 35279 5730 35313
rect 5664 35055 5680 35089
rect 5714 35055 5730 35089
rect 5554 34965 5570 34999
rect 5604 34965 5620 34999
rect 7031 34919 7484 34953
rect 5664 34853 5680 34887
rect 5714 34853 5730 34887
rect 5664 34691 5680 34725
rect 5714 34691 5730 34725
rect 7031 34625 7484 34659
rect 5554 34579 5570 34613
rect 5604 34579 5620 34613
rect 5664 34489 5680 34523
rect 5714 34489 5730 34523
rect 5664 34265 5680 34299
rect 5714 34265 5730 34299
rect 5554 34175 5570 34209
rect 5604 34175 5620 34209
rect 7031 34129 7484 34163
rect 5664 34063 5680 34097
rect 5714 34063 5730 34097
rect 5664 33901 5680 33935
rect 5714 33901 5730 33935
rect 7031 33835 7484 33869
rect 5554 33789 5570 33823
rect 5604 33789 5620 33823
rect 5664 33699 5680 33733
rect 5714 33699 5730 33733
rect 5664 33475 5680 33509
rect 5714 33475 5730 33509
rect 5554 33385 5570 33419
rect 5604 33385 5620 33419
rect 7031 33339 7484 33373
rect 5664 33273 5680 33307
rect 5714 33273 5730 33307
rect 5664 33111 5680 33145
rect 5714 33111 5730 33145
rect 7031 33045 7484 33079
rect 5554 32999 5570 33033
rect 5604 32999 5620 33033
rect 5664 32909 5680 32943
rect 5714 32909 5730 32943
rect 5664 32685 5680 32719
rect 5714 32685 5730 32719
rect 5554 32595 5570 32629
rect 5604 32595 5620 32629
rect 7031 32549 7484 32583
rect 5664 32483 5680 32517
rect 5714 32483 5730 32517
rect 5664 32321 5680 32355
rect 5714 32321 5730 32355
rect 7031 32255 7484 32289
rect 5554 32209 5570 32243
rect 5604 32209 5620 32243
rect 5664 32119 5680 32153
rect 5714 32119 5730 32153
rect 5664 31895 5680 31929
rect 5714 31895 5730 31929
rect 5554 31805 5570 31839
rect 5604 31805 5620 31839
rect 7031 31759 7484 31793
rect 5664 31693 5680 31727
rect 5714 31693 5730 31727
rect 5664 31531 5680 31565
rect 5714 31531 5730 31565
rect 7031 31465 7484 31499
rect 5554 31419 5570 31453
rect 5604 31419 5620 31453
rect 5664 31329 5680 31363
rect 5714 31329 5730 31363
rect 5664 31105 5680 31139
rect 5714 31105 5730 31139
rect 5554 31015 5570 31049
rect 5604 31015 5620 31049
rect 7031 30969 7484 31003
rect 5664 30903 5680 30937
rect 5714 30903 5730 30937
rect 5664 30741 5680 30775
rect 5714 30741 5730 30775
rect 7031 30675 7484 30709
rect 5554 30629 5570 30663
rect 5604 30629 5620 30663
rect 5664 30539 5680 30573
rect 5714 30539 5730 30573
rect 5664 30315 5680 30349
rect 5714 30315 5730 30349
rect 5554 30225 5570 30259
rect 5604 30225 5620 30259
rect 7031 30179 7484 30213
rect 5664 30113 5680 30147
rect 5714 30113 5730 30147
rect 5664 29951 5680 29985
rect 5714 29951 5730 29985
rect 7031 29885 7484 29919
rect 5554 29839 5570 29873
rect 5604 29839 5620 29873
rect 5664 29749 5680 29783
rect 5714 29749 5730 29783
rect 5664 29525 5680 29559
rect 5714 29525 5730 29559
rect 5554 29435 5570 29469
rect 5604 29435 5620 29469
rect 7031 29389 7484 29423
rect 5664 29323 5680 29357
rect 5714 29323 5730 29357
rect 5664 29161 5680 29195
rect 5714 29161 5730 29195
rect 7031 29095 7484 29129
rect 5554 29049 5570 29083
rect 5604 29049 5620 29083
rect 5664 28959 5680 28993
rect 5714 28959 5730 28993
rect 5664 28735 5680 28769
rect 5714 28735 5730 28769
rect 5554 28645 5570 28679
rect 5604 28645 5620 28679
rect 7031 28599 7484 28633
rect 5664 28533 5680 28567
rect 5714 28533 5730 28567
rect 5664 28371 5680 28405
rect 5714 28371 5730 28405
rect 7031 28305 7484 28339
rect 5554 28259 5570 28293
rect 5604 28259 5620 28293
rect 5664 28169 5680 28203
rect 5714 28169 5730 28203
rect 5664 27945 5680 27979
rect 5714 27945 5730 27979
rect 5554 27855 5570 27889
rect 5604 27855 5620 27889
rect 7031 27809 7484 27843
rect 5664 27743 5680 27777
rect 5714 27743 5730 27777
rect 5664 27581 5680 27615
rect 5714 27581 5730 27615
rect 7031 27515 7484 27549
rect 5554 27469 5570 27503
rect 5604 27469 5620 27503
rect 5664 27379 5680 27413
rect 5714 27379 5730 27413
rect 5664 27155 5680 27189
rect 5714 27155 5730 27189
rect 5554 27065 5570 27099
rect 5604 27065 5620 27099
rect 7031 27019 7484 27053
rect 5664 26953 5680 26987
rect 5714 26953 5730 26987
rect 5664 26791 5680 26825
rect 5714 26791 5730 26825
rect 7031 26725 7484 26759
rect 5554 26679 5570 26713
rect 5604 26679 5620 26713
rect 5664 26589 5680 26623
rect 5714 26589 5730 26623
rect 5664 26365 5680 26399
rect 5714 26365 5730 26399
rect 5554 26275 5570 26309
rect 5604 26275 5620 26309
rect 7031 26229 7484 26263
rect 5664 26163 5680 26197
rect 5714 26163 5730 26197
rect 5664 26001 5680 26035
rect 5714 26001 5730 26035
rect 7031 25935 7484 25969
rect 5554 25889 5570 25923
rect 5604 25889 5620 25923
rect 5664 25799 5680 25833
rect 5714 25799 5730 25833
rect 5664 25575 5680 25609
rect 5714 25575 5730 25609
rect 5554 25485 5570 25519
rect 5604 25485 5620 25519
rect 7031 25439 7484 25473
rect 5664 25373 5680 25407
rect 5714 25373 5730 25407
rect 5664 25211 5680 25245
rect 5714 25211 5730 25245
rect 7031 25145 7484 25179
rect 5554 25099 5570 25133
rect 5604 25099 5620 25133
rect 5664 25009 5680 25043
rect 5714 25009 5730 25043
rect 5664 24785 5680 24819
rect 5714 24785 5730 24819
rect 5554 24695 5570 24729
rect 5604 24695 5620 24729
rect 7031 24649 7484 24683
rect 5664 24583 5680 24617
rect 5714 24583 5730 24617
rect 5664 24421 5680 24455
rect 5714 24421 5730 24455
rect 7031 24355 7484 24389
rect 5554 24309 5570 24343
rect 5604 24309 5620 24343
rect 5664 24219 5680 24253
rect 5714 24219 5730 24253
rect 5664 23995 5680 24029
rect 5714 23995 5730 24029
rect 5554 23905 5570 23939
rect 5604 23905 5620 23939
rect 7031 23859 7484 23893
rect 5664 23793 5680 23827
rect 5714 23793 5730 23827
rect 5664 23631 5680 23665
rect 5714 23631 5730 23665
rect 7031 23565 7484 23599
rect 5554 23519 5570 23553
rect 5604 23519 5620 23553
rect 5664 23429 5680 23463
rect 5714 23429 5730 23463
rect 5664 23205 5680 23239
rect 5714 23205 5730 23239
rect 5554 23115 5570 23149
rect 5604 23115 5620 23149
rect 7031 23069 7484 23103
rect 5664 23003 5680 23037
rect 5714 23003 5730 23037
rect 5664 22841 5680 22875
rect 5714 22841 5730 22875
rect 7031 22775 7484 22809
rect 5554 22729 5570 22763
rect 5604 22729 5620 22763
rect 5664 22639 5680 22673
rect 5714 22639 5730 22673
rect 5664 22415 5680 22449
rect 5714 22415 5730 22449
rect 5554 22325 5570 22359
rect 5604 22325 5620 22359
rect 7031 22279 7484 22313
rect 5664 22213 5680 22247
rect 5714 22213 5730 22247
rect 5664 22051 5680 22085
rect 5714 22051 5730 22085
rect 7031 21985 7484 22019
rect 5554 21939 5570 21973
rect 5604 21939 5620 21973
rect 5664 21849 5680 21883
rect 5714 21849 5730 21883
rect 5664 21625 5680 21659
rect 5714 21625 5730 21659
rect 5554 21535 5570 21569
rect 5604 21535 5620 21569
rect 7031 21489 7484 21523
rect 5664 21423 5680 21457
rect 5714 21423 5730 21457
rect 5664 21261 5680 21295
rect 5714 21261 5730 21295
rect 7031 21195 7484 21229
rect 5554 21149 5570 21183
rect 5604 21149 5620 21183
rect 5664 21059 5680 21093
rect 5714 21059 5730 21093
rect 5664 20835 5680 20869
rect 5714 20835 5730 20869
rect 5554 20745 5570 20779
rect 5604 20745 5620 20779
rect 7031 20699 7484 20733
rect 5664 20633 5680 20667
rect 5714 20633 5730 20667
rect 5664 20471 5680 20505
rect 5714 20471 5730 20505
rect 7031 20405 7484 20439
rect 5554 20359 5570 20393
rect 5604 20359 5620 20393
rect 5664 20269 5680 20303
rect 5714 20269 5730 20303
rect 5664 20045 5680 20079
rect 5714 20045 5730 20079
rect 5554 19955 5570 19989
rect 5604 19955 5620 19989
rect 7031 19909 7484 19943
rect 5664 19843 5680 19877
rect 5714 19843 5730 19877
rect 5664 19681 5680 19715
rect 5714 19681 5730 19715
rect 7031 19615 7484 19649
rect 5554 19569 5570 19603
rect 5604 19569 5620 19603
rect 5664 19479 5680 19513
rect 5714 19479 5730 19513
rect 5664 19255 5680 19289
rect 5714 19255 5730 19289
rect 5554 19165 5570 19199
rect 5604 19165 5620 19199
rect 7031 19119 7484 19153
rect 5664 19053 5680 19087
rect 5714 19053 5730 19087
rect 5664 18891 5680 18925
rect 5714 18891 5730 18925
rect 7031 18825 7484 18859
rect 5554 18779 5570 18813
rect 5604 18779 5620 18813
rect 5664 18689 5680 18723
rect 5714 18689 5730 18723
rect 5664 18465 5680 18499
rect 5714 18465 5730 18499
rect 5554 18375 5570 18409
rect 5604 18375 5620 18409
rect 7031 18329 7484 18363
rect 5664 18263 5680 18297
rect 5714 18263 5730 18297
rect 5664 18101 5680 18135
rect 5714 18101 5730 18135
rect 7031 18035 7484 18069
rect 5554 17989 5570 18023
rect 5604 17989 5620 18023
rect 5664 17899 5680 17933
rect 5714 17899 5730 17933
rect 5664 17675 5680 17709
rect 5714 17675 5730 17709
rect 5554 17585 5570 17619
rect 5604 17585 5620 17619
rect 7031 17539 7484 17573
rect 5664 17473 5680 17507
rect 5714 17473 5730 17507
rect 5664 17311 5680 17345
rect 5714 17311 5730 17345
rect 7031 17245 7484 17279
rect 5554 17199 5570 17233
rect 5604 17199 5620 17233
rect 5664 17109 5680 17143
rect 5714 17109 5730 17143
rect 5664 16885 5680 16919
rect 5714 16885 5730 16919
rect 5554 16795 5570 16829
rect 5604 16795 5620 16829
rect 7031 16749 7484 16783
rect 5664 16683 5680 16717
rect 5714 16683 5730 16717
rect 5664 16521 5680 16555
rect 5714 16521 5730 16555
rect 7031 16455 7484 16489
rect 5554 16409 5570 16443
rect 5604 16409 5620 16443
rect 5664 16319 5680 16353
rect 5714 16319 5730 16353
rect 5664 16095 5680 16129
rect 5714 16095 5730 16129
rect 5554 16005 5570 16039
rect 5604 16005 5620 16039
rect 7031 15959 7484 15993
rect 5664 15893 5680 15927
rect 5714 15893 5730 15927
rect 5664 15731 5680 15765
rect 5714 15731 5730 15765
rect 7031 15665 7484 15699
rect 5554 15619 5570 15653
rect 5604 15619 5620 15653
rect 5664 15529 5680 15563
rect 5714 15529 5730 15563
rect 5664 15305 5680 15339
rect 5714 15305 5730 15339
rect 5554 15215 5570 15249
rect 5604 15215 5620 15249
rect 7031 15169 7484 15203
rect 5664 15103 5680 15137
rect 5714 15103 5730 15137
rect 5664 14941 5680 14975
rect 5714 14941 5730 14975
rect 7031 14875 7484 14909
rect 5554 14829 5570 14863
rect 5604 14829 5620 14863
rect 5664 14739 5680 14773
rect 5714 14739 5730 14773
rect 5664 14515 5680 14549
rect 5714 14515 5730 14549
rect 5554 14425 5570 14459
rect 5604 14425 5620 14459
rect 7031 14379 7484 14413
rect 5664 14313 5680 14347
rect 5714 14313 5730 14347
rect 5664 14151 5680 14185
rect 5714 14151 5730 14185
rect 7031 14085 7484 14119
rect 5554 14039 5570 14073
rect 5604 14039 5620 14073
rect 5664 13949 5680 13983
rect 5714 13949 5730 13983
rect 5664 13725 5680 13759
rect 5714 13725 5730 13759
rect 5554 13635 5570 13669
rect 5604 13635 5620 13669
rect 7031 13589 7484 13623
rect 5664 13523 5680 13557
rect 5714 13523 5730 13557
rect 5664 13361 5680 13395
rect 5714 13361 5730 13395
rect 7031 13295 7484 13329
rect 5554 13249 5570 13283
rect 5604 13249 5620 13283
rect 5664 13159 5680 13193
rect 5714 13159 5730 13193
rect 5664 12935 5680 12969
rect 5714 12935 5730 12969
rect 5554 12845 5570 12879
rect 5604 12845 5620 12879
rect 7031 12799 7484 12833
rect 5664 12733 5680 12767
rect 5714 12733 5730 12767
rect 5664 12571 5680 12605
rect 5714 12571 5730 12605
rect 7031 12505 7484 12539
rect 5554 12459 5570 12493
rect 5604 12459 5620 12493
rect 5664 12369 5680 12403
rect 5714 12369 5730 12403
rect 5664 12145 5680 12179
rect 5714 12145 5730 12179
rect 5554 12055 5570 12089
rect 5604 12055 5620 12089
rect 7031 12009 7484 12043
rect 5664 11943 5680 11977
rect 5714 11943 5730 11977
rect 5664 11781 5680 11815
rect 5714 11781 5730 11815
rect 7031 11715 7484 11749
rect 5554 11669 5570 11703
rect 5604 11669 5620 11703
rect 5664 11579 5680 11613
rect 5714 11579 5730 11613
rect 5664 11355 5680 11389
rect 5714 11355 5730 11389
rect 5554 11265 5570 11299
rect 5604 11265 5620 11299
rect 7031 11219 7484 11253
rect 5664 11153 5680 11187
rect 5714 11153 5730 11187
rect 5664 10991 5680 11025
rect 5714 10991 5730 11025
rect 7031 10925 7484 10959
rect 5554 10879 5570 10913
rect 5604 10879 5620 10913
rect 5664 10789 5680 10823
rect 5714 10789 5730 10823
rect 5664 10565 5680 10599
rect 5714 10565 5730 10599
rect 5554 10475 5570 10509
rect 5604 10475 5620 10509
rect 7031 10429 7484 10463
rect 5664 10363 5680 10397
rect 5714 10363 5730 10397
rect 5664 10201 5680 10235
rect 5714 10201 5730 10235
rect 7031 10135 7484 10169
rect 5554 10089 5570 10123
rect 5604 10089 5620 10123
rect 5664 9999 5680 10033
rect 5714 9999 5730 10033
rect 5664 9775 5680 9809
rect 5714 9775 5730 9809
rect 5554 9685 5570 9719
rect 5604 9685 5620 9719
rect 7031 9639 7484 9673
rect 5664 9573 5680 9607
rect 5714 9573 5730 9607
rect 5664 9411 5680 9445
rect 5714 9411 5730 9445
rect 7031 9345 7484 9379
rect 5554 9299 5570 9333
rect 5604 9299 5620 9333
rect 5664 9209 5680 9243
rect 5714 9209 5730 9243
rect 5664 8985 5680 9019
rect 5714 8985 5730 9019
rect 5554 8895 5570 8929
rect 5604 8895 5620 8929
rect 7031 8849 7484 8883
rect 5664 8783 5680 8817
rect 5714 8783 5730 8817
rect 5664 8621 5680 8655
rect 5714 8621 5730 8655
rect 7031 8555 7484 8589
rect 5554 8509 5570 8543
rect 5604 8509 5620 8543
rect 5664 8419 5680 8453
rect 5714 8419 5730 8453
rect 5664 8195 5680 8229
rect 5714 8195 5730 8229
rect 5554 8105 5570 8139
rect 5604 8105 5620 8139
rect 7031 8059 7484 8093
rect 5664 7993 5680 8027
rect 5714 7993 5730 8027
rect 5664 7831 5680 7865
rect 5714 7831 5730 7865
rect 4177 7765 4279 7799
rect 7031 7765 7484 7799
rect 4245 7551 4279 7765
rect 5554 7719 5570 7753
rect 5604 7719 5620 7753
rect 5664 7629 5680 7663
rect 5714 7629 5730 7663
rect 4245 7517 5471 7551
rect 5505 7517 5521 7551
rect 5664 7405 5680 7439
rect 5714 7405 5730 7439
rect 5554 7315 5570 7349
rect 5604 7315 5620 7349
rect 4177 7269 4279 7303
rect 7031 7269 7484 7303
rect 4245 7156 4279 7269
rect 5664 7203 5680 7237
rect 5714 7203 5730 7237
rect 4245 7122 5391 7156
rect 5425 7122 5441 7156
rect 5664 7041 5680 7075
rect 5714 7041 5730 7075
rect 4177 6975 4279 7009
rect 7031 6975 7484 7009
rect 4245 6761 4279 6975
rect 5554 6929 5570 6963
rect 5604 6929 5620 6963
rect 5664 6839 5680 6873
rect 5714 6839 5730 6873
rect 4245 6727 5311 6761
rect 5345 6727 5361 6761
rect 5664 6615 5680 6649
rect 5714 6615 5730 6649
rect 5554 6525 5570 6559
rect 5604 6525 5620 6559
rect 4177 6479 4279 6513
rect 7031 6479 7484 6513
rect 4245 6366 4279 6479
rect 5664 6413 5680 6447
rect 5714 6413 5730 6447
rect 4245 6332 5231 6366
rect 5265 6332 5281 6366
rect 5664 6251 5680 6285
rect 5714 6251 5730 6285
rect 4177 6185 4279 6219
rect 7031 6185 7484 6219
rect 4245 5971 4279 6185
rect 5554 6139 5570 6173
rect 5604 6139 5620 6173
rect 5664 6049 5680 6083
rect 5714 6049 5730 6083
rect 4245 5937 5151 5971
rect 5185 5937 5201 5971
rect 5664 5825 5680 5859
rect 5714 5825 5730 5859
rect 5554 5735 5570 5769
rect 5604 5735 5620 5769
rect 4177 5689 4279 5723
rect 7031 5689 7484 5723
rect 4245 5576 4279 5689
rect 5664 5623 5680 5657
rect 5714 5623 5730 5657
rect 4245 5542 5071 5576
rect 5105 5542 5121 5576
rect 5664 5461 5680 5495
rect 5714 5461 5730 5495
rect 4177 5395 4279 5429
rect 7031 5395 7484 5429
rect 4245 5181 4279 5395
rect 5554 5349 5570 5383
rect 5604 5349 5620 5383
rect 5664 5259 5680 5293
rect 5714 5259 5730 5293
rect 4245 5147 4991 5181
rect 5025 5147 5041 5181
rect 5664 5035 5680 5069
rect 5714 5035 5730 5069
rect 5554 4945 5570 4979
rect 5604 4945 5620 4979
rect 4177 4899 4279 4933
rect 7031 4899 7484 4933
rect 4245 4786 4279 4899
rect 5664 4833 5680 4867
rect 5714 4833 5730 4867
rect 4245 4752 4911 4786
rect 4945 4752 4961 4786
rect 5664 4671 5680 4705
rect 5714 4671 5730 4705
rect 7031 4605 7484 4639
rect 5554 4559 5570 4593
rect 5604 4559 5620 4593
rect 5664 4469 5680 4503
rect 5714 4469 5730 4503
rect 5664 4245 5680 4279
rect 5714 4245 5730 4279
rect 5554 4155 5570 4189
rect 5604 4155 5620 4189
rect 7031 4109 7484 4143
rect 5664 4043 5680 4077
rect 5714 4043 5730 4077
rect 5664 3881 5680 3915
rect 5714 3881 5730 3915
rect 4177 3815 4279 3849
rect 7031 3815 7484 3849
rect 4245 3601 4279 3815
rect 5554 3769 5570 3803
rect 5604 3769 5620 3803
rect 5664 3679 5680 3713
rect 5714 3679 5730 3713
rect 4245 3567 4831 3601
rect 4865 3567 4881 3601
rect 5664 3455 5680 3489
rect 5714 3455 5730 3489
rect 5554 3365 5570 3399
rect 5604 3365 5620 3399
rect 4177 3319 4279 3353
rect 7031 3319 7484 3353
rect 4245 3206 4279 3319
rect 5664 3253 5680 3287
rect 5714 3253 5730 3287
rect 4245 3172 4751 3206
rect 4785 3172 4801 3206
rect 5664 3091 5680 3125
rect 5714 3091 5730 3125
rect 4177 3025 4279 3059
rect 7031 3025 7484 3059
rect 4245 2811 4279 3025
rect 5554 2979 5570 3013
rect 5604 2979 5620 3013
rect 5664 2889 5680 2923
rect 5714 2889 5730 2923
rect 4245 2777 4671 2811
rect 4705 2777 4721 2811
rect 5664 2665 5680 2699
rect 5714 2665 5730 2699
rect 5554 2575 5570 2609
rect 5604 2575 5620 2609
rect 4177 2529 4279 2563
rect 7031 2529 7484 2563
rect 4245 2416 4279 2529
rect 5664 2463 5680 2497
rect 5714 2463 5730 2497
rect 4245 2382 4591 2416
rect 4625 2382 4641 2416
rect 5664 2301 5680 2335
rect 5714 2301 5730 2335
rect 7031 2235 7484 2269
rect 5554 2189 5570 2223
rect 5604 2189 5620 2223
rect 5664 2099 5680 2133
rect 5714 2099 5730 2133
rect 5664 1875 5680 1909
rect 5714 1875 5730 1909
rect 5554 1785 5570 1819
rect 5604 1785 5620 1819
rect 7031 1739 7484 1773
rect 5664 1673 5680 1707
rect 5714 1673 5730 1707
rect 5664 1511 5680 1545
rect 5714 1511 5730 1545
rect 4177 1445 4279 1479
rect 7031 1445 7484 1479
rect 4245 1231 4279 1445
rect 5554 1399 5570 1433
rect 5604 1399 5620 1433
rect 5664 1309 5680 1343
rect 5714 1309 5730 1343
rect 4245 1197 4511 1231
rect 4545 1197 4561 1231
rect 5664 1085 5680 1119
rect 5714 1085 5730 1119
rect 5554 995 5570 1029
rect 5604 995 5620 1029
rect 4177 949 4279 983
rect 7031 949 7484 983
rect 4245 836 4279 949
rect 5664 883 5680 917
rect 5714 883 5730 917
rect 4245 802 4431 836
rect 4465 802 4481 836
rect 5664 721 5680 755
rect 5714 721 5730 755
rect 4177 655 4279 689
rect 7031 655 7484 689
rect 4245 441 4279 655
rect 5554 609 5570 643
rect 5604 609 5620 643
rect 5664 519 5680 553
rect 5714 519 5730 553
rect 4245 407 4351 441
rect 4385 407 4401 441
rect 5664 295 5680 329
rect 5714 295 5730 329
rect 5554 205 5570 239
rect 5604 205 5620 239
rect 4177 159 4279 193
rect 7031 159 7484 193
rect 4245 46 4279 159
rect 5664 93 5680 127
rect 5714 93 5730 127
rect 4245 12 4271 46
rect 4305 12 4321 46
<< viali >>
rect 5680 50491 5714 50525
rect 5570 50379 5604 50413
rect 5680 50289 5714 50323
rect 5680 50065 5714 50099
rect 5570 49975 5604 50009
rect 5680 49863 5714 49897
rect 5680 49701 5714 49735
rect 5570 49589 5604 49623
rect 5680 49499 5714 49533
rect 5680 49275 5714 49309
rect 5570 49185 5604 49219
rect 5680 49073 5714 49107
rect 5680 48911 5714 48945
rect 5570 48799 5604 48833
rect 5680 48709 5714 48743
rect 5680 48485 5714 48519
rect 5570 48395 5604 48429
rect 5680 48283 5714 48317
rect 5680 48121 5714 48155
rect 5570 48009 5604 48043
rect 5680 47919 5714 47953
rect 5680 47695 5714 47729
rect 5570 47605 5604 47639
rect 5680 47493 5714 47527
rect 5680 47331 5714 47365
rect 5570 47219 5604 47253
rect 5680 47129 5714 47163
rect 5680 46905 5714 46939
rect 5570 46815 5604 46849
rect 5680 46703 5714 46737
rect 5680 46541 5714 46575
rect 5570 46429 5604 46463
rect 5680 46339 5714 46373
rect 5680 46115 5714 46149
rect 5570 46025 5604 46059
rect 5680 45913 5714 45947
rect 5680 45751 5714 45785
rect 5570 45639 5604 45673
rect 5680 45549 5714 45583
rect 5680 45325 5714 45359
rect 5570 45235 5604 45269
rect 5680 45123 5714 45157
rect 5680 44961 5714 44995
rect 5570 44849 5604 44883
rect 5680 44759 5714 44793
rect 5680 44535 5714 44569
rect 5570 44445 5604 44479
rect 5680 44333 5714 44367
rect 5680 44171 5714 44205
rect 5570 44059 5604 44093
rect 5680 43969 5714 44003
rect 5680 43745 5714 43779
rect 5570 43655 5604 43689
rect 5680 43543 5714 43577
rect 5680 43381 5714 43415
rect 5570 43269 5604 43303
rect 5680 43179 5714 43213
rect 5680 42955 5714 42989
rect 5570 42865 5604 42899
rect 5680 42753 5714 42787
rect 5680 42591 5714 42625
rect 5570 42479 5604 42513
rect 5680 42389 5714 42423
rect 5680 42165 5714 42199
rect 5570 42075 5604 42109
rect 5680 41963 5714 41997
rect 5680 41801 5714 41835
rect 5570 41689 5604 41723
rect 5680 41599 5714 41633
rect 5680 41375 5714 41409
rect 5570 41285 5604 41319
rect 5680 41173 5714 41207
rect 5680 41011 5714 41045
rect 5570 40899 5604 40933
rect 5680 40809 5714 40843
rect 5680 40585 5714 40619
rect 5570 40495 5604 40529
rect 5680 40383 5714 40417
rect 5680 40221 5714 40255
rect 5570 40109 5604 40143
rect 5680 40019 5714 40053
rect 5680 39795 5714 39829
rect 5570 39705 5604 39739
rect 5680 39593 5714 39627
rect 5680 39431 5714 39465
rect 5570 39319 5604 39353
rect 5680 39229 5714 39263
rect 5680 39005 5714 39039
rect 5570 38915 5604 38949
rect 5680 38803 5714 38837
rect 5680 38641 5714 38675
rect 5570 38529 5604 38563
rect 5680 38439 5714 38473
rect 5680 38215 5714 38249
rect 5570 38125 5604 38159
rect 5680 38013 5714 38047
rect 5680 37851 5714 37885
rect 5570 37739 5604 37773
rect 5680 37649 5714 37683
rect 5680 37425 5714 37459
rect 5570 37335 5604 37369
rect 5680 37223 5714 37257
rect 5680 37061 5714 37095
rect 5570 36949 5604 36983
rect 5680 36859 5714 36893
rect 5680 36635 5714 36669
rect 5570 36545 5604 36579
rect 5680 36433 5714 36467
rect 5680 36271 5714 36305
rect 5570 36159 5604 36193
rect 5680 36069 5714 36103
rect 5680 35845 5714 35879
rect 5570 35755 5604 35789
rect 5680 35643 5714 35677
rect 5680 35481 5714 35515
rect 5570 35369 5604 35403
rect 5680 35279 5714 35313
rect 5680 35055 5714 35089
rect 5570 34965 5604 34999
rect 5680 34853 5714 34887
rect 5680 34691 5714 34725
rect 5570 34579 5604 34613
rect 5680 34489 5714 34523
rect 5680 34265 5714 34299
rect 5570 34175 5604 34209
rect 5680 34063 5714 34097
rect 5680 33901 5714 33935
rect 5570 33789 5604 33823
rect 5680 33699 5714 33733
rect 5680 33475 5714 33509
rect 5570 33385 5604 33419
rect 5680 33273 5714 33307
rect 5680 33111 5714 33145
rect 5570 32999 5604 33033
rect 5680 32909 5714 32943
rect 5680 32685 5714 32719
rect 5570 32595 5604 32629
rect 5680 32483 5714 32517
rect 5680 32321 5714 32355
rect 5570 32209 5604 32243
rect 5680 32119 5714 32153
rect 5680 31895 5714 31929
rect 5570 31805 5604 31839
rect 5680 31693 5714 31727
rect 5680 31531 5714 31565
rect 5570 31419 5604 31453
rect 5680 31329 5714 31363
rect 5680 31105 5714 31139
rect 5570 31015 5604 31049
rect 5680 30903 5714 30937
rect 5680 30741 5714 30775
rect 5570 30629 5604 30663
rect 5680 30539 5714 30573
rect 5680 30315 5714 30349
rect 5570 30225 5604 30259
rect 5680 30113 5714 30147
rect 5680 29951 5714 29985
rect 5570 29839 5604 29873
rect 5680 29749 5714 29783
rect 5680 29525 5714 29559
rect 5570 29435 5604 29469
rect 5680 29323 5714 29357
rect 5680 29161 5714 29195
rect 5570 29049 5604 29083
rect 5680 28959 5714 28993
rect 5680 28735 5714 28769
rect 5570 28645 5604 28679
rect 5680 28533 5714 28567
rect 5680 28371 5714 28405
rect 5570 28259 5604 28293
rect 5680 28169 5714 28203
rect 5680 27945 5714 27979
rect 5570 27855 5604 27889
rect 5680 27743 5714 27777
rect 5680 27581 5714 27615
rect 5570 27469 5604 27503
rect 5680 27379 5714 27413
rect 5680 27155 5714 27189
rect 5570 27065 5604 27099
rect 5680 26953 5714 26987
rect 5680 26791 5714 26825
rect 5570 26679 5604 26713
rect 5680 26589 5714 26623
rect 5680 26365 5714 26399
rect 5570 26275 5604 26309
rect 5680 26163 5714 26197
rect 5680 26001 5714 26035
rect 5570 25889 5604 25923
rect 5680 25799 5714 25833
rect 5680 25575 5714 25609
rect 5570 25485 5604 25519
rect 5680 25373 5714 25407
rect 5680 25211 5714 25245
rect 5570 25099 5604 25133
rect 5680 25009 5714 25043
rect 5680 24785 5714 24819
rect 5570 24695 5604 24729
rect 5680 24583 5714 24617
rect 5680 24421 5714 24455
rect 5570 24309 5604 24343
rect 5680 24219 5714 24253
rect 5680 23995 5714 24029
rect 5570 23905 5604 23939
rect 5680 23793 5714 23827
rect 5680 23631 5714 23665
rect 5570 23519 5604 23553
rect 5680 23429 5714 23463
rect 5680 23205 5714 23239
rect 5570 23115 5604 23149
rect 5680 23003 5714 23037
rect 5680 22841 5714 22875
rect 5570 22729 5604 22763
rect 5680 22639 5714 22673
rect 5680 22415 5714 22449
rect 5570 22325 5604 22359
rect 5680 22213 5714 22247
rect 5680 22051 5714 22085
rect 5570 21939 5604 21973
rect 5680 21849 5714 21883
rect 5680 21625 5714 21659
rect 5570 21535 5604 21569
rect 5680 21423 5714 21457
rect 5680 21261 5714 21295
rect 5570 21149 5604 21183
rect 5680 21059 5714 21093
rect 5680 20835 5714 20869
rect 5570 20745 5604 20779
rect 5680 20633 5714 20667
rect 5680 20471 5714 20505
rect 5570 20359 5604 20393
rect 5680 20269 5714 20303
rect 5680 20045 5714 20079
rect 5570 19955 5604 19989
rect 5680 19843 5714 19877
rect 5680 19681 5714 19715
rect 5570 19569 5604 19603
rect 5680 19479 5714 19513
rect 5680 19255 5714 19289
rect 5570 19165 5604 19199
rect 5680 19053 5714 19087
rect 5680 18891 5714 18925
rect 5570 18779 5604 18813
rect 5680 18689 5714 18723
rect 5680 18465 5714 18499
rect 5570 18375 5604 18409
rect 5680 18263 5714 18297
rect 5680 18101 5714 18135
rect 5570 17989 5604 18023
rect 5680 17899 5714 17933
rect 5680 17675 5714 17709
rect 5570 17585 5604 17619
rect 5680 17473 5714 17507
rect 5680 17311 5714 17345
rect 5570 17199 5604 17233
rect 5680 17109 5714 17143
rect 5680 16885 5714 16919
rect 5570 16795 5604 16829
rect 5680 16683 5714 16717
rect 5680 16521 5714 16555
rect 5570 16409 5604 16443
rect 5680 16319 5714 16353
rect 5680 16095 5714 16129
rect 5570 16005 5604 16039
rect 5680 15893 5714 15927
rect 5680 15731 5714 15765
rect 5570 15619 5604 15653
rect 5680 15529 5714 15563
rect 5680 15305 5714 15339
rect 5570 15215 5604 15249
rect 5680 15103 5714 15137
rect 5680 14941 5714 14975
rect 5570 14829 5604 14863
rect 5680 14739 5714 14773
rect 5680 14515 5714 14549
rect 5570 14425 5604 14459
rect 5680 14313 5714 14347
rect 5680 14151 5714 14185
rect 5570 14039 5604 14073
rect 5680 13949 5714 13983
rect 5680 13725 5714 13759
rect 5570 13635 5604 13669
rect 5680 13523 5714 13557
rect 5680 13361 5714 13395
rect 5570 13249 5604 13283
rect 5680 13159 5714 13193
rect 5680 12935 5714 12969
rect 5570 12845 5604 12879
rect 5680 12733 5714 12767
rect 5680 12571 5714 12605
rect 5570 12459 5604 12493
rect 5680 12369 5714 12403
rect 5680 12145 5714 12179
rect 5570 12055 5604 12089
rect 5680 11943 5714 11977
rect 5680 11781 5714 11815
rect 5570 11669 5604 11703
rect 5680 11579 5714 11613
rect 5680 11355 5714 11389
rect 5570 11265 5604 11299
rect 5680 11153 5714 11187
rect 5680 10991 5714 11025
rect 5570 10879 5604 10913
rect 5680 10789 5714 10823
rect 5680 10565 5714 10599
rect 5570 10475 5604 10509
rect 5680 10363 5714 10397
rect 5680 10201 5714 10235
rect 5570 10089 5604 10123
rect 5680 9999 5714 10033
rect 5680 9775 5714 9809
rect 5570 9685 5604 9719
rect 5680 9573 5714 9607
rect 5680 9411 5714 9445
rect 5570 9299 5604 9333
rect 5680 9209 5714 9243
rect 5680 8985 5714 9019
rect 5570 8895 5604 8929
rect 5680 8783 5714 8817
rect 5680 8621 5714 8655
rect 5570 8509 5604 8543
rect 5680 8419 5714 8453
rect 5680 8195 5714 8229
rect 5570 8105 5604 8139
rect 5680 7993 5714 8027
rect 5680 7831 5714 7865
rect 5570 7719 5604 7753
rect 5680 7629 5714 7663
rect 5471 7517 5505 7551
rect 5680 7405 5714 7439
rect 5570 7315 5604 7349
rect 5680 7203 5714 7237
rect 5391 7122 5425 7156
rect 5680 7041 5714 7075
rect 5570 6929 5604 6963
rect 5680 6839 5714 6873
rect 5311 6727 5345 6761
rect 5680 6615 5714 6649
rect 5570 6525 5604 6559
rect 5680 6413 5714 6447
rect 5231 6332 5265 6366
rect 5680 6251 5714 6285
rect 5570 6139 5604 6173
rect 5680 6049 5714 6083
rect 5151 5937 5185 5971
rect 5680 5825 5714 5859
rect 5570 5735 5604 5769
rect 5680 5623 5714 5657
rect 5071 5542 5105 5576
rect 5680 5461 5714 5495
rect 5570 5349 5604 5383
rect 5680 5259 5714 5293
rect 4991 5147 5025 5181
rect 5680 5035 5714 5069
rect 5570 4945 5604 4979
rect 5680 4833 5714 4867
rect 4911 4752 4945 4786
rect 5680 4671 5714 4705
rect 5570 4559 5604 4593
rect 5680 4469 5714 4503
rect 5680 4245 5714 4279
rect 5570 4155 5604 4189
rect 5680 4043 5714 4077
rect 5680 3881 5714 3915
rect 5570 3769 5604 3803
rect 5680 3679 5714 3713
rect 4831 3567 4865 3601
rect 5680 3455 5714 3489
rect 5570 3365 5604 3399
rect 5680 3253 5714 3287
rect 4751 3172 4785 3206
rect 5680 3091 5714 3125
rect 5570 2979 5604 3013
rect 5680 2889 5714 2923
rect 4671 2777 4705 2811
rect 5680 2665 5714 2699
rect 5570 2575 5604 2609
rect 5680 2463 5714 2497
rect 4591 2382 4625 2416
rect 5680 2301 5714 2335
rect 5570 2189 5604 2223
rect 5680 2099 5714 2133
rect 5680 1875 5714 1909
rect 5570 1785 5604 1819
rect 5680 1673 5714 1707
rect 5680 1511 5714 1545
rect 5570 1399 5604 1433
rect 5680 1309 5714 1343
rect 4511 1197 4545 1231
rect 5680 1085 5714 1119
rect 5570 995 5604 1029
rect 5680 883 5714 917
rect 4431 802 4465 836
rect 5680 721 5714 755
rect 5570 609 5604 643
rect 5680 519 5714 553
rect 4351 407 4385 441
rect 5680 295 5714 329
rect 5570 205 5604 239
rect 5680 93 5714 127
rect 4271 12 4305 46
<< metal1 >>
rect 4274 49122 4302 50617
rect 4354 49750 4382 50617
rect 4434 49912 4462 50617
rect 4514 50540 4542 50617
rect 4502 50534 4554 50540
rect 4502 50476 4554 50482
rect 4422 49906 4474 49912
rect 4422 49848 4474 49854
rect 4342 49744 4394 49750
rect 4342 49686 4394 49692
rect 4262 49116 4314 49122
rect 4262 49058 4314 49064
rect 4274 47542 4302 49058
rect 4354 48170 4382 49686
rect 4434 48332 4462 49848
rect 4514 48960 4542 50476
rect 4502 48954 4554 48960
rect 4502 48896 4554 48902
rect 4422 48326 4474 48332
rect 4422 48268 4474 48274
rect 4342 48164 4394 48170
rect 4342 48106 4394 48112
rect 4262 47536 4314 47542
rect 4262 47478 4314 47484
rect 4274 45962 4302 47478
rect 4354 46590 4382 48106
rect 4434 46752 4462 48268
rect 4514 47380 4542 48896
rect 4502 47374 4554 47380
rect 4502 47316 4554 47322
rect 4422 46746 4474 46752
rect 4422 46688 4474 46694
rect 4342 46584 4394 46590
rect 4342 46526 4394 46532
rect 4262 45956 4314 45962
rect 4262 45898 4314 45904
rect 4274 44382 4302 45898
rect 4354 45010 4382 46526
rect 4434 45172 4462 46688
rect 4514 45800 4542 47316
rect 4502 45794 4554 45800
rect 4502 45736 4554 45742
rect 4422 45166 4474 45172
rect 4422 45108 4474 45114
rect 4342 45004 4394 45010
rect 4342 44946 4394 44952
rect 4262 44376 4314 44382
rect 4262 44318 4314 44324
rect 4274 42802 4302 44318
rect 4354 43430 4382 44946
rect 4434 43592 4462 45108
rect 4514 44220 4542 45736
rect 4594 45688 4622 50617
rect 4674 47268 4702 50617
rect 4754 48848 4782 50617
rect 4834 50428 4862 50617
rect 4822 50422 4874 50428
rect 4822 50364 4874 50370
rect 4834 50024 4862 50364
rect 4822 50018 4874 50024
rect 4822 49960 4874 49966
rect 4834 49638 4862 49960
rect 4822 49632 4874 49638
rect 4822 49574 4874 49580
rect 4834 49234 4862 49574
rect 4822 49228 4874 49234
rect 4822 49170 4874 49176
rect 4742 48842 4794 48848
rect 4742 48784 4794 48790
rect 4754 48444 4782 48784
rect 4742 48438 4794 48444
rect 4742 48380 4794 48386
rect 4754 48058 4782 48380
rect 4742 48052 4794 48058
rect 4742 47994 4794 48000
rect 4754 47654 4782 47994
rect 4742 47648 4794 47654
rect 4742 47590 4794 47596
rect 4662 47262 4714 47268
rect 4662 47204 4714 47210
rect 4674 46864 4702 47204
rect 4662 46858 4714 46864
rect 4662 46800 4714 46806
rect 4674 46478 4702 46800
rect 4662 46472 4714 46478
rect 4662 46414 4714 46420
rect 4674 46074 4702 46414
rect 4662 46068 4714 46074
rect 4662 46010 4714 46016
rect 4582 45682 4634 45688
rect 4582 45624 4634 45630
rect 4594 45284 4622 45624
rect 4582 45278 4634 45284
rect 4582 45220 4634 45226
rect 4594 44898 4622 45220
rect 4582 44892 4634 44898
rect 4582 44834 4634 44840
rect 4594 44494 4622 44834
rect 4582 44488 4634 44494
rect 4582 44430 4634 44436
rect 4502 44214 4554 44220
rect 4502 44156 4554 44162
rect 4422 43586 4474 43592
rect 4422 43528 4474 43534
rect 4342 43424 4394 43430
rect 4342 43366 4394 43372
rect 4262 42796 4314 42802
rect 4262 42738 4314 42744
rect 4274 41222 4302 42738
rect 4354 41850 4382 43366
rect 4434 42012 4462 43528
rect 4514 42640 4542 44156
rect 4502 42634 4554 42640
rect 4502 42576 4554 42582
rect 4422 42006 4474 42012
rect 4422 41948 4474 41954
rect 4342 41844 4394 41850
rect 4342 41786 4394 41792
rect 4262 41216 4314 41222
rect 4262 41158 4314 41164
rect 4274 39642 4302 41158
rect 4354 40270 4382 41786
rect 4434 40432 4462 41948
rect 4514 41060 4542 42576
rect 4502 41054 4554 41060
rect 4502 40996 4554 41002
rect 4422 40426 4474 40432
rect 4422 40368 4474 40374
rect 4342 40264 4394 40270
rect 4342 40206 4394 40212
rect 4262 39636 4314 39642
rect 4262 39578 4314 39584
rect 4274 38062 4302 39578
rect 4354 38690 4382 40206
rect 4434 38852 4462 40368
rect 4514 39480 4542 40996
rect 4502 39474 4554 39480
rect 4502 39416 4554 39422
rect 4422 38846 4474 38852
rect 4422 38788 4474 38794
rect 4342 38684 4394 38690
rect 4342 38626 4394 38632
rect 4262 38056 4314 38062
rect 4262 37998 4314 38004
rect 4274 36482 4302 37998
rect 4354 37110 4382 38626
rect 4434 37272 4462 38788
rect 4514 37900 4542 39416
rect 4594 39368 4622 44430
rect 4674 40948 4702 46010
rect 4754 42528 4782 47590
rect 4834 44108 4862 49170
rect 4822 44102 4874 44108
rect 4822 44044 4874 44050
rect 4834 43704 4862 44044
rect 4822 43698 4874 43704
rect 4822 43640 4874 43646
rect 4834 43318 4862 43640
rect 4822 43312 4874 43318
rect 4822 43254 4874 43260
rect 4834 42914 4862 43254
rect 4822 42908 4874 42914
rect 4822 42850 4874 42856
rect 4742 42522 4794 42528
rect 4742 42464 4794 42470
rect 4754 42124 4782 42464
rect 4742 42118 4794 42124
rect 4742 42060 4794 42066
rect 4754 41738 4782 42060
rect 4742 41732 4794 41738
rect 4742 41674 4794 41680
rect 4754 41334 4782 41674
rect 4742 41328 4794 41334
rect 4742 41270 4794 41276
rect 4662 40942 4714 40948
rect 4662 40884 4714 40890
rect 4674 40544 4702 40884
rect 4662 40538 4714 40544
rect 4662 40480 4714 40486
rect 4674 40158 4702 40480
rect 4662 40152 4714 40158
rect 4662 40094 4714 40100
rect 4674 39754 4702 40094
rect 4662 39748 4714 39754
rect 4662 39690 4714 39696
rect 4582 39362 4634 39368
rect 4582 39304 4634 39310
rect 4594 38964 4622 39304
rect 4582 38958 4634 38964
rect 4582 38900 4634 38906
rect 4594 38578 4622 38900
rect 4582 38572 4634 38578
rect 4582 38514 4634 38520
rect 4594 38174 4622 38514
rect 4582 38168 4634 38174
rect 4582 38110 4634 38116
rect 4502 37894 4554 37900
rect 4502 37836 4554 37842
rect 4422 37266 4474 37272
rect 4422 37208 4474 37214
rect 4342 37104 4394 37110
rect 4342 37046 4394 37052
rect 4262 36476 4314 36482
rect 4262 36418 4314 36424
rect 4274 34902 4302 36418
rect 4354 35530 4382 37046
rect 4434 35692 4462 37208
rect 4514 36320 4542 37836
rect 4502 36314 4554 36320
rect 4502 36256 4554 36262
rect 4422 35686 4474 35692
rect 4422 35628 4474 35634
rect 4342 35524 4394 35530
rect 4342 35466 4394 35472
rect 4262 34896 4314 34902
rect 4262 34838 4314 34844
rect 4274 33322 4302 34838
rect 4354 33950 4382 35466
rect 4434 34112 4462 35628
rect 4514 34740 4542 36256
rect 4502 34734 4554 34740
rect 4502 34676 4554 34682
rect 4422 34106 4474 34112
rect 4422 34048 4474 34054
rect 4342 33944 4394 33950
rect 4342 33886 4394 33892
rect 4262 33316 4314 33322
rect 4262 33258 4314 33264
rect 4274 31742 4302 33258
rect 4354 32370 4382 33886
rect 4434 32532 4462 34048
rect 4514 33160 4542 34676
rect 4502 33154 4554 33160
rect 4502 33096 4554 33102
rect 4422 32526 4474 32532
rect 4422 32468 4474 32474
rect 4342 32364 4394 32370
rect 4342 32306 4394 32312
rect 4262 31736 4314 31742
rect 4262 31678 4314 31684
rect 4274 30162 4302 31678
rect 4354 30790 4382 32306
rect 4434 30952 4462 32468
rect 4514 31580 4542 33096
rect 4594 33048 4622 38110
rect 4674 34628 4702 39690
rect 4754 36208 4782 41270
rect 4834 37788 4862 42850
rect 4822 37782 4874 37788
rect 4822 37724 4874 37730
rect 4834 37384 4862 37724
rect 4822 37378 4874 37384
rect 4822 37320 4874 37326
rect 4834 36998 4862 37320
rect 4822 36992 4874 36998
rect 4822 36934 4874 36940
rect 4834 36594 4862 36934
rect 4822 36588 4874 36594
rect 4822 36530 4874 36536
rect 4742 36202 4794 36208
rect 4742 36144 4794 36150
rect 4754 35804 4782 36144
rect 4742 35798 4794 35804
rect 4742 35740 4794 35746
rect 4754 35418 4782 35740
rect 4742 35412 4794 35418
rect 4742 35354 4794 35360
rect 4754 35014 4782 35354
rect 4742 35008 4794 35014
rect 4742 34950 4794 34956
rect 4662 34622 4714 34628
rect 4662 34564 4714 34570
rect 4674 34224 4702 34564
rect 4662 34218 4714 34224
rect 4662 34160 4714 34166
rect 4674 33838 4702 34160
rect 4662 33832 4714 33838
rect 4662 33774 4714 33780
rect 4674 33434 4702 33774
rect 4662 33428 4714 33434
rect 4662 33370 4714 33376
rect 4582 33042 4634 33048
rect 4582 32984 4634 32990
rect 4594 32644 4622 32984
rect 4582 32638 4634 32644
rect 4582 32580 4634 32586
rect 4594 32258 4622 32580
rect 4582 32252 4634 32258
rect 4582 32194 4634 32200
rect 4594 31854 4622 32194
rect 4582 31848 4634 31854
rect 4582 31790 4634 31796
rect 4502 31574 4554 31580
rect 4502 31516 4554 31522
rect 4422 30946 4474 30952
rect 4422 30888 4474 30894
rect 4342 30784 4394 30790
rect 4342 30726 4394 30732
rect 4262 30156 4314 30162
rect 4262 30098 4314 30104
rect 4274 28582 4302 30098
rect 4354 29210 4382 30726
rect 4434 29372 4462 30888
rect 4514 30000 4542 31516
rect 4502 29994 4554 30000
rect 4502 29936 4554 29942
rect 4422 29366 4474 29372
rect 4422 29308 4474 29314
rect 4342 29204 4394 29210
rect 4342 29146 4394 29152
rect 4262 28576 4314 28582
rect 4262 28518 4314 28524
rect 4274 27002 4302 28518
rect 4354 27630 4382 29146
rect 4434 27792 4462 29308
rect 4514 28420 4542 29936
rect 4502 28414 4554 28420
rect 4502 28356 4554 28362
rect 4422 27786 4474 27792
rect 4422 27728 4474 27734
rect 4342 27624 4394 27630
rect 4342 27566 4394 27572
rect 4262 26996 4314 27002
rect 4262 26938 4314 26944
rect 4274 25422 4302 26938
rect 4354 26050 4382 27566
rect 4434 26212 4462 27728
rect 4514 26840 4542 28356
rect 4502 26834 4554 26840
rect 4502 26776 4554 26782
rect 4422 26206 4474 26212
rect 4422 26148 4474 26154
rect 4342 26044 4394 26050
rect 4342 25986 4394 25992
rect 4262 25416 4314 25422
rect 4262 25358 4314 25364
rect 4274 23842 4302 25358
rect 4354 24470 4382 25986
rect 4434 24632 4462 26148
rect 4514 25260 4542 26776
rect 4594 26728 4622 31790
rect 4674 28308 4702 33370
rect 4754 29888 4782 34950
rect 4834 31468 4862 36530
rect 4822 31462 4874 31468
rect 4822 31404 4874 31410
rect 4834 31064 4862 31404
rect 4822 31058 4874 31064
rect 4822 31000 4874 31006
rect 4834 30678 4862 31000
rect 4822 30672 4874 30678
rect 4822 30614 4874 30620
rect 4834 30274 4862 30614
rect 4822 30268 4874 30274
rect 4822 30210 4874 30216
rect 4742 29882 4794 29888
rect 4742 29824 4794 29830
rect 4754 29484 4782 29824
rect 4742 29478 4794 29484
rect 4742 29420 4794 29426
rect 4754 29098 4782 29420
rect 4742 29092 4794 29098
rect 4742 29034 4794 29040
rect 4754 28694 4782 29034
rect 4742 28688 4794 28694
rect 4742 28630 4794 28636
rect 4662 28302 4714 28308
rect 4662 28244 4714 28250
rect 4674 27904 4702 28244
rect 4662 27898 4714 27904
rect 4662 27840 4714 27846
rect 4674 27518 4702 27840
rect 4662 27512 4714 27518
rect 4662 27454 4714 27460
rect 4674 27114 4702 27454
rect 4662 27108 4714 27114
rect 4662 27050 4714 27056
rect 4582 26722 4634 26728
rect 4582 26664 4634 26670
rect 4594 26324 4622 26664
rect 4582 26318 4634 26324
rect 4582 26260 4634 26266
rect 4594 25938 4622 26260
rect 4582 25932 4634 25938
rect 4582 25874 4634 25880
rect 4594 25534 4622 25874
rect 4582 25528 4634 25534
rect 4582 25470 4634 25476
rect 4502 25254 4554 25260
rect 4502 25196 4554 25202
rect 4422 24626 4474 24632
rect 4422 24568 4474 24574
rect 4342 24464 4394 24470
rect 4342 24406 4394 24412
rect 4262 23836 4314 23842
rect 4262 23778 4314 23784
rect 4274 22262 4302 23778
rect 4354 22890 4382 24406
rect 4434 23052 4462 24568
rect 4514 23680 4542 25196
rect 4502 23674 4554 23680
rect 4502 23616 4554 23622
rect 4422 23046 4474 23052
rect 4422 22988 4474 22994
rect 4342 22884 4394 22890
rect 4342 22826 4394 22832
rect 4262 22256 4314 22262
rect 4262 22198 4314 22204
rect 4274 20682 4302 22198
rect 4354 21310 4382 22826
rect 4434 21472 4462 22988
rect 4514 22100 4542 23616
rect 4502 22094 4554 22100
rect 4502 22036 4554 22042
rect 4422 21466 4474 21472
rect 4422 21408 4474 21414
rect 4342 21304 4394 21310
rect 4342 21246 4394 21252
rect 4262 20676 4314 20682
rect 4262 20618 4314 20624
rect 4274 19102 4302 20618
rect 4354 19730 4382 21246
rect 4434 19892 4462 21408
rect 4514 20520 4542 22036
rect 4502 20514 4554 20520
rect 4502 20456 4554 20462
rect 4422 19886 4474 19892
rect 4422 19828 4474 19834
rect 4342 19724 4394 19730
rect 4342 19666 4394 19672
rect 4262 19096 4314 19102
rect 4262 19038 4314 19044
rect 4274 17522 4302 19038
rect 4354 18150 4382 19666
rect 4434 18312 4462 19828
rect 4514 18940 4542 20456
rect 4594 20408 4622 25470
rect 4674 21988 4702 27050
rect 4754 23568 4782 28630
rect 4834 25148 4862 30210
rect 4822 25142 4874 25148
rect 4822 25084 4874 25090
rect 4834 24744 4862 25084
rect 4822 24738 4874 24744
rect 4822 24680 4874 24686
rect 4834 24358 4862 24680
rect 4822 24352 4874 24358
rect 4822 24294 4874 24300
rect 4834 23954 4862 24294
rect 4822 23948 4874 23954
rect 4822 23890 4874 23896
rect 4742 23562 4794 23568
rect 4742 23504 4794 23510
rect 4754 23164 4782 23504
rect 4742 23158 4794 23164
rect 4742 23100 4794 23106
rect 4754 22778 4782 23100
rect 4742 22772 4794 22778
rect 4742 22714 4794 22720
rect 4754 22374 4782 22714
rect 4742 22368 4794 22374
rect 4742 22310 4794 22316
rect 4662 21982 4714 21988
rect 4662 21924 4714 21930
rect 4674 21584 4702 21924
rect 4662 21578 4714 21584
rect 4662 21520 4714 21526
rect 4674 21198 4702 21520
rect 4662 21192 4714 21198
rect 4662 21134 4714 21140
rect 4674 20794 4702 21134
rect 4662 20788 4714 20794
rect 4662 20730 4714 20736
rect 4582 20402 4634 20408
rect 4582 20344 4634 20350
rect 4594 20004 4622 20344
rect 4582 19998 4634 20004
rect 4582 19940 4634 19946
rect 4594 19618 4622 19940
rect 4582 19612 4634 19618
rect 4582 19554 4634 19560
rect 4594 19214 4622 19554
rect 4582 19208 4634 19214
rect 4582 19150 4634 19156
rect 4502 18934 4554 18940
rect 4502 18876 4554 18882
rect 4422 18306 4474 18312
rect 4422 18248 4474 18254
rect 4342 18144 4394 18150
rect 4342 18086 4394 18092
rect 4262 17516 4314 17522
rect 4262 17458 4314 17464
rect 4274 15942 4302 17458
rect 4354 16570 4382 18086
rect 4434 16732 4462 18248
rect 4514 17360 4542 18876
rect 4502 17354 4554 17360
rect 4502 17296 4554 17302
rect 4422 16726 4474 16732
rect 4422 16668 4474 16674
rect 4342 16564 4394 16570
rect 4342 16506 4394 16512
rect 4262 15936 4314 15942
rect 4262 15878 4314 15884
rect 4274 14362 4302 15878
rect 4354 14990 4382 16506
rect 4434 15152 4462 16668
rect 4514 15780 4542 17296
rect 4502 15774 4554 15780
rect 4502 15716 4554 15722
rect 4422 15146 4474 15152
rect 4422 15088 4474 15094
rect 4342 14984 4394 14990
rect 4342 14926 4394 14932
rect 4262 14356 4314 14362
rect 4262 14298 4314 14304
rect 4274 12782 4302 14298
rect 4354 13410 4382 14926
rect 4434 13572 4462 15088
rect 4514 14200 4542 15716
rect 4502 14194 4554 14200
rect 4502 14136 4554 14142
rect 4422 13566 4474 13572
rect 4422 13508 4474 13514
rect 4342 13404 4394 13410
rect 4342 13346 4394 13352
rect 4262 12776 4314 12782
rect 4262 12718 4314 12724
rect 4274 11202 4302 12718
rect 4354 11830 4382 13346
rect 4434 11992 4462 13508
rect 4514 12620 4542 14136
rect 4594 14088 4622 19150
rect 4674 15668 4702 20730
rect 4754 17248 4782 22310
rect 4834 18828 4862 23890
rect 4822 18822 4874 18828
rect 4822 18764 4874 18770
rect 4834 18424 4862 18764
rect 4822 18418 4874 18424
rect 4822 18360 4874 18366
rect 4834 18038 4862 18360
rect 4822 18032 4874 18038
rect 4822 17974 4874 17980
rect 4834 17634 4862 17974
rect 4822 17628 4874 17634
rect 4822 17570 4874 17576
rect 4742 17242 4794 17248
rect 4742 17184 4794 17190
rect 4754 16844 4782 17184
rect 4742 16838 4794 16844
rect 4742 16780 4794 16786
rect 4754 16458 4782 16780
rect 4742 16452 4794 16458
rect 4742 16394 4794 16400
rect 4754 16054 4782 16394
rect 4742 16048 4794 16054
rect 4742 15990 4794 15996
rect 4662 15662 4714 15668
rect 4662 15604 4714 15610
rect 4674 15264 4702 15604
rect 4662 15258 4714 15264
rect 4662 15200 4714 15206
rect 4674 14878 4702 15200
rect 4662 14872 4714 14878
rect 4662 14814 4714 14820
rect 4674 14474 4702 14814
rect 4662 14468 4714 14474
rect 4662 14410 4714 14416
rect 4582 14082 4634 14088
rect 4582 14024 4634 14030
rect 4594 13684 4622 14024
rect 4582 13678 4634 13684
rect 4582 13620 4634 13626
rect 4594 13298 4622 13620
rect 4582 13292 4634 13298
rect 4582 13234 4634 13240
rect 4594 12894 4622 13234
rect 4582 12888 4634 12894
rect 4582 12830 4634 12836
rect 4502 12614 4554 12620
rect 4502 12556 4554 12562
rect 4422 11986 4474 11992
rect 4422 11928 4474 11934
rect 4342 11824 4394 11830
rect 4342 11766 4394 11772
rect 4262 11196 4314 11202
rect 4262 11138 4314 11144
rect 4274 9622 4302 11138
rect 4354 10250 4382 11766
rect 4434 10412 4462 11928
rect 4514 11040 4542 12556
rect 4502 11034 4554 11040
rect 4502 10976 4554 10982
rect 4422 10406 4474 10412
rect 4422 10348 4474 10354
rect 4342 10244 4394 10250
rect 4342 10186 4394 10192
rect 4262 9616 4314 9622
rect 4262 9558 4314 9564
rect 4274 8042 4302 9558
rect 4354 8670 4382 10186
rect 4434 8832 4462 10348
rect 4514 9460 4542 10976
rect 4502 9454 4554 9460
rect 4502 9396 4554 9402
rect 4422 8826 4474 8832
rect 4422 8768 4474 8774
rect 4342 8664 4394 8670
rect 4342 8606 4394 8612
rect 4262 8036 4314 8042
rect 4262 7978 4314 7984
rect 18 258 46 7929
rect 98 654 126 7929
rect 178 2628 206 7929
rect 258 3024 286 7929
rect 338 4998 366 7929
rect 418 5394 446 7929
rect 498 5788 526 7929
rect 4274 6462 4302 7978
rect 4354 7090 4382 8606
rect 4434 7252 4462 8768
rect 4514 7880 4542 9396
rect 4502 7874 4554 7880
rect 4502 7816 4554 7822
rect 4422 7246 4474 7252
rect 4422 7188 4474 7194
rect 4342 7084 4394 7090
rect 4342 7026 4394 7032
rect 4262 6456 4314 6462
rect 4262 6398 4314 6404
rect 486 5782 538 5788
rect 828 5730 834 5782
rect 886 5730 892 5782
rect 486 5724 538 5730
rect 406 5388 458 5394
rect 406 5330 458 5336
rect 326 4992 378 4998
rect 326 4934 378 4940
rect 246 3018 298 3024
rect 246 2960 298 2966
rect 166 2622 218 2628
rect 166 2564 218 2570
rect 86 648 138 654
rect 86 590 138 596
rect 6 252 58 258
rect 6 194 58 200
rect 18 29 46 194
rect 98 29 126 590
rect 178 29 206 2564
rect 258 29 286 2960
rect 338 29 366 4934
rect 418 29 446 5330
rect 498 29 526 5724
rect 748 5336 754 5388
rect 806 5336 812 5388
rect 668 4940 674 4992
rect 726 4940 732 4992
rect 4274 4882 4302 6398
rect 4354 5510 4382 7026
rect 4434 5672 4462 7188
rect 4514 6300 4542 7816
rect 4594 7768 4622 12830
rect 4674 9348 4702 14410
rect 4754 10928 4782 15990
rect 4834 12508 4862 17570
rect 4822 12502 4874 12508
rect 4822 12444 4874 12450
rect 4834 12104 4862 12444
rect 4822 12098 4874 12104
rect 4822 12040 4874 12046
rect 4834 11718 4862 12040
rect 4822 11712 4874 11718
rect 4822 11654 4874 11660
rect 4834 11314 4862 11654
rect 4822 11308 4874 11314
rect 4822 11250 4874 11256
rect 4742 10922 4794 10928
rect 4742 10864 4794 10870
rect 4754 10524 4782 10864
rect 4742 10518 4794 10524
rect 4742 10460 4794 10466
rect 4754 10138 4782 10460
rect 4742 10132 4794 10138
rect 4742 10074 4794 10080
rect 4754 9734 4782 10074
rect 4742 9728 4794 9734
rect 4742 9670 4794 9676
rect 4662 9342 4714 9348
rect 4662 9284 4714 9290
rect 4674 8944 4702 9284
rect 4662 8938 4714 8944
rect 4662 8880 4714 8886
rect 4674 8558 4702 8880
rect 4662 8552 4714 8558
rect 4662 8494 4714 8500
rect 4674 8154 4702 8494
rect 4662 8148 4714 8154
rect 4662 8090 4714 8096
rect 4582 7762 4634 7768
rect 4582 7704 4634 7710
rect 4594 7364 4622 7704
rect 4582 7358 4634 7364
rect 4582 7300 4634 7306
rect 4594 6978 4622 7300
rect 4582 6972 4634 6978
rect 4582 6914 4634 6920
rect 4594 6574 4622 6914
rect 4582 6568 4634 6574
rect 4582 6510 4634 6516
rect 4502 6294 4554 6300
rect 4502 6236 4554 6242
rect 4422 5666 4474 5672
rect 4422 5608 4474 5614
rect 4342 5504 4394 5510
rect 4342 5446 4394 5452
rect 4262 4876 4314 4882
rect 4262 4818 4314 4824
rect 4274 3302 4302 4818
rect 4354 3930 4382 5446
rect 4434 4092 4462 5608
rect 4514 4720 4542 6236
rect 4502 4714 4554 4720
rect 4502 4656 4554 4662
rect 4422 4086 4474 4092
rect 4422 4028 4474 4034
rect 4342 3924 4394 3930
rect 4342 3866 4394 3872
rect 4262 3296 4314 3302
rect 4262 3238 4314 3244
rect 1424 2966 1430 3018
rect 1482 2966 1488 3018
rect 1344 2570 1350 2622
rect 1402 2570 1408 2622
rect 4274 1722 4302 3238
rect 4354 2350 4382 3866
rect 4434 2512 4462 4028
rect 4514 3140 4542 4656
rect 4502 3134 4554 3140
rect 4502 3076 4554 3082
rect 4422 2506 4474 2512
rect 4422 2448 4474 2454
rect 4342 2344 4394 2350
rect 4342 2286 4394 2292
rect 4262 1716 4314 1722
rect 4262 1658 4314 1664
rect 1424 596 1430 648
rect 1482 596 1488 648
rect 1344 200 1350 252
rect 1402 200 1408 252
rect 4274 142 4302 1658
rect 4354 770 4382 2286
rect 4434 932 4462 2448
rect 4514 1560 4542 3076
rect 4594 2428 4622 6510
rect 4674 3028 4702 8090
rect 4754 4608 4782 9670
rect 4834 6188 4862 11250
rect 4822 6182 4874 6188
rect 4822 6124 4874 6130
rect 4834 5784 4862 6124
rect 4914 6098 4942 50617
rect 4994 12418 5022 50617
rect 5074 18738 5102 50617
rect 5154 25058 5182 50617
rect 5234 31378 5262 50617
rect 5314 37698 5342 50617
rect 5394 44018 5422 50617
rect 5474 50338 5502 50617
rect 5665 50482 5671 50534
rect 5723 50482 5729 50534
rect 5555 50370 5561 50422
rect 5613 50370 5619 50422
rect 5462 50332 5514 50338
rect 5665 50280 5671 50332
rect 5723 50280 5729 50332
rect 5462 50274 5514 50280
rect 5474 50114 5502 50274
rect 5802 50243 5848 50545
rect 6226 50243 6274 50603
rect 6658 50243 6706 50603
rect 5793 50191 5799 50243
rect 5851 50191 5857 50243
rect 6218 50191 6224 50243
rect 6276 50191 6282 50243
rect 6650 50191 6656 50243
rect 6708 50191 6714 50243
rect 7050 50220 7078 50589
rect 7322 50220 7350 50589
rect 5462 50108 5514 50114
rect 5665 50056 5671 50108
rect 5723 50056 5729 50108
rect 5462 50050 5514 50056
rect 5474 49548 5502 50050
rect 5555 49966 5561 50018
rect 5613 49966 5619 50018
rect 5665 49854 5671 49906
rect 5723 49854 5729 49906
rect 5802 49869 5848 50191
rect 5793 49817 5799 49869
rect 5851 49817 5857 49869
rect 5665 49692 5671 49744
rect 5723 49692 5729 49744
rect 5555 49580 5561 49632
rect 5613 49580 5619 49632
rect 5462 49542 5514 49548
rect 5665 49490 5671 49542
rect 5723 49490 5729 49542
rect 5462 49484 5514 49490
rect 5474 49324 5502 49484
rect 5802 49453 5848 49817
rect 6226 49811 6274 50191
rect 6658 49811 6706 50191
rect 7032 50168 7038 50220
rect 7090 50168 7096 50220
rect 7304 50168 7310 50220
rect 7362 50168 7368 50220
rect 7050 49825 7078 50168
rect 7322 49825 7350 50168
rect 6218 49759 6224 49811
rect 6276 49759 6282 49811
rect 6650 49759 6656 49811
rect 6708 49759 6714 49811
rect 7032 49773 7038 49825
rect 7090 49773 7096 49825
rect 7304 49773 7310 49825
rect 7362 49773 7368 49825
rect 6226 49453 6274 49759
rect 6658 49453 6706 49759
rect 5793 49401 5799 49453
rect 5851 49401 5857 49453
rect 6218 49401 6224 49453
rect 6276 49401 6282 49453
rect 6650 49401 6656 49453
rect 6708 49401 6714 49453
rect 7050 49430 7078 49773
rect 7322 49430 7350 49773
rect 5462 49318 5514 49324
rect 5665 49266 5671 49318
rect 5723 49266 5729 49318
rect 5462 49260 5514 49266
rect 5474 48758 5502 49260
rect 5555 49176 5561 49228
rect 5613 49176 5619 49228
rect 5665 49064 5671 49116
rect 5723 49064 5729 49116
rect 5802 49079 5848 49401
rect 5793 49027 5799 49079
rect 5851 49027 5857 49079
rect 5665 48902 5671 48954
rect 5723 48902 5729 48954
rect 5555 48790 5561 48842
rect 5613 48790 5619 48842
rect 5462 48752 5514 48758
rect 5665 48700 5671 48752
rect 5723 48700 5729 48752
rect 5462 48694 5514 48700
rect 5474 48534 5502 48694
rect 5802 48663 5848 49027
rect 6226 49021 6274 49401
rect 6658 49021 6706 49401
rect 7032 49378 7038 49430
rect 7090 49378 7096 49430
rect 7304 49378 7310 49430
rect 7362 49378 7368 49430
rect 7050 49035 7078 49378
rect 7322 49035 7350 49378
rect 6218 48969 6224 49021
rect 6276 48969 6282 49021
rect 6650 48969 6656 49021
rect 6708 48969 6714 49021
rect 7032 48983 7038 49035
rect 7090 48983 7096 49035
rect 7304 48983 7310 49035
rect 7362 48983 7368 49035
rect 6226 48663 6274 48969
rect 6658 48663 6706 48969
rect 5793 48611 5799 48663
rect 5851 48611 5857 48663
rect 6218 48611 6224 48663
rect 6276 48611 6282 48663
rect 6650 48611 6656 48663
rect 6708 48611 6714 48663
rect 7050 48640 7078 48983
rect 7322 48640 7350 48983
rect 5462 48528 5514 48534
rect 5665 48476 5671 48528
rect 5723 48476 5729 48528
rect 5462 48470 5514 48476
rect 5474 47968 5502 48470
rect 5555 48386 5561 48438
rect 5613 48386 5619 48438
rect 5665 48274 5671 48326
rect 5723 48274 5729 48326
rect 5802 48289 5848 48611
rect 5793 48237 5799 48289
rect 5851 48237 5857 48289
rect 5665 48112 5671 48164
rect 5723 48112 5729 48164
rect 5555 48000 5561 48052
rect 5613 48000 5619 48052
rect 5462 47962 5514 47968
rect 5665 47910 5671 47962
rect 5723 47910 5729 47962
rect 5462 47904 5514 47910
rect 5474 47744 5502 47904
rect 5802 47873 5848 48237
rect 6226 48231 6274 48611
rect 6658 48231 6706 48611
rect 7032 48588 7038 48640
rect 7090 48588 7096 48640
rect 7304 48588 7310 48640
rect 7362 48588 7368 48640
rect 7050 48245 7078 48588
rect 7322 48245 7350 48588
rect 6218 48179 6224 48231
rect 6276 48179 6282 48231
rect 6650 48179 6656 48231
rect 6708 48179 6714 48231
rect 7032 48193 7038 48245
rect 7090 48193 7096 48245
rect 7304 48193 7310 48245
rect 7362 48193 7368 48245
rect 6226 47873 6274 48179
rect 6658 47873 6706 48179
rect 5793 47821 5799 47873
rect 5851 47821 5857 47873
rect 6218 47821 6224 47873
rect 6276 47821 6282 47873
rect 6650 47821 6656 47873
rect 6708 47821 6714 47873
rect 7050 47850 7078 48193
rect 7322 47850 7350 48193
rect 5462 47738 5514 47744
rect 5665 47686 5671 47738
rect 5723 47686 5729 47738
rect 5462 47680 5514 47686
rect 5474 47178 5502 47680
rect 5555 47596 5561 47648
rect 5613 47596 5619 47648
rect 5665 47484 5671 47536
rect 5723 47484 5729 47536
rect 5802 47499 5848 47821
rect 5793 47447 5799 47499
rect 5851 47447 5857 47499
rect 5665 47322 5671 47374
rect 5723 47322 5729 47374
rect 5555 47210 5561 47262
rect 5613 47210 5619 47262
rect 5462 47172 5514 47178
rect 5665 47120 5671 47172
rect 5723 47120 5729 47172
rect 5462 47114 5514 47120
rect 5474 46954 5502 47114
rect 5802 47083 5848 47447
rect 6226 47441 6274 47821
rect 6658 47441 6706 47821
rect 7032 47798 7038 47850
rect 7090 47798 7096 47850
rect 7304 47798 7310 47850
rect 7362 47798 7368 47850
rect 7050 47455 7078 47798
rect 7322 47455 7350 47798
rect 6218 47389 6224 47441
rect 6276 47389 6282 47441
rect 6650 47389 6656 47441
rect 6708 47389 6714 47441
rect 7032 47403 7038 47455
rect 7090 47403 7096 47455
rect 7304 47403 7310 47455
rect 7362 47403 7368 47455
rect 6226 47083 6274 47389
rect 6658 47083 6706 47389
rect 5793 47031 5799 47083
rect 5851 47031 5857 47083
rect 6218 47031 6224 47083
rect 6276 47031 6282 47083
rect 6650 47031 6656 47083
rect 6708 47031 6714 47083
rect 7050 47060 7078 47403
rect 7322 47060 7350 47403
rect 5462 46948 5514 46954
rect 5665 46896 5671 46948
rect 5723 46896 5729 46948
rect 5462 46890 5514 46896
rect 5474 46388 5502 46890
rect 5555 46806 5561 46858
rect 5613 46806 5619 46858
rect 5665 46694 5671 46746
rect 5723 46694 5729 46746
rect 5802 46709 5848 47031
rect 5793 46657 5799 46709
rect 5851 46657 5857 46709
rect 5665 46532 5671 46584
rect 5723 46532 5729 46584
rect 5555 46420 5561 46472
rect 5613 46420 5619 46472
rect 5462 46382 5514 46388
rect 5665 46330 5671 46382
rect 5723 46330 5729 46382
rect 5462 46324 5514 46330
rect 5474 46164 5502 46324
rect 5802 46293 5848 46657
rect 6226 46651 6274 47031
rect 6658 46651 6706 47031
rect 7032 47008 7038 47060
rect 7090 47008 7096 47060
rect 7304 47008 7310 47060
rect 7362 47008 7368 47060
rect 7050 46665 7078 47008
rect 7322 46665 7350 47008
rect 6218 46599 6224 46651
rect 6276 46599 6282 46651
rect 6650 46599 6656 46651
rect 6708 46599 6714 46651
rect 7032 46613 7038 46665
rect 7090 46613 7096 46665
rect 7304 46613 7310 46665
rect 7362 46613 7368 46665
rect 6226 46293 6274 46599
rect 6658 46293 6706 46599
rect 5793 46241 5799 46293
rect 5851 46241 5857 46293
rect 6218 46241 6224 46293
rect 6276 46241 6282 46293
rect 6650 46241 6656 46293
rect 6708 46241 6714 46293
rect 7050 46270 7078 46613
rect 7322 46270 7350 46613
rect 5462 46158 5514 46164
rect 5665 46106 5671 46158
rect 5723 46106 5729 46158
rect 5462 46100 5514 46106
rect 5474 45598 5502 46100
rect 5555 46016 5561 46068
rect 5613 46016 5619 46068
rect 5665 45904 5671 45956
rect 5723 45904 5729 45956
rect 5802 45919 5848 46241
rect 5793 45867 5799 45919
rect 5851 45867 5857 45919
rect 5665 45742 5671 45794
rect 5723 45742 5729 45794
rect 5555 45630 5561 45682
rect 5613 45630 5619 45682
rect 5462 45592 5514 45598
rect 5665 45540 5671 45592
rect 5723 45540 5729 45592
rect 5462 45534 5514 45540
rect 5474 45374 5502 45534
rect 5802 45503 5848 45867
rect 6226 45861 6274 46241
rect 6658 45861 6706 46241
rect 7032 46218 7038 46270
rect 7090 46218 7096 46270
rect 7304 46218 7310 46270
rect 7362 46218 7368 46270
rect 7050 45875 7078 46218
rect 7322 45875 7350 46218
rect 6218 45809 6224 45861
rect 6276 45809 6282 45861
rect 6650 45809 6656 45861
rect 6708 45809 6714 45861
rect 7032 45823 7038 45875
rect 7090 45823 7096 45875
rect 7304 45823 7310 45875
rect 7362 45823 7368 45875
rect 6226 45503 6274 45809
rect 6658 45503 6706 45809
rect 5793 45451 5799 45503
rect 5851 45451 5857 45503
rect 6218 45451 6224 45503
rect 6276 45451 6282 45503
rect 6650 45451 6656 45503
rect 6708 45451 6714 45503
rect 7050 45480 7078 45823
rect 7322 45480 7350 45823
rect 5462 45368 5514 45374
rect 5665 45316 5671 45368
rect 5723 45316 5729 45368
rect 5462 45310 5514 45316
rect 5474 44808 5502 45310
rect 5555 45226 5561 45278
rect 5613 45226 5619 45278
rect 5665 45114 5671 45166
rect 5723 45114 5729 45166
rect 5802 45129 5848 45451
rect 5793 45077 5799 45129
rect 5851 45077 5857 45129
rect 5665 44952 5671 45004
rect 5723 44952 5729 45004
rect 5555 44840 5561 44892
rect 5613 44840 5619 44892
rect 5462 44802 5514 44808
rect 5665 44750 5671 44802
rect 5723 44750 5729 44802
rect 5462 44744 5514 44750
rect 5474 44584 5502 44744
rect 5802 44713 5848 45077
rect 6226 45071 6274 45451
rect 6658 45071 6706 45451
rect 7032 45428 7038 45480
rect 7090 45428 7096 45480
rect 7304 45428 7310 45480
rect 7362 45428 7368 45480
rect 7050 45085 7078 45428
rect 7322 45085 7350 45428
rect 6218 45019 6224 45071
rect 6276 45019 6282 45071
rect 6650 45019 6656 45071
rect 6708 45019 6714 45071
rect 7032 45033 7038 45085
rect 7090 45033 7096 45085
rect 7304 45033 7310 45085
rect 7362 45033 7368 45085
rect 6226 44713 6274 45019
rect 6658 44713 6706 45019
rect 5793 44661 5799 44713
rect 5851 44661 5857 44713
rect 6218 44661 6224 44713
rect 6276 44661 6282 44713
rect 6650 44661 6656 44713
rect 6708 44661 6714 44713
rect 7050 44690 7078 45033
rect 7322 44690 7350 45033
rect 5462 44578 5514 44584
rect 5665 44526 5671 44578
rect 5723 44526 5729 44578
rect 5462 44520 5514 44526
rect 5382 44012 5434 44018
rect 5382 43954 5434 43960
rect 5394 43794 5422 43954
rect 5382 43788 5434 43794
rect 5382 43730 5434 43736
rect 5394 43228 5422 43730
rect 5382 43222 5434 43228
rect 5382 43164 5434 43170
rect 5394 43004 5422 43164
rect 5382 42998 5434 43004
rect 5382 42940 5434 42946
rect 5394 42438 5422 42940
rect 5382 42432 5434 42438
rect 5382 42374 5434 42380
rect 5394 42214 5422 42374
rect 5382 42208 5434 42214
rect 5382 42150 5434 42156
rect 5394 41648 5422 42150
rect 5382 41642 5434 41648
rect 5382 41584 5434 41590
rect 5394 41424 5422 41584
rect 5382 41418 5434 41424
rect 5382 41360 5434 41366
rect 5394 40858 5422 41360
rect 5382 40852 5434 40858
rect 5382 40794 5434 40800
rect 5394 40634 5422 40794
rect 5382 40628 5434 40634
rect 5382 40570 5434 40576
rect 5394 40068 5422 40570
rect 5382 40062 5434 40068
rect 5382 40004 5434 40010
rect 5394 39844 5422 40004
rect 5382 39838 5434 39844
rect 5382 39780 5434 39786
rect 5394 39278 5422 39780
rect 5382 39272 5434 39278
rect 5382 39214 5434 39220
rect 5394 39054 5422 39214
rect 5382 39048 5434 39054
rect 5382 38990 5434 38996
rect 5394 38488 5422 38990
rect 5382 38482 5434 38488
rect 5382 38424 5434 38430
rect 5394 38264 5422 38424
rect 5382 38258 5434 38264
rect 5382 38200 5434 38206
rect 5302 37692 5354 37698
rect 5302 37634 5354 37640
rect 5314 37474 5342 37634
rect 5302 37468 5354 37474
rect 5302 37410 5354 37416
rect 5314 36908 5342 37410
rect 5302 36902 5354 36908
rect 5302 36844 5354 36850
rect 5314 36684 5342 36844
rect 5302 36678 5354 36684
rect 5302 36620 5354 36626
rect 5314 36118 5342 36620
rect 5302 36112 5354 36118
rect 5302 36054 5354 36060
rect 5314 35894 5342 36054
rect 5302 35888 5354 35894
rect 5302 35830 5354 35836
rect 5314 35328 5342 35830
rect 5302 35322 5354 35328
rect 5302 35264 5354 35270
rect 5314 35104 5342 35264
rect 5302 35098 5354 35104
rect 5302 35040 5354 35046
rect 5314 34538 5342 35040
rect 5302 34532 5354 34538
rect 5302 34474 5354 34480
rect 5314 34314 5342 34474
rect 5302 34308 5354 34314
rect 5302 34250 5354 34256
rect 5314 33748 5342 34250
rect 5302 33742 5354 33748
rect 5302 33684 5354 33690
rect 5314 33524 5342 33684
rect 5302 33518 5354 33524
rect 5302 33460 5354 33466
rect 5314 32958 5342 33460
rect 5302 32952 5354 32958
rect 5302 32894 5354 32900
rect 5314 32734 5342 32894
rect 5302 32728 5354 32734
rect 5302 32670 5354 32676
rect 5314 32168 5342 32670
rect 5302 32162 5354 32168
rect 5302 32104 5354 32110
rect 5314 31944 5342 32104
rect 5302 31938 5354 31944
rect 5302 31880 5354 31886
rect 5222 31372 5274 31378
rect 5222 31314 5274 31320
rect 5234 31154 5262 31314
rect 5222 31148 5274 31154
rect 5222 31090 5274 31096
rect 5234 30588 5262 31090
rect 5222 30582 5274 30588
rect 5222 30524 5274 30530
rect 5234 30364 5262 30524
rect 5222 30358 5274 30364
rect 5222 30300 5274 30306
rect 5234 29798 5262 30300
rect 5222 29792 5274 29798
rect 5222 29734 5274 29740
rect 5234 29574 5262 29734
rect 5222 29568 5274 29574
rect 5222 29510 5274 29516
rect 5234 29008 5262 29510
rect 5222 29002 5274 29008
rect 5222 28944 5274 28950
rect 5234 28784 5262 28944
rect 5222 28778 5274 28784
rect 5222 28720 5274 28726
rect 5234 28218 5262 28720
rect 5222 28212 5274 28218
rect 5222 28154 5274 28160
rect 5234 27994 5262 28154
rect 5222 27988 5274 27994
rect 5222 27930 5274 27936
rect 5234 27428 5262 27930
rect 5222 27422 5274 27428
rect 5222 27364 5274 27370
rect 5234 27204 5262 27364
rect 5222 27198 5274 27204
rect 5222 27140 5274 27146
rect 5234 26638 5262 27140
rect 5222 26632 5274 26638
rect 5222 26574 5274 26580
rect 5234 26414 5262 26574
rect 5222 26408 5274 26414
rect 5222 26350 5274 26356
rect 5234 25848 5262 26350
rect 5222 25842 5274 25848
rect 5222 25784 5274 25790
rect 5234 25624 5262 25784
rect 5222 25618 5274 25624
rect 5222 25560 5274 25566
rect 5142 25052 5194 25058
rect 5142 24994 5194 25000
rect 5154 24834 5182 24994
rect 5142 24828 5194 24834
rect 5142 24770 5194 24776
rect 5154 24268 5182 24770
rect 5142 24262 5194 24268
rect 5142 24204 5194 24210
rect 5154 24044 5182 24204
rect 5142 24038 5194 24044
rect 5142 23980 5194 23986
rect 5154 23478 5182 23980
rect 5142 23472 5194 23478
rect 5142 23414 5194 23420
rect 5154 23254 5182 23414
rect 5142 23248 5194 23254
rect 5142 23190 5194 23196
rect 5154 22688 5182 23190
rect 5142 22682 5194 22688
rect 5142 22624 5194 22630
rect 5154 22464 5182 22624
rect 5142 22458 5194 22464
rect 5142 22400 5194 22406
rect 5154 21898 5182 22400
rect 5142 21892 5194 21898
rect 5142 21834 5194 21840
rect 5154 21674 5182 21834
rect 5142 21668 5194 21674
rect 5142 21610 5194 21616
rect 5154 21108 5182 21610
rect 5142 21102 5194 21108
rect 5142 21044 5194 21050
rect 5154 20884 5182 21044
rect 5142 20878 5194 20884
rect 5142 20820 5194 20826
rect 5154 20318 5182 20820
rect 5142 20312 5194 20318
rect 5142 20254 5194 20260
rect 5154 20094 5182 20254
rect 5142 20088 5194 20094
rect 5142 20030 5194 20036
rect 5154 19528 5182 20030
rect 5142 19522 5194 19528
rect 5142 19464 5194 19470
rect 5154 19304 5182 19464
rect 5142 19298 5194 19304
rect 5142 19240 5194 19246
rect 5062 18732 5114 18738
rect 5062 18674 5114 18680
rect 5074 18514 5102 18674
rect 5062 18508 5114 18514
rect 5062 18450 5114 18456
rect 5074 17948 5102 18450
rect 5062 17942 5114 17948
rect 5062 17884 5114 17890
rect 5074 17724 5102 17884
rect 5062 17718 5114 17724
rect 5062 17660 5114 17666
rect 5074 17158 5102 17660
rect 5062 17152 5114 17158
rect 5062 17094 5114 17100
rect 5074 16934 5102 17094
rect 5062 16928 5114 16934
rect 5062 16870 5114 16876
rect 5074 16368 5102 16870
rect 5062 16362 5114 16368
rect 5062 16304 5114 16310
rect 5074 16144 5102 16304
rect 5062 16138 5114 16144
rect 5062 16080 5114 16086
rect 5074 15578 5102 16080
rect 5062 15572 5114 15578
rect 5062 15514 5114 15520
rect 5074 15354 5102 15514
rect 5062 15348 5114 15354
rect 5062 15290 5114 15296
rect 5074 14788 5102 15290
rect 5062 14782 5114 14788
rect 5062 14724 5114 14730
rect 5074 14564 5102 14724
rect 5062 14558 5114 14564
rect 5062 14500 5114 14506
rect 5074 13998 5102 14500
rect 5062 13992 5114 13998
rect 5062 13934 5114 13940
rect 5074 13774 5102 13934
rect 5062 13768 5114 13774
rect 5062 13710 5114 13716
rect 5074 13208 5102 13710
rect 5062 13202 5114 13208
rect 5062 13144 5114 13150
rect 5074 12984 5102 13144
rect 5062 12978 5114 12984
rect 5062 12920 5114 12926
rect 4982 12412 5034 12418
rect 4982 12354 5034 12360
rect 4994 12194 5022 12354
rect 4982 12188 5034 12194
rect 4982 12130 5034 12136
rect 4994 11628 5022 12130
rect 4982 11622 5034 11628
rect 4982 11564 5034 11570
rect 4994 11404 5022 11564
rect 4982 11398 5034 11404
rect 4982 11340 5034 11346
rect 4994 10838 5022 11340
rect 4982 10832 5034 10838
rect 4982 10774 5034 10780
rect 4994 10614 5022 10774
rect 4982 10608 5034 10614
rect 4982 10550 5034 10556
rect 4994 10048 5022 10550
rect 4982 10042 5034 10048
rect 4982 9984 5034 9990
rect 4994 9824 5022 9984
rect 4982 9818 5034 9824
rect 4982 9760 5034 9766
rect 4994 9258 5022 9760
rect 4982 9252 5034 9258
rect 4982 9194 5034 9200
rect 4994 9034 5022 9194
rect 4982 9028 5034 9034
rect 4982 8970 5034 8976
rect 4994 8468 5022 8970
rect 4982 8462 5034 8468
rect 4982 8404 5034 8410
rect 4994 8244 5022 8404
rect 4982 8238 5034 8244
rect 4982 8180 5034 8186
rect 4994 7678 5022 8180
rect 4982 7672 5034 7678
rect 4982 7614 5034 7620
rect 4994 7454 5022 7614
rect 4982 7448 5034 7454
rect 4982 7390 5034 7396
rect 4994 6888 5022 7390
rect 4982 6882 5034 6888
rect 4982 6824 5034 6830
rect 4994 6664 5022 6824
rect 4982 6658 5034 6664
rect 4982 6600 5034 6606
rect 4902 6092 4954 6098
rect 4902 6034 4954 6040
rect 4914 5874 4942 6034
rect 4902 5868 4954 5874
rect 4902 5810 4954 5816
rect 4822 5778 4874 5784
rect 4822 5720 4874 5726
rect 4834 5398 4862 5720
rect 4822 5392 4874 5398
rect 4822 5334 4874 5340
rect 4834 4994 4862 5334
rect 4914 5308 4942 5810
rect 4902 5302 4954 5308
rect 4902 5244 4954 5250
rect 4914 5084 4942 5244
rect 4994 5193 5022 6600
rect 5074 5588 5102 12920
rect 5154 5983 5182 19240
rect 5234 6378 5262 25560
rect 5314 6773 5342 31880
rect 5394 7168 5422 38200
rect 5474 7563 5502 44520
rect 5555 44436 5561 44488
rect 5613 44436 5619 44488
rect 5665 44324 5671 44376
rect 5723 44324 5729 44376
rect 5802 44339 5848 44661
rect 5793 44287 5799 44339
rect 5851 44287 5857 44339
rect 5665 44162 5671 44214
rect 5723 44162 5729 44214
rect 5555 44050 5561 44102
rect 5613 44050 5619 44102
rect 5665 43960 5671 44012
rect 5723 43960 5729 44012
rect 5802 43923 5848 44287
rect 6226 44281 6274 44661
rect 6658 44281 6706 44661
rect 7032 44638 7038 44690
rect 7090 44638 7096 44690
rect 7304 44638 7310 44690
rect 7362 44638 7368 44690
rect 7050 44295 7078 44638
rect 7322 44295 7350 44638
rect 6218 44229 6224 44281
rect 6276 44229 6282 44281
rect 6650 44229 6656 44281
rect 6708 44229 6714 44281
rect 7032 44243 7038 44295
rect 7090 44243 7096 44295
rect 7304 44243 7310 44295
rect 7362 44243 7368 44295
rect 6226 43923 6274 44229
rect 6658 43923 6706 44229
rect 5793 43871 5799 43923
rect 5851 43871 5857 43923
rect 6218 43871 6224 43923
rect 6276 43871 6282 43923
rect 6650 43871 6656 43923
rect 6708 43871 6714 43923
rect 7050 43900 7078 44243
rect 7322 43900 7350 44243
rect 5665 43736 5671 43788
rect 5723 43736 5729 43788
rect 5555 43646 5561 43698
rect 5613 43646 5619 43698
rect 5665 43534 5671 43586
rect 5723 43534 5729 43586
rect 5802 43549 5848 43871
rect 5793 43497 5799 43549
rect 5851 43497 5857 43549
rect 5665 43372 5671 43424
rect 5723 43372 5729 43424
rect 5555 43260 5561 43312
rect 5613 43260 5619 43312
rect 5665 43170 5671 43222
rect 5723 43170 5729 43222
rect 5802 43133 5848 43497
rect 6226 43491 6274 43871
rect 6658 43491 6706 43871
rect 7032 43848 7038 43900
rect 7090 43848 7096 43900
rect 7304 43848 7310 43900
rect 7362 43848 7368 43900
rect 7050 43505 7078 43848
rect 7322 43505 7350 43848
rect 6218 43439 6224 43491
rect 6276 43439 6282 43491
rect 6650 43439 6656 43491
rect 6708 43439 6714 43491
rect 7032 43453 7038 43505
rect 7090 43453 7096 43505
rect 7304 43453 7310 43505
rect 7362 43453 7368 43505
rect 6226 43133 6274 43439
rect 6658 43133 6706 43439
rect 5793 43081 5799 43133
rect 5851 43081 5857 43133
rect 6218 43081 6224 43133
rect 6276 43081 6282 43133
rect 6650 43081 6656 43133
rect 6708 43081 6714 43133
rect 7050 43110 7078 43453
rect 7322 43110 7350 43453
rect 5665 42946 5671 42998
rect 5723 42946 5729 42998
rect 5555 42856 5561 42908
rect 5613 42856 5619 42908
rect 5665 42744 5671 42796
rect 5723 42744 5729 42796
rect 5802 42759 5848 43081
rect 5793 42707 5799 42759
rect 5851 42707 5857 42759
rect 5665 42582 5671 42634
rect 5723 42582 5729 42634
rect 5555 42470 5561 42522
rect 5613 42470 5619 42522
rect 5665 42380 5671 42432
rect 5723 42380 5729 42432
rect 5802 42343 5848 42707
rect 6226 42701 6274 43081
rect 6658 42701 6706 43081
rect 7032 43058 7038 43110
rect 7090 43058 7096 43110
rect 7304 43058 7310 43110
rect 7362 43058 7368 43110
rect 7050 42715 7078 43058
rect 7322 42715 7350 43058
rect 6218 42649 6224 42701
rect 6276 42649 6282 42701
rect 6650 42649 6656 42701
rect 6708 42649 6714 42701
rect 7032 42663 7038 42715
rect 7090 42663 7096 42715
rect 7304 42663 7310 42715
rect 7362 42663 7368 42715
rect 6226 42343 6274 42649
rect 6658 42343 6706 42649
rect 5793 42291 5799 42343
rect 5851 42291 5857 42343
rect 6218 42291 6224 42343
rect 6276 42291 6282 42343
rect 6650 42291 6656 42343
rect 6708 42291 6714 42343
rect 7050 42320 7078 42663
rect 7322 42320 7350 42663
rect 5665 42156 5671 42208
rect 5723 42156 5729 42208
rect 5555 42066 5561 42118
rect 5613 42066 5619 42118
rect 5665 41954 5671 42006
rect 5723 41954 5729 42006
rect 5802 41969 5848 42291
rect 5793 41917 5799 41969
rect 5851 41917 5857 41969
rect 5665 41792 5671 41844
rect 5723 41792 5729 41844
rect 5555 41680 5561 41732
rect 5613 41680 5619 41732
rect 5665 41590 5671 41642
rect 5723 41590 5729 41642
rect 5802 41553 5848 41917
rect 6226 41911 6274 42291
rect 6658 41911 6706 42291
rect 7032 42268 7038 42320
rect 7090 42268 7096 42320
rect 7304 42268 7310 42320
rect 7362 42268 7368 42320
rect 7050 41925 7078 42268
rect 7322 41925 7350 42268
rect 6218 41859 6224 41911
rect 6276 41859 6282 41911
rect 6650 41859 6656 41911
rect 6708 41859 6714 41911
rect 7032 41873 7038 41925
rect 7090 41873 7096 41925
rect 7304 41873 7310 41925
rect 7362 41873 7368 41925
rect 6226 41553 6274 41859
rect 6658 41553 6706 41859
rect 5793 41501 5799 41553
rect 5851 41501 5857 41553
rect 6218 41501 6224 41553
rect 6276 41501 6282 41553
rect 6650 41501 6656 41553
rect 6708 41501 6714 41553
rect 7050 41530 7078 41873
rect 7322 41530 7350 41873
rect 5665 41366 5671 41418
rect 5723 41366 5729 41418
rect 5555 41276 5561 41328
rect 5613 41276 5619 41328
rect 5665 41164 5671 41216
rect 5723 41164 5729 41216
rect 5802 41179 5848 41501
rect 5793 41127 5799 41179
rect 5851 41127 5857 41179
rect 5665 41002 5671 41054
rect 5723 41002 5729 41054
rect 5555 40890 5561 40942
rect 5613 40890 5619 40942
rect 5665 40800 5671 40852
rect 5723 40800 5729 40852
rect 5802 40763 5848 41127
rect 6226 41121 6274 41501
rect 6658 41121 6706 41501
rect 7032 41478 7038 41530
rect 7090 41478 7096 41530
rect 7304 41478 7310 41530
rect 7362 41478 7368 41530
rect 7050 41135 7078 41478
rect 7322 41135 7350 41478
rect 6218 41069 6224 41121
rect 6276 41069 6282 41121
rect 6650 41069 6656 41121
rect 6708 41069 6714 41121
rect 7032 41083 7038 41135
rect 7090 41083 7096 41135
rect 7304 41083 7310 41135
rect 7362 41083 7368 41135
rect 6226 40763 6274 41069
rect 6658 40763 6706 41069
rect 5793 40711 5799 40763
rect 5851 40711 5857 40763
rect 6218 40711 6224 40763
rect 6276 40711 6282 40763
rect 6650 40711 6656 40763
rect 6708 40711 6714 40763
rect 7050 40740 7078 41083
rect 7322 40740 7350 41083
rect 5665 40576 5671 40628
rect 5723 40576 5729 40628
rect 5555 40486 5561 40538
rect 5613 40486 5619 40538
rect 5665 40374 5671 40426
rect 5723 40374 5729 40426
rect 5802 40389 5848 40711
rect 5793 40337 5799 40389
rect 5851 40337 5857 40389
rect 5665 40212 5671 40264
rect 5723 40212 5729 40264
rect 5555 40100 5561 40152
rect 5613 40100 5619 40152
rect 5665 40010 5671 40062
rect 5723 40010 5729 40062
rect 5802 39973 5848 40337
rect 6226 40331 6274 40711
rect 6658 40331 6706 40711
rect 7032 40688 7038 40740
rect 7090 40688 7096 40740
rect 7304 40688 7310 40740
rect 7362 40688 7368 40740
rect 7050 40345 7078 40688
rect 7322 40345 7350 40688
rect 6218 40279 6224 40331
rect 6276 40279 6282 40331
rect 6650 40279 6656 40331
rect 6708 40279 6714 40331
rect 7032 40293 7038 40345
rect 7090 40293 7096 40345
rect 7304 40293 7310 40345
rect 7362 40293 7368 40345
rect 6226 39973 6274 40279
rect 6658 39973 6706 40279
rect 5793 39921 5799 39973
rect 5851 39921 5857 39973
rect 6218 39921 6224 39973
rect 6276 39921 6282 39973
rect 6650 39921 6656 39973
rect 6708 39921 6714 39973
rect 7050 39950 7078 40293
rect 7322 39950 7350 40293
rect 5665 39786 5671 39838
rect 5723 39786 5729 39838
rect 5555 39696 5561 39748
rect 5613 39696 5619 39748
rect 5665 39584 5671 39636
rect 5723 39584 5729 39636
rect 5802 39599 5848 39921
rect 5793 39547 5799 39599
rect 5851 39547 5857 39599
rect 5665 39422 5671 39474
rect 5723 39422 5729 39474
rect 5555 39310 5561 39362
rect 5613 39310 5619 39362
rect 5665 39220 5671 39272
rect 5723 39220 5729 39272
rect 5802 39183 5848 39547
rect 6226 39541 6274 39921
rect 6658 39541 6706 39921
rect 7032 39898 7038 39950
rect 7090 39898 7096 39950
rect 7304 39898 7310 39950
rect 7362 39898 7368 39950
rect 7050 39555 7078 39898
rect 7322 39555 7350 39898
rect 6218 39489 6224 39541
rect 6276 39489 6282 39541
rect 6650 39489 6656 39541
rect 6708 39489 6714 39541
rect 7032 39503 7038 39555
rect 7090 39503 7096 39555
rect 7304 39503 7310 39555
rect 7362 39503 7368 39555
rect 6226 39183 6274 39489
rect 6658 39183 6706 39489
rect 5793 39131 5799 39183
rect 5851 39131 5857 39183
rect 6218 39131 6224 39183
rect 6276 39131 6282 39183
rect 6650 39131 6656 39183
rect 6708 39131 6714 39183
rect 7050 39160 7078 39503
rect 7322 39160 7350 39503
rect 5665 38996 5671 39048
rect 5723 38996 5729 39048
rect 5555 38906 5561 38958
rect 5613 38906 5619 38958
rect 5665 38794 5671 38846
rect 5723 38794 5729 38846
rect 5802 38809 5848 39131
rect 5793 38757 5799 38809
rect 5851 38757 5857 38809
rect 5665 38632 5671 38684
rect 5723 38632 5729 38684
rect 5555 38520 5561 38572
rect 5613 38520 5619 38572
rect 5665 38430 5671 38482
rect 5723 38430 5729 38482
rect 5802 38393 5848 38757
rect 6226 38751 6274 39131
rect 6658 38751 6706 39131
rect 7032 39108 7038 39160
rect 7090 39108 7096 39160
rect 7304 39108 7310 39160
rect 7362 39108 7368 39160
rect 7050 38765 7078 39108
rect 7322 38765 7350 39108
rect 6218 38699 6224 38751
rect 6276 38699 6282 38751
rect 6650 38699 6656 38751
rect 6708 38699 6714 38751
rect 7032 38713 7038 38765
rect 7090 38713 7096 38765
rect 7304 38713 7310 38765
rect 7362 38713 7368 38765
rect 6226 38393 6274 38699
rect 6658 38393 6706 38699
rect 5793 38341 5799 38393
rect 5851 38341 5857 38393
rect 6218 38341 6224 38393
rect 6276 38341 6282 38393
rect 6650 38341 6656 38393
rect 6708 38341 6714 38393
rect 7050 38370 7078 38713
rect 7322 38370 7350 38713
rect 5665 38206 5671 38258
rect 5723 38206 5729 38258
rect 5555 38116 5561 38168
rect 5613 38116 5619 38168
rect 5665 38004 5671 38056
rect 5723 38004 5729 38056
rect 5802 38019 5848 38341
rect 5793 37967 5799 38019
rect 5851 37967 5857 38019
rect 5665 37842 5671 37894
rect 5723 37842 5729 37894
rect 5555 37730 5561 37782
rect 5613 37730 5619 37782
rect 5665 37640 5671 37692
rect 5723 37640 5729 37692
rect 5802 37603 5848 37967
rect 6226 37961 6274 38341
rect 6658 37961 6706 38341
rect 7032 38318 7038 38370
rect 7090 38318 7096 38370
rect 7304 38318 7310 38370
rect 7362 38318 7368 38370
rect 7050 37975 7078 38318
rect 7322 37975 7350 38318
rect 6218 37909 6224 37961
rect 6276 37909 6282 37961
rect 6650 37909 6656 37961
rect 6708 37909 6714 37961
rect 7032 37923 7038 37975
rect 7090 37923 7096 37975
rect 7304 37923 7310 37975
rect 7362 37923 7368 37975
rect 6226 37603 6274 37909
rect 6658 37603 6706 37909
rect 5793 37551 5799 37603
rect 5851 37551 5857 37603
rect 6218 37551 6224 37603
rect 6276 37551 6282 37603
rect 6650 37551 6656 37603
rect 6708 37551 6714 37603
rect 7050 37580 7078 37923
rect 7322 37580 7350 37923
rect 5665 37416 5671 37468
rect 5723 37416 5729 37468
rect 5555 37326 5561 37378
rect 5613 37326 5619 37378
rect 5665 37214 5671 37266
rect 5723 37214 5729 37266
rect 5802 37229 5848 37551
rect 5793 37177 5799 37229
rect 5851 37177 5857 37229
rect 5665 37052 5671 37104
rect 5723 37052 5729 37104
rect 5555 36940 5561 36992
rect 5613 36940 5619 36992
rect 5665 36850 5671 36902
rect 5723 36850 5729 36902
rect 5802 36813 5848 37177
rect 6226 37171 6274 37551
rect 6658 37171 6706 37551
rect 7032 37528 7038 37580
rect 7090 37528 7096 37580
rect 7304 37528 7310 37580
rect 7362 37528 7368 37580
rect 7050 37185 7078 37528
rect 7322 37185 7350 37528
rect 6218 37119 6224 37171
rect 6276 37119 6282 37171
rect 6650 37119 6656 37171
rect 6708 37119 6714 37171
rect 7032 37133 7038 37185
rect 7090 37133 7096 37185
rect 7304 37133 7310 37185
rect 7362 37133 7368 37185
rect 6226 36813 6274 37119
rect 6658 36813 6706 37119
rect 5793 36761 5799 36813
rect 5851 36761 5857 36813
rect 6218 36761 6224 36813
rect 6276 36761 6282 36813
rect 6650 36761 6656 36813
rect 6708 36761 6714 36813
rect 7050 36790 7078 37133
rect 7322 36790 7350 37133
rect 5665 36626 5671 36678
rect 5723 36626 5729 36678
rect 5555 36536 5561 36588
rect 5613 36536 5619 36588
rect 5665 36424 5671 36476
rect 5723 36424 5729 36476
rect 5802 36439 5848 36761
rect 5793 36387 5799 36439
rect 5851 36387 5857 36439
rect 5665 36262 5671 36314
rect 5723 36262 5729 36314
rect 5555 36150 5561 36202
rect 5613 36150 5619 36202
rect 5665 36060 5671 36112
rect 5723 36060 5729 36112
rect 5802 36023 5848 36387
rect 6226 36381 6274 36761
rect 6658 36381 6706 36761
rect 7032 36738 7038 36790
rect 7090 36738 7096 36790
rect 7304 36738 7310 36790
rect 7362 36738 7368 36790
rect 7050 36395 7078 36738
rect 7322 36395 7350 36738
rect 6218 36329 6224 36381
rect 6276 36329 6282 36381
rect 6650 36329 6656 36381
rect 6708 36329 6714 36381
rect 7032 36343 7038 36395
rect 7090 36343 7096 36395
rect 7304 36343 7310 36395
rect 7362 36343 7368 36395
rect 6226 36023 6274 36329
rect 6658 36023 6706 36329
rect 5793 35971 5799 36023
rect 5851 35971 5857 36023
rect 6218 35971 6224 36023
rect 6276 35971 6282 36023
rect 6650 35971 6656 36023
rect 6708 35971 6714 36023
rect 7050 36000 7078 36343
rect 7322 36000 7350 36343
rect 5665 35836 5671 35888
rect 5723 35836 5729 35888
rect 5555 35746 5561 35798
rect 5613 35746 5619 35798
rect 5665 35634 5671 35686
rect 5723 35634 5729 35686
rect 5802 35649 5848 35971
rect 5793 35597 5799 35649
rect 5851 35597 5857 35649
rect 5665 35472 5671 35524
rect 5723 35472 5729 35524
rect 5555 35360 5561 35412
rect 5613 35360 5619 35412
rect 5665 35270 5671 35322
rect 5723 35270 5729 35322
rect 5802 35233 5848 35597
rect 6226 35591 6274 35971
rect 6658 35591 6706 35971
rect 7032 35948 7038 36000
rect 7090 35948 7096 36000
rect 7304 35948 7310 36000
rect 7362 35948 7368 36000
rect 7050 35605 7078 35948
rect 7322 35605 7350 35948
rect 6218 35539 6224 35591
rect 6276 35539 6282 35591
rect 6650 35539 6656 35591
rect 6708 35539 6714 35591
rect 7032 35553 7038 35605
rect 7090 35553 7096 35605
rect 7304 35553 7310 35605
rect 7362 35553 7368 35605
rect 6226 35233 6274 35539
rect 6658 35233 6706 35539
rect 5793 35181 5799 35233
rect 5851 35181 5857 35233
rect 6218 35181 6224 35233
rect 6276 35181 6282 35233
rect 6650 35181 6656 35233
rect 6708 35181 6714 35233
rect 7050 35210 7078 35553
rect 7322 35210 7350 35553
rect 5665 35046 5671 35098
rect 5723 35046 5729 35098
rect 5555 34956 5561 35008
rect 5613 34956 5619 35008
rect 5665 34844 5671 34896
rect 5723 34844 5729 34896
rect 5802 34859 5848 35181
rect 5793 34807 5799 34859
rect 5851 34807 5857 34859
rect 5665 34682 5671 34734
rect 5723 34682 5729 34734
rect 5555 34570 5561 34622
rect 5613 34570 5619 34622
rect 5665 34480 5671 34532
rect 5723 34480 5729 34532
rect 5802 34443 5848 34807
rect 6226 34801 6274 35181
rect 6658 34801 6706 35181
rect 7032 35158 7038 35210
rect 7090 35158 7096 35210
rect 7304 35158 7310 35210
rect 7362 35158 7368 35210
rect 7050 34815 7078 35158
rect 7322 34815 7350 35158
rect 6218 34749 6224 34801
rect 6276 34749 6282 34801
rect 6650 34749 6656 34801
rect 6708 34749 6714 34801
rect 7032 34763 7038 34815
rect 7090 34763 7096 34815
rect 7304 34763 7310 34815
rect 7362 34763 7368 34815
rect 6226 34443 6274 34749
rect 6658 34443 6706 34749
rect 5793 34391 5799 34443
rect 5851 34391 5857 34443
rect 6218 34391 6224 34443
rect 6276 34391 6282 34443
rect 6650 34391 6656 34443
rect 6708 34391 6714 34443
rect 7050 34420 7078 34763
rect 7322 34420 7350 34763
rect 5665 34256 5671 34308
rect 5723 34256 5729 34308
rect 5555 34166 5561 34218
rect 5613 34166 5619 34218
rect 5665 34054 5671 34106
rect 5723 34054 5729 34106
rect 5802 34069 5848 34391
rect 5793 34017 5799 34069
rect 5851 34017 5857 34069
rect 5665 33892 5671 33944
rect 5723 33892 5729 33944
rect 5555 33780 5561 33832
rect 5613 33780 5619 33832
rect 5665 33690 5671 33742
rect 5723 33690 5729 33742
rect 5802 33653 5848 34017
rect 6226 34011 6274 34391
rect 6658 34011 6706 34391
rect 7032 34368 7038 34420
rect 7090 34368 7096 34420
rect 7304 34368 7310 34420
rect 7362 34368 7368 34420
rect 7050 34025 7078 34368
rect 7322 34025 7350 34368
rect 6218 33959 6224 34011
rect 6276 33959 6282 34011
rect 6650 33959 6656 34011
rect 6708 33959 6714 34011
rect 7032 33973 7038 34025
rect 7090 33973 7096 34025
rect 7304 33973 7310 34025
rect 7362 33973 7368 34025
rect 6226 33653 6274 33959
rect 6658 33653 6706 33959
rect 5793 33601 5799 33653
rect 5851 33601 5857 33653
rect 6218 33601 6224 33653
rect 6276 33601 6282 33653
rect 6650 33601 6656 33653
rect 6708 33601 6714 33653
rect 7050 33630 7078 33973
rect 7322 33630 7350 33973
rect 5665 33466 5671 33518
rect 5723 33466 5729 33518
rect 5555 33376 5561 33428
rect 5613 33376 5619 33428
rect 5665 33264 5671 33316
rect 5723 33264 5729 33316
rect 5802 33279 5848 33601
rect 5793 33227 5799 33279
rect 5851 33227 5857 33279
rect 5665 33102 5671 33154
rect 5723 33102 5729 33154
rect 5555 32990 5561 33042
rect 5613 32990 5619 33042
rect 5665 32900 5671 32952
rect 5723 32900 5729 32952
rect 5802 32863 5848 33227
rect 6226 33221 6274 33601
rect 6658 33221 6706 33601
rect 7032 33578 7038 33630
rect 7090 33578 7096 33630
rect 7304 33578 7310 33630
rect 7362 33578 7368 33630
rect 7050 33235 7078 33578
rect 7322 33235 7350 33578
rect 6218 33169 6224 33221
rect 6276 33169 6282 33221
rect 6650 33169 6656 33221
rect 6708 33169 6714 33221
rect 7032 33183 7038 33235
rect 7090 33183 7096 33235
rect 7304 33183 7310 33235
rect 7362 33183 7368 33235
rect 6226 32863 6274 33169
rect 6658 32863 6706 33169
rect 5793 32811 5799 32863
rect 5851 32811 5857 32863
rect 6218 32811 6224 32863
rect 6276 32811 6282 32863
rect 6650 32811 6656 32863
rect 6708 32811 6714 32863
rect 7050 32840 7078 33183
rect 7322 32840 7350 33183
rect 5665 32676 5671 32728
rect 5723 32676 5729 32728
rect 5555 32586 5561 32638
rect 5613 32586 5619 32638
rect 5665 32474 5671 32526
rect 5723 32474 5729 32526
rect 5802 32489 5848 32811
rect 5793 32437 5799 32489
rect 5851 32437 5857 32489
rect 5665 32312 5671 32364
rect 5723 32312 5729 32364
rect 5555 32200 5561 32252
rect 5613 32200 5619 32252
rect 5665 32110 5671 32162
rect 5723 32110 5729 32162
rect 5802 32073 5848 32437
rect 6226 32431 6274 32811
rect 6658 32431 6706 32811
rect 7032 32788 7038 32840
rect 7090 32788 7096 32840
rect 7304 32788 7310 32840
rect 7362 32788 7368 32840
rect 7050 32445 7078 32788
rect 7322 32445 7350 32788
rect 6218 32379 6224 32431
rect 6276 32379 6282 32431
rect 6650 32379 6656 32431
rect 6708 32379 6714 32431
rect 7032 32393 7038 32445
rect 7090 32393 7096 32445
rect 7304 32393 7310 32445
rect 7362 32393 7368 32445
rect 6226 32073 6274 32379
rect 6658 32073 6706 32379
rect 5793 32021 5799 32073
rect 5851 32021 5857 32073
rect 6218 32021 6224 32073
rect 6276 32021 6282 32073
rect 6650 32021 6656 32073
rect 6708 32021 6714 32073
rect 7050 32050 7078 32393
rect 7322 32050 7350 32393
rect 5665 31886 5671 31938
rect 5723 31886 5729 31938
rect 5555 31796 5561 31848
rect 5613 31796 5619 31848
rect 5665 31684 5671 31736
rect 5723 31684 5729 31736
rect 5802 31699 5848 32021
rect 5793 31647 5799 31699
rect 5851 31647 5857 31699
rect 5665 31522 5671 31574
rect 5723 31522 5729 31574
rect 5555 31410 5561 31462
rect 5613 31410 5619 31462
rect 5665 31320 5671 31372
rect 5723 31320 5729 31372
rect 5802 31283 5848 31647
rect 6226 31641 6274 32021
rect 6658 31641 6706 32021
rect 7032 31998 7038 32050
rect 7090 31998 7096 32050
rect 7304 31998 7310 32050
rect 7362 31998 7368 32050
rect 7050 31655 7078 31998
rect 7322 31655 7350 31998
rect 6218 31589 6224 31641
rect 6276 31589 6282 31641
rect 6650 31589 6656 31641
rect 6708 31589 6714 31641
rect 7032 31603 7038 31655
rect 7090 31603 7096 31655
rect 7304 31603 7310 31655
rect 7362 31603 7368 31655
rect 6226 31283 6274 31589
rect 6658 31283 6706 31589
rect 5793 31231 5799 31283
rect 5851 31231 5857 31283
rect 6218 31231 6224 31283
rect 6276 31231 6282 31283
rect 6650 31231 6656 31283
rect 6708 31231 6714 31283
rect 7050 31260 7078 31603
rect 7322 31260 7350 31603
rect 5665 31096 5671 31148
rect 5723 31096 5729 31148
rect 5555 31006 5561 31058
rect 5613 31006 5619 31058
rect 5665 30894 5671 30946
rect 5723 30894 5729 30946
rect 5802 30909 5848 31231
rect 5793 30857 5799 30909
rect 5851 30857 5857 30909
rect 5665 30732 5671 30784
rect 5723 30732 5729 30784
rect 5555 30620 5561 30672
rect 5613 30620 5619 30672
rect 5665 30530 5671 30582
rect 5723 30530 5729 30582
rect 5802 30493 5848 30857
rect 6226 30851 6274 31231
rect 6658 30851 6706 31231
rect 7032 31208 7038 31260
rect 7090 31208 7096 31260
rect 7304 31208 7310 31260
rect 7362 31208 7368 31260
rect 7050 30865 7078 31208
rect 7322 30865 7350 31208
rect 6218 30799 6224 30851
rect 6276 30799 6282 30851
rect 6650 30799 6656 30851
rect 6708 30799 6714 30851
rect 7032 30813 7038 30865
rect 7090 30813 7096 30865
rect 7304 30813 7310 30865
rect 7362 30813 7368 30865
rect 6226 30493 6274 30799
rect 6658 30493 6706 30799
rect 5793 30441 5799 30493
rect 5851 30441 5857 30493
rect 6218 30441 6224 30493
rect 6276 30441 6282 30493
rect 6650 30441 6656 30493
rect 6708 30441 6714 30493
rect 7050 30470 7078 30813
rect 7322 30470 7350 30813
rect 5665 30306 5671 30358
rect 5723 30306 5729 30358
rect 5555 30216 5561 30268
rect 5613 30216 5619 30268
rect 5665 30104 5671 30156
rect 5723 30104 5729 30156
rect 5802 30119 5848 30441
rect 5793 30067 5799 30119
rect 5851 30067 5857 30119
rect 5665 29942 5671 29994
rect 5723 29942 5729 29994
rect 5555 29830 5561 29882
rect 5613 29830 5619 29882
rect 5665 29740 5671 29792
rect 5723 29740 5729 29792
rect 5802 29703 5848 30067
rect 6226 30061 6274 30441
rect 6658 30061 6706 30441
rect 7032 30418 7038 30470
rect 7090 30418 7096 30470
rect 7304 30418 7310 30470
rect 7362 30418 7368 30470
rect 7050 30075 7078 30418
rect 7322 30075 7350 30418
rect 6218 30009 6224 30061
rect 6276 30009 6282 30061
rect 6650 30009 6656 30061
rect 6708 30009 6714 30061
rect 7032 30023 7038 30075
rect 7090 30023 7096 30075
rect 7304 30023 7310 30075
rect 7362 30023 7368 30075
rect 6226 29703 6274 30009
rect 6658 29703 6706 30009
rect 5793 29651 5799 29703
rect 5851 29651 5857 29703
rect 6218 29651 6224 29703
rect 6276 29651 6282 29703
rect 6650 29651 6656 29703
rect 6708 29651 6714 29703
rect 7050 29680 7078 30023
rect 7322 29680 7350 30023
rect 5665 29516 5671 29568
rect 5723 29516 5729 29568
rect 5555 29426 5561 29478
rect 5613 29426 5619 29478
rect 5665 29314 5671 29366
rect 5723 29314 5729 29366
rect 5802 29329 5848 29651
rect 5793 29277 5799 29329
rect 5851 29277 5857 29329
rect 5665 29152 5671 29204
rect 5723 29152 5729 29204
rect 5555 29040 5561 29092
rect 5613 29040 5619 29092
rect 5665 28950 5671 29002
rect 5723 28950 5729 29002
rect 5802 28913 5848 29277
rect 6226 29271 6274 29651
rect 6658 29271 6706 29651
rect 7032 29628 7038 29680
rect 7090 29628 7096 29680
rect 7304 29628 7310 29680
rect 7362 29628 7368 29680
rect 7050 29285 7078 29628
rect 7322 29285 7350 29628
rect 6218 29219 6224 29271
rect 6276 29219 6282 29271
rect 6650 29219 6656 29271
rect 6708 29219 6714 29271
rect 7032 29233 7038 29285
rect 7090 29233 7096 29285
rect 7304 29233 7310 29285
rect 7362 29233 7368 29285
rect 6226 28913 6274 29219
rect 6658 28913 6706 29219
rect 5793 28861 5799 28913
rect 5851 28861 5857 28913
rect 6218 28861 6224 28913
rect 6276 28861 6282 28913
rect 6650 28861 6656 28913
rect 6708 28861 6714 28913
rect 7050 28890 7078 29233
rect 7322 28890 7350 29233
rect 5665 28726 5671 28778
rect 5723 28726 5729 28778
rect 5555 28636 5561 28688
rect 5613 28636 5619 28688
rect 5665 28524 5671 28576
rect 5723 28524 5729 28576
rect 5802 28539 5848 28861
rect 5793 28487 5799 28539
rect 5851 28487 5857 28539
rect 5665 28362 5671 28414
rect 5723 28362 5729 28414
rect 5555 28250 5561 28302
rect 5613 28250 5619 28302
rect 5665 28160 5671 28212
rect 5723 28160 5729 28212
rect 5802 28123 5848 28487
rect 6226 28481 6274 28861
rect 6658 28481 6706 28861
rect 7032 28838 7038 28890
rect 7090 28838 7096 28890
rect 7304 28838 7310 28890
rect 7362 28838 7368 28890
rect 7050 28495 7078 28838
rect 7322 28495 7350 28838
rect 6218 28429 6224 28481
rect 6276 28429 6282 28481
rect 6650 28429 6656 28481
rect 6708 28429 6714 28481
rect 7032 28443 7038 28495
rect 7090 28443 7096 28495
rect 7304 28443 7310 28495
rect 7362 28443 7368 28495
rect 6226 28123 6274 28429
rect 6658 28123 6706 28429
rect 5793 28071 5799 28123
rect 5851 28071 5857 28123
rect 6218 28071 6224 28123
rect 6276 28071 6282 28123
rect 6650 28071 6656 28123
rect 6708 28071 6714 28123
rect 7050 28100 7078 28443
rect 7322 28100 7350 28443
rect 5665 27936 5671 27988
rect 5723 27936 5729 27988
rect 5555 27846 5561 27898
rect 5613 27846 5619 27898
rect 5665 27734 5671 27786
rect 5723 27734 5729 27786
rect 5802 27749 5848 28071
rect 5793 27697 5799 27749
rect 5851 27697 5857 27749
rect 5665 27572 5671 27624
rect 5723 27572 5729 27624
rect 5555 27460 5561 27512
rect 5613 27460 5619 27512
rect 5665 27370 5671 27422
rect 5723 27370 5729 27422
rect 5802 27333 5848 27697
rect 6226 27691 6274 28071
rect 6658 27691 6706 28071
rect 7032 28048 7038 28100
rect 7090 28048 7096 28100
rect 7304 28048 7310 28100
rect 7362 28048 7368 28100
rect 7050 27705 7078 28048
rect 7322 27705 7350 28048
rect 6218 27639 6224 27691
rect 6276 27639 6282 27691
rect 6650 27639 6656 27691
rect 6708 27639 6714 27691
rect 7032 27653 7038 27705
rect 7090 27653 7096 27705
rect 7304 27653 7310 27705
rect 7362 27653 7368 27705
rect 6226 27333 6274 27639
rect 6658 27333 6706 27639
rect 5793 27281 5799 27333
rect 5851 27281 5857 27333
rect 6218 27281 6224 27333
rect 6276 27281 6282 27333
rect 6650 27281 6656 27333
rect 6708 27281 6714 27333
rect 7050 27310 7078 27653
rect 7322 27310 7350 27653
rect 5665 27146 5671 27198
rect 5723 27146 5729 27198
rect 5555 27056 5561 27108
rect 5613 27056 5619 27108
rect 5665 26944 5671 26996
rect 5723 26944 5729 26996
rect 5802 26959 5848 27281
rect 5793 26907 5799 26959
rect 5851 26907 5857 26959
rect 5665 26782 5671 26834
rect 5723 26782 5729 26834
rect 5555 26670 5561 26722
rect 5613 26670 5619 26722
rect 5665 26580 5671 26632
rect 5723 26580 5729 26632
rect 5802 26543 5848 26907
rect 6226 26901 6274 27281
rect 6658 26901 6706 27281
rect 7032 27258 7038 27310
rect 7090 27258 7096 27310
rect 7304 27258 7310 27310
rect 7362 27258 7368 27310
rect 7050 26915 7078 27258
rect 7322 26915 7350 27258
rect 6218 26849 6224 26901
rect 6276 26849 6282 26901
rect 6650 26849 6656 26901
rect 6708 26849 6714 26901
rect 7032 26863 7038 26915
rect 7090 26863 7096 26915
rect 7304 26863 7310 26915
rect 7362 26863 7368 26915
rect 6226 26543 6274 26849
rect 6658 26543 6706 26849
rect 5793 26491 5799 26543
rect 5851 26491 5857 26543
rect 6218 26491 6224 26543
rect 6276 26491 6282 26543
rect 6650 26491 6656 26543
rect 6708 26491 6714 26543
rect 7050 26520 7078 26863
rect 7322 26520 7350 26863
rect 5665 26356 5671 26408
rect 5723 26356 5729 26408
rect 5555 26266 5561 26318
rect 5613 26266 5619 26318
rect 5665 26154 5671 26206
rect 5723 26154 5729 26206
rect 5802 26169 5848 26491
rect 5793 26117 5799 26169
rect 5851 26117 5857 26169
rect 5665 25992 5671 26044
rect 5723 25992 5729 26044
rect 5555 25880 5561 25932
rect 5613 25880 5619 25932
rect 5665 25790 5671 25842
rect 5723 25790 5729 25842
rect 5802 25753 5848 26117
rect 6226 26111 6274 26491
rect 6658 26111 6706 26491
rect 7032 26468 7038 26520
rect 7090 26468 7096 26520
rect 7304 26468 7310 26520
rect 7362 26468 7368 26520
rect 7050 26125 7078 26468
rect 7322 26125 7350 26468
rect 6218 26059 6224 26111
rect 6276 26059 6282 26111
rect 6650 26059 6656 26111
rect 6708 26059 6714 26111
rect 7032 26073 7038 26125
rect 7090 26073 7096 26125
rect 7304 26073 7310 26125
rect 7362 26073 7368 26125
rect 6226 25753 6274 26059
rect 6658 25753 6706 26059
rect 5793 25701 5799 25753
rect 5851 25701 5857 25753
rect 6218 25701 6224 25753
rect 6276 25701 6282 25753
rect 6650 25701 6656 25753
rect 6708 25701 6714 25753
rect 7050 25730 7078 26073
rect 7322 25730 7350 26073
rect 5665 25566 5671 25618
rect 5723 25566 5729 25618
rect 5555 25476 5561 25528
rect 5613 25476 5619 25528
rect 5665 25364 5671 25416
rect 5723 25364 5729 25416
rect 5802 25379 5848 25701
rect 5793 25327 5799 25379
rect 5851 25327 5857 25379
rect 5665 25202 5671 25254
rect 5723 25202 5729 25254
rect 5555 25090 5561 25142
rect 5613 25090 5619 25142
rect 5665 25000 5671 25052
rect 5723 25000 5729 25052
rect 5802 24963 5848 25327
rect 6226 25321 6274 25701
rect 6658 25321 6706 25701
rect 7032 25678 7038 25730
rect 7090 25678 7096 25730
rect 7304 25678 7310 25730
rect 7362 25678 7368 25730
rect 7050 25335 7078 25678
rect 7322 25335 7350 25678
rect 6218 25269 6224 25321
rect 6276 25269 6282 25321
rect 6650 25269 6656 25321
rect 6708 25269 6714 25321
rect 7032 25283 7038 25335
rect 7090 25283 7096 25335
rect 7304 25283 7310 25335
rect 7362 25283 7368 25335
rect 6226 24963 6274 25269
rect 6658 24963 6706 25269
rect 5793 24911 5799 24963
rect 5851 24911 5857 24963
rect 6218 24911 6224 24963
rect 6276 24911 6282 24963
rect 6650 24911 6656 24963
rect 6708 24911 6714 24963
rect 7050 24940 7078 25283
rect 7322 24940 7350 25283
rect 5665 24776 5671 24828
rect 5723 24776 5729 24828
rect 5555 24686 5561 24738
rect 5613 24686 5619 24738
rect 5665 24574 5671 24626
rect 5723 24574 5729 24626
rect 5802 24589 5848 24911
rect 5793 24537 5799 24589
rect 5851 24537 5857 24589
rect 5665 24412 5671 24464
rect 5723 24412 5729 24464
rect 5555 24300 5561 24352
rect 5613 24300 5619 24352
rect 5665 24210 5671 24262
rect 5723 24210 5729 24262
rect 5802 24173 5848 24537
rect 6226 24531 6274 24911
rect 6658 24531 6706 24911
rect 7032 24888 7038 24940
rect 7090 24888 7096 24940
rect 7304 24888 7310 24940
rect 7362 24888 7368 24940
rect 7050 24545 7078 24888
rect 7322 24545 7350 24888
rect 6218 24479 6224 24531
rect 6276 24479 6282 24531
rect 6650 24479 6656 24531
rect 6708 24479 6714 24531
rect 7032 24493 7038 24545
rect 7090 24493 7096 24545
rect 7304 24493 7310 24545
rect 7362 24493 7368 24545
rect 6226 24173 6274 24479
rect 6658 24173 6706 24479
rect 5793 24121 5799 24173
rect 5851 24121 5857 24173
rect 6218 24121 6224 24173
rect 6276 24121 6282 24173
rect 6650 24121 6656 24173
rect 6708 24121 6714 24173
rect 7050 24150 7078 24493
rect 7322 24150 7350 24493
rect 5665 23986 5671 24038
rect 5723 23986 5729 24038
rect 5555 23896 5561 23948
rect 5613 23896 5619 23948
rect 5665 23784 5671 23836
rect 5723 23784 5729 23836
rect 5802 23799 5848 24121
rect 5793 23747 5799 23799
rect 5851 23747 5857 23799
rect 5665 23622 5671 23674
rect 5723 23622 5729 23674
rect 5555 23510 5561 23562
rect 5613 23510 5619 23562
rect 5665 23420 5671 23472
rect 5723 23420 5729 23472
rect 5802 23383 5848 23747
rect 6226 23741 6274 24121
rect 6658 23741 6706 24121
rect 7032 24098 7038 24150
rect 7090 24098 7096 24150
rect 7304 24098 7310 24150
rect 7362 24098 7368 24150
rect 7050 23755 7078 24098
rect 7322 23755 7350 24098
rect 6218 23689 6224 23741
rect 6276 23689 6282 23741
rect 6650 23689 6656 23741
rect 6708 23689 6714 23741
rect 7032 23703 7038 23755
rect 7090 23703 7096 23755
rect 7304 23703 7310 23755
rect 7362 23703 7368 23755
rect 6226 23383 6274 23689
rect 6658 23383 6706 23689
rect 5793 23331 5799 23383
rect 5851 23331 5857 23383
rect 6218 23331 6224 23383
rect 6276 23331 6282 23383
rect 6650 23331 6656 23383
rect 6708 23331 6714 23383
rect 7050 23360 7078 23703
rect 7322 23360 7350 23703
rect 5665 23196 5671 23248
rect 5723 23196 5729 23248
rect 5555 23106 5561 23158
rect 5613 23106 5619 23158
rect 5665 22994 5671 23046
rect 5723 22994 5729 23046
rect 5802 23009 5848 23331
rect 5793 22957 5799 23009
rect 5851 22957 5857 23009
rect 5665 22832 5671 22884
rect 5723 22832 5729 22884
rect 5555 22720 5561 22772
rect 5613 22720 5619 22772
rect 5665 22630 5671 22682
rect 5723 22630 5729 22682
rect 5802 22593 5848 22957
rect 6226 22951 6274 23331
rect 6658 22951 6706 23331
rect 7032 23308 7038 23360
rect 7090 23308 7096 23360
rect 7304 23308 7310 23360
rect 7362 23308 7368 23360
rect 7050 22965 7078 23308
rect 7322 22965 7350 23308
rect 6218 22899 6224 22951
rect 6276 22899 6282 22951
rect 6650 22899 6656 22951
rect 6708 22899 6714 22951
rect 7032 22913 7038 22965
rect 7090 22913 7096 22965
rect 7304 22913 7310 22965
rect 7362 22913 7368 22965
rect 6226 22593 6274 22899
rect 6658 22593 6706 22899
rect 5793 22541 5799 22593
rect 5851 22541 5857 22593
rect 6218 22541 6224 22593
rect 6276 22541 6282 22593
rect 6650 22541 6656 22593
rect 6708 22541 6714 22593
rect 7050 22570 7078 22913
rect 7322 22570 7350 22913
rect 5665 22406 5671 22458
rect 5723 22406 5729 22458
rect 5555 22316 5561 22368
rect 5613 22316 5619 22368
rect 5665 22204 5671 22256
rect 5723 22204 5729 22256
rect 5802 22219 5848 22541
rect 5793 22167 5799 22219
rect 5851 22167 5857 22219
rect 5665 22042 5671 22094
rect 5723 22042 5729 22094
rect 5555 21930 5561 21982
rect 5613 21930 5619 21982
rect 5665 21840 5671 21892
rect 5723 21840 5729 21892
rect 5802 21803 5848 22167
rect 6226 22161 6274 22541
rect 6658 22161 6706 22541
rect 7032 22518 7038 22570
rect 7090 22518 7096 22570
rect 7304 22518 7310 22570
rect 7362 22518 7368 22570
rect 7050 22175 7078 22518
rect 7322 22175 7350 22518
rect 6218 22109 6224 22161
rect 6276 22109 6282 22161
rect 6650 22109 6656 22161
rect 6708 22109 6714 22161
rect 7032 22123 7038 22175
rect 7090 22123 7096 22175
rect 7304 22123 7310 22175
rect 7362 22123 7368 22175
rect 6226 21803 6274 22109
rect 6658 21803 6706 22109
rect 5793 21751 5799 21803
rect 5851 21751 5857 21803
rect 6218 21751 6224 21803
rect 6276 21751 6282 21803
rect 6650 21751 6656 21803
rect 6708 21751 6714 21803
rect 7050 21780 7078 22123
rect 7322 21780 7350 22123
rect 5665 21616 5671 21668
rect 5723 21616 5729 21668
rect 5555 21526 5561 21578
rect 5613 21526 5619 21578
rect 5665 21414 5671 21466
rect 5723 21414 5729 21466
rect 5802 21429 5848 21751
rect 5793 21377 5799 21429
rect 5851 21377 5857 21429
rect 5665 21252 5671 21304
rect 5723 21252 5729 21304
rect 5555 21140 5561 21192
rect 5613 21140 5619 21192
rect 5665 21050 5671 21102
rect 5723 21050 5729 21102
rect 5802 21013 5848 21377
rect 6226 21371 6274 21751
rect 6658 21371 6706 21751
rect 7032 21728 7038 21780
rect 7090 21728 7096 21780
rect 7304 21728 7310 21780
rect 7362 21728 7368 21780
rect 7050 21385 7078 21728
rect 7322 21385 7350 21728
rect 6218 21319 6224 21371
rect 6276 21319 6282 21371
rect 6650 21319 6656 21371
rect 6708 21319 6714 21371
rect 7032 21333 7038 21385
rect 7090 21333 7096 21385
rect 7304 21333 7310 21385
rect 7362 21333 7368 21385
rect 6226 21013 6274 21319
rect 6658 21013 6706 21319
rect 5793 20961 5799 21013
rect 5851 20961 5857 21013
rect 6218 20961 6224 21013
rect 6276 20961 6282 21013
rect 6650 20961 6656 21013
rect 6708 20961 6714 21013
rect 7050 20990 7078 21333
rect 7322 20990 7350 21333
rect 5665 20826 5671 20878
rect 5723 20826 5729 20878
rect 5555 20736 5561 20788
rect 5613 20736 5619 20788
rect 5665 20624 5671 20676
rect 5723 20624 5729 20676
rect 5802 20639 5848 20961
rect 5793 20587 5799 20639
rect 5851 20587 5857 20639
rect 5665 20462 5671 20514
rect 5723 20462 5729 20514
rect 5555 20350 5561 20402
rect 5613 20350 5619 20402
rect 5665 20260 5671 20312
rect 5723 20260 5729 20312
rect 5802 20223 5848 20587
rect 6226 20581 6274 20961
rect 6658 20581 6706 20961
rect 7032 20938 7038 20990
rect 7090 20938 7096 20990
rect 7304 20938 7310 20990
rect 7362 20938 7368 20990
rect 7050 20595 7078 20938
rect 7322 20595 7350 20938
rect 6218 20529 6224 20581
rect 6276 20529 6282 20581
rect 6650 20529 6656 20581
rect 6708 20529 6714 20581
rect 7032 20543 7038 20595
rect 7090 20543 7096 20595
rect 7304 20543 7310 20595
rect 7362 20543 7368 20595
rect 6226 20223 6274 20529
rect 6658 20223 6706 20529
rect 5793 20171 5799 20223
rect 5851 20171 5857 20223
rect 6218 20171 6224 20223
rect 6276 20171 6282 20223
rect 6650 20171 6656 20223
rect 6708 20171 6714 20223
rect 7050 20200 7078 20543
rect 7322 20200 7350 20543
rect 5665 20036 5671 20088
rect 5723 20036 5729 20088
rect 5555 19946 5561 19998
rect 5613 19946 5619 19998
rect 5665 19834 5671 19886
rect 5723 19834 5729 19886
rect 5802 19849 5848 20171
rect 5793 19797 5799 19849
rect 5851 19797 5857 19849
rect 5665 19672 5671 19724
rect 5723 19672 5729 19724
rect 5555 19560 5561 19612
rect 5613 19560 5619 19612
rect 5665 19470 5671 19522
rect 5723 19470 5729 19522
rect 5802 19433 5848 19797
rect 6226 19791 6274 20171
rect 6658 19791 6706 20171
rect 7032 20148 7038 20200
rect 7090 20148 7096 20200
rect 7304 20148 7310 20200
rect 7362 20148 7368 20200
rect 7050 19805 7078 20148
rect 7322 19805 7350 20148
rect 6218 19739 6224 19791
rect 6276 19739 6282 19791
rect 6650 19739 6656 19791
rect 6708 19739 6714 19791
rect 7032 19753 7038 19805
rect 7090 19753 7096 19805
rect 7304 19753 7310 19805
rect 7362 19753 7368 19805
rect 6226 19433 6274 19739
rect 6658 19433 6706 19739
rect 5793 19381 5799 19433
rect 5851 19381 5857 19433
rect 6218 19381 6224 19433
rect 6276 19381 6282 19433
rect 6650 19381 6656 19433
rect 6708 19381 6714 19433
rect 7050 19410 7078 19753
rect 7322 19410 7350 19753
rect 5665 19246 5671 19298
rect 5723 19246 5729 19298
rect 5555 19156 5561 19208
rect 5613 19156 5619 19208
rect 5665 19044 5671 19096
rect 5723 19044 5729 19096
rect 5802 19059 5848 19381
rect 5793 19007 5799 19059
rect 5851 19007 5857 19059
rect 5665 18882 5671 18934
rect 5723 18882 5729 18934
rect 5555 18770 5561 18822
rect 5613 18770 5619 18822
rect 5665 18680 5671 18732
rect 5723 18680 5729 18732
rect 5802 18643 5848 19007
rect 6226 19001 6274 19381
rect 6658 19001 6706 19381
rect 7032 19358 7038 19410
rect 7090 19358 7096 19410
rect 7304 19358 7310 19410
rect 7362 19358 7368 19410
rect 7050 19015 7078 19358
rect 7322 19015 7350 19358
rect 6218 18949 6224 19001
rect 6276 18949 6282 19001
rect 6650 18949 6656 19001
rect 6708 18949 6714 19001
rect 7032 18963 7038 19015
rect 7090 18963 7096 19015
rect 7304 18963 7310 19015
rect 7362 18963 7368 19015
rect 6226 18643 6274 18949
rect 6658 18643 6706 18949
rect 5793 18591 5799 18643
rect 5851 18591 5857 18643
rect 6218 18591 6224 18643
rect 6276 18591 6282 18643
rect 6650 18591 6656 18643
rect 6708 18591 6714 18643
rect 7050 18620 7078 18963
rect 7322 18620 7350 18963
rect 5665 18456 5671 18508
rect 5723 18456 5729 18508
rect 5555 18366 5561 18418
rect 5613 18366 5619 18418
rect 5665 18254 5671 18306
rect 5723 18254 5729 18306
rect 5802 18269 5848 18591
rect 5793 18217 5799 18269
rect 5851 18217 5857 18269
rect 5665 18092 5671 18144
rect 5723 18092 5729 18144
rect 5555 17980 5561 18032
rect 5613 17980 5619 18032
rect 5665 17890 5671 17942
rect 5723 17890 5729 17942
rect 5802 17853 5848 18217
rect 6226 18211 6274 18591
rect 6658 18211 6706 18591
rect 7032 18568 7038 18620
rect 7090 18568 7096 18620
rect 7304 18568 7310 18620
rect 7362 18568 7368 18620
rect 7050 18225 7078 18568
rect 7322 18225 7350 18568
rect 6218 18159 6224 18211
rect 6276 18159 6282 18211
rect 6650 18159 6656 18211
rect 6708 18159 6714 18211
rect 7032 18173 7038 18225
rect 7090 18173 7096 18225
rect 7304 18173 7310 18225
rect 7362 18173 7368 18225
rect 6226 17853 6274 18159
rect 6658 17853 6706 18159
rect 5793 17801 5799 17853
rect 5851 17801 5857 17853
rect 6218 17801 6224 17853
rect 6276 17801 6282 17853
rect 6650 17801 6656 17853
rect 6708 17801 6714 17853
rect 7050 17830 7078 18173
rect 7322 17830 7350 18173
rect 5665 17666 5671 17718
rect 5723 17666 5729 17718
rect 5555 17576 5561 17628
rect 5613 17576 5619 17628
rect 5665 17464 5671 17516
rect 5723 17464 5729 17516
rect 5802 17479 5848 17801
rect 5793 17427 5799 17479
rect 5851 17427 5857 17479
rect 5665 17302 5671 17354
rect 5723 17302 5729 17354
rect 5555 17190 5561 17242
rect 5613 17190 5619 17242
rect 5665 17100 5671 17152
rect 5723 17100 5729 17152
rect 5802 17063 5848 17427
rect 6226 17421 6274 17801
rect 6658 17421 6706 17801
rect 7032 17778 7038 17830
rect 7090 17778 7096 17830
rect 7304 17778 7310 17830
rect 7362 17778 7368 17830
rect 7050 17435 7078 17778
rect 7322 17435 7350 17778
rect 6218 17369 6224 17421
rect 6276 17369 6282 17421
rect 6650 17369 6656 17421
rect 6708 17369 6714 17421
rect 7032 17383 7038 17435
rect 7090 17383 7096 17435
rect 7304 17383 7310 17435
rect 7362 17383 7368 17435
rect 6226 17063 6274 17369
rect 6658 17063 6706 17369
rect 5793 17011 5799 17063
rect 5851 17011 5857 17063
rect 6218 17011 6224 17063
rect 6276 17011 6282 17063
rect 6650 17011 6656 17063
rect 6708 17011 6714 17063
rect 7050 17040 7078 17383
rect 7322 17040 7350 17383
rect 5665 16876 5671 16928
rect 5723 16876 5729 16928
rect 5555 16786 5561 16838
rect 5613 16786 5619 16838
rect 5665 16674 5671 16726
rect 5723 16674 5729 16726
rect 5802 16689 5848 17011
rect 5793 16637 5799 16689
rect 5851 16637 5857 16689
rect 5665 16512 5671 16564
rect 5723 16512 5729 16564
rect 5555 16400 5561 16452
rect 5613 16400 5619 16452
rect 5665 16310 5671 16362
rect 5723 16310 5729 16362
rect 5802 16273 5848 16637
rect 6226 16631 6274 17011
rect 6658 16631 6706 17011
rect 7032 16988 7038 17040
rect 7090 16988 7096 17040
rect 7304 16988 7310 17040
rect 7362 16988 7368 17040
rect 7050 16645 7078 16988
rect 7322 16645 7350 16988
rect 6218 16579 6224 16631
rect 6276 16579 6282 16631
rect 6650 16579 6656 16631
rect 6708 16579 6714 16631
rect 7032 16593 7038 16645
rect 7090 16593 7096 16645
rect 7304 16593 7310 16645
rect 7362 16593 7368 16645
rect 6226 16273 6274 16579
rect 6658 16273 6706 16579
rect 5793 16221 5799 16273
rect 5851 16221 5857 16273
rect 6218 16221 6224 16273
rect 6276 16221 6282 16273
rect 6650 16221 6656 16273
rect 6708 16221 6714 16273
rect 7050 16250 7078 16593
rect 7322 16250 7350 16593
rect 5665 16086 5671 16138
rect 5723 16086 5729 16138
rect 5555 15996 5561 16048
rect 5613 15996 5619 16048
rect 5665 15884 5671 15936
rect 5723 15884 5729 15936
rect 5802 15899 5848 16221
rect 5793 15847 5799 15899
rect 5851 15847 5857 15899
rect 5665 15722 5671 15774
rect 5723 15722 5729 15774
rect 5555 15610 5561 15662
rect 5613 15610 5619 15662
rect 5665 15520 5671 15572
rect 5723 15520 5729 15572
rect 5802 15483 5848 15847
rect 6226 15841 6274 16221
rect 6658 15841 6706 16221
rect 7032 16198 7038 16250
rect 7090 16198 7096 16250
rect 7304 16198 7310 16250
rect 7362 16198 7368 16250
rect 7050 15855 7078 16198
rect 7322 15855 7350 16198
rect 6218 15789 6224 15841
rect 6276 15789 6282 15841
rect 6650 15789 6656 15841
rect 6708 15789 6714 15841
rect 7032 15803 7038 15855
rect 7090 15803 7096 15855
rect 7304 15803 7310 15855
rect 7362 15803 7368 15855
rect 6226 15483 6274 15789
rect 6658 15483 6706 15789
rect 5793 15431 5799 15483
rect 5851 15431 5857 15483
rect 6218 15431 6224 15483
rect 6276 15431 6282 15483
rect 6650 15431 6656 15483
rect 6708 15431 6714 15483
rect 7050 15460 7078 15803
rect 7322 15460 7350 15803
rect 5665 15296 5671 15348
rect 5723 15296 5729 15348
rect 5555 15206 5561 15258
rect 5613 15206 5619 15258
rect 5665 15094 5671 15146
rect 5723 15094 5729 15146
rect 5802 15109 5848 15431
rect 5793 15057 5799 15109
rect 5851 15057 5857 15109
rect 5665 14932 5671 14984
rect 5723 14932 5729 14984
rect 5555 14820 5561 14872
rect 5613 14820 5619 14872
rect 5665 14730 5671 14782
rect 5723 14730 5729 14782
rect 5802 14693 5848 15057
rect 6226 15051 6274 15431
rect 6658 15051 6706 15431
rect 7032 15408 7038 15460
rect 7090 15408 7096 15460
rect 7304 15408 7310 15460
rect 7362 15408 7368 15460
rect 7050 15065 7078 15408
rect 7322 15065 7350 15408
rect 6218 14999 6224 15051
rect 6276 14999 6282 15051
rect 6650 14999 6656 15051
rect 6708 14999 6714 15051
rect 7032 15013 7038 15065
rect 7090 15013 7096 15065
rect 7304 15013 7310 15065
rect 7362 15013 7368 15065
rect 6226 14693 6274 14999
rect 6658 14693 6706 14999
rect 5793 14641 5799 14693
rect 5851 14641 5857 14693
rect 6218 14641 6224 14693
rect 6276 14641 6282 14693
rect 6650 14641 6656 14693
rect 6708 14641 6714 14693
rect 7050 14670 7078 15013
rect 7322 14670 7350 15013
rect 5665 14506 5671 14558
rect 5723 14506 5729 14558
rect 5555 14416 5561 14468
rect 5613 14416 5619 14468
rect 5665 14304 5671 14356
rect 5723 14304 5729 14356
rect 5802 14319 5848 14641
rect 5793 14267 5799 14319
rect 5851 14267 5857 14319
rect 5665 14142 5671 14194
rect 5723 14142 5729 14194
rect 5555 14030 5561 14082
rect 5613 14030 5619 14082
rect 5665 13940 5671 13992
rect 5723 13940 5729 13992
rect 5802 13903 5848 14267
rect 6226 14261 6274 14641
rect 6658 14261 6706 14641
rect 7032 14618 7038 14670
rect 7090 14618 7096 14670
rect 7304 14618 7310 14670
rect 7362 14618 7368 14670
rect 7050 14275 7078 14618
rect 7322 14275 7350 14618
rect 6218 14209 6224 14261
rect 6276 14209 6282 14261
rect 6650 14209 6656 14261
rect 6708 14209 6714 14261
rect 7032 14223 7038 14275
rect 7090 14223 7096 14275
rect 7304 14223 7310 14275
rect 7362 14223 7368 14275
rect 6226 13903 6274 14209
rect 6658 13903 6706 14209
rect 5793 13851 5799 13903
rect 5851 13851 5857 13903
rect 6218 13851 6224 13903
rect 6276 13851 6282 13903
rect 6650 13851 6656 13903
rect 6708 13851 6714 13903
rect 7050 13880 7078 14223
rect 7322 13880 7350 14223
rect 5665 13716 5671 13768
rect 5723 13716 5729 13768
rect 5555 13626 5561 13678
rect 5613 13626 5619 13678
rect 5665 13514 5671 13566
rect 5723 13514 5729 13566
rect 5802 13529 5848 13851
rect 5793 13477 5799 13529
rect 5851 13477 5857 13529
rect 5665 13352 5671 13404
rect 5723 13352 5729 13404
rect 5555 13240 5561 13292
rect 5613 13240 5619 13292
rect 5665 13150 5671 13202
rect 5723 13150 5729 13202
rect 5802 13113 5848 13477
rect 6226 13471 6274 13851
rect 6658 13471 6706 13851
rect 7032 13828 7038 13880
rect 7090 13828 7096 13880
rect 7304 13828 7310 13880
rect 7362 13828 7368 13880
rect 7050 13485 7078 13828
rect 7322 13485 7350 13828
rect 6218 13419 6224 13471
rect 6276 13419 6282 13471
rect 6650 13419 6656 13471
rect 6708 13419 6714 13471
rect 7032 13433 7038 13485
rect 7090 13433 7096 13485
rect 7304 13433 7310 13485
rect 7362 13433 7368 13485
rect 6226 13113 6274 13419
rect 6658 13113 6706 13419
rect 5793 13061 5799 13113
rect 5851 13061 5857 13113
rect 6218 13061 6224 13113
rect 6276 13061 6282 13113
rect 6650 13061 6656 13113
rect 6708 13061 6714 13113
rect 7050 13090 7078 13433
rect 7322 13090 7350 13433
rect 5665 12926 5671 12978
rect 5723 12926 5729 12978
rect 5555 12836 5561 12888
rect 5613 12836 5619 12888
rect 5665 12724 5671 12776
rect 5723 12724 5729 12776
rect 5802 12739 5848 13061
rect 5793 12687 5799 12739
rect 5851 12687 5857 12739
rect 5665 12562 5671 12614
rect 5723 12562 5729 12614
rect 5555 12450 5561 12502
rect 5613 12450 5619 12502
rect 5665 12360 5671 12412
rect 5723 12360 5729 12412
rect 5802 12323 5848 12687
rect 6226 12681 6274 13061
rect 6658 12681 6706 13061
rect 7032 13038 7038 13090
rect 7090 13038 7096 13090
rect 7304 13038 7310 13090
rect 7362 13038 7368 13090
rect 7050 12695 7078 13038
rect 7322 12695 7350 13038
rect 6218 12629 6224 12681
rect 6276 12629 6282 12681
rect 6650 12629 6656 12681
rect 6708 12629 6714 12681
rect 7032 12643 7038 12695
rect 7090 12643 7096 12695
rect 7304 12643 7310 12695
rect 7362 12643 7368 12695
rect 6226 12323 6274 12629
rect 6658 12323 6706 12629
rect 5793 12271 5799 12323
rect 5851 12271 5857 12323
rect 6218 12271 6224 12323
rect 6276 12271 6282 12323
rect 6650 12271 6656 12323
rect 6708 12271 6714 12323
rect 7050 12300 7078 12643
rect 7322 12300 7350 12643
rect 5665 12136 5671 12188
rect 5723 12136 5729 12188
rect 5555 12046 5561 12098
rect 5613 12046 5619 12098
rect 5665 11934 5671 11986
rect 5723 11934 5729 11986
rect 5802 11949 5848 12271
rect 5793 11897 5799 11949
rect 5851 11897 5857 11949
rect 5665 11772 5671 11824
rect 5723 11772 5729 11824
rect 5555 11660 5561 11712
rect 5613 11660 5619 11712
rect 5665 11570 5671 11622
rect 5723 11570 5729 11622
rect 5802 11533 5848 11897
rect 6226 11891 6274 12271
rect 6658 11891 6706 12271
rect 7032 12248 7038 12300
rect 7090 12248 7096 12300
rect 7304 12248 7310 12300
rect 7362 12248 7368 12300
rect 7050 11905 7078 12248
rect 7322 11905 7350 12248
rect 6218 11839 6224 11891
rect 6276 11839 6282 11891
rect 6650 11839 6656 11891
rect 6708 11839 6714 11891
rect 7032 11853 7038 11905
rect 7090 11853 7096 11905
rect 7304 11853 7310 11905
rect 7362 11853 7368 11905
rect 6226 11533 6274 11839
rect 6658 11533 6706 11839
rect 5793 11481 5799 11533
rect 5851 11481 5857 11533
rect 6218 11481 6224 11533
rect 6276 11481 6282 11533
rect 6650 11481 6656 11533
rect 6708 11481 6714 11533
rect 7050 11510 7078 11853
rect 7322 11510 7350 11853
rect 5665 11346 5671 11398
rect 5723 11346 5729 11398
rect 5555 11256 5561 11308
rect 5613 11256 5619 11308
rect 5665 11144 5671 11196
rect 5723 11144 5729 11196
rect 5802 11159 5848 11481
rect 5793 11107 5799 11159
rect 5851 11107 5857 11159
rect 5665 10982 5671 11034
rect 5723 10982 5729 11034
rect 5555 10870 5561 10922
rect 5613 10870 5619 10922
rect 5665 10780 5671 10832
rect 5723 10780 5729 10832
rect 5802 10743 5848 11107
rect 6226 11101 6274 11481
rect 6658 11101 6706 11481
rect 7032 11458 7038 11510
rect 7090 11458 7096 11510
rect 7304 11458 7310 11510
rect 7362 11458 7368 11510
rect 7050 11115 7078 11458
rect 7322 11115 7350 11458
rect 6218 11049 6224 11101
rect 6276 11049 6282 11101
rect 6650 11049 6656 11101
rect 6708 11049 6714 11101
rect 7032 11063 7038 11115
rect 7090 11063 7096 11115
rect 7304 11063 7310 11115
rect 7362 11063 7368 11115
rect 6226 10743 6274 11049
rect 6658 10743 6706 11049
rect 5793 10691 5799 10743
rect 5851 10691 5857 10743
rect 6218 10691 6224 10743
rect 6276 10691 6282 10743
rect 6650 10691 6656 10743
rect 6708 10691 6714 10743
rect 7050 10720 7078 11063
rect 7322 10720 7350 11063
rect 5665 10556 5671 10608
rect 5723 10556 5729 10608
rect 5555 10466 5561 10518
rect 5613 10466 5619 10518
rect 5665 10354 5671 10406
rect 5723 10354 5729 10406
rect 5802 10369 5848 10691
rect 5793 10317 5799 10369
rect 5851 10317 5857 10369
rect 5665 10192 5671 10244
rect 5723 10192 5729 10244
rect 5555 10080 5561 10132
rect 5613 10080 5619 10132
rect 5665 9990 5671 10042
rect 5723 9990 5729 10042
rect 5802 9953 5848 10317
rect 6226 10311 6274 10691
rect 6658 10311 6706 10691
rect 7032 10668 7038 10720
rect 7090 10668 7096 10720
rect 7304 10668 7310 10720
rect 7362 10668 7368 10720
rect 7050 10325 7078 10668
rect 7322 10325 7350 10668
rect 6218 10259 6224 10311
rect 6276 10259 6282 10311
rect 6650 10259 6656 10311
rect 6708 10259 6714 10311
rect 7032 10273 7038 10325
rect 7090 10273 7096 10325
rect 7304 10273 7310 10325
rect 7362 10273 7368 10325
rect 6226 9953 6274 10259
rect 6658 9953 6706 10259
rect 5793 9901 5799 9953
rect 5851 9901 5857 9953
rect 6218 9901 6224 9953
rect 6276 9901 6282 9953
rect 6650 9901 6656 9953
rect 6708 9901 6714 9953
rect 7050 9930 7078 10273
rect 7322 9930 7350 10273
rect 5665 9766 5671 9818
rect 5723 9766 5729 9818
rect 5555 9676 5561 9728
rect 5613 9676 5619 9728
rect 5665 9564 5671 9616
rect 5723 9564 5729 9616
rect 5802 9579 5848 9901
rect 5793 9527 5799 9579
rect 5851 9527 5857 9579
rect 5665 9402 5671 9454
rect 5723 9402 5729 9454
rect 5555 9290 5561 9342
rect 5613 9290 5619 9342
rect 5665 9200 5671 9252
rect 5723 9200 5729 9252
rect 5802 9163 5848 9527
rect 6226 9521 6274 9901
rect 6658 9521 6706 9901
rect 7032 9878 7038 9930
rect 7090 9878 7096 9930
rect 7304 9878 7310 9930
rect 7362 9878 7368 9930
rect 7050 9535 7078 9878
rect 7322 9535 7350 9878
rect 6218 9469 6224 9521
rect 6276 9469 6282 9521
rect 6650 9469 6656 9521
rect 6708 9469 6714 9521
rect 7032 9483 7038 9535
rect 7090 9483 7096 9535
rect 7304 9483 7310 9535
rect 7362 9483 7368 9535
rect 6226 9163 6274 9469
rect 6658 9163 6706 9469
rect 5793 9111 5799 9163
rect 5851 9111 5857 9163
rect 6218 9111 6224 9163
rect 6276 9111 6282 9163
rect 6650 9111 6656 9163
rect 6708 9111 6714 9163
rect 7050 9140 7078 9483
rect 7322 9140 7350 9483
rect 5665 8976 5671 9028
rect 5723 8976 5729 9028
rect 5555 8886 5561 8938
rect 5613 8886 5619 8938
rect 5665 8774 5671 8826
rect 5723 8774 5729 8826
rect 5802 8789 5848 9111
rect 5793 8737 5799 8789
rect 5851 8737 5857 8789
rect 5665 8612 5671 8664
rect 5723 8612 5729 8664
rect 5555 8500 5561 8552
rect 5613 8500 5619 8552
rect 5665 8410 5671 8462
rect 5723 8410 5729 8462
rect 5802 8373 5848 8737
rect 6226 8731 6274 9111
rect 6658 8731 6706 9111
rect 7032 9088 7038 9140
rect 7090 9088 7096 9140
rect 7304 9088 7310 9140
rect 7362 9088 7368 9140
rect 7050 8745 7078 9088
rect 7322 8745 7350 9088
rect 6218 8679 6224 8731
rect 6276 8679 6282 8731
rect 6650 8679 6656 8731
rect 6708 8679 6714 8731
rect 7032 8693 7038 8745
rect 7090 8693 7096 8745
rect 7304 8693 7310 8745
rect 7362 8693 7368 8745
rect 6226 8373 6274 8679
rect 6658 8373 6706 8679
rect 5793 8321 5799 8373
rect 5851 8321 5857 8373
rect 6218 8321 6224 8373
rect 6276 8321 6282 8373
rect 6650 8321 6656 8373
rect 6708 8321 6714 8373
rect 7050 8350 7078 8693
rect 7322 8350 7350 8693
rect 5665 8186 5671 8238
rect 5723 8186 5729 8238
rect 5555 8096 5561 8148
rect 5613 8096 5619 8148
rect 5665 7984 5671 8036
rect 5723 7984 5729 8036
rect 5802 7999 5848 8321
rect 5793 7947 5799 7999
rect 5851 7947 5857 7999
rect 5665 7822 5671 7874
rect 5723 7822 5729 7874
rect 5555 7710 5561 7762
rect 5613 7710 5619 7762
rect 5665 7620 5671 7672
rect 5723 7620 5729 7672
rect 5802 7583 5848 7947
rect 6226 7941 6274 8321
rect 6658 7941 6706 8321
rect 7032 8298 7038 8350
rect 7090 8298 7096 8350
rect 7304 8298 7310 8350
rect 7362 8298 7368 8350
rect 7050 7955 7078 8298
rect 7322 7955 7350 8298
rect 6218 7889 6224 7941
rect 6276 7889 6282 7941
rect 6650 7889 6656 7941
rect 6708 7889 6714 7941
rect 7032 7903 7038 7955
rect 7090 7903 7096 7955
rect 7304 7903 7310 7955
rect 7362 7903 7368 7955
rect 6226 7583 6274 7889
rect 6658 7583 6706 7889
rect 5465 7551 5511 7563
rect 5465 7517 5471 7551
rect 5505 7517 5511 7551
rect 5793 7531 5799 7583
rect 5851 7531 5857 7583
rect 6218 7531 6224 7583
rect 6276 7531 6282 7583
rect 6650 7531 6656 7583
rect 6708 7531 6714 7583
rect 7050 7560 7078 7903
rect 7322 7560 7350 7903
rect 5465 7505 5511 7517
rect 5385 7156 5431 7168
rect 5385 7122 5391 7156
rect 5425 7122 5431 7156
rect 5385 7110 5431 7122
rect 5305 6761 5351 6773
rect 5305 6727 5311 6761
rect 5345 6727 5351 6761
rect 5305 6715 5351 6727
rect 5225 6366 5271 6378
rect 5225 6332 5231 6366
rect 5265 6332 5271 6366
rect 5225 6320 5271 6332
rect 5145 5971 5191 5983
rect 5145 5937 5151 5971
rect 5185 5937 5191 5971
rect 5145 5925 5191 5937
rect 5065 5576 5111 5588
rect 5065 5542 5071 5576
rect 5105 5542 5111 5576
rect 5065 5530 5111 5542
rect 4985 5181 5031 5193
rect 4985 5147 4991 5181
rect 5025 5147 5031 5181
rect 4985 5135 5031 5147
rect 4902 5078 4954 5084
rect 4902 5020 4954 5026
rect 4822 4988 4874 4994
rect 4822 4930 4874 4936
rect 4742 4602 4794 4608
rect 4742 4544 4794 4550
rect 4754 4204 4782 4544
rect 4742 4198 4794 4204
rect 4742 4140 4794 4146
rect 4754 3818 4782 4140
rect 4742 3812 4794 3818
rect 4742 3754 4794 3760
rect 4754 3414 4782 3754
rect 4834 3613 4862 4930
rect 4914 4798 4942 5020
rect 4905 4786 4951 4798
rect 4905 4752 4911 4786
rect 4945 4752 4951 4786
rect 4905 4740 4951 4752
rect 4914 4518 4942 4740
rect 4902 4512 4954 4518
rect 4902 4454 4954 4460
rect 4914 4294 4942 4454
rect 4902 4288 4954 4294
rect 4902 4230 4954 4236
rect 4914 3728 4942 4230
rect 4902 3722 4954 3728
rect 4902 3664 4954 3670
rect 4825 3601 4871 3613
rect 4825 3567 4831 3601
rect 4865 3567 4871 3601
rect 4825 3555 4871 3567
rect 4742 3408 4794 3414
rect 4742 3350 4794 3356
rect 4754 3218 4782 3350
rect 4745 3206 4791 3218
rect 4745 3172 4751 3206
rect 4785 3172 4791 3206
rect 4745 3160 4791 3172
rect 4662 3022 4714 3028
rect 4662 2964 4714 2970
rect 4674 2823 4702 2964
rect 4665 2811 4711 2823
rect 4665 2777 4671 2811
rect 4705 2777 4711 2811
rect 4665 2765 4711 2777
rect 4674 2624 4702 2765
rect 4662 2618 4714 2624
rect 4662 2560 4714 2566
rect 4585 2416 4631 2428
rect 4585 2382 4591 2416
rect 4625 2382 4631 2416
rect 4585 2370 4631 2382
rect 4502 1554 4554 1560
rect 4502 1496 4554 1502
rect 4514 1243 4542 1496
rect 4594 1448 4622 2370
rect 4674 2238 4702 2560
rect 4662 2232 4714 2238
rect 4662 2174 4714 2180
rect 4674 1834 4702 2174
rect 4662 1828 4714 1834
rect 4662 1770 4714 1776
rect 4582 1442 4634 1448
rect 4582 1384 4634 1390
rect 4505 1231 4551 1243
rect 4505 1197 4511 1231
rect 4545 1197 4551 1231
rect 4505 1185 4551 1197
rect 4422 926 4474 932
rect 4422 868 4474 874
rect 4434 848 4462 868
rect 4425 836 4471 848
rect 4425 802 4431 836
rect 4465 802 4471 836
rect 4425 790 4471 802
rect 4342 764 4394 770
rect 4342 706 4394 712
rect 4354 453 4382 706
rect 4345 441 4391 453
rect 4345 407 4351 441
rect 4385 407 4391 441
rect 4345 395 4391 407
rect 4262 136 4314 142
rect 4262 78 4314 84
rect 4274 58 4302 78
rect 4265 46 4311 58
rect 4265 12 4271 46
rect 4305 12 4311 46
rect 4354 29 4382 395
rect 4434 29 4462 790
rect 4514 29 4542 1185
rect 4594 1044 4622 1384
rect 4582 1038 4634 1044
rect 4582 980 4634 986
rect 4594 658 4622 980
rect 4582 652 4634 658
rect 4582 594 4634 600
rect 4594 254 4622 594
rect 4582 248 4634 254
rect 4582 190 4634 196
rect 4594 29 4622 190
rect 4674 29 4702 1770
rect 4754 29 4782 3160
rect 4834 29 4862 3555
rect 4914 3504 4942 3664
rect 4902 3498 4954 3504
rect 4902 3440 4954 3446
rect 4914 2938 4942 3440
rect 4902 2932 4954 2938
rect 4902 2874 4954 2880
rect 4914 2714 4942 2874
rect 4902 2708 4954 2714
rect 4902 2650 4954 2656
rect 4914 2148 4942 2650
rect 4902 2142 4954 2148
rect 4902 2084 4954 2090
rect 4914 1924 4942 2084
rect 4902 1918 4954 1924
rect 4902 1860 4954 1866
rect 4914 1358 4942 1860
rect 4902 1352 4954 1358
rect 4902 1294 4954 1300
rect 4914 1134 4942 1294
rect 4902 1128 4954 1134
rect 4902 1070 4954 1076
rect 4914 568 4942 1070
rect 4902 562 4954 568
rect 4902 504 4954 510
rect 4914 344 4942 504
rect 4902 338 4954 344
rect 4902 280 4954 286
rect 4914 29 4942 280
rect 4994 29 5022 5135
rect 5074 29 5102 5530
rect 5154 29 5182 5925
rect 5234 29 5262 6320
rect 5314 29 5342 6715
rect 5394 29 5422 7110
rect 5474 29 5502 7505
rect 5665 7396 5671 7448
rect 5723 7396 5729 7448
rect 5555 7306 5561 7358
rect 5613 7306 5619 7358
rect 5665 7194 5671 7246
rect 5723 7194 5729 7246
rect 5802 7209 5848 7531
rect 5793 7157 5799 7209
rect 5851 7157 5857 7209
rect 5665 7032 5671 7084
rect 5723 7032 5729 7084
rect 5555 6920 5561 6972
rect 5613 6920 5619 6972
rect 5665 6830 5671 6882
rect 5723 6830 5729 6882
rect 5802 6793 5848 7157
rect 6226 7151 6274 7531
rect 6658 7151 6706 7531
rect 7032 7508 7038 7560
rect 7090 7508 7096 7560
rect 7304 7508 7310 7560
rect 7362 7508 7368 7560
rect 7050 7165 7078 7508
rect 7322 7165 7350 7508
rect 6218 7099 6224 7151
rect 6276 7099 6282 7151
rect 6650 7099 6656 7151
rect 6708 7099 6714 7151
rect 7032 7113 7038 7165
rect 7090 7113 7096 7165
rect 7304 7113 7310 7165
rect 7362 7113 7368 7165
rect 6226 6793 6274 7099
rect 6658 6793 6706 7099
rect 5793 6741 5799 6793
rect 5851 6741 5857 6793
rect 6218 6741 6224 6793
rect 6276 6741 6282 6793
rect 6650 6741 6656 6793
rect 6708 6741 6714 6793
rect 7050 6770 7078 7113
rect 7322 6770 7350 7113
rect 5665 6606 5671 6658
rect 5723 6606 5729 6658
rect 5555 6516 5561 6568
rect 5613 6516 5619 6568
rect 5665 6404 5671 6456
rect 5723 6404 5729 6456
rect 5802 6419 5848 6741
rect 5793 6367 5799 6419
rect 5851 6367 5857 6419
rect 5665 6242 5671 6294
rect 5723 6242 5729 6294
rect 5555 6130 5561 6182
rect 5613 6130 5619 6182
rect 5665 6040 5671 6092
rect 5723 6040 5729 6092
rect 5802 6003 5848 6367
rect 6226 6361 6274 6741
rect 6658 6361 6706 6741
rect 7032 6718 7038 6770
rect 7090 6718 7096 6770
rect 7304 6718 7310 6770
rect 7362 6718 7368 6770
rect 7050 6375 7078 6718
rect 7322 6375 7350 6718
rect 6218 6309 6224 6361
rect 6276 6309 6282 6361
rect 6650 6309 6656 6361
rect 6708 6309 6714 6361
rect 7032 6323 7038 6375
rect 7090 6323 7096 6375
rect 7304 6323 7310 6375
rect 7362 6323 7368 6375
rect 6226 6003 6274 6309
rect 6658 6003 6706 6309
rect 5793 5951 5799 6003
rect 5851 5951 5857 6003
rect 6218 5951 6224 6003
rect 6276 5951 6282 6003
rect 6650 5951 6656 6003
rect 6708 5951 6714 6003
rect 7050 5980 7078 6323
rect 7322 5980 7350 6323
rect 5665 5816 5671 5868
rect 5723 5816 5729 5868
rect 5555 5726 5561 5778
rect 5613 5726 5619 5778
rect 5665 5614 5671 5666
rect 5723 5614 5729 5666
rect 5802 5629 5848 5951
rect 5793 5577 5799 5629
rect 5851 5577 5857 5629
rect 5665 5452 5671 5504
rect 5723 5452 5729 5504
rect 5555 5340 5561 5392
rect 5613 5340 5619 5392
rect 5665 5250 5671 5302
rect 5723 5250 5729 5302
rect 5802 5213 5848 5577
rect 6226 5571 6274 5951
rect 6658 5571 6706 5951
rect 7032 5928 7038 5980
rect 7090 5928 7096 5980
rect 7304 5928 7310 5980
rect 7362 5928 7368 5980
rect 7050 5585 7078 5928
rect 7322 5585 7350 5928
rect 6218 5519 6224 5571
rect 6276 5519 6282 5571
rect 6650 5519 6656 5571
rect 6708 5519 6714 5571
rect 7032 5533 7038 5585
rect 7090 5533 7096 5585
rect 7304 5533 7310 5585
rect 7362 5533 7368 5585
rect 6226 5213 6274 5519
rect 6658 5213 6706 5519
rect 5793 5161 5799 5213
rect 5851 5161 5857 5213
rect 6218 5161 6224 5213
rect 6276 5161 6282 5213
rect 6650 5161 6656 5213
rect 6708 5161 6714 5213
rect 7050 5190 7078 5533
rect 7322 5190 7350 5533
rect 5665 5026 5671 5078
rect 5723 5026 5729 5078
rect 5555 4936 5561 4988
rect 5613 4936 5619 4988
rect 5665 4824 5671 4876
rect 5723 4824 5729 4876
rect 5802 4839 5848 5161
rect 5793 4787 5799 4839
rect 5851 4787 5857 4839
rect 5665 4662 5671 4714
rect 5723 4662 5729 4714
rect 5555 4550 5561 4602
rect 5613 4550 5619 4602
rect 5665 4460 5671 4512
rect 5723 4460 5729 4512
rect 5802 4423 5848 4787
rect 6226 4781 6274 5161
rect 6658 4781 6706 5161
rect 7032 5138 7038 5190
rect 7090 5138 7096 5190
rect 7304 5138 7310 5190
rect 7362 5138 7368 5190
rect 7050 4795 7078 5138
rect 7322 4795 7350 5138
rect 6218 4729 6224 4781
rect 6276 4729 6282 4781
rect 6650 4729 6656 4781
rect 6708 4729 6714 4781
rect 7032 4743 7038 4795
rect 7090 4743 7096 4795
rect 7304 4743 7310 4795
rect 7362 4743 7368 4795
rect 6226 4423 6274 4729
rect 6658 4423 6706 4729
rect 5793 4371 5799 4423
rect 5851 4371 5857 4423
rect 6218 4371 6224 4423
rect 6276 4371 6282 4423
rect 6650 4371 6656 4423
rect 6708 4371 6714 4423
rect 7050 4400 7078 4743
rect 7322 4400 7350 4743
rect 5665 4236 5671 4288
rect 5723 4236 5729 4288
rect 5555 4146 5561 4198
rect 5613 4146 5619 4198
rect 5665 4034 5671 4086
rect 5723 4034 5729 4086
rect 5802 4049 5848 4371
rect 5793 3997 5799 4049
rect 5851 3997 5857 4049
rect 5665 3872 5671 3924
rect 5723 3872 5729 3924
rect 5555 3760 5561 3812
rect 5613 3760 5619 3812
rect 5665 3670 5671 3722
rect 5723 3670 5729 3722
rect 5802 3633 5848 3997
rect 6226 3991 6274 4371
rect 6658 3991 6706 4371
rect 7032 4348 7038 4400
rect 7090 4348 7096 4400
rect 7304 4348 7310 4400
rect 7362 4348 7368 4400
rect 7050 4005 7078 4348
rect 7322 4005 7350 4348
rect 6218 3939 6224 3991
rect 6276 3939 6282 3991
rect 6650 3939 6656 3991
rect 6708 3939 6714 3991
rect 7032 3953 7038 4005
rect 7090 3953 7096 4005
rect 7304 3953 7310 4005
rect 7362 3953 7368 4005
rect 6226 3633 6274 3939
rect 6658 3633 6706 3939
rect 5793 3581 5799 3633
rect 5851 3581 5857 3633
rect 6218 3581 6224 3633
rect 6276 3581 6282 3633
rect 6650 3581 6656 3633
rect 6708 3581 6714 3633
rect 7050 3610 7078 3953
rect 7322 3610 7350 3953
rect 5665 3446 5671 3498
rect 5723 3446 5729 3498
rect 5555 3356 5561 3408
rect 5613 3356 5619 3408
rect 5665 3244 5671 3296
rect 5723 3244 5729 3296
rect 5802 3259 5848 3581
rect 5793 3207 5799 3259
rect 5851 3207 5857 3259
rect 5665 3082 5671 3134
rect 5723 3082 5729 3134
rect 5555 2970 5561 3022
rect 5613 2970 5619 3022
rect 5665 2880 5671 2932
rect 5723 2880 5729 2932
rect 5802 2843 5848 3207
rect 6226 3201 6274 3581
rect 6658 3201 6706 3581
rect 7032 3558 7038 3610
rect 7090 3558 7096 3610
rect 7304 3558 7310 3610
rect 7362 3558 7368 3610
rect 7050 3215 7078 3558
rect 7322 3215 7350 3558
rect 6218 3149 6224 3201
rect 6276 3149 6282 3201
rect 6650 3149 6656 3201
rect 6708 3149 6714 3201
rect 7032 3163 7038 3215
rect 7090 3163 7096 3215
rect 7304 3163 7310 3215
rect 7362 3163 7368 3215
rect 6226 2843 6274 3149
rect 6658 2843 6706 3149
rect 5793 2791 5799 2843
rect 5851 2791 5857 2843
rect 6218 2791 6224 2843
rect 6276 2791 6282 2843
rect 6650 2791 6656 2843
rect 6708 2791 6714 2843
rect 7050 2820 7078 3163
rect 7322 2820 7350 3163
rect 5665 2656 5671 2708
rect 5723 2656 5729 2708
rect 5555 2566 5561 2618
rect 5613 2566 5619 2618
rect 5665 2454 5671 2506
rect 5723 2454 5729 2506
rect 5802 2469 5848 2791
rect 5793 2417 5799 2469
rect 5851 2417 5857 2469
rect 5665 2292 5671 2344
rect 5723 2292 5729 2344
rect 5555 2180 5561 2232
rect 5613 2180 5619 2232
rect 5665 2090 5671 2142
rect 5723 2090 5729 2142
rect 5802 2053 5848 2417
rect 6226 2411 6274 2791
rect 6658 2411 6706 2791
rect 7032 2768 7038 2820
rect 7090 2768 7096 2820
rect 7304 2768 7310 2820
rect 7362 2768 7368 2820
rect 7050 2425 7078 2768
rect 7322 2425 7350 2768
rect 6218 2359 6224 2411
rect 6276 2359 6282 2411
rect 6650 2359 6656 2411
rect 6708 2359 6714 2411
rect 7032 2373 7038 2425
rect 7090 2373 7096 2425
rect 7304 2373 7310 2425
rect 7362 2373 7368 2425
rect 6226 2053 6274 2359
rect 6658 2053 6706 2359
rect 5793 2001 5799 2053
rect 5851 2001 5857 2053
rect 6218 2001 6224 2053
rect 6276 2001 6282 2053
rect 6650 2001 6656 2053
rect 6708 2001 6714 2053
rect 7050 2030 7078 2373
rect 7322 2030 7350 2373
rect 5665 1866 5671 1918
rect 5723 1866 5729 1918
rect 5555 1776 5561 1828
rect 5613 1776 5619 1828
rect 5665 1664 5671 1716
rect 5723 1664 5729 1716
rect 5802 1679 5848 2001
rect 5793 1627 5799 1679
rect 5851 1627 5857 1679
rect 5665 1502 5671 1554
rect 5723 1502 5729 1554
rect 5555 1390 5561 1442
rect 5613 1390 5619 1442
rect 5665 1300 5671 1352
rect 5723 1300 5729 1352
rect 5802 1263 5848 1627
rect 6226 1621 6274 2001
rect 6658 1621 6706 2001
rect 7032 1978 7038 2030
rect 7090 1978 7096 2030
rect 7304 1978 7310 2030
rect 7362 1978 7368 2030
rect 7050 1635 7078 1978
rect 7322 1635 7350 1978
rect 6218 1569 6224 1621
rect 6276 1569 6282 1621
rect 6650 1569 6656 1621
rect 6708 1569 6714 1621
rect 7032 1583 7038 1635
rect 7090 1583 7096 1635
rect 7304 1583 7310 1635
rect 7362 1583 7368 1635
rect 6226 1263 6274 1569
rect 6658 1263 6706 1569
rect 5793 1211 5799 1263
rect 5851 1211 5857 1263
rect 6218 1211 6224 1263
rect 6276 1211 6282 1263
rect 6650 1211 6656 1263
rect 6708 1211 6714 1263
rect 7050 1240 7078 1583
rect 7322 1240 7350 1583
rect 5665 1076 5671 1128
rect 5723 1076 5729 1128
rect 5555 986 5561 1038
rect 5613 986 5619 1038
rect 5665 874 5671 926
rect 5723 874 5729 926
rect 5802 889 5848 1211
rect 5793 837 5799 889
rect 5851 837 5857 889
rect 5665 712 5671 764
rect 5723 712 5729 764
rect 5555 600 5561 652
rect 5613 600 5619 652
rect 5665 510 5671 562
rect 5723 510 5729 562
rect 5802 473 5848 837
rect 6226 831 6274 1211
rect 6658 831 6706 1211
rect 7032 1188 7038 1240
rect 7090 1188 7096 1240
rect 7304 1188 7310 1240
rect 7362 1188 7368 1240
rect 7050 845 7078 1188
rect 7322 845 7350 1188
rect 6218 779 6224 831
rect 6276 779 6282 831
rect 6650 779 6656 831
rect 6708 779 6714 831
rect 7032 793 7038 845
rect 7090 793 7096 845
rect 7304 793 7310 845
rect 7362 793 7368 845
rect 6226 473 6274 779
rect 6658 473 6706 779
rect 5793 421 5799 473
rect 5851 421 5857 473
rect 6218 421 6224 473
rect 6276 421 6282 473
rect 6650 421 6656 473
rect 6708 421 6714 473
rect 7050 450 7078 793
rect 7322 450 7350 793
rect 5665 286 5671 338
rect 5723 286 5729 338
rect 5555 196 5561 248
rect 5613 196 5619 248
rect 5665 84 5671 136
rect 5723 84 5729 136
rect 5802 13 5848 421
rect 6226 71 6274 421
rect 6658 71 6706 421
rect 7032 398 7038 450
rect 7090 398 7096 450
rect 7304 398 7310 450
rect 7362 398 7368 450
rect 7050 57 7078 398
rect 7322 57 7350 398
rect 4265 0 4311 12
<< via1 >>
rect 4502 50482 4554 50534
rect 4422 49854 4474 49906
rect 4342 49692 4394 49744
rect 4262 49064 4314 49116
rect 4502 48902 4554 48954
rect 4422 48274 4474 48326
rect 4342 48112 4394 48164
rect 4262 47484 4314 47536
rect 4502 47322 4554 47374
rect 4422 46694 4474 46746
rect 4342 46532 4394 46584
rect 4262 45904 4314 45956
rect 4502 45742 4554 45794
rect 4422 45114 4474 45166
rect 4342 44952 4394 45004
rect 4262 44324 4314 44376
rect 4822 50370 4874 50422
rect 4822 49966 4874 50018
rect 4822 49580 4874 49632
rect 4822 49176 4874 49228
rect 4742 48790 4794 48842
rect 4742 48386 4794 48438
rect 4742 48000 4794 48052
rect 4742 47596 4794 47648
rect 4662 47210 4714 47262
rect 4662 46806 4714 46858
rect 4662 46420 4714 46472
rect 4662 46016 4714 46068
rect 4582 45630 4634 45682
rect 4582 45226 4634 45278
rect 4582 44840 4634 44892
rect 4582 44436 4634 44488
rect 4502 44162 4554 44214
rect 4422 43534 4474 43586
rect 4342 43372 4394 43424
rect 4262 42744 4314 42796
rect 4502 42582 4554 42634
rect 4422 41954 4474 42006
rect 4342 41792 4394 41844
rect 4262 41164 4314 41216
rect 4502 41002 4554 41054
rect 4422 40374 4474 40426
rect 4342 40212 4394 40264
rect 4262 39584 4314 39636
rect 4502 39422 4554 39474
rect 4422 38794 4474 38846
rect 4342 38632 4394 38684
rect 4262 38004 4314 38056
rect 4822 44050 4874 44102
rect 4822 43646 4874 43698
rect 4822 43260 4874 43312
rect 4822 42856 4874 42908
rect 4742 42470 4794 42522
rect 4742 42066 4794 42118
rect 4742 41680 4794 41732
rect 4742 41276 4794 41328
rect 4662 40890 4714 40942
rect 4662 40486 4714 40538
rect 4662 40100 4714 40152
rect 4662 39696 4714 39748
rect 4582 39310 4634 39362
rect 4582 38906 4634 38958
rect 4582 38520 4634 38572
rect 4582 38116 4634 38168
rect 4502 37842 4554 37894
rect 4422 37214 4474 37266
rect 4342 37052 4394 37104
rect 4262 36424 4314 36476
rect 4502 36262 4554 36314
rect 4422 35634 4474 35686
rect 4342 35472 4394 35524
rect 4262 34844 4314 34896
rect 4502 34682 4554 34734
rect 4422 34054 4474 34106
rect 4342 33892 4394 33944
rect 4262 33264 4314 33316
rect 4502 33102 4554 33154
rect 4422 32474 4474 32526
rect 4342 32312 4394 32364
rect 4262 31684 4314 31736
rect 4822 37730 4874 37782
rect 4822 37326 4874 37378
rect 4822 36940 4874 36992
rect 4822 36536 4874 36588
rect 4742 36150 4794 36202
rect 4742 35746 4794 35798
rect 4742 35360 4794 35412
rect 4742 34956 4794 35008
rect 4662 34570 4714 34622
rect 4662 34166 4714 34218
rect 4662 33780 4714 33832
rect 4662 33376 4714 33428
rect 4582 32990 4634 33042
rect 4582 32586 4634 32638
rect 4582 32200 4634 32252
rect 4582 31796 4634 31848
rect 4502 31522 4554 31574
rect 4422 30894 4474 30946
rect 4342 30732 4394 30784
rect 4262 30104 4314 30156
rect 4502 29942 4554 29994
rect 4422 29314 4474 29366
rect 4342 29152 4394 29204
rect 4262 28524 4314 28576
rect 4502 28362 4554 28414
rect 4422 27734 4474 27786
rect 4342 27572 4394 27624
rect 4262 26944 4314 26996
rect 4502 26782 4554 26834
rect 4422 26154 4474 26206
rect 4342 25992 4394 26044
rect 4262 25364 4314 25416
rect 4822 31410 4874 31462
rect 4822 31006 4874 31058
rect 4822 30620 4874 30672
rect 4822 30216 4874 30268
rect 4742 29830 4794 29882
rect 4742 29426 4794 29478
rect 4742 29040 4794 29092
rect 4742 28636 4794 28688
rect 4662 28250 4714 28302
rect 4662 27846 4714 27898
rect 4662 27460 4714 27512
rect 4662 27056 4714 27108
rect 4582 26670 4634 26722
rect 4582 26266 4634 26318
rect 4582 25880 4634 25932
rect 4582 25476 4634 25528
rect 4502 25202 4554 25254
rect 4422 24574 4474 24626
rect 4342 24412 4394 24464
rect 4262 23784 4314 23836
rect 4502 23622 4554 23674
rect 4422 22994 4474 23046
rect 4342 22832 4394 22884
rect 4262 22204 4314 22256
rect 4502 22042 4554 22094
rect 4422 21414 4474 21466
rect 4342 21252 4394 21304
rect 4262 20624 4314 20676
rect 4502 20462 4554 20514
rect 4422 19834 4474 19886
rect 4342 19672 4394 19724
rect 4262 19044 4314 19096
rect 4822 25090 4874 25142
rect 4822 24686 4874 24738
rect 4822 24300 4874 24352
rect 4822 23896 4874 23948
rect 4742 23510 4794 23562
rect 4742 23106 4794 23158
rect 4742 22720 4794 22772
rect 4742 22316 4794 22368
rect 4662 21930 4714 21982
rect 4662 21526 4714 21578
rect 4662 21140 4714 21192
rect 4662 20736 4714 20788
rect 4582 20350 4634 20402
rect 4582 19946 4634 19998
rect 4582 19560 4634 19612
rect 4582 19156 4634 19208
rect 4502 18882 4554 18934
rect 4422 18254 4474 18306
rect 4342 18092 4394 18144
rect 4262 17464 4314 17516
rect 4502 17302 4554 17354
rect 4422 16674 4474 16726
rect 4342 16512 4394 16564
rect 4262 15884 4314 15936
rect 4502 15722 4554 15774
rect 4422 15094 4474 15146
rect 4342 14932 4394 14984
rect 4262 14304 4314 14356
rect 4502 14142 4554 14194
rect 4422 13514 4474 13566
rect 4342 13352 4394 13404
rect 4262 12724 4314 12776
rect 4822 18770 4874 18822
rect 4822 18366 4874 18418
rect 4822 17980 4874 18032
rect 4822 17576 4874 17628
rect 4742 17190 4794 17242
rect 4742 16786 4794 16838
rect 4742 16400 4794 16452
rect 4742 15996 4794 16048
rect 4662 15610 4714 15662
rect 4662 15206 4714 15258
rect 4662 14820 4714 14872
rect 4662 14416 4714 14468
rect 4582 14030 4634 14082
rect 4582 13626 4634 13678
rect 4582 13240 4634 13292
rect 4582 12836 4634 12888
rect 4502 12562 4554 12614
rect 4422 11934 4474 11986
rect 4342 11772 4394 11824
rect 4262 11144 4314 11196
rect 4502 10982 4554 11034
rect 4422 10354 4474 10406
rect 4342 10192 4394 10244
rect 4262 9564 4314 9616
rect 4502 9402 4554 9454
rect 4422 8774 4474 8826
rect 4342 8612 4394 8664
rect 4262 7984 4314 8036
rect 4502 7822 4554 7874
rect 4422 7194 4474 7246
rect 4342 7032 4394 7084
rect 4262 6404 4314 6456
rect 486 5730 538 5782
rect 834 5730 886 5782
rect 406 5336 458 5388
rect 326 4940 378 4992
rect 246 2966 298 3018
rect 166 2570 218 2622
rect 86 596 138 648
rect 6 200 58 252
rect 754 5336 806 5388
rect 674 4940 726 4992
rect 4822 12450 4874 12502
rect 4822 12046 4874 12098
rect 4822 11660 4874 11712
rect 4822 11256 4874 11308
rect 4742 10870 4794 10922
rect 4742 10466 4794 10518
rect 4742 10080 4794 10132
rect 4742 9676 4794 9728
rect 4662 9290 4714 9342
rect 4662 8886 4714 8938
rect 4662 8500 4714 8552
rect 4662 8096 4714 8148
rect 4582 7710 4634 7762
rect 4582 7306 4634 7358
rect 4582 6920 4634 6972
rect 4582 6516 4634 6568
rect 4502 6242 4554 6294
rect 4422 5614 4474 5666
rect 4342 5452 4394 5504
rect 4262 4824 4314 4876
rect 4502 4662 4554 4714
rect 4422 4034 4474 4086
rect 4342 3872 4394 3924
rect 4262 3244 4314 3296
rect 1430 2966 1482 3018
rect 1350 2570 1402 2622
rect 4502 3082 4554 3134
rect 4422 2454 4474 2506
rect 4342 2292 4394 2344
rect 4262 1664 4314 1716
rect 1430 596 1482 648
rect 1350 200 1402 252
rect 4822 6130 4874 6182
rect 5671 50525 5723 50534
rect 5671 50491 5680 50525
rect 5680 50491 5714 50525
rect 5714 50491 5723 50525
rect 5671 50482 5723 50491
rect 5561 50413 5613 50422
rect 5561 50379 5570 50413
rect 5570 50379 5604 50413
rect 5604 50379 5613 50413
rect 5561 50370 5613 50379
rect 5462 50280 5514 50332
rect 5671 50323 5723 50332
rect 5671 50289 5680 50323
rect 5680 50289 5714 50323
rect 5714 50289 5723 50323
rect 5671 50280 5723 50289
rect 5799 50191 5851 50243
rect 6224 50191 6276 50243
rect 6656 50191 6708 50243
rect 5462 50056 5514 50108
rect 5671 50099 5723 50108
rect 5671 50065 5680 50099
rect 5680 50065 5714 50099
rect 5714 50065 5723 50099
rect 5671 50056 5723 50065
rect 5561 50009 5613 50018
rect 5561 49975 5570 50009
rect 5570 49975 5604 50009
rect 5604 49975 5613 50009
rect 5561 49966 5613 49975
rect 5671 49897 5723 49906
rect 5671 49863 5680 49897
rect 5680 49863 5714 49897
rect 5714 49863 5723 49897
rect 5671 49854 5723 49863
rect 5799 49817 5851 49869
rect 5671 49735 5723 49744
rect 5671 49701 5680 49735
rect 5680 49701 5714 49735
rect 5714 49701 5723 49735
rect 5671 49692 5723 49701
rect 5561 49623 5613 49632
rect 5561 49589 5570 49623
rect 5570 49589 5604 49623
rect 5604 49589 5613 49623
rect 5561 49580 5613 49589
rect 5462 49490 5514 49542
rect 5671 49533 5723 49542
rect 5671 49499 5680 49533
rect 5680 49499 5714 49533
rect 5714 49499 5723 49533
rect 5671 49490 5723 49499
rect 7038 50168 7090 50220
rect 7310 50168 7362 50220
rect 6224 49759 6276 49811
rect 6656 49759 6708 49811
rect 7038 49773 7090 49825
rect 7310 49773 7362 49825
rect 5799 49401 5851 49453
rect 6224 49401 6276 49453
rect 6656 49401 6708 49453
rect 5462 49266 5514 49318
rect 5671 49309 5723 49318
rect 5671 49275 5680 49309
rect 5680 49275 5714 49309
rect 5714 49275 5723 49309
rect 5671 49266 5723 49275
rect 5561 49219 5613 49228
rect 5561 49185 5570 49219
rect 5570 49185 5604 49219
rect 5604 49185 5613 49219
rect 5561 49176 5613 49185
rect 5671 49107 5723 49116
rect 5671 49073 5680 49107
rect 5680 49073 5714 49107
rect 5714 49073 5723 49107
rect 5671 49064 5723 49073
rect 5799 49027 5851 49079
rect 5671 48945 5723 48954
rect 5671 48911 5680 48945
rect 5680 48911 5714 48945
rect 5714 48911 5723 48945
rect 5671 48902 5723 48911
rect 5561 48833 5613 48842
rect 5561 48799 5570 48833
rect 5570 48799 5604 48833
rect 5604 48799 5613 48833
rect 5561 48790 5613 48799
rect 5462 48700 5514 48752
rect 5671 48743 5723 48752
rect 5671 48709 5680 48743
rect 5680 48709 5714 48743
rect 5714 48709 5723 48743
rect 5671 48700 5723 48709
rect 7038 49378 7090 49430
rect 7310 49378 7362 49430
rect 6224 48969 6276 49021
rect 6656 48969 6708 49021
rect 7038 48983 7090 49035
rect 7310 48983 7362 49035
rect 5799 48611 5851 48663
rect 6224 48611 6276 48663
rect 6656 48611 6708 48663
rect 5462 48476 5514 48528
rect 5671 48519 5723 48528
rect 5671 48485 5680 48519
rect 5680 48485 5714 48519
rect 5714 48485 5723 48519
rect 5671 48476 5723 48485
rect 5561 48429 5613 48438
rect 5561 48395 5570 48429
rect 5570 48395 5604 48429
rect 5604 48395 5613 48429
rect 5561 48386 5613 48395
rect 5671 48317 5723 48326
rect 5671 48283 5680 48317
rect 5680 48283 5714 48317
rect 5714 48283 5723 48317
rect 5671 48274 5723 48283
rect 5799 48237 5851 48289
rect 5671 48155 5723 48164
rect 5671 48121 5680 48155
rect 5680 48121 5714 48155
rect 5714 48121 5723 48155
rect 5671 48112 5723 48121
rect 5561 48043 5613 48052
rect 5561 48009 5570 48043
rect 5570 48009 5604 48043
rect 5604 48009 5613 48043
rect 5561 48000 5613 48009
rect 5462 47910 5514 47962
rect 5671 47953 5723 47962
rect 5671 47919 5680 47953
rect 5680 47919 5714 47953
rect 5714 47919 5723 47953
rect 5671 47910 5723 47919
rect 7038 48588 7090 48640
rect 7310 48588 7362 48640
rect 6224 48179 6276 48231
rect 6656 48179 6708 48231
rect 7038 48193 7090 48245
rect 7310 48193 7362 48245
rect 5799 47821 5851 47873
rect 6224 47821 6276 47873
rect 6656 47821 6708 47873
rect 5462 47686 5514 47738
rect 5671 47729 5723 47738
rect 5671 47695 5680 47729
rect 5680 47695 5714 47729
rect 5714 47695 5723 47729
rect 5671 47686 5723 47695
rect 5561 47639 5613 47648
rect 5561 47605 5570 47639
rect 5570 47605 5604 47639
rect 5604 47605 5613 47639
rect 5561 47596 5613 47605
rect 5671 47527 5723 47536
rect 5671 47493 5680 47527
rect 5680 47493 5714 47527
rect 5714 47493 5723 47527
rect 5671 47484 5723 47493
rect 5799 47447 5851 47499
rect 5671 47365 5723 47374
rect 5671 47331 5680 47365
rect 5680 47331 5714 47365
rect 5714 47331 5723 47365
rect 5671 47322 5723 47331
rect 5561 47253 5613 47262
rect 5561 47219 5570 47253
rect 5570 47219 5604 47253
rect 5604 47219 5613 47253
rect 5561 47210 5613 47219
rect 5462 47120 5514 47172
rect 5671 47163 5723 47172
rect 5671 47129 5680 47163
rect 5680 47129 5714 47163
rect 5714 47129 5723 47163
rect 5671 47120 5723 47129
rect 7038 47798 7090 47850
rect 7310 47798 7362 47850
rect 6224 47389 6276 47441
rect 6656 47389 6708 47441
rect 7038 47403 7090 47455
rect 7310 47403 7362 47455
rect 5799 47031 5851 47083
rect 6224 47031 6276 47083
rect 6656 47031 6708 47083
rect 5462 46896 5514 46948
rect 5671 46939 5723 46948
rect 5671 46905 5680 46939
rect 5680 46905 5714 46939
rect 5714 46905 5723 46939
rect 5671 46896 5723 46905
rect 5561 46849 5613 46858
rect 5561 46815 5570 46849
rect 5570 46815 5604 46849
rect 5604 46815 5613 46849
rect 5561 46806 5613 46815
rect 5671 46737 5723 46746
rect 5671 46703 5680 46737
rect 5680 46703 5714 46737
rect 5714 46703 5723 46737
rect 5671 46694 5723 46703
rect 5799 46657 5851 46709
rect 5671 46575 5723 46584
rect 5671 46541 5680 46575
rect 5680 46541 5714 46575
rect 5714 46541 5723 46575
rect 5671 46532 5723 46541
rect 5561 46463 5613 46472
rect 5561 46429 5570 46463
rect 5570 46429 5604 46463
rect 5604 46429 5613 46463
rect 5561 46420 5613 46429
rect 5462 46330 5514 46382
rect 5671 46373 5723 46382
rect 5671 46339 5680 46373
rect 5680 46339 5714 46373
rect 5714 46339 5723 46373
rect 5671 46330 5723 46339
rect 7038 47008 7090 47060
rect 7310 47008 7362 47060
rect 6224 46599 6276 46651
rect 6656 46599 6708 46651
rect 7038 46613 7090 46665
rect 7310 46613 7362 46665
rect 5799 46241 5851 46293
rect 6224 46241 6276 46293
rect 6656 46241 6708 46293
rect 5462 46106 5514 46158
rect 5671 46149 5723 46158
rect 5671 46115 5680 46149
rect 5680 46115 5714 46149
rect 5714 46115 5723 46149
rect 5671 46106 5723 46115
rect 5561 46059 5613 46068
rect 5561 46025 5570 46059
rect 5570 46025 5604 46059
rect 5604 46025 5613 46059
rect 5561 46016 5613 46025
rect 5671 45947 5723 45956
rect 5671 45913 5680 45947
rect 5680 45913 5714 45947
rect 5714 45913 5723 45947
rect 5671 45904 5723 45913
rect 5799 45867 5851 45919
rect 5671 45785 5723 45794
rect 5671 45751 5680 45785
rect 5680 45751 5714 45785
rect 5714 45751 5723 45785
rect 5671 45742 5723 45751
rect 5561 45673 5613 45682
rect 5561 45639 5570 45673
rect 5570 45639 5604 45673
rect 5604 45639 5613 45673
rect 5561 45630 5613 45639
rect 5462 45540 5514 45592
rect 5671 45583 5723 45592
rect 5671 45549 5680 45583
rect 5680 45549 5714 45583
rect 5714 45549 5723 45583
rect 5671 45540 5723 45549
rect 7038 46218 7090 46270
rect 7310 46218 7362 46270
rect 6224 45809 6276 45861
rect 6656 45809 6708 45861
rect 7038 45823 7090 45875
rect 7310 45823 7362 45875
rect 5799 45451 5851 45503
rect 6224 45451 6276 45503
rect 6656 45451 6708 45503
rect 5462 45316 5514 45368
rect 5671 45359 5723 45368
rect 5671 45325 5680 45359
rect 5680 45325 5714 45359
rect 5714 45325 5723 45359
rect 5671 45316 5723 45325
rect 5561 45269 5613 45278
rect 5561 45235 5570 45269
rect 5570 45235 5604 45269
rect 5604 45235 5613 45269
rect 5561 45226 5613 45235
rect 5671 45157 5723 45166
rect 5671 45123 5680 45157
rect 5680 45123 5714 45157
rect 5714 45123 5723 45157
rect 5671 45114 5723 45123
rect 5799 45077 5851 45129
rect 5671 44995 5723 45004
rect 5671 44961 5680 44995
rect 5680 44961 5714 44995
rect 5714 44961 5723 44995
rect 5671 44952 5723 44961
rect 5561 44883 5613 44892
rect 5561 44849 5570 44883
rect 5570 44849 5604 44883
rect 5604 44849 5613 44883
rect 5561 44840 5613 44849
rect 5462 44750 5514 44802
rect 5671 44793 5723 44802
rect 5671 44759 5680 44793
rect 5680 44759 5714 44793
rect 5714 44759 5723 44793
rect 5671 44750 5723 44759
rect 7038 45428 7090 45480
rect 7310 45428 7362 45480
rect 6224 45019 6276 45071
rect 6656 45019 6708 45071
rect 7038 45033 7090 45085
rect 7310 45033 7362 45085
rect 5799 44661 5851 44713
rect 6224 44661 6276 44713
rect 6656 44661 6708 44713
rect 5462 44526 5514 44578
rect 5671 44569 5723 44578
rect 5671 44535 5680 44569
rect 5680 44535 5714 44569
rect 5714 44535 5723 44569
rect 5671 44526 5723 44535
rect 5382 43960 5434 44012
rect 5382 43736 5434 43788
rect 5382 43170 5434 43222
rect 5382 42946 5434 42998
rect 5382 42380 5434 42432
rect 5382 42156 5434 42208
rect 5382 41590 5434 41642
rect 5382 41366 5434 41418
rect 5382 40800 5434 40852
rect 5382 40576 5434 40628
rect 5382 40010 5434 40062
rect 5382 39786 5434 39838
rect 5382 39220 5434 39272
rect 5382 38996 5434 39048
rect 5382 38430 5434 38482
rect 5382 38206 5434 38258
rect 5302 37640 5354 37692
rect 5302 37416 5354 37468
rect 5302 36850 5354 36902
rect 5302 36626 5354 36678
rect 5302 36060 5354 36112
rect 5302 35836 5354 35888
rect 5302 35270 5354 35322
rect 5302 35046 5354 35098
rect 5302 34480 5354 34532
rect 5302 34256 5354 34308
rect 5302 33690 5354 33742
rect 5302 33466 5354 33518
rect 5302 32900 5354 32952
rect 5302 32676 5354 32728
rect 5302 32110 5354 32162
rect 5302 31886 5354 31938
rect 5222 31320 5274 31372
rect 5222 31096 5274 31148
rect 5222 30530 5274 30582
rect 5222 30306 5274 30358
rect 5222 29740 5274 29792
rect 5222 29516 5274 29568
rect 5222 28950 5274 29002
rect 5222 28726 5274 28778
rect 5222 28160 5274 28212
rect 5222 27936 5274 27988
rect 5222 27370 5274 27422
rect 5222 27146 5274 27198
rect 5222 26580 5274 26632
rect 5222 26356 5274 26408
rect 5222 25790 5274 25842
rect 5222 25566 5274 25618
rect 5142 25000 5194 25052
rect 5142 24776 5194 24828
rect 5142 24210 5194 24262
rect 5142 23986 5194 24038
rect 5142 23420 5194 23472
rect 5142 23196 5194 23248
rect 5142 22630 5194 22682
rect 5142 22406 5194 22458
rect 5142 21840 5194 21892
rect 5142 21616 5194 21668
rect 5142 21050 5194 21102
rect 5142 20826 5194 20878
rect 5142 20260 5194 20312
rect 5142 20036 5194 20088
rect 5142 19470 5194 19522
rect 5142 19246 5194 19298
rect 5062 18680 5114 18732
rect 5062 18456 5114 18508
rect 5062 17890 5114 17942
rect 5062 17666 5114 17718
rect 5062 17100 5114 17152
rect 5062 16876 5114 16928
rect 5062 16310 5114 16362
rect 5062 16086 5114 16138
rect 5062 15520 5114 15572
rect 5062 15296 5114 15348
rect 5062 14730 5114 14782
rect 5062 14506 5114 14558
rect 5062 13940 5114 13992
rect 5062 13716 5114 13768
rect 5062 13150 5114 13202
rect 5062 12926 5114 12978
rect 4982 12360 5034 12412
rect 4982 12136 5034 12188
rect 4982 11570 5034 11622
rect 4982 11346 5034 11398
rect 4982 10780 5034 10832
rect 4982 10556 5034 10608
rect 4982 9990 5034 10042
rect 4982 9766 5034 9818
rect 4982 9200 5034 9252
rect 4982 8976 5034 9028
rect 4982 8410 5034 8462
rect 4982 8186 5034 8238
rect 4982 7620 5034 7672
rect 4982 7396 5034 7448
rect 4982 6830 5034 6882
rect 4982 6606 5034 6658
rect 4902 6040 4954 6092
rect 4902 5816 4954 5868
rect 4822 5726 4874 5778
rect 4822 5340 4874 5392
rect 4902 5250 4954 5302
rect 5561 44479 5613 44488
rect 5561 44445 5570 44479
rect 5570 44445 5604 44479
rect 5604 44445 5613 44479
rect 5561 44436 5613 44445
rect 5671 44367 5723 44376
rect 5671 44333 5680 44367
rect 5680 44333 5714 44367
rect 5714 44333 5723 44367
rect 5671 44324 5723 44333
rect 5799 44287 5851 44339
rect 5671 44205 5723 44214
rect 5671 44171 5680 44205
rect 5680 44171 5714 44205
rect 5714 44171 5723 44205
rect 5671 44162 5723 44171
rect 5561 44093 5613 44102
rect 5561 44059 5570 44093
rect 5570 44059 5604 44093
rect 5604 44059 5613 44093
rect 5561 44050 5613 44059
rect 5671 44003 5723 44012
rect 5671 43969 5680 44003
rect 5680 43969 5714 44003
rect 5714 43969 5723 44003
rect 5671 43960 5723 43969
rect 7038 44638 7090 44690
rect 7310 44638 7362 44690
rect 6224 44229 6276 44281
rect 6656 44229 6708 44281
rect 7038 44243 7090 44295
rect 7310 44243 7362 44295
rect 5799 43871 5851 43923
rect 6224 43871 6276 43923
rect 6656 43871 6708 43923
rect 5671 43779 5723 43788
rect 5671 43745 5680 43779
rect 5680 43745 5714 43779
rect 5714 43745 5723 43779
rect 5671 43736 5723 43745
rect 5561 43689 5613 43698
rect 5561 43655 5570 43689
rect 5570 43655 5604 43689
rect 5604 43655 5613 43689
rect 5561 43646 5613 43655
rect 5671 43577 5723 43586
rect 5671 43543 5680 43577
rect 5680 43543 5714 43577
rect 5714 43543 5723 43577
rect 5671 43534 5723 43543
rect 5799 43497 5851 43549
rect 5671 43415 5723 43424
rect 5671 43381 5680 43415
rect 5680 43381 5714 43415
rect 5714 43381 5723 43415
rect 5671 43372 5723 43381
rect 5561 43303 5613 43312
rect 5561 43269 5570 43303
rect 5570 43269 5604 43303
rect 5604 43269 5613 43303
rect 5561 43260 5613 43269
rect 5671 43213 5723 43222
rect 5671 43179 5680 43213
rect 5680 43179 5714 43213
rect 5714 43179 5723 43213
rect 5671 43170 5723 43179
rect 7038 43848 7090 43900
rect 7310 43848 7362 43900
rect 6224 43439 6276 43491
rect 6656 43439 6708 43491
rect 7038 43453 7090 43505
rect 7310 43453 7362 43505
rect 5799 43081 5851 43133
rect 6224 43081 6276 43133
rect 6656 43081 6708 43133
rect 5671 42989 5723 42998
rect 5671 42955 5680 42989
rect 5680 42955 5714 42989
rect 5714 42955 5723 42989
rect 5671 42946 5723 42955
rect 5561 42899 5613 42908
rect 5561 42865 5570 42899
rect 5570 42865 5604 42899
rect 5604 42865 5613 42899
rect 5561 42856 5613 42865
rect 5671 42787 5723 42796
rect 5671 42753 5680 42787
rect 5680 42753 5714 42787
rect 5714 42753 5723 42787
rect 5671 42744 5723 42753
rect 5799 42707 5851 42759
rect 5671 42625 5723 42634
rect 5671 42591 5680 42625
rect 5680 42591 5714 42625
rect 5714 42591 5723 42625
rect 5671 42582 5723 42591
rect 5561 42513 5613 42522
rect 5561 42479 5570 42513
rect 5570 42479 5604 42513
rect 5604 42479 5613 42513
rect 5561 42470 5613 42479
rect 5671 42423 5723 42432
rect 5671 42389 5680 42423
rect 5680 42389 5714 42423
rect 5714 42389 5723 42423
rect 5671 42380 5723 42389
rect 7038 43058 7090 43110
rect 7310 43058 7362 43110
rect 6224 42649 6276 42701
rect 6656 42649 6708 42701
rect 7038 42663 7090 42715
rect 7310 42663 7362 42715
rect 5799 42291 5851 42343
rect 6224 42291 6276 42343
rect 6656 42291 6708 42343
rect 5671 42199 5723 42208
rect 5671 42165 5680 42199
rect 5680 42165 5714 42199
rect 5714 42165 5723 42199
rect 5671 42156 5723 42165
rect 5561 42109 5613 42118
rect 5561 42075 5570 42109
rect 5570 42075 5604 42109
rect 5604 42075 5613 42109
rect 5561 42066 5613 42075
rect 5671 41997 5723 42006
rect 5671 41963 5680 41997
rect 5680 41963 5714 41997
rect 5714 41963 5723 41997
rect 5671 41954 5723 41963
rect 5799 41917 5851 41969
rect 5671 41835 5723 41844
rect 5671 41801 5680 41835
rect 5680 41801 5714 41835
rect 5714 41801 5723 41835
rect 5671 41792 5723 41801
rect 5561 41723 5613 41732
rect 5561 41689 5570 41723
rect 5570 41689 5604 41723
rect 5604 41689 5613 41723
rect 5561 41680 5613 41689
rect 5671 41633 5723 41642
rect 5671 41599 5680 41633
rect 5680 41599 5714 41633
rect 5714 41599 5723 41633
rect 5671 41590 5723 41599
rect 7038 42268 7090 42320
rect 7310 42268 7362 42320
rect 6224 41859 6276 41911
rect 6656 41859 6708 41911
rect 7038 41873 7090 41925
rect 7310 41873 7362 41925
rect 5799 41501 5851 41553
rect 6224 41501 6276 41553
rect 6656 41501 6708 41553
rect 5671 41409 5723 41418
rect 5671 41375 5680 41409
rect 5680 41375 5714 41409
rect 5714 41375 5723 41409
rect 5671 41366 5723 41375
rect 5561 41319 5613 41328
rect 5561 41285 5570 41319
rect 5570 41285 5604 41319
rect 5604 41285 5613 41319
rect 5561 41276 5613 41285
rect 5671 41207 5723 41216
rect 5671 41173 5680 41207
rect 5680 41173 5714 41207
rect 5714 41173 5723 41207
rect 5671 41164 5723 41173
rect 5799 41127 5851 41179
rect 5671 41045 5723 41054
rect 5671 41011 5680 41045
rect 5680 41011 5714 41045
rect 5714 41011 5723 41045
rect 5671 41002 5723 41011
rect 5561 40933 5613 40942
rect 5561 40899 5570 40933
rect 5570 40899 5604 40933
rect 5604 40899 5613 40933
rect 5561 40890 5613 40899
rect 5671 40843 5723 40852
rect 5671 40809 5680 40843
rect 5680 40809 5714 40843
rect 5714 40809 5723 40843
rect 5671 40800 5723 40809
rect 7038 41478 7090 41530
rect 7310 41478 7362 41530
rect 6224 41069 6276 41121
rect 6656 41069 6708 41121
rect 7038 41083 7090 41135
rect 7310 41083 7362 41135
rect 5799 40711 5851 40763
rect 6224 40711 6276 40763
rect 6656 40711 6708 40763
rect 5671 40619 5723 40628
rect 5671 40585 5680 40619
rect 5680 40585 5714 40619
rect 5714 40585 5723 40619
rect 5671 40576 5723 40585
rect 5561 40529 5613 40538
rect 5561 40495 5570 40529
rect 5570 40495 5604 40529
rect 5604 40495 5613 40529
rect 5561 40486 5613 40495
rect 5671 40417 5723 40426
rect 5671 40383 5680 40417
rect 5680 40383 5714 40417
rect 5714 40383 5723 40417
rect 5671 40374 5723 40383
rect 5799 40337 5851 40389
rect 5671 40255 5723 40264
rect 5671 40221 5680 40255
rect 5680 40221 5714 40255
rect 5714 40221 5723 40255
rect 5671 40212 5723 40221
rect 5561 40143 5613 40152
rect 5561 40109 5570 40143
rect 5570 40109 5604 40143
rect 5604 40109 5613 40143
rect 5561 40100 5613 40109
rect 5671 40053 5723 40062
rect 5671 40019 5680 40053
rect 5680 40019 5714 40053
rect 5714 40019 5723 40053
rect 5671 40010 5723 40019
rect 7038 40688 7090 40740
rect 7310 40688 7362 40740
rect 6224 40279 6276 40331
rect 6656 40279 6708 40331
rect 7038 40293 7090 40345
rect 7310 40293 7362 40345
rect 5799 39921 5851 39973
rect 6224 39921 6276 39973
rect 6656 39921 6708 39973
rect 5671 39829 5723 39838
rect 5671 39795 5680 39829
rect 5680 39795 5714 39829
rect 5714 39795 5723 39829
rect 5671 39786 5723 39795
rect 5561 39739 5613 39748
rect 5561 39705 5570 39739
rect 5570 39705 5604 39739
rect 5604 39705 5613 39739
rect 5561 39696 5613 39705
rect 5671 39627 5723 39636
rect 5671 39593 5680 39627
rect 5680 39593 5714 39627
rect 5714 39593 5723 39627
rect 5671 39584 5723 39593
rect 5799 39547 5851 39599
rect 5671 39465 5723 39474
rect 5671 39431 5680 39465
rect 5680 39431 5714 39465
rect 5714 39431 5723 39465
rect 5671 39422 5723 39431
rect 5561 39353 5613 39362
rect 5561 39319 5570 39353
rect 5570 39319 5604 39353
rect 5604 39319 5613 39353
rect 5561 39310 5613 39319
rect 5671 39263 5723 39272
rect 5671 39229 5680 39263
rect 5680 39229 5714 39263
rect 5714 39229 5723 39263
rect 5671 39220 5723 39229
rect 7038 39898 7090 39950
rect 7310 39898 7362 39950
rect 6224 39489 6276 39541
rect 6656 39489 6708 39541
rect 7038 39503 7090 39555
rect 7310 39503 7362 39555
rect 5799 39131 5851 39183
rect 6224 39131 6276 39183
rect 6656 39131 6708 39183
rect 5671 39039 5723 39048
rect 5671 39005 5680 39039
rect 5680 39005 5714 39039
rect 5714 39005 5723 39039
rect 5671 38996 5723 39005
rect 5561 38949 5613 38958
rect 5561 38915 5570 38949
rect 5570 38915 5604 38949
rect 5604 38915 5613 38949
rect 5561 38906 5613 38915
rect 5671 38837 5723 38846
rect 5671 38803 5680 38837
rect 5680 38803 5714 38837
rect 5714 38803 5723 38837
rect 5671 38794 5723 38803
rect 5799 38757 5851 38809
rect 5671 38675 5723 38684
rect 5671 38641 5680 38675
rect 5680 38641 5714 38675
rect 5714 38641 5723 38675
rect 5671 38632 5723 38641
rect 5561 38563 5613 38572
rect 5561 38529 5570 38563
rect 5570 38529 5604 38563
rect 5604 38529 5613 38563
rect 5561 38520 5613 38529
rect 5671 38473 5723 38482
rect 5671 38439 5680 38473
rect 5680 38439 5714 38473
rect 5714 38439 5723 38473
rect 5671 38430 5723 38439
rect 7038 39108 7090 39160
rect 7310 39108 7362 39160
rect 6224 38699 6276 38751
rect 6656 38699 6708 38751
rect 7038 38713 7090 38765
rect 7310 38713 7362 38765
rect 5799 38341 5851 38393
rect 6224 38341 6276 38393
rect 6656 38341 6708 38393
rect 5671 38249 5723 38258
rect 5671 38215 5680 38249
rect 5680 38215 5714 38249
rect 5714 38215 5723 38249
rect 5671 38206 5723 38215
rect 5561 38159 5613 38168
rect 5561 38125 5570 38159
rect 5570 38125 5604 38159
rect 5604 38125 5613 38159
rect 5561 38116 5613 38125
rect 5671 38047 5723 38056
rect 5671 38013 5680 38047
rect 5680 38013 5714 38047
rect 5714 38013 5723 38047
rect 5671 38004 5723 38013
rect 5799 37967 5851 38019
rect 5671 37885 5723 37894
rect 5671 37851 5680 37885
rect 5680 37851 5714 37885
rect 5714 37851 5723 37885
rect 5671 37842 5723 37851
rect 5561 37773 5613 37782
rect 5561 37739 5570 37773
rect 5570 37739 5604 37773
rect 5604 37739 5613 37773
rect 5561 37730 5613 37739
rect 5671 37683 5723 37692
rect 5671 37649 5680 37683
rect 5680 37649 5714 37683
rect 5714 37649 5723 37683
rect 5671 37640 5723 37649
rect 7038 38318 7090 38370
rect 7310 38318 7362 38370
rect 6224 37909 6276 37961
rect 6656 37909 6708 37961
rect 7038 37923 7090 37975
rect 7310 37923 7362 37975
rect 5799 37551 5851 37603
rect 6224 37551 6276 37603
rect 6656 37551 6708 37603
rect 5671 37459 5723 37468
rect 5671 37425 5680 37459
rect 5680 37425 5714 37459
rect 5714 37425 5723 37459
rect 5671 37416 5723 37425
rect 5561 37369 5613 37378
rect 5561 37335 5570 37369
rect 5570 37335 5604 37369
rect 5604 37335 5613 37369
rect 5561 37326 5613 37335
rect 5671 37257 5723 37266
rect 5671 37223 5680 37257
rect 5680 37223 5714 37257
rect 5714 37223 5723 37257
rect 5671 37214 5723 37223
rect 5799 37177 5851 37229
rect 5671 37095 5723 37104
rect 5671 37061 5680 37095
rect 5680 37061 5714 37095
rect 5714 37061 5723 37095
rect 5671 37052 5723 37061
rect 5561 36983 5613 36992
rect 5561 36949 5570 36983
rect 5570 36949 5604 36983
rect 5604 36949 5613 36983
rect 5561 36940 5613 36949
rect 5671 36893 5723 36902
rect 5671 36859 5680 36893
rect 5680 36859 5714 36893
rect 5714 36859 5723 36893
rect 5671 36850 5723 36859
rect 7038 37528 7090 37580
rect 7310 37528 7362 37580
rect 6224 37119 6276 37171
rect 6656 37119 6708 37171
rect 7038 37133 7090 37185
rect 7310 37133 7362 37185
rect 5799 36761 5851 36813
rect 6224 36761 6276 36813
rect 6656 36761 6708 36813
rect 5671 36669 5723 36678
rect 5671 36635 5680 36669
rect 5680 36635 5714 36669
rect 5714 36635 5723 36669
rect 5671 36626 5723 36635
rect 5561 36579 5613 36588
rect 5561 36545 5570 36579
rect 5570 36545 5604 36579
rect 5604 36545 5613 36579
rect 5561 36536 5613 36545
rect 5671 36467 5723 36476
rect 5671 36433 5680 36467
rect 5680 36433 5714 36467
rect 5714 36433 5723 36467
rect 5671 36424 5723 36433
rect 5799 36387 5851 36439
rect 5671 36305 5723 36314
rect 5671 36271 5680 36305
rect 5680 36271 5714 36305
rect 5714 36271 5723 36305
rect 5671 36262 5723 36271
rect 5561 36193 5613 36202
rect 5561 36159 5570 36193
rect 5570 36159 5604 36193
rect 5604 36159 5613 36193
rect 5561 36150 5613 36159
rect 5671 36103 5723 36112
rect 5671 36069 5680 36103
rect 5680 36069 5714 36103
rect 5714 36069 5723 36103
rect 5671 36060 5723 36069
rect 7038 36738 7090 36790
rect 7310 36738 7362 36790
rect 6224 36329 6276 36381
rect 6656 36329 6708 36381
rect 7038 36343 7090 36395
rect 7310 36343 7362 36395
rect 5799 35971 5851 36023
rect 6224 35971 6276 36023
rect 6656 35971 6708 36023
rect 5671 35879 5723 35888
rect 5671 35845 5680 35879
rect 5680 35845 5714 35879
rect 5714 35845 5723 35879
rect 5671 35836 5723 35845
rect 5561 35789 5613 35798
rect 5561 35755 5570 35789
rect 5570 35755 5604 35789
rect 5604 35755 5613 35789
rect 5561 35746 5613 35755
rect 5671 35677 5723 35686
rect 5671 35643 5680 35677
rect 5680 35643 5714 35677
rect 5714 35643 5723 35677
rect 5671 35634 5723 35643
rect 5799 35597 5851 35649
rect 5671 35515 5723 35524
rect 5671 35481 5680 35515
rect 5680 35481 5714 35515
rect 5714 35481 5723 35515
rect 5671 35472 5723 35481
rect 5561 35403 5613 35412
rect 5561 35369 5570 35403
rect 5570 35369 5604 35403
rect 5604 35369 5613 35403
rect 5561 35360 5613 35369
rect 5671 35313 5723 35322
rect 5671 35279 5680 35313
rect 5680 35279 5714 35313
rect 5714 35279 5723 35313
rect 5671 35270 5723 35279
rect 7038 35948 7090 36000
rect 7310 35948 7362 36000
rect 6224 35539 6276 35591
rect 6656 35539 6708 35591
rect 7038 35553 7090 35605
rect 7310 35553 7362 35605
rect 5799 35181 5851 35233
rect 6224 35181 6276 35233
rect 6656 35181 6708 35233
rect 5671 35089 5723 35098
rect 5671 35055 5680 35089
rect 5680 35055 5714 35089
rect 5714 35055 5723 35089
rect 5671 35046 5723 35055
rect 5561 34999 5613 35008
rect 5561 34965 5570 34999
rect 5570 34965 5604 34999
rect 5604 34965 5613 34999
rect 5561 34956 5613 34965
rect 5671 34887 5723 34896
rect 5671 34853 5680 34887
rect 5680 34853 5714 34887
rect 5714 34853 5723 34887
rect 5671 34844 5723 34853
rect 5799 34807 5851 34859
rect 5671 34725 5723 34734
rect 5671 34691 5680 34725
rect 5680 34691 5714 34725
rect 5714 34691 5723 34725
rect 5671 34682 5723 34691
rect 5561 34613 5613 34622
rect 5561 34579 5570 34613
rect 5570 34579 5604 34613
rect 5604 34579 5613 34613
rect 5561 34570 5613 34579
rect 5671 34523 5723 34532
rect 5671 34489 5680 34523
rect 5680 34489 5714 34523
rect 5714 34489 5723 34523
rect 5671 34480 5723 34489
rect 7038 35158 7090 35210
rect 7310 35158 7362 35210
rect 6224 34749 6276 34801
rect 6656 34749 6708 34801
rect 7038 34763 7090 34815
rect 7310 34763 7362 34815
rect 5799 34391 5851 34443
rect 6224 34391 6276 34443
rect 6656 34391 6708 34443
rect 5671 34299 5723 34308
rect 5671 34265 5680 34299
rect 5680 34265 5714 34299
rect 5714 34265 5723 34299
rect 5671 34256 5723 34265
rect 5561 34209 5613 34218
rect 5561 34175 5570 34209
rect 5570 34175 5604 34209
rect 5604 34175 5613 34209
rect 5561 34166 5613 34175
rect 5671 34097 5723 34106
rect 5671 34063 5680 34097
rect 5680 34063 5714 34097
rect 5714 34063 5723 34097
rect 5671 34054 5723 34063
rect 5799 34017 5851 34069
rect 5671 33935 5723 33944
rect 5671 33901 5680 33935
rect 5680 33901 5714 33935
rect 5714 33901 5723 33935
rect 5671 33892 5723 33901
rect 5561 33823 5613 33832
rect 5561 33789 5570 33823
rect 5570 33789 5604 33823
rect 5604 33789 5613 33823
rect 5561 33780 5613 33789
rect 5671 33733 5723 33742
rect 5671 33699 5680 33733
rect 5680 33699 5714 33733
rect 5714 33699 5723 33733
rect 5671 33690 5723 33699
rect 7038 34368 7090 34420
rect 7310 34368 7362 34420
rect 6224 33959 6276 34011
rect 6656 33959 6708 34011
rect 7038 33973 7090 34025
rect 7310 33973 7362 34025
rect 5799 33601 5851 33653
rect 6224 33601 6276 33653
rect 6656 33601 6708 33653
rect 5671 33509 5723 33518
rect 5671 33475 5680 33509
rect 5680 33475 5714 33509
rect 5714 33475 5723 33509
rect 5671 33466 5723 33475
rect 5561 33419 5613 33428
rect 5561 33385 5570 33419
rect 5570 33385 5604 33419
rect 5604 33385 5613 33419
rect 5561 33376 5613 33385
rect 5671 33307 5723 33316
rect 5671 33273 5680 33307
rect 5680 33273 5714 33307
rect 5714 33273 5723 33307
rect 5671 33264 5723 33273
rect 5799 33227 5851 33279
rect 5671 33145 5723 33154
rect 5671 33111 5680 33145
rect 5680 33111 5714 33145
rect 5714 33111 5723 33145
rect 5671 33102 5723 33111
rect 5561 33033 5613 33042
rect 5561 32999 5570 33033
rect 5570 32999 5604 33033
rect 5604 32999 5613 33033
rect 5561 32990 5613 32999
rect 5671 32943 5723 32952
rect 5671 32909 5680 32943
rect 5680 32909 5714 32943
rect 5714 32909 5723 32943
rect 5671 32900 5723 32909
rect 7038 33578 7090 33630
rect 7310 33578 7362 33630
rect 6224 33169 6276 33221
rect 6656 33169 6708 33221
rect 7038 33183 7090 33235
rect 7310 33183 7362 33235
rect 5799 32811 5851 32863
rect 6224 32811 6276 32863
rect 6656 32811 6708 32863
rect 5671 32719 5723 32728
rect 5671 32685 5680 32719
rect 5680 32685 5714 32719
rect 5714 32685 5723 32719
rect 5671 32676 5723 32685
rect 5561 32629 5613 32638
rect 5561 32595 5570 32629
rect 5570 32595 5604 32629
rect 5604 32595 5613 32629
rect 5561 32586 5613 32595
rect 5671 32517 5723 32526
rect 5671 32483 5680 32517
rect 5680 32483 5714 32517
rect 5714 32483 5723 32517
rect 5671 32474 5723 32483
rect 5799 32437 5851 32489
rect 5671 32355 5723 32364
rect 5671 32321 5680 32355
rect 5680 32321 5714 32355
rect 5714 32321 5723 32355
rect 5671 32312 5723 32321
rect 5561 32243 5613 32252
rect 5561 32209 5570 32243
rect 5570 32209 5604 32243
rect 5604 32209 5613 32243
rect 5561 32200 5613 32209
rect 5671 32153 5723 32162
rect 5671 32119 5680 32153
rect 5680 32119 5714 32153
rect 5714 32119 5723 32153
rect 5671 32110 5723 32119
rect 7038 32788 7090 32840
rect 7310 32788 7362 32840
rect 6224 32379 6276 32431
rect 6656 32379 6708 32431
rect 7038 32393 7090 32445
rect 7310 32393 7362 32445
rect 5799 32021 5851 32073
rect 6224 32021 6276 32073
rect 6656 32021 6708 32073
rect 5671 31929 5723 31938
rect 5671 31895 5680 31929
rect 5680 31895 5714 31929
rect 5714 31895 5723 31929
rect 5671 31886 5723 31895
rect 5561 31839 5613 31848
rect 5561 31805 5570 31839
rect 5570 31805 5604 31839
rect 5604 31805 5613 31839
rect 5561 31796 5613 31805
rect 5671 31727 5723 31736
rect 5671 31693 5680 31727
rect 5680 31693 5714 31727
rect 5714 31693 5723 31727
rect 5671 31684 5723 31693
rect 5799 31647 5851 31699
rect 5671 31565 5723 31574
rect 5671 31531 5680 31565
rect 5680 31531 5714 31565
rect 5714 31531 5723 31565
rect 5671 31522 5723 31531
rect 5561 31453 5613 31462
rect 5561 31419 5570 31453
rect 5570 31419 5604 31453
rect 5604 31419 5613 31453
rect 5561 31410 5613 31419
rect 5671 31363 5723 31372
rect 5671 31329 5680 31363
rect 5680 31329 5714 31363
rect 5714 31329 5723 31363
rect 5671 31320 5723 31329
rect 7038 31998 7090 32050
rect 7310 31998 7362 32050
rect 6224 31589 6276 31641
rect 6656 31589 6708 31641
rect 7038 31603 7090 31655
rect 7310 31603 7362 31655
rect 5799 31231 5851 31283
rect 6224 31231 6276 31283
rect 6656 31231 6708 31283
rect 5671 31139 5723 31148
rect 5671 31105 5680 31139
rect 5680 31105 5714 31139
rect 5714 31105 5723 31139
rect 5671 31096 5723 31105
rect 5561 31049 5613 31058
rect 5561 31015 5570 31049
rect 5570 31015 5604 31049
rect 5604 31015 5613 31049
rect 5561 31006 5613 31015
rect 5671 30937 5723 30946
rect 5671 30903 5680 30937
rect 5680 30903 5714 30937
rect 5714 30903 5723 30937
rect 5671 30894 5723 30903
rect 5799 30857 5851 30909
rect 5671 30775 5723 30784
rect 5671 30741 5680 30775
rect 5680 30741 5714 30775
rect 5714 30741 5723 30775
rect 5671 30732 5723 30741
rect 5561 30663 5613 30672
rect 5561 30629 5570 30663
rect 5570 30629 5604 30663
rect 5604 30629 5613 30663
rect 5561 30620 5613 30629
rect 5671 30573 5723 30582
rect 5671 30539 5680 30573
rect 5680 30539 5714 30573
rect 5714 30539 5723 30573
rect 5671 30530 5723 30539
rect 7038 31208 7090 31260
rect 7310 31208 7362 31260
rect 6224 30799 6276 30851
rect 6656 30799 6708 30851
rect 7038 30813 7090 30865
rect 7310 30813 7362 30865
rect 5799 30441 5851 30493
rect 6224 30441 6276 30493
rect 6656 30441 6708 30493
rect 5671 30349 5723 30358
rect 5671 30315 5680 30349
rect 5680 30315 5714 30349
rect 5714 30315 5723 30349
rect 5671 30306 5723 30315
rect 5561 30259 5613 30268
rect 5561 30225 5570 30259
rect 5570 30225 5604 30259
rect 5604 30225 5613 30259
rect 5561 30216 5613 30225
rect 5671 30147 5723 30156
rect 5671 30113 5680 30147
rect 5680 30113 5714 30147
rect 5714 30113 5723 30147
rect 5671 30104 5723 30113
rect 5799 30067 5851 30119
rect 5671 29985 5723 29994
rect 5671 29951 5680 29985
rect 5680 29951 5714 29985
rect 5714 29951 5723 29985
rect 5671 29942 5723 29951
rect 5561 29873 5613 29882
rect 5561 29839 5570 29873
rect 5570 29839 5604 29873
rect 5604 29839 5613 29873
rect 5561 29830 5613 29839
rect 5671 29783 5723 29792
rect 5671 29749 5680 29783
rect 5680 29749 5714 29783
rect 5714 29749 5723 29783
rect 5671 29740 5723 29749
rect 7038 30418 7090 30470
rect 7310 30418 7362 30470
rect 6224 30009 6276 30061
rect 6656 30009 6708 30061
rect 7038 30023 7090 30075
rect 7310 30023 7362 30075
rect 5799 29651 5851 29703
rect 6224 29651 6276 29703
rect 6656 29651 6708 29703
rect 5671 29559 5723 29568
rect 5671 29525 5680 29559
rect 5680 29525 5714 29559
rect 5714 29525 5723 29559
rect 5671 29516 5723 29525
rect 5561 29469 5613 29478
rect 5561 29435 5570 29469
rect 5570 29435 5604 29469
rect 5604 29435 5613 29469
rect 5561 29426 5613 29435
rect 5671 29357 5723 29366
rect 5671 29323 5680 29357
rect 5680 29323 5714 29357
rect 5714 29323 5723 29357
rect 5671 29314 5723 29323
rect 5799 29277 5851 29329
rect 5671 29195 5723 29204
rect 5671 29161 5680 29195
rect 5680 29161 5714 29195
rect 5714 29161 5723 29195
rect 5671 29152 5723 29161
rect 5561 29083 5613 29092
rect 5561 29049 5570 29083
rect 5570 29049 5604 29083
rect 5604 29049 5613 29083
rect 5561 29040 5613 29049
rect 5671 28993 5723 29002
rect 5671 28959 5680 28993
rect 5680 28959 5714 28993
rect 5714 28959 5723 28993
rect 5671 28950 5723 28959
rect 7038 29628 7090 29680
rect 7310 29628 7362 29680
rect 6224 29219 6276 29271
rect 6656 29219 6708 29271
rect 7038 29233 7090 29285
rect 7310 29233 7362 29285
rect 5799 28861 5851 28913
rect 6224 28861 6276 28913
rect 6656 28861 6708 28913
rect 5671 28769 5723 28778
rect 5671 28735 5680 28769
rect 5680 28735 5714 28769
rect 5714 28735 5723 28769
rect 5671 28726 5723 28735
rect 5561 28679 5613 28688
rect 5561 28645 5570 28679
rect 5570 28645 5604 28679
rect 5604 28645 5613 28679
rect 5561 28636 5613 28645
rect 5671 28567 5723 28576
rect 5671 28533 5680 28567
rect 5680 28533 5714 28567
rect 5714 28533 5723 28567
rect 5671 28524 5723 28533
rect 5799 28487 5851 28539
rect 5671 28405 5723 28414
rect 5671 28371 5680 28405
rect 5680 28371 5714 28405
rect 5714 28371 5723 28405
rect 5671 28362 5723 28371
rect 5561 28293 5613 28302
rect 5561 28259 5570 28293
rect 5570 28259 5604 28293
rect 5604 28259 5613 28293
rect 5561 28250 5613 28259
rect 5671 28203 5723 28212
rect 5671 28169 5680 28203
rect 5680 28169 5714 28203
rect 5714 28169 5723 28203
rect 5671 28160 5723 28169
rect 7038 28838 7090 28890
rect 7310 28838 7362 28890
rect 6224 28429 6276 28481
rect 6656 28429 6708 28481
rect 7038 28443 7090 28495
rect 7310 28443 7362 28495
rect 5799 28071 5851 28123
rect 6224 28071 6276 28123
rect 6656 28071 6708 28123
rect 5671 27979 5723 27988
rect 5671 27945 5680 27979
rect 5680 27945 5714 27979
rect 5714 27945 5723 27979
rect 5671 27936 5723 27945
rect 5561 27889 5613 27898
rect 5561 27855 5570 27889
rect 5570 27855 5604 27889
rect 5604 27855 5613 27889
rect 5561 27846 5613 27855
rect 5671 27777 5723 27786
rect 5671 27743 5680 27777
rect 5680 27743 5714 27777
rect 5714 27743 5723 27777
rect 5671 27734 5723 27743
rect 5799 27697 5851 27749
rect 5671 27615 5723 27624
rect 5671 27581 5680 27615
rect 5680 27581 5714 27615
rect 5714 27581 5723 27615
rect 5671 27572 5723 27581
rect 5561 27503 5613 27512
rect 5561 27469 5570 27503
rect 5570 27469 5604 27503
rect 5604 27469 5613 27503
rect 5561 27460 5613 27469
rect 5671 27413 5723 27422
rect 5671 27379 5680 27413
rect 5680 27379 5714 27413
rect 5714 27379 5723 27413
rect 5671 27370 5723 27379
rect 7038 28048 7090 28100
rect 7310 28048 7362 28100
rect 6224 27639 6276 27691
rect 6656 27639 6708 27691
rect 7038 27653 7090 27705
rect 7310 27653 7362 27705
rect 5799 27281 5851 27333
rect 6224 27281 6276 27333
rect 6656 27281 6708 27333
rect 5671 27189 5723 27198
rect 5671 27155 5680 27189
rect 5680 27155 5714 27189
rect 5714 27155 5723 27189
rect 5671 27146 5723 27155
rect 5561 27099 5613 27108
rect 5561 27065 5570 27099
rect 5570 27065 5604 27099
rect 5604 27065 5613 27099
rect 5561 27056 5613 27065
rect 5671 26987 5723 26996
rect 5671 26953 5680 26987
rect 5680 26953 5714 26987
rect 5714 26953 5723 26987
rect 5671 26944 5723 26953
rect 5799 26907 5851 26959
rect 5671 26825 5723 26834
rect 5671 26791 5680 26825
rect 5680 26791 5714 26825
rect 5714 26791 5723 26825
rect 5671 26782 5723 26791
rect 5561 26713 5613 26722
rect 5561 26679 5570 26713
rect 5570 26679 5604 26713
rect 5604 26679 5613 26713
rect 5561 26670 5613 26679
rect 5671 26623 5723 26632
rect 5671 26589 5680 26623
rect 5680 26589 5714 26623
rect 5714 26589 5723 26623
rect 5671 26580 5723 26589
rect 7038 27258 7090 27310
rect 7310 27258 7362 27310
rect 6224 26849 6276 26901
rect 6656 26849 6708 26901
rect 7038 26863 7090 26915
rect 7310 26863 7362 26915
rect 5799 26491 5851 26543
rect 6224 26491 6276 26543
rect 6656 26491 6708 26543
rect 5671 26399 5723 26408
rect 5671 26365 5680 26399
rect 5680 26365 5714 26399
rect 5714 26365 5723 26399
rect 5671 26356 5723 26365
rect 5561 26309 5613 26318
rect 5561 26275 5570 26309
rect 5570 26275 5604 26309
rect 5604 26275 5613 26309
rect 5561 26266 5613 26275
rect 5671 26197 5723 26206
rect 5671 26163 5680 26197
rect 5680 26163 5714 26197
rect 5714 26163 5723 26197
rect 5671 26154 5723 26163
rect 5799 26117 5851 26169
rect 5671 26035 5723 26044
rect 5671 26001 5680 26035
rect 5680 26001 5714 26035
rect 5714 26001 5723 26035
rect 5671 25992 5723 26001
rect 5561 25923 5613 25932
rect 5561 25889 5570 25923
rect 5570 25889 5604 25923
rect 5604 25889 5613 25923
rect 5561 25880 5613 25889
rect 5671 25833 5723 25842
rect 5671 25799 5680 25833
rect 5680 25799 5714 25833
rect 5714 25799 5723 25833
rect 5671 25790 5723 25799
rect 7038 26468 7090 26520
rect 7310 26468 7362 26520
rect 6224 26059 6276 26111
rect 6656 26059 6708 26111
rect 7038 26073 7090 26125
rect 7310 26073 7362 26125
rect 5799 25701 5851 25753
rect 6224 25701 6276 25753
rect 6656 25701 6708 25753
rect 5671 25609 5723 25618
rect 5671 25575 5680 25609
rect 5680 25575 5714 25609
rect 5714 25575 5723 25609
rect 5671 25566 5723 25575
rect 5561 25519 5613 25528
rect 5561 25485 5570 25519
rect 5570 25485 5604 25519
rect 5604 25485 5613 25519
rect 5561 25476 5613 25485
rect 5671 25407 5723 25416
rect 5671 25373 5680 25407
rect 5680 25373 5714 25407
rect 5714 25373 5723 25407
rect 5671 25364 5723 25373
rect 5799 25327 5851 25379
rect 5671 25245 5723 25254
rect 5671 25211 5680 25245
rect 5680 25211 5714 25245
rect 5714 25211 5723 25245
rect 5671 25202 5723 25211
rect 5561 25133 5613 25142
rect 5561 25099 5570 25133
rect 5570 25099 5604 25133
rect 5604 25099 5613 25133
rect 5561 25090 5613 25099
rect 5671 25043 5723 25052
rect 5671 25009 5680 25043
rect 5680 25009 5714 25043
rect 5714 25009 5723 25043
rect 5671 25000 5723 25009
rect 7038 25678 7090 25730
rect 7310 25678 7362 25730
rect 6224 25269 6276 25321
rect 6656 25269 6708 25321
rect 7038 25283 7090 25335
rect 7310 25283 7362 25335
rect 5799 24911 5851 24963
rect 6224 24911 6276 24963
rect 6656 24911 6708 24963
rect 5671 24819 5723 24828
rect 5671 24785 5680 24819
rect 5680 24785 5714 24819
rect 5714 24785 5723 24819
rect 5671 24776 5723 24785
rect 5561 24729 5613 24738
rect 5561 24695 5570 24729
rect 5570 24695 5604 24729
rect 5604 24695 5613 24729
rect 5561 24686 5613 24695
rect 5671 24617 5723 24626
rect 5671 24583 5680 24617
rect 5680 24583 5714 24617
rect 5714 24583 5723 24617
rect 5671 24574 5723 24583
rect 5799 24537 5851 24589
rect 5671 24455 5723 24464
rect 5671 24421 5680 24455
rect 5680 24421 5714 24455
rect 5714 24421 5723 24455
rect 5671 24412 5723 24421
rect 5561 24343 5613 24352
rect 5561 24309 5570 24343
rect 5570 24309 5604 24343
rect 5604 24309 5613 24343
rect 5561 24300 5613 24309
rect 5671 24253 5723 24262
rect 5671 24219 5680 24253
rect 5680 24219 5714 24253
rect 5714 24219 5723 24253
rect 5671 24210 5723 24219
rect 7038 24888 7090 24940
rect 7310 24888 7362 24940
rect 6224 24479 6276 24531
rect 6656 24479 6708 24531
rect 7038 24493 7090 24545
rect 7310 24493 7362 24545
rect 5799 24121 5851 24173
rect 6224 24121 6276 24173
rect 6656 24121 6708 24173
rect 5671 24029 5723 24038
rect 5671 23995 5680 24029
rect 5680 23995 5714 24029
rect 5714 23995 5723 24029
rect 5671 23986 5723 23995
rect 5561 23939 5613 23948
rect 5561 23905 5570 23939
rect 5570 23905 5604 23939
rect 5604 23905 5613 23939
rect 5561 23896 5613 23905
rect 5671 23827 5723 23836
rect 5671 23793 5680 23827
rect 5680 23793 5714 23827
rect 5714 23793 5723 23827
rect 5671 23784 5723 23793
rect 5799 23747 5851 23799
rect 5671 23665 5723 23674
rect 5671 23631 5680 23665
rect 5680 23631 5714 23665
rect 5714 23631 5723 23665
rect 5671 23622 5723 23631
rect 5561 23553 5613 23562
rect 5561 23519 5570 23553
rect 5570 23519 5604 23553
rect 5604 23519 5613 23553
rect 5561 23510 5613 23519
rect 5671 23463 5723 23472
rect 5671 23429 5680 23463
rect 5680 23429 5714 23463
rect 5714 23429 5723 23463
rect 5671 23420 5723 23429
rect 7038 24098 7090 24150
rect 7310 24098 7362 24150
rect 6224 23689 6276 23741
rect 6656 23689 6708 23741
rect 7038 23703 7090 23755
rect 7310 23703 7362 23755
rect 5799 23331 5851 23383
rect 6224 23331 6276 23383
rect 6656 23331 6708 23383
rect 5671 23239 5723 23248
rect 5671 23205 5680 23239
rect 5680 23205 5714 23239
rect 5714 23205 5723 23239
rect 5671 23196 5723 23205
rect 5561 23149 5613 23158
rect 5561 23115 5570 23149
rect 5570 23115 5604 23149
rect 5604 23115 5613 23149
rect 5561 23106 5613 23115
rect 5671 23037 5723 23046
rect 5671 23003 5680 23037
rect 5680 23003 5714 23037
rect 5714 23003 5723 23037
rect 5671 22994 5723 23003
rect 5799 22957 5851 23009
rect 5671 22875 5723 22884
rect 5671 22841 5680 22875
rect 5680 22841 5714 22875
rect 5714 22841 5723 22875
rect 5671 22832 5723 22841
rect 5561 22763 5613 22772
rect 5561 22729 5570 22763
rect 5570 22729 5604 22763
rect 5604 22729 5613 22763
rect 5561 22720 5613 22729
rect 5671 22673 5723 22682
rect 5671 22639 5680 22673
rect 5680 22639 5714 22673
rect 5714 22639 5723 22673
rect 5671 22630 5723 22639
rect 7038 23308 7090 23360
rect 7310 23308 7362 23360
rect 6224 22899 6276 22951
rect 6656 22899 6708 22951
rect 7038 22913 7090 22965
rect 7310 22913 7362 22965
rect 5799 22541 5851 22593
rect 6224 22541 6276 22593
rect 6656 22541 6708 22593
rect 5671 22449 5723 22458
rect 5671 22415 5680 22449
rect 5680 22415 5714 22449
rect 5714 22415 5723 22449
rect 5671 22406 5723 22415
rect 5561 22359 5613 22368
rect 5561 22325 5570 22359
rect 5570 22325 5604 22359
rect 5604 22325 5613 22359
rect 5561 22316 5613 22325
rect 5671 22247 5723 22256
rect 5671 22213 5680 22247
rect 5680 22213 5714 22247
rect 5714 22213 5723 22247
rect 5671 22204 5723 22213
rect 5799 22167 5851 22219
rect 5671 22085 5723 22094
rect 5671 22051 5680 22085
rect 5680 22051 5714 22085
rect 5714 22051 5723 22085
rect 5671 22042 5723 22051
rect 5561 21973 5613 21982
rect 5561 21939 5570 21973
rect 5570 21939 5604 21973
rect 5604 21939 5613 21973
rect 5561 21930 5613 21939
rect 5671 21883 5723 21892
rect 5671 21849 5680 21883
rect 5680 21849 5714 21883
rect 5714 21849 5723 21883
rect 5671 21840 5723 21849
rect 7038 22518 7090 22570
rect 7310 22518 7362 22570
rect 6224 22109 6276 22161
rect 6656 22109 6708 22161
rect 7038 22123 7090 22175
rect 7310 22123 7362 22175
rect 5799 21751 5851 21803
rect 6224 21751 6276 21803
rect 6656 21751 6708 21803
rect 5671 21659 5723 21668
rect 5671 21625 5680 21659
rect 5680 21625 5714 21659
rect 5714 21625 5723 21659
rect 5671 21616 5723 21625
rect 5561 21569 5613 21578
rect 5561 21535 5570 21569
rect 5570 21535 5604 21569
rect 5604 21535 5613 21569
rect 5561 21526 5613 21535
rect 5671 21457 5723 21466
rect 5671 21423 5680 21457
rect 5680 21423 5714 21457
rect 5714 21423 5723 21457
rect 5671 21414 5723 21423
rect 5799 21377 5851 21429
rect 5671 21295 5723 21304
rect 5671 21261 5680 21295
rect 5680 21261 5714 21295
rect 5714 21261 5723 21295
rect 5671 21252 5723 21261
rect 5561 21183 5613 21192
rect 5561 21149 5570 21183
rect 5570 21149 5604 21183
rect 5604 21149 5613 21183
rect 5561 21140 5613 21149
rect 5671 21093 5723 21102
rect 5671 21059 5680 21093
rect 5680 21059 5714 21093
rect 5714 21059 5723 21093
rect 5671 21050 5723 21059
rect 7038 21728 7090 21780
rect 7310 21728 7362 21780
rect 6224 21319 6276 21371
rect 6656 21319 6708 21371
rect 7038 21333 7090 21385
rect 7310 21333 7362 21385
rect 5799 20961 5851 21013
rect 6224 20961 6276 21013
rect 6656 20961 6708 21013
rect 5671 20869 5723 20878
rect 5671 20835 5680 20869
rect 5680 20835 5714 20869
rect 5714 20835 5723 20869
rect 5671 20826 5723 20835
rect 5561 20779 5613 20788
rect 5561 20745 5570 20779
rect 5570 20745 5604 20779
rect 5604 20745 5613 20779
rect 5561 20736 5613 20745
rect 5671 20667 5723 20676
rect 5671 20633 5680 20667
rect 5680 20633 5714 20667
rect 5714 20633 5723 20667
rect 5671 20624 5723 20633
rect 5799 20587 5851 20639
rect 5671 20505 5723 20514
rect 5671 20471 5680 20505
rect 5680 20471 5714 20505
rect 5714 20471 5723 20505
rect 5671 20462 5723 20471
rect 5561 20393 5613 20402
rect 5561 20359 5570 20393
rect 5570 20359 5604 20393
rect 5604 20359 5613 20393
rect 5561 20350 5613 20359
rect 5671 20303 5723 20312
rect 5671 20269 5680 20303
rect 5680 20269 5714 20303
rect 5714 20269 5723 20303
rect 5671 20260 5723 20269
rect 7038 20938 7090 20990
rect 7310 20938 7362 20990
rect 6224 20529 6276 20581
rect 6656 20529 6708 20581
rect 7038 20543 7090 20595
rect 7310 20543 7362 20595
rect 5799 20171 5851 20223
rect 6224 20171 6276 20223
rect 6656 20171 6708 20223
rect 5671 20079 5723 20088
rect 5671 20045 5680 20079
rect 5680 20045 5714 20079
rect 5714 20045 5723 20079
rect 5671 20036 5723 20045
rect 5561 19989 5613 19998
rect 5561 19955 5570 19989
rect 5570 19955 5604 19989
rect 5604 19955 5613 19989
rect 5561 19946 5613 19955
rect 5671 19877 5723 19886
rect 5671 19843 5680 19877
rect 5680 19843 5714 19877
rect 5714 19843 5723 19877
rect 5671 19834 5723 19843
rect 5799 19797 5851 19849
rect 5671 19715 5723 19724
rect 5671 19681 5680 19715
rect 5680 19681 5714 19715
rect 5714 19681 5723 19715
rect 5671 19672 5723 19681
rect 5561 19603 5613 19612
rect 5561 19569 5570 19603
rect 5570 19569 5604 19603
rect 5604 19569 5613 19603
rect 5561 19560 5613 19569
rect 5671 19513 5723 19522
rect 5671 19479 5680 19513
rect 5680 19479 5714 19513
rect 5714 19479 5723 19513
rect 5671 19470 5723 19479
rect 7038 20148 7090 20200
rect 7310 20148 7362 20200
rect 6224 19739 6276 19791
rect 6656 19739 6708 19791
rect 7038 19753 7090 19805
rect 7310 19753 7362 19805
rect 5799 19381 5851 19433
rect 6224 19381 6276 19433
rect 6656 19381 6708 19433
rect 5671 19289 5723 19298
rect 5671 19255 5680 19289
rect 5680 19255 5714 19289
rect 5714 19255 5723 19289
rect 5671 19246 5723 19255
rect 5561 19199 5613 19208
rect 5561 19165 5570 19199
rect 5570 19165 5604 19199
rect 5604 19165 5613 19199
rect 5561 19156 5613 19165
rect 5671 19087 5723 19096
rect 5671 19053 5680 19087
rect 5680 19053 5714 19087
rect 5714 19053 5723 19087
rect 5671 19044 5723 19053
rect 5799 19007 5851 19059
rect 5671 18925 5723 18934
rect 5671 18891 5680 18925
rect 5680 18891 5714 18925
rect 5714 18891 5723 18925
rect 5671 18882 5723 18891
rect 5561 18813 5613 18822
rect 5561 18779 5570 18813
rect 5570 18779 5604 18813
rect 5604 18779 5613 18813
rect 5561 18770 5613 18779
rect 5671 18723 5723 18732
rect 5671 18689 5680 18723
rect 5680 18689 5714 18723
rect 5714 18689 5723 18723
rect 5671 18680 5723 18689
rect 7038 19358 7090 19410
rect 7310 19358 7362 19410
rect 6224 18949 6276 19001
rect 6656 18949 6708 19001
rect 7038 18963 7090 19015
rect 7310 18963 7362 19015
rect 5799 18591 5851 18643
rect 6224 18591 6276 18643
rect 6656 18591 6708 18643
rect 5671 18499 5723 18508
rect 5671 18465 5680 18499
rect 5680 18465 5714 18499
rect 5714 18465 5723 18499
rect 5671 18456 5723 18465
rect 5561 18409 5613 18418
rect 5561 18375 5570 18409
rect 5570 18375 5604 18409
rect 5604 18375 5613 18409
rect 5561 18366 5613 18375
rect 5671 18297 5723 18306
rect 5671 18263 5680 18297
rect 5680 18263 5714 18297
rect 5714 18263 5723 18297
rect 5671 18254 5723 18263
rect 5799 18217 5851 18269
rect 5671 18135 5723 18144
rect 5671 18101 5680 18135
rect 5680 18101 5714 18135
rect 5714 18101 5723 18135
rect 5671 18092 5723 18101
rect 5561 18023 5613 18032
rect 5561 17989 5570 18023
rect 5570 17989 5604 18023
rect 5604 17989 5613 18023
rect 5561 17980 5613 17989
rect 5671 17933 5723 17942
rect 5671 17899 5680 17933
rect 5680 17899 5714 17933
rect 5714 17899 5723 17933
rect 5671 17890 5723 17899
rect 7038 18568 7090 18620
rect 7310 18568 7362 18620
rect 6224 18159 6276 18211
rect 6656 18159 6708 18211
rect 7038 18173 7090 18225
rect 7310 18173 7362 18225
rect 5799 17801 5851 17853
rect 6224 17801 6276 17853
rect 6656 17801 6708 17853
rect 5671 17709 5723 17718
rect 5671 17675 5680 17709
rect 5680 17675 5714 17709
rect 5714 17675 5723 17709
rect 5671 17666 5723 17675
rect 5561 17619 5613 17628
rect 5561 17585 5570 17619
rect 5570 17585 5604 17619
rect 5604 17585 5613 17619
rect 5561 17576 5613 17585
rect 5671 17507 5723 17516
rect 5671 17473 5680 17507
rect 5680 17473 5714 17507
rect 5714 17473 5723 17507
rect 5671 17464 5723 17473
rect 5799 17427 5851 17479
rect 5671 17345 5723 17354
rect 5671 17311 5680 17345
rect 5680 17311 5714 17345
rect 5714 17311 5723 17345
rect 5671 17302 5723 17311
rect 5561 17233 5613 17242
rect 5561 17199 5570 17233
rect 5570 17199 5604 17233
rect 5604 17199 5613 17233
rect 5561 17190 5613 17199
rect 5671 17143 5723 17152
rect 5671 17109 5680 17143
rect 5680 17109 5714 17143
rect 5714 17109 5723 17143
rect 5671 17100 5723 17109
rect 7038 17778 7090 17830
rect 7310 17778 7362 17830
rect 6224 17369 6276 17421
rect 6656 17369 6708 17421
rect 7038 17383 7090 17435
rect 7310 17383 7362 17435
rect 5799 17011 5851 17063
rect 6224 17011 6276 17063
rect 6656 17011 6708 17063
rect 5671 16919 5723 16928
rect 5671 16885 5680 16919
rect 5680 16885 5714 16919
rect 5714 16885 5723 16919
rect 5671 16876 5723 16885
rect 5561 16829 5613 16838
rect 5561 16795 5570 16829
rect 5570 16795 5604 16829
rect 5604 16795 5613 16829
rect 5561 16786 5613 16795
rect 5671 16717 5723 16726
rect 5671 16683 5680 16717
rect 5680 16683 5714 16717
rect 5714 16683 5723 16717
rect 5671 16674 5723 16683
rect 5799 16637 5851 16689
rect 5671 16555 5723 16564
rect 5671 16521 5680 16555
rect 5680 16521 5714 16555
rect 5714 16521 5723 16555
rect 5671 16512 5723 16521
rect 5561 16443 5613 16452
rect 5561 16409 5570 16443
rect 5570 16409 5604 16443
rect 5604 16409 5613 16443
rect 5561 16400 5613 16409
rect 5671 16353 5723 16362
rect 5671 16319 5680 16353
rect 5680 16319 5714 16353
rect 5714 16319 5723 16353
rect 5671 16310 5723 16319
rect 7038 16988 7090 17040
rect 7310 16988 7362 17040
rect 6224 16579 6276 16631
rect 6656 16579 6708 16631
rect 7038 16593 7090 16645
rect 7310 16593 7362 16645
rect 5799 16221 5851 16273
rect 6224 16221 6276 16273
rect 6656 16221 6708 16273
rect 5671 16129 5723 16138
rect 5671 16095 5680 16129
rect 5680 16095 5714 16129
rect 5714 16095 5723 16129
rect 5671 16086 5723 16095
rect 5561 16039 5613 16048
rect 5561 16005 5570 16039
rect 5570 16005 5604 16039
rect 5604 16005 5613 16039
rect 5561 15996 5613 16005
rect 5671 15927 5723 15936
rect 5671 15893 5680 15927
rect 5680 15893 5714 15927
rect 5714 15893 5723 15927
rect 5671 15884 5723 15893
rect 5799 15847 5851 15899
rect 5671 15765 5723 15774
rect 5671 15731 5680 15765
rect 5680 15731 5714 15765
rect 5714 15731 5723 15765
rect 5671 15722 5723 15731
rect 5561 15653 5613 15662
rect 5561 15619 5570 15653
rect 5570 15619 5604 15653
rect 5604 15619 5613 15653
rect 5561 15610 5613 15619
rect 5671 15563 5723 15572
rect 5671 15529 5680 15563
rect 5680 15529 5714 15563
rect 5714 15529 5723 15563
rect 5671 15520 5723 15529
rect 7038 16198 7090 16250
rect 7310 16198 7362 16250
rect 6224 15789 6276 15841
rect 6656 15789 6708 15841
rect 7038 15803 7090 15855
rect 7310 15803 7362 15855
rect 5799 15431 5851 15483
rect 6224 15431 6276 15483
rect 6656 15431 6708 15483
rect 5671 15339 5723 15348
rect 5671 15305 5680 15339
rect 5680 15305 5714 15339
rect 5714 15305 5723 15339
rect 5671 15296 5723 15305
rect 5561 15249 5613 15258
rect 5561 15215 5570 15249
rect 5570 15215 5604 15249
rect 5604 15215 5613 15249
rect 5561 15206 5613 15215
rect 5671 15137 5723 15146
rect 5671 15103 5680 15137
rect 5680 15103 5714 15137
rect 5714 15103 5723 15137
rect 5671 15094 5723 15103
rect 5799 15057 5851 15109
rect 5671 14975 5723 14984
rect 5671 14941 5680 14975
rect 5680 14941 5714 14975
rect 5714 14941 5723 14975
rect 5671 14932 5723 14941
rect 5561 14863 5613 14872
rect 5561 14829 5570 14863
rect 5570 14829 5604 14863
rect 5604 14829 5613 14863
rect 5561 14820 5613 14829
rect 5671 14773 5723 14782
rect 5671 14739 5680 14773
rect 5680 14739 5714 14773
rect 5714 14739 5723 14773
rect 5671 14730 5723 14739
rect 7038 15408 7090 15460
rect 7310 15408 7362 15460
rect 6224 14999 6276 15051
rect 6656 14999 6708 15051
rect 7038 15013 7090 15065
rect 7310 15013 7362 15065
rect 5799 14641 5851 14693
rect 6224 14641 6276 14693
rect 6656 14641 6708 14693
rect 5671 14549 5723 14558
rect 5671 14515 5680 14549
rect 5680 14515 5714 14549
rect 5714 14515 5723 14549
rect 5671 14506 5723 14515
rect 5561 14459 5613 14468
rect 5561 14425 5570 14459
rect 5570 14425 5604 14459
rect 5604 14425 5613 14459
rect 5561 14416 5613 14425
rect 5671 14347 5723 14356
rect 5671 14313 5680 14347
rect 5680 14313 5714 14347
rect 5714 14313 5723 14347
rect 5671 14304 5723 14313
rect 5799 14267 5851 14319
rect 5671 14185 5723 14194
rect 5671 14151 5680 14185
rect 5680 14151 5714 14185
rect 5714 14151 5723 14185
rect 5671 14142 5723 14151
rect 5561 14073 5613 14082
rect 5561 14039 5570 14073
rect 5570 14039 5604 14073
rect 5604 14039 5613 14073
rect 5561 14030 5613 14039
rect 5671 13983 5723 13992
rect 5671 13949 5680 13983
rect 5680 13949 5714 13983
rect 5714 13949 5723 13983
rect 5671 13940 5723 13949
rect 7038 14618 7090 14670
rect 7310 14618 7362 14670
rect 6224 14209 6276 14261
rect 6656 14209 6708 14261
rect 7038 14223 7090 14275
rect 7310 14223 7362 14275
rect 5799 13851 5851 13903
rect 6224 13851 6276 13903
rect 6656 13851 6708 13903
rect 5671 13759 5723 13768
rect 5671 13725 5680 13759
rect 5680 13725 5714 13759
rect 5714 13725 5723 13759
rect 5671 13716 5723 13725
rect 5561 13669 5613 13678
rect 5561 13635 5570 13669
rect 5570 13635 5604 13669
rect 5604 13635 5613 13669
rect 5561 13626 5613 13635
rect 5671 13557 5723 13566
rect 5671 13523 5680 13557
rect 5680 13523 5714 13557
rect 5714 13523 5723 13557
rect 5671 13514 5723 13523
rect 5799 13477 5851 13529
rect 5671 13395 5723 13404
rect 5671 13361 5680 13395
rect 5680 13361 5714 13395
rect 5714 13361 5723 13395
rect 5671 13352 5723 13361
rect 5561 13283 5613 13292
rect 5561 13249 5570 13283
rect 5570 13249 5604 13283
rect 5604 13249 5613 13283
rect 5561 13240 5613 13249
rect 5671 13193 5723 13202
rect 5671 13159 5680 13193
rect 5680 13159 5714 13193
rect 5714 13159 5723 13193
rect 5671 13150 5723 13159
rect 7038 13828 7090 13880
rect 7310 13828 7362 13880
rect 6224 13419 6276 13471
rect 6656 13419 6708 13471
rect 7038 13433 7090 13485
rect 7310 13433 7362 13485
rect 5799 13061 5851 13113
rect 6224 13061 6276 13113
rect 6656 13061 6708 13113
rect 5671 12969 5723 12978
rect 5671 12935 5680 12969
rect 5680 12935 5714 12969
rect 5714 12935 5723 12969
rect 5671 12926 5723 12935
rect 5561 12879 5613 12888
rect 5561 12845 5570 12879
rect 5570 12845 5604 12879
rect 5604 12845 5613 12879
rect 5561 12836 5613 12845
rect 5671 12767 5723 12776
rect 5671 12733 5680 12767
rect 5680 12733 5714 12767
rect 5714 12733 5723 12767
rect 5671 12724 5723 12733
rect 5799 12687 5851 12739
rect 5671 12605 5723 12614
rect 5671 12571 5680 12605
rect 5680 12571 5714 12605
rect 5714 12571 5723 12605
rect 5671 12562 5723 12571
rect 5561 12493 5613 12502
rect 5561 12459 5570 12493
rect 5570 12459 5604 12493
rect 5604 12459 5613 12493
rect 5561 12450 5613 12459
rect 5671 12403 5723 12412
rect 5671 12369 5680 12403
rect 5680 12369 5714 12403
rect 5714 12369 5723 12403
rect 5671 12360 5723 12369
rect 7038 13038 7090 13090
rect 7310 13038 7362 13090
rect 6224 12629 6276 12681
rect 6656 12629 6708 12681
rect 7038 12643 7090 12695
rect 7310 12643 7362 12695
rect 5799 12271 5851 12323
rect 6224 12271 6276 12323
rect 6656 12271 6708 12323
rect 5671 12179 5723 12188
rect 5671 12145 5680 12179
rect 5680 12145 5714 12179
rect 5714 12145 5723 12179
rect 5671 12136 5723 12145
rect 5561 12089 5613 12098
rect 5561 12055 5570 12089
rect 5570 12055 5604 12089
rect 5604 12055 5613 12089
rect 5561 12046 5613 12055
rect 5671 11977 5723 11986
rect 5671 11943 5680 11977
rect 5680 11943 5714 11977
rect 5714 11943 5723 11977
rect 5671 11934 5723 11943
rect 5799 11897 5851 11949
rect 5671 11815 5723 11824
rect 5671 11781 5680 11815
rect 5680 11781 5714 11815
rect 5714 11781 5723 11815
rect 5671 11772 5723 11781
rect 5561 11703 5613 11712
rect 5561 11669 5570 11703
rect 5570 11669 5604 11703
rect 5604 11669 5613 11703
rect 5561 11660 5613 11669
rect 5671 11613 5723 11622
rect 5671 11579 5680 11613
rect 5680 11579 5714 11613
rect 5714 11579 5723 11613
rect 5671 11570 5723 11579
rect 7038 12248 7090 12300
rect 7310 12248 7362 12300
rect 6224 11839 6276 11891
rect 6656 11839 6708 11891
rect 7038 11853 7090 11905
rect 7310 11853 7362 11905
rect 5799 11481 5851 11533
rect 6224 11481 6276 11533
rect 6656 11481 6708 11533
rect 5671 11389 5723 11398
rect 5671 11355 5680 11389
rect 5680 11355 5714 11389
rect 5714 11355 5723 11389
rect 5671 11346 5723 11355
rect 5561 11299 5613 11308
rect 5561 11265 5570 11299
rect 5570 11265 5604 11299
rect 5604 11265 5613 11299
rect 5561 11256 5613 11265
rect 5671 11187 5723 11196
rect 5671 11153 5680 11187
rect 5680 11153 5714 11187
rect 5714 11153 5723 11187
rect 5671 11144 5723 11153
rect 5799 11107 5851 11159
rect 5671 11025 5723 11034
rect 5671 10991 5680 11025
rect 5680 10991 5714 11025
rect 5714 10991 5723 11025
rect 5671 10982 5723 10991
rect 5561 10913 5613 10922
rect 5561 10879 5570 10913
rect 5570 10879 5604 10913
rect 5604 10879 5613 10913
rect 5561 10870 5613 10879
rect 5671 10823 5723 10832
rect 5671 10789 5680 10823
rect 5680 10789 5714 10823
rect 5714 10789 5723 10823
rect 5671 10780 5723 10789
rect 7038 11458 7090 11510
rect 7310 11458 7362 11510
rect 6224 11049 6276 11101
rect 6656 11049 6708 11101
rect 7038 11063 7090 11115
rect 7310 11063 7362 11115
rect 5799 10691 5851 10743
rect 6224 10691 6276 10743
rect 6656 10691 6708 10743
rect 5671 10599 5723 10608
rect 5671 10565 5680 10599
rect 5680 10565 5714 10599
rect 5714 10565 5723 10599
rect 5671 10556 5723 10565
rect 5561 10509 5613 10518
rect 5561 10475 5570 10509
rect 5570 10475 5604 10509
rect 5604 10475 5613 10509
rect 5561 10466 5613 10475
rect 5671 10397 5723 10406
rect 5671 10363 5680 10397
rect 5680 10363 5714 10397
rect 5714 10363 5723 10397
rect 5671 10354 5723 10363
rect 5799 10317 5851 10369
rect 5671 10235 5723 10244
rect 5671 10201 5680 10235
rect 5680 10201 5714 10235
rect 5714 10201 5723 10235
rect 5671 10192 5723 10201
rect 5561 10123 5613 10132
rect 5561 10089 5570 10123
rect 5570 10089 5604 10123
rect 5604 10089 5613 10123
rect 5561 10080 5613 10089
rect 5671 10033 5723 10042
rect 5671 9999 5680 10033
rect 5680 9999 5714 10033
rect 5714 9999 5723 10033
rect 5671 9990 5723 9999
rect 7038 10668 7090 10720
rect 7310 10668 7362 10720
rect 6224 10259 6276 10311
rect 6656 10259 6708 10311
rect 7038 10273 7090 10325
rect 7310 10273 7362 10325
rect 5799 9901 5851 9953
rect 6224 9901 6276 9953
rect 6656 9901 6708 9953
rect 5671 9809 5723 9818
rect 5671 9775 5680 9809
rect 5680 9775 5714 9809
rect 5714 9775 5723 9809
rect 5671 9766 5723 9775
rect 5561 9719 5613 9728
rect 5561 9685 5570 9719
rect 5570 9685 5604 9719
rect 5604 9685 5613 9719
rect 5561 9676 5613 9685
rect 5671 9607 5723 9616
rect 5671 9573 5680 9607
rect 5680 9573 5714 9607
rect 5714 9573 5723 9607
rect 5671 9564 5723 9573
rect 5799 9527 5851 9579
rect 5671 9445 5723 9454
rect 5671 9411 5680 9445
rect 5680 9411 5714 9445
rect 5714 9411 5723 9445
rect 5671 9402 5723 9411
rect 5561 9333 5613 9342
rect 5561 9299 5570 9333
rect 5570 9299 5604 9333
rect 5604 9299 5613 9333
rect 5561 9290 5613 9299
rect 5671 9243 5723 9252
rect 5671 9209 5680 9243
rect 5680 9209 5714 9243
rect 5714 9209 5723 9243
rect 5671 9200 5723 9209
rect 7038 9878 7090 9930
rect 7310 9878 7362 9930
rect 6224 9469 6276 9521
rect 6656 9469 6708 9521
rect 7038 9483 7090 9535
rect 7310 9483 7362 9535
rect 5799 9111 5851 9163
rect 6224 9111 6276 9163
rect 6656 9111 6708 9163
rect 5671 9019 5723 9028
rect 5671 8985 5680 9019
rect 5680 8985 5714 9019
rect 5714 8985 5723 9019
rect 5671 8976 5723 8985
rect 5561 8929 5613 8938
rect 5561 8895 5570 8929
rect 5570 8895 5604 8929
rect 5604 8895 5613 8929
rect 5561 8886 5613 8895
rect 5671 8817 5723 8826
rect 5671 8783 5680 8817
rect 5680 8783 5714 8817
rect 5714 8783 5723 8817
rect 5671 8774 5723 8783
rect 5799 8737 5851 8789
rect 5671 8655 5723 8664
rect 5671 8621 5680 8655
rect 5680 8621 5714 8655
rect 5714 8621 5723 8655
rect 5671 8612 5723 8621
rect 5561 8543 5613 8552
rect 5561 8509 5570 8543
rect 5570 8509 5604 8543
rect 5604 8509 5613 8543
rect 5561 8500 5613 8509
rect 5671 8453 5723 8462
rect 5671 8419 5680 8453
rect 5680 8419 5714 8453
rect 5714 8419 5723 8453
rect 5671 8410 5723 8419
rect 7038 9088 7090 9140
rect 7310 9088 7362 9140
rect 6224 8679 6276 8731
rect 6656 8679 6708 8731
rect 7038 8693 7090 8745
rect 7310 8693 7362 8745
rect 5799 8321 5851 8373
rect 6224 8321 6276 8373
rect 6656 8321 6708 8373
rect 5671 8229 5723 8238
rect 5671 8195 5680 8229
rect 5680 8195 5714 8229
rect 5714 8195 5723 8229
rect 5671 8186 5723 8195
rect 5561 8139 5613 8148
rect 5561 8105 5570 8139
rect 5570 8105 5604 8139
rect 5604 8105 5613 8139
rect 5561 8096 5613 8105
rect 5671 8027 5723 8036
rect 5671 7993 5680 8027
rect 5680 7993 5714 8027
rect 5714 7993 5723 8027
rect 5671 7984 5723 7993
rect 5799 7947 5851 7999
rect 5671 7865 5723 7874
rect 5671 7831 5680 7865
rect 5680 7831 5714 7865
rect 5714 7831 5723 7865
rect 5671 7822 5723 7831
rect 5561 7753 5613 7762
rect 5561 7719 5570 7753
rect 5570 7719 5604 7753
rect 5604 7719 5613 7753
rect 5561 7710 5613 7719
rect 5671 7663 5723 7672
rect 5671 7629 5680 7663
rect 5680 7629 5714 7663
rect 5714 7629 5723 7663
rect 5671 7620 5723 7629
rect 7038 8298 7090 8350
rect 7310 8298 7362 8350
rect 6224 7889 6276 7941
rect 6656 7889 6708 7941
rect 7038 7903 7090 7955
rect 7310 7903 7362 7955
rect 5799 7531 5851 7583
rect 6224 7531 6276 7583
rect 6656 7531 6708 7583
rect 4902 5026 4954 5078
rect 4822 4936 4874 4988
rect 4742 4550 4794 4602
rect 4742 4146 4794 4198
rect 4742 3760 4794 3812
rect 4902 4460 4954 4512
rect 4902 4236 4954 4288
rect 4902 3670 4954 3722
rect 4742 3356 4794 3408
rect 4662 2970 4714 3022
rect 4662 2566 4714 2618
rect 4502 1502 4554 1554
rect 4662 2180 4714 2232
rect 4662 1776 4714 1828
rect 4582 1390 4634 1442
rect 4422 874 4474 926
rect 4342 712 4394 764
rect 4262 84 4314 136
rect 4582 986 4634 1038
rect 4582 600 4634 652
rect 4582 196 4634 248
rect 4902 3446 4954 3498
rect 4902 2880 4954 2932
rect 4902 2656 4954 2708
rect 4902 2090 4954 2142
rect 4902 1866 4954 1918
rect 4902 1300 4954 1352
rect 4902 1076 4954 1128
rect 4902 510 4954 562
rect 4902 286 4954 338
rect 5671 7439 5723 7448
rect 5671 7405 5680 7439
rect 5680 7405 5714 7439
rect 5714 7405 5723 7439
rect 5671 7396 5723 7405
rect 5561 7349 5613 7358
rect 5561 7315 5570 7349
rect 5570 7315 5604 7349
rect 5604 7315 5613 7349
rect 5561 7306 5613 7315
rect 5671 7237 5723 7246
rect 5671 7203 5680 7237
rect 5680 7203 5714 7237
rect 5714 7203 5723 7237
rect 5671 7194 5723 7203
rect 5799 7157 5851 7209
rect 5671 7075 5723 7084
rect 5671 7041 5680 7075
rect 5680 7041 5714 7075
rect 5714 7041 5723 7075
rect 5671 7032 5723 7041
rect 5561 6963 5613 6972
rect 5561 6929 5570 6963
rect 5570 6929 5604 6963
rect 5604 6929 5613 6963
rect 5561 6920 5613 6929
rect 5671 6873 5723 6882
rect 5671 6839 5680 6873
rect 5680 6839 5714 6873
rect 5714 6839 5723 6873
rect 5671 6830 5723 6839
rect 7038 7508 7090 7560
rect 7310 7508 7362 7560
rect 6224 7099 6276 7151
rect 6656 7099 6708 7151
rect 7038 7113 7090 7165
rect 7310 7113 7362 7165
rect 5799 6741 5851 6793
rect 6224 6741 6276 6793
rect 6656 6741 6708 6793
rect 5671 6649 5723 6658
rect 5671 6615 5680 6649
rect 5680 6615 5714 6649
rect 5714 6615 5723 6649
rect 5671 6606 5723 6615
rect 5561 6559 5613 6568
rect 5561 6525 5570 6559
rect 5570 6525 5604 6559
rect 5604 6525 5613 6559
rect 5561 6516 5613 6525
rect 5671 6447 5723 6456
rect 5671 6413 5680 6447
rect 5680 6413 5714 6447
rect 5714 6413 5723 6447
rect 5671 6404 5723 6413
rect 5799 6367 5851 6419
rect 5671 6285 5723 6294
rect 5671 6251 5680 6285
rect 5680 6251 5714 6285
rect 5714 6251 5723 6285
rect 5671 6242 5723 6251
rect 5561 6173 5613 6182
rect 5561 6139 5570 6173
rect 5570 6139 5604 6173
rect 5604 6139 5613 6173
rect 5561 6130 5613 6139
rect 5671 6083 5723 6092
rect 5671 6049 5680 6083
rect 5680 6049 5714 6083
rect 5714 6049 5723 6083
rect 5671 6040 5723 6049
rect 7038 6718 7090 6770
rect 7310 6718 7362 6770
rect 6224 6309 6276 6361
rect 6656 6309 6708 6361
rect 7038 6323 7090 6375
rect 7310 6323 7362 6375
rect 5799 5951 5851 6003
rect 6224 5951 6276 6003
rect 6656 5951 6708 6003
rect 5671 5859 5723 5868
rect 5671 5825 5680 5859
rect 5680 5825 5714 5859
rect 5714 5825 5723 5859
rect 5671 5816 5723 5825
rect 5561 5769 5613 5778
rect 5561 5735 5570 5769
rect 5570 5735 5604 5769
rect 5604 5735 5613 5769
rect 5561 5726 5613 5735
rect 5671 5657 5723 5666
rect 5671 5623 5680 5657
rect 5680 5623 5714 5657
rect 5714 5623 5723 5657
rect 5671 5614 5723 5623
rect 5799 5577 5851 5629
rect 5671 5495 5723 5504
rect 5671 5461 5680 5495
rect 5680 5461 5714 5495
rect 5714 5461 5723 5495
rect 5671 5452 5723 5461
rect 5561 5383 5613 5392
rect 5561 5349 5570 5383
rect 5570 5349 5604 5383
rect 5604 5349 5613 5383
rect 5561 5340 5613 5349
rect 5671 5293 5723 5302
rect 5671 5259 5680 5293
rect 5680 5259 5714 5293
rect 5714 5259 5723 5293
rect 5671 5250 5723 5259
rect 7038 5928 7090 5980
rect 7310 5928 7362 5980
rect 6224 5519 6276 5571
rect 6656 5519 6708 5571
rect 7038 5533 7090 5585
rect 7310 5533 7362 5585
rect 5799 5161 5851 5213
rect 6224 5161 6276 5213
rect 6656 5161 6708 5213
rect 5671 5069 5723 5078
rect 5671 5035 5680 5069
rect 5680 5035 5714 5069
rect 5714 5035 5723 5069
rect 5671 5026 5723 5035
rect 5561 4979 5613 4988
rect 5561 4945 5570 4979
rect 5570 4945 5604 4979
rect 5604 4945 5613 4979
rect 5561 4936 5613 4945
rect 5671 4867 5723 4876
rect 5671 4833 5680 4867
rect 5680 4833 5714 4867
rect 5714 4833 5723 4867
rect 5671 4824 5723 4833
rect 5799 4787 5851 4839
rect 5671 4705 5723 4714
rect 5671 4671 5680 4705
rect 5680 4671 5714 4705
rect 5714 4671 5723 4705
rect 5671 4662 5723 4671
rect 5561 4593 5613 4602
rect 5561 4559 5570 4593
rect 5570 4559 5604 4593
rect 5604 4559 5613 4593
rect 5561 4550 5613 4559
rect 5671 4503 5723 4512
rect 5671 4469 5680 4503
rect 5680 4469 5714 4503
rect 5714 4469 5723 4503
rect 5671 4460 5723 4469
rect 7038 5138 7090 5190
rect 7310 5138 7362 5190
rect 6224 4729 6276 4781
rect 6656 4729 6708 4781
rect 7038 4743 7090 4795
rect 7310 4743 7362 4795
rect 5799 4371 5851 4423
rect 6224 4371 6276 4423
rect 6656 4371 6708 4423
rect 5671 4279 5723 4288
rect 5671 4245 5680 4279
rect 5680 4245 5714 4279
rect 5714 4245 5723 4279
rect 5671 4236 5723 4245
rect 5561 4189 5613 4198
rect 5561 4155 5570 4189
rect 5570 4155 5604 4189
rect 5604 4155 5613 4189
rect 5561 4146 5613 4155
rect 5671 4077 5723 4086
rect 5671 4043 5680 4077
rect 5680 4043 5714 4077
rect 5714 4043 5723 4077
rect 5671 4034 5723 4043
rect 5799 3997 5851 4049
rect 5671 3915 5723 3924
rect 5671 3881 5680 3915
rect 5680 3881 5714 3915
rect 5714 3881 5723 3915
rect 5671 3872 5723 3881
rect 5561 3803 5613 3812
rect 5561 3769 5570 3803
rect 5570 3769 5604 3803
rect 5604 3769 5613 3803
rect 5561 3760 5613 3769
rect 5671 3713 5723 3722
rect 5671 3679 5680 3713
rect 5680 3679 5714 3713
rect 5714 3679 5723 3713
rect 5671 3670 5723 3679
rect 7038 4348 7090 4400
rect 7310 4348 7362 4400
rect 6224 3939 6276 3991
rect 6656 3939 6708 3991
rect 7038 3953 7090 4005
rect 7310 3953 7362 4005
rect 5799 3581 5851 3633
rect 6224 3581 6276 3633
rect 6656 3581 6708 3633
rect 5671 3489 5723 3498
rect 5671 3455 5680 3489
rect 5680 3455 5714 3489
rect 5714 3455 5723 3489
rect 5671 3446 5723 3455
rect 5561 3399 5613 3408
rect 5561 3365 5570 3399
rect 5570 3365 5604 3399
rect 5604 3365 5613 3399
rect 5561 3356 5613 3365
rect 5671 3287 5723 3296
rect 5671 3253 5680 3287
rect 5680 3253 5714 3287
rect 5714 3253 5723 3287
rect 5671 3244 5723 3253
rect 5799 3207 5851 3259
rect 5671 3125 5723 3134
rect 5671 3091 5680 3125
rect 5680 3091 5714 3125
rect 5714 3091 5723 3125
rect 5671 3082 5723 3091
rect 5561 3013 5613 3022
rect 5561 2979 5570 3013
rect 5570 2979 5604 3013
rect 5604 2979 5613 3013
rect 5561 2970 5613 2979
rect 5671 2923 5723 2932
rect 5671 2889 5680 2923
rect 5680 2889 5714 2923
rect 5714 2889 5723 2923
rect 5671 2880 5723 2889
rect 7038 3558 7090 3610
rect 7310 3558 7362 3610
rect 6224 3149 6276 3201
rect 6656 3149 6708 3201
rect 7038 3163 7090 3215
rect 7310 3163 7362 3215
rect 5799 2791 5851 2843
rect 6224 2791 6276 2843
rect 6656 2791 6708 2843
rect 5671 2699 5723 2708
rect 5671 2665 5680 2699
rect 5680 2665 5714 2699
rect 5714 2665 5723 2699
rect 5671 2656 5723 2665
rect 5561 2609 5613 2618
rect 5561 2575 5570 2609
rect 5570 2575 5604 2609
rect 5604 2575 5613 2609
rect 5561 2566 5613 2575
rect 5671 2497 5723 2506
rect 5671 2463 5680 2497
rect 5680 2463 5714 2497
rect 5714 2463 5723 2497
rect 5671 2454 5723 2463
rect 5799 2417 5851 2469
rect 5671 2335 5723 2344
rect 5671 2301 5680 2335
rect 5680 2301 5714 2335
rect 5714 2301 5723 2335
rect 5671 2292 5723 2301
rect 5561 2223 5613 2232
rect 5561 2189 5570 2223
rect 5570 2189 5604 2223
rect 5604 2189 5613 2223
rect 5561 2180 5613 2189
rect 5671 2133 5723 2142
rect 5671 2099 5680 2133
rect 5680 2099 5714 2133
rect 5714 2099 5723 2133
rect 5671 2090 5723 2099
rect 7038 2768 7090 2820
rect 7310 2768 7362 2820
rect 6224 2359 6276 2411
rect 6656 2359 6708 2411
rect 7038 2373 7090 2425
rect 7310 2373 7362 2425
rect 5799 2001 5851 2053
rect 6224 2001 6276 2053
rect 6656 2001 6708 2053
rect 5671 1909 5723 1918
rect 5671 1875 5680 1909
rect 5680 1875 5714 1909
rect 5714 1875 5723 1909
rect 5671 1866 5723 1875
rect 5561 1819 5613 1828
rect 5561 1785 5570 1819
rect 5570 1785 5604 1819
rect 5604 1785 5613 1819
rect 5561 1776 5613 1785
rect 5671 1707 5723 1716
rect 5671 1673 5680 1707
rect 5680 1673 5714 1707
rect 5714 1673 5723 1707
rect 5671 1664 5723 1673
rect 5799 1627 5851 1679
rect 5671 1545 5723 1554
rect 5671 1511 5680 1545
rect 5680 1511 5714 1545
rect 5714 1511 5723 1545
rect 5671 1502 5723 1511
rect 5561 1433 5613 1442
rect 5561 1399 5570 1433
rect 5570 1399 5604 1433
rect 5604 1399 5613 1433
rect 5561 1390 5613 1399
rect 5671 1343 5723 1352
rect 5671 1309 5680 1343
rect 5680 1309 5714 1343
rect 5714 1309 5723 1343
rect 5671 1300 5723 1309
rect 7038 1978 7090 2030
rect 7310 1978 7362 2030
rect 6224 1569 6276 1621
rect 6656 1569 6708 1621
rect 7038 1583 7090 1635
rect 7310 1583 7362 1635
rect 5799 1211 5851 1263
rect 6224 1211 6276 1263
rect 6656 1211 6708 1263
rect 5671 1119 5723 1128
rect 5671 1085 5680 1119
rect 5680 1085 5714 1119
rect 5714 1085 5723 1119
rect 5671 1076 5723 1085
rect 5561 1029 5613 1038
rect 5561 995 5570 1029
rect 5570 995 5604 1029
rect 5604 995 5613 1029
rect 5561 986 5613 995
rect 5671 917 5723 926
rect 5671 883 5680 917
rect 5680 883 5714 917
rect 5714 883 5723 917
rect 5671 874 5723 883
rect 5799 837 5851 889
rect 5671 755 5723 764
rect 5671 721 5680 755
rect 5680 721 5714 755
rect 5714 721 5723 755
rect 5671 712 5723 721
rect 5561 643 5613 652
rect 5561 609 5570 643
rect 5570 609 5604 643
rect 5604 609 5613 643
rect 5561 600 5613 609
rect 5671 553 5723 562
rect 5671 519 5680 553
rect 5680 519 5714 553
rect 5714 519 5723 553
rect 5671 510 5723 519
rect 7038 1188 7090 1240
rect 7310 1188 7362 1240
rect 6224 779 6276 831
rect 6656 779 6708 831
rect 7038 793 7090 845
rect 7310 793 7362 845
rect 5799 421 5851 473
rect 6224 421 6276 473
rect 6656 421 6708 473
rect 5671 329 5723 338
rect 5671 295 5680 329
rect 5680 295 5714 329
rect 5714 295 5723 329
rect 5671 286 5723 295
rect 5561 239 5613 248
rect 5561 205 5570 239
rect 5570 205 5604 239
rect 5604 205 5613 239
rect 5561 196 5613 205
rect 5671 127 5723 136
rect 5671 93 5680 127
rect 5680 93 5714 127
rect 5714 93 5723 127
rect 5671 84 5723 93
rect 7038 398 7090 450
rect 7310 398 7362 450
<< metal2 >>
rect 4496 50482 4502 50534
rect 4554 50522 4560 50534
rect 5665 50522 5671 50534
rect 4554 50494 5671 50522
rect 4554 50482 4560 50494
rect 5665 50482 5671 50494
rect 5723 50482 5729 50534
rect 4816 50370 4822 50422
rect 4874 50410 4880 50422
rect 5555 50410 5561 50422
rect 4874 50382 5561 50410
rect 4874 50370 4880 50382
rect 5555 50370 5561 50382
rect 5613 50370 5619 50422
rect 5456 50280 5462 50332
rect 5514 50320 5520 50332
rect 5665 50320 5671 50332
rect 5514 50292 5671 50320
rect 5514 50280 5520 50292
rect 5665 50280 5671 50292
rect 5723 50280 5729 50332
rect 5797 50245 5853 50254
rect 5797 50180 5853 50189
rect 6222 50245 6278 50254
rect 6222 50180 6278 50189
rect 6654 50245 6710 50254
rect 6654 50180 6710 50189
rect 7036 50222 7092 50231
rect 7036 50157 7092 50166
rect 7308 50222 7364 50231
rect 7308 50157 7364 50166
rect 5456 50056 5462 50108
rect 5514 50096 5520 50108
rect 5665 50096 5671 50108
rect 5514 50068 5671 50096
rect 5514 50056 5520 50068
rect 5665 50056 5671 50068
rect 5723 50056 5729 50108
rect 4816 49966 4822 50018
rect 4874 50006 4880 50018
rect 5555 50006 5561 50018
rect 4874 49978 5561 50006
rect 4874 49966 4880 49978
rect 5555 49966 5561 49978
rect 5613 49966 5619 50018
rect 4416 49854 4422 49906
rect 4474 49894 4480 49906
rect 5665 49894 5671 49906
rect 4474 49866 5671 49894
rect 4474 49854 4480 49866
rect 5665 49854 5671 49866
rect 5723 49854 5729 49906
rect 5797 49871 5853 49880
rect 7036 49827 7092 49836
rect 5797 49806 5853 49815
rect 6222 49813 6278 49822
rect 6222 49748 6278 49757
rect 6654 49813 6710 49822
rect 7036 49762 7092 49771
rect 7308 49827 7364 49836
rect 7308 49762 7364 49771
rect 6654 49748 6710 49757
rect 4336 49692 4342 49744
rect 4394 49732 4400 49744
rect 5665 49732 5671 49744
rect 4394 49704 5671 49732
rect 4394 49692 4400 49704
rect 5665 49692 5671 49704
rect 5723 49692 5729 49744
rect 4816 49580 4822 49632
rect 4874 49620 4880 49632
rect 5555 49620 5561 49632
rect 4874 49592 5561 49620
rect 4874 49580 4880 49592
rect 5555 49580 5561 49592
rect 5613 49580 5619 49632
rect 5456 49490 5462 49542
rect 5514 49530 5520 49542
rect 5665 49530 5671 49542
rect 5514 49502 5671 49530
rect 5514 49490 5520 49502
rect 5665 49490 5671 49502
rect 5723 49490 5729 49542
rect 5797 49455 5853 49464
rect 5797 49390 5853 49399
rect 6222 49455 6278 49464
rect 6222 49390 6278 49399
rect 6654 49455 6710 49464
rect 6654 49390 6710 49399
rect 7036 49432 7092 49441
rect 7036 49367 7092 49376
rect 7308 49432 7364 49441
rect 7308 49367 7364 49376
rect 5456 49266 5462 49318
rect 5514 49306 5520 49318
rect 5665 49306 5671 49318
rect 5514 49278 5671 49306
rect 5514 49266 5520 49278
rect 5665 49266 5671 49278
rect 5723 49266 5729 49318
rect 4816 49176 4822 49228
rect 4874 49216 4880 49228
rect 5555 49216 5561 49228
rect 4874 49188 5561 49216
rect 4874 49176 4880 49188
rect 5555 49176 5561 49188
rect 5613 49176 5619 49228
rect 4256 49064 4262 49116
rect 4314 49104 4320 49116
rect 5665 49104 5671 49116
rect 4314 49076 5671 49104
rect 4314 49064 4320 49076
rect 5665 49064 5671 49076
rect 5723 49064 5729 49116
rect 5797 49081 5853 49090
rect 7036 49037 7092 49046
rect 5797 49016 5853 49025
rect 6222 49023 6278 49032
rect 6222 48958 6278 48967
rect 6654 49023 6710 49032
rect 7036 48972 7092 48981
rect 7308 49037 7364 49046
rect 7308 48972 7364 48981
rect 6654 48958 6710 48967
rect 4496 48902 4502 48954
rect 4554 48942 4560 48954
rect 5665 48942 5671 48954
rect 4554 48914 5671 48942
rect 4554 48902 4560 48914
rect 5665 48902 5671 48914
rect 5723 48902 5729 48954
rect 4736 48790 4742 48842
rect 4794 48830 4800 48842
rect 5555 48830 5561 48842
rect 4794 48802 5561 48830
rect 4794 48790 4800 48802
rect 5555 48790 5561 48802
rect 5613 48790 5619 48842
rect 5456 48700 5462 48752
rect 5514 48740 5520 48752
rect 5665 48740 5671 48752
rect 5514 48712 5671 48740
rect 5514 48700 5520 48712
rect 5665 48700 5671 48712
rect 5723 48700 5729 48752
rect 5797 48665 5853 48674
rect 5797 48600 5853 48609
rect 6222 48665 6278 48674
rect 6222 48600 6278 48609
rect 6654 48665 6710 48674
rect 6654 48600 6710 48609
rect 7036 48642 7092 48651
rect 7036 48577 7092 48586
rect 7308 48642 7364 48651
rect 7308 48577 7364 48586
rect 5456 48476 5462 48528
rect 5514 48516 5520 48528
rect 5665 48516 5671 48528
rect 5514 48488 5671 48516
rect 5514 48476 5520 48488
rect 5665 48476 5671 48488
rect 5723 48476 5729 48528
rect 4736 48386 4742 48438
rect 4794 48426 4800 48438
rect 5555 48426 5561 48438
rect 4794 48398 5561 48426
rect 4794 48386 4800 48398
rect 5555 48386 5561 48398
rect 5613 48386 5619 48438
rect 4416 48274 4422 48326
rect 4474 48314 4480 48326
rect 5665 48314 5671 48326
rect 4474 48286 5671 48314
rect 4474 48274 4480 48286
rect 5665 48274 5671 48286
rect 5723 48274 5729 48326
rect 5797 48291 5853 48300
rect 7036 48247 7092 48256
rect 5797 48226 5853 48235
rect 6222 48233 6278 48242
rect 6222 48168 6278 48177
rect 6654 48233 6710 48242
rect 7036 48182 7092 48191
rect 7308 48247 7364 48256
rect 7308 48182 7364 48191
rect 6654 48168 6710 48177
rect 4336 48112 4342 48164
rect 4394 48152 4400 48164
rect 5665 48152 5671 48164
rect 4394 48124 5671 48152
rect 4394 48112 4400 48124
rect 5665 48112 5671 48124
rect 5723 48112 5729 48164
rect 4736 48000 4742 48052
rect 4794 48040 4800 48052
rect 5555 48040 5561 48052
rect 4794 48012 5561 48040
rect 4794 48000 4800 48012
rect 5555 48000 5561 48012
rect 5613 48000 5619 48052
rect 5456 47910 5462 47962
rect 5514 47950 5520 47962
rect 5665 47950 5671 47962
rect 5514 47922 5671 47950
rect 5514 47910 5520 47922
rect 5665 47910 5671 47922
rect 5723 47910 5729 47962
rect 5797 47875 5853 47884
rect 5797 47810 5853 47819
rect 6222 47875 6278 47884
rect 6222 47810 6278 47819
rect 6654 47875 6710 47884
rect 6654 47810 6710 47819
rect 7036 47852 7092 47861
rect 7036 47787 7092 47796
rect 7308 47852 7364 47861
rect 7308 47787 7364 47796
rect 5456 47686 5462 47738
rect 5514 47726 5520 47738
rect 5665 47726 5671 47738
rect 5514 47698 5671 47726
rect 5514 47686 5520 47698
rect 5665 47686 5671 47698
rect 5723 47686 5729 47738
rect 4736 47596 4742 47648
rect 4794 47636 4800 47648
rect 5555 47636 5561 47648
rect 4794 47608 5561 47636
rect 4794 47596 4800 47608
rect 5555 47596 5561 47608
rect 5613 47596 5619 47648
rect 4256 47484 4262 47536
rect 4314 47524 4320 47536
rect 5665 47524 5671 47536
rect 4314 47496 5671 47524
rect 4314 47484 4320 47496
rect 5665 47484 5671 47496
rect 5723 47484 5729 47536
rect 5797 47501 5853 47510
rect 7036 47457 7092 47466
rect 5797 47436 5853 47445
rect 6222 47443 6278 47452
rect 6222 47378 6278 47387
rect 6654 47443 6710 47452
rect 7036 47392 7092 47401
rect 7308 47457 7364 47466
rect 7308 47392 7364 47401
rect 6654 47378 6710 47387
rect 4496 47322 4502 47374
rect 4554 47362 4560 47374
rect 5665 47362 5671 47374
rect 4554 47334 5671 47362
rect 4554 47322 4560 47334
rect 5665 47322 5671 47334
rect 5723 47322 5729 47374
rect 4656 47210 4662 47262
rect 4714 47250 4720 47262
rect 5555 47250 5561 47262
rect 4714 47222 5561 47250
rect 4714 47210 4720 47222
rect 5555 47210 5561 47222
rect 5613 47210 5619 47262
rect 5456 47120 5462 47172
rect 5514 47160 5520 47172
rect 5665 47160 5671 47172
rect 5514 47132 5671 47160
rect 5514 47120 5520 47132
rect 5665 47120 5671 47132
rect 5723 47120 5729 47172
rect 5797 47085 5853 47094
rect 5797 47020 5853 47029
rect 6222 47085 6278 47094
rect 6222 47020 6278 47029
rect 6654 47085 6710 47094
rect 6654 47020 6710 47029
rect 7036 47062 7092 47071
rect 7036 46997 7092 47006
rect 7308 47062 7364 47071
rect 7308 46997 7364 47006
rect 5456 46896 5462 46948
rect 5514 46936 5520 46948
rect 5665 46936 5671 46948
rect 5514 46908 5671 46936
rect 5514 46896 5520 46908
rect 5665 46896 5671 46908
rect 5723 46896 5729 46948
rect 4656 46806 4662 46858
rect 4714 46846 4720 46858
rect 5555 46846 5561 46858
rect 4714 46818 5561 46846
rect 4714 46806 4720 46818
rect 5555 46806 5561 46818
rect 5613 46806 5619 46858
rect 4416 46694 4422 46746
rect 4474 46734 4480 46746
rect 5665 46734 5671 46746
rect 4474 46706 5671 46734
rect 4474 46694 4480 46706
rect 5665 46694 5671 46706
rect 5723 46694 5729 46746
rect 5797 46711 5853 46720
rect 7036 46667 7092 46676
rect 5797 46646 5853 46655
rect 6222 46653 6278 46662
rect 6222 46588 6278 46597
rect 6654 46653 6710 46662
rect 7036 46602 7092 46611
rect 7308 46667 7364 46676
rect 7308 46602 7364 46611
rect 6654 46588 6710 46597
rect 4336 46532 4342 46584
rect 4394 46572 4400 46584
rect 5665 46572 5671 46584
rect 4394 46544 5671 46572
rect 4394 46532 4400 46544
rect 5665 46532 5671 46544
rect 5723 46532 5729 46584
rect 4656 46420 4662 46472
rect 4714 46460 4720 46472
rect 5555 46460 5561 46472
rect 4714 46432 5561 46460
rect 4714 46420 4720 46432
rect 5555 46420 5561 46432
rect 5613 46420 5619 46472
rect 5456 46330 5462 46382
rect 5514 46370 5520 46382
rect 5665 46370 5671 46382
rect 5514 46342 5671 46370
rect 5514 46330 5520 46342
rect 5665 46330 5671 46342
rect 5723 46330 5729 46382
rect 5797 46295 5853 46304
rect 5797 46230 5853 46239
rect 6222 46295 6278 46304
rect 6222 46230 6278 46239
rect 6654 46295 6710 46304
rect 6654 46230 6710 46239
rect 7036 46272 7092 46281
rect 7036 46207 7092 46216
rect 7308 46272 7364 46281
rect 7308 46207 7364 46216
rect 5456 46106 5462 46158
rect 5514 46146 5520 46158
rect 5665 46146 5671 46158
rect 5514 46118 5671 46146
rect 5514 46106 5520 46118
rect 5665 46106 5671 46118
rect 5723 46106 5729 46158
rect 4656 46016 4662 46068
rect 4714 46056 4720 46068
rect 5555 46056 5561 46068
rect 4714 46028 5561 46056
rect 4714 46016 4720 46028
rect 5555 46016 5561 46028
rect 5613 46016 5619 46068
rect 4256 45904 4262 45956
rect 4314 45944 4320 45956
rect 5665 45944 5671 45956
rect 4314 45916 5671 45944
rect 4314 45904 4320 45916
rect 5665 45904 5671 45916
rect 5723 45904 5729 45956
rect 5797 45921 5853 45930
rect 7036 45877 7092 45886
rect 5797 45856 5853 45865
rect 6222 45863 6278 45872
rect 6222 45798 6278 45807
rect 6654 45863 6710 45872
rect 7036 45812 7092 45821
rect 7308 45877 7364 45886
rect 7308 45812 7364 45821
rect 6654 45798 6710 45807
rect 4496 45742 4502 45794
rect 4554 45782 4560 45794
rect 5665 45782 5671 45794
rect 4554 45754 5671 45782
rect 4554 45742 4560 45754
rect 5665 45742 5671 45754
rect 5723 45742 5729 45794
rect 4576 45630 4582 45682
rect 4634 45670 4640 45682
rect 5555 45670 5561 45682
rect 4634 45642 5561 45670
rect 4634 45630 4640 45642
rect 5555 45630 5561 45642
rect 5613 45630 5619 45682
rect 5456 45540 5462 45592
rect 5514 45580 5520 45592
rect 5665 45580 5671 45592
rect 5514 45552 5671 45580
rect 5514 45540 5520 45552
rect 5665 45540 5671 45552
rect 5723 45540 5729 45592
rect 5797 45505 5853 45514
rect 5797 45440 5853 45449
rect 6222 45505 6278 45514
rect 6222 45440 6278 45449
rect 6654 45505 6710 45514
rect 6654 45440 6710 45449
rect 7036 45482 7092 45491
rect 7036 45417 7092 45426
rect 7308 45482 7364 45491
rect 7308 45417 7364 45426
rect 5456 45316 5462 45368
rect 5514 45356 5520 45368
rect 5665 45356 5671 45368
rect 5514 45328 5671 45356
rect 5514 45316 5520 45328
rect 5665 45316 5671 45328
rect 5723 45316 5729 45368
rect 4576 45226 4582 45278
rect 4634 45266 4640 45278
rect 5555 45266 5561 45278
rect 4634 45238 5561 45266
rect 4634 45226 4640 45238
rect 5555 45226 5561 45238
rect 5613 45226 5619 45278
rect 4416 45114 4422 45166
rect 4474 45154 4480 45166
rect 5665 45154 5671 45166
rect 4474 45126 5671 45154
rect 4474 45114 4480 45126
rect 5665 45114 5671 45126
rect 5723 45114 5729 45166
rect 5797 45131 5853 45140
rect 7036 45087 7092 45096
rect 5797 45066 5853 45075
rect 6222 45073 6278 45082
rect 6222 45008 6278 45017
rect 6654 45073 6710 45082
rect 7036 45022 7092 45031
rect 7308 45087 7364 45096
rect 7308 45022 7364 45031
rect 6654 45008 6710 45017
rect 4336 44952 4342 45004
rect 4394 44992 4400 45004
rect 5665 44992 5671 45004
rect 4394 44964 5671 44992
rect 4394 44952 4400 44964
rect 5665 44952 5671 44964
rect 5723 44952 5729 45004
rect 4576 44840 4582 44892
rect 4634 44880 4640 44892
rect 5555 44880 5561 44892
rect 4634 44852 5561 44880
rect 4634 44840 4640 44852
rect 5555 44840 5561 44852
rect 5613 44840 5619 44892
rect 5456 44750 5462 44802
rect 5514 44790 5520 44802
rect 5665 44790 5671 44802
rect 5514 44762 5671 44790
rect 5514 44750 5520 44762
rect 5665 44750 5671 44762
rect 5723 44750 5729 44802
rect 5797 44715 5853 44724
rect 5797 44650 5853 44659
rect 6222 44715 6278 44724
rect 6222 44650 6278 44659
rect 6654 44715 6710 44724
rect 6654 44650 6710 44659
rect 7036 44692 7092 44701
rect 7036 44627 7092 44636
rect 7308 44692 7364 44701
rect 7308 44627 7364 44636
rect 5456 44526 5462 44578
rect 5514 44566 5520 44578
rect 5665 44566 5671 44578
rect 5514 44538 5671 44566
rect 5514 44526 5520 44538
rect 5665 44526 5671 44538
rect 5723 44526 5729 44578
rect 4576 44436 4582 44488
rect 4634 44476 4640 44488
rect 5555 44476 5561 44488
rect 4634 44448 5561 44476
rect 4634 44436 4640 44448
rect 5555 44436 5561 44448
rect 5613 44436 5619 44488
rect 4256 44324 4262 44376
rect 4314 44364 4320 44376
rect 5665 44364 5671 44376
rect 4314 44336 5671 44364
rect 4314 44324 4320 44336
rect 5665 44324 5671 44336
rect 5723 44324 5729 44376
rect 5797 44341 5853 44350
rect 7036 44297 7092 44306
rect 5797 44276 5853 44285
rect 6222 44283 6278 44292
rect 6222 44218 6278 44227
rect 6654 44283 6710 44292
rect 7036 44232 7092 44241
rect 7308 44297 7364 44306
rect 7308 44232 7364 44241
rect 6654 44218 6710 44227
rect 4496 44162 4502 44214
rect 4554 44202 4560 44214
rect 5665 44202 5671 44214
rect 4554 44174 5671 44202
rect 4554 44162 4560 44174
rect 5665 44162 5671 44174
rect 5723 44162 5729 44214
rect 4816 44050 4822 44102
rect 4874 44090 4880 44102
rect 5555 44090 5561 44102
rect 4874 44062 5561 44090
rect 4874 44050 4880 44062
rect 5555 44050 5561 44062
rect 5613 44050 5619 44102
rect 5376 43960 5382 44012
rect 5434 44000 5440 44012
rect 5665 44000 5671 44012
rect 5434 43972 5671 44000
rect 5434 43960 5440 43972
rect 5665 43960 5671 43972
rect 5723 43960 5729 44012
rect 5797 43925 5853 43934
rect 5797 43860 5853 43869
rect 6222 43925 6278 43934
rect 6222 43860 6278 43869
rect 6654 43925 6710 43934
rect 6654 43860 6710 43869
rect 7036 43902 7092 43911
rect 7036 43837 7092 43846
rect 7308 43902 7364 43911
rect 7308 43837 7364 43846
rect 5376 43736 5382 43788
rect 5434 43776 5440 43788
rect 5665 43776 5671 43788
rect 5434 43748 5671 43776
rect 5434 43736 5440 43748
rect 5665 43736 5671 43748
rect 5723 43736 5729 43788
rect 4816 43646 4822 43698
rect 4874 43686 4880 43698
rect 5555 43686 5561 43698
rect 4874 43658 5561 43686
rect 4874 43646 4880 43658
rect 5555 43646 5561 43658
rect 5613 43646 5619 43698
rect 4416 43534 4422 43586
rect 4474 43574 4480 43586
rect 5665 43574 5671 43586
rect 4474 43546 5671 43574
rect 4474 43534 4480 43546
rect 5665 43534 5671 43546
rect 5723 43534 5729 43586
rect 5797 43551 5853 43560
rect 7036 43507 7092 43516
rect 5797 43486 5853 43495
rect 6222 43493 6278 43502
rect 6222 43428 6278 43437
rect 6654 43493 6710 43502
rect 7036 43442 7092 43451
rect 7308 43507 7364 43516
rect 7308 43442 7364 43451
rect 6654 43428 6710 43437
rect 4336 43372 4342 43424
rect 4394 43412 4400 43424
rect 5665 43412 5671 43424
rect 4394 43384 5671 43412
rect 4394 43372 4400 43384
rect 5665 43372 5671 43384
rect 5723 43372 5729 43424
rect 4816 43260 4822 43312
rect 4874 43300 4880 43312
rect 5555 43300 5561 43312
rect 4874 43272 5561 43300
rect 4874 43260 4880 43272
rect 5555 43260 5561 43272
rect 5613 43260 5619 43312
rect 5376 43170 5382 43222
rect 5434 43210 5440 43222
rect 5665 43210 5671 43222
rect 5434 43182 5671 43210
rect 5434 43170 5440 43182
rect 5665 43170 5671 43182
rect 5723 43170 5729 43222
rect 5797 43135 5853 43144
rect 5797 43070 5853 43079
rect 6222 43135 6278 43144
rect 6222 43070 6278 43079
rect 6654 43135 6710 43144
rect 6654 43070 6710 43079
rect 7036 43112 7092 43121
rect 7036 43047 7092 43056
rect 7308 43112 7364 43121
rect 7308 43047 7364 43056
rect 5376 42946 5382 42998
rect 5434 42986 5440 42998
rect 5665 42986 5671 42998
rect 5434 42958 5671 42986
rect 5434 42946 5440 42958
rect 5665 42946 5671 42958
rect 5723 42946 5729 42998
rect 4816 42856 4822 42908
rect 4874 42896 4880 42908
rect 5555 42896 5561 42908
rect 4874 42868 5561 42896
rect 4874 42856 4880 42868
rect 5555 42856 5561 42868
rect 5613 42856 5619 42908
rect 4256 42744 4262 42796
rect 4314 42784 4320 42796
rect 5665 42784 5671 42796
rect 4314 42756 5671 42784
rect 4314 42744 4320 42756
rect 5665 42744 5671 42756
rect 5723 42744 5729 42796
rect 5797 42761 5853 42770
rect 7036 42717 7092 42726
rect 5797 42696 5853 42705
rect 6222 42703 6278 42712
rect 6222 42638 6278 42647
rect 6654 42703 6710 42712
rect 7036 42652 7092 42661
rect 7308 42717 7364 42726
rect 7308 42652 7364 42661
rect 6654 42638 6710 42647
rect 4496 42582 4502 42634
rect 4554 42622 4560 42634
rect 5665 42622 5671 42634
rect 4554 42594 5671 42622
rect 4554 42582 4560 42594
rect 5665 42582 5671 42594
rect 5723 42582 5729 42634
rect 4736 42470 4742 42522
rect 4794 42510 4800 42522
rect 5555 42510 5561 42522
rect 4794 42482 5561 42510
rect 4794 42470 4800 42482
rect 5555 42470 5561 42482
rect 5613 42470 5619 42522
rect 5376 42380 5382 42432
rect 5434 42420 5440 42432
rect 5665 42420 5671 42432
rect 5434 42392 5671 42420
rect 5434 42380 5440 42392
rect 5665 42380 5671 42392
rect 5723 42380 5729 42432
rect 5797 42345 5853 42354
rect 5797 42280 5853 42289
rect 6222 42345 6278 42354
rect 6222 42280 6278 42289
rect 6654 42345 6710 42354
rect 6654 42280 6710 42289
rect 7036 42322 7092 42331
rect 7036 42257 7092 42266
rect 7308 42322 7364 42331
rect 7308 42257 7364 42266
rect 5376 42156 5382 42208
rect 5434 42196 5440 42208
rect 5665 42196 5671 42208
rect 5434 42168 5671 42196
rect 5434 42156 5440 42168
rect 5665 42156 5671 42168
rect 5723 42156 5729 42208
rect 4736 42066 4742 42118
rect 4794 42106 4800 42118
rect 5555 42106 5561 42118
rect 4794 42078 5561 42106
rect 4794 42066 4800 42078
rect 5555 42066 5561 42078
rect 5613 42066 5619 42118
rect 4416 41954 4422 42006
rect 4474 41994 4480 42006
rect 5665 41994 5671 42006
rect 4474 41966 5671 41994
rect 4474 41954 4480 41966
rect 5665 41954 5671 41966
rect 5723 41954 5729 42006
rect 5797 41971 5853 41980
rect 7036 41927 7092 41936
rect 5797 41906 5853 41915
rect 6222 41913 6278 41922
rect 6222 41848 6278 41857
rect 6654 41913 6710 41922
rect 7036 41862 7092 41871
rect 7308 41927 7364 41936
rect 7308 41862 7364 41871
rect 6654 41848 6710 41857
rect 4336 41792 4342 41844
rect 4394 41832 4400 41844
rect 5665 41832 5671 41844
rect 4394 41804 5671 41832
rect 4394 41792 4400 41804
rect 5665 41792 5671 41804
rect 5723 41792 5729 41844
rect 4736 41680 4742 41732
rect 4794 41720 4800 41732
rect 5555 41720 5561 41732
rect 4794 41692 5561 41720
rect 4794 41680 4800 41692
rect 5555 41680 5561 41692
rect 5613 41680 5619 41732
rect 5376 41590 5382 41642
rect 5434 41630 5440 41642
rect 5665 41630 5671 41642
rect 5434 41602 5671 41630
rect 5434 41590 5440 41602
rect 5665 41590 5671 41602
rect 5723 41590 5729 41642
rect 5797 41555 5853 41564
rect 5797 41490 5853 41499
rect 6222 41555 6278 41564
rect 6222 41490 6278 41499
rect 6654 41555 6710 41564
rect 6654 41490 6710 41499
rect 7036 41532 7092 41541
rect 7036 41467 7092 41476
rect 7308 41532 7364 41541
rect 7308 41467 7364 41476
rect 5376 41366 5382 41418
rect 5434 41406 5440 41418
rect 5665 41406 5671 41418
rect 5434 41378 5671 41406
rect 5434 41366 5440 41378
rect 5665 41366 5671 41378
rect 5723 41366 5729 41418
rect 4736 41276 4742 41328
rect 4794 41316 4800 41328
rect 5555 41316 5561 41328
rect 4794 41288 5561 41316
rect 4794 41276 4800 41288
rect 5555 41276 5561 41288
rect 5613 41276 5619 41328
rect 4256 41164 4262 41216
rect 4314 41204 4320 41216
rect 5665 41204 5671 41216
rect 4314 41176 5671 41204
rect 4314 41164 4320 41176
rect 5665 41164 5671 41176
rect 5723 41164 5729 41216
rect 5797 41181 5853 41190
rect 7036 41137 7092 41146
rect 5797 41116 5853 41125
rect 6222 41123 6278 41132
rect 6222 41058 6278 41067
rect 6654 41123 6710 41132
rect 7036 41072 7092 41081
rect 7308 41137 7364 41146
rect 7308 41072 7364 41081
rect 6654 41058 6710 41067
rect 4496 41002 4502 41054
rect 4554 41042 4560 41054
rect 5665 41042 5671 41054
rect 4554 41014 5671 41042
rect 4554 41002 4560 41014
rect 5665 41002 5671 41014
rect 5723 41002 5729 41054
rect 4656 40890 4662 40942
rect 4714 40930 4720 40942
rect 5555 40930 5561 40942
rect 4714 40902 5561 40930
rect 4714 40890 4720 40902
rect 5555 40890 5561 40902
rect 5613 40890 5619 40942
rect 5376 40800 5382 40852
rect 5434 40840 5440 40852
rect 5665 40840 5671 40852
rect 5434 40812 5671 40840
rect 5434 40800 5440 40812
rect 5665 40800 5671 40812
rect 5723 40800 5729 40852
rect 5797 40765 5853 40774
rect 5797 40700 5853 40709
rect 6222 40765 6278 40774
rect 6222 40700 6278 40709
rect 6654 40765 6710 40774
rect 6654 40700 6710 40709
rect 7036 40742 7092 40751
rect 7036 40677 7092 40686
rect 7308 40742 7364 40751
rect 7308 40677 7364 40686
rect 5376 40576 5382 40628
rect 5434 40616 5440 40628
rect 5665 40616 5671 40628
rect 5434 40588 5671 40616
rect 5434 40576 5440 40588
rect 5665 40576 5671 40588
rect 5723 40576 5729 40628
rect 4656 40486 4662 40538
rect 4714 40526 4720 40538
rect 5555 40526 5561 40538
rect 4714 40498 5561 40526
rect 4714 40486 4720 40498
rect 5555 40486 5561 40498
rect 5613 40486 5619 40538
rect 4416 40374 4422 40426
rect 4474 40414 4480 40426
rect 5665 40414 5671 40426
rect 4474 40386 5671 40414
rect 4474 40374 4480 40386
rect 5665 40374 5671 40386
rect 5723 40374 5729 40426
rect 5797 40391 5853 40400
rect 7036 40347 7092 40356
rect 5797 40326 5853 40335
rect 6222 40333 6278 40342
rect 6222 40268 6278 40277
rect 6654 40333 6710 40342
rect 7036 40282 7092 40291
rect 7308 40347 7364 40356
rect 7308 40282 7364 40291
rect 6654 40268 6710 40277
rect 4336 40212 4342 40264
rect 4394 40252 4400 40264
rect 5665 40252 5671 40264
rect 4394 40224 5671 40252
rect 4394 40212 4400 40224
rect 5665 40212 5671 40224
rect 5723 40212 5729 40264
rect 4656 40100 4662 40152
rect 4714 40140 4720 40152
rect 5555 40140 5561 40152
rect 4714 40112 5561 40140
rect 4714 40100 4720 40112
rect 5555 40100 5561 40112
rect 5613 40100 5619 40152
rect 5376 40010 5382 40062
rect 5434 40050 5440 40062
rect 5665 40050 5671 40062
rect 5434 40022 5671 40050
rect 5434 40010 5440 40022
rect 5665 40010 5671 40022
rect 5723 40010 5729 40062
rect 5797 39975 5853 39984
rect 5797 39910 5853 39919
rect 6222 39975 6278 39984
rect 6222 39910 6278 39919
rect 6654 39975 6710 39984
rect 6654 39910 6710 39919
rect 7036 39952 7092 39961
rect 7036 39887 7092 39896
rect 7308 39952 7364 39961
rect 7308 39887 7364 39896
rect 5376 39786 5382 39838
rect 5434 39826 5440 39838
rect 5665 39826 5671 39838
rect 5434 39798 5671 39826
rect 5434 39786 5440 39798
rect 5665 39786 5671 39798
rect 5723 39786 5729 39838
rect 4656 39696 4662 39748
rect 4714 39736 4720 39748
rect 5555 39736 5561 39748
rect 4714 39708 5561 39736
rect 4714 39696 4720 39708
rect 5555 39696 5561 39708
rect 5613 39696 5619 39748
rect 4256 39584 4262 39636
rect 4314 39624 4320 39636
rect 5665 39624 5671 39636
rect 4314 39596 5671 39624
rect 4314 39584 4320 39596
rect 5665 39584 5671 39596
rect 5723 39584 5729 39636
rect 5797 39601 5853 39610
rect 7036 39557 7092 39566
rect 5797 39536 5853 39545
rect 6222 39543 6278 39552
rect 6222 39478 6278 39487
rect 6654 39543 6710 39552
rect 7036 39492 7092 39501
rect 7308 39557 7364 39566
rect 7308 39492 7364 39501
rect 6654 39478 6710 39487
rect 4496 39422 4502 39474
rect 4554 39462 4560 39474
rect 5665 39462 5671 39474
rect 4554 39434 5671 39462
rect 4554 39422 4560 39434
rect 5665 39422 5671 39434
rect 5723 39422 5729 39474
rect 4576 39310 4582 39362
rect 4634 39350 4640 39362
rect 5555 39350 5561 39362
rect 4634 39322 5561 39350
rect 4634 39310 4640 39322
rect 5555 39310 5561 39322
rect 5613 39310 5619 39362
rect 5376 39220 5382 39272
rect 5434 39260 5440 39272
rect 5665 39260 5671 39272
rect 5434 39232 5671 39260
rect 5434 39220 5440 39232
rect 5665 39220 5671 39232
rect 5723 39220 5729 39272
rect 5797 39185 5853 39194
rect 5797 39120 5853 39129
rect 6222 39185 6278 39194
rect 6222 39120 6278 39129
rect 6654 39185 6710 39194
rect 6654 39120 6710 39129
rect 7036 39162 7092 39171
rect 7036 39097 7092 39106
rect 7308 39162 7364 39171
rect 7308 39097 7364 39106
rect 5376 38996 5382 39048
rect 5434 39036 5440 39048
rect 5665 39036 5671 39048
rect 5434 39008 5671 39036
rect 5434 38996 5440 39008
rect 5665 38996 5671 39008
rect 5723 38996 5729 39048
rect 4576 38906 4582 38958
rect 4634 38946 4640 38958
rect 5555 38946 5561 38958
rect 4634 38918 5561 38946
rect 4634 38906 4640 38918
rect 5555 38906 5561 38918
rect 5613 38906 5619 38958
rect 4416 38794 4422 38846
rect 4474 38834 4480 38846
rect 5665 38834 5671 38846
rect 4474 38806 5671 38834
rect 4474 38794 4480 38806
rect 5665 38794 5671 38806
rect 5723 38794 5729 38846
rect 5797 38811 5853 38820
rect 7036 38767 7092 38776
rect 5797 38746 5853 38755
rect 6222 38753 6278 38762
rect 6222 38688 6278 38697
rect 6654 38753 6710 38762
rect 7036 38702 7092 38711
rect 7308 38767 7364 38776
rect 7308 38702 7364 38711
rect 6654 38688 6710 38697
rect 4336 38632 4342 38684
rect 4394 38672 4400 38684
rect 5665 38672 5671 38684
rect 4394 38644 5671 38672
rect 4394 38632 4400 38644
rect 5665 38632 5671 38644
rect 5723 38632 5729 38684
rect 4576 38520 4582 38572
rect 4634 38560 4640 38572
rect 5555 38560 5561 38572
rect 4634 38532 5561 38560
rect 4634 38520 4640 38532
rect 5555 38520 5561 38532
rect 5613 38520 5619 38572
rect 5376 38430 5382 38482
rect 5434 38470 5440 38482
rect 5665 38470 5671 38482
rect 5434 38442 5671 38470
rect 5434 38430 5440 38442
rect 5665 38430 5671 38442
rect 5723 38430 5729 38482
rect 5797 38395 5853 38404
rect 5797 38330 5853 38339
rect 6222 38395 6278 38404
rect 6222 38330 6278 38339
rect 6654 38395 6710 38404
rect 6654 38330 6710 38339
rect 7036 38372 7092 38381
rect 7036 38307 7092 38316
rect 7308 38372 7364 38381
rect 7308 38307 7364 38316
rect 5376 38206 5382 38258
rect 5434 38246 5440 38258
rect 5665 38246 5671 38258
rect 5434 38218 5671 38246
rect 5434 38206 5440 38218
rect 5665 38206 5671 38218
rect 5723 38206 5729 38258
rect 4576 38116 4582 38168
rect 4634 38156 4640 38168
rect 5555 38156 5561 38168
rect 4634 38128 5561 38156
rect 4634 38116 4640 38128
rect 5555 38116 5561 38128
rect 5613 38116 5619 38168
rect 4256 38004 4262 38056
rect 4314 38044 4320 38056
rect 5665 38044 5671 38056
rect 4314 38016 5671 38044
rect 4314 38004 4320 38016
rect 5665 38004 5671 38016
rect 5723 38004 5729 38056
rect 5797 38021 5853 38030
rect 7036 37977 7092 37986
rect 5797 37956 5853 37965
rect 6222 37963 6278 37972
rect 6222 37898 6278 37907
rect 6654 37963 6710 37972
rect 7036 37912 7092 37921
rect 7308 37977 7364 37986
rect 7308 37912 7364 37921
rect 6654 37898 6710 37907
rect 4496 37842 4502 37894
rect 4554 37882 4560 37894
rect 5665 37882 5671 37894
rect 4554 37854 5671 37882
rect 4554 37842 4560 37854
rect 5665 37842 5671 37854
rect 5723 37842 5729 37894
rect 4816 37730 4822 37782
rect 4874 37770 4880 37782
rect 5555 37770 5561 37782
rect 4874 37742 5561 37770
rect 4874 37730 4880 37742
rect 5555 37730 5561 37742
rect 5613 37730 5619 37782
rect 5296 37640 5302 37692
rect 5354 37680 5360 37692
rect 5665 37680 5671 37692
rect 5354 37652 5671 37680
rect 5354 37640 5360 37652
rect 5665 37640 5671 37652
rect 5723 37640 5729 37692
rect 5797 37605 5853 37614
rect 5797 37540 5853 37549
rect 6222 37605 6278 37614
rect 6222 37540 6278 37549
rect 6654 37605 6710 37614
rect 6654 37540 6710 37549
rect 7036 37582 7092 37591
rect 7036 37517 7092 37526
rect 7308 37582 7364 37591
rect 7308 37517 7364 37526
rect 5296 37416 5302 37468
rect 5354 37456 5360 37468
rect 5665 37456 5671 37468
rect 5354 37428 5671 37456
rect 5354 37416 5360 37428
rect 5665 37416 5671 37428
rect 5723 37416 5729 37468
rect 4816 37326 4822 37378
rect 4874 37366 4880 37378
rect 5555 37366 5561 37378
rect 4874 37338 5561 37366
rect 4874 37326 4880 37338
rect 5555 37326 5561 37338
rect 5613 37326 5619 37378
rect 4416 37214 4422 37266
rect 4474 37254 4480 37266
rect 5665 37254 5671 37266
rect 4474 37226 5671 37254
rect 4474 37214 4480 37226
rect 5665 37214 5671 37226
rect 5723 37214 5729 37266
rect 5797 37231 5853 37240
rect 7036 37187 7092 37196
rect 5797 37166 5853 37175
rect 6222 37173 6278 37182
rect 6222 37108 6278 37117
rect 6654 37173 6710 37182
rect 7036 37122 7092 37131
rect 7308 37187 7364 37196
rect 7308 37122 7364 37131
rect 6654 37108 6710 37117
rect 4336 37052 4342 37104
rect 4394 37092 4400 37104
rect 5665 37092 5671 37104
rect 4394 37064 5671 37092
rect 4394 37052 4400 37064
rect 5665 37052 5671 37064
rect 5723 37052 5729 37104
rect 4816 36940 4822 36992
rect 4874 36980 4880 36992
rect 5555 36980 5561 36992
rect 4874 36952 5561 36980
rect 4874 36940 4880 36952
rect 5555 36940 5561 36952
rect 5613 36940 5619 36992
rect 5296 36850 5302 36902
rect 5354 36890 5360 36902
rect 5665 36890 5671 36902
rect 5354 36862 5671 36890
rect 5354 36850 5360 36862
rect 5665 36850 5671 36862
rect 5723 36850 5729 36902
rect 5797 36815 5853 36824
rect 5797 36750 5853 36759
rect 6222 36815 6278 36824
rect 6222 36750 6278 36759
rect 6654 36815 6710 36824
rect 6654 36750 6710 36759
rect 7036 36792 7092 36801
rect 7036 36727 7092 36736
rect 7308 36792 7364 36801
rect 7308 36727 7364 36736
rect 5296 36626 5302 36678
rect 5354 36666 5360 36678
rect 5665 36666 5671 36678
rect 5354 36638 5671 36666
rect 5354 36626 5360 36638
rect 5665 36626 5671 36638
rect 5723 36626 5729 36678
rect 4816 36536 4822 36588
rect 4874 36576 4880 36588
rect 5555 36576 5561 36588
rect 4874 36548 5561 36576
rect 4874 36536 4880 36548
rect 5555 36536 5561 36548
rect 5613 36536 5619 36588
rect 4256 36424 4262 36476
rect 4314 36464 4320 36476
rect 5665 36464 5671 36476
rect 4314 36436 5671 36464
rect 4314 36424 4320 36436
rect 5665 36424 5671 36436
rect 5723 36424 5729 36476
rect 5797 36441 5853 36450
rect 7036 36397 7092 36406
rect 5797 36376 5853 36385
rect 6222 36383 6278 36392
rect 6222 36318 6278 36327
rect 6654 36383 6710 36392
rect 7036 36332 7092 36341
rect 7308 36397 7364 36406
rect 7308 36332 7364 36341
rect 6654 36318 6710 36327
rect 4496 36262 4502 36314
rect 4554 36302 4560 36314
rect 5665 36302 5671 36314
rect 4554 36274 5671 36302
rect 4554 36262 4560 36274
rect 5665 36262 5671 36274
rect 5723 36262 5729 36314
rect 4736 36150 4742 36202
rect 4794 36190 4800 36202
rect 5555 36190 5561 36202
rect 4794 36162 5561 36190
rect 4794 36150 4800 36162
rect 5555 36150 5561 36162
rect 5613 36150 5619 36202
rect 5296 36060 5302 36112
rect 5354 36100 5360 36112
rect 5665 36100 5671 36112
rect 5354 36072 5671 36100
rect 5354 36060 5360 36072
rect 5665 36060 5671 36072
rect 5723 36060 5729 36112
rect 5797 36025 5853 36034
rect 5797 35960 5853 35969
rect 6222 36025 6278 36034
rect 6222 35960 6278 35969
rect 6654 36025 6710 36034
rect 6654 35960 6710 35969
rect 7036 36002 7092 36011
rect 7036 35937 7092 35946
rect 7308 36002 7364 36011
rect 7308 35937 7364 35946
rect 5296 35836 5302 35888
rect 5354 35876 5360 35888
rect 5665 35876 5671 35888
rect 5354 35848 5671 35876
rect 5354 35836 5360 35848
rect 5665 35836 5671 35848
rect 5723 35836 5729 35888
rect 4736 35746 4742 35798
rect 4794 35786 4800 35798
rect 5555 35786 5561 35798
rect 4794 35758 5561 35786
rect 4794 35746 4800 35758
rect 5555 35746 5561 35758
rect 5613 35746 5619 35798
rect 4416 35634 4422 35686
rect 4474 35674 4480 35686
rect 5665 35674 5671 35686
rect 4474 35646 5671 35674
rect 4474 35634 4480 35646
rect 5665 35634 5671 35646
rect 5723 35634 5729 35686
rect 5797 35651 5853 35660
rect 7036 35607 7092 35616
rect 5797 35586 5853 35595
rect 6222 35593 6278 35602
rect 6222 35528 6278 35537
rect 6654 35593 6710 35602
rect 7036 35542 7092 35551
rect 7308 35607 7364 35616
rect 7308 35542 7364 35551
rect 6654 35528 6710 35537
rect 4336 35472 4342 35524
rect 4394 35512 4400 35524
rect 5665 35512 5671 35524
rect 4394 35484 5671 35512
rect 4394 35472 4400 35484
rect 5665 35472 5671 35484
rect 5723 35472 5729 35524
rect 4736 35360 4742 35412
rect 4794 35400 4800 35412
rect 5555 35400 5561 35412
rect 4794 35372 5561 35400
rect 4794 35360 4800 35372
rect 5555 35360 5561 35372
rect 5613 35360 5619 35412
rect 5296 35270 5302 35322
rect 5354 35310 5360 35322
rect 5665 35310 5671 35322
rect 5354 35282 5671 35310
rect 5354 35270 5360 35282
rect 5665 35270 5671 35282
rect 5723 35270 5729 35322
rect 5797 35235 5853 35244
rect 5797 35170 5853 35179
rect 6222 35235 6278 35244
rect 6222 35170 6278 35179
rect 6654 35235 6710 35244
rect 6654 35170 6710 35179
rect 7036 35212 7092 35221
rect 7036 35147 7092 35156
rect 7308 35212 7364 35221
rect 7308 35147 7364 35156
rect 5296 35046 5302 35098
rect 5354 35086 5360 35098
rect 5665 35086 5671 35098
rect 5354 35058 5671 35086
rect 5354 35046 5360 35058
rect 5665 35046 5671 35058
rect 5723 35046 5729 35098
rect 4736 34956 4742 35008
rect 4794 34996 4800 35008
rect 5555 34996 5561 35008
rect 4794 34968 5561 34996
rect 4794 34956 4800 34968
rect 5555 34956 5561 34968
rect 5613 34956 5619 35008
rect 4256 34844 4262 34896
rect 4314 34884 4320 34896
rect 5665 34884 5671 34896
rect 4314 34856 5671 34884
rect 4314 34844 4320 34856
rect 5665 34844 5671 34856
rect 5723 34844 5729 34896
rect 5797 34861 5853 34870
rect 7036 34817 7092 34826
rect 5797 34796 5853 34805
rect 6222 34803 6278 34812
rect 6222 34738 6278 34747
rect 6654 34803 6710 34812
rect 7036 34752 7092 34761
rect 7308 34817 7364 34826
rect 7308 34752 7364 34761
rect 6654 34738 6710 34747
rect 4496 34682 4502 34734
rect 4554 34722 4560 34734
rect 5665 34722 5671 34734
rect 4554 34694 5671 34722
rect 4554 34682 4560 34694
rect 5665 34682 5671 34694
rect 5723 34682 5729 34734
rect 4656 34570 4662 34622
rect 4714 34610 4720 34622
rect 5555 34610 5561 34622
rect 4714 34582 5561 34610
rect 4714 34570 4720 34582
rect 5555 34570 5561 34582
rect 5613 34570 5619 34622
rect 5296 34480 5302 34532
rect 5354 34520 5360 34532
rect 5665 34520 5671 34532
rect 5354 34492 5671 34520
rect 5354 34480 5360 34492
rect 5665 34480 5671 34492
rect 5723 34480 5729 34532
rect 5797 34445 5853 34454
rect 5797 34380 5853 34389
rect 6222 34445 6278 34454
rect 6222 34380 6278 34389
rect 6654 34445 6710 34454
rect 6654 34380 6710 34389
rect 7036 34422 7092 34431
rect 7036 34357 7092 34366
rect 7308 34422 7364 34431
rect 7308 34357 7364 34366
rect 5296 34256 5302 34308
rect 5354 34296 5360 34308
rect 5665 34296 5671 34308
rect 5354 34268 5671 34296
rect 5354 34256 5360 34268
rect 5665 34256 5671 34268
rect 5723 34256 5729 34308
rect 4656 34166 4662 34218
rect 4714 34206 4720 34218
rect 5555 34206 5561 34218
rect 4714 34178 5561 34206
rect 4714 34166 4720 34178
rect 5555 34166 5561 34178
rect 5613 34166 5619 34218
rect 4416 34054 4422 34106
rect 4474 34094 4480 34106
rect 5665 34094 5671 34106
rect 4474 34066 5671 34094
rect 4474 34054 4480 34066
rect 5665 34054 5671 34066
rect 5723 34054 5729 34106
rect 5797 34071 5853 34080
rect 7036 34027 7092 34036
rect 5797 34006 5853 34015
rect 6222 34013 6278 34022
rect 6222 33948 6278 33957
rect 6654 34013 6710 34022
rect 7036 33962 7092 33971
rect 7308 34027 7364 34036
rect 7308 33962 7364 33971
rect 6654 33948 6710 33957
rect 4336 33892 4342 33944
rect 4394 33932 4400 33944
rect 5665 33932 5671 33944
rect 4394 33904 5671 33932
rect 4394 33892 4400 33904
rect 5665 33892 5671 33904
rect 5723 33892 5729 33944
rect 4656 33780 4662 33832
rect 4714 33820 4720 33832
rect 5555 33820 5561 33832
rect 4714 33792 5561 33820
rect 4714 33780 4720 33792
rect 5555 33780 5561 33792
rect 5613 33780 5619 33832
rect 5296 33690 5302 33742
rect 5354 33730 5360 33742
rect 5665 33730 5671 33742
rect 5354 33702 5671 33730
rect 5354 33690 5360 33702
rect 5665 33690 5671 33702
rect 5723 33690 5729 33742
rect 5797 33655 5853 33664
rect 5797 33590 5853 33599
rect 6222 33655 6278 33664
rect 6222 33590 6278 33599
rect 6654 33655 6710 33664
rect 6654 33590 6710 33599
rect 7036 33632 7092 33641
rect 7036 33567 7092 33576
rect 7308 33632 7364 33641
rect 7308 33567 7364 33576
rect 5296 33466 5302 33518
rect 5354 33506 5360 33518
rect 5665 33506 5671 33518
rect 5354 33478 5671 33506
rect 5354 33466 5360 33478
rect 5665 33466 5671 33478
rect 5723 33466 5729 33518
rect 4656 33376 4662 33428
rect 4714 33416 4720 33428
rect 5555 33416 5561 33428
rect 4714 33388 5561 33416
rect 4714 33376 4720 33388
rect 5555 33376 5561 33388
rect 5613 33376 5619 33428
rect 4256 33264 4262 33316
rect 4314 33304 4320 33316
rect 5665 33304 5671 33316
rect 4314 33276 5671 33304
rect 4314 33264 4320 33276
rect 5665 33264 5671 33276
rect 5723 33264 5729 33316
rect 5797 33281 5853 33290
rect 7036 33237 7092 33246
rect 5797 33216 5853 33225
rect 6222 33223 6278 33232
rect 6222 33158 6278 33167
rect 6654 33223 6710 33232
rect 7036 33172 7092 33181
rect 7308 33237 7364 33246
rect 7308 33172 7364 33181
rect 6654 33158 6710 33167
rect 4496 33102 4502 33154
rect 4554 33142 4560 33154
rect 5665 33142 5671 33154
rect 4554 33114 5671 33142
rect 4554 33102 4560 33114
rect 5665 33102 5671 33114
rect 5723 33102 5729 33154
rect 4576 32990 4582 33042
rect 4634 33030 4640 33042
rect 5555 33030 5561 33042
rect 4634 33002 5561 33030
rect 4634 32990 4640 33002
rect 5555 32990 5561 33002
rect 5613 32990 5619 33042
rect 5296 32900 5302 32952
rect 5354 32940 5360 32952
rect 5665 32940 5671 32952
rect 5354 32912 5671 32940
rect 5354 32900 5360 32912
rect 5665 32900 5671 32912
rect 5723 32900 5729 32952
rect 5797 32865 5853 32874
rect 5797 32800 5853 32809
rect 6222 32865 6278 32874
rect 6222 32800 6278 32809
rect 6654 32865 6710 32874
rect 6654 32800 6710 32809
rect 7036 32842 7092 32851
rect 7036 32777 7092 32786
rect 7308 32842 7364 32851
rect 7308 32777 7364 32786
rect 5296 32676 5302 32728
rect 5354 32716 5360 32728
rect 5665 32716 5671 32728
rect 5354 32688 5671 32716
rect 5354 32676 5360 32688
rect 5665 32676 5671 32688
rect 5723 32676 5729 32728
rect 4576 32586 4582 32638
rect 4634 32626 4640 32638
rect 5555 32626 5561 32638
rect 4634 32598 5561 32626
rect 4634 32586 4640 32598
rect 5555 32586 5561 32598
rect 5613 32586 5619 32638
rect 4416 32474 4422 32526
rect 4474 32514 4480 32526
rect 5665 32514 5671 32526
rect 4474 32486 5671 32514
rect 4474 32474 4480 32486
rect 5665 32474 5671 32486
rect 5723 32474 5729 32526
rect 5797 32491 5853 32500
rect 7036 32447 7092 32456
rect 5797 32426 5853 32435
rect 6222 32433 6278 32442
rect 6222 32368 6278 32377
rect 6654 32433 6710 32442
rect 7036 32382 7092 32391
rect 7308 32447 7364 32456
rect 7308 32382 7364 32391
rect 6654 32368 6710 32377
rect 4336 32312 4342 32364
rect 4394 32352 4400 32364
rect 5665 32352 5671 32364
rect 4394 32324 5671 32352
rect 4394 32312 4400 32324
rect 5665 32312 5671 32324
rect 5723 32312 5729 32364
rect 4576 32200 4582 32252
rect 4634 32240 4640 32252
rect 5555 32240 5561 32252
rect 4634 32212 5561 32240
rect 4634 32200 4640 32212
rect 5555 32200 5561 32212
rect 5613 32200 5619 32252
rect 5296 32110 5302 32162
rect 5354 32150 5360 32162
rect 5665 32150 5671 32162
rect 5354 32122 5671 32150
rect 5354 32110 5360 32122
rect 5665 32110 5671 32122
rect 5723 32110 5729 32162
rect 5797 32075 5853 32084
rect 5797 32010 5853 32019
rect 6222 32075 6278 32084
rect 6222 32010 6278 32019
rect 6654 32075 6710 32084
rect 6654 32010 6710 32019
rect 7036 32052 7092 32061
rect 7036 31987 7092 31996
rect 7308 32052 7364 32061
rect 7308 31987 7364 31996
rect 5296 31886 5302 31938
rect 5354 31926 5360 31938
rect 5665 31926 5671 31938
rect 5354 31898 5671 31926
rect 5354 31886 5360 31898
rect 5665 31886 5671 31898
rect 5723 31886 5729 31938
rect 4576 31796 4582 31848
rect 4634 31836 4640 31848
rect 5555 31836 5561 31848
rect 4634 31808 5561 31836
rect 4634 31796 4640 31808
rect 5555 31796 5561 31808
rect 5613 31796 5619 31848
rect 4256 31684 4262 31736
rect 4314 31724 4320 31736
rect 5665 31724 5671 31736
rect 4314 31696 5671 31724
rect 4314 31684 4320 31696
rect 5665 31684 5671 31696
rect 5723 31684 5729 31736
rect 5797 31701 5853 31710
rect 7036 31657 7092 31666
rect 5797 31636 5853 31645
rect 6222 31643 6278 31652
rect 6222 31578 6278 31587
rect 6654 31643 6710 31652
rect 7036 31592 7092 31601
rect 7308 31657 7364 31666
rect 7308 31592 7364 31601
rect 6654 31578 6710 31587
rect 4496 31522 4502 31574
rect 4554 31562 4560 31574
rect 5665 31562 5671 31574
rect 4554 31534 5671 31562
rect 4554 31522 4560 31534
rect 5665 31522 5671 31534
rect 5723 31522 5729 31574
rect 4816 31410 4822 31462
rect 4874 31450 4880 31462
rect 5555 31450 5561 31462
rect 4874 31422 5561 31450
rect 4874 31410 4880 31422
rect 5555 31410 5561 31422
rect 5613 31410 5619 31462
rect 5216 31320 5222 31372
rect 5274 31360 5280 31372
rect 5665 31360 5671 31372
rect 5274 31332 5671 31360
rect 5274 31320 5280 31332
rect 5665 31320 5671 31332
rect 5723 31320 5729 31372
rect 5797 31285 5853 31294
rect 5797 31220 5853 31229
rect 6222 31285 6278 31294
rect 6222 31220 6278 31229
rect 6654 31285 6710 31294
rect 6654 31220 6710 31229
rect 7036 31262 7092 31271
rect 7036 31197 7092 31206
rect 7308 31262 7364 31271
rect 7308 31197 7364 31206
rect 5216 31096 5222 31148
rect 5274 31136 5280 31148
rect 5665 31136 5671 31148
rect 5274 31108 5671 31136
rect 5274 31096 5280 31108
rect 5665 31096 5671 31108
rect 5723 31096 5729 31148
rect 4816 31006 4822 31058
rect 4874 31046 4880 31058
rect 5555 31046 5561 31058
rect 4874 31018 5561 31046
rect 4874 31006 4880 31018
rect 5555 31006 5561 31018
rect 5613 31006 5619 31058
rect 4416 30894 4422 30946
rect 4474 30934 4480 30946
rect 5665 30934 5671 30946
rect 4474 30906 5671 30934
rect 4474 30894 4480 30906
rect 5665 30894 5671 30906
rect 5723 30894 5729 30946
rect 5797 30911 5853 30920
rect 7036 30867 7092 30876
rect 5797 30846 5853 30855
rect 6222 30853 6278 30862
rect 6222 30788 6278 30797
rect 6654 30853 6710 30862
rect 7036 30802 7092 30811
rect 7308 30867 7364 30876
rect 7308 30802 7364 30811
rect 6654 30788 6710 30797
rect 4336 30732 4342 30784
rect 4394 30772 4400 30784
rect 5665 30772 5671 30784
rect 4394 30744 5671 30772
rect 4394 30732 4400 30744
rect 5665 30732 5671 30744
rect 5723 30732 5729 30784
rect 4816 30620 4822 30672
rect 4874 30660 4880 30672
rect 5555 30660 5561 30672
rect 4874 30632 5561 30660
rect 4874 30620 4880 30632
rect 5555 30620 5561 30632
rect 5613 30620 5619 30672
rect 5216 30530 5222 30582
rect 5274 30570 5280 30582
rect 5665 30570 5671 30582
rect 5274 30542 5671 30570
rect 5274 30530 5280 30542
rect 5665 30530 5671 30542
rect 5723 30530 5729 30582
rect 5797 30495 5853 30504
rect 5797 30430 5853 30439
rect 6222 30495 6278 30504
rect 6222 30430 6278 30439
rect 6654 30495 6710 30504
rect 6654 30430 6710 30439
rect 7036 30472 7092 30481
rect 7036 30407 7092 30416
rect 7308 30472 7364 30481
rect 7308 30407 7364 30416
rect 5216 30306 5222 30358
rect 5274 30346 5280 30358
rect 5665 30346 5671 30358
rect 5274 30318 5671 30346
rect 5274 30306 5280 30318
rect 5665 30306 5671 30318
rect 5723 30306 5729 30358
rect 4816 30216 4822 30268
rect 4874 30256 4880 30268
rect 5555 30256 5561 30268
rect 4874 30228 5561 30256
rect 4874 30216 4880 30228
rect 5555 30216 5561 30228
rect 5613 30216 5619 30268
rect 4256 30104 4262 30156
rect 4314 30144 4320 30156
rect 5665 30144 5671 30156
rect 4314 30116 5671 30144
rect 4314 30104 4320 30116
rect 5665 30104 5671 30116
rect 5723 30104 5729 30156
rect 5797 30121 5853 30130
rect 7036 30077 7092 30086
rect 5797 30056 5853 30065
rect 6222 30063 6278 30072
rect 6222 29998 6278 30007
rect 6654 30063 6710 30072
rect 7036 30012 7092 30021
rect 7308 30077 7364 30086
rect 7308 30012 7364 30021
rect 6654 29998 6710 30007
rect 4496 29942 4502 29994
rect 4554 29982 4560 29994
rect 5665 29982 5671 29994
rect 4554 29954 5671 29982
rect 4554 29942 4560 29954
rect 5665 29942 5671 29954
rect 5723 29942 5729 29994
rect 4736 29830 4742 29882
rect 4794 29870 4800 29882
rect 5555 29870 5561 29882
rect 4794 29842 5561 29870
rect 4794 29830 4800 29842
rect 5555 29830 5561 29842
rect 5613 29830 5619 29882
rect 5216 29740 5222 29792
rect 5274 29780 5280 29792
rect 5665 29780 5671 29792
rect 5274 29752 5671 29780
rect 5274 29740 5280 29752
rect 5665 29740 5671 29752
rect 5723 29740 5729 29792
rect 5797 29705 5853 29714
rect 5797 29640 5853 29649
rect 6222 29705 6278 29714
rect 6222 29640 6278 29649
rect 6654 29705 6710 29714
rect 6654 29640 6710 29649
rect 7036 29682 7092 29691
rect 7036 29617 7092 29626
rect 7308 29682 7364 29691
rect 7308 29617 7364 29626
rect 5216 29516 5222 29568
rect 5274 29556 5280 29568
rect 5665 29556 5671 29568
rect 5274 29528 5671 29556
rect 5274 29516 5280 29528
rect 5665 29516 5671 29528
rect 5723 29516 5729 29568
rect 4736 29426 4742 29478
rect 4794 29466 4800 29478
rect 5555 29466 5561 29478
rect 4794 29438 5561 29466
rect 4794 29426 4800 29438
rect 5555 29426 5561 29438
rect 5613 29426 5619 29478
rect 4416 29314 4422 29366
rect 4474 29354 4480 29366
rect 5665 29354 5671 29366
rect 4474 29326 5671 29354
rect 4474 29314 4480 29326
rect 5665 29314 5671 29326
rect 5723 29314 5729 29366
rect 5797 29331 5853 29340
rect 7036 29287 7092 29296
rect 5797 29266 5853 29275
rect 6222 29273 6278 29282
rect 6222 29208 6278 29217
rect 6654 29273 6710 29282
rect 7036 29222 7092 29231
rect 7308 29287 7364 29296
rect 7308 29222 7364 29231
rect 6654 29208 6710 29217
rect 4336 29152 4342 29204
rect 4394 29192 4400 29204
rect 5665 29192 5671 29204
rect 4394 29164 5671 29192
rect 4394 29152 4400 29164
rect 5665 29152 5671 29164
rect 5723 29152 5729 29204
rect 4736 29040 4742 29092
rect 4794 29080 4800 29092
rect 5555 29080 5561 29092
rect 4794 29052 5561 29080
rect 4794 29040 4800 29052
rect 5555 29040 5561 29052
rect 5613 29040 5619 29092
rect 5216 28950 5222 29002
rect 5274 28990 5280 29002
rect 5665 28990 5671 29002
rect 5274 28962 5671 28990
rect 5274 28950 5280 28962
rect 5665 28950 5671 28962
rect 5723 28950 5729 29002
rect 5797 28915 5853 28924
rect 5797 28850 5853 28859
rect 6222 28915 6278 28924
rect 6222 28850 6278 28859
rect 6654 28915 6710 28924
rect 6654 28850 6710 28859
rect 7036 28892 7092 28901
rect 7036 28827 7092 28836
rect 7308 28892 7364 28901
rect 7308 28827 7364 28836
rect 5216 28726 5222 28778
rect 5274 28766 5280 28778
rect 5665 28766 5671 28778
rect 5274 28738 5671 28766
rect 5274 28726 5280 28738
rect 5665 28726 5671 28738
rect 5723 28726 5729 28778
rect 4736 28636 4742 28688
rect 4794 28676 4800 28688
rect 5555 28676 5561 28688
rect 4794 28648 5561 28676
rect 4794 28636 4800 28648
rect 5555 28636 5561 28648
rect 5613 28636 5619 28688
rect 4256 28524 4262 28576
rect 4314 28564 4320 28576
rect 5665 28564 5671 28576
rect 4314 28536 5671 28564
rect 4314 28524 4320 28536
rect 5665 28524 5671 28536
rect 5723 28524 5729 28576
rect 5797 28541 5853 28550
rect 7036 28497 7092 28506
rect 5797 28476 5853 28485
rect 6222 28483 6278 28492
rect 6222 28418 6278 28427
rect 6654 28483 6710 28492
rect 7036 28432 7092 28441
rect 7308 28497 7364 28506
rect 7308 28432 7364 28441
rect 6654 28418 6710 28427
rect 4496 28362 4502 28414
rect 4554 28402 4560 28414
rect 5665 28402 5671 28414
rect 4554 28374 5671 28402
rect 4554 28362 4560 28374
rect 5665 28362 5671 28374
rect 5723 28362 5729 28414
rect 4656 28250 4662 28302
rect 4714 28290 4720 28302
rect 5555 28290 5561 28302
rect 4714 28262 5561 28290
rect 4714 28250 4720 28262
rect 5555 28250 5561 28262
rect 5613 28250 5619 28302
rect 5216 28160 5222 28212
rect 5274 28200 5280 28212
rect 5665 28200 5671 28212
rect 5274 28172 5671 28200
rect 5274 28160 5280 28172
rect 5665 28160 5671 28172
rect 5723 28160 5729 28212
rect 5797 28125 5853 28134
rect 5797 28060 5853 28069
rect 6222 28125 6278 28134
rect 6222 28060 6278 28069
rect 6654 28125 6710 28134
rect 6654 28060 6710 28069
rect 7036 28102 7092 28111
rect 7036 28037 7092 28046
rect 7308 28102 7364 28111
rect 7308 28037 7364 28046
rect 5216 27936 5222 27988
rect 5274 27976 5280 27988
rect 5665 27976 5671 27988
rect 5274 27948 5671 27976
rect 5274 27936 5280 27948
rect 5665 27936 5671 27948
rect 5723 27936 5729 27988
rect 4656 27846 4662 27898
rect 4714 27886 4720 27898
rect 5555 27886 5561 27898
rect 4714 27858 5561 27886
rect 4714 27846 4720 27858
rect 5555 27846 5561 27858
rect 5613 27846 5619 27898
rect 4416 27734 4422 27786
rect 4474 27774 4480 27786
rect 5665 27774 5671 27786
rect 4474 27746 5671 27774
rect 4474 27734 4480 27746
rect 5665 27734 5671 27746
rect 5723 27734 5729 27786
rect 5797 27751 5853 27760
rect 7036 27707 7092 27716
rect 5797 27686 5853 27695
rect 6222 27693 6278 27702
rect 6222 27628 6278 27637
rect 6654 27693 6710 27702
rect 7036 27642 7092 27651
rect 7308 27707 7364 27716
rect 7308 27642 7364 27651
rect 6654 27628 6710 27637
rect 4336 27572 4342 27624
rect 4394 27612 4400 27624
rect 5665 27612 5671 27624
rect 4394 27584 5671 27612
rect 4394 27572 4400 27584
rect 5665 27572 5671 27584
rect 5723 27572 5729 27624
rect 4656 27460 4662 27512
rect 4714 27500 4720 27512
rect 5555 27500 5561 27512
rect 4714 27472 5561 27500
rect 4714 27460 4720 27472
rect 5555 27460 5561 27472
rect 5613 27460 5619 27512
rect 5216 27370 5222 27422
rect 5274 27410 5280 27422
rect 5665 27410 5671 27422
rect 5274 27382 5671 27410
rect 5274 27370 5280 27382
rect 5665 27370 5671 27382
rect 5723 27370 5729 27422
rect 5797 27335 5853 27344
rect 5797 27270 5853 27279
rect 6222 27335 6278 27344
rect 6222 27270 6278 27279
rect 6654 27335 6710 27344
rect 6654 27270 6710 27279
rect 7036 27312 7092 27321
rect 7036 27247 7092 27256
rect 7308 27312 7364 27321
rect 7308 27247 7364 27256
rect 5216 27146 5222 27198
rect 5274 27186 5280 27198
rect 5665 27186 5671 27198
rect 5274 27158 5671 27186
rect 5274 27146 5280 27158
rect 5665 27146 5671 27158
rect 5723 27146 5729 27198
rect 4656 27056 4662 27108
rect 4714 27096 4720 27108
rect 5555 27096 5561 27108
rect 4714 27068 5561 27096
rect 4714 27056 4720 27068
rect 5555 27056 5561 27068
rect 5613 27056 5619 27108
rect 4256 26944 4262 26996
rect 4314 26984 4320 26996
rect 5665 26984 5671 26996
rect 4314 26956 5671 26984
rect 4314 26944 4320 26956
rect 5665 26944 5671 26956
rect 5723 26944 5729 26996
rect 5797 26961 5853 26970
rect 7036 26917 7092 26926
rect 5797 26896 5853 26905
rect 6222 26903 6278 26912
rect 6222 26838 6278 26847
rect 6654 26903 6710 26912
rect 7036 26852 7092 26861
rect 7308 26917 7364 26926
rect 7308 26852 7364 26861
rect 6654 26838 6710 26847
rect 4496 26782 4502 26834
rect 4554 26822 4560 26834
rect 5665 26822 5671 26834
rect 4554 26794 5671 26822
rect 4554 26782 4560 26794
rect 5665 26782 5671 26794
rect 5723 26782 5729 26834
rect 4576 26670 4582 26722
rect 4634 26710 4640 26722
rect 5555 26710 5561 26722
rect 4634 26682 5561 26710
rect 4634 26670 4640 26682
rect 5555 26670 5561 26682
rect 5613 26670 5619 26722
rect 5216 26580 5222 26632
rect 5274 26620 5280 26632
rect 5665 26620 5671 26632
rect 5274 26592 5671 26620
rect 5274 26580 5280 26592
rect 5665 26580 5671 26592
rect 5723 26580 5729 26632
rect 5797 26545 5853 26554
rect 5797 26480 5853 26489
rect 6222 26545 6278 26554
rect 6222 26480 6278 26489
rect 6654 26545 6710 26554
rect 6654 26480 6710 26489
rect 7036 26522 7092 26531
rect 7036 26457 7092 26466
rect 7308 26522 7364 26531
rect 7308 26457 7364 26466
rect 5216 26356 5222 26408
rect 5274 26396 5280 26408
rect 5665 26396 5671 26408
rect 5274 26368 5671 26396
rect 5274 26356 5280 26368
rect 5665 26356 5671 26368
rect 5723 26356 5729 26408
rect 4576 26266 4582 26318
rect 4634 26306 4640 26318
rect 5555 26306 5561 26318
rect 4634 26278 5561 26306
rect 4634 26266 4640 26278
rect 5555 26266 5561 26278
rect 5613 26266 5619 26318
rect 4416 26154 4422 26206
rect 4474 26194 4480 26206
rect 5665 26194 5671 26206
rect 4474 26166 5671 26194
rect 4474 26154 4480 26166
rect 5665 26154 5671 26166
rect 5723 26154 5729 26206
rect 5797 26171 5853 26180
rect 7036 26127 7092 26136
rect 5797 26106 5853 26115
rect 6222 26113 6278 26122
rect 6222 26048 6278 26057
rect 6654 26113 6710 26122
rect 7036 26062 7092 26071
rect 7308 26127 7364 26136
rect 7308 26062 7364 26071
rect 6654 26048 6710 26057
rect 4336 25992 4342 26044
rect 4394 26032 4400 26044
rect 5665 26032 5671 26044
rect 4394 26004 5671 26032
rect 4394 25992 4400 26004
rect 5665 25992 5671 26004
rect 5723 25992 5729 26044
rect 4576 25880 4582 25932
rect 4634 25920 4640 25932
rect 5555 25920 5561 25932
rect 4634 25892 5561 25920
rect 4634 25880 4640 25892
rect 5555 25880 5561 25892
rect 5613 25880 5619 25932
rect 5216 25790 5222 25842
rect 5274 25830 5280 25842
rect 5665 25830 5671 25842
rect 5274 25802 5671 25830
rect 5274 25790 5280 25802
rect 5665 25790 5671 25802
rect 5723 25790 5729 25842
rect 5797 25755 5853 25764
rect 5797 25690 5853 25699
rect 6222 25755 6278 25764
rect 6222 25690 6278 25699
rect 6654 25755 6710 25764
rect 6654 25690 6710 25699
rect 7036 25732 7092 25741
rect 7036 25667 7092 25676
rect 7308 25732 7364 25741
rect 7308 25667 7364 25676
rect 5216 25566 5222 25618
rect 5274 25606 5280 25618
rect 5665 25606 5671 25618
rect 5274 25578 5671 25606
rect 5274 25566 5280 25578
rect 5665 25566 5671 25578
rect 5723 25566 5729 25618
rect 4576 25476 4582 25528
rect 4634 25516 4640 25528
rect 5555 25516 5561 25528
rect 4634 25488 5561 25516
rect 4634 25476 4640 25488
rect 5555 25476 5561 25488
rect 5613 25476 5619 25528
rect 4256 25364 4262 25416
rect 4314 25404 4320 25416
rect 5665 25404 5671 25416
rect 4314 25376 5671 25404
rect 4314 25364 4320 25376
rect 5665 25364 5671 25376
rect 5723 25364 5729 25416
rect 5797 25381 5853 25390
rect 7036 25337 7092 25346
rect 5797 25316 5853 25325
rect 6222 25323 6278 25332
rect 6222 25258 6278 25267
rect 6654 25323 6710 25332
rect 7036 25272 7092 25281
rect 7308 25337 7364 25346
rect 7308 25272 7364 25281
rect 6654 25258 6710 25267
rect 4496 25202 4502 25254
rect 4554 25242 4560 25254
rect 5665 25242 5671 25254
rect 4554 25214 5671 25242
rect 4554 25202 4560 25214
rect 5665 25202 5671 25214
rect 5723 25202 5729 25254
rect 4816 25090 4822 25142
rect 4874 25130 4880 25142
rect 5555 25130 5561 25142
rect 4874 25102 5561 25130
rect 4874 25090 4880 25102
rect 5555 25090 5561 25102
rect 5613 25090 5619 25142
rect 5136 25000 5142 25052
rect 5194 25040 5200 25052
rect 5665 25040 5671 25052
rect 5194 25012 5671 25040
rect 5194 25000 5200 25012
rect 5665 25000 5671 25012
rect 5723 25000 5729 25052
rect 5797 24965 5853 24974
rect 5797 24900 5853 24909
rect 6222 24965 6278 24974
rect 6222 24900 6278 24909
rect 6654 24965 6710 24974
rect 6654 24900 6710 24909
rect 7036 24942 7092 24951
rect 7036 24877 7092 24886
rect 7308 24942 7364 24951
rect 7308 24877 7364 24886
rect 5136 24776 5142 24828
rect 5194 24816 5200 24828
rect 5665 24816 5671 24828
rect 5194 24788 5671 24816
rect 5194 24776 5200 24788
rect 5665 24776 5671 24788
rect 5723 24776 5729 24828
rect 4816 24686 4822 24738
rect 4874 24726 4880 24738
rect 5555 24726 5561 24738
rect 4874 24698 5561 24726
rect 4874 24686 4880 24698
rect 5555 24686 5561 24698
rect 5613 24686 5619 24738
rect 4416 24574 4422 24626
rect 4474 24614 4480 24626
rect 5665 24614 5671 24626
rect 4474 24586 5671 24614
rect 4474 24574 4480 24586
rect 5665 24574 5671 24586
rect 5723 24574 5729 24626
rect 5797 24591 5853 24600
rect 7036 24547 7092 24556
rect 5797 24526 5853 24535
rect 6222 24533 6278 24542
rect 6222 24468 6278 24477
rect 6654 24533 6710 24542
rect 7036 24482 7092 24491
rect 7308 24547 7364 24556
rect 7308 24482 7364 24491
rect 6654 24468 6710 24477
rect 4336 24412 4342 24464
rect 4394 24452 4400 24464
rect 5665 24452 5671 24464
rect 4394 24424 5671 24452
rect 4394 24412 4400 24424
rect 5665 24412 5671 24424
rect 5723 24412 5729 24464
rect 4816 24300 4822 24352
rect 4874 24340 4880 24352
rect 5555 24340 5561 24352
rect 4874 24312 5561 24340
rect 4874 24300 4880 24312
rect 5555 24300 5561 24312
rect 5613 24300 5619 24352
rect 5136 24210 5142 24262
rect 5194 24250 5200 24262
rect 5665 24250 5671 24262
rect 5194 24222 5671 24250
rect 5194 24210 5200 24222
rect 5665 24210 5671 24222
rect 5723 24210 5729 24262
rect 5797 24175 5853 24184
rect 5797 24110 5853 24119
rect 6222 24175 6278 24184
rect 6222 24110 6278 24119
rect 6654 24175 6710 24184
rect 6654 24110 6710 24119
rect 7036 24152 7092 24161
rect 7036 24087 7092 24096
rect 7308 24152 7364 24161
rect 7308 24087 7364 24096
rect 5136 23986 5142 24038
rect 5194 24026 5200 24038
rect 5665 24026 5671 24038
rect 5194 23998 5671 24026
rect 5194 23986 5200 23998
rect 5665 23986 5671 23998
rect 5723 23986 5729 24038
rect 4816 23896 4822 23948
rect 4874 23936 4880 23948
rect 5555 23936 5561 23948
rect 4874 23908 5561 23936
rect 4874 23896 4880 23908
rect 5555 23896 5561 23908
rect 5613 23896 5619 23948
rect 4256 23784 4262 23836
rect 4314 23824 4320 23836
rect 5665 23824 5671 23836
rect 4314 23796 5671 23824
rect 4314 23784 4320 23796
rect 5665 23784 5671 23796
rect 5723 23784 5729 23836
rect 5797 23801 5853 23810
rect 7036 23757 7092 23766
rect 5797 23736 5853 23745
rect 6222 23743 6278 23752
rect 6222 23678 6278 23687
rect 6654 23743 6710 23752
rect 7036 23692 7092 23701
rect 7308 23757 7364 23766
rect 7308 23692 7364 23701
rect 6654 23678 6710 23687
rect 4496 23622 4502 23674
rect 4554 23662 4560 23674
rect 5665 23662 5671 23674
rect 4554 23634 5671 23662
rect 4554 23622 4560 23634
rect 5665 23622 5671 23634
rect 5723 23622 5729 23674
rect 4736 23510 4742 23562
rect 4794 23550 4800 23562
rect 5555 23550 5561 23562
rect 4794 23522 5561 23550
rect 4794 23510 4800 23522
rect 5555 23510 5561 23522
rect 5613 23510 5619 23562
rect 5136 23420 5142 23472
rect 5194 23460 5200 23472
rect 5665 23460 5671 23472
rect 5194 23432 5671 23460
rect 5194 23420 5200 23432
rect 5665 23420 5671 23432
rect 5723 23420 5729 23472
rect 5797 23385 5853 23394
rect 5797 23320 5853 23329
rect 6222 23385 6278 23394
rect 6222 23320 6278 23329
rect 6654 23385 6710 23394
rect 6654 23320 6710 23329
rect 7036 23362 7092 23371
rect 7036 23297 7092 23306
rect 7308 23362 7364 23371
rect 7308 23297 7364 23306
rect 5136 23196 5142 23248
rect 5194 23236 5200 23248
rect 5665 23236 5671 23248
rect 5194 23208 5671 23236
rect 5194 23196 5200 23208
rect 5665 23196 5671 23208
rect 5723 23196 5729 23248
rect 4736 23106 4742 23158
rect 4794 23146 4800 23158
rect 5555 23146 5561 23158
rect 4794 23118 5561 23146
rect 4794 23106 4800 23118
rect 5555 23106 5561 23118
rect 5613 23106 5619 23158
rect 4416 22994 4422 23046
rect 4474 23034 4480 23046
rect 5665 23034 5671 23046
rect 4474 23006 5671 23034
rect 4474 22994 4480 23006
rect 5665 22994 5671 23006
rect 5723 22994 5729 23046
rect 5797 23011 5853 23020
rect 7036 22967 7092 22976
rect 5797 22946 5853 22955
rect 6222 22953 6278 22962
rect 6222 22888 6278 22897
rect 6654 22953 6710 22962
rect 7036 22902 7092 22911
rect 7308 22967 7364 22976
rect 7308 22902 7364 22911
rect 6654 22888 6710 22897
rect 4336 22832 4342 22884
rect 4394 22872 4400 22884
rect 5665 22872 5671 22884
rect 4394 22844 5671 22872
rect 4394 22832 4400 22844
rect 5665 22832 5671 22844
rect 5723 22832 5729 22884
rect 4736 22720 4742 22772
rect 4794 22760 4800 22772
rect 5555 22760 5561 22772
rect 4794 22732 5561 22760
rect 4794 22720 4800 22732
rect 5555 22720 5561 22732
rect 5613 22720 5619 22772
rect 5136 22630 5142 22682
rect 5194 22670 5200 22682
rect 5665 22670 5671 22682
rect 5194 22642 5671 22670
rect 5194 22630 5200 22642
rect 5665 22630 5671 22642
rect 5723 22630 5729 22682
rect 5797 22595 5853 22604
rect 5797 22530 5853 22539
rect 6222 22595 6278 22604
rect 6222 22530 6278 22539
rect 6654 22595 6710 22604
rect 6654 22530 6710 22539
rect 7036 22572 7092 22581
rect 7036 22507 7092 22516
rect 7308 22572 7364 22581
rect 7308 22507 7364 22516
rect 5136 22406 5142 22458
rect 5194 22446 5200 22458
rect 5665 22446 5671 22458
rect 5194 22418 5671 22446
rect 5194 22406 5200 22418
rect 5665 22406 5671 22418
rect 5723 22406 5729 22458
rect 4736 22316 4742 22368
rect 4794 22356 4800 22368
rect 5555 22356 5561 22368
rect 4794 22328 5561 22356
rect 4794 22316 4800 22328
rect 5555 22316 5561 22328
rect 5613 22316 5619 22368
rect 4256 22204 4262 22256
rect 4314 22244 4320 22256
rect 5665 22244 5671 22256
rect 4314 22216 5671 22244
rect 4314 22204 4320 22216
rect 5665 22204 5671 22216
rect 5723 22204 5729 22256
rect 5797 22221 5853 22230
rect 7036 22177 7092 22186
rect 5797 22156 5853 22165
rect 6222 22163 6278 22172
rect 6222 22098 6278 22107
rect 6654 22163 6710 22172
rect 7036 22112 7092 22121
rect 7308 22177 7364 22186
rect 7308 22112 7364 22121
rect 6654 22098 6710 22107
rect 4496 22042 4502 22094
rect 4554 22082 4560 22094
rect 5665 22082 5671 22094
rect 4554 22054 5671 22082
rect 4554 22042 4560 22054
rect 5665 22042 5671 22054
rect 5723 22042 5729 22094
rect 4656 21930 4662 21982
rect 4714 21970 4720 21982
rect 5555 21970 5561 21982
rect 4714 21942 5561 21970
rect 4714 21930 4720 21942
rect 5555 21930 5561 21942
rect 5613 21930 5619 21982
rect 5136 21840 5142 21892
rect 5194 21880 5200 21892
rect 5665 21880 5671 21892
rect 5194 21852 5671 21880
rect 5194 21840 5200 21852
rect 5665 21840 5671 21852
rect 5723 21840 5729 21892
rect 5797 21805 5853 21814
rect 5797 21740 5853 21749
rect 6222 21805 6278 21814
rect 6222 21740 6278 21749
rect 6654 21805 6710 21814
rect 6654 21740 6710 21749
rect 7036 21782 7092 21791
rect 7036 21717 7092 21726
rect 7308 21782 7364 21791
rect 7308 21717 7364 21726
rect 5136 21616 5142 21668
rect 5194 21656 5200 21668
rect 5665 21656 5671 21668
rect 5194 21628 5671 21656
rect 5194 21616 5200 21628
rect 5665 21616 5671 21628
rect 5723 21616 5729 21668
rect 4656 21526 4662 21578
rect 4714 21566 4720 21578
rect 5555 21566 5561 21578
rect 4714 21538 5561 21566
rect 4714 21526 4720 21538
rect 5555 21526 5561 21538
rect 5613 21526 5619 21578
rect 4416 21414 4422 21466
rect 4474 21454 4480 21466
rect 5665 21454 5671 21466
rect 4474 21426 5671 21454
rect 4474 21414 4480 21426
rect 5665 21414 5671 21426
rect 5723 21414 5729 21466
rect 5797 21431 5853 21440
rect 7036 21387 7092 21396
rect 5797 21366 5853 21375
rect 6222 21373 6278 21382
rect 6222 21308 6278 21317
rect 6654 21373 6710 21382
rect 7036 21322 7092 21331
rect 7308 21387 7364 21396
rect 7308 21322 7364 21331
rect 6654 21308 6710 21317
rect 4336 21252 4342 21304
rect 4394 21292 4400 21304
rect 5665 21292 5671 21304
rect 4394 21264 5671 21292
rect 4394 21252 4400 21264
rect 5665 21252 5671 21264
rect 5723 21252 5729 21304
rect 4656 21140 4662 21192
rect 4714 21180 4720 21192
rect 5555 21180 5561 21192
rect 4714 21152 5561 21180
rect 4714 21140 4720 21152
rect 5555 21140 5561 21152
rect 5613 21140 5619 21192
rect 5136 21050 5142 21102
rect 5194 21090 5200 21102
rect 5665 21090 5671 21102
rect 5194 21062 5671 21090
rect 5194 21050 5200 21062
rect 5665 21050 5671 21062
rect 5723 21050 5729 21102
rect 5797 21015 5853 21024
rect 5797 20950 5853 20959
rect 6222 21015 6278 21024
rect 6222 20950 6278 20959
rect 6654 21015 6710 21024
rect 6654 20950 6710 20959
rect 7036 20992 7092 21001
rect 7036 20927 7092 20936
rect 7308 20992 7364 21001
rect 7308 20927 7364 20936
rect 5136 20826 5142 20878
rect 5194 20866 5200 20878
rect 5665 20866 5671 20878
rect 5194 20838 5671 20866
rect 5194 20826 5200 20838
rect 5665 20826 5671 20838
rect 5723 20826 5729 20878
rect 4656 20736 4662 20788
rect 4714 20776 4720 20788
rect 5555 20776 5561 20788
rect 4714 20748 5561 20776
rect 4714 20736 4720 20748
rect 5555 20736 5561 20748
rect 5613 20736 5619 20788
rect 4256 20624 4262 20676
rect 4314 20664 4320 20676
rect 5665 20664 5671 20676
rect 4314 20636 5671 20664
rect 4314 20624 4320 20636
rect 5665 20624 5671 20636
rect 5723 20624 5729 20676
rect 5797 20641 5853 20650
rect 7036 20597 7092 20606
rect 5797 20576 5853 20585
rect 6222 20583 6278 20592
rect 6222 20518 6278 20527
rect 6654 20583 6710 20592
rect 7036 20532 7092 20541
rect 7308 20597 7364 20606
rect 7308 20532 7364 20541
rect 6654 20518 6710 20527
rect 4496 20462 4502 20514
rect 4554 20502 4560 20514
rect 5665 20502 5671 20514
rect 4554 20474 5671 20502
rect 4554 20462 4560 20474
rect 5665 20462 5671 20474
rect 5723 20462 5729 20514
rect 4576 20350 4582 20402
rect 4634 20390 4640 20402
rect 5555 20390 5561 20402
rect 4634 20362 5561 20390
rect 4634 20350 4640 20362
rect 5555 20350 5561 20362
rect 5613 20350 5619 20402
rect 5136 20260 5142 20312
rect 5194 20300 5200 20312
rect 5665 20300 5671 20312
rect 5194 20272 5671 20300
rect 5194 20260 5200 20272
rect 5665 20260 5671 20272
rect 5723 20260 5729 20312
rect 5797 20225 5853 20234
rect 5797 20160 5853 20169
rect 6222 20225 6278 20234
rect 6222 20160 6278 20169
rect 6654 20225 6710 20234
rect 6654 20160 6710 20169
rect 7036 20202 7092 20211
rect 7036 20137 7092 20146
rect 7308 20202 7364 20211
rect 7308 20137 7364 20146
rect 5136 20036 5142 20088
rect 5194 20076 5200 20088
rect 5665 20076 5671 20088
rect 5194 20048 5671 20076
rect 5194 20036 5200 20048
rect 5665 20036 5671 20048
rect 5723 20036 5729 20088
rect 4576 19946 4582 19998
rect 4634 19986 4640 19998
rect 5555 19986 5561 19998
rect 4634 19958 5561 19986
rect 4634 19946 4640 19958
rect 5555 19946 5561 19958
rect 5613 19946 5619 19998
rect 4416 19834 4422 19886
rect 4474 19874 4480 19886
rect 5665 19874 5671 19886
rect 4474 19846 5671 19874
rect 4474 19834 4480 19846
rect 5665 19834 5671 19846
rect 5723 19834 5729 19886
rect 5797 19851 5853 19860
rect 7036 19807 7092 19816
rect 5797 19786 5853 19795
rect 6222 19793 6278 19802
rect 6222 19728 6278 19737
rect 6654 19793 6710 19802
rect 7036 19742 7092 19751
rect 7308 19807 7364 19816
rect 7308 19742 7364 19751
rect 6654 19728 6710 19737
rect 4336 19672 4342 19724
rect 4394 19712 4400 19724
rect 5665 19712 5671 19724
rect 4394 19684 5671 19712
rect 4394 19672 4400 19684
rect 5665 19672 5671 19684
rect 5723 19672 5729 19724
rect 4576 19560 4582 19612
rect 4634 19600 4640 19612
rect 5555 19600 5561 19612
rect 4634 19572 5561 19600
rect 4634 19560 4640 19572
rect 5555 19560 5561 19572
rect 5613 19560 5619 19612
rect 5136 19470 5142 19522
rect 5194 19510 5200 19522
rect 5665 19510 5671 19522
rect 5194 19482 5671 19510
rect 5194 19470 5200 19482
rect 5665 19470 5671 19482
rect 5723 19470 5729 19522
rect 5797 19435 5853 19444
rect 5797 19370 5853 19379
rect 6222 19435 6278 19444
rect 6222 19370 6278 19379
rect 6654 19435 6710 19444
rect 6654 19370 6710 19379
rect 7036 19412 7092 19421
rect 7036 19347 7092 19356
rect 7308 19412 7364 19421
rect 7308 19347 7364 19356
rect 5136 19246 5142 19298
rect 5194 19286 5200 19298
rect 5665 19286 5671 19298
rect 5194 19258 5671 19286
rect 5194 19246 5200 19258
rect 5665 19246 5671 19258
rect 5723 19246 5729 19298
rect 4576 19156 4582 19208
rect 4634 19196 4640 19208
rect 5555 19196 5561 19208
rect 4634 19168 5561 19196
rect 4634 19156 4640 19168
rect 5555 19156 5561 19168
rect 5613 19156 5619 19208
rect 4256 19044 4262 19096
rect 4314 19084 4320 19096
rect 5665 19084 5671 19096
rect 4314 19056 5671 19084
rect 4314 19044 4320 19056
rect 5665 19044 5671 19056
rect 5723 19044 5729 19096
rect 5797 19061 5853 19070
rect 7036 19017 7092 19026
rect 5797 18996 5853 19005
rect 6222 19003 6278 19012
rect 6222 18938 6278 18947
rect 6654 19003 6710 19012
rect 7036 18952 7092 18961
rect 7308 19017 7364 19026
rect 7308 18952 7364 18961
rect 6654 18938 6710 18947
rect 4496 18882 4502 18934
rect 4554 18922 4560 18934
rect 5665 18922 5671 18934
rect 4554 18894 5671 18922
rect 4554 18882 4560 18894
rect 5665 18882 5671 18894
rect 5723 18882 5729 18934
rect 4816 18770 4822 18822
rect 4874 18810 4880 18822
rect 5555 18810 5561 18822
rect 4874 18782 5561 18810
rect 4874 18770 4880 18782
rect 5555 18770 5561 18782
rect 5613 18770 5619 18822
rect 5056 18680 5062 18732
rect 5114 18720 5120 18732
rect 5665 18720 5671 18732
rect 5114 18692 5671 18720
rect 5114 18680 5120 18692
rect 5665 18680 5671 18692
rect 5723 18680 5729 18732
rect 5797 18645 5853 18654
rect 5797 18580 5853 18589
rect 6222 18645 6278 18654
rect 6222 18580 6278 18589
rect 6654 18645 6710 18654
rect 6654 18580 6710 18589
rect 7036 18622 7092 18631
rect 7036 18557 7092 18566
rect 7308 18622 7364 18631
rect 7308 18557 7364 18566
rect 5056 18456 5062 18508
rect 5114 18496 5120 18508
rect 5665 18496 5671 18508
rect 5114 18468 5671 18496
rect 5114 18456 5120 18468
rect 5665 18456 5671 18468
rect 5723 18456 5729 18508
rect 4816 18366 4822 18418
rect 4874 18406 4880 18418
rect 5555 18406 5561 18418
rect 4874 18378 5561 18406
rect 4874 18366 4880 18378
rect 5555 18366 5561 18378
rect 5613 18366 5619 18418
rect 4416 18254 4422 18306
rect 4474 18294 4480 18306
rect 5665 18294 5671 18306
rect 4474 18266 5671 18294
rect 4474 18254 4480 18266
rect 5665 18254 5671 18266
rect 5723 18254 5729 18306
rect 5797 18271 5853 18280
rect 7036 18227 7092 18236
rect 5797 18206 5853 18215
rect 6222 18213 6278 18222
rect 6222 18148 6278 18157
rect 6654 18213 6710 18222
rect 7036 18162 7092 18171
rect 7308 18227 7364 18236
rect 7308 18162 7364 18171
rect 6654 18148 6710 18157
rect 4336 18092 4342 18144
rect 4394 18132 4400 18144
rect 5665 18132 5671 18144
rect 4394 18104 5671 18132
rect 4394 18092 4400 18104
rect 5665 18092 5671 18104
rect 5723 18092 5729 18144
rect 4816 17980 4822 18032
rect 4874 18020 4880 18032
rect 5555 18020 5561 18032
rect 4874 17992 5561 18020
rect 4874 17980 4880 17992
rect 5555 17980 5561 17992
rect 5613 17980 5619 18032
rect 5056 17890 5062 17942
rect 5114 17930 5120 17942
rect 5665 17930 5671 17942
rect 5114 17902 5671 17930
rect 5114 17890 5120 17902
rect 5665 17890 5671 17902
rect 5723 17890 5729 17942
rect 5797 17855 5853 17864
rect 5797 17790 5853 17799
rect 6222 17855 6278 17864
rect 6222 17790 6278 17799
rect 6654 17855 6710 17864
rect 6654 17790 6710 17799
rect 7036 17832 7092 17841
rect 7036 17767 7092 17776
rect 7308 17832 7364 17841
rect 7308 17767 7364 17776
rect 5056 17666 5062 17718
rect 5114 17706 5120 17718
rect 5665 17706 5671 17718
rect 5114 17678 5671 17706
rect 5114 17666 5120 17678
rect 5665 17666 5671 17678
rect 5723 17666 5729 17718
rect 4816 17576 4822 17628
rect 4874 17616 4880 17628
rect 5555 17616 5561 17628
rect 4874 17588 5561 17616
rect 4874 17576 4880 17588
rect 5555 17576 5561 17588
rect 5613 17576 5619 17628
rect 4256 17464 4262 17516
rect 4314 17504 4320 17516
rect 5665 17504 5671 17516
rect 4314 17476 5671 17504
rect 4314 17464 4320 17476
rect 5665 17464 5671 17476
rect 5723 17464 5729 17516
rect 5797 17481 5853 17490
rect 7036 17437 7092 17446
rect 5797 17416 5853 17425
rect 6222 17423 6278 17432
rect 6222 17358 6278 17367
rect 6654 17423 6710 17432
rect 7036 17372 7092 17381
rect 7308 17437 7364 17446
rect 7308 17372 7364 17381
rect 6654 17358 6710 17367
rect 4496 17302 4502 17354
rect 4554 17342 4560 17354
rect 5665 17342 5671 17354
rect 4554 17314 5671 17342
rect 4554 17302 4560 17314
rect 5665 17302 5671 17314
rect 5723 17302 5729 17354
rect 4736 17190 4742 17242
rect 4794 17230 4800 17242
rect 5555 17230 5561 17242
rect 4794 17202 5561 17230
rect 4794 17190 4800 17202
rect 5555 17190 5561 17202
rect 5613 17190 5619 17242
rect 5056 17100 5062 17152
rect 5114 17140 5120 17152
rect 5665 17140 5671 17152
rect 5114 17112 5671 17140
rect 5114 17100 5120 17112
rect 5665 17100 5671 17112
rect 5723 17100 5729 17152
rect 5797 17065 5853 17074
rect 5797 17000 5853 17009
rect 6222 17065 6278 17074
rect 6222 17000 6278 17009
rect 6654 17065 6710 17074
rect 6654 17000 6710 17009
rect 7036 17042 7092 17051
rect 7036 16977 7092 16986
rect 7308 17042 7364 17051
rect 7308 16977 7364 16986
rect 5056 16876 5062 16928
rect 5114 16916 5120 16928
rect 5665 16916 5671 16928
rect 5114 16888 5671 16916
rect 5114 16876 5120 16888
rect 5665 16876 5671 16888
rect 5723 16876 5729 16928
rect 4736 16786 4742 16838
rect 4794 16826 4800 16838
rect 5555 16826 5561 16838
rect 4794 16798 5561 16826
rect 4794 16786 4800 16798
rect 5555 16786 5561 16798
rect 5613 16786 5619 16838
rect 4416 16674 4422 16726
rect 4474 16714 4480 16726
rect 5665 16714 5671 16726
rect 4474 16686 5671 16714
rect 4474 16674 4480 16686
rect 5665 16674 5671 16686
rect 5723 16674 5729 16726
rect 5797 16691 5853 16700
rect 7036 16647 7092 16656
rect 5797 16626 5853 16635
rect 6222 16633 6278 16642
rect 6222 16568 6278 16577
rect 6654 16633 6710 16642
rect 7036 16582 7092 16591
rect 7308 16647 7364 16656
rect 7308 16582 7364 16591
rect 6654 16568 6710 16577
rect 4336 16512 4342 16564
rect 4394 16552 4400 16564
rect 5665 16552 5671 16564
rect 4394 16524 5671 16552
rect 4394 16512 4400 16524
rect 5665 16512 5671 16524
rect 5723 16512 5729 16564
rect 4736 16400 4742 16452
rect 4794 16440 4800 16452
rect 5555 16440 5561 16452
rect 4794 16412 5561 16440
rect 4794 16400 4800 16412
rect 5555 16400 5561 16412
rect 5613 16400 5619 16452
rect 5056 16310 5062 16362
rect 5114 16350 5120 16362
rect 5665 16350 5671 16362
rect 5114 16322 5671 16350
rect 5114 16310 5120 16322
rect 5665 16310 5671 16322
rect 5723 16310 5729 16362
rect 5797 16275 5853 16284
rect 5797 16210 5853 16219
rect 6222 16275 6278 16284
rect 6222 16210 6278 16219
rect 6654 16275 6710 16284
rect 6654 16210 6710 16219
rect 7036 16252 7092 16261
rect 7036 16187 7092 16196
rect 7308 16252 7364 16261
rect 7308 16187 7364 16196
rect 5056 16086 5062 16138
rect 5114 16126 5120 16138
rect 5665 16126 5671 16138
rect 5114 16098 5671 16126
rect 5114 16086 5120 16098
rect 5665 16086 5671 16098
rect 5723 16086 5729 16138
rect 4736 15996 4742 16048
rect 4794 16036 4800 16048
rect 5555 16036 5561 16048
rect 4794 16008 5561 16036
rect 4794 15996 4800 16008
rect 5555 15996 5561 16008
rect 5613 15996 5619 16048
rect 4256 15884 4262 15936
rect 4314 15924 4320 15936
rect 5665 15924 5671 15936
rect 4314 15896 5671 15924
rect 4314 15884 4320 15896
rect 5665 15884 5671 15896
rect 5723 15884 5729 15936
rect 5797 15901 5853 15910
rect 7036 15857 7092 15866
rect 5797 15836 5853 15845
rect 6222 15843 6278 15852
rect 6222 15778 6278 15787
rect 6654 15843 6710 15852
rect 7036 15792 7092 15801
rect 7308 15857 7364 15866
rect 7308 15792 7364 15801
rect 6654 15778 6710 15787
rect 4496 15722 4502 15774
rect 4554 15762 4560 15774
rect 5665 15762 5671 15774
rect 4554 15734 5671 15762
rect 4554 15722 4560 15734
rect 5665 15722 5671 15734
rect 5723 15722 5729 15774
rect 4656 15610 4662 15662
rect 4714 15650 4720 15662
rect 5555 15650 5561 15662
rect 4714 15622 5561 15650
rect 4714 15610 4720 15622
rect 5555 15610 5561 15622
rect 5613 15610 5619 15662
rect 5056 15520 5062 15572
rect 5114 15560 5120 15572
rect 5665 15560 5671 15572
rect 5114 15532 5671 15560
rect 5114 15520 5120 15532
rect 5665 15520 5671 15532
rect 5723 15520 5729 15572
rect 5797 15485 5853 15494
rect 5797 15420 5853 15429
rect 6222 15485 6278 15494
rect 6222 15420 6278 15429
rect 6654 15485 6710 15494
rect 6654 15420 6710 15429
rect 7036 15462 7092 15471
rect 7036 15397 7092 15406
rect 7308 15462 7364 15471
rect 7308 15397 7364 15406
rect 5056 15296 5062 15348
rect 5114 15336 5120 15348
rect 5665 15336 5671 15348
rect 5114 15308 5671 15336
rect 5114 15296 5120 15308
rect 5665 15296 5671 15308
rect 5723 15296 5729 15348
rect 4656 15206 4662 15258
rect 4714 15246 4720 15258
rect 5555 15246 5561 15258
rect 4714 15218 5561 15246
rect 4714 15206 4720 15218
rect 5555 15206 5561 15218
rect 5613 15206 5619 15258
rect 4416 15094 4422 15146
rect 4474 15134 4480 15146
rect 5665 15134 5671 15146
rect 4474 15106 5671 15134
rect 4474 15094 4480 15106
rect 5665 15094 5671 15106
rect 5723 15094 5729 15146
rect 5797 15111 5853 15120
rect 7036 15067 7092 15076
rect 5797 15046 5853 15055
rect 6222 15053 6278 15062
rect 6222 14988 6278 14997
rect 6654 15053 6710 15062
rect 7036 15002 7092 15011
rect 7308 15067 7364 15076
rect 7308 15002 7364 15011
rect 6654 14988 6710 14997
rect 4336 14932 4342 14984
rect 4394 14972 4400 14984
rect 5665 14972 5671 14984
rect 4394 14944 5671 14972
rect 4394 14932 4400 14944
rect 5665 14932 5671 14944
rect 5723 14932 5729 14984
rect 4656 14820 4662 14872
rect 4714 14860 4720 14872
rect 5555 14860 5561 14872
rect 4714 14832 5561 14860
rect 4714 14820 4720 14832
rect 5555 14820 5561 14832
rect 5613 14820 5619 14872
rect 5056 14730 5062 14782
rect 5114 14770 5120 14782
rect 5665 14770 5671 14782
rect 5114 14742 5671 14770
rect 5114 14730 5120 14742
rect 5665 14730 5671 14742
rect 5723 14730 5729 14782
rect 5797 14695 5853 14704
rect 5797 14630 5853 14639
rect 6222 14695 6278 14704
rect 6222 14630 6278 14639
rect 6654 14695 6710 14704
rect 6654 14630 6710 14639
rect 7036 14672 7092 14681
rect 7036 14607 7092 14616
rect 7308 14672 7364 14681
rect 7308 14607 7364 14616
rect 5056 14506 5062 14558
rect 5114 14546 5120 14558
rect 5665 14546 5671 14558
rect 5114 14518 5671 14546
rect 5114 14506 5120 14518
rect 5665 14506 5671 14518
rect 5723 14506 5729 14558
rect 4656 14416 4662 14468
rect 4714 14456 4720 14468
rect 5555 14456 5561 14468
rect 4714 14428 5561 14456
rect 4714 14416 4720 14428
rect 5555 14416 5561 14428
rect 5613 14416 5619 14468
rect 4256 14304 4262 14356
rect 4314 14344 4320 14356
rect 5665 14344 5671 14356
rect 4314 14316 5671 14344
rect 4314 14304 4320 14316
rect 5665 14304 5671 14316
rect 5723 14304 5729 14356
rect 5797 14321 5853 14330
rect 7036 14277 7092 14286
rect 5797 14256 5853 14265
rect 6222 14263 6278 14272
rect 6222 14198 6278 14207
rect 6654 14263 6710 14272
rect 7036 14212 7092 14221
rect 7308 14277 7364 14286
rect 7308 14212 7364 14221
rect 6654 14198 6710 14207
rect 4496 14142 4502 14194
rect 4554 14182 4560 14194
rect 5665 14182 5671 14194
rect 4554 14154 5671 14182
rect 4554 14142 4560 14154
rect 5665 14142 5671 14154
rect 5723 14142 5729 14194
rect 4576 14030 4582 14082
rect 4634 14070 4640 14082
rect 5555 14070 5561 14082
rect 4634 14042 5561 14070
rect 4634 14030 4640 14042
rect 5555 14030 5561 14042
rect 5613 14030 5619 14082
rect 5056 13940 5062 13992
rect 5114 13980 5120 13992
rect 5665 13980 5671 13992
rect 5114 13952 5671 13980
rect 5114 13940 5120 13952
rect 5665 13940 5671 13952
rect 5723 13940 5729 13992
rect 5797 13905 5853 13914
rect 5797 13840 5853 13849
rect 6222 13905 6278 13914
rect 6222 13840 6278 13849
rect 6654 13905 6710 13914
rect 6654 13840 6710 13849
rect 7036 13882 7092 13891
rect 7036 13817 7092 13826
rect 7308 13882 7364 13891
rect 7308 13817 7364 13826
rect 5056 13716 5062 13768
rect 5114 13756 5120 13768
rect 5665 13756 5671 13768
rect 5114 13728 5671 13756
rect 5114 13716 5120 13728
rect 5665 13716 5671 13728
rect 5723 13716 5729 13768
rect 4576 13626 4582 13678
rect 4634 13666 4640 13678
rect 5555 13666 5561 13678
rect 4634 13638 5561 13666
rect 4634 13626 4640 13638
rect 5555 13626 5561 13638
rect 5613 13626 5619 13678
rect 4416 13514 4422 13566
rect 4474 13554 4480 13566
rect 5665 13554 5671 13566
rect 4474 13526 5671 13554
rect 4474 13514 4480 13526
rect 5665 13514 5671 13526
rect 5723 13514 5729 13566
rect 5797 13531 5853 13540
rect 7036 13487 7092 13496
rect 5797 13466 5853 13475
rect 6222 13473 6278 13482
rect 6222 13408 6278 13417
rect 6654 13473 6710 13482
rect 7036 13422 7092 13431
rect 7308 13487 7364 13496
rect 7308 13422 7364 13431
rect 6654 13408 6710 13417
rect 4336 13352 4342 13404
rect 4394 13392 4400 13404
rect 5665 13392 5671 13404
rect 4394 13364 5671 13392
rect 4394 13352 4400 13364
rect 5665 13352 5671 13364
rect 5723 13352 5729 13404
rect 4576 13240 4582 13292
rect 4634 13280 4640 13292
rect 5555 13280 5561 13292
rect 4634 13252 5561 13280
rect 4634 13240 4640 13252
rect 5555 13240 5561 13252
rect 5613 13240 5619 13292
rect 5056 13150 5062 13202
rect 5114 13190 5120 13202
rect 5665 13190 5671 13202
rect 5114 13162 5671 13190
rect 5114 13150 5120 13162
rect 5665 13150 5671 13162
rect 5723 13150 5729 13202
rect 5797 13115 5853 13124
rect 5797 13050 5853 13059
rect 6222 13115 6278 13124
rect 6222 13050 6278 13059
rect 6654 13115 6710 13124
rect 6654 13050 6710 13059
rect 7036 13092 7092 13101
rect 7036 13027 7092 13036
rect 7308 13092 7364 13101
rect 7308 13027 7364 13036
rect 5056 12926 5062 12978
rect 5114 12966 5120 12978
rect 5665 12966 5671 12978
rect 5114 12938 5671 12966
rect 5114 12926 5120 12938
rect 5665 12926 5671 12938
rect 5723 12926 5729 12978
rect 4576 12836 4582 12888
rect 4634 12876 4640 12888
rect 5555 12876 5561 12888
rect 4634 12848 5561 12876
rect 4634 12836 4640 12848
rect 5555 12836 5561 12848
rect 5613 12836 5619 12888
rect 4256 12724 4262 12776
rect 4314 12764 4320 12776
rect 5665 12764 5671 12776
rect 4314 12736 5671 12764
rect 4314 12724 4320 12736
rect 5665 12724 5671 12736
rect 5723 12724 5729 12776
rect 5797 12741 5853 12750
rect 7036 12697 7092 12706
rect 5797 12676 5853 12685
rect 6222 12683 6278 12692
rect 6222 12618 6278 12627
rect 6654 12683 6710 12692
rect 7036 12632 7092 12641
rect 7308 12697 7364 12706
rect 7308 12632 7364 12641
rect 6654 12618 6710 12627
rect 4496 12562 4502 12614
rect 4554 12602 4560 12614
rect 5665 12602 5671 12614
rect 4554 12574 5671 12602
rect 4554 12562 4560 12574
rect 5665 12562 5671 12574
rect 5723 12562 5729 12614
rect 4816 12450 4822 12502
rect 4874 12490 4880 12502
rect 5555 12490 5561 12502
rect 4874 12462 5561 12490
rect 4874 12450 4880 12462
rect 5555 12450 5561 12462
rect 5613 12450 5619 12502
rect 4976 12360 4982 12412
rect 5034 12400 5040 12412
rect 5665 12400 5671 12412
rect 5034 12372 5671 12400
rect 5034 12360 5040 12372
rect 5665 12360 5671 12372
rect 5723 12360 5729 12412
rect 5797 12325 5853 12334
rect 5797 12260 5853 12269
rect 6222 12325 6278 12334
rect 6222 12260 6278 12269
rect 6654 12325 6710 12334
rect 6654 12260 6710 12269
rect 7036 12302 7092 12311
rect 7036 12237 7092 12246
rect 7308 12302 7364 12311
rect 7308 12237 7364 12246
rect 4976 12136 4982 12188
rect 5034 12176 5040 12188
rect 5665 12176 5671 12188
rect 5034 12148 5671 12176
rect 5034 12136 5040 12148
rect 5665 12136 5671 12148
rect 5723 12136 5729 12188
rect 4816 12046 4822 12098
rect 4874 12086 4880 12098
rect 5555 12086 5561 12098
rect 4874 12058 5561 12086
rect 4874 12046 4880 12058
rect 5555 12046 5561 12058
rect 5613 12046 5619 12098
rect 4416 11934 4422 11986
rect 4474 11974 4480 11986
rect 5665 11974 5671 11986
rect 4474 11946 5671 11974
rect 4474 11934 4480 11946
rect 5665 11934 5671 11946
rect 5723 11934 5729 11986
rect 5797 11951 5853 11960
rect 7036 11907 7092 11916
rect 5797 11886 5853 11895
rect 6222 11893 6278 11902
rect 6222 11828 6278 11837
rect 6654 11893 6710 11902
rect 7036 11842 7092 11851
rect 7308 11907 7364 11916
rect 7308 11842 7364 11851
rect 6654 11828 6710 11837
rect 4336 11772 4342 11824
rect 4394 11812 4400 11824
rect 5665 11812 5671 11824
rect 4394 11784 5671 11812
rect 4394 11772 4400 11784
rect 5665 11772 5671 11784
rect 5723 11772 5729 11824
rect 4816 11660 4822 11712
rect 4874 11700 4880 11712
rect 5555 11700 5561 11712
rect 4874 11672 5561 11700
rect 4874 11660 4880 11672
rect 5555 11660 5561 11672
rect 5613 11660 5619 11712
rect 4976 11570 4982 11622
rect 5034 11610 5040 11622
rect 5665 11610 5671 11622
rect 5034 11582 5671 11610
rect 5034 11570 5040 11582
rect 5665 11570 5671 11582
rect 5723 11570 5729 11622
rect 5797 11535 5853 11544
rect 5797 11470 5853 11479
rect 6222 11535 6278 11544
rect 6222 11470 6278 11479
rect 6654 11535 6710 11544
rect 6654 11470 6710 11479
rect 7036 11512 7092 11521
rect 7036 11447 7092 11456
rect 7308 11512 7364 11521
rect 7308 11447 7364 11456
rect 4976 11346 4982 11398
rect 5034 11386 5040 11398
rect 5665 11386 5671 11398
rect 5034 11358 5671 11386
rect 5034 11346 5040 11358
rect 5665 11346 5671 11358
rect 5723 11346 5729 11398
rect 4816 11256 4822 11308
rect 4874 11296 4880 11308
rect 5555 11296 5561 11308
rect 4874 11268 5561 11296
rect 4874 11256 4880 11268
rect 5555 11256 5561 11268
rect 5613 11256 5619 11308
rect 4256 11144 4262 11196
rect 4314 11184 4320 11196
rect 5665 11184 5671 11196
rect 4314 11156 5671 11184
rect 4314 11144 4320 11156
rect 5665 11144 5671 11156
rect 5723 11144 5729 11196
rect 5797 11161 5853 11170
rect 7036 11117 7092 11126
rect 5797 11096 5853 11105
rect 6222 11103 6278 11112
rect 6222 11038 6278 11047
rect 6654 11103 6710 11112
rect 7036 11052 7092 11061
rect 7308 11117 7364 11126
rect 7308 11052 7364 11061
rect 6654 11038 6710 11047
rect 4496 10982 4502 11034
rect 4554 11022 4560 11034
rect 5665 11022 5671 11034
rect 4554 10994 5671 11022
rect 4554 10982 4560 10994
rect 5665 10982 5671 10994
rect 5723 10982 5729 11034
rect 4736 10870 4742 10922
rect 4794 10910 4800 10922
rect 5555 10910 5561 10922
rect 4794 10882 5561 10910
rect 4794 10870 4800 10882
rect 5555 10870 5561 10882
rect 5613 10870 5619 10922
rect 4976 10780 4982 10832
rect 5034 10820 5040 10832
rect 5665 10820 5671 10832
rect 5034 10792 5671 10820
rect 5034 10780 5040 10792
rect 5665 10780 5671 10792
rect 5723 10780 5729 10832
rect 5797 10745 5853 10754
rect 5797 10680 5853 10689
rect 6222 10745 6278 10754
rect 6222 10680 6278 10689
rect 6654 10745 6710 10754
rect 6654 10680 6710 10689
rect 7036 10722 7092 10731
rect 7036 10657 7092 10666
rect 7308 10722 7364 10731
rect 7308 10657 7364 10666
rect 4976 10556 4982 10608
rect 5034 10596 5040 10608
rect 5665 10596 5671 10608
rect 5034 10568 5671 10596
rect 5034 10556 5040 10568
rect 5665 10556 5671 10568
rect 5723 10556 5729 10608
rect 4736 10466 4742 10518
rect 4794 10506 4800 10518
rect 5555 10506 5561 10518
rect 4794 10478 5561 10506
rect 4794 10466 4800 10478
rect 5555 10466 5561 10478
rect 5613 10466 5619 10518
rect 4416 10354 4422 10406
rect 4474 10394 4480 10406
rect 5665 10394 5671 10406
rect 4474 10366 5671 10394
rect 4474 10354 4480 10366
rect 5665 10354 5671 10366
rect 5723 10354 5729 10406
rect 5797 10371 5853 10380
rect 7036 10327 7092 10336
rect 5797 10306 5853 10315
rect 6222 10313 6278 10322
rect 6222 10248 6278 10257
rect 6654 10313 6710 10322
rect 7036 10262 7092 10271
rect 7308 10327 7364 10336
rect 7308 10262 7364 10271
rect 6654 10248 6710 10257
rect 4336 10192 4342 10244
rect 4394 10232 4400 10244
rect 5665 10232 5671 10244
rect 4394 10204 5671 10232
rect 4394 10192 4400 10204
rect 5665 10192 5671 10204
rect 5723 10192 5729 10244
rect 4736 10080 4742 10132
rect 4794 10120 4800 10132
rect 5555 10120 5561 10132
rect 4794 10092 5561 10120
rect 4794 10080 4800 10092
rect 5555 10080 5561 10092
rect 5613 10080 5619 10132
rect 4976 9990 4982 10042
rect 5034 10030 5040 10042
rect 5665 10030 5671 10042
rect 5034 10002 5671 10030
rect 5034 9990 5040 10002
rect 5665 9990 5671 10002
rect 5723 9990 5729 10042
rect 5797 9955 5853 9964
rect 5797 9890 5853 9899
rect 6222 9955 6278 9964
rect 6222 9890 6278 9899
rect 6654 9955 6710 9964
rect 6654 9890 6710 9899
rect 7036 9932 7092 9941
rect 7036 9867 7092 9876
rect 7308 9932 7364 9941
rect 7308 9867 7364 9876
rect 4976 9766 4982 9818
rect 5034 9806 5040 9818
rect 5665 9806 5671 9818
rect 5034 9778 5671 9806
rect 5034 9766 5040 9778
rect 5665 9766 5671 9778
rect 5723 9766 5729 9818
rect 4736 9676 4742 9728
rect 4794 9716 4800 9728
rect 5555 9716 5561 9728
rect 4794 9688 5561 9716
rect 4794 9676 4800 9688
rect 5555 9676 5561 9688
rect 5613 9676 5619 9728
rect 4256 9564 4262 9616
rect 4314 9604 4320 9616
rect 5665 9604 5671 9616
rect 4314 9576 5671 9604
rect 4314 9564 4320 9576
rect 5665 9564 5671 9576
rect 5723 9564 5729 9616
rect 5797 9581 5853 9590
rect 7036 9537 7092 9546
rect 5797 9516 5853 9525
rect 6222 9523 6278 9532
rect 6222 9458 6278 9467
rect 6654 9523 6710 9532
rect 7036 9472 7092 9481
rect 7308 9537 7364 9546
rect 7308 9472 7364 9481
rect 6654 9458 6710 9467
rect 4496 9402 4502 9454
rect 4554 9442 4560 9454
rect 5665 9442 5671 9454
rect 4554 9414 5671 9442
rect 4554 9402 4560 9414
rect 5665 9402 5671 9414
rect 5723 9402 5729 9454
rect 4656 9290 4662 9342
rect 4714 9330 4720 9342
rect 5555 9330 5561 9342
rect 4714 9302 5561 9330
rect 4714 9290 4720 9302
rect 5555 9290 5561 9302
rect 5613 9290 5619 9342
rect 4976 9200 4982 9252
rect 5034 9240 5040 9252
rect 5665 9240 5671 9252
rect 5034 9212 5671 9240
rect 5034 9200 5040 9212
rect 5665 9200 5671 9212
rect 5723 9200 5729 9252
rect 5797 9165 5853 9174
rect 5797 9100 5853 9109
rect 6222 9165 6278 9174
rect 6222 9100 6278 9109
rect 6654 9165 6710 9174
rect 6654 9100 6710 9109
rect 7036 9142 7092 9151
rect 7036 9077 7092 9086
rect 7308 9142 7364 9151
rect 7308 9077 7364 9086
rect 4976 8976 4982 9028
rect 5034 9016 5040 9028
rect 5665 9016 5671 9028
rect 5034 8988 5671 9016
rect 5034 8976 5040 8988
rect 5665 8976 5671 8988
rect 5723 8976 5729 9028
rect 4656 8886 4662 8938
rect 4714 8926 4720 8938
rect 5555 8926 5561 8938
rect 4714 8898 5561 8926
rect 4714 8886 4720 8898
rect 5555 8886 5561 8898
rect 5613 8886 5619 8938
rect 4416 8774 4422 8826
rect 4474 8814 4480 8826
rect 5665 8814 5671 8826
rect 4474 8786 5671 8814
rect 4474 8774 4480 8786
rect 5665 8774 5671 8786
rect 5723 8774 5729 8826
rect 5797 8791 5853 8800
rect 7036 8747 7092 8756
rect 5797 8726 5853 8735
rect 6222 8733 6278 8742
rect 6222 8668 6278 8677
rect 6654 8733 6710 8742
rect 7036 8682 7092 8691
rect 7308 8747 7364 8756
rect 7308 8682 7364 8691
rect 6654 8668 6710 8677
rect 4336 8612 4342 8664
rect 4394 8652 4400 8664
rect 5665 8652 5671 8664
rect 4394 8624 5671 8652
rect 4394 8612 4400 8624
rect 5665 8612 5671 8624
rect 5723 8612 5729 8664
rect 4656 8500 4662 8552
rect 4714 8540 4720 8552
rect 5555 8540 5561 8552
rect 4714 8512 5561 8540
rect 4714 8500 4720 8512
rect 5555 8500 5561 8512
rect 5613 8500 5619 8552
rect 4976 8410 4982 8462
rect 5034 8450 5040 8462
rect 5665 8450 5671 8462
rect 5034 8422 5671 8450
rect 5034 8410 5040 8422
rect 5665 8410 5671 8422
rect 5723 8410 5729 8462
rect 5797 8375 5853 8384
rect 5797 8310 5853 8319
rect 6222 8375 6278 8384
rect 6222 8310 6278 8319
rect 6654 8375 6710 8384
rect 6654 8310 6710 8319
rect 7036 8352 7092 8361
rect 7036 8287 7092 8296
rect 7308 8352 7364 8361
rect 7308 8287 7364 8296
rect 4976 8186 4982 8238
rect 5034 8226 5040 8238
rect 5665 8226 5671 8238
rect 5034 8198 5671 8226
rect 5034 8186 5040 8198
rect 5665 8186 5671 8198
rect 5723 8186 5729 8238
rect 4656 8096 4662 8148
rect 4714 8136 4720 8148
rect 5555 8136 5561 8148
rect 4714 8108 5561 8136
rect 4714 8096 4720 8108
rect 5555 8096 5561 8108
rect 5613 8096 5619 8148
rect 4256 7984 4262 8036
rect 4314 8024 4320 8036
rect 5665 8024 5671 8036
rect 4314 7996 5671 8024
rect 4314 7984 4320 7996
rect 5665 7984 5671 7996
rect 5723 7984 5729 8036
rect 5797 8001 5853 8010
rect 7036 7957 7092 7966
rect 5797 7936 5853 7945
rect 6222 7943 6278 7952
rect 6222 7878 6278 7887
rect 6654 7943 6710 7952
rect 7036 7892 7092 7901
rect 7308 7957 7364 7966
rect 7308 7892 7364 7901
rect 6654 7878 6710 7887
rect 4496 7822 4502 7874
rect 4554 7862 4560 7874
rect 5665 7862 5671 7874
rect 4554 7834 5671 7862
rect 4554 7822 4560 7834
rect 5665 7822 5671 7834
rect 5723 7822 5729 7874
rect 4576 7710 4582 7762
rect 4634 7750 4640 7762
rect 5555 7750 5561 7762
rect 4634 7722 5561 7750
rect 4634 7710 4640 7722
rect 5555 7710 5561 7722
rect 5613 7710 5619 7762
rect 4976 7620 4982 7672
rect 5034 7660 5040 7672
rect 5665 7660 5671 7672
rect 5034 7632 5671 7660
rect 5034 7620 5040 7632
rect 5665 7620 5671 7632
rect 5723 7620 5729 7672
rect 5797 7585 5853 7594
rect 5797 7520 5853 7529
rect 6222 7585 6278 7594
rect 6222 7520 6278 7529
rect 6654 7585 6710 7594
rect 6654 7520 6710 7529
rect 7036 7562 7092 7571
rect 7036 7497 7092 7506
rect 7308 7562 7364 7571
rect 7308 7497 7364 7506
rect 4976 7396 4982 7448
rect 5034 7436 5040 7448
rect 5665 7436 5671 7448
rect 5034 7408 5671 7436
rect 5034 7396 5040 7408
rect 5665 7396 5671 7408
rect 5723 7396 5729 7448
rect 4576 7306 4582 7358
rect 4634 7346 4640 7358
rect 5555 7346 5561 7358
rect 4634 7318 5561 7346
rect 4634 7306 4640 7318
rect 5555 7306 5561 7318
rect 5613 7306 5619 7358
rect 4416 7194 4422 7246
rect 4474 7234 4480 7246
rect 5665 7234 5671 7246
rect 4474 7206 5671 7234
rect 4474 7194 4480 7206
rect 5665 7194 5671 7206
rect 5723 7194 5729 7246
rect 5797 7211 5853 7220
rect 7036 7167 7092 7176
rect 5797 7146 5853 7155
rect 6222 7153 6278 7162
rect 6222 7088 6278 7097
rect 6654 7153 6710 7162
rect 7036 7102 7092 7111
rect 7308 7167 7364 7176
rect 7308 7102 7364 7111
rect 6654 7088 6710 7097
rect 4336 7032 4342 7084
rect 4394 7072 4400 7084
rect 5665 7072 5671 7084
rect 4394 7044 5671 7072
rect 4394 7032 4400 7044
rect 5665 7032 5671 7044
rect 5723 7032 5729 7084
rect 4576 6920 4582 6972
rect 4634 6960 4640 6972
rect 5555 6960 5561 6972
rect 4634 6932 5561 6960
rect 4634 6920 4640 6932
rect 5555 6920 5561 6932
rect 5613 6920 5619 6972
rect 4976 6830 4982 6882
rect 5034 6870 5040 6882
rect 5665 6870 5671 6882
rect 5034 6842 5671 6870
rect 5034 6830 5040 6842
rect 5665 6830 5671 6842
rect 5723 6830 5729 6882
rect 5797 6795 5853 6804
rect 5797 6730 5853 6739
rect 6222 6795 6278 6804
rect 6222 6730 6278 6739
rect 6654 6795 6710 6804
rect 6654 6730 6710 6739
rect 7036 6772 7092 6781
rect 7036 6707 7092 6716
rect 7308 6772 7364 6781
rect 7308 6707 7364 6716
rect 4976 6606 4982 6658
rect 5034 6646 5040 6658
rect 5665 6646 5671 6658
rect 5034 6618 5671 6646
rect 5034 6606 5040 6618
rect 5665 6606 5671 6618
rect 5723 6606 5729 6658
rect 4576 6516 4582 6568
rect 4634 6556 4640 6568
rect 5555 6556 5561 6568
rect 4634 6528 5561 6556
rect 4634 6516 4640 6528
rect 5555 6516 5561 6528
rect 5613 6516 5619 6568
rect 4256 6404 4262 6456
rect 4314 6444 4320 6456
rect 5665 6444 5671 6456
rect 4314 6416 5671 6444
rect 4314 6404 4320 6416
rect 5665 6404 5671 6416
rect 5723 6404 5729 6456
rect 5797 6421 5853 6430
rect 7036 6377 7092 6386
rect 5797 6356 5853 6365
rect 6222 6363 6278 6372
rect 6222 6298 6278 6307
rect 6654 6363 6710 6372
rect 7036 6312 7092 6321
rect 7308 6377 7364 6386
rect 7308 6312 7364 6321
rect 6654 6298 6710 6307
rect 4496 6242 4502 6294
rect 4554 6282 4560 6294
rect 5665 6282 5671 6294
rect 4554 6254 5671 6282
rect 4554 6242 4560 6254
rect 5665 6242 5671 6254
rect 5723 6242 5729 6294
rect 4816 6130 4822 6182
rect 4874 6170 4880 6182
rect 5555 6170 5561 6182
rect 4874 6142 5561 6170
rect 4874 6130 4880 6142
rect 5555 6130 5561 6142
rect 5613 6130 5619 6182
rect 4896 6040 4902 6092
rect 4954 6080 4960 6092
rect 5665 6080 5671 6092
rect 4954 6052 5671 6080
rect 4954 6040 4960 6052
rect 5665 6040 5671 6052
rect 5723 6040 5729 6092
rect 5797 6005 5853 6014
rect 5797 5940 5853 5949
rect 6222 6005 6278 6014
rect 6222 5940 6278 5949
rect 6654 6005 6710 6014
rect 6654 5940 6710 5949
rect 7036 5982 7092 5991
rect 7036 5917 7092 5926
rect 7308 5982 7364 5991
rect 7308 5917 7364 5926
rect 4896 5816 4902 5868
rect 4954 5856 4960 5868
rect 5665 5856 5671 5868
rect 4954 5828 5671 5856
rect 4954 5816 4960 5828
rect 5665 5816 5671 5828
rect 5723 5816 5729 5868
rect 834 5782 886 5788
rect 480 5730 486 5782
rect 538 5770 544 5782
rect 538 5742 834 5770
rect 538 5730 544 5742
rect 834 5724 886 5730
rect 4816 5726 4822 5778
rect 4874 5766 4880 5778
rect 5555 5766 5561 5778
rect 4874 5738 5561 5766
rect 4874 5726 4880 5738
rect 5555 5726 5561 5738
rect 5613 5726 5619 5778
rect 4416 5614 4422 5666
rect 4474 5654 4480 5666
rect 5665 5654 5671 5666
rect 4474 5626 5671 5654
rect 4474 5614 4480 5626
rect 5665 5614 5671 5626
rect 5723 5614 5729 5666
rect 5797 5631 5853 5640
rect 7036 5587 7092 5596
rect 5797 5566 5853 5575
rect 6222 5573 6278 5582
rect 6222 5508 6278 5517
rect 6654 5573 6710 5582
rect 7036 5522 7092 5531
rect 7308 5587 7364 5596
rect 7308 5522 7364 5531
rect 6654 5508 6710 5517
rect 4336 5452 4342 5504
rect 4394 5492 4400 5504
rect 5665 5492 5671 5504
rect 4394 5464 5671 5492
rect 4394 5452 4400 5464
rect 5665 5452 5671 5464
rect 5723 5452 5729 5504
rect 754 5388 806 5394
rect 400 5336 406 5388
rect 458 5376 464 5388
rect 458 5348 754 5376
rect 458 5336 464 5348
rect 4816 5340 4822 5392
rect 4874 5380 4880 5392
rect 5555 5380 5561 5392
rect 4874 5352 5561 5380
rect 4874 5340 4880 5352
rect 5555 5340 5561 5352
rect 5613 5340 5619 5392
rect 754 5330 806 5336
rect 4896 5250 4902 5302
rect 4954 5290 4960 5302
rect 5665 5290 5671 5302
rect 4954 5262 5671 5290
rect 4954 5250 4960 5262
rect 5665 5250 5671 5262
rect 5723 5250 5729 5302
rect 5797 5215 5853 5224
rect 5797 5150 5853 5159
rect 6222 5215 6278 5224
rect 6222 5150 6278 5159
rect 6654 5215 6710 5224
rect 6654 5150 6710 5159
rect 7036 5192 7092 5201
rect 7036 5127 7092 5136
rect 7308 5192 7364 5201
rect 7308 5127 7364 5136
rect 4896 5026 4902 5078
rect 4954 5066 4960 5078
rect 5665 5066 5671 5078
rect 4954 5038 5671 5066
rect 4954 5026 4960 5038
rect 5665 5026 5671 5038
rect 5723 5026 5729 5078
rect 674 4992 726 4998
rect 320 4940 326 4992
rect 378 4980 384 4992
rect 378 4952 674 4980
rect 378 4940 384 4952
rect 674 4934 726 4940
rect 4816 4936 4822 4988
rect 4874 4976 4880 4988
rect 5555 4976 5561 4988
rect 4874 4948 5561 4976
rect 4874 4936 4880 4948
rect 5555 4936 5561 4948
rect 5613 4936 5619 4988
rect 4256 4824 4262 4876
rect 4314 4864 4320 4876
rect 5665 4864 5671 4876
rect 4314 4836 5671 4864
rect 4314 4824 4320 4836
rect 5665 4824 5671 4836
rect 5723 4824 5729 4876
rect 5797 4841 5853 4850
rect 7036 4797 7092 4806
rect 5797 4776 5853 4785
rect 6222 4783 6278 4792
rect 6222 4718 6278 4727
rect 6654 4783 6710 4792
rect 7036 4732 7092 4741
rect 7308 4797 7364 4806
rect 7308 4732 7364 4741
rect 6654 4718 6710 4727
rect 4496 4662 4502 4714
rect 4554 4702 4560 4714
rect 5665 4702 5671 4714
rect 4554 4674 5671 4702
rect 4554 4662 4560 4674
rect 5665 4662 5671 4674
rect 5723 4662 5729 4714
rect 4736 4550 4742 4602
rect 4794 4590 4800 4602
rect 5555 4590 5561 4602
rect 4794 4562 5561 4590
rect 4794 4550 4800 4562
rect 5555 4550 5561 4562
rect 5613 4550 5619 4602
rect 4896 4460 4902 4512
rect 4954 4500 4960 4512
rect 5665 4500 5671 4512
rect 4954 4472 5671 4500
rect 4954 4460 4960 4472
rect 5665 4460 5671 4472
rect 5723 4460 5729 4512
rect 5797 4425 5853 4434
rect 5797 4360 5853 4369
rect 6222 4425 6278 4434
rect 6222 4360 6278 4369
rect 6654 4425 6710 4434
rect 6654 4360 6710 4369
rect 7036 4402 7092 4411
rect 7036 4337 7092 4346
rect 7308 4402 7364 4411
rect 7308 4337 7364 4346
rect 4896 4236 4902 4288
rect 4954 4276 4960 4288
rect 5665 4276 5671 4288
rect 4954 4248 5671 4276
rect 4954 4236 4960 4248
rect 5665 4236 5671 4248
rect 5723 4236 5729 4288
rect 4736 4146 4742 4198
rect 4794 4186 4800 4198
rect 5555 4186 5561 4198
rect 4794 4158 5561 4186
rect 4794 4146 4800 4158
rect 5555 4146 5561 4158
rect 5613 4146 5619 4198
rect 4416 4034 4422 4086
rect 4474 4074 4480 4086
rect 5665 4074 5671 4086
rect 4474 4046 5671 4074
rect 4474 4034 4480 4046
rect 5665 4034 5671 4046
rect 5723 4034 5729 4086
rect 5797 4051 5853 4060
rect 7036 4007 7092 4016
rect 5797 3986 5853 3995
rect 6222 3993 6278 4002
rect 6222 3928 6278 3937
rect 6654 3993 6710 4002
rect 7036 3942 7092 3951
rect 7308 4007 7364 4016
rect 7308 3942 7364 3951
rect 6654 3928 6710 3937
rect 4336 3872 4342 3924
rect 4394 3912 4400 3924
rect 5665 3912 5671 3924
rect 4394 3884 5671 3912
rect 4394 3872 4400 3884
rect 5665 3872 5671 3884
rect 5723 3872 5729 3924
rect 4736 3760 4742 3812
rect 4794 3800 4800 3812
rect 5555 3800 5561 3812
rect 4794 3772 5561 3800
rect 4794 3760 4800 3772
rect 5555 3760 5561 3772
rect 5613 3760 5619 3812
rect 4896 3670 4902 3722
rect 4954 3710 4960 3722
rect 5665 3710 5671 3722
rect 4954 3682 5671 3710
rect 4954 3670 4960 3682
rect 5665 3670 5671 3682
rect 5723 3670 5729 3722
rect 5797 3635 5853 3644
rect 5797 3570 5853 3579
rect 6222 3635 6278 3644
rect 6222 3570 6278 3579
rect 6654 3635 6710 3644
rect 6654 3570 6710 3579
rect 7036 3612 7092 3621
rect 7036 3547 7092 3556
rect 7308 3612 7364 3621
rect 7308 3547 7364 3556
rect 4896 3446 4902 3498
rect 4954 3486 4960 3498
rect 5665 3486 5671 3498
rect 4954 3458 5671 3486
rect 4954 3446 4960 3458
rect 5665 3446 5671 3458
rect 5723 3446 5729 3498
rect 4736 3356 4742 3408
rect 4794 3396 4800 3408
rect 5555 3396 5561 3408
rect 4794 3368 5561 3396
rect 4794 3356 4800 3368
rect 5555 3356 5561 3368
rect 5613 3356 5619 3408
rect 4256 3244 4262 3296
rect 4314 3284 4320 3296
rect 5665 3284 5671 3296
rect 4314 3256 5671 3284
rect 4314 3244 4320 3256
rect 5665 3244 5671 3256
rect 5723 3244 5729 3296
rect 5797 3261 5853 3270
rect 7036 3217 7092 3226
rect 5797 3196 5853 3205
rect 6222 3203 6278 3212
rect 6222 3138 6278 3147
rect 6654 3203 6710 3212
rect 7036 3152 7092 3161
rect 7308 3217 7364 3226
rect 7308 3152 7364 3161
rect 6654 3138 6710 3147
rect 4496 3082 4502 3134
rect 4554 3122 4560 3134
rect 5665 3122 5671 3134
rect 4554 3094 5671 3122
rect 4554 3082 4560 3094
rect 5665 3082 5671 3094
rect 5723 3082 5729 3134
rect 1430 3018 1482 3024
rect 240 2966 246 3018
rect 298 3006 304 3018
rect 298 2978 1430 3006
rect 298 2966 304 2978
rect 4656 2970 4662 3022
rect 4714 3010 4720 3022
rect 5555 3010 5561 3022
rect 4714 2982 5561 3010
rect 4714 2970 4720 2982
rect 5555 2970 5561 2982
rect 5613 2970 5619 3022
rect 1430 2960 1482 2966
rect 4896 2880 4902 2932
rect 4954 2920 4960 2932
rect 5665 2920 5671 2932
rect 4954 2892 5671 2920
rect 4954 2880 4960 2892
rect 5665 2880 5671 2892
rect 5723 2880 5729 2932
rect 5797 2845 5853 2854
rect 5797 2780 5853 2789
rect 6222 2845 6278 2854
rect 6222 2780 6278 2789
rect 6654 2845 6710 2854
rect 6654 2780 6710 2789
rect 7036 2822 7092 2831
rect 7036 2757 7092 2766
rect 7308 2822 7364 2831
rect 7308 2757 7364 2766
rect 4896 2656 4902 2708
rect 4954 2696 4960 2708
rect 5665 2696 5671 2708
rect 4954 2668 5671 2696
rect 4954 2656 4960 2668
rect 5665 2656 5671 2668
rect 5723 2656 5729 2708
rect 1350 2622 1402 2628
rect 160 2570 166 2622
rect 218 2610 224 2622
rect 218 2582 1350 2610
rect 218 2570 224 2582
rect 1350 2564 1402 2570
rect 4656 2566 4662 2618
rect 4714 2606 4720 2618
rect 5555 2606 5561 2618
rect 4714 2578 5561 2606
rect 4714 2566 4720 2578
rect 5555 2566 5561 2578
rect 5613 2566 5619 2618
rect 4416 2454 4422 2506
rect 4474 2494 4480 2506
rect 5665 2494 5671 2506
rect 4474 2466 5671 2494
rect 4474 2454 4480 2466
rect 5665 2454 5671 2466
rect 5723 2454 5729 2506
rect 5797 2471 5853 2480
rect 7036 2427 7092 2436
rect 5797 2406 5853 2415
rect 6222 2413 6278 2422
rect 6222 2348 6278 2357
rect 6654 2413 6710 2422
rect 7036 2362 7092 2371
rect 7308 2427 7364 2436
rect 7308 2362 7364 2371
rect 6654 2348 6710 2357
rect 4336 2292 4342 2344
rect 4394 2332 4400 2344
rect 5665 2332 5671 2344
rect 4394 2304 5671 2332
rect 4394 2292 4400 2304
rect 5665 2292 5671 2304
rect 5723 2292 5729 2344
rect 4656 2180 4662 2232
rect 4714 2220 4720 2232
rect 5555 2220 5561 2232
rect 4714 2192 5561 2220
rect 4714 2180 4720 2192
rect 5555 2180 5561 2192
rect 5613 2180 5619 2232
rect 4896 2090 4902 2142
rect 4954 2130 4960 2142
rect 5665 2130 5671 2142
rect 4954 2102 5671 2130
rect 4954 2090 4960 2102
rect 5665 2090 5671 2102
rect 5723 2090 5729 2142
rect 5797 2055 5853 2064
rect 5797 1990 5853 1999
rect 6222 2055 6278 2064
rect 6222 1990 6278 1999
rect 6654 2055 6710 2064
rect 6654 1990 6710 1999
rect 7036 2032 7092 2041
rect 7036 1967 7092 1976
rect 7308 2032 7364 2041
rect 7308 1967 7364 1976
rect 4896 1866 4902 1918
rect 4954 1906 4960 1918
rect 5665 1906 5671 1918
rect 4954 1878 5671 1906
rect 4954 1866 4960 1878
rect 5665 1866 5671 1878
rect 5723 1866 5729 1918
rect 4656 1776 4662 1828
rect 4714 1816 4720 1828
rect 5555 1816 5561 1828
rect 4714 1788 5561 1816
rect 4714 1776 4720 1788
rect 5555 1776 5561 1788
rect 5613 1776 5619 1828
rect 4256 1664 4262 1716
rect 4314 1704 4320 1716
rect 5665 1704 5671 1716
rect 4314 1676 5671 1704
rect 4314 1664 4320 1676
rect 5665 1664 5671 1676
rect 5723 1664 5729 1716
rect 5797 1681 5853 1690
rect 7036 1637 7092 1646
rect 5797 1616 5853 1625
rect 6222 1623 6278 1632
rect 6222 1558 6278 1567
rect 6654 1623 6710 1632
rect 7036 1572 7092 1581
rect 7308 1637 7364 1646
rect 7308 1572 7364 1581
rect 6654 1558 6710 1567
rect 4496 1502 4502 1554
rect 4554 1542 4560 1554
rect 5665 1542 5671 1554
rect 4554 1514 5671 1542
rect 4554 1502 4560 1514
rect 5665 1502 5671 1514
rect 5723 1502 5729 1554
rect 4576 1390 4582 1442
rect 4634 1430 4640 1442
rect 5555 1430 5561 1442
rect 4634 1402 5561 1430
rect 4634 1390 4640 1402
rect 5555 1390 5561 1402
rect 5613 1390 5619 1442
rect 4896 1300 4902 1352
rect 4954 1340 4960 1352
rect 5665 1340 5671 1352
rect 4954 1312 5671 1340
rect 4954 1300 4960 1312
rect 5665 1300 5671 1312
rect 5723 1300 5729 1352
rect 5797 1265 5853 1274
rect 5797 1200 5853 1209
rect 6222 1265 6278 1274
rect 6222 1200 6278 1209
rect 6654 1265 6710 1274
rect 6654 1200 6710 1209
rect 7036 1242 7092 1251
rect 7036 1177 7092 1186
rect 7308 1242 7364 1251
rect 7308 1177 7364 1186
rect 4896 1076 4902 1128
rect 4954 1116 4960 1128
rect 5665 1116 5671 1128
rect 4954 1088 5671 1116
rect 4954 1076 4960 1088
rect 5665 1076 5671 1088
rect 5723 1076 5729 1128
rect 4576 986 4582 1038
rect 4634 1026 4640 1038
rect 5555 1026 5561 1038
rect 4634 998 5561 1026
rect 4634 986 4640 998
rect 5555 986 5561 998
rect 5613 986 5619 1038
rect 4416 874 4422 926
rect 4474 914 4480 926
rect 5665 914 5671 926
rect 4474 886 5671 914
rect 4474 874 4480 886
rect 5665 874 5671 886
rect 5723 874 5729 926
rect 5797 891 5853 900
rect 7036 847 7092 856
rect 5797 826 5853 835
rect 6222 833 6278 842
rect 6222 768 6278 777
rect 6654 833 6710 842
rect 7036 782 7092 791
rect 7308 847 7364 856
rect 7308 782 7364 791
rect 6654 768 6710 777
rect 4336 712 4342 764
rect 4394 752 4400 764
rect 5665 752 5671 764
rect 4394 724 5671 752
rect 4394 712 4400 724
rect 5665 712 5671 724
rect 5723 712 5729 764
rect 1430 648 1482 654
rect 80 596 86 648
rect 138 636 144 648
rect 138 608 1430 636
rect 138 596 144 608
rect 4576 600 4582 652
rect 4634 640 4640 652
rect 5555 640 5561 652
rect 4634 612 5561 640
rect 4634 600 4640 612
rect 5555 600 5561 612
rect 5613 600 5619 652
rect 1430 590 1482 596
rect 4896 510 4902 562
rect 4954 550 4960 562
rect 5665 550 5671 562
rect 4954 522 5671 550
rect 4954 510 4960 522
rect 5665 510 5671 522
rect 5723 510 5729 562
rect 5797 475 5853 484
rect 5797 410 5853 419
rect 6222 475 6278 484
rect 6222 410 6278 419
rect 6654 475 6710 484
rect 6654 410 6710 419
rect 7036 452 7092 461
rect 7036 387 7092 396
rect 7308 452 7364 461
rect 7308 387 7364 396
rect 4896 286 4902 338
rect 4954 326 4960 338
rect 5665 326 5671 338
rect 4954 298 5671 326
rect 4954 286 4960 298
rect 5665 286 5671 298
rect 5723 286 5729 338
rect 1350 252 1402 258
rect 0 200 6 252
rect 58 240 64 252
rect 58 212 1350 240
rect 58 200 64 212
rect 1350 194 1402 200
rect 4576 196 4582 248
rect 4634 236 4640 248
rect 5555 236 5561 248
rect 4634 208 5561 236
rect 4634 196 4640 208
rect 5555 196 5561 208
rect 5613 196 5619 248
rect 4256 84 4262 136
rect 4314 124 4320 136
rect 5665 124 5671 136
rect 4314 96 5671 124
rect 4314 84 4320 96
rect 5665 84 5671 96
rect 5723 84 5729 136
<< via2 >>
rect 5797 50243 5853 50245
rect 5797 50191 5799 50243
rect 5799 50191 5851 50243
rect 5851 50191 5853 50243
rect 5797 50189 5853 50191
rect 6222 50243 6278 50245
rect 6222 50191 6224 50243
rect 6224 50191 6276 50243
rect 6276 50191 6278 50243
rect 6222 50189 6278 50191
rect 6654 50243 6710 50245
rect 6654 50191 6656 50243
rect 6656 50191 6708 50243
rect 6708 50191 6710 50243
rect 6654 50189 6710 50191
rect 7036 50220 7092 50222
rect 7036 50168 7038 50220
rect 7038 50168 7090 50220
rect 7090 50168 7092 50220
rect 7036 50166 7092 50168
rect 7308 50220 7364 50222
rect 7308 50168 7310 50220
rect 7310 50168 7362 50220
rect 7362 50168 7364 50220
rect 7308 50166 7364 50168
rect 5797 49869 5853 49871
rect 5797 49817 5799 49869
rect 5799 49817 5851 49869
rect 5851 49817 5853 49869
rect 7036 49825 7092 49827
rect 5797 49815 5853 49817
rect 6222 49811 6278 49813
rect 6222 49759 6224 49811
rect 6224 49759 6276 49811
rect 6276 49759 6278 49811
rect 6222 49757 6278 49759
rect 6654 49811 6710 49813
rect 6654 49759 6656 49811
rect 6656 49759 6708 49811
rect 6708 49759 6710 49811
rect 7036 49773 7038 49825
rect 7038 49773 7090 49825
rect 7090 49773 7092 49825
rect 7036 49771 7092 49773
rect 7308 49825 7364 49827
rect 7308 49773 7310 49825
rect 7310 49773 7362 49825
rect 7362 49773 7364 49825
rect 7308 49771 7364 49773
rect 6654 49757 6710 49759
rect 5797 49453 5853 49455
rect 5797 49401 5799 49453
rect 5799 49401 5851 49453
rect 5851 49401 5853 49453
rect 5797 49399 5853 49401
rect 6222 49453 6278 49455
rect 6222 49401 6224 49453
rect 6224 49401 6276 49453
rect 6276 49401 6278 49453
rect 6222 49399 6278 49401
rect 6654 49453 6710 49455
rect 6654 49401 6656 49453
rect 6656 49401 6708 49453
rect 6708 49401 6710 49453
rect 6654 49399 6710 49401
rect 7036 49430 7092 49432
rect 7036 49378 7038 49430
rect 7038 49378 7090 49430
rect 7090 49378 7092 49430
rect 7036 49376 7092 49378
rect 7308 49430 7364 49432
rect 7308 49378 7310 49430
rect 7310 49378 7362 49430
rect 7362 49378 7364 49430
rect 7308 49376 7364 49378
rect 5797 49079 5853 49081
rect 5797 49027 5799 49079
rect 5799 49027 5851 49079
rect 5851 49027 5853 49079
rect 7036 49035 7092 49037
rect 5797 49025 5853 49027
rect 6222 49021 6278 49023
rect 6222 48969 6224 49021
rect 6224 48969 6276 49021
rect 6276 48969 6278 49021
rect 6222 48967 6278 48969
rect 6654 49021 6710 49023
rect 6654 48969 6656 49021
rect 6656 48969 6708 49021
rect 6708 48969 6710 49021
rect 7036 48983 7038 49035
rect 7038 48983 7090 49035
rect 7090 48983 7092 49035
rect 7036 48981 7092 48983
rect 7308 49035 7364 49037
rect 7308 48983 7310 49035
rect 7310 48983 7362 49035
rect 7362 48983 7364 49035
rect 7308 48981 7364 48983
rect 6654 48967 6710 48969
rect 5797 48663 5853 48665
rect 5797 48611 5799 48663
rect 5799 48611 5851 48663
rect 5851 48611 5853 48663
rect 5797 48609 5853 48611
rect 6222 48663 6278 48665
rect 6222 48611 6224 48663
rect 6224 48611 6276 48663
rect 6276 48611 6278 48663
rect 6222 48609 6278 48611
rect 6654 48663 6710 48665
rect 6654 48611 6656 48663
rect 6656 48611 6708 48663
rect 6708 48611 6710 48663
rect 6654 48609 6710 48611
rect 7036 48640 7092 48642
rect 7036 48588 7038 48640
rect 7038 48588 7090 48640
rect 7090 48588 7092 48640
rect 7036 48586 7092 48588
rect 7308 48640 7364 48642
rect 7308 48588 7310 48640
rect 7310 48588 7362 48640
rect 7362 48588 7364 48640
rect 7308 48586 7364 48588
rect 5797 48289 5853 48291
rect 5797 48237 5799 48289
rect 5799 48237 5851 48289
rect 5851 48237 5853 48289
rect 7036 48245 7092 48247
rect 5797 48235 5853 48237
rect 6222 48231 6278 48233
rect 6222 48179 6224 48231
rect 6224 48179 6276 48231
rect 6276 48179 6278 48231
rect 6222 48177 6278 48179
rect 6654 48231 6710 48233
rect 6654 48179 6656 48231
rect 6656 48179 6708 48231
rect 6708 48179 6710 48231
rect 7036 48193 7038 48245
rect 7038 48193 7090 48245
rect 7090 48193 7092 48245
rect 7036 48191 7092 48193
rect 7308 48245 7364 48247
rect 7308 48193 7310 48245
rect 7310 48193 7362 48245
rect 7362 48193 7364 48245
rect 7308 48191 7364 48193
rect 6654 48177 6710 48179
rect 5797 47873 5853 47875
rect 5797 47821 5799 47873
rect 5799 47821 5851 47873
rect 5851 47821 5853 47873
rect 5797 47819 5853 47821
rect 6222 47873 6278 47875
rect 6222 47821 6224 47873
rect 6224 47821 6276 47873
rect 6276 47821 6278 47873
rect 6222 47819 6278 47821
rect 6654 47873 6710 47875
rect 6654 47821 6656 47873
rect 6656 47821 6708 47873
rect 6708 47821 6710 47873
rect 6654 47819 6710 47821
rect 7036 47850 7092 47852
rect 7036 47798 7038 47850
rect 7038 47798 7090 47850
rect 7090 47798 7092 47850
rect 7036 47796 7092 47798
rect 7308 47850 7364 47852
rect 7308 47798 7310 47850
rect 7310 47798 7362 47850
rect 7362 47798 7364 47850
rect 7308 47796 7364 47798
rect 5797 47499 5853 47501
rect 5797 47447 5799 47499
rect 5799 47447 5851 47499
rect 5851 47447 5853 47499
rect 7036 47455 7092 47457
rect 5797 47445 5853 47447
rect 6222 47441 6278 47443
rect 6222 47389 6224 47441
rect 6224 47389 6276 47441
rect 6276 47389 6278 47441
rect 6222 47387 6278 47389
rect 6654 47441 6710 47443
rect 6654 47389 6656 47441
rect 6656 47389 6708 47441
rect 6708 47389 6710 47441
rect 7036 47403 7038 47455
rect 7038 47403 7090 47455
rect 7090 47403 7092 47455
rect 7036 47401 7092 47403
rect 7308 47455 7364 47457
rect 7308 47403 7310 47455
rect 7310 47403 7362 47455
rect 7362 47403 7364 47455
rect 7308 47401 7364 47403
rect 6654 47387 6710 47389
rect 5797 47083 5853 47085
rect 5797 47031 5799 47083
rect 5799 47031 5851 47083
rect 5851 47031 5853 47083
rect 5797 47029 5853 47031
rect 6222 47083 6278 47085
rect 6222 47031 6224 47083
rect 6224 47031 6276 47083
rect 6276 47031 6278 47083
rect 6222 47029 6278 47031
rect 6654 47083 6710 47085
rect 6654 47031 6656 47083
rect 6656 47031 6708 47083
rect 6708 47031 6710 47083
rect 6654 47029 6710 47031
rect 7036 47060 7092 47062
rect 7036 47008 7038 47060
rect 7038 47008 7090 47060
rect 7090 47008 7092 47060
rect 7036 47006 7092 47008
rect 7308 47060 7364 47062
rect 7308 47008 7310 47060
rect 7310 47008 7362 47060
rect 7362 47008 7364 47060
rect 7308 47006 7364 47008
rect 5797 46709 5853 46711
rect 5797 46657 5799 46709
rect 5799 46657 5851 46709
rect 5851 46657 5853 46709
rect 7036 46665 7092 46667
rect 5797 46655 5853 46657
rect 6222 46651 6278 46653
rect 6222 46599 6224 46651
rect 6224 46599 6276 46651
rect 6276 46599 6278 46651
rect 6222 46597 6278 46599
rect 6654 46651 6710 46653
rect 6654 46599 6656 46651
rect 6656 46599 6708 46651
rect 6708 46599 6710 46651
rect 7036 46613 7038 46665
rect 7038 46613 7090 46665
rect 7090 46613 7092 46665
rect 7036 46611 7092 46613
rect 7308 46665 7364 46667
rect 7308 46613 7310 46665
rect 7310 46613 7362 46665
rect 7362 46613 7364 46665
rect 7308 46611 7364 46613
rect 6654 46597 6710 46599
rect 5797 46293 5853 46295
rect 5797 46241 5799 46293
rect 5799 46241 5851 46293
rect 5851 46241 5853 46293
rect 5797 46239 5853 46241
rect 6222 46293 6278 46295
rect 6222 46241 6224 46293
rect 6224 46241 6276 46293
rect 6276 46241 6278 46293
rect 6222 46239 6278 46241
rect 6654 46293 6710 46295
rect 6654 46241 6656 46293
rect 6656 46241 6708 46293
rect 6708 46241 6710 46293
rect 6654 46239 6710 46241
rect 7036 46270 7092 46272
rect 7036 46218 7038 46270
rect 7038 46218 7090 46270
rect 7090 46218 7092 46270
rect 7036 46216 7092 46218
rect 7308 46270 7364 46272
rect 7308 46218 7310 46270
rect 7310 46218 7362 46270
rect 7362 46218 7364 46270
rect 7308 46216 7364 46218
rect 5797 45919 5853 45921
rect 5797 45867 5799 45919
rect 5799 45867 5851 45919
rect 5851 45867 5853 45919
rect 7036 45875 7092 45877
rect 5797 45865 5853 45867
rect 6222 45861 6278 45863
rect 6222 45809 6224 45861
rect 6224 45809 6276 45861
rect 6276 45809 6278 45861
rect 6222 45807 6278 45809
rect 6654 45861 6710 45863
rect 6654 45809 6656 45861
rect 6656 45809 6708 45861
rect 6708 45809 6710 45861
rect 7036 45823 7038 45875
rect 7038 45823 7090 45875
rect 7090 45823 7092 45875
rect 7036 45821 7092 45823
rect 7308 45875 7364 45877
rect 7308 45823 7310 45875
rect 7310 45823 7362 45875
rect 7362 45823 7364 45875
rect 7308 45821 7364 45823
rect 6654 45807 6710 45809
rect 5797 45503 5853 45505
rect 5797 45451 5799 45503
rect 5799 45451 5851 45503
rect 5851 45451 5853 45503
rect 5797 45449 5853 45451
rect 6222 45503 6278 45505
rect 6222 45451 6224 45503
rect 6224 45451 6276 45503
rect 6276 45451 6278 45503
rect 6222 45449 6278 45451
rect 6654 45503 6710 45505
rect 6654 45451 6656 45503
rect 6656 45451 6708 45503
rect 6708 45451 6710 45503
rect 6654 45449 6710 45451
rect 7036 45480 7092 45482
rect 7036 45428 7038 45480
rect 7038 45428 7090 45480
rect 7090 45428 7092 45480
rect 7036 45426 7092 45428
rect 7308 45480 7364 45482
rect 7308 45428 7310 45480
rect 7310 45428 7362 45480
rect 7362 45428 7364 45480
rect 7308 45426 7364 45428
rect 5797 45129 5853 45131
rect 5797 45077 5799 45129
rect 5799 45077 5851 45129
rect 5851 45077 5853 45129
rect 7036 45085 7092 45087
rect 5797 45075 5853 45077
rect 6222 45071 6278 45073
rect 6222 45019 6224 45071
rect 6224 45019 6276 45071
rect 6276 45019 6278 45071
rect 6222 45017 6278 45019
rect 6654 45071 6710 45073
rect 6654 45019 6656 45071
rect 6656 45019 6708 45071
rect 6708 45019 6710 45071
rect 7036 45033 7038 45085
rect 7038 45033 7090 45085
rect 7090 45033 7092 45085
rect 7036 45031 7092 45033
rect 7308 45085 7364 45087
rect 7308 45033 7310 45085
rect 7310 45033 7362 45085
rect 7362 45033 7364 45085
rect 7308 45031 7364 45033
rect 6654 45017 6710 45019
rect 5797 44713 5853 44715
rect 5797 44661 5799 44713
rect 5799 44661 5851 44713
rect 5851 44661 5853 44713
rect 5797 44659 5853 44661
rect 6222 44713 6278 44715
rect 6222 44661 6224 44713
rect 6224 44661 6276 44713
rect 6276 44661 6278 44713
rect 6222 44659 6278 44661
rect 6654 44713 6710 44715
rect 6654 44661 6656 44713
rect 6656 44661 6708 44713
rect 6708 44661 6710 44713
rect 6654 44659 6710 44661
rect 7036 44690 7092 44692
rect 7036 44638 7038 44690
rect 7038 44638 7090 44690
rect 7090 44638 7092 44690
rect 7036 44636 7092 44638
rect 7308 44690 7364 44692
rect 7308 44638 7310 44690
rect 7310 44638 7362 44690
rect 7362 44638 7364 44690
rect 7308 44636 7364 44638
rect 5797 44339 5853 44341
rect 5797 44287 5799 44339
rect 5799 44287 5851 44339
rect 5851 44287 5853 44339
rect 7036 44295 7092 44297
rect 5797 44285 5853 44287
rect 6222 44281 6278 44283
rect 6222 44229 6224 44281
rect 6224 44229 6276 44281
rect 6276 44229 6278 44281
rect 6222 44227 6278 44229
rect 6654 44281 6710 44283
rect 6654 44229 6656 44281
rect 6656 44229 6708 44281
rect 6708 44229 6710 44281
rect 7036 44243 7038 44295
rect 7038 44243 7090 44295
rect 7090 44243 7092 44295
rect 7036 44241 7092 44243
rect 7308 44295 7364 44297
rect 7308 44243 7310 44295
rect 7310 44243 7362 44295
rect 7362 44243 7364 44295
rect 7308 44241 7364 44243
rect 6654 44227 6710 44229
rect 5797 43923 5853 43925
rect 5797 43871 5799 43923
rect 5799 43871 5851 43923
rect 5851 43871 5853 43923
rect 5797 43869 5853 43871
rect 6222 43923 6278 43925
rect 6222 43871 6224 43923
rect 6224 43871 6276 43923
rect 6276 43871 6278 43923
rect 6222 43869 6278 43871
rect 6654 43923 6710 43925
rect 6654 43871 6656 43923
rect 6656 43871 6708 43923
rect 6708 43871 6710 43923
rect 6654 43869 6710 43871
rect 7036 43900 7092 43902
rect 7036 43848 7038 43900
rect 7038 43848 7090 43900
rect 7090 43848 7092 43900
rect 7036 43846 7092 43848
rect 7308 43900 7364 43902
rect 7308 43848 7310 43900
rect 7310 43848 7362 43900
rect 7362 43848 7364 43900
rect 7308 43846 7364 43848
rect 5797 43549 5853 43551
rect 5797 43497 5799 43549
rect 5799 43497 5851 43549
rect 5851 43497 5853 43549
rect 7036 43505 7092 43507
rect 5797 43495 5853 43497
rect 6222 43491 6278 43493
rect 6222 43439 6224 43491
rect 6224 43439 6276 43491
rect 6276 43439 6278 43491
rect 6222 43437 6278 43439
rect 6654 43491 6710 43493
rect 6654 43439 6656 43491
rect 6656 43439 6708 43491
rect 6708 43439 6710 43491
rect 7036 43453 7038 43505
rect 7038 43453 7090 43505
rect 7090 43453 7092 43505
rect 7036 43451 7092 43453
rect 7308 43505 7364 43507
rect 7308 43453 7310 43505
rect 7310 43453 7362 43505
rect 7362 43453 7364 43505
rect 7308 43451 7364 43453
rect 6654 43437 6710 43439
rect 5797 43133 5853 43135
rect 5797 43081 5799 43133
rect 5799 43081 5851 43133
rect 5851 43081 5853 43133
rect 5797 43079 5853 43081
rect 6222 43133 6278 43135
rect 6222 43081 6224 43133
rect 6224 43081 6276 43133
rect 6276 43081 6278 43133
rect 6222 43079 6278 43081
rect 6654 43133 6710 43135
rect 6654 43081 6656 43133
rect 6656 43081 6708 43133
rect 6708 43081 6710 43133
rect 6654 43079 6710 43081
rect 7036 43110 7092 43112
rect 7036 43058 7038 43110
rect 7038 43058 7090 43110
rect 7090 43058 7092 43110
rect 7036 43056 7092 43058
rect 7308 43110 7364 43112
rect 7308 43058 7310 43110
rect 7310 43058 7362 43110
rect 7362 43058 7364 43110
rect 7308 43056 7364 43058
rect 5797 42759 5853 42761
rect 5797 42707 5799 42759
rect 5799 42707 5851 42759
rect 5851 42707 5853 42759
rect 7036 42715 7092 42717
rect 5797 42705 5853 42707
rect 6222 42701 6278 42703
rect 6222 42649 6224 42701
rect 6224 42649 6276 42701
rect 6276 42649 6278 42701
rect 6222 42647 6278 42649
rect 6654 42701 6710 42703
rect 6654 42649 6656 42701
rect 6656 42649 6708 42701
rect 6708 42649 6710 42701
rect 7036 42663 7038 42715
rect 7038 42663 7090 42715
rect 7090 42663 7092 42715
rect 7036 42661 7092 42663
rect 7308 42715 7364 42717
rect 7308 42663 7310 42715
rect 7310 42663 7362 42715
rect 7362 42663 7364 42715
rect 7308 42661 7364 42663
rect 6654 42647 6710 42649
rect 5797 42343 5853 42345
rect 5797 42291 5799 42343
rect 5799 42291 5851 42343
rect 5851 42291 5853 42343
rect 5797 42289 5853 42291
rect 6222 42343 6278 42345
rect 6222 42291 6224 42343
rect 6224 42291 6276 42343
rect 6276 42291 6278 42343
rect 6222 42289 6278 42291
rect 6654 42343 6710 42345
rect 6654 42291 6656 42343
rect 6656 42291 6708 42343
rect 6708 42291 6710 42343
rect 6654 42289 6710 42291
rect 7036 42320 7092 42322
rect 7036 42268 7038 42320
rect 7038 42268 7090 42320
rect 7090 42268 7092 42320
rect 7036 42266 7092 42268
rect 7308 42320 7364 42322
rect 7308 42268 7310 42320
rect 7310 42268 7362 42320
rect 7362 42268 7364 42320
rect 7308 42266 7364 42268
rect 5797 41969 5853 41971
rect 5797 41917 5799 41969
rect 5799 41917 5851 41969
rect 5851 41917 5853 41969
rect 7036 41925 7092 41927
rect 5797 41915 5853 41917
rect 6222 41911 6278 41913
rect 6222 41859 6224 41911
rect 6224 41859 6276 41911
rect 6276 41859 6278 41911
rect 6222 41857 6278 41859
rect 6654 41911 6710 41913
rect 6654 41859 6656 41911
rect 6656 41859 6708 41911
rect 6708 41859 6710 41911
rect 7036 41873 7038 41925
rect 7038 41873 7090 41925
rect 7090 41873 7092 41925
rect 7036 41871 7092 41873
rect 7308 41925 7364 41927
rect 7308 41873 7310 41925
rect 7310 41873 7362 41925
rect 7362 41873 7364 41925
rect 7308 41871 7364 41873
rect 6654 41857 6710 41859
rect 5797 41553 5853 41555
rect 5797 41501 5799 41553
rect 5799 41501 5851 41553
rect 5851 41501 5853 41553
rect 5797 41499 5853 41501
rect 6222 41553 6278 41555
rect 6222 41501 6224 41553
rect 6224 41501 6276 41553
rect 6276 41501 6278 41553
rect 6222 41499 6278 41501
rect 6654 41553 6710 41555
rect 6654 41501 6656 41553
rect 6656 41501 6708 41553
rect 6708 41501 6710 41553
rect 6654 41499 6710 41501
rect 7036 41530 7092 41532
rect 7036 41478 7038 41530
rect 7038 41478 7090 41530
rect 7090 41478 7092 41530
rect 7036 41476 7092 41478
rect 7308 41530 7364 41532
rect 7308 41478 7310 41530
rect 7310 41478 7362 41530
rect 7362 41478 7364 41530
rect 7308 41476 7364 41478
rect 5797 41179 5853 41181
rect 5797 41127 5799 41179
rect 5799 41127 5851 41179
rect 5851 41127 5853 41179
rect 7036 41135 7092 41137
rect 5797 41125 5853 41127
rect 6222 41121 6278 41123
rect 6222 41069 6224 41121
rect 6224 41069 6276 41121
rect 6276 41069 6278 41121
rect 6222 41067 6278 41069
rect 6654 41121 6710 41123
rect 6654 41069 6656 41121
rect 6656 41069 6708 41121
rect 6708 41069 6710 41121
rect 7036 41083 7038 41135
rect 7038 41083 7090 41135
rect 7090 41083 7092 41135
rect 7036 41081 7092 41083
rect 7308 41135 7364 41137
rect 7308 41083 7310 41135
rect 7310 41083 7362 41135
rect 7362 41083 7364 41135
rect 7308 41081 7364 41083
rect 6654 41067 6710 41069
rect 5797 40763 5853 40765
rect 5797 40711 5799 40763
rect 5799 40711 5851 40763
rect 5851 40711 5853 40763
rect 5797 40709 5853 40711
rect 6222 40763 6278 40765
rect 6222 40711 6224 40763
rect 6224 40711 6276 40763
rect 6276 40711 6278 40763
rect 6222 40709 6278 40711
rect 6654 40763 6710 40765
rect 6654 40711 6656 40763
rect 6656 40711 6708 40763
rect 6708 40711 6710 40763
rect 6654 40709 6710 40711
rect 7036 40740 7092 40742
rect 7036 40688 7038 40740
rect 7038 40688 7090 40740
rect 7090 40688 7092 40740
rect 7036 40686 7092 40688
rect 7308 40740 7364 40742
rect 7308 40688 7310 40740
rect 7310 40688 7362 40740
rect 7362 40688 7364 40740
rect 7308 40686 7364 40688
rect 5797 40389 5853 40391
rect 5797 40337 5799 40389
rect 5799 40337 5851 40389
rect 5851 40337 5853 40389
rect 7036 40345 7092 40347
rect 5797 40335 5853 40337
rect 6222 40331 6278 40333
rect 6222 40279 6224 40331
rect 6224 40279 6276 40331
rect 6276 40279 6278 40331
rect 6222 40277 6278 40279
rect 6654 40331 6710 40333
rect 6654 40279 6656 40331
rect 6656 40279 6708 40331
rect 6708 40279 6710 40331
rect 7036 40293 7038 40345
rect 7038 40293 7090 40345
rect 7090 40293 7092 40345
rect 7036 40291 7092 40293
rect 7308 40345 7364 40347
rect 7308 40293 7310 40345
rect 7310 40293 7362 40345
rect 7362 40293 7364 40345
rect 7308 40291 7364 40293
rect 6654 40277 6710 40279
rect 5797 39973 5853 39975
rect 5797 39921 5799 39973
rect 5799 39921 5851 39973
rect 5851 39921 5853 39973
rect 5797 39919 5853 39921
rect 6222 39973 6278 39975
rect 6222 39921 6224 39973
rect 6224 39921 6276 39973
rect 6276 39921 6278 39973
rect 6222 39919 6278 39921
rect 6654 39973 6710 39975
rect 6654 39921 6656 39973
rect 6656 39921 6708 39973
rect 6708 39921 6710 39973
rect 6654 39919 6710 39921
rect 7036 39950 7092 39952
rect 7036 39898 7038 39950
rect 7038 39898 7090 39950
rect 7090 39898 7092 39950
rect 7036 39896 7092 39898
rect 7308 39950 7364 39952
rect 7308 39898 7310 39950
rect 7310 39898 7362 39950
rect 7362 39898 7364 39950
rect 7308 39896 7364 39898
rect 5797 39599 5853 39601
rect 5797 39547 5799 39599
rect 5799 39547 5851 39599
rect 5851 39547 5853 39599
rect 7036 39555 7092 39557
rect 5797 39545 5853 39547
rect 6222 39541 6278 39543
rect 6222 39489 6224 39541
rect 6224 39489 6276 39541
rect 6276 39489 6278 39541
rect 6222 39487 6278 39489
rect 6654 39541 6710 39543
rect 6654 39489 6656 39541
rect 6656 39489 6708 39541
rect 6708 39489 6710 39541
rect 7036 39503 7038 39555
rect 7038 39503 7090 39555
rect 7090 39503 7092 39555
rect 7036 39501 7092 39503
rect 7308 39555 7364 39557
rect 7308 39503 7310 39555
rect 7310 39503 7362 39555
rect 7362 39503 7364 39555
rect 7308 39501 7364 39503
rect 6654 39487 6710 39489
rect 5797 39183 5853 39185
rect 5797 39131 5799 39183
rect 5799 39131 5851 39183
rect 5851 39131 5853 39183
rect 5797 39129 5853 39131
rect 6222 39183 6278 39185
rect 6222 39131 6224 39183
rect 6224 39131 6276 39183
rect 6276 39131 6278 39183
rect 6222 39129 6278 39131
rect 6654 39183 6710 39185
rect 6654 39131 6656 39183
rect 6656 39131 6708 39183
rect 6708 39131 6710 39183
rect 6654 39129 6710 39131
rect 7036 39160 7092 39162
rect 7036 39108 7038 39160
rect 7038 39108 7090 39160
rect 7090 39108 7092 39160
rect 7036 39106 7092 39108
rect 7308 39160 7364 39162
rect 7308 39108 7310 39160
rect 7310 39108 7362 39160
rect 7362 39108 7364 39160
rect 7308 39106 7364 39108
rect 5797 38809 5853 38811
rect 5797 38757 5799 38809
rect 5799 38757 5851 38809
rect 5851 38757 5853 38809
rect 7036 38765 7092 38767
rect 5797 38755 5853 38757
rect 6222 38751 6278 38753
rect 6222 38699 6224 38751
rect 6224 38699 6276 38751
rect 6276 38699 6278 38751
rect 6222 38697 6278 38699
rect 6654 38751 6710 38753
rect 6654 38699 6656 38751
rect 6656 38699 6708 38751
rect 6708 38699 6710 38751
rect 7036 38713 7038 38765
rect 7038 38713 7090 38765
rect 7090 38713 7092 38765
rect 7036 38711 7092 38713
rect 7308 38765 7364 38767
rect 7308 38713 7310 38765
rect 7310 38713 7362 38765
rect 7362 38713 7364 38765
rect 7308 38711 7364 38713
rect 6654 38697 6710 38699
rect 5797 38393 5853 38395
rect 5797 38341 5799 38393
rect 5799 38341 5851 38393
rect 5851 38341 5853 38393
rect 5797 38339 5853 38341
rect 6222 38393 6278 38395
rect 6222 38341 6224 38393
rect 6224 38341 6276 38393
rect 6276 38341 6278 38393
rect 6222 38339 6278 38341
rect 6654 38393 6710 38395
rect 6654 38341 6656 38393
rect 6656 38341 6708 38393
rect 6708 38341 6710 38393
rect 6654 38339 6710 38341
rect 7036 38370 7092 38372
rect 7036 38318 7038 38370
rect 7038 38318 7090 38370
rect 7090 38318 7092 38370
rect 7036 38316 7092 38318
rect 7308 38370 7364 38372
rect 7308 38318 7310 38370
rect 7310 38318 7362 38370
rect 7362 38318 7364 38370
rect 7308 38316 7364 38318
rect 5797 38019 5853 38021
rect 5797 37967 5799 38019
rect 5799 37967 5851 38019
rect 5851 37967 5853 38019
rect 7036 37975 7092 37977
rect 5797 37965 5853 37967
rect 6222 37961 6278 37963
rect 6222 37909 6224 37961
rect 6224 37909 6276 37961
rect 6276 37909 6278 37961
rect 6222 37907 6278 37909
rect 6654 37961 6710 37963
rect 6654 37909 6656 37961
rect 6656 37909 6708 37961
rect 6708 37909 6710 37961
rect 7036 37923 7038 37975
rect 7038 37923 7090 37975
rect 7090 37923 7092 37975
rect 7036 37921 7092 37923
rect 7308 37975 7364 37977
rect 7308 37923 7310 37975
rect 7310 37923 7362 37975
rect 7362 37923 7364 37975
rect 7308 37921 7364 37923
rect 6654 37907 6710 37909
rect 5797 37603 5853 37605
rect 5797 37551 5799 37603
rect 5799 37551 5851 37603
rect 5851 37551 5853 37603
rect 5797 37549 5853 37551
rect 6222 37603 6278 37605
rect 6222 37551 6224 37603
rect 6224 37551 6276 37603
rect 6276 37551 6278 37603
rect 6222 37549 6278 37551
rect 6654 37603 6710 37605
rect 6654 37551 6656 37603
rect 6656 37551 6708 37603
rect 6708 37551 6710 37603
rect 6654 37549 6710 37551
rect 7036 37580 7092 37582
rect 7036 37528 7038 37580
rect 7038 37528 7090 37580
rect 7090 37528 7092 37580
rect 7036 37526 7092 37528
rect 7308 37580 7364 37582
rect 7308 37528 7310 37580
rect 7310 37528 7362 37580
rect 7362 37528 7364 37580
rect 7308 37526 7364 37528
rect 5797 37229 5853 37231
rect 5797 37177 5799 37229
rect 5799 37177 5851 37229
rect 5851 37177 5853 37229
rect 7036 37185 7092 37187
rect 5797 37175 5853 37177
rect 6222 37171 6278 37173
rect 6222 37119 6224 37171
rect 6224 37119 6276 37171
rect 6276 37119 6278 37171
rect 6222 37117 6278 37119
rect 6654 37171 6710 37173
rect 6654 37119 6656 37171
rect 6656 37119 6708 37171
rect 6708 37119 6710 37171
rect 7036 37133 7038 37185
rect 7038 37133 7090 37185
rect 7090 37133 7092 37185
rect 7036 37131 7092 37133
rect 7308 37185 7364 37187
rect 7308 37133 7310 37185
rect 7310 37133 7362 37185
rect 7362 37133 7364 37185
rect 7308 37131 7364 37133
rect 6654 37117 6710 37119
rect 5797 36813 5853 36815
rect 5797 36761 5799 36813
rect 5799 36761 5851 36813
rect 5851 36761 5853 36813
rect 5797 36759 5853 36761
rect 6222 36813 6278 36815
rect 6222 36761 6224 36813
rect 6224 36761 6276 36813
rect 6276 36761 6278 36813
rect 6222 36759 6278 36761
rect 6654 36813 6710 36815
rect 6654 36761 6656 36813
rect 6656 36761 6708 36813
rect 6708 36761 6710 36813
rect 6654 36759 6710 36761
rect 7036 36790 7092 36792
rect 7036 36738 7038 36790
rect 7038 36738 7090 36790
rect 7090 36738 7092 36790
rect 7036 36736 7092 36738
rect 7308 36790 7364 36792
rect 7308 36738 7310 36790
rect 7310 36738 7362 36790
rect 7362 36738 7364 36790
rect 7308 36736 7364 36738
rect 5797 36439 5853 36441
rect 5797 36387 5799 36439
rect 5799 36387 5851 36439
rect 5851 36387 5853 36439
rect 7036 36395 7092 36397
rect 5797 36385 5853 36387
rect 6222 36381 6278 36383
rect 6222 36329 6224 36381
rect 6224 36329 6276 36381
rect 6276 36329 6278 36381
rect 6222 36327 6278 36329
rect 6654 36381 6710 36383
rect 6654 36329 6656 36381
rect 6656 36329 6708 36381
rect 6708 36329 6710 36381
rect 7036 36343 7038 36395
rect 7038 36343 7090 36395
rect 7090 36343 7092 36395
rect 7036 36341 7092 36343
rect 7308 36395 7364 36397
rect 7308 36343 7310 36395
rect 7310 36343 7362 36395
rect 7362 36343 7364 36395
rect 7308 36341 7364 36343
rect 6654 36327 6710 36329
rect 5797 36023 5853 36025
rect 5797 35971 5799 36023
rect 5799 35971 5851 36023
rect 5851 35971 5853 36023
rect 5797 35969 5853 35971
rect 6222 36023 6278 36025
rect 6222 35971 6224 36023
rect 6224 35971 6276 36023
rect 6276 35971 6278 36023
rect 6222 35969 6278 35971
rect 6654 36023 6710 36025
rect 6654 35971 6656 36023
rect 6656 35971 6708 36023
rect 6708 35971 6710 36023
rect 6654 35969 6710 35971
rect 7036 36000 7092 36002
rect 7036 35948 7038 36000
rect 7038 35948 7090 36000
rect 7090 35948 7092 36000
rect 7036 35946 7092 35948
rect 7308 36000 7364 36002
rect 7308 35948 7310 36000
rect 7310 35948 7362 36000
rect 7362 35948 7364 36000
rect 7308 35946 7364 35948
rect 5797 35649 5853 35651
rect 5797 35597 5799 35649
rect 5799 35597 5851 35649
rect 5851 35597 5853 35649
rect 7036 35605 7092 35607
rect 5797 35595 5853 35597
rect 6222 35591 6278 35593
rect 6222 35539 6224 35591
rect 6224 35539 6276 35591
rect 6276 35539 6278 35591
rect 6222 35537 6278 35539
rect 6654 35591 6710 35593
rect 6654 35539 6656 35591
rect 6656 35539 6708 35591
rect 6708 35539 6710 35591
rect 7036 35553 7038 35605
rect 7038 35553 7090 35605
rect 7090 35553 7092 35605
rect 7036 35551 7092 35553
rect 7308 35605 7364 35607
rect 7308 35553 7310 35605
rect 7310 35553 7362 35605
rect 7362 35553 7364 35605
rect 7308 35551 7364 35553
rect 6654 35537 6710 35539
rect 5797 35233 5853 35235
rect 5797 35181 5799 35233
rect 5799 35181 5851 35233
rect 5851 35181 5853 35233
rect 5797 35179 5853 35181
rect 6222 35233 6278 35235
rect 6222 35181 6224 35233
rect 6224 35181 6276 35233
rect 6276 35181 6278 35233
rect 6222 35179 6278 35181
rect 6654 35233 6710 35235
rect 6654 35181 6656 35233
rect 6656 35181 6708 35233
rect 6708 35181 6710 35233
rect 6654 35179 6710 35181
rect 7036 35210 7092 35212
rect 7036 35158 7038 35210
rect 7038 35158 7090 35210
rect 7090 35158 7092 35210
rect 7036 35156 7092 35158
rect 7308 35210 7364 35212
rect 7308 35158 7310 35210
rect 7310 35158 7362 35210
rect 7362 35158 7364 35210
rect 7308 35156 7364 35158
rect 5797 34859 5853 34861
rect 5797 34807 5799 34859
rect 5799 34807 5851 34859
rect 5851 34807 5853 34859
rect 7036 34815 7092 34817
rect 5797 34805 5853 34807
rect 6222 34801 6278 34803
rect 6222 34749 6224 34801
rect 6224 34749 6276 34801
rect 6276 34749 6278 34801
rect 6222 34747 6278 34749
rect 6654 34801 6710 34803
rect 6654 34749 6656 34801
rect 6656 34749 6708 34801
rect 6708 34749 6710 34801
rect 7036 34763 7038 34815
rect 7038 34763 7090 34815
rect 7090 34763 7092 34815
rect 7036 34761 7092 34763
rect 7308 34815 7364 34817
rect 7308 34763 7310 34815
rect 7310 34763 7362 34815
rect 7362 34763 7364 34815
rect 7308 34761 7364 34763
rect 6654 34747 6710 34749
rect 5797 34443 5853 34445
rect 5797 34391 5799 34443
rect 5799 34391 5851 34443
rect 5851 34391 5853 34443
rect 5797 34389 5853 34391
rect 6222 34443 6278 34445
rect 6222 34391 6224 34443
rect 6224 34391 6276 34443
rect 6276 34391 6278 34443
rect 6222 34389 6278 34391
rect 6654 34443 6710 34445
rect 6654 34391 6656 34443
rect 6656 34391 6708 34443
rect 6708 34391 6710 34443
rect 6654 34389 6710 34391
rect 7036 34420 7092 34422
rect 7036 34368 7038 34420
rect 7038 34368 7090 34420
rect 7090 34368 7092 34420
rect 7036 34366 7092 34368
rect 7308 34420 7364 34422
rect 7308 34368 7310 34420
rect 7310 34368 7362 34420
rect 7362 34368 7364 34420
rect 7308 34366 7364 34368
rect 5797 34069 5853 34071
rect 5797 34017 5799 34069
rect 5799 34017 5851 34069
rect 5851 34017 5853 34069
rect 7036 34025 7092 34027
rect 5797 34015 5853 34017
rect 6222 34011 6278 34013
rect 6222 33959 6224 34011
rect 6224 33959 6276 34011
rect 6276 33959 6278 34011
rect 6222 33957 6278 33959
rect 6654 34011 6710 34013
rect 6654 33959 6656 34011
rect 6656 33959 6708 34011
rect 6708 33959 6710 34011
rect 7036 33973 7038 34025
rect 7038 33973 7090 34025
rect 7090 33973 7092 34025
rect 7036 33971 7092 33973
rect 7308 34025 7364 34027
rect 7308 33973 7310 34025
rect 7310 33973 7362 34025
rect 7362 33973 7364 34025
rect 7308 33971 7364 33973
rect 6654 33957 6710 33959
rect 5797 33653 5853 33655
rect 5797 33601 5799 33653
rect 5799 33601 5851 33653
rect 5851 33601 5853 33653
rect 5797 33599 5853 33601
rect 6222 33653 6278 33655
rect 6222 33601 6224 33653
rect 6224 33601 6276 33653
rect 6276 33601 6278 33653
rect 6222 33599 6278 33601
rect 6654 33653 6710 33655
rect 6654 33601 6656 33653
rect 6656 33601 6708 33653
rect 6708 33601 6710 33653
rect 6654 33599 6710 33601
rect 7036 33630 7092 33632
rect 7036 33578 7038 33630
rect 7038 33578 7090 33630
rect 7090 33578 7092 33630
rect 7036 33576 7092 33578
rect 7308 33630 7364 33632
rect 7308 33578 7310 33630
rect 7310 33578 7362 33630
rect 7362 33578 7364 33630
rect 7308 33576 7364 33578
rect 5797 33279 5853 33281
rect 5797 33227 5799 33279
rect 5799 33227 5851 33279
rect 5851 33227 5853 33279
rect 7036 33235 7092 33237
rect 5797 33225 5853 33227
rect 6222 33221 6278 33223
rect 6222 33169 6224 33221
rect 6224 33169 6276 33221
rect 6276 33169 6278 33221
rect 6222 33167 6278 33169
rect 6654 33221 6710 33223
rect 6654 33169 6656 33221
rect 6656 33169 6708 33221
rect 6708 33169 6710 33221
rect 7036 33183 7038 33235
rect 7038 33183 7090 33235
rect 7090 33183 7092 33235
rect 7036 33181 7092 33183
rect 7308 33235 7364 33237
rect 7308 33183 7310 33235
rect 7310 33183 7362 33235
rect 7362 33183 7364 33235
rect 7308 33181 7364 33183
rect 6654 33167 6710 33169
rect 5797 32863 5853 32865
rect 5797 32811 5799 32863
rect 5799 32811 5851 32863
rect 5851 32811 5853 32863
rect 5797 32809 5853 32811
rect 6222 32863 6278 32865
rect 6222 32811 6224 32863
rect 6224 32811 6276 32863
rect 6276 32811 6278 32863
rect 6222 32809 6278 32811
rect 6654 32863 6710 32865
rect 6654 32811 6656 32863
rect 6656 32811 6708 32863
rect 6708 32811 6710 32863
rect 6654 32809 6710 32811
rect 7036 32840 7092 32842
rect 7036 32788 7038 32840
rect 7038 32788 7090 32840
rect 7090 32788 7092 32840
rect 7036 32786 7092 32788
rect 7308 32840 7364 32842
rect 7308 32788 7310 32840
rect 7310 32788 7362 32840
rect 7362 32788 7364 32840
rect 7308 32786 7364 32788
rect 5797 32489 5853 32491
rect 5797 32437 5799 32489
rect 5799 32437 5851 32489
rect 5851 32437 5853 32489
rect 7036 32445 7092 32447
rect 5797 32435 5853 32437
rect 6222 32431 6278 32433
rect 6222 32379 6224 32431
rect 6224 32379 6276 32431
rect 6276 32379 6278 32431
rect 6222 32377 6278 32379
rect 6654 32431 6710 32433
rect 6654 32379 6656 32431
rect 6656 32379 6708 32431
rect 6708 32379 6710 32431
rect 7036 32393 7038 32445
rect 7038 32393 7090 32445
rect 7090 32393 7092 32445
rect 7036 32391 7092 32393
rect 7308 32445 7364 32447
rect 7308 32393 7310 32445
rect 7310 32393 7362 32445
rect 7362 32393 7364 32445
rect 7308 32391 7364 32393
rect 6654 32377 6710 32379
rect 5797 32073 5853 32075
rect 5797 32021 5799 32073
rect 5799 32021 5851 32073
rect 5851 32021 5853 32073
rect 5797 32019 5853 32021
rect 6222 32073 6278 32075
rect 6222 32021 6224 32073
rect 6224 32021 6276 32073
rect 6276 32021 6278 32073
rect 6222 32019 6278 32021
rect 6654 32073 6710 32075
rect 6654 32021 6656 32073
rect 6656 32021 6708 32073
rect 6708 32021 6710 32073
rect 6654 32019 6710 32021
rect 7036 32050 7092 32052
rect 7036 31998 7038 32050
rect 7038 31998 7090 32050
rect 7090 31998 7092 32050
rect 7036 31996 7092 31998
rect 7308 32050 7364 32052
rect 7308 31998 7310 32050
rect 7310 31998 7362 32050
rect 7362 31998 7364 32050
rect 7308 31996 7364 31998
rect 5797 31699 5853 31701
rect 5797 31647 5799 31699
rect 5799 31647 5851 31699
rect 5851 31647 5853 31699
rect 7036 31655 7092 31657
rect 5797 31645 5853 31647
rect 6222 31641 6278 31643
rect 6222 31589 6224 31641
rect 6224 31589 6276 31641
rect 6276 31589 6278 31641
rect 6222 31587 6278 31589
rect 6654 31641 6710 31643
rect 6654 31589 6656 31641
rect 6656 31589 6708 31641
rect 6708 31589 6710 31641
rect 7036 31603 7038 31655
rect 7038 31603 7090 31655
rect 7090 31603 7092 31655
rect 7036 31601 7092 31603
rect 7308 31655 7364 31657
rect 7308 31603 7310 31655
rect 7310 31603 7362 31655
rect 7362 31603 7364 31655
rect 7308 31601 7364 31603
rect 6654 31587 6710 31589
rect 5797 31283 5853 31285
rect 5797 31231 5799 31283
rect 5799 31231 5851 31283
rect 5851 31231 5853 31283
rect 5797 31229 5853 31231
rect 6222 31283 6278 31285
rect 6222 31231 6224 31283
rect 6224 31231 6276 31283
rect 6276 31231 6278 31283
rect 6222 31229 6278 31231
rect 6654 31283 6710 31285
rect 6654 31231 6656 31283
rect 6656 31231 6708 31283
rect 6708 31231 6710 31283
rect 6654 31229 6710 31231
rect 7036 31260 7092 31262
rect 7036 31208 7038 31260
rect 7038 31208 7090 31260
rect 7090 31208 7092 31260
rect 7036 31206 7092 31208
rect 7308 31260 7364 31262
rect 7308 31208 7310 31260
rect 7310 31208 7362 31260
rect 7362 31208 7364 31260
rect 7308 31206 7364 31208
rect 5797 30909 5853 30911
rect 5797 30857 5799 30909
rect 5799 30857 5851 30909
rect 5851 30857 5853 30909
rect 7036 30865 7092 30867
rect 5797 30855 5853 30857
rect 6222 30851 6278 30853
rect 6222 30799 6224 30851
rect 6224 30799 6276 30851
rect 6276 30799 6278 30851
rect 6222 30797 6278 30799
rect 6654 30851 6710 30853
rect 6654 30799 6656 30851
rect 6656 30799 6708 30851
rect 6708 30799 6710 30851
rect 7036 30813 7038 30865
rect 7038 30813 7090 30865
rect 7090 30813 7092 30865
rect 7036 30811 7092 30813
rect 7308 30865 7364 30867
rect 7308 30813 7310 30865
rect 7310 30813 7362 30865
rect 7362 30813 7364 30865
rect 7308 30811 7364 30813
rect 6654 30797 6710 30799
rect 5797 30493 5853 30495
rect 5797 30441 5799 30493
rect 5799 30441 5851 30493
rect 5851 30441 5853 30493
rect 5797 30439 5853 30441
rect 6222 30493 6278 30495
rect 6222 30441 6224 30493
rect 6224 30441 6276 30493
rect 6276 30441 6278 30493
rect 6222 30439 6278 30441
rect 6654 30493 6710 30495
rect 6654 30441 6656 30493
rect 6656 30441 6708 30493
rect 6708 30441 6710 30493
rect 6654 30439 6710 30441
rect 7036 30470 7092 30472
rect 7036 30418 7038 30470
rect 7038 30418 7090 30470
rect 7090 30418 7092 30470
rect 7036 30416 7092 30418
rect 7308 30470 7364 30472
rect 7308 30418 7310 30470
rect 7310 30418 7362 30470
rect 7362 30418 7364 30470
rect 7308 30416 7364 30418
rect 5797 30119 5853 30121
rect 5797 30067 5799 30119
rect 5799 30067 5851 30119
rect 5851 30067 5853 30119
rect 7036 30075 7092 30077
rect 5797 30065 5853 30067
rect 6222 30061 6278 30063
rect 6222 30009 6224 30061
rect 6224 30009 6276 30061
rect 6276 30009 6278 30061
rect 6222 30007 6278 30009
rect 6654 30061 6710 30063
rect 6654 30009 6656 30061
rect 6656 30009 6708 30061
rect 6708 30009 6710 30061
rect 7036 30023 7038 30075
rect 7038 30023 7090 30075
rect 7090 30023 7092 30075
rect 7036 30021 7092 30023
rect 7308 30075 7364 30077
rect 7308 30023 7310 30075
rect 7310 30023 7362 30075
rect 7362 30023 7364 30075
rect 7308 30021 7364 30023
rect 6654 30007 6710 30009
rect 5797 29703 5853 29705
rect 5797 29651 5799 29703
rect 5799 29651 5851 29703
rect 5851 29651 5853 29703
rect 5797 29649 5853 29651
rect 6222 29703 6278 29705
rect 6222 29651 6224 29703
rect 6224 29651 6276 29703
rect 6276 29651 6278 29703
rect 6222 29649 6278 29651
rect 6654 29703 6710 29705
rect 6654 29651 6656 29703
rect 6656 29651 6708 29703
rect 6708 29651 6710 29703
rect 6654 29649 6710 29651
rect 7036 29680 7092 29682
rect 7036 29628 7038 29680
rect 7038 29628 7090 29680
rect 7090 29628 7092 29680
rect 7036 29626 7092 29628
rect 7308 29680 7364 29682
rect 7308 29628 7310 29680
rect 7310 29628 7362 29680
rect 7362 29628 7364 29680
rect 7308 29626 7364 29628
rect 5797 29329 5853 29331
rect 5797 29277 5799 29329
rect 5799 29277 5851 29329
rect 5851 29277 5853 29329
rect 7036 29285 7092 29287
rect 5797 29275 5853 29277
rect 6222 29271 6278 29273
rect 6222 29219 6224 29271
rect 6224 29219 6276 29271
rect 6276 29219 6278 29271
rect 6222 29217 6278 29219
rect 6654 29271 6710 29273
rect 6654 29219 6656 29271
rect 6656 29219 6708 29271
rect 6708 29219 6710 29271
rect 7036 29233 7038 29285
rect 7038 29233 7090 29285
rect 7090 29233 7092 29285
rect 7036 29231 7092 29233
rect 7308 29285 7364 29287
rect 7308 29233 7310 29285
rect 7310 29233 7362 29285
rect 7362 29233 7364 29285
rect 7308 29231 7364 29233
rect 6654 29217 6710 29219
rect 5797 28913 5853 28915
rect 5797 28861 5799 28913
rect 5799 28861 5851 28913
rect 5851 28861 5853 28913
rect 5797 28859 5853 28861
rect 6222 28913 6278 28915
rect 6222 28861 6224 28913
rect 6224 28861 6276 28913
rect 6276 28861 6278 28913
rect 6222 28859 6278 28861
rect 6654 28913 6710 28915
rect 6654 28861 6656 28913
rect 6656 28861 6708 28913
rect 6708 28861 6710 28913
rect 6654 28859 6710 28861
rect 7036 28890 7092 28892
rect 7036 28838 7038 28890
rect 7038 28838 7090 28890
rect 7090 28838 7092 28890
rect 7036 28836 7092 28838
rect 7308 28890 7364 28892
rect 7308 28838 7310 28890
rect 7310 28838 7362 28890
rect 7362 28838 7364 28890
rect 7308 28836 7364 28838
rect 5797 28539 5853 28541
rect 5797 28487 5799 28539
rect 5799 28487 5851 28539
rect 5851 28487 5853 28539
rect 7036 28495 7092 28497
rect 5797 28485 5853 28487
rect 6222 28481 6278 28483
rect 6222 28429 6224 28481
rect 6224 28429 6276 28481
rect 6276 28429 6278 28481
rect 6222 28427 6278 28429
rect 6654 28481 6710 28483
rect 6654 28429 6656 28481
rect 6656 28429 6708 28481
rect 6708 28429 6710 28481
rect 7036 28443 7038 28495
rect 7038 28443 7090 28495
rect 7090 28443 7092 28495
rect 7036 28441 7092 28443
rect 7308 28495 7364 28497
rect 7308 28443 7310 28495
rect 7310 28443 7362 28495
rect 7362 28443 7364 28495
rect 7308 28441 7364 28443
rect 6654 28427 6710 28429
rect 5797 28123 5853 28125
rect 5797 28071 5799 28123
rect 5799 28071 5851 28123
rect 5851 28071 5853 28123
rect 5797 28069 5853 28071
rect 6222 28123 6278 28125
rect 6222 28071 6224 28123
rect 6224 28071 6276 28123
rect 6276 28071 6278 28123
rect 6222 28069 6278 28071
rect 6654 28123 6710 28125
rect 6654 28071 6656 28123
rect 6656 28071 6708 28123
rect 6708 28071 6710 28123
rect 6654 28069 6710 28071
rect 7036 28100 7092 28102
rect 7036 28048 7038 28100
rect 7038 28048 7090 28100
rect 7090 28048 7092 28100
rect 7036 28046 7092 28048
rect 7308 28100 7364 28102
rect 7308 28048 7310 28100
rect 7310 28048 7362 28100
rect 7362 28048 7364 28100
rect 7308 28046 7364 28048
rect 5797 27749 5853 27751
rect 5797 27697 5799 27749
rect 5799 27697 5851 27749
rect 5851 27697 5853 27749
rect 7036 27705 7092 27707
rect 5797 27695 5853 27697
rect 6222 27691 6278 27693
rect 6222 27639 6224 27691
rect 6224 27639 6276 27691
rect 6276 27639 6278 27691
rect 6222 27637 6278 27639
rect 6654 27691 6710 27693
rect 6654 27639 6656 27691
rect 6656 27639 6708 27691
rect 6708 27639 6710 27691
rect 7036 27653 7038 27705
rect 7038 27653 7090 27705
rect 7090 27653 7092 27705
rect 7036 27651 7092 27653
rect 7308 27705 7364 27707
rect 7308 27653 7310 27705
rect 7310 27653 7362 27705
rect 7362 27653 7364 27705
rect 7308 27651 7364 27653
rect 6654 27637 6710 27639
rect 5797 27333 5853 27335
rect 5797 27281 5799 27333
rect 5799 27281 5851 27333
rect 5851 27281 5853 27333
rect 5797 27279 5853 27281
rect 6222 27333 6278 27335
rect 6222 27281 6224 27333
rect 6224 27281 6276 27333
rect 6276 27281 6278 27333
rect 6222 27279 6278 27281
rect 6654 27333 6710 27335
rect 6654 27281 6656 27333
rect 6656 27281 6708 27333
rect 6708 27281 6710 27333
rect 6654 27279 6710 27281
rect 7036 27310 7092 27312
rect 7036 27258 7038 27310
rect 7038 27258 7090 27310
rect 7090 27258 7092 27310
rect 7036 27256 7092 27258
rect 7308 27310 7364 27312
rect 7308 27258 7310 27310
rect 7310 27258 7362 27310
rect 7362 27258 7364 27310
rect 7308 27256 7364 27258
rect 5797 26959 5853 26961
rect 5797 26907 5799 26959
rect 5799 26907 5851 26959
rect 5851 26907 5853 26959
rect 7036 26915 7092 26917
rect 5797 26905 5853 26907
rect 6222 26901 6278 26903
rect 6222 26849 6224 26901
rect 6224 26849 6276 26901
rect 6276 26849 6278 26901
rect 6222 26847 6278 26849
rect 6654 26901 6710 26903
rect 6654 26849 6656 26901
rect 6656 26849 6708 26901
rect 6708 26849 6710 26901
rect 7036 26863 7038 26915
rect 7038 26863 7090 26915
rect 7090 26863 7092 26915
rect 7036 26861 7092 26863
rect 7308 26915 7364 26917
rect 7308 26863 7310 26915
rect 7310 26863 7362 26915
rect 7362 26863 7364 26915
rect 7308 26861 7364 26863
rect 6654 26847 6710 26849
rect 5797 26543 5853 26545
rect 5797 26491 5799 26543
rect 5799 26491 5851 26543
rect 5851 26491 5853 26543
rect 5797 26489 5853 26491
rect 6222 26543 6278 26545
rect 6222 26491 6224 26543
rect 6224 26491 6276 26543
rect 6276 26491 6278 26543
rect 6222 26489 6278 26491
rect 6654 26543 6710 26545
rect 6654 26491 6656 26543
rect 6656 26491 6708 26543
rect 6708 26491 6710 26543
rect 6654 26489 6710 26491
rect 7036 26520 7092 26522
rect 7036 26468 7038 26520
rect 7038 26468 7090 26520
rect 7090 26468 7092 26520
rect 7036 26466 7092 26468
rect 7308 26520 7364 26522
rect 7308 26468 7310 26520
rect 7310 26468 7362 26520
rect 7362 26468 7364 26520
rect 7308 26466 7364 26468
rect 5797 26169 5853 26171
rect 5797 26117 5799 26169
rect 5799 26117 5851 26169
rect 5851 26117 5853 26169
rect 7036 26125 7092 26127
rect 5797 26115 5853 26117
rect 6222 26111 6278 26113
rect 6222 26059 6224 26111
rect 6224 26059 6276 26111
rect 6276 26059 6278 26111
rect 6222 26057 6278 26059
rect 6654 26111 6710 26113
rect 6654 26059 6656 26111
rect 6656 26059 6708 26111
rect 6708 26059 6710 26111
rect 7036 26073 7038 26125
rect 7038 26073 7090 26125
rect 7090 26073 7092 26125
rect 7036 26071 7092 26073
rect 7308 26125 7364 26127
rect 7308 26073 7310 26125
rect 7310 26073 7362 26125
rect 7362 26073 7364 26125
rect 7308 26071 7364 26073
rect 6654 26057 6710 26059
rect 5797 25753 5853 25755
rect 5797 25701 5799 25753
rect 5799 25701 5851 25753
rect 5851 25701 5853 25753
rect 5797 25699 5853 25701
rect 6222 25753 6278 25755
rect 6222 25701 6224 25753
rect 6224 25701 6276 25753
rect 6276 25701 6278 25753
rect 6222 25699 6278 25701
rect 6654 25753 6710 25755
rect 6654 25701 6656 25753
rect 6656 25701 6708 25753
rect 6708 25701 6710 25753
rect 6654 25699 6710 25701
rect 7036 25730 7092 25732
rect 7036 25678 7038 25730
rect 7038 25678 7090 25730
rect 7090 25678 7092 25730
rect 7036 25676 7092 25678
rect 7308 25730 7364 25732
rect 7308 25678 7310 25730
rect 7310 25678 7362 25730
rect 7362 25678 7364 25730
rect 7308 25676 7364 25678
rect 5797 25379 5853 25381
rect 5797 25327 5799 25379
rect 5799 25327 5851 25379
rect 5851 25327 5853 25379
rect 7036 25335 7092 25337
rect 5797 25325 5853 25327
rect 6222 25321 6278 25323
rect 6222 25269 6224 25321
rect 6224 25269 6276 25321
rect 6276 25269 6278 25321
rect 6222 25267 6278 25269
rect 6654 25321 6710 25323
rect 6654 25269 6656 25321
rect 6656 25269 6708 25321
rect 6708 25269 6710 25321
rect 7036 25283 7038 25335
rect 7038 25283 7090 25335
rect 7090 25283 7092 25335
rect 7036 25281 7092 25283
rect 7308 25335 7364 25337
rect 7308 25283 7310 25335
rect 7310 25283 7362 25335
rect 7362 25283 7364 25335
rect 7308 25281 7364 25283
rect 6654 25267 6710 25269
rect 5797 24963 5853 24965
rect 5797 24911 5799 24963
rect 5799 24911 5851 24963
rect 5851 24911 5853 24963
rect 5797 24909 5853 24911
rect 6222 24963 6278 24965
rect 6222 24911 6224 24963
rect 6224 24911 6276 24963
rect 6276 24911 6278 24963
rect 6222 24909 6278 24911
rect 6654 24963 6710 24965
rect 6654 24911 6656 24963
rect 6656 24911 6708 24963
rect 6708 24911 6710 24963
rect 6654 24909 6710 24911
rect 7036 24940 7092 24942
rect 7036 24888 7038 24940
rect 7038 24888 7090 24940
rect 7090 24888 7092 24940
rect 7036 24886 7092 24888
rect 7308 24940 7364 24942
rect 7308 24888 7310 24940
rect 7310 24888 7362 24940
rect 7362 24888 7364 24940
rect 7308 24886 7364 24888
rect 5797 24589 5853 24591
rect 5797 24537 5799 24589
rect 5799 24537 5851 24589
rect 5851 24537 5853 24589
rect 7036 24545 7092 24547
rect 5797 24535 5853 24537
rect 6222 24531 6278 24533
rect 6222 24479 6224 24531
rect 6224 24479 6276 24531
rect 6276 24479 6278 24531
rect 6222 24477 6278 24479
rect 6654 24531 6710 24533
rect 6654 24479 6656 24531
rect 6656 24479 6708 24531
rect 6708 24479 6710 24531
rect 7036 24493 7038 24545
rect 7038 24493 7090 24545
rect 7090 24493 7092 24545
rect 7036 24491 7092 24493
rect 7308 24545 7364 24547
rect 7308 24493 7310 24545
rect 7310 24493 7362 24545
rect 7362 24493 7364 24545
rect 7308 24491 7364 24493
rect 6654 24477 6710 24479
rect 5797 24173 5853 24175
rect 5797 24121 5799 24173
rect 5799 24121 5851 24173
rect 5851 24121 5853 24173
rect 5797 24119 5853 24121
rect 6222 24173 6278 24175
rect 6222 24121 6224 24173
rect 6224 24121 6276 24173
rect 6276 24121 6278 24173
rect 6222 24119 6278 24121
rect 6654 24173 6710 24175
rect 6654 24121 6656 24173
rect 6656 24121 6708 24173
rect 6708 24121 6710 24173
rect 6654 24119 6710 24121
rect 7036 24150 7092 24152
rect 7036 24098 7038 24150
rect 7038 24098 7090 24150
rect 7090 24098 7092 24150
rect 7036 24096 7092 24098
rect 7308 24150 7364 24152
rect 7308 24098 7310 24150
rect 7310 24098 7362 24150
rect 7362 24098 7364 24150
rect 7308 24096 7364 24098
rect 5797 23799 5853 23801
rect 5797 23747 5799 23799
rect 5799 23747 5851 23799
rect 5851 23747 5853 23799
rect 7036 23755 7092 23757
rect 5797 23745 5853 23747
rect 6222 23741 6278 23743
rect 6222 23689 6224 23741
rect 6224 23689 6276 23741
rect 6276 23689 6278 23741
rect 6222 23687 6278 23689
rect 6654 23741 6710 23743
rect 6654 23689 6656 23741
rect 6656 23689 6708 23741
rect 6708 23689 6710 23741
rect 7036 23703 7038 23755
rect 7038 23703 7090 23755
rect 7090 23703 7092 23755
rect 7036 23701 7092 23703
rect 7308 23755 7364 23757
rect 7308 23703 7310 23755
rect 7310 23703 7362 23755
rect 7362 23703 7364 23755
rect 7308 23701 7364 23703
rect 6654 23687 6710 23689
rect 5797 23383 5853 23385
rect 5797 23331 5799 23383
rect 5799 23331 5851 23383
rect 5851 23331 5853 23383
rect 5797 23329 5853 23331
rect 6222 23383 6278 23385
rect 6222 23331 6224 23383
rect 6224 23331 6276 23383
rect 6276 23331 6278 23383
rect 6222 23329 6278 23331
rect 6654 23383 6710 23385
rect 6654 23331 6656 23383
rect 6656 23331 6708 23383
rect 6708 23331 6710 23383
rect 6654 23329 6710 23331
rect 7036 23360 7092 23362
rect 7036 23308 7038 23360
rect 7038 23308 7090 23360
rect 7090 23308 7092 23360
rect 7036 23306 7092 23308
rect 7308 23360 7364 23362
rect 7308 23308 7310 23360
rect 7310 23308 7362 23360
rect 7362 23308 7364 23360
rect 7308 23306 7364 23308
rect 5797 23009 5853 23011
rect 5797 22957 5799 23009
rect 5799 22957 5851 23009
rect 5851 22957 5853 23009
rect 7036 22965 7092 22967
rect 5797 22955 5853 22957
rect 6222 22951 6278 22953
rect 6222 22899 6224 22951
rect 6224 22899 6276 22951
rect 6276 22899 6278 22951
rect 6222 22897 6278 22899
rect 6654 22951 6710 22953
rect 6654 22899 6656 22951
rect 6656 22899 6708 22951
rect 6708 22899 6710 22951
rect 7036 22913 7038 22965
rect 7038 22913 7090 22965
rect 7090 22913 7092 22965
rect 7036 22911 7092 22913
rect 7308 22965 7364 22967
rect 7308 22913 7310 22965
rect 7310 22913 7362 22965
rect 7362 22913 7364 22965
rect 7308 22911 7364 22913
rect 6654 22897 6710 22899
rect 5797 22593 5853 22595
rect 5797 22541 5799 22593
rect 5799 22541 5851 22593
rect 5851 22541 5853 22593
rect 5797 22539 5853 22541
rect 6222 22593 6278 22595
rect 6222 22541 6224 22593
rect 6224 22541 6276 22593
rect 6276 22541 6278 22593
rect 6222 22539 6278 22541
rect 6654 22593 6710 22595
rect 6654 22541 6656 22593
rect 6656 22541 6708 22593
rect 6708 22541 6710 22593
rect 6654 22539 6710 22541
rect 7036 22570 7092 22572
rect 7036 22518 7038 22570
rect 7038 22518 7090 22570
rect 7090 22518 7092 22570
rect 7036 22516 7092 22518
rect 7308 22570 7364 22572
rect 7308 22518 7310 22570
rect 7310 22518 7362 22570
rect 7362 22518 7364 22570
rect 7308 22516 7364 22518
rect 5797 22219 5853 22221
rect 5797 22167 5799 22219
rect 5799 22167 5851 22219
rect 5851 22167 5853 22219
rect 7036 22175 7092 22177
rect 5797 22165 5853 22167
rect 6222 22161 6278 22163
rect 6222 22109 6224 22161
rect 6224 22109 6276 22161
rect 6276 22109 6278 22161
rect 6222 22107 6278 22109
rect 6654 22161 6710 22163
rect 6654 22109 6656 22161
rect 6656 22109 6708 22161
rect 6708 22109 6710 22161
rect 7036 22123 7038 22175
rect 7038 22123 7090 22175
rect 7090 22123 7092 22175
rect 7036 22121 7092 22123
rect 7308 22175 7364 22177
rect 7308 22123 7310 22175
rect 7310 22123 7362 22175
rect 7362 22123 7364 22175
rect 7308 22121 7364 22123
rect 6654 22107 6710 22109
rect 5797 21803 5853 21805
rect 5797 21751 5799 21803
rect 5799 21751 5851 21803
rect 5851 21751 5853 21803
rect 5797 21749 5853 21751
rect 6222 21803 6278 21805
rect 6222 21751 6224 21803
rect 6224 21751 6276 21803
rect 6276 21751 6278 21803
rect 6222 21749 6278 21751
rect 6654 21803 6710 21805
rect 6654 21751 6656 21803
rect 6656 21751 6708 21803
rect 6708 21751 6710 21803
rect 6654 21749 6710 21751
rect 7036 21780 7092 21782
rect 7036 21728 7038 21780
rect 7038 21728 7090 21780
rect 7090 21728 7092 21780
rect 7036 21726 7092 21728
rect 7308 21780 7364 21782
rect 7308 21728 7310 21780
rect 7310 21728 7362 21780
rect 7362 21728 7364 21780
rect 7308 21726 7364 21728
rect 5797 21429 5853 21431
rect 5797 21377 5799 21429
rect 5799 21377 5851 21429
rect 5851 21377 5853 21429
rect 7036 21385 7092 21387
rect 5797 21375 5853 21377
rect 6222 21371 6278 21373
rect 6222 21319 6224 21371
rect 6224 21319 6276 21371
rect 6276 21319 6278 21371
rect 6222 21317 6278 21319
rect 6654 21371 6710 21373
rect 6654 21319 6656 21371
rect 6656 21319 6708 21371
rect 6708 21319 6710 21371
rect 7036 21333 7038 21385
rect 7038 21333 7090 21385
rect 7090 21333 7092 21385
rect 7036 21331 7092 21333
rect 7308 21385 7364 21387
rect 7308 21333 7310 21385
rect 7310 21333 7362 21385
rect 7362 21333 7364 21385
rect 7308 21331 7364 21333
rect 6654 21317 6710 21319
rect 5797 21013 5853 21015
rect 5797 20961 5799 21013
rect 5799 20961 5851 21013
rect 5851 20961 5853 21013
rect 5797 20959 5853 20961
rect 6222 21013 6278 21015
rect 6222 20961 6224 21013
rect 6224 20961 6276 21013
rect 6276 20961 6278 21013
rect 6222 20959 6278 20961
rect 6654 21013 6710 21015
rect 6654 20961 6656 21013
rect 6656 20961 6708 21013
rect 6708 20961 6710 21013
rect 6654 20959 6710 20961
rect 7036 20990 7092 20992
rect 7036 20938 7038 20990
rect 7038 20938 7090 20990
rect 7090 20938 7092 20990
rect 7036 20936 7092 20938
rect 7308 20990 7364 20992
rect 7308 20938 7310 20990
rect 7310 20938 7362 20990
rect 7362 20938 7364 20990
rect 7308 20936 7364 20938
rect 5797 20639 5853 20641
rect 5797 20587 5799 20639
rect 5799 20587 5851 20639
rect 5851 20587 5853 20639
rect 7036 20595 7092 20597
rect 5797 20585 5853 20587
rect 6222 20581 6278 20583
rect 6222 20529 6224 20581
rect 6224 20529 6276 20581
rect 6276 20529 6278 20581
rect 6222 20527 6278 20529
rect 6654 20581 6710 20583
rect 6654 20529 6656 20581
rect 6656 20529 6708 20581
rect 6708 20529 6710 20581
rect 7036 20543 7038 20595
rect 7038 20543 7090 20595
rect 7090 20543 7092 20595
rect 7036 20541 7092 20543
rect 7308 20595 7364 20597
rect 7308 20543 7310 20595
rect 7310 20543 7362 20595
rect 7362 20543 7364 20595
rect 7308 20541 7364 20543
rect 6654 20527 6710 20529
rect 5797 20223 5853 20225
rect 5797 20171 5799 20223
rect 5799 20171 5851 20223
rect 5851 20171 5853 20223
rect 5797 20169 5853 20171
rect 6222 20223 6278 20225
rect 6222 20171 6224 20223
rect 6224 20171 6276 20223
rect 6276 20171 6278 20223
rect 6222 20169 6278 20171
rect 6654 20223 6710 20225
rect 6654 20171 6656 20223
rect 6656 20171 6708 20223
rect 6708 20171 6710 20223
rect 6654 20169 6710 20171
rect 7036 20200 7092 20202
rect 7036 20148 7038 20200
rect 7038 20148 7090 20200
rect 7090 20148 7092 20200
rect 7036 20146 7092 20148
rect 7308 20200 7364 20202
rect 7308 20148 7310 20200
rect 7310 20148 7362 20200
rect 7362 20148 7364 20200
rect 7308 20146 7364 20148
rect 5797 19849 5853 19851
rect 5797 19797 5799 19849
rect 5799 19797 5851 19849
rect 5851 19797 5853 19849
rect 7036 19805 7092 19807
rect 5797 19795 5853 19797
rect 6222 19791 6278 19793
rect 6222 19739 6224 19791
rect 6224 19739 6276 19791
rect 6276 19739 6278 19791
rect 6222 19737 6278 19739
rect 6654 19791 6710 19793
rect 6654 19739 6656 19791
rect 6656 19739 6708 19791
rect 6708 19739 6710 19791
rect 7036 19753 7038 19805
rect 7038 19753 7090 19805
rect 7090 19753 7092 19805
rect 7036 19751 7092 19753
rect 7308 19805 7364 19807
rect 7308 19753 7310 19805
rect 7310 19753 7362 19805
rect 7362 19753 7364 19805
rect 7308 19751 7364 19753
rect 6654 19737 6710 19739
rect 5797 19433 5853 19435
rect 5797 19381 5799 19433
rect 5799 19381 5851 19433
rect 5851 19381 5853 19433
rect 5797 19379 5853 19381
rect 6222 19433 6278 19435
rect 6222 19381 6224 19433
rect 6224 19381 6276 19433
rect 6276 19381 6278 19433
rect 6222 19379 6278 19381
rect 6654 19433 6710 19435
rect 6654 19381 6656 19433
rect 6656 19381 6708 19433
rect 6708 19381 6710 19433
rect 6654 19379 6710 19381
rect 7036 19410 7092 19412
rect 7036 19358 7038 19410
rect 7038 19358 7090 19410
rect 7090 19358 7092 19410
rect 7036 19356 7092 19358
rect 7308 19410 7364 19412
rect 7308 19358 7310 19410
rect 7310 19358 7362 19410
rect 7362 19358 7364 19410
rect 7308 19356 7364 19358
rect 5797 19059 5853 19061
rect 5797 19007 5799 19059
rect 5799 19007 5851 19059
rect 5851 19007 5853 19059
rect 7036 19015 7092 19017
rect 5797 19005 5853 19007
rect 6222 19001 6278 19003
rect 6222 18949 6224 19001
rect 6224 18949 6276 19001
rect 6276 18949 6278 19001
rect 6222 18947 6278 18949
rect 6654 19001 6710 19003
rect 6654 18949 6656 19001
rect 6656 18949 6708 19001
rect 6708 18949 6710 19001
rect 7036 18963 7038 19015
rect 7038 18963 7090 19015
rect 7090 18963 7092 19015
rect 7036 18961 7092 18963
rect 7308 19015 7364 19017
rect 7308 18963 7310 19015
rect 7310 18963 7362 19015
rect 7362 18963 7364 19015
rect 7308 18961 7364 18963
rect 6654 18947 6710 18949
rect 5797 18643 5853 18645
rect 5797 18591 5799 18643
rect 5799 18591 5851 18643
rect 5851 18591 5853 18643
rect 5797 18589 5853 18591
rect 6222 18643 6278 18645
rect 6222 18591 6224 18643
rect 6224 18591 6276 18643
rect 6276 18591 6278 18643
rect 6222 18589 6278 18591
rect 6654 18643 6710 18645
rect 6654 18591 6656 18643
rect 6656 18591 6708 18643
rect 6708 18591 6710 18643
rect 6654 18589 6710 18591
rect 7036 18620 7092 18622
rect 7036 18568 7038 18620
rect 7038 18568 7090 18620
rect 7090 18568 7092 18620
rect 7036 18566 7092 18568
rect 7308 18620 7364 18622
rect 7308 18568 7310 18620
rect 7310 18568 7362 18620
rect 7362 18568 7364 18620
rect 7308 18566 7364 18568
rect 5797 18269 5853 18271
rect 5797 18217 5799 18269
rect 5799 18217 5851 18269
rect 5851 18217 5853 18269
rect 7036 18225 7092 18227
rect 5797 18215 5853 18217
rect 6222 18211 6278 18213
rect 6222 18159 6224 18211
rect 6224 18159 6276 18211
rect 6276 18159 6278 18211
rect 6222 18157 6278 18159
rect 6654 18211 6710 18213
rect 6654 18159 6656 18211
rect 6656 18159 6708 18211
rect 6708 18159 6710 18211
rect 7036 18173 7038 18225
rect 7038 18173 7090 18225
rect 7090 18173 7092 18225
rect 7036 18171 7092 18173
rect 7308 18225 7364 18227
rect 7308 18173 7310 18225
rect 7310 18173 7362 18225
rect 7362 18173 7364 18225
rect 7308 18171 7364 18173
rect 6654 18157 6710 18159
rect 5797 17853 5853 17855
rect 5797 17801 5799 17853
rect 5799 17801 5851 17853
rect 5851 17801 5853 17853
rect 5797 17799 5853 17801
rect 6222 17853 6278 17855
rect 6222 17801 6224 17853
rect 6224 17801 6276 17853
rect 6276 17801 6278 17853
rect 6222 17799 6278 17801
rect 6654 17853 6710 17855
rect 6654 17801 6656 17853
rect 6656 17801 6708 17853
rect 6708 17801 6710 17853
rect 6654 17799 6710 17801
rect 7036 17830 7092 17832
rect 7036 17778 7038 17830
rect 7038 17778 7090 17830
rect 7090 17778 7092 17830
rect 7036 17776 7092 17778
rect 7308 17830 7364 17832
rect 7308 17778 7310 17830
rect 7310 17778 7362 17830
rect 7362 17778 7364 17830
rect 7308 17776 7364 17778
rect 5797 17479 5853 17481
rect 5797 17427 5799 17479
rect 5799 17427 5851 17479
rect 5851 17427 5853 17479
rect 7036 17435 7092 17437
rect 5797 17425 5853 17427
rect 6222 17421 6278 17423
rect 6222 17369 6224 17421
rect 6224 17369 6276 17421
rect 6276 17369 6278 17421
rect 6222 17367 6278 17369
rect 6654 17421 6710 17423
rect 6654 17369 6656 17421
rect 6656 17369 6708 17421
rect 6708 17369 6710 17421
rect 7036 17383 7038 17435
rect 7038 17383 7090 17435
rect 7090 17383 7092 17435
rect 7036 17381 7092 17383
rect 7308 17435 7364 17437
rect 7308 17383 7310 17435
rect 7310 17383 7362 17435
rect 7362 17383 7364 17435
rect 7308 17381 7364 17383
rect 6654 17367 6710 17369
rect 5797 17063 5853 17065
rect 5797 17011 5799 17063
rect 5799 17011 5851 17063
rect 5851 17011 5853 17063
rect 5797 17009 5853 17011
rect 6222 17063 6278 17065
rect 6222 17011 6224 17063
rect 6224 17011 6276 17063
rect 6276 17011 6278 17063
rect 6222 17009 6278 17011
rect 6654 17063 6710 17065
rect 6654 17011 6656 17063
rect 6656 17011 6708 17063
rect 6708 17011 6710 17063
rect 6654 17009 6710 17011
rect 7036 17040 7092 17042
rect 7036 16988 7038 17040
rect 7038 16988 7090 17040
rect 7090 16988 7092 17040
rect 7036 16986 7092 16988
rect 7308 17040 7364 17042
rect 7308 16988 7310 17040
rect 7310 16988 7362 17040
rect 7362 16988 7364 17040
rect 7308 16986 7364 16988
rect 5797 16689 5853 16691
rect 5797 16637 5799 16689
rect 5799 16637 5851 16689
rect 5851 16637 5853 16689
rect 7036 16645 7092 16647
rect 5797 16635 5853 16637
rect 6222 16631 6278 16633
rect 6222 16579 6224 16631
rect 6224 16579 6276 16631
rect 6276 16579 6278 16631
rect 6222 16577 6278 16579
rect 6654 16631 6710 16633
rect 6654 16579 6656 16631
rect 6656 16579 6708 16631
rect 6708 16579 6710 16631
rect 7036 16593 7038 16645
rect 7038 16593 7090 16645
rect 7090 16593 7092 16645
rect 7036 16591 7092 16593
rect 7308 16645 7364 16647
rect 7308 16593 7310 16645
rect 7310 16593 7362 16645
rect 7362 16593 7364 16645
rect 7308 16591 7364 16593
rect 6654 16577 6710 16579
rect 5797 16273 5853 16275
rect 5797 16221 5799 16273
rect 5799 16221 5851 16273
rect 5851 16221 5853 16273
rect 5797 16219 5853 16221
rect 6222 16273 6278 16275
rect 6222 16221 6224 16273
rect 6224 16221 6276 16273
rect 6276 16221 6278 16273
rect 6222 16219 6278 16221
rect 6654 16273 6710 16275
rect 6654 16221 6656 16273
rect 6656 16221 6708 16273
rect 6708 16221 6710 16273
rect 6654 16219 6710 16221
rect 7036 16250 7092 16252
rect 7036 16198 7038 16250
rect 7038 16198 7090 16250
rect 7090 16198 7092 16250
rect 7036 16196 7092 16198
rect 7308 16250 7364 16252
rect 7308 16198 7310 16250
rect 7310 16198 7362 16250
rect 7362 16198 7364 16250
rect 7308 16196 7364 16198
rect 5797 15899 5853 15901
rect 5797 15847 5799 15899
rect 5799 15847 5851 15899
rect 5851 15847 5853 15899
rect 7036 15855 7092 15857
rect 5797 15845 5853 15847
rect 6222 15841 6278 15843
rect 6222 15789 6224 15841
rect 6224 15789 6276 15841
rect 6276 15789 6278 15841
rect 6222 15787 6278 15789
rect 6654 15841 6710 15843
rect 6654 15789 6656 15841
rect 6656 15789 6708 15841
rect 6708 15789 6710 15841
rect 7036 15803 7038 15855
rect 7038 15803 7090 15855
rect 7090 15803 7092 15855
rect 7036 15801 7092 15803
rect 7308 15855 7364 15857
rect 7308 15803 7310 15855
rect 7310 15803 7362 15855
rect 7362 15803 7364 15855
rect 7308 15801 7364 15803
rect 6654 15787 6710 15789
rect 5797 15483 5853 15485
rect 5797 15431 5799 15483
rect 5799 15431 5851 15483
rect 5851 15431 5853 15483
rect 5797 15429 5853 15431
rect 6222 15483 6278 15485
rect 6222 15431 6224 15483
rect 6224 15431 6276 15483
rect 6276 15431 6278 15483
rect 6222 15429 6278 15431
rect 6654 15483 6710 15485
rect 6654 15431 6656 15483
rect 6656 15431 6708 15483
rect 6708 15431 6710 15483
rect 6654 15429 6710 15431
rect 7036 15460 7092 15462
rect 7036 15408 7038 15460
rect 7038 15408 7090 15460
rect 7090 15408 7092 15460
rect 7036 15406 7092 15408
rect 7308 15460 7364 15462
rect 7308 15408 7310 15460
rect 7310 15408 7362 15460
rect 7362 15408 7364 15460
rect 7308 15406 7364 15408
rect 5797 15109 5853 15111
rect 5797 15057 5799 15109
rect 5799 15057 5851 15109
rect 5851 15057 5853 15109
rect 7036 15065 7092 15067
rect 5797 15055 5853 15057
rect 6222 15051 6278 15053
rect 6222 14999 6224 15051
rect 6224 14999 6276 15051
rect 6276 14999 6278 15051
rect 6222 14997 6278 14999
rect 6654 15051 6710 15053
rect 6654 14999 6656 15051
rect 6656 14999 6708 15051
rect 6708 14999 6710 15051
rect 7036 15013 7038 15065
rect 7038 15013 7090 15065
rect 7090 15013 7092 15065
rect 7036 15011 7092 15013
rect 7308 15065 7364 15067
rect 7308 15013 7310 15065
rect 7310 15013 7362 15065
rect 7362 15013 7364 15065
rect 7308 15011 7364 15013
rect 6654 14997 6710 14999
rect 5797 14693 5853 14695
rect 5797 14641 5799 14693
rect 5799 14641 5851 14693
rect 5851 14641 5853 14693
rect 5797 14639 5853 14641
rect 6222 14693 6278 14695
rect 6222 14641 6224 14693
rect 6224 14641 6276 14693
rect 6276 14641 6278 14693
rect 6222 14639 6278 14641
rect 6654 14693 6710 14695
rect 6654 14641 6656 14693
rect 6656 14641 6708 14693
rect 6708 14641 6710 14693
rect 6654 14639 6710 14641
rect 7036 14670 7092 14672
rect 7036 14618 7038 14670
rect 7038 14618 7090 14670
rect 7090 14618 7092 14670
rect 7036 14616 7092 14618
rect 7308 14670 7364 14672
rect 7308 14618 7310 14670
rect 7310 14618 7362 14670
rect 7362 14618 7364 14670
rect 7308 14616 7364 14618
rect 5797 14319 5853 14321
rect 5797 14267 5799 14319
rect 5799 14267 5851 14319
rect 5851 14267 5853 14319
rect 7036 14275 7092 14277
rect 5797 14265 5853 14267
rect 6222 14261 6278 14263
rect 6222 14209 6224 14261
rect 6224 14209 6276 14261
rect 6276 14209 6278 14261
rect 6222 14207 6278 14209
rect 6654 14261 6710 14263
rect 6654 14209 6656 14261
rect 6656 14209 6708 14261
rect 6708 14209 6710 14261
rect 7036 14223 7038 14275
rect 7038 14223 7090 14275
rect 7090 14223 7092 14275
rect 7036 14221 7092 14223
rect 7308 14275 7364 14277
rect 7308 14223 7310 14275
rect 7310 14223 7362 14275
rect 7362 14223 7364 14275
rect 7308 14221 7364 14223
rect 6654 14207 6710 14209
rect 5797 13903 5853 13905
rect 5797 13851 5799 13903
rect 5799 13851 5851 13903
rect 5851 13851 5853 13903
rect 5797 13849 5853 13851
rect 6222 13903 6278 13905
rect 6222 13851 6224 13903
rect 6224 13851 6276 13903
rect 6276 13851 6278 13903
rect 6222 13849 6278 13851
rect 6654 13903 6710 13905
rect 6654 13851 6656 13903
rect 6656 13851 6708 13903
rect 6708 13851 6710 13903
rect 6654 13849 6710 13851
rect 7036 13880 7092 13882
rect 7036 13828 7038 13880
rect 7038 13828 7090 13880
rect 7090 13828 7092 13880
rect 7036 13826 7092 13828
rect 7308 13880 7364 13882
rect 7308 13828 7310 13880
rect 7310 13828 7362 13880
rect 7362 13828 7364 13880
rect 7308 13826 7364 13828
rect 5797 13529 5853 13531
rect 5797 13477 5799 13529
rect 5799 13477 5851 13529
rect 5851 13477 5853 13529
rect 7036 13485 7092 13487
rect 5797 13475 5853 13477
rect 6222 13471 6278 13473
rect 6222 13419 6224 13471
rect 6224 13419 6276 13471
rect 6276 13419 6278 13471
rect 6222 13417 6278 13419
rect 6654 13471 6710 13473
rect 6654 13419 6656 13471
rect 6656 13419 6708 13471
rect 6708 13419 6710 13471
rect 7036 13433 7038 13485
rect 7038 13433 7090 13485
rect 7090 13433 7092 13485
rect 7036 13431 7092 13433
rect 7308 13485 7364 13487
rect 7308 13433 7310 13485
rect 7310 13433 7362 13485
rect 7362 13433 7364 13485
rect 7308 13431 7364 13433
rect 6654 13417 6710 13419
rect 5797 13113 5853 13115
rect 5797 13061 5799 13113
rect 5799 13061 5851 13113
rect 5851 13061 5853 13113
rect 5797 13059 5853 13061
rect 6222 13113 6278 13115
rect 6222 13061 6224 13113
rect 6224 13061 6276 13113
rect 6276 13061 6278 13113
rect 6222 13059 6278 13061
rect 6654 13113 6710 13115
rect 6654 13061 6656 13113
rect 6656 13061 6708 13113
rect 6708 13061 6710 13113
rect 6654 13059 6710 13061
rect 7036 13090 7092 13092
rect 7036 13038 7038 13090
rect 7038 13038 7090 13090
rect 7090 13038 7092 13090
rect 7036 13036 7092 13038
rect 7308 13090 7364 13092
rect 7308 13038 7310 13090
rect 7310 13038 7362 13090
rect 7362 13038 7364 13090
rect 7308 13036 7364 13038
rect 5797 12739 5853 12741
rect 5797 12687 5799 12739
rect 5799 12687 5851 12739
rect 5851 12687 5853 12739
rect 7036 12695 7092 12697
rect 5797 12685 5853 12687
rect 6222 12681 6278 12683
rect 6222 12629 6224 12681
rect 6224 12629 6276 12681
rect 6276 12629 6278 12681
rect 6222 12627 6278 12629
rect 6654 12681 6710 12683
rect 6654 12629 6656 12681
rect 6656 12629 6708 12681
rect 6708 12629 6710 12681
rect 7036 12643 7038 12695
rect 7038 12643 7090 12695
rect 7090 12643 7092 12695
rect 7036 12641 7092 12643
rect 7308 12695 7364 12697
rect 7308 12643 7310 12695
rect 7310 12643 7362 12695
rect 7362 12643 7364 12695
rect 7308 12641 7364 12643
rect 6654 12627 6710 12629
rect 5797 12323 5853 12325
rect 5797 12271 5799 12323
rect 5799 12271 5851 12323
rect 5851 12271 5853 12323
rect 5797 12269 5853 12271
rect 6222 12323 6278 12325
rect 6222 12271 6224 12323
rect 6224 12271 6276 12323
rect 6276 12271 6278 12323
rect 6222 12269 6278 12271
rect 6654 12323 6710 12325
rect 6654 12271 6656 12323
rect 6656 12271 6708 12323
rect 6708 12271 6710 12323
rect 6654 12269 6710 12271
rect 7036 12300 7092 12302
rect 7036 12248 7038 12300
rect 7038 12248 7090 12300
rect 7090 12248 7092 12300
rect 7036 12246 7092 12248
rect 7308 12300 7364 12302
rect 7308 12248 7310 12300
rect 7310 12248 7362 12300
rect 7362 12248 7364 12300
rect 7308 12246 7364 12248
rect 5797 11949 5853 11951
rect 5797 11897 5799 11949
rect 5799 11897 5851 11949
rect 5851 11897 5853 11949
rect 7036 11905 7092 11907
rect 5797 11895 5853 11897
rect 6222 11891 6278 11893
rect 6222 11839 6224 11891
rect 6224 11839 6276 11891
rect 6276 11839 6278 11891
rect 6222 11837 6278 11839
rect 6654 11891 6710 11893
rect 6654 11839 6656 11891
rect 6656 11839 6708 11891
rect 6708 11839 6710 11891
rect 7036 11853 7038 11905
rect 7038 11853 7090 11905
rect 7090 11853 7092 11905
rect 7036 11851 7092 11853
rect 7308 11905 7364 11907
rect 7308 11853 7310 11905
rect 7310 11853 7362 11905
rect 7362 11853 7364 11905
rect 7308 11851 7364 11853
rect 6654 11837 6710 11839
rect 5797 11533 5853 11535
rect 5797 11481 5799 11533
rect 5799 11481 5851 11533
rect 5851 11481 5853 11533
rect 5797 11479 5853 11481
rect 6222 11533 6278 11535
rect 6222 11481 6224 11533
rect 6224 11481 6276 11533
rect 6276 11481 6278 11533
rect 6222 11479 6278 11481
rect 6654 11533 6710 11535
rect 6654 11481 6656 11533
rect 6656 11481 6708 11533
rect 6708 11481 6710 11533
rect 6654 11479 6710 11481
rect 7036 11510 7092 11512
rect 7036 11458 7038 11510
rect 7038 11458 7090 11510
rect 7090 11458 7092 11510
rect 7036 11456 7092 11458
rect 7308 11510 7364 11512
rect 7308 11458 7310 11510
rect 7310 11458 7362 11510
rect 7362 11458 7364 11510
rect 7308 11456 7364 11458
rect 5797 11159 5853 11161
rect 5797 11107 5799 11159
rect 5799 11107 5851 11159
rect 5851 11107 5853 11159
rect 7036 11115 7092 11117
rect 5797 11105 5853 11107
rect 6222 11101 6278 11103
rect 6222 11049 6224 11101
rect 6224 11049 6276 11101
rect 6276 11049 6278 11101
rect 6222 11047 6278 11049
rect 6654 11101 6710 11103
rect 6654 11049 6656 11101
rect 6656 11049 6708 11101
rect 6708 11049 6710 11101
rect 7036 11063 7038 11115
rect 7038 11063 7090 11115
rect 7090 11063 7092 11115
rect 7036 11061 7092 11063
rect 7308 11115 7364 11117
rect 7308 11063 7310 11115
rect 7310 11063 7362 11115
rect 7362 11063 7364 11115
rect 7308 11061 7364 11063
rect 6654 11047 6710 11049
rect 5797 10743 5853 10745
rect 5797 10691 5799 10743
rect 5799 10691 5851 10743
rect 5851 10691 5853 10743
rect 5797 10689 5853 10691
rect 6222 10743 6278 10745
rect 6222 10691 6224 10743
rect 6224 10691 6276 10743
rect 6276 10691 6278 10743
rect 6222 10689 6278 10691
rect 6654 10743 6710 10745
rect 6654 10691 6656 10743
rect 6656 10691 6708 10743
rect 6708 10691 6710 10743
rect 6654 10689 6710 10691
rect 7036 10720 7092 10722
rect 7036 10668 7038 10720
rect 7038 10668 7090 10720
rect 7090 10668 7092 10720
rect 7036 10666 7092 10668
rect 7308 10720 7364 10722
rect 7308 10668 7310 10720
rect 7310 10668 7362 10720
rect 7362 10668 7364 10720
rect 7308 10666 7364 10668
rect 5797 10369 5853 10371
rect 5797 10317 5799 10369
rect 5799 10317 5851 10369
rect 5851 10317 5853 10369
rect 7036 10325 7092 10327
rect 5797 10315 5853 10317
rect 6222 10311 6278 10313
rect 6222 10259 6224 10311
rect 6224 10259 6276 10311
rect 6276 10259 6278 10311
rect 6222 10257 6278 10259
rect 6654 10311 6710 10313
rect 6654 10259 6656 10311
rect 6656 10259 6708 10311
rect 6708 10259 6710 10311
rect 7036 10273 7038 10325
rect 7038 10273 7090 10325
rect 7090 10273 7092 10325
rect 7036 10271 7092 10273
rect 7308 10325 7364 10327
rect 7308 10273 7310 10325
rect 7310 10273 7362 10325
rect 7362 10273 7364 10325
rect 7308 10271 7364 10273
rect 6654 10257 6710 10259
rect 5797 9953 5853 9955
rect 5797 9901 5799 9953
rect 5799 9901 5851 9953
rect 5851 9901 5853 9953
rect 5797 9899 5853 9901
rect 6222 9953 6278 9955
rect 6222 9901 6224 9953
rect 6224 9901 6276 9953
rect 6276 9901 6278 9953
rect 6222 9899 6278 9901
rect 6654 9953 6710 9955
rect 6654 9901 6656 9953
rect 6656 9901 6708 9953
rect 6708 9901 6710 9953
rect 6654 9899 6710 9901
rect 7036 9930 7092 9932
rect 7036 9878 7038 9930
rect 7038 9878 7090 9930
rect 7090 9878 7092 9930
rect 7036 9876 7092 9878
rect 7308 9930 7364 9932
rect 7308 9878 7310 9930
rect 7310 9878 7362 9930
rect 7362 9878 7364 9930
rect 7308 9876 7364 9878
rect 5797 9579 5853 9581
rect 5797 9527 5799 9579
rect 5799 9527 5851 9579
rect 5851 9527 5853 9579
rect 7036 9535 7092 9537
rect 5797 9525 5853 9527
rect 6222 9521 6278 9523
rect 6222 9469 6224 9521
rect 6224 9469 6276 9521
rect 6276 9469 6278 9521
rect 6222 9467 6278 9469
rect 6654 9521 6710 9523
rect 6654 9469 6656 9521
rect 6656 9469 6708 9521
rect 6708 9469 6710 9521
rect 7036 9483 7038 9535
rect 7038 9483 7090 9535
rect 7090 9483 7092 9535
rect 7036 9481 7092 9483
rect 7308 9535 7364 9537
rect 7308 9483 7310 9535
rect 7310 9483 7362 9535
rect 7362 9483 7364 9535
rect 7308 9481 7364 9483
rect 6654 9467 6710 9469
rect 5797 9163 5853 9165
rect 5797 9111 5799 9163
rect 5799 9111 5851 9163
rect 5851 9111 5853 9163
rect 5797 9109 5853 9111
rect 6222 9163 6278 9165
rect 6222 9111 6224 9163
rect 6224 9111 6276 9163
rect 6276 9111 6278 9163
rect 6222 9109 6278 9111
rect 6654 9163 6710 9165
rect 6654 9111 6656 9163
rect 6656 9111 6708 9163
rect 6708 9111 6710 9163
rect 6654 9109 6710 9111
rect 7036 9140 7092 9142
rect 7036 9088 7038 9140
rect 7038 9088 7090 9140
rect 7090 9088 7092 9140
rect 7036 9086 7092 9088
rect 7308 9140 7364 9142
rect 7308 9088 7310 9140
rect 7310 9088 7362 9140
rect 7362 9088 7364 9140
rect 7308 9086 7364 9088
rect 5797 8789 5853 8791
rect 5797 8737 5799 8789
rect 5799 8737 5851 8789
rect 5851 8737 5853 8789
rect 7036 8745 7092 8747
rect 5797 8735 5853 8737
rect 6222 8731 6278 8733
rect 6222 8679 6224 8731
rect 6224 8679 6276 8731
rect 6276 8679 6278 8731
rect 6222 8677 6278 8679
rect 6654 8731 6710 8733
rect 6654 8679 6656 8731
rect 6656 8679 6708 8731
rect 6708 8679 6710 8731
rect 7036 8693 7038 8745
rect 7038 8693 7090 8745
rect 7090 8693 7092 8745
rect 7036 8691 7092 8693
rect 7308 8745 7364 8747
rect 7308 8693 7310 8745
rect 7310 8693 7362 8745
rect 7362 8693 7364 8745
rect 7308 8691 7364 8693
rect 6654 8677 6710 8679
rect 5797 8373 5853 8375
rect 5797 8321 5799 8373
rect 5799 8321 5851 8373
rect 5851 8321 5853 8373
rect 5797 8319 5853 8321
rect 6222 8373 6278 8375
rect 6222 8321 6224 8373
rect 6224 8321 6276 8373
rect 6276 8321 6278 8373
rect 6222 8319 6278 8321
rect 6654 8373 6710 8375
rect 6654 8321 6656 8373
rect 6656 8321 6708 8373
rect 6708 8321 6710 8373
rect 6654 8319 6710 8321
rect 7036 8350 7092 8352
rect 7036 8298 7038 8350
rect 7038 8298 7090 8350
rect 7090 8298 7092 8350
rect 7036 8296 7092 8298
rect 7308 8350 7364 8352
rect 7308 8298 7310 8350
rect 7310 8298 7362 8350
rect 7362 8298 7364 8350
rect 7308 8296 7364 8298
rect 5797 7999 5853 8001
rect 5797 7947 5799 7999
rect 5799 7947 5851 7999
rect 5851 7947 5853 7999
rect 7036 7955 7092 7957
rect 5797 7945 5853 7947
rect 6222 7941 6278 7943
rect 6222 7889 6224 7941
rect 6224 7889 6276 7941
rect 6276 7889 6278 7941
rect 6222 7887 6278 7889
rect 6654 7941 6710 7943
rect 6654 7889 6656 7941
rect 6656 7889 6708 7941
rect 6708 7889 6710 7941
rect 7036 7903 7038 7955
rect 7038 7903 7090 7955
rect 7090 7903 7092 7955
rect 7036 7901 7092 7903
rect 7308 7955 7364 7957
rect 7308 7903 7310 7955
rect 7310 7903 7362 7955
rect 7362 7903 7364 7955
rect 7308 7901 7364 7903
rect 6654 7887 6710 7889
rect 5797 7583 5853 7585
rect 5797 7531 5799 7583
rect 5799 7531 5851 7583
rect 5851 7531 5853 7583
rect 5797 7529 5853 7531
rect 6222 7583 6278 7585
rect 6222 7531 6224 7583
rect 6224 7531 6276 7583
rect 6276 7531 6278 7583
rect 6222 7529 6278 7531
rect 6654 7583 6710 7585
rect 6654 7531 6656 7583
rect 6656 7531 6708 7583
rect 6708 7531 6710 7583
rect 6654 7529 6710 7531
rect 7036 7560 7092 7562
rect 7036 7508 7038 7560
rect 7038 7508 7090 7560
rect 7090 7508 7092 7560
rect 7036 7506 7092 7508
rect 7308 7560 7364 7562
rect 7308 7508 7310 7560
rect 7310 7508 7362 7560
rect 7362 7508 7364 7560
rect 7308 7506 7364 7508
rect 5797 7209 5853 7211
rect 5797 7157 5799 7209
rect 5799 7157 5851 7209
rect 5851 7157 5853 7209
rect 7036 7165 7092 7167
rect 5797 7155 5853 7157
rect 6222 7151 6278 7153
rect 6222 7099 6224 7151
rect 6224 7099 6276 7151
rect 6276 7099 6278 7151
rect 6222 7097 6278 7099
rect 6654 7151 6710 7153
rect 6654 7099 6656 7151
rect 6656 7099 6708 7151
rect 6708 7099 6710 7151
rect 7036 7113 7038 7165
rect 7038 7113 7090 7165
rect 7090 7113 7092 7165
rect 7036 7111 7092 7113
rect 7308 7165 7364 7167
rect 7308 7113 7310 7165
rect 7310 7113 7362 7165
rect 7362 7113 7364 7165
rect 7308 7111 7364 7113
rect 6654 7097 6710 7099
rect 5797 6793 5853 6795
rect 5797 6741 5799 6793
rect 5799 6741 5851 6793
rect 5851 6741 5853 6793
rect 5797 6739 5853 6741
rect 6222 6793 6278 6795
rect 6222 6741 6224 6793
rect 6224 6741 6276 6793
rect 6276 6741 6278 6793
rect 6222 6739 6278 6741
rect 6654 6793 6710 6795
rect 6654 6741 6656 6793
rect 6656 6741 6708 6793
rect 6708 6741 6710 6793
rect 6654 6739 6710 6741
rect 7036 6770 7092 6772
rect 7036 6718 7038 6770
rect 7038 6718 7090 6770
rect 7090 6718 7092 6770
rect 7036 6716 7092 6718
rect 7308 6770 7364 6772
rect 7308 6718 7310 6770
rect 7310 6718 7362 6770
rect 7362 6718 7364 6770
rect 7308 6716 7364 6718
rect 5797 6419 5853 6421
rect 5797 6367 5799 6419
rect 5799 6367 5851 6419
rect 5851 6367 5853 6419
rect 7036 6375 7092 6377
rect 5797 6365 5853 6367
rect 6222 6361 6278 6363
rect 6222 6309 6224 6361
rect 6224 6309 6276 6361
rect 6276 6309 6278 6361
rect 6222 6307 6278 6309
rect 6654 6361 6710 6363
rect 6654 6309 6656 6361
rect 6656 6309 6708 6361
rect 6708 6309 6710 6361
rect 7036 6323 7038 6375
rect 7038 6323 7090 6375
rect 7090 6323 7092 6375
rect 7036 6321 7092 6323
rect 7308 6375 7364 6377
rect 7308 6323 7310 6375
rect 7310 6323 7362 6375
rect 7362 6323 7364 6375
rect 7308 6321 7364 6323
rect 6654 6307 6710 6309
rect 5797 6003 5853 6005
rect 5797 5951 5799 6003
rect 5799 5951 5851 6003
rect 5851 5951 5853 6003
rect 5797 5949 5853 5951
rect 6222 6003 6278 6005
rect 6222 5951 6224 6003
rect 6224 5951 6276 6003
rect 6276 5951 6278 6003
rect 6222 5949 6278 5951
rect 6654 6003 6710 6005
rect 6654 5951 6656 6003
rect 6656 5951 6708 6003
rect 6708 5951 6710 6003
rect 6654 5949 6710 5951
rect 7036 5980 7092 5982
rect 7036 5928 7038 5980
rect 7038 5928 7090 5980
rect 7090 5928 7092 5980
rect 7036 5926 7092 5928
rect 7308 5980 7364 5982
rect 7308 5928 7310 5980
rect 7310 5928 7362 5980
rect 7362 5928 7364 5980
rect 7308 5926 7364 5928
rect 5797 5629 5853 5631
rect 5797 5577 5799 5629
rect 5799 5577 5851 5629
rect 5851 5577 5853 5629
rect 7036 5585 7092 5587
rect 5797 5575 5853 5577
rect 6222 5571 6278 5573
rect 6222 5519 6224 5571
rect 6224 5519 6276 5571
rect 6276 5519 6278 5571
rect 6222 5517 6278 5519
rect 6654 5571 6710 5573
rect 6654 5519 6656 5571
rect 6656 5519 6708 5571
rect 6708 5519 6710 5571
rect 7036 5533 7038 5585
rect 7038 5533 7090 5585
rect 7090 5533 7092 5585
rect 7036 5531 7092 5533
rect 7308 5585 7364 5587
rect 7308 5533 7310 5585
rect 7310 5533 7362 5585
rect 7362 5533 7364 5585
rect 7308 5531 7364 5533
rect 6654 5517 6710 5519
rect 5797 5213 5853 5215
rect 5797 5161 5799 5213
rect 5799 5161 5851 5213
rect 5851 5161 5853 5213
rect 5797 5159 5853 5161
rect 6222 5213 6278 5215
rect 6222 5161 6224 5213
rect 6224 5161 6276 5213
rect 6276 5161 6278 5213
rect 6222 5159 6278 5161
rect 6654 5213 6710 5215
rect 6654 5161 6656 5213
rect 6656 5161 6708 5213
rect 6708 5161 6710 5213
rect 6654 5159 6710 5161
rect 7036 5190 7092 5192
rect 7036 5138 7038 5190
rect 7038 5138 7090 5190
rect 7090 5138 7092 5190
rect 7036 5136 7092 5138
rect 7308 5190 7364 5192
rect 7308 5138 7310 5190
rect 7310 5138 7362 5190
rect 7362 5138 7364 5190
rect 7308 5136 7364 5138
rect 5797 4839 5853 4841
rect 5797 4787 5799 4839
rect 5799 4787 5851 4839
rect 5851 4787 5853 4839
rect 7036 4795 7092 4797
rect 5797 4785 5853 4787
rect 6222 4781 6278 4783
rect 6222 4729 6224 4781
rect 6224 4729 6276 4781
rect 6276 4729 6278 4781
rect 6222 4727 6278 4729
rect 6654 4781 6710 4783
rect 6654 4729 6656 4781
rect 6656 4729 6708 4781
rect 6708 4729 6710 4781
rect 7036 4743 7038 4795
rect 7038 4743 7090 4795
rect 7090 4743 7092 4795
rect 7036 4741 7092 4743
rect 7308 4795 7364 4797
rect 7308 4743 7310 4795
rect 7310 4743 7362 4795
rect 7362 4743 7364 4795
rect 7308 4741 7364 4743
rect 6654 4727 6710 4729
rect 5797 4423 5853 4425
rect 5797 4371 5799 4423
rect 5799 4371 5851 4423
rect 5851 4371 5853 4423
rect 5797 4369 5853 4371
rect 6222 4423 6278 4425
rect 6222 4371 6224 4423
rect 6224 4371 6276 4423
rect 6276 4371 6278 4423
rect 6222 4369 6278 4371
rect 6654 4423 6710 4425
rect 6654 4371 6656 4423
rect 6656 4371 6708 4423
rect 6708 4371 6710 4423
rect 6654 4369 6710 4371
rect 7036 4400 7092 4402
rect 7036 4348 7038 4400
rect 7038 4348 7090 4400
rect 7090 4348 7092 4400
rect 7036 4346 7092 4348
rect 7308 4400 7364 4402
rect 7308 4348 7310 4400
rect 7310 4348 7362 4400
rect 7362 4348 7364 4400
rect 7308 4346 7364 4348
rect 5797 4049 5853 4051
rect 5797 3997 5799 4049
rect 5799 3997 5851 4049
rect 5851 3997 5853 4049
rect 7036 4005 7092 4007
rect 5797 3995 5853 3997
rect 6222 3991 6278 3993
rect 6222 3939 6224 3991
rect 6224 3939 6276 3991
rect 6276 3939 6278 3991
rect 6222 3937 6278 3939
rect 6654 3991 6710 3993
rect 6654 3939 6656 3991
rect 6656 3939 6708 3991
rect 6708 3939 6710 3991
rect 7036 3953 7038 4005
rect 7038 3953 7090 4005
rect 7090 3953 7092 4005
rect 7036 3951 7092 3953
rect 7308 4005 7364 4007
rect 7308 3953 7310 4005
rect 7310 3953 7362 4005
rect 7362 3953 7364 4005
rect 7308 3951 7364 3953
rect 6654 3937 6710 3939
rect 5797 3633 5853 3635
rect 5797 3581 5799 3633
rect 5799 3581 5851 3633
rect 5851 3581 5853 3633
rect 5797 3579 5853 3581
rect 6222 3633 6278 3635
rect 6222 3581 6224 3633
rect 6224 3581 6276 3633
rect 6276 3581 6278 3633
rect 6222 3579 6278 3581
rect 6654 3633 6710 3635
rect 6654 3581 6656 3633
rect 6656 3581 6708 3633
rect 6708 3581 6710 3633
rect 6654 3579 6710 3581
rect 7036 3610 7092 3612
rect 7036 3558 7038 3610
rect 7038 3558 7090 3610
rect 7090 3558 7092 3610
rect 7036 3556 7092 3558
rect 7308 3610 7364 3612
rect 7308 3558 7310 3610
rect 7310 3558 7362 3610
rect 7362 3558 7364 3610
rect 7308 3556 7364 3558
rect 5797 3259 5853 3261
rect 5797 3207 5799 3259
rect 5799 3207 5851 3259
rect 5851 3207 5853 3259
rect 7036 3215 7092 3217
rect 5797 3205 5853 3207
rect 6222 3201 6278 3203
rect 6222 3149 6224 3201
rect 6224 3149 6276 3201
rect 6276 3149 6278 3201
rect 6222 3147 6278 3149
rect 6654 3201 6710 3203
rect 6654 3149 6656 3201
rect 6656 3149 6708 3201
rect 6708 3149 6710 3201
rect 7036 3163 7038 3215
rect 7038 3163 7090 3215
rect 7090 3163 7092 3215
rect 7036 3161 7092 3163
rect 7308 3215 7364 3217
rect 7308 3163 7310 3215
rect 7310 3163 7362 3215
rect 7362 3163 7364 3215
rect 7308 3161 7364 3163
rect 6654 3147 6710 3149
rect 5797 2843 5853 2845
rect 5797 2791 5799 2843
rect 5799 2791 5851 2843
rect 5851 2791 5853 2843
rect 5797 2789 5853 2791
rect 6222 2843 6278 2845
rect 6222 2791 6224 2843
rect 6224 2791 6276 2843
rect 6276 2791 6278 2843
rect 6222 2789 6278 2791
rect 6654 2843 6710 2845
rect 6654 2791 6656 2843
rect 6656 2791 6708 2843
rect 6708 2791 6710 2843
rect 6654 2789 6710 2791
rect 7036 2820 7092 2822
rect 7036 2768 7038 2820
rect 7038 2768 7090 2820
rect 7090 2768 7092 2820
rect 7036 2766 7092 2768
rect 7308 2820 7364 2822
rect 7308 2768 7310 2820
rect 7310 2768 7362 2820
rect 7362 2768 7364 2820
rect 7308 2766 7364 2768
rect 5797 2469 5853 2471
rect 5797 2417 5799 2469
rect 5799 2417 5851 2469
rect 5851 2417 5853 2469
rect 7036 2425 7092 2427
rect 5797 2415 5853 2417
rect 6222 2411 6278 2413
rect 6222 2359 6224 2411
rect 6224 2359 6276 2411
rect 6276 2359 6278 2411
rect 6222 2357 6278 2359
rect 6654 2411 6710 2413
rect 6654 2359 6656 2411
rect 6656 2359 6708 2411
rect 6708 2359 6710 2411
rect 7036 2373 7038 2425
rect 7038 2373 7090 2425
rect 7090 2373 7092 2425
rect 7036 2371 7092 2373
rect 7308 2425 7364 2427
rect 7308 2373 7310 2425
rect 7310 2373 7362 2425
rect 7362 2373 7364 2425
rect 7308 2371 7364 2373
rect 6654 2357 6710 2359
rect 5797 2053 5853 2055
rect 5797 2001 5799 2053
rect 5799 2001 5851 2053
rect 5851 2001 5853 2053
rect 5797 1999 5853 2001
rect 6222 2053 6278 2055
rect 6222 2001 6224 2053
rect 6224 2001 6276 2053
rect 6276 2001 6278 2053
rect 6222 1999 6278 2001
rect 6654 2053 6710 2055
rect 6654 2001 6656 2053
rect 6656 2001 6708 2053
rect 6708 2001 6710 2053
rect 6654 1999 6710 2001
rect 7036 2030 7092 2032
rect 7036 1978 7038 2030
rect 7038 1978 7090 2030
rect 7090 1978 7092 2030
rect 7036 1976 7092 1978
rect 7308 2030 7364 2032
rect 7308 1978 7310 2030
rect 7310 1978 7362 2030
rect 7362 1978 7364 2030
rect 7308 1976 7364 1978
rect 5797 1679 5853 1681
rect 5797 1627 5799 1679
rect 5799 1627 5851 1679
rect 5851 1627 5853 1679
rect 7036 1635 7092 1637
rect 5797 1625 5853 1627
rect 6222 1621 6278 1623
rect 6222 1569 6224 1621
rect 6224 1569 6276 1621
rect 6276 1569 6278 1621
rect 6222 1567 6278 1569
rect 6654 1621 6710 1623
rect 6654 1569 6656 1621
rect 6656 1569 6708 1621
rect 6708 1569 6710 1621
rect 7036 1583 7038 1635
rect 7038 1583 7090 1635
rect 7090 1583 7092 1635
rect 7036 1581 7092 1583
rect 7308 1635 7364 1637
rect 7308 1583 7310 1635
rect 7310 1583 7362 1635
rect 7362 1583 7364 1635
rect 7308 1581 7364 1583
rect 6654 1567 6710 1569
rect 5797 1263 5853 1265
rect 5797 1211 5799 1263
rect 5799 1211 5851 1263
rect 5851 1211 5853 1263
rect 5797 1209 5853 1211
rect 6222 1263 6278 1265
rect 6222 1211 6224 1263
rect 6224 1211 6276 1263
rect 6276 1211 6278 1263
rect 6222 1209 6278 1211
rect 6654 1263 6710 1265
rect 6654 1211 6656 1263
rect 6656 1211 6708 1263
rect 6708 1211 6710 1263
rect 6654 1209 6710 1211
rect 7036 1240 7092 1242
rect 7036 1188 7038 1240
rect 7038 1188 7090 1240
rect 7090 1188 7092 1240
rect 7036 1186 7092 1188
rect 7308 1240 7364 1242
rect 7308 1188 7310 1240
rect 7310 1188 7362 1240
rect 7362 1188 7364 1240
rect 7308 1186 7364 1188
rect 5797 889 5853 891
rect 5797 837 5799 889
rect 5799 837 5851 889
rect 5851 837 5853 889
rect 7036 845 7092 847
rect 5797 835 5853 837
rect 6222 831 6278 833
rect 6222 779 6224 831
rect 6224 779 6276 831
rect 6276 779 6278 831
rect 6222 777 6278 779
rect 6654 831 6710 833
rect 6654 779 6656 831
rect 6656 779 6708 831
rect 6708 779 6710 831
rect 7036 793 7038 845
rect 7038 793 7090 845
rect 7090 793 7092 845
rect 7036 791 7092 793
rect 7308 845 7364 847
rect 7308 793 7310 845
rect 7310 793 7362 845
rect 7362 793 7364 845
rect 7308 791 7364 793
rect 6654 777 6710 779
rect 5797 473 5853 475
rect 5797 421 5799 473
rect 5799 421 5851 473
rect 5851 421 5853 473
rect 5797 419 5853 421
rect 6222 473 6278 475
rect 6222 421 6224 473
rect 6224 421 6276 473
rect 6276 421 6278 473
rect 6222 419 6278 421
rect 6654 473 6710 475
rect 6654 421 6656 473
rect 6656 421 6708 473
rect 6708 421 6710 473
rect 6654 419 6710 421
rect 7036 450 7092 452
rect 7036 398 7038 450
rect 7038 398 7090 450
rect 7090 398 7092 450
rect 7036 396 7092 398
rect 7308 450 7364 452
rect 7308 398 7310 450
rect 7310 398 7362 450
rect 7362 398 7364 450
rect 7308 396 7364 398
<< metal3 >>
rect 5776 50245 5874 50266
rect 5776 50189 5797 50245
rect 5853 50189 5874 50245
rect 5776 50168 5874 50189
rect 6201 50245 6299 50266
rect 6201 50189 6222 50245
rect 6278 50189 6299 50245
rect 6201 50168 6299 50189
rect 6633 50245 6731 50266
rect 6633 50189 6654 50245
rect 6710 50189 6731 50245
rect 6633 50168 6731 50189
rect 7015 50222 7113 50243
rect 7015 50166 7036 50222
rect 7092 50166 7113 50222
rect 7015 50145 7113 50166
rect 7287 50222 7385 50243
rect 7287 50166 7308 50222
rect 7364 50166 7385 50222
rect 7287 50145 7385 50166
rect 5776 49871 5874 49892
rect 5776 49815 5797 49871
rect 5853 49815 5874 49871
rect 5776 49794 5874 49815
rect 6201 49813 6299 49834
rect 6201 49757 6222 49813
rect 6278 49757 6299 49813
rect 6201 49736 6299 49757
rect 6633 49813 6731 49834
rect 6633 49757 6654 49813
rect 6710 49757 6731 49813
rect 6633 49736 6731 49757
rect 7015 49827 7113 49848
rect 7015 49771 7036 49827
rect 7092 49771 7113 49827
rect 7015 49750 7113 49771
rect 7287 49827 7385 49848
rect 7287 49771 7308 49827
rect 7364 49771 7385 49827
rect 7287 49750 7385 49771
rect 5776 49455 5874 49476
rect 5776 49399 5797 49455
rect 5853 49399 5874 49455
rect 5776 49378 5874 49399
rect 6201 49455 6299 49476
rect 6201 49399 6222 49455
rect 6278 49399 6299 49455
rect 6201 49378 6299 49399
rect 6633 49455 6731 49476
rect 6633 49399 6654 49455
rect 6710 49399 6731 49455
rect 6633 49378 6731 49399
rect 7015 49432 7113 49453
rect 7015 49376 7036 49432
rect 7092 49376 7113 49432
rect 7015 49355 7113 49376
rect 7287 49432 7382 49453
rect 7287 49376 7308 49432
rect 7364 49376 7382 49432
rect 7287 49355 7382 49376
rect 5776 49081 5874 49102
rect 5776 49025 5797 49081
rect 5853 49025 5874 49081
rect 5776 49004 5874 49025
rect 6201 49023 6299 49044
rect 6201 48967 6222 49023
rect 6278 48967 6299 49023
rect 6201 48946 6299 48967
rect 6633 49023 6731 49044
rect 6633 48967 6654 49023
rect 6710 48967 6731 49023
rect 6633 48946 6731 48967
rect 7015 49037 7113 49058
rect 7015 48981 7036 49037
rect 7092 48981 7113 49037
rect 7015 48960 7113 48981
rect 7287 49037 7385 49058
rect 7287 48981 7308 49037
rect 7364 48981 7385 49037
rect 7287 48960 7385 48981
rect 5776 48665 5874 48686
rect 5776 48609 5797 48665
rect 5853 48609 5874 48665
rect 5776 48588 5874 48609
rect 6201 48665 6299 48686
rect 6201 48609 6222 48665
rect 6278 48609 6299 48665
rect 6201 48588 6299 48609
rect 6633 48665 6731 48686
rect 6633 48609 6654 48665
rect 6710 48609 6731 48665
rect 6633 48588 6731 48609
rect 7015 48642 7113 48663
rect 7015 48586 7036 48642
rect 7092 48586 7113 48642
rect 7015 48565 7113 48586
rect 7287 48642 7385 48663
rect 7287 48586 7308 48642
rect 7364 48586 7385 48642
rect 7287 48565 7385 48586
rect 5776 48291 5874 48312
rect 5776 48235 5797 48291
rect 5853 48235 5874 48291
rect 5776 48214 5874 48235
rect 6201 48233 6299 48254
rect 6201 48177 6222 48233
rect 6278 48177 6299 48233
rect 6201 48156 6299 48177
rect 6633 48233 6731 48254
rect 6633 48177 6654 48233
rect 6710 48177 6731 48233
rect 6633 48156 6731 48177
rect 7015 48247 7113 48268
rect 7015 48191 7036 48247
rect 7092 48191 7113 48247
rect 7015 48170 7113 48191
rect 7287 48247 7385 48268
rect 7287 48191 7308 48247
rect 7364 48191 7385 48247
rect 7287 48170 7385 48191
rect 5776 47875 5874 47896
rect 5776 47819 5797 47875
rect 5853 47819 5874 47875
rect 5776 47798 5874 47819
rect 6201 47875 6299 47896
rect 6201 47819 6222 47875
rect 6278 47819 6299 47875
rect 6201 47798 6299 47819
rect 6633 47875 6731 47896
rect 6633 47819 6654 47875
rect 6710 47819 6731 47875
rect 6633 47798 6731 47819
rect 7015 47852 7113 47873
rect 7015 47796 7036 47852
rect 7092 47796 7113 47852
rect 7015 47775 7113 47796
rect 7287 47852 7385 47873
rect 7287 47796 7308 47852
rect 7364 47796 7385 47852
rect 7287 47775 7385 47796
rect 5776 47501 5874 47522
rect 5776 47445 5797 47501
rect 5853 47445 5874 47501
rect 5776 47424 5874 47445
rect 6201 47443 6299 47464
rect 6201 47387 6222 47443
rect 6278 47387 6299 47443
rect 6201 47366 6299 47387
rect 6633 47443 6731 47464
rect 6633 47387 6654 47443
rect 6710 47387 6731 47443
rect 6633 47366 6731 47387
rect 7015 47457 7113 47478
rect 7015 47401 7036 47457
rect 7092 47401 7113 47457
rect 7015 47380 7113 47401
rect 7287 47457 7385 47478
rect 7287 47401 7308 47457
rect 7364 47401 7385 47457
rect 7287 47380 7385 47401
rect 5776 47085 5874 47106
rect 5776 47029 5797 47085
rect 5853 47029 5874 47085
rect 5776 47008 5874 47029
rect 6201 47085 6299 47106
rect 6201 47029 6222 47085
rect 6278 47029 6299 47085
rect 6201 47008 6299 47029
rect 6633 47085 6731 47106
rect 6633 47029 6654 47085
rect 6710 47029 6731 47085
rect 6633 47008 6731 47029
rect 7015 47062 7113 47083
rect 7015 47006 7036 47062
rect 7092 47006 7113 47062
rect 7015 46985 7113 47006
rect 7287 47062 7385 47083
rect 7287 47006 7308 47062
rect 7364 47006 7385 47062
rect 7287 46985 7385 47006
rect 5776 46711 5874 46732
rect 5776 46655 5797 46711
rect 5853 46655 5874 46711
rect 5776 46634 5874 46655
rect 6201 46653 6299 46674
rect 6201 46597 6222 46653
rect 6278 46597 6299 46653
rect 6201 46576 6299 46597
rect 6633 46653 6731 46674
rect 6633 46597 6654 46653
rect 6710 46597 6731 46653
rect 6633 46576 6731 46597
rect 7015 46667 7113 46688
rect 7015 46611 7036 46667
rect 7092 46611 7113 46667
rect 7015 46590 7113 46611
rect 7287 46667 7385 46688
rect 7287 46611 7308 46667
rect 7364 46611 7385 46667
rect 7287 46590 7385 46611
rect 5776 46295 5874 46316
rect 5776 46239 5797 46295
rect 5853 46239 5874 46295
rect 5776 46218 5874 46239
rect 6201 46295 6299 46316
rect 6201 46239 6222 46295
rect 6278 46239 6299 46295
rect 6201 46218 6299 46239
rect 6633 46295 6731 46316
rect 6633 46239 6654 46295
rect 6710 46239 6731 46295
rect 6633 46218 6731 46239
rect 7015 46272 7113 46293
rect 7015 46216 7036 46272
rect 7092 46216 7113 46272
rect 7015 46195 7113 46216
rect 7287 46272 7385 46293
rect 7287 46216 7308 46272
rect 7364 46216 7385 46272
rect 7287 46195 7385 46216
rect 5776 45921 5874 45942
rect 5776 45865 5797 45921
rect 5853 45865 5874 45921
rect 5776 45844 5874 45865
rect 6201 45863 6299 45884
rect 6201 45807 6222 45863
rect 6278 45807 6299 45863
rect 6201 45786 6299 45807
rect 6633 45863 6731 45884
rect 6633 45807 6654 45863
rect 6710 45807 6731 45863
rect 6633 45786 6731 45807
rect 7015 45877 7113 45898
rect 7015 45821 7036 45877
rect 7092 45821 7113 45877
rect 7015 45800 7113 45821
rect 7287 45877 7385 45898
rect 7287 45821 7308 45877
rect 7364 45821 7385 45877
rect 7287 45800 7385 45821
rect 5776 45505 5874 45526
rect 5776 45449 5797 45505
rect 5853 45449 5874 45505
rect 5776 45428 5874 45449
rect 6201 45505 6299 45526
rect 6201 45449 6222 45505
rect 6278 45449 6299 45505
rect 6201 45428 6299 45449
rect 6633 45505 6731 45526
rect 6633 45449 6654 45505
rect 6710 45449 6731 45505
rect 6633 45428 6731 45449
rect 7015 45482 7113 45503
rect 7015 45426 7036 45482
rect 7092 45426 7113 45482
rect 7015 45405 7113 45426
rect 7287 45482 7385 45503
rect 7287 45426 7308 45482
rect 7364 45426 7385 45482
rect 7287 45405 7385 45426
rect 5776 45131 5874 45152
rect 5776 45075 5797 45131
rect 5853 45075 5874 45131
rect 5776 45054 5874 45075
rect 6201 45073 6299 45094
rect 6201 45017 6222 45073
rect 6278 45017 6299 45073
rect 6201 44996 6299 45017
rect 6633 45073 6731 45094
rect 6633 45017 6654 45073
rect 6710 45017 6731 45073
rect 6633 44996 6731 45017
rect 7015 45087 7113 45108
rect 7015 45031 7036 45087
rect 7092 45031 7113 45087
rect 7015 45010 7113 45031
rect 7287 45087 7385 45108
rect 7287 45031 7308 45087
rect 7364 45031 7385 45087
rect 7287 45010 7385 45031
rect 5776 44715 5874 44736
rect 5776 44659 5797 44715
rect 5853 44659 5874 44715
rect 5776 44638 5874 44659
rect 6201 44715 6299 44736
rect 6201 44659 6222 44715
rect 6278 44659 6299 44715
rect 6201 44638 6299 44659
rect 6633 44715 6731 44736
rect 6633 44659 6654 44715
rect 6710 44659 6731 44715
rect 6633 44638 6731 44659
rect 7015 44692 7113 44713
rect 7015 44636 7036 44692
rect 7092 44636 7113 44692
rect 7015 44615 7113 44636
rect 7287 44692 7385 44713
rect 7287 44636 7308 44692
rect 7364 44636 7385 44692
rect 7287 44615 7385 44636
rect 5776 44341 5874 44362
rect 5776 44285 5797 44341
rect 5853 44285 5874 44341
rect 5776 44264 5874 44285
rect 6201 44283 6299 44304
rect 6201 44227 6222 44283
rect 6278 44227 6299 44283
rect 6201 44206 6299 44227
rect 6633 44283 6731 44304
rect 6633 44227 6654 44283
rect 6710 44227 6731 44283
rect 6633 44206 6731 44227
rect 7015 44297 7113 44318
rect 7015 44241 7036 44297
rect 7092 44241 7113 44297
rect 7015 44220 7113 44241
rect 7287 44297 7385 44318
rect 7287 44241 7308 44297
rect 7364 44241 7385 44297
rect 7287 44220 7385 44241
rect 5776 43925 5874 43946
rect 5776 43869 5797 43925
rect 5853 43869 5874 43925
rect 5776 43848 5874 43869
rect 6201 43925 6299 43946
rect 6201 43869 6222 43925
rect 6278 43869 6299 43925
rect 6201 43848 6299 43869
rect 6633 43925 6731 43946
rect 6633 43869 6654 43925
rect 6710 43869 6731 43925
rect 6633 43848 6731 43869
rect 7015 43902 7113 43923
rect 7015 43846 7036 43902
rect 7092 43846 7113 43902
rect 7015 43825 7113 43846
rect 7287 43902 7385 43923
rect 7287 43846 7308 43902
rect 7364 43846 7385 43902
rect 7287 43825 7385 43846
rect 5776 43551 5874 43572
rect 5776 43495 5797 43551
rect 5853 43495 5874 43551
rect 5776 43474 5874 43495
rect 6201 43493 6299 43514
rect 6201 43437 6222 43493
rect 6278 43437 6299 43493
rect 6201 43416 6299 43437
rect 6633 43493 6731 43514
rect 6633 43437 6654 43493
rect 6710 43437 6731 43493
rect 6633 43416 6731 43437
rect 7015 43507 7113 43528
rect 7015 43451 7036 43507
rect 7092 43451 7113 43507
rect 7015 43430 7113 43451
rect 7287 43507 7385 43528
rect 7287 43451 7308 43507
rect 7364 43451 7385 43507
rect 7287 43430 7385 43451
rect 5776 43135 5874 43156
rect 5776 43079 5797 43135
rect 5853 43079 5874 43135
rect 5776 43058 5874 43079
rect 6201 43135 6299 43156
rect 6201 43079 6222 43135
rect 6278 43079 6299 43135
rect 6201 43058 6299 43079
rect 6633 43135 6731 43156
rect 6633 43079 6654 43135
rect 6710 43079 6731 43135
rect 6633 43058 6731 43079
rect 7015 43112 7113 43133
rect 7015 43056 7036 43112
rect 7092 43056 7113 43112
rect 7015 43035 7113 43056
rect 7287 43112 7385 43133
rect 7287 43056 7308 43112
rect 7364 43056 7385 43112
rect 7287 43035 7385 43056
rect 5776 42761 5874 42782
rect 5776 42705 5797 42761
rect 5853 42705 5874 42761
rect 5776 42684 5874 42705
rect 6201 42703 6299 42724
rect 6201 42647 6222 42703
rect 6278 42647 6299 42703
rect 6201 42626 6299 42647
rect 6633 42703 6731 42724
rect 6633 42647 6654 42703
rect 6710 42647 6731 42703
rect 6633 42626 6731 42647
rect 7015 42717 7113 42738
rect 7015 42661 7036 42717
rect 7092 42661 7113 42717
rect 7015 42640 7113 42661
rect 7287 42717 7385 42738
rect 7287 42661 7308 42717
rect 7364 42661 7385 42717
rect 7287 42640 7385 42661
rect 5776 42345 5874 42366
rect 5776 42289 5797 42345
rect 5853 42289 5874 42345
rect 5776 42268 5874 42289
rect 6201 42345 6299 42366
rect 6201 42289 6222 42345
rect 6278 42289 6299 42345
rect 6201 42268 6299 42289
rect 6633 42345 6731 42366
rect 6633 42289 6654 42345
rect 6710 42289 6731 42345
rect 6633 42268 6731 42289
rect 7015 42322 7113 42343
rect 7015 42266 7036 42322
rect 7092 42266 7113 42322
rect 7015 42245 7113 42266
rect 7287 42322 7385 42343
rect 7287 42266 7308 42322
rect 7364 42266 7385 42322
rect 7287 42245 7385 42266
rect 5776 41971 5874 41992
rect 5776 41915 5797 41971
rect 5853 41915 5874 41971
rect 5776 41894 5874 41915
rect 6201 41913 6299 41934
rect 6201 41857 6222 41913
rect 6278 41857 6299 41913
rect 6201 41836 6299 41857
rect 6633 41913 6731 41934
rect 6633 41857 6654 41913
rect 6710 41857 6731 41913
rect 6633 41836 6731 41857
rect 7015 41927 7113 41948
rect 7015 41871 7036 41927
rect 7092 41871 7113 41927
rect 7015 41850 7113 41871
rect 7287 41927 7385 41948
rect 7287 41871 7308 41927
rect 7364 41871 7385 41927
rect 7287 41850 7385 41871
rect 5776 41555 5874 41576
rect 5776 41499 5797 41555
rect 5853 41499 5874 41555
rect 5776 41478 5874 41499
rect 6201 41555 6299 41576
rect 6201 41499 6222 41555
rect 6278 41499 6299 41555
rect 6201 41478 6299 41499
rect 6633 41555 6731 41576
rect 6633 41499 6654 41555
rect 6710 41499 6731 41555
rect 6633 41478 6731 41499
rect 7015 41532 7113 41553
rect 7015 41476 7036 41532
rect 7092 41476 7113 41532
rect 7015 41455 7113 41476
rect 7287 41532 7385 41553
rect 7287 41476 7308 41532
rect 7364 41476 7385 41532
rect 7287 41455 7385 41476
rect 5776 41181 5874 41202
rect 5776 41125 5797 41181
rect 5853 41125 5874 41181
rect 5776 41104 5874 41125
rect 6201 41123 6299 41144
rect 6201 41067 6222 41123
rect 6278 41067 6299 41123
rect 6201 41046 6299 41067
rect 6633 41123 6731 41144
rect 6633 41067 6654 41123
rect 6710 41067 6731 41123
rect 6633 41046 6731 41067
rect 7015 41137 7113 41158
rect 7015 41081 7036 41137
rect 7092 41081 7113 41137
rect 7015 41060 7113 41081
rect 7287 41137 7385 41158
rect 7287 41081 7308 41137
rect 7364 41081 7385 41137
rect 7287 41060 7385 41081
rect 5776 40765 5874 40786
rect 5776 40709 5797 40765
rect 5853 40709 5874 40765
rect 5776 40688 5874 40709
rect 6201 40765 6299 40786
rect 6201 40709 6222 40765
rect 6278 40709 6299 40765
rect 6201 40688 6299 40709
rect 6633 40765 6731 40786
rect 6633 40709 6654 40765
rect 6710 40709 6731 40765
rect 6633 40688 6731 40709
rect 7015 40742 7113 40763
rect 7015 40686 7036 40742
rect 7092 40686 7113 40742
rect 7015 40665 7113 40686
rect 7287 40742 7385 40763
rect 7287 40686 7308 40742
rect 7364 40686 7385 40742
rect 7287 40665 7385 40686
rect 5776 40391 5874 40412
rect 5776 40335 5797 40391
rect 5853 40335 5874 40391
rect 5776 40314 5874 40335
rect 6201 40333 6299 40354
rect 6201 40277 6222 40333
rect 6278 40277 6299 40333
rect 6201 40256 6299 40277
rect 6633 40333 6731 40354
rect 6633 40277 6654 40333
rect 6710 40277 6731 40333
rect 6633 40256 6731 40277
rect 7015 40347 7113 40368
rect 7015 40291 7036 40347
rect 7092 40291 7113 40347
rect 7015 40270 7113 40291
rect 7287 40347 7385 40368
rect 7287 40291 7308 40347
rect 7364 40291 7385 40347
rect 7287 40270 7385 40291
rect 5776 39975 5874 39996
rect 5776 39919 5797 39975
rect 5853 39919 5874 39975
rect 5776 39898 5874 39919
rect 6201 39975 6299 39996
rect 6201 39919 6222 39975
rect 6278 39919 6299 39975
rect 6201 39898 6299 39919
rect 6633 39975 6731 39996
rect 6633 39919 6654 39975
rect 6710 39919 6731 39975
rect 6633 39898 6731 39919
rect 7015 39952 7113 39973
rect 7015 39896 7036 39952
rect 7092 39896 7113 39952
rect 7015 39875 7113 39896
rect 7287 39952 7385 39973
rect 7287 39896 7308 39952
rect 7364 39896 7385 39952
rect 7287 39875 7385 39896
rect 5776 39601 5874 39622
rect 5776 39545 5797 39601
rect 5853 39545 5874 39601
rect 5776 39524 5874 39545
rect 6201 39543 6299 39564
rect 6201 39487 6222 39543
rect 6278 39487 6299 39543
rect 6201 39466 6299 39487
rect 6633 39543 6731 39564
rect 6633 39487 6654 39543
rect 6710 39487 6731 39543
rect 6633 39466 6731 39487
rect 7015 39557 7113 39578
rect 7015 39501 7036 39557
rect 7092 39501 7113 39557
rect 7015 39480 7113 39501
rect 7287 39557 7385 39578
rect 7287 39501 7308 39557
rect 7364 39501 7385 39557
rect 7287 39480 7385 39501
rect 5776 39185 5874 39206
rect 5776 39129 5797 39185
rect 5853 39129 5874 39185
rect 5776 39108 5874 39129
rect 6201 39185 6299 39206
rect 6201 39129 6222 39185
rect 6278 39129 6299 39185
rect 6201 39108 6299 39129
rect 6633 39185 6731 39206
rect 6633 39129 6654 39185
rect 6710 39129 6731 39185
rect 6633 39108 6731 39129
rect 7015 39162 7113 39183
rect 7015 39106 7036 39162
rect 7092 39106 7113 39162
rect 7015 39085 7113 39106
rect 7287 39162 7385 39183
rect 7287 39106 7308 39162
rect 7364 39106 7385 39162
rect 7287 39085 7385 39106
rect 5776 38811 5874 38832
rect 5776 38755 5797 38811
rect 5853 38755 5874 38811
rect 5776 38734 5874 38755
rect 6201 38753 6299 38774
rect 6201 38697 6222 38753
rect 6278 38697 6299 38753
rect 6201 38676 6299 38697
rect 6633 38753 6731 38774
rect 6633 38697 6654 38753
rect 6710 38697 6731 38753
rect 6633 38676 6731 38697
rect 7015 38767 7113 38788
rect 7015 38711 7036 38767
rect 7092 38711 7113 38767
rect 7015 38690 7113 38711
rect 7287 38767 7385 38788
rect 7287 38711 7308 38767
rect 7364 38711 7385 38767
rect 7287 38690 7385 38711
rect 5776 38395 5874 38416
rect 5776 38339 5797 38395
rect 5853 38339 5874 38395
rect 5776 38318 5874 38339
rect 6201 38395 6299 38416
rect 6201 38339 6222 38395
rect 6278 38339 6299 38395
rect 6201 38318 6299 38339
rect 6633 38395 6731 38416
rect 6633 38339 6654 38395
rect 6710 38339 6731 38395
rect 6633 38318 6731 38339
rect 7015 38372 7113 38393
rect 7015 38316 7036 38372
rect 7092 38316 7113 38372
rect 7015 38295 7113 38316
rect 7287 38372 7385 38393
rect 7287 38316 7308 38372
rect 7364 38316 7385 38372
rect 7287 38295 7385 38316
rect 5776 38021 5874 38042
rect 5776 37965 5797 38021
rect 5853 37965 5874 38021
rect 5776 37944 5874 37965
rect 6201 37963 6299 37984
rect 6201 37907 6222 37963
rect 6278 37907 6299 37963
rect 6201 37886 6299 37907
rect 6633 37963 6731 37984
rect 6633 37907 6654 37963
rect 6710 37907 6731 37963
rect 6633 37886 6731 37907
rect 7015 37977 7113 37998
rect 7015 37921 7036 37977
rect 7092 37921 7113 37977
rect 7015 37900 7113 37921
rect 7287 37977 7385 37998
rect 7287 37921 7308 37977
rect 7364 37921 7385 37977
rect 7287 37900 7385 37921
rect 5776 37605 5874 37626
rect 5776 37549 5797 37605
rect 5853 37549 5874 37605
rect 5776 37528 5874 37549
rect 6201 37605 6299 37626
rect 6201 37549 6222 37605
rect 6278 37549 6299 37605
rect 6201 37528 6299 37549
rect 6633 37605 6731 37626
rect 6633 37549 6654 37605
rect 6710 37549 6731 37605
rect 6633 37528 6731 37549
rect 7015 37582 7113 37603
rect 7015 37526 7036 37582
rect 7092 37526 7113 37582
rect 7015 37505 7113 37526
rect 7287 37582 7385 37603
rect 7287 37526 7308 37582
rect 7364 37526 7385 37582
rect 7287 37505 7385 37526
rect 5776 37231 5874 37252
rect 5776 37175 5797 37231
rect 5853 37175 5874 37231
rect 5776 37154 5874 37175
rect 6201 37173 6299 37194
rect 6201 37117 6222 37173
rect 6278 37117 6299 37173
rect 6201 37096 6299 37117
rect 6633 37173 6731 37194
rect 6633 37117 6654 37173
rect 6710 37117 6731 37173
rect 6633 37096 6731 37117
rect 7015 37187 7113 37208
rect 7015 37131 7036 37187
rect 7092 37131 7113 37187
rect 7015 37110 7113 37131
rect 7287 37187 7385 37208
rect 7287 37131 7308 37187
rect 7364 37131 7385 37187
rect 7287 37110 7385 37131
rect 5776 36815 5874 36836
rect 5776 36759 5797 36815
rect 5853 36759 5874 36815
rect 5776 36738 5874 36759
rect 6201 36815 6299 36836
rect 6201 36759 6222 36815
rect 6278 36759 6299 36815
rect 6201 36738 6299 36759
rect 6633 36815 6731 36836
rect 6633 36759 6654 36815
rect 6710 36759 6731 36815
rect 6633 36738 6731 36759
rect 7015 36792 7113 36813
rect 7015 36736 7036 36792
rect 7092 36736 7113 36792
rect 7015 36715 7113 36736
rect 7287 36792 7385 36813
rect 7287 36736 7308 36792
rect 7364 36736 7385 36792
rect 7287 36715 7385 36736
rect 5776 36441 5874 36462
rect 5776 36385 5797 36441
rect 5853 36385 5874 36441
rect 5776 36364 5874 36385
rect 6201 36383 6299 36404
rect 6201 36327 6222 36383
rect 6278 36327 6299 36383
rect 6201 36306 6299 36327
rect 6633 36383 6731 36404
rect 6633 36327 6654 36383
rect 6710 36327 6731 36383
rect 6633 36306 6731 36327
rect 7015 36397 7113 36418
rect 7015 36341 7036 36397
rect 7092 36341 7113 36397
rect 7015 36320 7113 36341
rect 7287 36397 7385 36418
rect 7287 36341 7308 36397
rect 7364 36341 7385 36397
rect 7287 36320 7385 36341
rect 5776 36025 5874 36046
rect 5776 35969 5797 36025
rect 5853 35969 5874 36025
rect 5776 35948 5874 35969
rect 6201 36025 6299 36046
rect 6201 35969 6222 36025
rect 6278 35969 6299 36025
rect 6201 35948 6299 35969
rect 6633 36025 6731 36046
rect 6633 35969 6654 36025
rect 6710 35969 6731 36025
rect 6633 35948 6731 35969
rect 7015 36002 7113 36023
rect 7015 35946 7036 36002
rect 7092 35946 7113 36002
rect 7015 35925 7113 35946
rect 7287 36002 7385 36023
rect 7287 35946 7308 36002
rect 7364 35946 7385 36002
rect 7287 35925 7385 35946
rect 5776 35651 5874 35672
rect 5776 35595 5797 35651
rect 5853 35595 5874 35651
rect 5776 35574 5874 35595
rect 6201 35593 6299 35614
rect 6201 35537 6222 35593
rect 6278 35537 6299 35593
rect 6201 35516 6299 35537
rect 6633 35593 6731 35614
rect 6633 35537 6654 35593
rect 6710 35537 6731 35593
rect 6633 35516 6731 35537
rect 7015 35607 7113 35628
rect 7015 35551 7036 35607
rect 7092 35551 7113 35607
rect 7015 35530 7113 35551
rect 7287 35607 7385 35628
rect 7287 35551 7308 35607
rect 7364 35551 7385 35607
rect 7287 35530 7385 35551
rect 5776 35235 5874 35256
rect 5776 35179 5797 35235
rect 5853 35179 5874 35235
rect 5776 35158 5874 35179
rect 6201 35235 6299 35256
rect 6201 35179 6222 35235
rect 6278 35179 6299 35235
rect 6201 35158 6299 35179
rect 6633 35235 6731 35256
rect 6633 35179 6654 35235
rect 6710 35179 6731 35235
rect 6633 35158 6731 35179
rect 7015 35212 7113 35233
rect 7015 35156 7036 35212
rect 7092 35156 7113 35212
rect 7015 35135 7113 35156
rect 7287 35212 7385 35233
rect 7287 35156 7308 35212
rect 7364 35156 7385 35212
rect 7287 35135 7385 35156
rect 5776 34861 5874 34882
rect 5776 34805 5797 34861
rect 5853 34805 5874 34861
rect 5776 34784 5874 34805
rect 6201 34803 6299 34824
rect 6201 34747 6222 34803
rect 6278 34747 6299 34803
rect 6201 34726 6299 34747
rect 6633 34803 6731 34824
rect 6633 34747 6654 34803
rect 6710 34747 6731 34803
rect 6633 34726 6731 34747
rect 7015 34817 7113 34838
rect 7015 34761 7036 34817
rect 7092 34761 7113 34817
rect 7015 34740 7113 34761
rect 7287 34817 7385 34838
rect 7287 34761 7308 34817
rect 7364 34761 7385 34817
rect 7287 34740 7385 34761
rect 5776 34445 5874 34466
rect 5776 34389 5797 34445
rect 5853 34389 5874 34445
rect 5776 34368 5874 34389
rect 6201 34445 6299 34466
rect 6201 34389 6222 34445
rect 6278 34389 6299 34445
rect 6201 34368 6299 34389
rect 6633 34445 6731 34466
rect 6633 34389 6654 34445
rect 6710 34389 6731 34445
rect 6633 34368 6731 34389
rect 7015 34422 7113 34443
rect 7015 34366 7036 34422
rect 7092 34366 7113 34422
rect 7015 34345 7113 34366
rect 7287 34422 7385 34443
rect 7287 34366 7308 34422
rect 7364 34366 7385 34422
rect 7287 34345 7385 34366
rect 5776 34071 5874 34092
rect 5776 34015 5797 34071
rect 5853 34015 5874 34071
rect 5776 33994 5874 34015
rect 6201 34013 6299 34034
rect 6201 33957 6222 34013
rect 6278 33957 6299 34013
rect 6201 33936 6299 33957
rect 6633 34013 6731 34034
rect 6633 33957 6654 34013
rect 6710 33957 6731 34013
rect 6633 33936 6731 33957
rect 7015 34027 7113 34048
rect 7015 33971 7036 34027
rect 7092 33971 7113 34027
rect 7015 33950 7113 33971
rect 7287 34027 7385 34048
rect 7287 33971 7308 34027
rect 7364 33971 7385 34027
rect 7287 33950 7385 33971
rect 5776 33655 5874 33676
rect 5776 33599 5797 33655
rect 5853 33599 5874 33655
rect 5776 33578 5874 33599
rect 6201 33655 6299 33676
rect 6201 33599 6222 33655
rect 6278 33599 6299 33655
rect 6201 33578 6299 33599
rect 6633 33655 6731 33676
rect 6633 33599 6654 33655
rect 6710 33599 6731 33655
rect 6633 33578 6731 33599
rect 7015 33632 7113 33653
rect 7015 33576 7036 33632
rect 7092 33576 7113 33632
rect 7015 33555 7113 33576
rect 7287 33632 7385 33653
rect 7287 33576 7308 33632
rect 7364 33576 7385 33632
rect 7287 33555 7385 33576
rect 5776 33281 5874 33302
rect 5776 33225 5797 33281
rect 5853 33225 5874 33281
rect 5776 33204 5874 33225
rect 6201 33223 6299 33244
rect 6201 33167 6222 33223
rect 6278 33167 6299 33223
rect 6201 33146 6299 33167
rect 6633 33223 6731 33244
rect 6633 33167 6654 33223
rect 6710 33167 6731 33223
rect 6633 33146 6731 33167
rect 7015 33237 7113 33258
rect 7015 33181 7036 33237
rect 7092 33181 7113 33237
rect 7015 33160 7113 33181
rect 7287 33237 7385 33258
rect 7287 33181 7308 33237
rect 7364 33181 7385 33237
rect 7287 33160 7385 33181
rect 5776 32865 5874 32886
rect 5776 32809 5797 32865
rect 5853 32809 5874 32865
rect 5776 32788 5874 32809
rect 6201 32865 6299 32886
rect 6201 32809 6222 32865
rect 6278 32809 6299 32865
rect 6201 32788 6299 32809
rect 6633 32865 6731 32886
rect 6633 32809 6654 32865
rect 6710 32809 6731 32865
rect 6633 32788 6731 32809
rect 7015 32842 7113 32863
rect 7015 32786 7036 32842
rect 7092 32786 7113 32842
rect 7015 32765 7113 32786
rect 7287 32842 7385 32863
rect 7287 32786 7308 32842
rect 7364 32786 7385 32842
rect 7287 32765 7385 32786
rect 5776 32491 5874 32512
rect 5776 32435 5797 32491
rect 5853 32435 5874 32491
rect 5776 32414 5874 32435
rect 6201 32433 6299 32454
rect 6201 32377 6222 32433
rect 6278 32377 6299 32433
rect 6201 32356 6299 32377
rect 6633 32433 6731 32454
rect 6633 32377 6654 32433
rect 6710 32377 6731 32433
rect 6633 32356 6731 32377
rect 7015 32447 7113 32468
rect 7015 32391 7036 32447
rect 7092 32391 7113 32447
rect 7015 32370 7113 32391
rect 7287 32447 7385 32468
rect 7287 32391 7308 32447
rect 7364 32391 7385 32447
rect 7287 32370 7385 32391
rect 5776 32075 5874 32096
rect 5776 32019 5797 32075
rect 5853 32019 5874 32075
rect 5776 31998 5874 32019
rect 6201 32075 6299 32096
rect 6201 32019 6222 32075
rect 6278 32019 6299 32075
rect 6201 31998 6299 32019
rect 6633 32075 6731 32096
rect 6633 32019 6654 32075
rect 6710 32019 6731 32075
rect 6633 31998 6731 32019
rect 7015 32052 7113 32073
rect 7015 31996 7036 32052
rect 7092 31996 7113 32052
rect 7015 31975 7113 31996
rect 7287 32052 7385 32073
rect 7287 31996 7308 32052
rect 7364 31996 7385 32052
rect 7287 31975 7385 31996
rect 5776 31701 5874 31722
rect 5776 31645 5797 31701
rect 5853 31645 5874 31701
rect 5776 31624 5874 31645
rect 6201 31643 6299 31664
rect 6201 31587 6222 31643
rect 6278 31587 6299 31643
rect 6201 31566 6299 31587
rect 6633 31643 6731 31664
rect 6633 31587 6654 31643
rect 6710 31587 6731 31643
rect 6633 31566 6731 31587
rect 7015 31657 7113 31678
rect 7015 31601 7036 31657
rect 7092 31601 7113 31657
rect 7015 31580 7113 31601
rect 7287 31657 7385 31678
rect 7287 31601 7308 31657
rect 7364 31601 7385 31657
rect 7287 31580 7385 31601
rect 5776 31285 5874 31306
rect 5776 31229 5797 31285
rect 5853 31229 5874 31285
rect 5776 31208 5874 31229
rect 6201 31285 6299 31306
rect 6201 31229 6222 31285
rect 6278 31229 6299 31285
rect 6201 31208 6299 31229
rect 6633 31285 6731 31306
rect 6633 31229 6654 31285
rect 6710 31229 6731 31285
rect 6633 31208 6731 31229
rect 7015 31262 7113 31283
rect 7015 31206 7036 31262
rect 7092 31206 7113 31262
rect 7015 31185 7113 31206
rect 7287 31262 7385 31283
rect 7287 31206 7308 31262
rect 7364 31206 7385 31262
rect 7287 31185 7385 31206
rect 5776 30911 5874 30932
rect 5776 30855 5797 30911
rect 5853 30855 5874 30911
rect 5776 30834 5874 30855
rect 6201 30853 6299 30874
rect 6201 30797 6222 30853
rect 6278 30797 6299 30853
rect 6201 30776 6299 30797
rect 6633 30853 6731 30874
rect 6633 30797 6654 30853
rect 6710 30797 6731 30853
rect 6633 30776 6731 30797
rect 7015 30867 7113 30888
rect 7015 30811 7036 30867
rect 7092 30811 7113 30867
rect 7015 30790 7113 30811
rect 7287 30867 7385 30888
rect 7287 30811 7308 30867
rect 7364 30811 7385 30867
rect 7287 30790 7385 30811
rect 5776 30495 5874 30516
rect 5776 30439 5797 30495
rect 5853 30439 5874 30495
rect 5776 30418 5874 30439
rect 6201 30495 6299 30516
rect 6201 30439 6222 30495
rect 6278 30439 6299 30495
rect 6201 30418 6299 30439
rect 6633 30495 6731 30516
rect 6633 30439 6654 30495
rect 6710 30439 6731 30495
rect 6633 30418 6731 30439
rect 7015 30472 7113 30493
rect 7015 30416 7036 30472
rect 7092 30416 7113 30472
rect 7015 30395 7113 30416
rect 7287 30472 7385 30493
rect 7287 30416 7308 30472
rect 7364 30416 7385 30472
rect 7287 30395 7385 30416
rect 5776 30121 5874 30142
rect 5776 30065 5797 30121
rect 5853 30065 5874 30121
rect 5776 30044 5874 30065
rect 6201 30063 6299 30084
rect 6201 30007 6222 30063
rect 6278 30007 6299 30063
rect 6201 29986 6299 30007
rect 6633 30063 6731 30084
rect 6633 30007 6654 30063
rect 6710 30007 6731 30063
rect 6633 29986 6731 30007
rect 7015 30077 7113 30098
rect 7015 30021 7036 30077
rect 7092 30021 7113 30077
rect 7015 30000 7113 30021
rect 7287 30077 7385 30098
rect 7287 30021 7308 30077
rect 7364 30021 7385 30077
rect 7287 30000 7385 30021
rect 5776 29705 5874 29726
rect 5776 29649 5797 29705
rect 5853 29649 5874 29705
rect 5776 29628 5874 29649
rect 6201 29705 6299 29726
rect 6201 29649 6222 29705
rect 6278 29649 6299 29705
rect 6201 29628 6299 29649
rect 6633 29705 6731 29726
rect 6633 29649 6654 29705
rect 6710 29649 6731 29705
rect 6633 29628 6731 29649
rect 7015 29682 7113 29703
rect 7015 29626 7036 29682
rect 7092 29626 7113 29682
rect 7015 29605 7113 29626
rect 7287 29682 7385 29703
rect 7287 29626 7308 29682
rect 7364 29626 7385 29682
rect 7287 29605 7385 29626
rect 5776 29331 5874 29352
rect 5776 29275 5797 29331
rect 5853 29275 5874 29331
rect 5776 29254 5874 29275
rect 6201 29273 6299 29294
rect 6201 29217 6222 29273
rect 6278 29217 6299 29273
rect 6201 29196 6299 29217
rect 6633 29273 6731 29294
rect 6633 29217 6654 29273
rect 6710 29217 6731 29273
rect 6633 29196 6731 29217
rect 7015 29287 7113 29308
rect 7015 29231 7036 29287
rect 7092 29231 7113 29287
rect 7015 29210 7113 29231
rect 7287 29287 7385 29308
rect 7287 29231 7308 29287
rect 7364 29231 7385 29287
rect 7287 29210 7385 29231
rect 5776 28915 5874 28936
rect 5776 28859 5797 28915
rect 5853 28859 5874 28915
rect 5776 28838 5874 28859
rect 6201 28915 6299 28936
rect 6201 28859 6222 28915
rect 6278 28859 6299 28915
rect 6201 28838 6299 28859
rect 6633 28915 6731 28936
rect 6633 28859 6654 28915
rect 6710 28859 6731 28915
rect 6633 28838 6731 28859
rect 7015 28892 7113 28913
rect 7015 28836 7036 28892
rect 7092 28836 7113 28892
rect 7015 28815 7113 28836
rect 7287 28892 7385 28913
rect 7287 28836 7308 28892
rect 7364 28836 7385 28892
rect 7287 28815 7385 28836
rect 5776 28541 5874 28562
rect 5776 28485 5797 28541
rect 5853 28485 5874 28541
rect 5776 28464 5874 28485
rect 6201 28483 6299 28504
rect 6201 28427 6222 28483
rect 6278 28427 6299 28483
rect 6201 28406 6299 28427
rect 6633 28483 6731 28504
rect 6633 28427 6654 28483
rect 6710 28427 6731 28483
rect 6633 28406 6731 28427
rect 7015 28497 7113 28518
rect 7015 28441 7036 28497
rect 7092 28441 7113 28497
rect 7015 28420 7113 28441
rect 7287 28497 7385 28518
rect 7287 28441 7308 28497
rect 7364 28441 7385 28497
rect 7287 28420 7385 28441
rect 5776 28125 5874 28146
rect 5776 28069 5797 28125
rect 5853 28069 5874 28125
rect 5776 28048 5874 28069
rect 6201 28125 6299 28146
rect 6201 28069 6222 28125
rect 6278 28069 6299 28125
rect 6201 28048 6299 28069
rect 6633 28125 6731 28146
rect 6633 28069 6654 28125
rect 6710 28069 6731 28125
rect 6633 28048 6731 28069
rect 7015 28102 7113 28123
rect 7015 28046 7036 28102
rect 7092 28046 7113 28102
rect 7015 28025 7113 28046
rect 7287 28102 7385 28123
rect 7287 28046 7308 28102
rect 7364 28046 7385 28102
rect 7287 28025 7385 28046
rect 5776 27751 5874 27772
rect 5776 27695 5797 27751
rect 5853 27695 5874 27751
rect 5776 27674 5874 27695
rect 6201 27693 6299 27714
rect 6201 27637 6222 27693
rect 6278 27637 6299 27693
rect 6201 27616 6299 27637
rect 6633 27693 6731 27714
rect 6633 27637 6654 27693
rect 6710 27637 6731 27693
rect 6633 27616 6731 27637
rect 7015 27707 7113 27728
rect 7015 27651 7036 27707
rect 7092 27651 7113 27707
rect 7015 27630 7113 27651
rect 7287 27707 7385 27728
rect 7287 27651 7308 27707
rect 7364 27651 7385 27707
rect 7287 27630 7385 27651
rect 5776 27335 5874 27356
rect 5776 27279 5797 27335
rect 5853 27279 5874 27335
rect 5776 27258 5874 27279
rect 6201 27335 6299 27356
rect 6201 27279 6222 27335
rect 6278 27279 6299 27335
rect 6201 27258 6299 27279
rect 6633 27335 6731 27356
rect 6633 27279 6654 27335
rect 6710 27279 6731 27335
rect 6633 27258 6731 27279
rect 7015 27312 7113 27333
rect 7015 27256 7036 27312
rect 7092 27256 7113 27312
rect 7015 27235 7113 27256
rect 7287 27312 7385 27333
rect 7287 27256 7308 27312
rect 7364 27256 7385 27312
rect 7287 27235 7385 27256
rect 5776 26961 5874 26982
rect 5776 26905 5797 26961
rect 5853 26905 5874 26961
rect 5776 26884 5874 26905
rect 6201 26903 6299 26924
rect 6201 26847 6222 26903
rect 6278 26847 6299 26903
rect 6201 26826 6299 26847
rect 6633 26903 6731 26924
rect 6633 26847 6654 26903
rect 6710 26847 6731 26903
rect 6633 26826 6731 26847
rect 7015 26917 7113 26938
rect 7015 26861 7036 26917
rect 7092 26861 7113 26917
rect 7015 26840 7113 26861
rect 7287 26917 7385 26938
rect 7287 26861 7308 26917
rect 7364 26861 7385 26917
rect 7287 26840 7385 26861
rect 5776 26545 5874 26566
rect 5776 26489 5797 26545
rect 5853 26489 5874 26545
rect 5776 26468 5874 26489
rect 6201 26545 6299 26566
rect 6201 26489 6222 26545
rect 6278 26489 6299 26545
rect 6201 26468 6299 26489
rect 6633 26545 6731 26566
rect 6633 26489 6654 26545
rect 6710 26489 6731 26545
rect 6633 26468 6731 26489
rect 7015 26522 7113 26543
rect 7015 26466 7036 26522
rect 7092 26466 7113 26522
rect 7015 26445 7113 26466
rect 7287 26522 7385 26543
rect 7287 26466 7308 26522
rect 7364 26466 7385 26522
rect 7287 26445 7385 26466
rect 5776 26171 5874 26192
rect 5776 26115 5797 26171
rect 5853 26115 5874 26171
rect 5776 26094 5874 26115
rect 6201 26113 6299 26134
rect 6201 26057 6222 26113
rect 6278 26057 6299 26113
rect 6201 26036 6299 26057
rect 6633 26113 6731 26134
rect 6633 26057 6654 26113
rect 6710 26057 6731 26113
rect 6633 26036 6731 26057
rect 7015 26127 7113 26148
rect 7015 26071 7036 26127
rect 7092 26071 7113 26127
rect 7015 26050 7113 26071
rect 7287 26127 7385 26148
rect 7287 26071 7308 26127
rect 7364 26071 7385 26127
rect 7287 26050 7385 26071
rect 5776 25755 5874 25776
rect 5776 25699 5797 25755
rect 5853 25699 5874 25755
rect 5776 25678 5874 25699
rect 6201 25755 6299 25776
rect 6201 25699 6222 25755
rect 6278 25699 6299 25755
rect 6201 25678 6299 25699
rect 6633 25755 6731 25776
rect 6633 25699 6654 25755
rect 6710 25699 6731 25755
rect 6633 25678 6731 25699
rect 7015 25732 7113 25753
rect 7015 25676 7036 25732
rect 7092 25676 7113 25732
rect 7015 25655 7113 25676
rect 7287 25732 7385 25753
rect 7287 25676 7308 25732
rect 7364 25676 7385 25732
rect 7287 25655 7385 25676
rect 5776 25381 5874 25402
rect 5776 25325 5797 25381
rect 5853 25325 5874 25381
rect 5776 25304 5874 25325
rect 6201 25323 6299 25344
rect 6201 25267 6222 25323
rect 6278 25267 6299 25323
rect 6201 25246 6299 25267
rect 6633 25323 6731 25344
rect 6633 25267 6654 25323
rect 6710 25267 6731 25323
rect 6633 25246 6731 25267
rect 7015 25337 7113 25358
rect 7015 25281 7036 25337
rect 7092 25281 7113 25337
rect 7015 25260 7113 25281
rect 7287 25337 7385 25358
rect 7287 25281 7308 25337
rect 7364 25281 7385 25337
rect 7287 25260 7385 25281
rect 5776 24965 5874 24986
rect 5776 24909 5797 24965
rect 5853 24909 5874 24965
rect 5776 24888 5874 24909
rect 6201 24965 6299 24986
rect 6201 24909 6222 24965
rect 6278 24909 6299 24965
rect 6201 24888 6299 24909
rect 6633 24965 6731 24986
rect 6633 24909 6654 24965
rect 6710 24909 6731 24965
rect 6633 24888 6731 24909
rect 7015 24942 7113 24963
rect 7015 24886 7036 24942
rect 7092 24886 7113 24942
rect 7015 24865 7113 24886
rect 7287 24942 7385 24963
rect 7287 24886 7308 24942
rect 7364 24886 7385 24942
rect 7287 24865 7385 24886
rect 5776 24591 5874 24612
rect 5776 24535 5797 24591
rect 5853 24535 5874 24591
rect 5776 24514 5874 24535
rect 6201 24533 6299 24554
rect 6201 24477 6222 24533
rect 6278 24477 6299 24533
rect 6201 24456 6299 24477
rect 6633 24533 6731 24554
rect 6633 24477 6654 24533
rect 6710 24477 6731 24533
rect 6633 24456 6731 24477
rect 7015 24547 7113 24568
rect 7015 24491 7036 24547
rect 7092 24491 7113 24547
rect 7015 24470 7113 24491
rect 7287 24547 7385 24568
rect 7287 24491 7308 24547
rect 7364 24491 7385 24547
rect 7287 24470 7385 24491
rect 5776 24175 5874 24196
rect 5776 24119 5797 24175
rect 5853 24119 5874 24175
rect 5776 24098 5874 24119
rect 6201 24175 6299 24196
rect 6201 24119 6222 24175
rect 6278 24119 6299 24175
rect 6201 24098 6299 24119
rect 6633 24175 6731 24196
rect 6633 24119 6654 24175
rect 6710 24119 6731 24175
rect 6633 24098 6731 24119
rect 7015 24152 7113 24173
rect 7015 24096 7036 24152
rect 7092 24096 7113 24152
rect 7015 24075 7113 24096
rect 7287 24152 7385 24173
rect 7287 24096 7308 24152
rect 7364 24096 7385 24152
rect 7287 24075 7385 24096
rect 5776 23801 5874 23822
rect 5776 23745 5797 23801
rect 5853 23745 5874 23801
rect 5776 23724 5874 23745
rect 6201 23743 6299 23764
rect 6201 23687 6222 23743
rect 6278 23687 6299 23743
rect 6201 23666 6299 23687
rect 6633 23743 6731 23764
rect 6633 23687 6654 23743
rect 6710 23687 6731 23743
rect 6633 23666 6731 23687
rect 7015 23757 7113 23778
rect 7015 23701 7036 23757
rect 7092 23701 7113 23757
rect 7015 23680 7113 23701
rect 7287 23757 7385 23778
rect 7287 23701 7308 23757
rect 7364 23701 7385 23757
rect 7287 23680 7385 23701
rect 5776 23385 5874 23406
rect 5776 23329 5797 23385
rect 5853 23329 5874 23385
rect 5776 23308 5874 23329
rect 6201 23385 6299 23406
rect 6201 23329 6222 23385
rect 6278 23329 6299 23385
rect 6201 23308 6299 23329
rect 6633 23385 6731 23406
rect 6633 23329 6654 23385
rect 6710 23329 6731 23385
rect 6633 23308 6731 23329
rect 7015 23362 7113 23383
rect 7015 23306 7036 23362
rect 7092 23306 7113 23362
rect 7015 23285 7113 23306
rect 7287 23362 7385 23383
rect 7287 23306 7308 23362
rect 7364 23306 7385 23362
rect 7287 23285 7385 23306
rect 5776 23011 5874 23032
rect 5776 22955 5797 23011
rect 5853 22955 5874 23011
rect 5776 22934 5874 22955
rect 6201 22953 6299 22974
rect 6201 22897 6222 22953
rect 6278 22897 6299 22953
rect 6201 22876 6299 22897
rect 6633 22953 6731 22974
rect 6633 22897 6654 22953
rect 6710 22897 6731 22953
rect 6633 22876 6731 22897
rect 7015 22967 7113 22988
rect 7015 22911 7036 22967
rect 7092 22911 7113 22967
rect 7015 22890 7113 22911
rect 7287 22967 7385 22988
rect 7287 22911 7308 22967
rect 7364 22911 7385 22967
rect 7287 22890 7385 22911
rect 5776 22595 5874 22616
rect 5776 22539 5797 22595
rect 5853 22539 5874 22595
rect 5776 22518 5874 22539
rect 6201 22595 6299 22616
rect 6201 22539 6222 22595
rect 6278 22539 6299 22595
rect 6201 22518 6299 22539
rect 6633 22595 6731 22616
rect 6633 22539 6654 22595
rect 6710 22539 6731 22595
rect 6633 22518 6731 22539
rect 7015 22572 7113 22593
rect 7015 22516 7036 22572
rect 7092 22516 7113 22572
rect 7015 22495 7113 22516
rect 7287 22572 7385 22593
rect 7287 22516 7308 22572
rect 7364 22516 7385 22572
rect 7287 22495 7385 22516
rect 5776 22221 5874 22242
rect 5776 22165 5797 22221
rect 5853 22165 5874 22221
rect 5776 22144 5874 22165
rect 6201 22163 6299 22184
rect 6201 22107 6222 22163
rect 6278 22107 6299 22163
rect 6201 22086 6299 22107
rect 6633 22163 6731 22184
rect 6633 22107 6654 22163
rect 6710 22107 6731 22163
rect 6633 22086 6731 22107
rect 7015 22177 7113 22198
rect 7015 22121 7036 22177
rect 7092 22121 7113 22177
rect 7015 22100 7113 22121
rect 7287 22177 7385 22198
rect 7287 22121 7308 22177
rect 7364 22121 7385 22177
rect 7287 22100 7385 22121
rect 5776 21805 5874 21826
rect 5776 21749 5797 21805
rect 5853 21749 5874 21805
rect 5776 21728 5874 21749
rect 6201 21805 6299 21826
rect 6201 21749 6222 21805
rect 6278 21749 6299 21805
rect 6201 21728 6299 21749
rect 6633 21805 6731 21826
rect 6633 21749 6654 21805
rect 6710 21749 6731 21805
rect 6633 21728 6731 21749
rect 7015 21782 7113 21803
rect 7015 21726 7036 21782
rect 7092 21726 7113 21782
rect 7015 21705 7113 21726
rect 7287 21782 7385 21803
rect 7287 21726 7308 21782
rect 7364 21726 7385 21782
rect 7287 21705 7385 21726
rect 5776 21431 5874 21452
rect 5776 21375 5797 21431
rect 5853 21375 5874 21431
rect 5776 21354 5874 21375
rect 6201 21373 6299 21394
rect 6201 21317 6222 21373
rect 6278 21317 6299 21373
rect 6201 21296 6299 21317
rect 6633 21373 6731 21394
rect 6633 21317 6654 21373
rect 6710 21317 6731 21373
rect 6633 21296 6731 21317
rect 7015 21387 7113 21408
rect 7015 21331 7036 21387
rect 7092 21331 7113 21387
rect 7015 21310 7113 21331
rect 7287 21387 7385 21408
rect 7287 21331 7308 21387
rect 7364 21331 7385 21387
rect 7287 21310 7385 21331
rect 5776 21015 5874 21036
rect 5776 20959 5797 21015
rect 5853 20959 5874 21015
rect 5776 20938 5874 20959
rect 6201 21015 6299 21036
rect 6201 20959 6222 21015
rect 6278 20959 6299 21015
rect 6201 20938 6299 20959
rect 6633 21015 6731 21036
rect 6633 20959 6654 21015
rect 6710 20959 6731 21015
rect 6633 20938 6731 20959
rect 7015 20992 7113 21013
rect 7015 20936 7036 20992
rect 7092 20936 7113 20992
rect 7015 20915 7113 20936
rect 7287 20992 7385 21013
rect 7287 20936 7308 20992
rect 7364 20936 7385 20992
rect 7287 20915 7385 20936
rect 5776 20641 5874 20662
rect 5776 20585 5797 20641
rect 5853 20585 5874 20641
rect 5776 20564 5874 20585
rect 6201 20583 6299 20604
rect 6201 20527 6222 20583
rect 6278 20527 6299 20583
rect 6201 20506 6299 20527
rect 6633 20583 6731 20604
rect 6633 20527 6654 20583
rect 6710 20527 6731 20583
rect 6633 20506 6731 20527
rect 7015 20597 7113 20618
rect 7015 20541 7036 20597
rect 7092 20541 7113 20597
rect 7015 20520 7113 20541
rect 7287 20597 7385 20618
rect 7287 20541 7308 20597
rect 7364 20541 7385 20597
rect 7287 20520 7385 20541
rect 5776 20225 5874 20246
rect 5776 20169 5797 20225
rect 5853 20169 5874 20225
rect 5776 20148 5874 20169
rect 6201 20225 6299 20246
rect 6201 20169 6222 20225
rect 6278 20169 6299 20225
rect 6201 20148 6299 20169
rect 6633 20225 6731 20246
rect 6633 20169 6654 20225
rect 6710 20169 6731 20225
rect 6633 20148 6731 20169
rect 7015 20202 7113 20223
rect 7015 20146 7036 20202
rect 7092 20146 7113 20202
rect 7015 20125 7113 20146
rect 7287 20202 7385 20223
rect 7287 20146 7308 20202
rect 7364 20146 7385 20202
rect 7287 20125 7385 20146
rect 5776 19851 5874 19872
rect 5776 19795 5797 19851
rect 5853 19795 5874 19851
rect 5776 19774 5874 19795
rect 6201 19793 6299 19814
rect 6201 19737 6222 19793
rect 6278 19737 6299 19793
rect 6201 19716 6299 19737
rect 6633 19793 6731 19814
rect 6633 19737 6654 19793
rect 6710 19737 6731 19793
rect 6633 19716 6731 19737
rect 7015 19807 7113 19828
rect 7015 19751 7036 19807
rect 7092 19751 7113 19807
rect 7015 19730 7113 19751
rect 7287 19807 7385 19828
rect 7287 19751 7308 19807
rect 7364 19751 7385 19807
rect 7287 19730 7385 19751
rect 5776 19435 5874 19456
rect 5776 19379 5797 19435
rect 5853 19379 5874 19435
rect 5776 19358 5874 19379
rect 6201 19435 6299 19456
rect 6201 19379 6222 19435
rect 6278 19379 6299 19435
rect 6201 19358 6299 19379
rect 6633 19435 6731 19456
rect 6633 19379 6654 19435
rect 6710 19379 6731 19435
rect 6633 19358 6731 19379
rect 7015 19412 7113 19433
rect 7015 19356 7036 19412
rect 7092 19356 7113 19412
rect 7015 19335 7113 19356
rect 7287 19412 7385 19433
rect 7287 19356 7308 19412
rect 7364 19356 7385 19412
rect 7287 19335 7385 19356
rect 5776 19061 5874 19082
rect 5776 19005 5797 19061
rect 5853 19005 5874 19061
rect 5776 18984 5874 19005
rect 6201 19003 6299 19024
rect 6201 18947 6222 19003
rect 6278 18947 6299 19003
rect 6201 18926 6299 18947
rect 6633 19003 6731 19024
rect 6633 18947 6654 19003
rect 6710 18947 6731 19003
rect 6633 18926 6731 18947
rect 7015 19017 7113 19038
rect 7015 18961 7036 19017
rect 7092 18961 7113 19017
rect 7015 18940 7113 18961
rect 7287 19017 7385 19038
rect 7287 18961 7308 19017
rect 7364 18961 7385 19017
rect 7287 18940 7385 18961
rect 5776 18645 5874 18666
rect 5776 18589 5797 18645
rect 5853 18589 5874 18645
rect 5776 18568 5874 18589
rect 6201 18645 6299 18666
rect 6201 18589 6222 18645
rect 6278 18589 6299 18645
rect 6201 18568 6299 18589
rect 6633 18645 6731 18666
rect 6633 18589 6654 18645
rect 6710 18589 6731 18645
rect 6633 18568 6731 18589
rect 7015 18622 7113 18643
rect 7015 18566 7036 18622
rect 7092 18566 7113 18622
rect 7015 18545 7113 18566
rect 7287 18622 7385 18643
rect 7287 18566 7308 18622
rect 7364 18566 7385 18622
rect 7287 18545 7385 18566
rect 5776 18271 5874 18292
rect 5776 18215 5797 18271
rect 5853 18215 5874 18271
rect 5776 18194 5874 18215
rect 6201 18213 6299 18234
rect 6201 18157 6222 18213
rect 6278 18157 6299 18213
rect 6201 18136 6299 18157
rect 6633 18213 6731 18234
rect 6633 18157 6654 18213
rect 6710 18157 6731 18213
rect 6633 18136 6731 18157
rect 7015 18227 7113 18248
rect 7015 18171 7036 18227
rect 7092 18171 7113 18227
rect 7015 18150 7113 18171
rect 7287 18227 7385 18248
rect 7287 18171 7308 18227
rect 7364 18171 7385 18227
rect 7287 18150 7385 18171
rect 5776 17855 5874 17876
rect 5776 17799 5797 17855
rect 5853 17799 5874 17855
rect 5776 17778 5874 17799
rect 6201 17855 6299 17876
rect 6201 17799 6222 17855
rect 6278 17799 6299 17855
rect 6201 17778 6299 17799
rect 6633 17855 6731 17876
rect 6633 17799 6654 17855
rect 6710 17799 6731 17855
rect 6633 17778 6731 17799
rect 7015 17832 7113 17853
rect 7015 17776 7036 17832
rect 7092 17776 7113 17832
rect 7015 17755 7113 17776
rect 7287 17832 7385 17853
rect 7287 17776 7308 17832
rect 7364 17776 7385 17832
rect 7287 17755 7385 17776
rect 5776 17481 5874 17502
rect 5776 17425 5797 17481
rect 5853 17425 5874 17481
rect 5776 17404 5874 17425
rect 6201 17423 6299 17444
rect 6201 17367 6222 17423
rect 6278 17367 6299 17423
rect 6201 17346 6299 17367
rect 6633 17423 6731 17444
rect 6633 17367 6654 17423
rect 6710 17367 6731 17423
rect 6633 17346 6731 17367
rect 7015 17437 7113 17458
rect 7015 17381 7036 17437
rect 7092 17381 7113 17437
rect 7015 17360 7113 17381
rect 7287 17437 7385 17458
rect 7287 17381 7308 17437
rect 7364 17381 7385 17437
rect 7287 17360 7385 17381
rect 5776 17065 5874 17086
rect 5776 17009 5797 17065
rect 5853 17009 5874 17065
rect 5776 16988 5874 17009
rect 6201 17065 6299 17086
rect 6201 17009 6222 17065
rect 6278 17009 6299 17065
rect 6201 16988 6299 17009
rect 6633 17065 6731 17086
rect 6633 17009 6654 17065
rect 6710 17009 6731 17065
rect 6633 16988 6731 17009
rect 7015 17042 7113 17063
rect 7015 16986 7036 17042
rect 7092 16986 7113 17042
rect 7015 16965 7113 16986
rect 7287 17042 7382 17063
rect 7287 16986 7308 17042
rect 7364 16986 7382 17042
rect 7287 16965 7382 16986
rect 5776 16691 5874 16712
rect 5776 16635 5797 16691
rect 5853 16635 5874 16691
rect 5776 16614 5874 16635
rect 6201 16633 6299 16654
rect 6201 16577 6222 16633
rect 6278 16577 6299 16633
rect 6201 16556 6299 16577
rect 6633 16633 6731 16654
rect 6633 16577 6654 16633
rect 6710 16577 6731 16633
rect 6633 16556 6731 16577
rect 7015 16647 7113 16668
rect 7015 16591 7036 16647
rect 7092 16591 7113 16647
rect 7015 16570 7113 16591
rect 7287 16647 7385 16668
rect 7287 16591 7308 16647
rect 7364 16591 7385 16647
rect 7287 16570 7385 16591
rect 5776 16275 5874 16296
rect 5776 16219 5797 16275
rect 5853 16219 5874 16275
rect 5776 16198 5874 16219
rect 6201 16275 6299 16296
rect 6201 16219 6222 16275
rect 6278 16219 6299 16275
rect 6201 16198 6299 16219
rect 6633 16275 6731 16296
rect 6633 16219 6654 16275
rect 6710 16219 6731 16275
rect 6633 16198 6731 16219
rect 7015 16252 7113 16273
rect 7015 16196 7036 16252
rect 7092 16196 7113 16252
rect 7015 16175 7113 16196
rect 7287 16252 7385 16273
rect 7287 16196 7308 16252
rect 7364 16196 7385 16252
rect 7287 16175 7385 16196
rect 5776 15901 5874 15922
rect 5776 15845 5797 15901
rect 5853 15845 5874 15901
rect 5776 15824 5874 15845
rect 6201 15843 6299 15864
rect 6201 15787 6222 15843
rect 6278 15787 6299 15843
rect 6201 15766 6299 15787
rect 6633 15843 6731 15864
rect 6633 15787 6654 15843
rect 6710 15787 6731 15843
rect 6633 15766 6731 15787
rect 7015 15857 7113 15878
rect 7015 15801 7036 15857
rect 7092 15801 7113 15857
rect 7015 15780 7113 15801
rect 7287 15857 7385 15878
rect 7287 15801 7308 15857
rect 7364 15801 7385 15857
rect 7287 15780 7385 15801
rect 5776 15485 5874 15506
rect 5776 15429 5797 15485
rect 5853 15429 5874 15485
rect 5776 15408 5874 15429
rect 6201 15485 6299 15506
rect 6201 15429 6222 15485
rect 6278 15429 6299 15485
rect 6201 15408 6299 15429
rect 6633 15485 6731 15506
rect 6633 15429 6654 15485
rect 6710 15429 6731 15485
rect 6633 15408 6731 15429
rect 7015 15462 7113 15483
rect 7015 15406 7036 15462
rect 7092 15406 7113 15462
rect 7015 15385 7113 15406
rect 7287 15462 7385 15483
rect 7287 15406 7308 15462
rect 7364 15406 7385 15462
rect 7287 15385 7385 15406
rect 5776 15111 5874 15132
rect 5776 15055 5797 15111
rect 5853 15055 5874 15111
rect 5776 15034 5874 15055
rect 6201 15053 6299 15074
rect 6201 14997 6222 15053
rect 6278 14997 6299 15053
rect 6201 14976 6299 14997
rect 6633 15053 6731 15074
rect 6633 14997 6654 15053
rect 6710 14997 6731 15053
rect 6633 14976 6731 14997
rect 7015 15067 7113 15088
rect 7015 15011 7036 15067
rect 7092 15011 7113 15067
rect 7015 14990 7113 15011
rect 7287 15067 7385 15088
rect 7287 15011 7308 15067
rect 7364 15011 7385 15067
rect 7287 14990 7385 15011
rect 5776 14695 5874 14716
rect 5776 14639 5797 14695
rect 5853 14639 5874 14695
rect 5776 14618 5874 14639
rect 6201 14695 6299 14716
rect 6201 14639 6222 14695
rect 6278 14639 6299 14695
rect 6201 14618 6299 14639
rect 6633 14695 6731 14716
rect 6633 14639 6654 14695
rect 6710 14639 6731 14695
rect 6633 14618 6731 14639
rect 7015 14672 7113 14693
rect 7015 14616 7036 14672
rect 7092 14616 7113 14672
rect 7015 14595 7113 14616
rect 7287 14672 7385 14693
rect 7287 14616 7308 14672
rect 7364 14616 7385 14672
rect 7287 14595 7385 14616
rect 5776 14321 5874 14342
rect 5776 14265 5797 14321
rect 5853 14265 5874 14321
rect 5776 14244 5874 14265
rect 6201 14263 6299 14284
rect 6201 14207 6222 14263
rect 6278 14207 6299 14263
rect 6201 14186 6299 14207
rect 6633 14263 6731 14284
rect 6633 14207 6654 14263
rect 6710 14207 6731 14263
rect 6633 14186 6731 14207
rect 7015 14277 7113 14298
rect 7015 14221 7036 14277
rect 7092 14221 7113 14277
rect 7015 14200 7113 14221
rect 7287 14277 7385 14298
rect 7287 14221 7308 14277
rect 7364 14221 7385 14277
rect 7287 14200 7385 14221
rect 5776 13905 5874 13926
rect 5776 13849 5797 13905
rect 5853 13849 5874 13905
rect 5776 13828 5874 13849
rect 6201 13905 6299 13926
rect 6201 13849 6222 13905
rect 6278 13849 6299 13905
rect 6201 13828 6299 13849
rect 6633 13905 6731 13926
rect 6633 13849 6654 13905
rect 6710 13849 6731 13905
rect 6633 13828 6731 13849
rect 7015 13882 7113 13903
rect 7015 13826 7036 13882
rect 7092 13826 7113 13882
rect 7015 13805 7113 13826
rect 7287 13882 7385 13903
rect 7287 13826 7308 13882
rect 7364 13826 7385 13882
rect 7287 13805 7385 13826
rect 5776 13531 5874 13552
rect 5776 13475 5797 13531
rect 5853 13475 5874 13531
rect 5776 13454 5874 13475
rect 6201 13473 6299 13494
rect 6201 13417 6222 13473
rect 6278 13417 6299 13473
rect 6201 13396 6299 13417
rect 6633 13473 6731 13494
rect 6633 13417 6654 13473
rect 6710 13417 6731 13473
rect 6633 13396 6731 13417
rect 7015 13487 7113 13508
rect 7015 13431 7036 13487
rect 7092 13431 7113 13487
rect 7015 13410 7113 13431
rect 7287 13487 7385 13508
rect 7287 13431 7308 13487
rect 7364 13431 7385 13487
rect 7287 13410 7385 13431
rect 5776 13115 5874 13136
rect 5776 13059 5797 13115
rect 5853 13059 5874 13115
rect 5776 13038 5874 13059
rect 6201 13115 6299 13136
rect 6201 13059 6222 13115
rect 6278 13059 6299 13115
rect 6201 13038 6299 13059
rect 6633 13115 6731 13136
rect 6633 13059 6654 13115
rect 6710 13059 6731 13115
rect 6633 13038 6731 13059
rect 7015 13092 7113 13113
rect 7015 13036 7036 13092
rect 7092 13036 7113 13092
rect 7015 13015 7113 13036
rect 7287 13092 7385 13113
rect 7287 13036 7308 13092
rect 7364 13036 7385 13092
rect 7287 13015 7385 13036
rect 5776 12741 5874 12762
rect 5776 12685 5797 12741
rect 5853 12685 5874 12741
rect 5776 12664 5874 12685
rect 6201 12683 6299 12704
rect 6201 12627 6222 12683
rect 6278 12627 6299 12683
rect 6201 12606 6299 12627
rect 6633 12683 6731 12704
rect 6633 12627 6654 12683
rect 6710 12627 6731 12683
rect 6633 12606 6731 12627
rect 7015 12697 7113 12718
rect 7015 12641 7036 12697
rect 7092 12641 7113 12697
rect 7015 12620 7113 12641
rect 7287 12697 7385 12718
rect 7287 12641 7308 12697
rect 7364 12641 7385 12697
rect 7287 12620 7385 12641
rect 5776 12325 5874 12346
rect 5776 12269 5797 12325
rect 5853 12269 5874 12325
rect 5776 12248 5874 12269
rect 6201 12325 6299 12346
rect 6201 12269 6222 12325
rect 6278 12269 6299 12325
rect 6201 12248 6299 12269
rect 6633 12325 6731 12346
rect 6633 12269 6654 12325
rect 6710 12269 6731 12325
rect 6633 12248 6731 12269
rect 7015 12302 7113 12323
rect 7015 12246 7036 12302
rect 7092 12246 7113 12302
rect 7015 12225 7113 12246
rect 7287 12302 7385 12323
rect 7287 12246 7308 12302
rect 7364 12246 7385 12302
rect 7287 12225 7385 12246
rect 5776 11951 5874 11972
rect 5776 11895 5797 11951
rect 5853 11895 5874 11951
rect 5776 11874 5874 11895
rect 6201 11893 6299 11914
rect 6201 11837 6222 11893
rect 6278 11837 6299 11893
rect 6201 11816 6299 11837
rect 6633 11893 6731 11914
rect 6633 11837 6654 11893
rect 6710 11837 6731 11893
rect 6633 11816 6731 11837
rect 7015 11907 7113 11928
rect 7015 11851 7036 11907
rect 7092 11851 7113 11907
rect 7015 11830 7113 11851
rect 7287 11907 7385 11928
rect 7287 11851 7308 11907
rect 7364 11851 7385 11907
rect 7287 11830 7385 11851
rect 5776 11535 5874 11556
rect 5776 11479 5797 11535
rect 5853 11479 5874 11535
rect 5776 11458 5874 11479
rect 6201 11535 6299 11556
rect 6201 11479 6222 11535
rect 6278 11479 6299 11535
rect 6201 11458 6299 11479
rect 6633 11535 6731 11556
rect 6633 11479 6654 11535
rect 6710 11479 6731 11535
rect 6633 11458 6731 11479
rect 7015 11512 7113 11533
rect 7015 11456 7036 11512
rect 7092 11456 7113 11512
rect 7015 11435 7113 11456
rect 7287 11512 7385 11533
rect 7287 11456 7308 11512
rect 7364 11456 7385 11512
rect 7287 11435 7385 11456
rect 5776 11161 5874 11182
rect 5776 11105 5797 11161
rect 5853 11105 5874 11161
rect 5776 11084 5874 11105
rect 6201 11103 6299 11124
rect 6201 11047 6222 11103
rect 6278 11047 6299 11103
rect 6201 11026 6299 11047
rect 6633 11103 6731 11124
rect 6633 11047 6654 11103
rect 6710 11047 6731 11103
rect 6633 11026 6731 11047
rect 7015 11117 7113 11138
rect 7015 11061 7036 11117
rect 7092 11061 7113 11117
rect 7015 11040 7113 11061
rect 7287 11117 7385 11138
rect 7287 11061 7308 11117
rect 7364 11061 7385 11117
rect 7287 11040 7385 11061
rect 5776 10745 5874 10766
rect 5776 10689 5797 10745
rect 5853 10689 5874 10745
rect 5776 10668 5874 10689
rect 6201 10745 6299 10766
rect 6201 10689 6222 10745
rect 6278 10689 6299 10745
rect 6201 10668 6299 10689
rect 6633 10745 6731 10766
rect 6633 10689 6654 10745
rect 6710 10689 6731 10745
rect 6633 10668 6731 10689
rect 7015 10722 7113 10743
rect 7015 10666 7036 10722
rect 7092 10666 7113 10722
rect 7015 10645 7113 10666
rect 7287 10722 7385 10743
rect 7287 10666 7308 10722
rect 7364 10666 7385 10722
rect 7287 10645 7385 10666
rect 5776 10371 5874 10392
rect 5776 10315 5797 10371
rect 5853 10315 5874 10371
rect 5776 10294 5874 10315
rect 6201 10313 6299 10334
rect 6201 10257 6222 10313
rect 6278 10257 6299 10313
rect 6201 10236 6299 10257
rect 6633 10313 6731 10334
rect 6633 10257 6654 10313
rect 6710 10257 6731 10313
rect 6633 10236 6731 10257
rect 7015 10327 7113 10348
rect 7015 10271 7036 10327
rect 7092 10271 7113 10327
rect 7015 10250 7113 10271
rect 7287 10327 7385 10348
rect 7287 10271 7308 10327
rect 7364 10271 7385 10327
rect 7287 10250 7385 10271
rect 5776 9955 5874 9976
rect 5776 9899 5797 9955
rect 5853 9899 5874 9955
rect 5776 9878 5874 9899
rect 6201 9955 6299 9976
rect 6201 9899 6222 9955
rect 6278 9899 6299 9955
rect 6201 9878 6299 9899
rect 6633 9955 6731 9976
rect 6633 9899 6654 9955
rect 6710 9899 6731 9955
rect 6633 9878 6731 9899
rect 7015 9932 7113 9953
rect 7015 9876 7036 9932
rect 7092 9876 7113 9932
rect 7015 9855 7113 9876
rect 7287 9932 7385 9953
rect 7287 9876 7308 9932
rect 7364 9876 7385 9932
rect 7287 9855 7385 9876
rect 5776 9581 5874 9602
rect 5776 9525 5797 9581
rect 5853 9525 5874 9581
rect 5776 9504 5874 9525
rect 6201 9523 6299 9544
rect 6201 9467 6222 9523
rect 6278 9467 6299 9523
rect 6201 9446 6299 9467
rect 6633 9523 6731 9544
rect 6633 9467 6654 9523
rect 6710 9467 6731 9523
rect 6633 9446 6731 9467
rect 7015 9537 7113 9558
rect 7015 9481 7036 9537
rect 7092 9481 7113 9537
rect 7015 9460 7113 9481
rect 7287 9537 7385 9558
rect 7287 9481 7308 9537
rect 7364 9481 7385 9537
rect 7287 9460 7385 9481
rect 5776 9165 5874 9186
rect 5776 9109 5797 9165
rect 5853 9109 5874 9165
rect 5776 9088 5874 9109
rect 6201 9165 6299 9186
rect 6201 9109 6222 9165
rect 6278 9109 6299 9165
rect 6201 9088 6299 9109
rect 6633 9165 6731 9186
rect 6633 9109 6654 9165
rect 6710 9109 6731 9165
rect 6633 9088 6731 9109
rect 7015 9142 7113 9163
rect 7015 9086 7036 9142
rect 7092 9086 7113 9142
rect 7015 9065 7113 9086
rect 7287 9142 7385 9163
rect 7287 9086 7308 9142
rect 7364 9086 7385 9142
rect 7287 9065 7385 9086
rect 5776 8791 5874 8812
rect 5776 8735 5797 8791
rect 5853 8735 5874 8791
rect 5776 8714 5874 8735
rect 6201 8733 6299 8754
rect 6201 8677 6222 8733
rect 6278 8677 6299 8733
rect 6201 8656 6299 8677
rect 6633 8733 6731 8754
rect 6633 8677 6654 8733
rect 6710 8677 6731 8733
rect 6633 8656 6731 8677
rect 7015 8747 7113 8768
rect 7015 8691 7036 8747
rect 7092 8691 7113 8747
rect 7015 8670 7113 8691
rect 7287 8747 7385 8768
rect 7287 8691 7308 8747
rect 7364 8691 7385 8747
rect 7287 8670 7385 8691
rect 5776 8375 5874 8396
rect 5776 8319 5797 8375
rect 5853 8319 5874 8375
rect 5776 8298 5874 8319
rect 6201 8375 6299 8396
rect 6201 8319 6222 8375
rect 6278 8319 6299 8375
rect 6201 8298 6299 8319
rect 6633 8375 6731 8396
rect 6633 8319 6654 8375
rect 6710 8319 6731 8375
rect 6633 8298 6731 8319
rect 7015 8352 7113 8373
rect 7015 8296 7036 8352
rect 7092 8296 7113 8352
rect 7015 8275 7113 8296
rect 7287 8352 7385 8373
rect 7287 8296 7308 8352
rect 7364 8296 7385 8352
rect 7287 8275 7385 8296
rect 5776 8001 5874 8022
rect 5776 7945 5797 8001
rect 5853 7945 5874 8001
rect 5776 7924 5874 7945
rect 6201 7943 6299 7964
rect 6201 7887 6222 7943
rect 6278 7887 6299 7943
rect 6201 7866 6299 7887
rect 6633 7943 6731 7964
rect 6633 7887 6654 7943
rect 6710 7887 6731 7943
rect 6633 7866 6731 7887
rect 7015 7957 7113 7978
rect 7015 7901 7036 7957
rect 7092 7901 7113 7957
rect 7015 7880 7113 7901
rect 7287 7957 7385 7978
rect 7287 7901 7308 7957
rect 7364 7901 7385 7957
rect 7287 7880 7385 7901
rect 2486 7508 2584 7606
rect 2911 7508 3009 7606
rect 3343 7508 3441 7606
rect 5776 7585 5874 7606
rect 3725 7485 3823 7583
rect 3997 7485 4095 7583
rect 5776 7529 5797 7585
rect 5853 7529 5874 7585
rect 5776 7508 5874 7529
rect 6201 7585 6299 7606
rect 6201 7529 6222 7585
rect 6278 7529 6299 7585
rect 6201 7508 6299 7529
rect 6633 7585 6731 7606
rect 6633 7529 6654 7585
rect 6710 7529 6731 7585
rect 6633 7508 6731 7529
rect 7015 7562 7113 7583
rect 7015 7506 7036 7562
rect 7092 7506 7113 7562
rect 7015 7485 7113 7506
rect 7287 7562 7385 7583
rect 7287 7506 7308 7562
rect 7364 7506 7385 7562
rect 7287 7485 7385 7506
rect 5776 7211 5874 7232
rect 5776 7155 5797 7211
rect 5853 7155 5874 7211
rect 5776 7134 5874 7155
rect 6201 7153 6299 7174
rect 6201 7097 6222 7153
rect 6278 7097 6299 7153
rect 6201 7076 6299 7097
rect 6633 7153 6731 7174
rect 6633 7097 6654 7153
rect 6710 7097 6731 7153
rect 6633 7076 6731 7097
rect 7015 7167 7113 7188
rect 7015 7111 7036 7167
rect 7092 7111 7113 7167
rect 7015 7090 7113 7111
rect 7287 7167 7385 7188
rect 7287 7111 7308 7167
rect 7364 7111 7385 7167
rect 7287 7090 7385 7111
rect 2486 6718 2584 6816
rect 2911 6718 3009 6816
rect 3343 6718 3441 6816
rect 5776 6795 5874 6816
rect 3725 6695 3823 6793
rect 3997 6695 4095 6793
rect 5776 6739 5797 6795
rect 5853 6739 5874 6795
rect 5776 6718 5874 6739
rect 6201 6795 6299 6816
rect 6201 6739 6222 6795
rect 6278 6739 6299 6795
rect 6201 6718 6299 6739
rect 6633 6795 6731 6816
rect 6633 6739 6654 6795
rect 6710 6739 6731 6795
rect 6633 6718 6731 6739
rect 7015 6772 7113 6793
rect 7015 6716 7036 6772
rect 7092 6716 7113 6772
rect 7015 6695 7113 6716
rect 7287 6772 7385 6793
rect 7287 6716 7308 6772
rect 7364 6716 7385 6772
rect 7287 6695 7385 6716
rect 5776 6421 5874 6442
rect 5776 6365 5797 6421
rect 5853 6365 5874 6421
rect 5776 6344 5874 6365
rect 6201 6363 6299 6384
rect 6201 6307 6222 6363
rect 6278 6307 6299 6363
rect 6201 6286 6299 6307
rect 6633 6363 6731 6384
rect 6633 6307 6654 6363
rect 6710 6307 6731 6363
rect 6633 6286 6731 6307
rect 7015 6377 7113 6398
rect 7015 6321 7036 6377
rect 7092 6321 7113 6377
rect 7015 6300 7113 6321
rect 7287 6377 7385 6398
rect 7287 6321 7308 6377
rect 7364 6321 7385 6377
rect 7287 6300 7385 6321
rect 2486 5928 2584 6026
rect 2911 5928 3009 6026
rect 3343 5928 3441 6026
rect 5776 6005 5874 6026
rect 3725 5905 3823 6003
rect 3997 5905 4095 6003
rect 5776 5949 5797 6005
rect 5853 5949 5874 6005
rect 5776 5928 5874 5949
rect 6201 6005 6299 6026
rect 6201 5949 6222 6005
rect 6278 5949 6299 6005
rect 6201 5928 6299 5949
rect 6633 6005 6731 6026
rect 6633 5949 6654 6005
rect 6710 5949 6731 6005
rect 6633 5928 6731 5949
rect 7015 5982 7113 6003
rect 7015 5926 7036 5982
rect 7092 5926 7113 5982
rect 7015 5905 7113 5926
rect 7287 5982 7385 6003
rect 7287 5926 7308 5982
rect 7364 5926 7385 5982
rect 7287 5905 7385 5926
rect 5776 5631 5874 5652
rect 5776 5575 5797 5631
rect 5853 5575 5874 5631
rect 5776 5554 5874 5575
rect 6201 5573 6299 5594
rect 6201 5517 6222 5573
rect 6278 5517 6299 5573
rect 6201 5496 6299 5517
rect 6633 5573 6731 5594
rect 6633 5517 6654 5573
rect 6710 5517 6731 5573
rect 6633 5496 6731 5517
rect 7015 5587 7113 5608
rect 7015 5531 7036 5587
rect 7092 5531 7113 5587
rect 7015 5510 7113 5531
rect 7287 5587 7385 5608
rect 7287 5531 7308 5587
rect 7364 5531 7385 5587
rect 7287 5510 7385 5531
rect 1155 5115 1253 5213
rect 1427 5115 1525 5213
rect 2486 5138 2584 5236
rect 2911 5138 3009 5236
rect 3343 5138 3441 5236
rect 5776 5215 5874 5236
rect 3725 5115 3823 5213
rect 3997 5115 4095 5213
rect 5776 5159 5797 5215
rect 5853 5159 5874 5215
rect 5776 5138 5874 5159
rect 6201 5215 6299 5236
rect 6201 5159 6222 5215
rect 6278 5159 6299 5215
rect 6201 5138 6299 5159
rect 6633 5215 6731 5236
rect 6633 5159 6654 5215
rect 6710 5159 6731 5215
rect 6633 5138 6731 5159
rect 7015 5192 7113 5213
rect 7015 5136 7036 5192
rect 7092 5136 7113 5192
rect 7015 5115 7113 5136
rect 7287 5192 7385 5213
rect 7287 5136 7308 5192
rect 7364 5136 7385 5192
rect 7287 5115 7385 5136
rect 5776 4841 5874 4862
rect 5776 4785 5797 4841
rect 5853 4785 5874 4841
rect 5776 4764 5874 4785
rect 6201 4783 6299 4804
rect 6201 4727 6222 4783
rect 6278 4727 6299 4783
rect 6201 4706 6299 4727
rect 6633 4783 6731 4804
rect 6633 4727 6654 4783
rect 6710 4727 6731 4783
rect 6633 4706 6731 4727
rect 7015 4797 7113 4818
rect 7015 4741 7036 4797
rect 7092 4741 7113 4797
rect 7015 4720 7113 4741
rect 7287 4797 7385 4818
rect 7287 4741 7308 4797
rect 7364 4741 7385 4797
rect 7287 4720 7385 4741
rect 5776 4425 5874 4446
rect 5776 4369 5797 4425
rect 5853 4369 5874 4425
rect 5776 4348 5874 4369
rect 6201 4425 6299 4446
rect 6201 4369 6222 4425
rect 6278 4369 6299 4425
rect 6201 4348 6299 4369
rect 6633 4425 6731 4446
rect 6633 4369 6654 4425
rect 6710 4369 6731 4425
rect 6633 4348 6731 4369
rect 7015 4402 7113 4423
rect 7015 4346 7036 4402
rect 7092 4346 7113 4402
rect 7015 4325 7113 4346
rect 7287 4402 7385 4423
rect 7287 4346 7308 4402
rect 7364 4346 7385 4402
rect 7287 4325 7385 4346
rect 5776 4051 5874 4072
rect 5776 3995 5797 4051
rect 5853 3995 5874 4051
rect 5776 3974 5874 3995
rect 6201 3993 6299 4014
rect 6201 3937 6222 3993
rect 6278 3937 6299 3993
rect 6201 3916 6299 3937
rect 6633 3993 6731 4014
rect 6633 3937 6654 3993
rect 6710 3937 6731 3993
rect 6633 3916 6731 3937
rect 7015 4007 7113 4028
rect 7015 3951 7036 4007
rect 7092 3951 7113 4007
rect 7015 3930 7113 3951
rect 7287 4007 7385 4028
rect 7287 3951 7308 4007
rect 7364 3951 7385 4007
rect 7287 3930 7385 3951
rect 2921 3542 3019 3640
rect 3346 3542 3444 3640
rect 5776 3635 5874 3656
rect 3725 3535 3823 3633
rect 3997 3535 4095 3633
rect 5776 3579 5797 3635
rect 5853 3579 5874 3635
rect 5776 3558 5874 3579
rect 6201 3635 6299 3656
rect 6201 3579 6222 3635
rect 6278 3579 6299 3635
rect 6201 3558 6299 3579
rect 6633 3635 6731 3656
rect 6633 3579 6654 3635
rect 6710 3579 6731 3635
rect 6633 3558 6731 3579
rect 7015 3612 7113 3633
rect 7015 3556 7036 3612
rect 7092 3556 7113 3612
rect 7015 3535 7113 3556
rect 7287 3612 7385 3633
rect 7287 3556 7308 3612
rect 7364 3556 7385 3612
rect 7287 3535 7385 3556
rect 5776 3261 5874 3282
rect 5776 3205 5797 3261
rect 5853 3205 5874 3261
rect 5776 3184 5874 3205
rect 6201 3203 6299 3224
rect 6201 3147 6222 3203
rect 6278 3147 6299 3203
rect 6201 3126 6299 3147
rect 6633 3203 6731 3224
rect 6633 3147 6654 3203
rect 6710 3147 6731 3203
rect 6633 3126 6731 3147
rect 7015 3217 7113 3238
rect 7015 3161 7036 3217
rect 7092 3161 7113 3217
rect 7015 3140 7113 3161
rect 7287 3217 7385 3238
rect 7287 3161 7308 3217
rect 7364 3161 7385 3217
rect 7287 3140 7385 3161
rect 1751 2745 1849 2843
rect 2023 2745 2121 2843
rect 2921 2752 3019 2850
rect 3346 2752 3444 2850
rect 5776 2845 5874 2866
rect 3725 2745 3823 2843
rect 3997 2745 4095 2843
rect 5776 2789 5797 2845
rect 5853 2789 5874 2845
rect 5776 2768 5874 2789
rect 6201 2845 6299 2866
rect 6201 2789 6222 2845
rect 6278 2789 6299 2845
rect 6201 2768 6299 2789
rect 6633 2845 6731 2866
rect 6633 2789 6654 2845
rect 6710 2789 6731 2845
rect 6633 2768 6731 2789
rect 7015 2822 7113 2843
rect 7015 2766 7036 2822
rect 7092 2766 7113 2822
rect 7015 2745 7113 2766
rect 7287 2822 7385 2843
rect 7287 2766 7308 2822
rect 7364 2766 7385 2822
rect 7287 2745 7385 2766
rect 5776 2471 5874 2492
rect 5776 2415 5797 2471
rect 5853 2415 5874 2471
rect 5776 2394 5874 2415
rect 6201 2413 6299 2434
rect 6201 2357 6222 2413
rect 6278 2357 6299 2413
rect 6201 2336 6299 2357
rect 6633 2413 6731 2434
rect 6633 2357 6654 2413
rect 6710 2357 6731 2413
rect 6633 2336 6731 2357
rect 7015 2427 7113 2448
rect 7015 2371 7036 2427
rect 7092 2371 7113 2427
rect 7015 2350 7113 2371
rect 7287 2427 7385 2448
rect 7287 2371 7308 2427
rect 7364 2371 7385 2427
rect 7287 2350 7385 2371
rect 5776 2055 5874 2076
rect 5776 1999 5797 2055
rect 5853 1999 5874 2055
rect 5776 1978 5874 1999
rect 6201 2055 6299 2076
rect 6201 1999 6222 2055
rect 6278 1999 6299 2055
rect 6201 1978 6299 1999
rect 6633 2055 6731 2076
rect 6633 1999 6654 2055
rect 6710 1999 6731 2055
rect 6633 1978 6731 1999
rect 7015 2032 7113 2053
rect 7015 1976 7036 2032
rect 7092 1976 7113 2032
rect 7015 1955 7113 1976
rect 7287 2032 7385 2053
rect 7287 1976 7308 2032
rect 7364 1976 7385 2032
rect 7287 1955 7385 1976
rect 5776 1681 5874 1702
rect 5776 1625 5797 1681
rect 5853 1625 5874 1681
rect 5776 1604 5874 1625
rect 6201 1623 6299 1644
rect 6201 1567 6222 1623
rect 6278 1567 6299 1623
rect 6201 1546 6299 1567
rect 6633 1623 6731 1644
rect 6633 1567 6654 1623
rect 6710 1567 6731 1623
rect 6633 1546 6731 1567
rect 7015 1637 7113 1658
rect 7015 1581 7036 1637
rect 7092 1581 7113 1637
rect 7015 1560 7113 1581
rect 7287 1637 7385 1658
rect 7287 1581 7308 1637
rect 7364 1581 7385 1637
rect 7287 1560 7385 1581
rect 2921 1172 3019 1270
rect 3346 1172 3444 1270
rect 5776 1265 5874 1286
rect 3725 1165 3823 1263
rect 3997 1165 4095 1263
rect 5776 1209 5797 1265
rect 5853 1209 5874 1265
rect 5776 1188 5874 1209
rect 6201 1265 6299 1286
rect 6201 1209 6222 1265
rect 6278 1209 6299 1265
rect 6201 1188 6299 1209
rect 6633 1265 6731 1286
rect 6633 1209 6654 1265
rect 6710 1209 6731 1265
rect 6633 1188 6731 1209
rect 7015 1242 7113 1263
rect 7015 1186 7036 1242
rect 7092 1186 7113 1242
rect 7015 1165 7113 1186
rect 7287 1242 7385 1263
rect 7287 1186 7308 1242
rect 7364 1186 7385 1242
rect 7287 1165 7385 1186
rect 5776 891 5874 912
rect 5776 835 5797 891
rect 5853 835 5874 891
rect 5776 814 5874 835
rect 6201 833 6299 854
rect 6201 777 6222 833
rect 6278 777 6299 833
rect 6201 756 6299 777
rect 6633 833 6731 854
rect 6633 777 6654 833
rect 6710 777 6731 833
rect 6633 756 6731 777
rect 7015 847 7113 868
rect 7015 791 7036 847
rect 7092 791 7113 847
rect 7015 770 7113 791
rect 7287 847 7385 868
rect 7287 791 7308 847
rect 7364 791 7385 847
rect 7287 770 7385 791
rect 1751 375 1849 473
rect 2023 375 2121 473
rect 2921 382 3019 480
rect 3346 382 3444 480
rect 5776 475 5874 496
rect 3725 375 3823 473
rect 3997 375 4095 473
rect 5776 419 5797 475
rect 5853 419 5874 475
rect 5776 398 5874 419
rect 6201 475 6299 496
rect 6201 419 6222 475
rect 6278 419 6299 475
rect 6201 398 6299 419
rect 6633 475 6731 496
rect 6633 419 6654 475
rect 6710 419 6731 475
rect 6633 398 6731 419
rect 7015 452 7113 473
rect 7015 396 7036 452
rect 7092 396 7113 452
rect 7015 375 7113 396
rect 7287 452 7385 473
rect 7287 396 7308 452
rect 7364 396 7385 452
rect 7287 375 7385 396
use and3_dec  and3_dec_0
timestamp 1707688321
transform 1 0 5554 0 -1 5559
box 0 -60 1948 490
use and3_dec  and3_dec_1
timestamp 1707688321
transform 1 0 5554 0 1 4769
box 0 -60 1948 490
use and3_dec  and3_dec_2
timestamp 1707688321
transform 1 0 5554 0 -1 4769
box 0 -60 1948 490
use and3_dec  and3_dec_3
timestamp 1707688321
transform 1 0 5554 0 1 3979
box 0 -60 1948 490
use and3_dec  and3_dec_4
timestamp 1707688321
transform 1 0 5554 0 -1 3979
box 0 -60 1948 490
use and3_dec  and3_dec_5
timestamp 1707688321
transform 1 0 5554 0 1 3189
box 0 -60 1948 490
use and3_dec  and3_dec_6
timestamp 1707688321
transform 1 0 5554 0 -1 3189
box 0 -60 1948 490
use and3_dec  and3_dec_7
timestamp 1707688321
transform 1 0 5554 0 1 2399
box 0 -60 1948 490
use and3_dec  and3_dec_8
timestamp 1707688321
transform 1 0 5554 0 -1 2399
box 0 -60 1948 490
use and3_dec  and3_dec_9
timestamp 1707688321
transform 1 0 5554 0 1 1609
box 0 -60 1948 490
use and3_dec  and3_dec_10
timestamp 1707688321
transform 1 0 5554 0 -1 1609
box 0 -60 1948 490
use and3_dec  and3_dec_11
timestamp 1707688321
transform 1 0 5554 0 1 819
box 0 -60 1948 490
use and3_dec  and3_dec_12
timestamp 1707688321
transform 1 0 5554 0 -1 819
box 0 -60 1948 490
use and3_dec  and3_dec_13
timestamp 1707688321
transform 1 0 5554 0 1 29
box 0 -60 1948 490
use and3_dec  and3_dec_14
timestamp 1707688321
transform 1 0 5554 0 -1 7139
box 0 -60 1948 490
use and3_dec  and3_dec_15
timestamp 1707688321
transform 1 0 5554 0 1 6349
box 0 -60 1948 490
use and3_dec  and3_dec_16
timestamp 1707688321
transform 1 0 5554 0 1 11879
box 0 -60 1948 490
use and3_dec  and3_dec_17
timestamp 1707688321
transform 1 0 5554 0 -1 11879
box 0 -60 1948 490
use and3_dec  and3_dec_18
timestamp 1707688321
transform 1 0 5554 0 1 11089
box 0 -60 1948 490
use and3_dec  and3_dec_19
timestamp 1707688321
transform 1 0 5554 0 -1 11089
box 0 -60 1948 490
use and3_dec  and3_dec_20
timestamp 1707688321
transform 1 0 5554 0 1 10299
box 0 -60 1948 490
use and3_dec  and3_dec_21
timestamp 1707688321
transform 1 0 5554 0 -1 10299
box 0 -60 1948 490
use and3_dec  and3_dec_22
timestamp 1707688321
transform 1 0 5554 0 1 9509
box 0 -60 1948 490
use and3_dec  and3_dec_23
timestamp 1707688321
transform 1 0 5554 0 -1 9509
box 0 -60 1948 490
use and3_dec  and3_dec_24
timestamp 1707688321
transform 1 0 5554 0 1 8719
box 0 -60 1948 490
use and3_dec  and3_dec_25
timestamp 1707688321
transform 1 0 5554 0 -1 8719
box 0 -60 1948 490
use and3_dec  and3_dec_26
timestamp 1707688321
transform 1 0 5554 0 1 7929
box 0 -60 1948 490
use and3_dec  and3_dec_27
timestamp 1707688321
transform 1 0 5554 0 -1 7929
box 0 -60 1948 490
use and3_dec  and3_dec_28
timestamp 1707688321
transform 1 0 5554 0 1 7139
box 0 -60 1948 490
use and3_dec  and3_dec_29
timestamp 1707688321
transform 1 0 5554 0 -1 6349
box 0 -60 1948 490
use and3_dec  and3_dec_30
timestamp 1707688321
transform 1 0 5554 0 1 5559
box 0 -60 1948 490
use and3_dec  and3_dec_31
timestamp 1707688321
transform 1 0 5554 0 1 18989
box 0 -60 1948 490
use and3_dec  and3_dec_32
timestamp 1707688321
transform 1 0 5554 0 -1 18989
box 0 -60 1948 490
use and3_dec  and3_dec_33
timestamp 1707688321
transform 1 0 5554 0 1 18199
box 0 -60 1948 490
use and3_dec  and3_dec_34
timestamp 1707688321
transform 1 0 5554 0 -1 18199
box 0 -60 1948 490
use and3_dec  and3_dec_35
timestamp 1707688321
transform 1 0 5554 0 1 17409
box 0 -60 1948 490
use and3_dec  and3_dec_36
timestamp 1707688321
transform 1 0 5554 0 -1 17409
box 0 -60 1948 490
use and3_dec  and3_dec_37
timestamp 1707688321
transform 1 0 5554 0 1 16619
box 0 -60 1948 490
use and3_dec  and3_dec_38
timestamp 1707688321
transform 1 0 5554 0 -1 16619
box 0 -60 1948 490
use and3_dec  and3_dec_39
timestamp 1707688321
transform 1 0 5554 0 1 15829
box 0 -60 1948 490
use and3_dec  and3_dec_40
timestamp 1707688321
transform 1 0 5554 0 -1 15829
box 0 -60 1948 490
use and3_dec  and3_dec_41
timestamp 1707688321
transform 1 0 5554 0 1 15039
box 0 -60 1948 490
use and3_dec  and3_dec_42
timestamp 1707688321
transform 1 0 5554 0 -1 15039
box 0 -60 1948 490
use and3_dec  and3_dec_43
timestamp 1707688321
transform 1 0 5554 0 1 14249
box 0 -60 1948 490
use and3_dec  and3_dec_44
timestamp 1707688321
transform 1 0 5554 0 -1 14249
box 0 -60 1948 490
use and3_dec  and3_dec_45
timestamp 1707688321
transform 1 0 5554 0 1 13459
box 0 -60 1948 490
use and3_dec  and3_dec_46
timestamp 1707688321
transform 1 0 5554 0 -1 13459
box 0 -60 1948 490
use and3_dec  and3_dec_47
timestamp 1707688321
transform 1 0 5554 0 1 24519
box 0 -60 1948 490
use and3_dec  and3_dec_48
timestamp 1707688321
transform 1 0 5554 0 -1 24519
box 0 -60 1948 490
use and3_dec  and3_dec_49
timestamp 1707688321
transform 1 0 5554 0 1 23729
box 0 -60 1948 490
use and3_dec  and3_dec_50
timestamp 1707688321
transform 1 0 5554 0 -1 23729
box 0 -60 1948 490
use and3_dec  and3_dec_51
timestamp 1707688321
transform 1 0 5554 0 1 22939
box 0 -60 1948 490
use and3_dec  and3_dec_52
timestamp 1707688321
transform 1 0 5554 0 -1 22939
box 0 -60 1948 490
use and3_dec  and3_dec_53
timestamp 1707688321
transform 1 0 5554 0 1 22149
box 0 -60 1948 490
use and3_dec  and3_dec_54
timestamp 1707688321
transform 1 0 5554 0 -1 22149
box 0 -60 1948 490
use and3_dec  and3_dec_55
timestamp 1707688321
transform 1 0 5554 0 1 21359
box 0 -60 1948 490
use and3_dec  and3_dec_56
timestamp 1707688321
transform 1 0 5554 0 -1 21359
box 0 -60 1948 490
use and3_dec  and3_dec_57
timestamp 1707688321
transform 1 0 5554 0 1 20569
box 0 -60 1948 490
use and3_dec  and3_dec_58
timestamp 1707688321
transform 1 0 5554 0 -1 20569
box 0 -60 1948 490
use and3_dec  and3_dec_59
timestamp 1707688321
transform 1 0 5554 0 1 19779
box 0 -60 1948 490
use and3_dec  and3_dec_60
timestamp 1707688321
transform 1 0 5554 0 -1 19779
box 0 -60 1948 490
use and3_dec  and3_dec_61
timestamp 1707688321
transform 1 0 5554 0 1 12669
box 0 -60 1948 490
use and3_dec  and3_dec_62
timestamp 1707688321
transform 1 0 5554 0 -1 12669
box 0 -60 1948 490
use and3_dec  and3_dec_63
timestamp 1707688321
transform 1 0 5554 0 1 27679
box 0 -60 1948 490
use and3_dec  and3_dec_64
timestamp 1707688321
transform 1 0 5554 0 -1 27679
box 0 -60 1948 490
use and3_dec  and3_dec_65
timestamp 1707688321
transform 1 0 5554 0 1 26889
box 0 -60 1948 490
use and3_dec  and3_dec_66
timestamp 1707688321
transform 1 0 5554 0 -1 26889
box 0 -60 1948 490
use and3_dec  and3_dec_67
timestamp 1707688321
transform 1 0 5554 0 1 26099
box 0 -60 1948 490
use and3_dec  and3_dec_68
timestamp 1707688321
transform 1 0 5554 0 -1 26099
box 0 -60 1948 490
use and3_dec  and3_dec_69
timestamp 1707688321
transform 1 0 5554 0 -1 33999
box 0 -60 1948 490
use and3_dec  and3_dec_70
timestamp 1707688321
transform 1 0 5554 0 1 33209
box 0 -60 1948 490
use and3_dec  and3_dec_71
timestamp 1707688321
transform 1 0 5554 0 -1 33209
box 0 -60 1948 490
use and3_dec  and3_dec_72
timestamp 1707688321
transform 1 0 5554 0 1 32419
box 0 -60 1948 490
use and3_dec  and3_dec_73
timestamp 1707688321
transform 1 0 5554 0 -1 32419
box 0 -60 1948 490
use and3_dec  and3_dec_74
timestamp 1707688321
transform 1 0 5554 0 1 37159
box 0 -60 1948 490
use and3_dec  and3_dec_75
timestamp 1707688321
transform 1 0 5554 0 -1 37159
box 0 -60 1948 490
use and3_dec  and3_dec_76
timestamp 1707688321
transform 1 0 5554 0 1 36369
box 0 -60 1948 490
use and3_dec  and3_dec_77
timestamp 1707688321
transform 1 0 5554 0 -1 36369
box 0 -60 1948 490
use and3_dec  and3_dec_78
timestamp 1707688321
transform 1 0 5554 0 1 35579
box 0 -60 1948 490
use and3_dec  and3_dec_79
timestamp 1707688321
transform 1 0 5554 0 1 31629
box 0 -60 1948 490
use and3_dec  and3_dec_80
timestamp 1707688321
transform 1 0 5554 0 -1 31629
box 0 -60 1948 490
use and3_dec  and3_dec_81
timestamp 1707688321
transform 1 0 5554 0 1 30839
box 0 -60 1948 490
use and3_dec  and3_dec_82
timestamp 1707688321
transform 1 0 5554 0 -1 30839
box 0 -60 1948 490
use and3_dec  and3_dec_83
timestamp 1707688321
transform 1 0 5554 0 -1 35579
box 0 -60 1948 490
use and3_dec  and3_dec_84
timestamp 1707688321
transform 1 0 5554 0 1 34789
box 0 -60 1948 490
use and3_dec  and3_dec_85
timestamp 1707688321
transform 1 0 5554 0 -1 34789
box 0 -60 1948 490
use and3_dec  and3_dec_86
timestamp 1707688321
transform 1 0 5554 0 1 33999
box 0 -60 1948 490
use and3_dec  and3_dec_87
timestamp 1707688321
transform 1 0 5554 0 1 30049
box 0 -60 1948 490
use and3_dec  and3_dec_88
timestamp 1707688321
transform 1 0 5554 0 -1 30049
box 0 -60 1948 490
use and3_dec  and3_dec_89
timestamp 1707688321
transform 1 0 5554 0 1 29259
box 0 -60 1948 490
use and3_dec  and3_dec_90
timestamp 1707688321
transform 1 0 5554 0 -1 29259
box 0 -60 1948 490
use and3_dec  and3_dec_91
timestamp 1707688321
transform 1 0 5554 0 1 28469
box 0 -60 1948 490
use and3_dec  and3_dec_92
timestamp 1707688321
transform 1 0 5554 0 -1 28469
box 0 -60 1948 490
use and3_dec  and3_dec_93
timestamp 1707688321
transform 1 0 5554 0 1 42689
box 0 -60 1948 490
use and3_dec  and3_dec_94
timestamp 1707688321
transform 1 0 5554 0 -1 42689
box 0 -60 1948 490
use and3_dec  and3_dec_95
timestamp 1707688321
transform 1 0 5554 0 1 41899
box 0 -60 1948 490
use and3_dec  and3_dec_96
timestamp 1707688321
transform 1 0 5554 0 -1 41899
box 0 -60 1948 490
use and3_dec  and3_dec_97
timestamp 1707688321
transform 1 0 5554 0 1 41109
box 0 -60 1948 490
use and3_dec  and3_dec_98
timestamp 1707688321
transform 1 0 5554 0 -1 41109
box 0 -60 1948 490
use and3_dec  and3_dec_99
timestamp 1707688321
transform 1 0 5554 0 1 40319
box 0 -60 1948 490
use and3_dec  and3_dec_100
timestamp 1707688321
transform 1 0 5554 0 -1 40319
box 0 -60 1948 490
use and3_dec  and3_dec_101
timestamp 1707688321
transform 1 0 5554 0 1 39529
box 0 -60 1948 490
use and3_dec  and3_dec_102
timestamp 1707688321
transform 1 0 5554 0 -1 39529
box 0 -60 1948 490
use and3_dec  and3_dec_103
timestamp 1707688321
transform 1 0 5554 0 1 38739
box 0 -60 1948 490
use and3_dec  and3_dec_104
timestamp 1707688321
transform 1 0 5554 0 -1 38739
box 0 -60 1948 490
use and3_dec  and3_dec_105
timestamp 1707688321
transform 1 0 5554 0 -1 50589
box 0 -60 1948 490
use and3_dec  and3_dec_106
timestamp 1707688321
transform 1 0 5554 0 1 49799
box 0 -60 1948 490
use and3_dec  and3_dec_107
timestamp 1707688321
transform 1 0 5554 0 -1 49799
box 0 -60 1948 490
use and3_dec  and3_dec_108
timestamp 1707688321
transform 1 0 5554 0 1 49009
box 0 -60 1948 490
use and3_dec  and3_dec_109
timestamp 1707688321
transform 1 0 5554 0 -1 49009
box 0 -60 1948 490
use and3_dec  and3_dec_110
timestamp 1707688321
transform 1 0 5554 0 1 48219
box 0 -60 1948 490
use and3_dec  and3_dec_111
timestamp 1707688321
transform 1 0 5554 0 -1 48219
box 0 -60 1948 490
use and3_dec  and3_dec_112
timestamp 1707688321
transform 1 0 5554 0 1 47429
box 0 -60 1948 490
use and3_dec  and3_dec_113
timestamp 1707688321
transform 1 0 5554 0 -1 47429
box 0 -60 1948 490
use and3_dec  and3_dec_114
timestamp 1707688321
transform 1 0 5554 0 1 46639
box 0 -60 1948 490
use and3_dec  and3_dec_115
timestamp 1707688321
transform 1 0 5554 0 -1 46639
box 0 -60 1948 490
use and3_dec  and3_dec_116
timestamp 1707688321
transform 1 0 5554 0 1 45849
box 0 -60 1948 490
use and3_dec  and3_dec_117
timestamp 1707688321
transform 1 0 5554 0 -1 45849
box 0 -60 1948 490
use and3_dec  and3_dec_118
timestamp 1707688321
transform 1 0 5554 0 1 45059
box 0 -60 1948 490
use and3_dec  and3_dec_119
timestamp 1707688321
transform 1 0 5554 0 -1 45059
box 0 -60 1948 490
use and3_dec  and3_dec_120
timestamp 1707688321
transform 1 0 5554 0 1 44269
box 0 -60 1948 490
use and3_dec  and3_dec_121
timestamp 1707688321
transform 1 0 5554 0 -1 44269
box 0 -60 1948 490
use and3_dec  and3_dec_122
timestamp 1707688321
transform 1 0 5554 0 1 43479
box 0 -60 1948 490
use and3_dec  and3_dec_123
timestamp 1707688321
transform 1 0 5554 0 -1 43479
box 0 -60 1948 490
use and3_dec  and3_dec_124
timestamp 1707688321
transform 1 0 5554 0 1 37949
box 0 -60 1948 490
use and3_dec  and3_dec_125
timestamp 1707688321
transform 1 0 5554 0 -1 37949
box 0 -60 1948 490
use and3_dec  and3_dec_126
timestamp 1707688321
transform 1 0 5554 0 1 25309
box 0 -60 1948 490
use and3_dec  and3_dec_127
timestamp 1707688321
transform 1 0 5554 0 -1 25309
box 0 -60 1948 490
use contact_8  contact_8_0
timestamp 1707688321
transform 1 0 7304 0 1 1577
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1707688321
transform 1 0 7304 0 1 2367
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1707688321
transform 1 0 7304 0 1 787
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1707688321
transform 1 0 7304 0 1 1972
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1707688321
transform 1 0 7304 0 1 2762
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1707688321
transform 1 0 7304 0 1 1182
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1707688321
transform 1 0 7304 0 1 392
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1707688321
transform 1 0 6650 0 1 2353
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1707688321
transform 1 0 6650 0 1 773
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1707688321
transform 1 0 6650 0 1 2785
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1707688321
transform 1 0 6650 0 1 1995
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1707688321
transform 1 0 6650 0 1 1563
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1707688321
transform 1 0 6650 0 1 415
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1707688321
transform 1 0 6650 0 1 1205
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1707688321
transform 1 0 7032 0 1 2367
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1707688321
transform 1 0 7032 0 1 1972
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1707688321
transform 1 0 7032 0 1 1577
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1707688321
transform 1 0 7032 0 1 1182
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1707688321
transform 1 0 7032 0 1 787
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1707688321
transform 1 0 7032 0 1 392
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1707688321
transform 1 0 7032 0 1 2762
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1707688321
transform 1 0 6218 0 1 1563
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1707688321
transform 1 0 6218 0 1 1205
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1707688321
transform 1 0 6218 0 1 773
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1707688321
transform 1 0 6218 0 1 415
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1707688321
transform 1 0 6218 0 1 2785
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1707688321
transform 1 0 6218 0 1 2353
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1707688321
transform 1 0 6218 0 1 1995
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1707688321
transform 1 0 5793 0 1 2785
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1707688321
transform 1 0 5793 0 1 2411
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1707688321
transform 1 0 5793 0 1 1995
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1707688321
transform 1 0 5793 0 1 1621
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1707688321
transform 1 0 5793 0 1 1205
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1707688321
transform 1 0 5793 0 1 831
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1707688321
transform 1 0 5793 0 1 415
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1707688321
transform 1 0 5793 0 1 5945
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1707688321
transform 1 0 5793 0 1 5571
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1707688321
transform 1 0 5793 0 1 5155
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1707688321
transform 1 0 5793 0 1 4781
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1707688321
transform 1 0 5793 0 1 4365
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1707688321
transform 1 0 5793 0 1 3991
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1707688321
transform 1 0 5793 0 1 3575
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1707688321
transform 1 0 5793 0 1 3201
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1707688321
transform 1 0 6218 0 1 5945
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1707688321
transform 1 0 6218 0 1 5513
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1707688321
transform 1 0 6218 0 1 5155
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1707688321
transform 1 0 6218 0 1 4723
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1707688321
transform 1 0 6218 0 1 4365
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1707688321
transform 1 0 6218 0 1 3933
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1707688321
transform 1 0 6218 0 1 3575
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1707688321
transform 1 0 6218 0 1 3143
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1707688321
transform 1 0 6650 0 1 3575
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1707688321
transform 1 0 6650 0 1 5155
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1707688321
transform 1 0 6650 0 1 5945
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1707688321
transform 1 0 6650 0 1 4365
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1707688321
transform 1 0 6650 0 1 3143
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1707688321
transform 1 0 6650 0 1 3933
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1707688321
transform 1 0 6650 0 1 4723
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1707688321
transform 1 0 6650 0 1 5513
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1707688321
transform 1 0 7304 0 1 3947
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1707688321
transform 1 0 7304 0 1 5132
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1707688321
transform 1 0 7304 0 1 3552
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1707688321
transform 1 0 7304 0 1 4342
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1707688321
transform 1 0 7304 0 1 3157
box 0 0 1 1
use contact_8  contact_8_64
timestamp 1707688321
transform 1 0 7304 0 1 5922
box 0 0 1 1
use contact_8  contact_8_65
timestamp 1707688321
transform 1 0 7304 0 1 4737
box 0 0 1 1
use contact_8  contact_8_66
timestamp 1707688321
transform 1 0 7304 0 1 5527
box 0 0 1 1
use contact_8  contact_8_67
timestamp 1707688321
transform 1 0 7032 0 1 4342
box 0 0 1 1
use contact_8  contact_8_68
timestamp 1707688321
transform 1 0 7032 0 1 3947
box 0 0 1 1
use contact_8  contact_8_69
timestamp 1707688321
transform 1 0 7032 0 1 3552
box 0 0 1 1
use contact_8  contact_8_70
timestamp 1707688321
transform 1 0 7032 0 1 3157
box 0 0 1 1
use contact_8  contact_8_71
timestamp 1707688321
transform 1 0 7032 0 1 5922
box 0 0 1 1
use contact_8  contact_8_72
timestamp 1707688321
transform 1 0 7032 0 1 5527
box 0 0 1 1
use contact_8  contact_8_73
timestamp 1707688321
transform 1 0 7032 0 1 5132
box 0 0 1 1
use contact_8  contact_8_74
timestamp 1707688321
transform 1 0 7032 0 1 4737
box 0 0 1 1
use contact_8  contact_8_75
timestamp 1707688321
transform 1 0 7032 0 1 9082
box 0 0 1 1
use contact_8  contact_8_76
timestamp 1707688321
transform 1 0 7304 0 1 6317
box 0 0 1 1
use contact_8  contact_8_77
timestamp 1707688321
transform 1 0 7304 0 1 9082
box 0 0 1 1
use contact_8  contact_8_78
timestamp 1707688321
transform 1 0 7304 0 1 7502
box 0 0 1 1
use contact_8  contact_8_79
timestamp 1707688321
transform 1 0 7304 0 1 8687
box 0 0 1 1
use contact_8  contact_8_80
timestamp 1707688321
transform 1 0 7304 0 1 6712
box 0 0 1 1
use contact_8  contact_8_81
timestamp 1707688321
transform 1 0 7304 0 1 8292
box 0 0 1 1
use contact_8  contact_8_82
timestamp 1707688321
transform 1 0 7304 0 1 7107
box 0 0 1 1
use contact_8  contact_8_83
timestamp 1707688321
transform 1 0 7304 0 1 7897
box 0 0 1 1
use contact_8  contact_8_84
timestamp 1707688321
transform 1 0 6650 0 1 7883
box 0 0 1 1
use contact_8  contact_8_85
timestamp 1707688321
transform 1 0 6650 0 1 7525
box 0 0 1 1
use contact_8  contact_8_86
timestamp 1707688321
transform 1 0 6650 0 1 7093
box 0 0 1 1
use contact_8  contact_8_87
timestamp 1707688321
transform 1 0 6650 0 1 6735
box 0 0 1 1
use contact_8  contact_8_88
timestamp 1707688321
transform 1 0 6650 0 1 9105
box 0 0 1 1
use contact_8  contact_8_89
timestamp 1707688321
transform 1 0 6650 0 1 8673
box 0 0 1 1
use contact_8  contact_8_90
timestamp 1707688321
transform 1 0 6650 0 1 8315
box 0 0 1 1
use contact_8  contact_8_91
timestamp 1707688321
transform 1 0 7032 0 1 8687
box 0 0 1 1
use contact_8  contact_8_92
timestamp 1707688321
transform 1 0 7032 0 1 8292
box 0 0 1 1
use contact_8  contact_8_93
timestamp 1707688321
transform 1 0 7032 0 1 7897
box 0 0 1 1
use contact_8  contact_8_94
timestamp 1707688321
transform 1 0 7032 0 1 7502
box 0 0 1 1
use contact_8  contact_8_95
timestamp 1707688321
transform 1 0 7032 0 1 7107
box 0 0 1 1
use contact_8  contact_8_96
timestamp 1707688321
transform 1 0 7032 0 1 6712
box 0 0 1 1
use contact_8  contact_8_97
timestamp 1707688321
transform 1 0 7032 0 1 6317
box 0 0 1 1
use contact_8  contact_8_98
timestamp 1707688321
transform 1 0 6218 0 1 6735
box 0 0 1 1
use contact_8  contact_8_99
timestamp 1707688321
transform 1 0 6218 0 1 8315
box 0 0 1 1
use contact_8  contact_8_100
timestamp 1707688321
transform 1 0 6218 0 1 7525
box 0 0 1 1
use contact_8  contact_8_101
timestamp 1707688321
transform 1 0 6218 0 1 9105
box 0 0 1 1
use contact_8  contact_8_102
timestamp 1707688321
transform 1 0 6218 0 1 7093
box 0 0 1 1
use contact_8  contact_8_103
timestamp 1707688321
transform 1 0 6218 0 1 7883
box 0 0 1 1
use contact_8  contact_8_104
timestamp 1707688321
transform 1 0 6218 0 1 8673
box 0 0 1 1
use contact_8  contact_8_105
timestamp 1707688321
transform 1 0 5793 0 1 9105
box 0 0 1 1
use contact_8  contact_8_106
timestamp 1707688321
transform 1 0 5793 0 1 8731
box 0 0 1 1
use contact_8  contact_8_107
timestamp 1707688321
transform 1 0 5793 0 1 8315
box 0 0 1 1
use contact_8  contact_8_108
timestamp 1707688321
transform 1 0 5793 0 1 7941
box 0 0 1 1
use contact_8  contact_8_109
timestamp 1707688321
transform 1 0 5793 0 1 7525
box 0 0 1 1
use contact_8  contact_8_110
timestamp 1707688321
transform 1 0 5793 0 1 7151
box 0 0 1 1
use contact_8  contact_8_111
timestamp 1707688321
transform 1 0 5793 0 1 6735
box 0 0 1 1
use contact_8  contact_8_112
timestamp 1707688321
transform 1 0 5793 0 1 6361
box 0 0 1 1
use contact_8  contact_8_113
timestamp 1707688321
transform 1 0 5793 0 1 12265
box 0 0 1 1
use contact_8  contact_8_114
timestamp 1707688321
transform 1 0 5793 0 1 11891
box 0 0 1 1
use contact_8  contact_8_115
timestamp 1707688321
transform 1 0 5793 0 1 11475
box 0 0 1 1
use contact_8  contact_8_116
timestamp 1707688321
transform 1 0 5793 0 1 11101
box 0 0 1 1
use contact_8  contact_8_117
timestamp 1707688321
transform 1 0 5793 0 1 10685
box 0 0 1 1
use contact_8  contact_8_118
timestamp 1707688321
transform 1 0 5793 0 1 10311
box 0 0 1 1
use contact_8  contact_8_119
timestamp 1707688321
transform 1 0 5793 0 1 9895
box 0 0 1 1
use contact_8  contact_8_120
timestamp 1707688321
transform 1 0 5793 0 1 9521
box 0 0 1 1
use contact_8  contact_8_121
timestamp 1707688321
transform 1 0 6218 0 1 10253
box 0 0 1 1
use contact_8  contact_8_122
timestamp 1707688321
transform 1 0 6218 0 1 9895
box 0 0 1 1
use contact_8  contact_8_123
timestamp 1707688321
transform 1 0 6218 0 1 10685
box 0 0 1 1
use contact_8  contact_8_124
timestamp 1707688321
transform 1 0 6218 0 1 12265
box 0 0 1 1
use contact_8  contact_8_125
timestamp 1707688321
transform 1 0 6218 0 1 11833
box 0 0 1 1
use contact_8  contact_8_126
timestamp 1707688321
transform 1 0 6218 0 1 11475
box 0 0 1 1
use contact_8  contact_8_127
timestamp 1707688321
transform 1 0 6218 0 1 11043
box 0 0 1 1
use contact_8  contact_8_128
timestamp 1707688321
transform 1 0 7032 0 1 9477
box 0 0 1 1
use contact_8  contact_8_129
timestamp 1707688321
transform 1 0 6650 0 1 9895
box 0 0 1 1
use contact_8  contact_8_130
timestamp 1707688321
transform 1 0 6650 0 1 11043
box 0 0 1 1
use contact_8  contact_8_131
timestamp 1707688321
transform 1 0 6650 0 1 12265
box 0 0 1 1
use contact_8  contact_8_132
timestamp 1707688321
transform 1 0 6650 0 1 10253
box 0 0 1 1
use contact_8  contact_8_133
timestamp 1707688321
transform 1 0 6650 0 1 11833
box 0 0 1 1
use contact_8  contact_8_134
timestamp 1707688321
transform 1 0 6650 0 1 10685
box 0 0 1 1
use contact_8  contact_8_135
timestamp 1707688321
transform 1 0 6650 0 1 11475
box 0 0 1 1
use contact_8  contact_8_136
timestamp 1707688321
transform 1 0 7304 0 1 12242
box 0 0 1 1
use contact_8  contact_8_137
timestamp 1707688321
transform 1 0 7304 0 1 11847
box 0 0 1 1
use contact_8  contact_8_138
timestamp 1707688321
transform 1 0 7304 0 1 11452
box 0 0 1 1
use contact_8  contact_8_139
timestamp 1707688321
transform 1 0 7304 0 1 11057
box 0 0 1 1
use contact_8  contact_8_140
timestamp 1707688321
transform 1 0 7304 0 1 10662
box 0 0 1 1
use contact_8  contact_8_141
timestamp 1707688321
transform 1 0 7304 0 1 10267
box 0 0 1 1
use contact_8  contact_8_142
timestamp 1707688321
transform 1 0 7304 0 1 9872
box 0 0 1 1
use contact_8  contact_8_143
timestamp 1707688321
transform 1 0 7304 0 1 9477
box 0 0 1 1
use contact_8  contact_8_144
timestamp 1707688321
transform 1 0 7032 0 1 12242
box 0 0 1 1
use contact_8  contact_8_145
timestamp 1707688321
transform 1 0 7032 0 1 11847
box 0 0 1 1
use contact_8  contact_8_146
timestamp 1707688321
transform 1 0 7032 0 1 11452
box 0 0 1 1
use contact_8  contact_8_147
timestamp 1707688321
transform 1 0 7032 0 1 11057
box 0 0 1 1
use contact_8  contact_8_148
timestamp 1707688321
transform 1 0 7032 0 1 10662
box 0 0 1 1
use contact_8  contact_8_149
timestamp 1707688321
transform 1 0 7032 0 1 10267
box 0 0 1 1
use contact_8  contact_8_150
timestamp 1707688321
transform 1 0 7032 0 1 9872
box 0 0 1 1
use contact_8  contact_8_151
timestamp 1707688321
transform 1 0 6218 0 1 9463
box 0 0 1 1
use contact_8  contact_8_152
timestamp 1707688321
transform 1 0 6650 0 1 9463
box 0 0 1 1
use contact_8  contact_8_153
timestamp 1707688321
transform 1 0 6218 0 1 6303
box 0 0 1 1
use contact_8  contact_8_154
timestamp 1707688321
transform 1 0 6650 0 1 6303
box 0 0 1 1
use contact_8  contact_8_155
timestamp 1707688321
transform 1 0 1344 0 1 194
box 0 0 1 1
use contact_8  contact_8_156
timestamp 1707688321
transform 1 0 828 0 1 5724
box 0 0 1 1
use contact_8  contact_8_157
timestamp 1707688321
transform 1 0 748 0 1 5330
box 0 0 1 1
use contact_8  contact_8_158
timestamp 1707688321
transform 1 0 668 0 1 4934
box 0 0 1 1
use contact_8  contact_8_159
timestamp 1707688321
transform 1 0 1424 0 1 2960
box 0 0 1 1
use contact_8  contact_8_160
timestamp 1707688321
transform 1 0 1344 0 1 2564
box 0 0 1 1
use contact_8  contact_8_161
timestamp 1707688321
transform 1 0 1424 0 1 590
box 0 0 1 1
use contact_8  contact_8_162
timestamp 1707688321
transform 1 0 7304 0 1 14612
box 0 0 1 1
use contact_8  contact_8_163
timestamp 1707688321
transform 1 0 7304 0 1 14217
box 0 0 1 1
use contact_8  contact_8_164
timestamp 1707688321
transform 1 0 6650 0 1 13413
box 0 0 1 1
use contact_8  contact_8_165
timestamp 1707688321
transform 1 0 6650 0 1 14635
box 0 0 1 1
use contact_8  contact_8_166
timestamp 1707688321
transform 1 0 6650 0 1 15425
box 0 0 1 1
use contact_8  contact_8_167
timestamp 1707688321
transform 1 0 6650 0 1 14203
box 0 0 1 1
use contact_8  contact_8_168
timestamp 1707688321
transform 1 0 6650 0 1 13055
box 0 0 1 1
use contact_8  contact_8_169
timestamp 1707688321
transform 1 0 6650 0 1 13845
box 0 0 1 1
use contact_8  contact_8_170
timestamp 1707688321
transform 1 0 6650 0 1 14993
box 0 0 1 1
use contact_8  contact_8_171
timestamp 1707688321
transform 1 0 7032 0 1 14612
box 0 0 1 1
use contact_8  contact_8_172
timestamp 1707688321
transform 1 0 7032 0 1 13427
box 0 0 1 1
use contact_8  contact_8_173
timestamp 1707688321
transform 1 0 7032 0 1 15402
box 0 0 1 1
use contact_8  contact_8_174
timestamp 1707688321
transform 1 0 7032 0 1 15007
box 0 0 1 1
use contact_8  contact_8_175
timestamp 1707688321
transform 1 0 7032 0 1 13032
box 0 0 1 1
use contact_8  contact_8_176
timestamp 1707688321
transform 1 0 7032 0 1 13822
box 0 0 1 1
use contact_8  contact_8_177
timestamp 1707688321
transform 1 0 7032 0 1 14217
box 0 0 1 1
use contact_8  contact_8_178
timestamp 1707688321
transform 1 0 7304 0 1 15007
box 0 0 1 1
use contact_8  contact_8_179
timestamp 1707688321
transform 1 0 7304 0 1 13427
box 0 0 1 1
use contact_8  contact_8_180
timestamp 1707688321
transform 1 0 7304 0 1 13032
box 0 0 1 1
use contact_8  contact_8_181
timestamp 1707688321
transform 1 0 7304 0 1 15402
box 0 0 1 1
use contact_8  contact_8_182
timestamp 1707688321
transform 1 0 7304 0 1 13822
box 0 0 1 1
use contact_8  contact_8_183
timestamp 1707688321
transform 1 0 5793 0 1 13055
box 0 0 1 1
use contact_8  contact_8_184
timestamp 1707688321
transform 1 0 5793 0 1 12681
box 0 0 1 1
use contact_8  contact_8_185
timestamp 1707688321
transform 1 0 5793 0 1 13471
box 0 0 1 1
use contact_8  contact_8_186
timestamp 1707688321
transform 1 0 5793 0 1 15425
box 0 0 1 1
use contact_8  contact_8_187
timestamp 1707688321
transform 1 0 5793 0 1 15051
box 0 0 1 1
use contact_8  contact_8_188
timestamp 1707688321
transform 1 0 5793 0 1 14635
box 0 0 1 1
use contact_8  contact_8_189
timestamp 1707688321
transform 1 0 5793 0 1 14261
box 0 0 1 1
use contact_8  contact_8_190
timestamp 1707688321
transform 1 0 5793 0 1 13845
box 0 0 1 1
use contact_8  contact_8_191
timestamp 1707688321
transform 1 0 6218 0 1 13055
box 0 0 1 1
use contact_8  contact_8_192
timestamp 1707688321
transform 1 0 6218 0 1 15425
box 0 0 1 1
use contact_8  contact_8_193
timestamp 1707688321
transform 1 0 6218 0 1 14993
box 0 0 1 1
use contact_8  contact_8_194
timestamp 1707688321
transform 1 0 6218 0 1 14635
box 0 0 1 1
use contact_8  contact_8_195
timestamp 1707688321
transform 1 0 6218 0 1 14203
box 0 0 1 1
use contact_8  contact_8_196
timestamp 1707688321
transform 1 0 6218 0 1 13845
box 0 0 1 1
use contact_8  contact_8_197
timestamp 1707688321
transform 1 0 6218 0 1 13413
box 0 0 1 1
use contact_8  contact_8_198
timestamp 1707688321
transform 1 0 5793 0 1 18585
box 0 0 1 1
use contact_8  contact_8_199
timestamp 1707688321
transform 1 0 5793 0 1 18211
box 0 0 1 1
use contact_8  contact_8_200
timestamp 1707688321
transform 1 0 5793 0 1 17795
box 0 0 1 1
use contact_8  contact_8_201
timestamp 1707688321
transform 1 0 5793 0 1 17421
box 0 0 1 1
use contact_8  contact_8_202
timestamp 1707688321
transform 1 0 5793 0 1 17005
box 0 0 1 1
use contact_8  contact_8_203
timestamp 1707688321
transform 1 0 5793 0 1 16631
box 0 0 1 1
use contact_8  contact_8_204
timestamp 1707688321
transform 1 0 5793 0 1 16215
box 0 0 1 1
use contact_8  contact_8_205
timestamp 1707688321
transform 1 0 5793 0 1 15841
box 0 0 1 1
use contact_8  contact_8_206
timestamp 1707688321
transform 1 0 6218 0 1 18585
box 0 0 1 1
use contact_8  contact_8_207
timestamp 1707688321
transform 1 0 6218 0 1 18153
box 0 0 1 1
use contact_8  contact_8_208
timestamp 1707688321
transform 1 0 6218 0 1 17795
box 0 0 1 1
use contact_8  contact_8_209
timestamp 1707688321
transform 1 0 6218 0 1 17363
box 0 0 1 1
use contact_8  contact_8_210
timestamp 1707688321
transform 1 0 6218 0 1 17005
box 0 0 1 1
use contact_8  contact_8_211
timestamp 1707688321
transform 1 0 6218 0 1 16573
box 0 0 1 1
use contact_8  contact_8_212
timestamp 1707688321
transform 1 0 6218 0 1 16215
box 0 0 1 1
use contact_8  contact_8_213
timestamp 1707688321
transform 1 0 7032 0 1 18562
box 0 0 1 1
use contact_8  contact_8_214
timestamp 1707688321
transform 1 0 6650 0 1 16215
box 0 0 1 1
use contact_8  contact_8_215
timestamp 1707688321
transform 1 0 6650 0 1 17005
box 0 0 1 1
use contact_8  contact_8_216
timestamp 1707688321
transform 1 0 6650 0 1 18153
box 0 0 1 1
use contact_8  contact_8_217
timestamp 1707688321
transform 1 0 6650 0 1 17363
box 0 0 1 1
use contact_8  contact_8_218
timestamp 1707688321
transform 1 0 6650 0 1 16573
box 0 0 1 1
use contact_8  contact_8_219
timestamp 1707688321
transform 1 0 6650 0 1 17795
box 0 0 1 1
use contact_8  contact_8_220
timestamp 1707688321
transform 1 0 6650 0 1 18585
box 0 0 1 1
use contact_8  contact_8_221
timestamp 1707688321
transform 1 0 7304 0 1 16587
box 0 0 1 1
use contact_8  contact_8_222
timestamp 1707688321
transform 1 0 7304 0 1 18167
box 0 0 1 1
use contact_8  contact_8_223
timestamp 1707688321
transform 1 0 7304 0 1 16982
box 0 0 1 1
use contact_8  contact_8_224
timestamp 1707688321
transform 1 0 7304 0 1 17772
box 0 0 1 1
use contact_8  contact_8_225
timestamp 1707688321
transform 1 0 7304 0 1 16192
box 0 0 1 1
use contact_8  contact_8_226
timestamp 1707688321
transform 1 0 7304 0 1 17377
box 0 0 1 1
use contact_8  contact_8_227
timestamp 1707688321
transform 1 0 7304 0 1 18562
box 0 0 1 1
use contact_8  contact_8_228
timestamp 1707688321
transform 1 0 7032 0 1 17772
box 0 0 1 1
use contact_8  contact_8_229
timestamp 1707688321
transform 1 0 7032 0 1 17377
box 0 0 1 1
use contact_8  contact_8_230
timestamp 1707688321
transform 1 0 7032 0 1 16982
box 0 0 1 1
use contact_8  contact_8_231
timestamp 1707688321
transform 1 0 7032 0 1 16587
box 0 0 1 1
use contact_8  contact_8_232
timestamp 1707688321
transform 1 0 7032 0 1 16192
box 0 0 1 1
use contact_8  contact_8_233
timestamp 1707688321
transform 1 0 7032 0 1 18167
box 0 0 1 1
use contact_8  contact_8_234
timestamp 1707688321
transform 1 0 6218 0 1 15783
box 0 0 1 1
use contact_8  contact_8_235
timestamp 1707688321
transform 1 0 7032 0 1 15797
box 0 0 1 1
use contact_8  contact_8_236
timestamp 1707688321
transform 1 0 6650 0 1 15783
box 0 0 1 1
use contact_8  contact_8_237
timestamp 1707688321
transform 1 0 7304 0 1 15797
box 0 0 1 1
use contact_8  contact_8_238
timestamp 1707688321
transform 1 0 7032 0 1 21327
box 0 0 1 1
use contact_8  contact_8_239
timestamp 1707688321
transform 1 0 7032 0 1 20932
box 0 0 1 1
use contact_8  contact_8_240
timestamp 1707688321
transform 1 0 7032 0 1 20537
box 0 0 1 1
use contact_8  contact_8_241
timestamp 1707688321
transform 1 0 7032 0 1 20142
box 0 0 1 1
use contact_8  contact_8_242
timestamp 1707688321
transform 1 0 7032 0 1 19747
box 0 0 1 1
use contact_8  contact_8_243
timestamp 1707688321
transform 1 0 7304 0 1 20537
box 0 0 1 1
use contact_8  contact_8_244
timestamp 1707688321
transform 1 0 7304 0 1 19352
box 0 0 1 1
use contact_8  contact_8_245
timestamp 1707688321
transform 1 0 7304 0 1 20142
box 0 0 1 1
use contact_8  contact_8_246
timestamp 1707688321
transform 1 0 7304 0 1 21722
box 0 0 1 1
use contact_8  contact_8_247
timestamp 1707688321
transform 1 0 7304 0 1 21327
box 0 0 1 1
use contact_8  contact_8_248
timestamp 1707688321
transform 1 0 7304 0 1 19747
box 0 0 1 1
use contact_8  contact_8_249
timestamp 1707688321
transform 1 0 7304 0 1 20932
box 0 0 1 1
use contact_8  contact_8_250
timestamp 1707688321
transform 1 0 6650 0 1 20523
box 0 0 1 1
use contact_8  contact_8_251
timestamp 1707688321
transform 1 0 6650 0 1 20165
box 0 0 1 1
use contact_8  contact_8_252
timestamp 1707688321
transform 1 0 6650 0 1 19733
box 0 0 1 1
use contact_8  contact_8_253
timestamp 1707688321
transform 1 0 6650 0 1 19375
box 0 0 1 1
use contact_8  contact_8_254
timestamp 1707688321
transform 1 0 6650 0 1 21745
box 0 0 1 1
use contact_8  contact_8_255
timestamp 1707688321
transform 1 0 6650 0 1 21313
box 0 0 1 1
use contact_8  contact_8_256
timestamp 1707688321
transform 1 0 6650 0 1 20955
box 0 0 1 1
use contact_8  contact_8_257
timestamp 1707688321
transform 1 0 7032 0 1 19352
box 0 0 1 1
use contact_8  contact_8_258
timestamp 1707688321
transform 1 0 7032 0 1 21722
box 0 0 1 1
use contact_8  contact_8_259
timestamp 1707688321
transform 1 0 6218 0 1 20523
box 0 0 1 1
use contact_8  contact_8_260
timestamp 1707688321
transform 1 0 6218 0 1 20955
box 0 0 1 1
use contact_8  contact_8_261
timestamp 1707688321
transform 1 0 6218 0 1 20165
box 0 0 1 1
use contact_8  contact_8_262
timestamp 1707688321
transform 1 0 6218 0 1 19375
box 0 0 1 1
use contact_8  contact_8_263
timestamp 1707688321
transform 1 0 6218 0 1 21745
box 0 0 1 1
use contact_8  contact_8_264
timestamp 1707688321
transform 1 0 6218 0 1 21313
box 0 0 1 1
use contact_8  contact_8_265
timestamp 1707688321
transform 1 0 6218 0 1 19733
box 0 0 1 1
use contact_8  contact_8_266
timestamp 1707688321
transform 1 0 5793 0 1 19001
box 0 0 1 1
use contact_8  contact_8_267
timestamp 1707688321
transform 1 0 5793 0 1 20955
box 0 0 1 1
use contact_8  contact_8_268
timestamp 1707688321
transform 1 0 5793 0 1 19375
box 0 0 1 1
use contact_8  contact_8_269
timestamp 1707688321
transform 1 0 5793 0 1 20581
box 0 0 1 1
use contact_8  contact_8_270
timestamp 1707688321
transform 1 0 5793 0 1 19791
box 0 0 1 1
use contact_8  contact_8_271
timestamp 1707688321
transform 1 0 5793 0 1 20165
box 0 0 1 1
use contact_8  contact_8_272
timestamp 1707688321
transform 1 0 5793 0 1 21745
box 0 0 1 1
use contact_8  contact_8_273
timestamp 1707688321
transform 1 0 5793 0 1 21371
box 0 0 1 1
use contact_8  contact_8_274
timestamp 1707688321
transform 1 0 5793 0 1 22951
box 0 0 1 1
use contact_8  contact_8_275
timestamp 1707688321
transform 1 0 5793 0 1 24905
box 0 0 1 1
use contact_8  contact_8_276
timestamp 1707688321
transform 1 0 5793 0 1 22535
box 0 0 1 1
use contact_8  contact_8_277
timestamp 1707688321
transform 1 0 5793 0 1 24531
box 0 0 1 1
use contact_8  contact_8_278
timestamp 1707688321
transform 1 0 5793 0 1 24115
box 0 0 1 1
use contact_8  contact_8_279
timestamp 1707688321
transform 1 0 5793 0 1 23741
box 0 0 1 1
use contact_8  contact_8_280
timestamp 1707688321
transform 1 0 5793 0 1 22161
box 0 0 1 1
use contact_8  contact_8_281
timestamp 1707688321
transform 1 0 5793 0 1 23325
box 0 0 1 1
use contact_8  contact_8_282
timestamp 1707688321
transform 1 0 6218 0 1 22893
box 0 0 1 1
use contact_8  contact_8_283
timestamp 1707688321
transform 1 0 6218 0 1 22535
box 0 0 1 1
use contact_8  contact_8_284
timestamp 1707688321
transform 1 0 6218 0 1 23683
box 0 0 1 1
use contact_8  contact_8_285
timestamp 1707688321
transform 1 0 6218 0 1 24905
box 0 0 1 1
use contact_8  contact_8_286
timestamp 1707688321
transform 1 0 6218 0 1 23325
box 0 0 1 1
use contact_8  contact_8_287
timestamp 1707688321
transform 1 0 6218 0 1 24115
box 0 0 1 1
use contact_8  contact_8_288
timestamp 1707688321
transform 1 0 6218 0 1 24473
box 0 0 1 1
use contact_8  contact_8_289
timestamp 1707688321
transform 1 0 7032 0 1 22512
box 0 0 1 1
use contact_8  contact_8_290
timestamp 1707688321
transform 1 0 6650 0 1 24115
box 0 0 1 1
use contact_8  contact_8_291
timestamp 1707688321
transform 1 0 6650 0 1 22535
box 0 0 1 1
use contact_8  contact_8_292
timestamp 1707688321
transform 1 0 6650 0 1 23683
box 0 0 1 1
use contact_8  contact_8_293
timestamp 1707688321
transform 1 0 6650 0 1 23325
box 0 0 1 1
use contact_8  contact_8_294
timestamp 1707688321
transform 1 0 6650 0 1 24473
box 0 0 1 1
use contact_8  contact_8_295
timestamp 1707688321
transform 1 0 6650 0 1 22893
box 0 0 1 1
use contact_8  contact_8_296
timestamp 1707688321
transform 1 0 6650 0 1 24905
box 0 0 1 1
use contact_8  contact_8_297
timestamp 1707688321
transform 1 0 7304 0 1 24092
box 0 0 1 1
use contact_8  contact_8_298
timestamp 1707688321
transform 1 0 7304 0 1 23302
box 0 0 1 1
use contact_8  contact_8_299
timestamp 1707688321
transform 1 0 7304 0 1 23697
box 0 0 1 1
use contact_8  contact_8_300
timestamp 1707688321
transform 1 0 7304 0 1 22907
box 0 0 1 1
use contact_8  contact_8_301
timestamp 1707688321
transform 1 0 7304 0 1 22512
box 0 0 1 1
use contact_8  contact_8_302
timestamp 1707688321
transform 1 0 7304 0 1 24882
box 0 0 1 1
use contact_8  contact_8_303
timestamp 1707688321
transform 1 0 7304 0 1 24487
box 0 0 1 1
use contact_8  contact_8_304
timestamp 1707688321
transform 1 0 7032 0 1 24882
box 0 0 1 1
use contact_8  contact_8_305
timestamp 1707688321
transform 1 0 7032 0 1 24487
box 0 0 1 1
use contact_8  contact_8_306
timestamp 1707688321
transform 1 0 7032 0 1 24092
box 0 0 1 1
use contact_8  contact_8_307
timestamp 1707688321
transform 1 0 7032 0 1 23697
box 0 0 1 1
use contact_8  contact_8_308
timestamp 1707688321
transform 1 0 7032 0 1 23302
box 0 0 1 1
use contact_8  contact_8_309
timestamp 1707688321
transform 1 0 7032 0 1 22907
box 0 0 1 1
use contact_8  contact_8_310
timestamp 1707688321
transform 1 0 6218 0 1 22103
box 0 0 1 1
use contact_8  contact_8_311
timestamp 1707688321
transform 1 0 7032 0 1 22117
box 0 0 1 1
use contact_8  contact_8_312
timestamp 1707688321
transform 1 0 6650 0 1 22103
box 0 0 1 1
use contact_8  contact_8_313
timestamp 1707688321
transform 1 0 7304 0 1 22117
box 0 0 1 1
use contact_8  contact_8_314
timestamp 1707688321
transform 1 0 6218 0 1 18943
box 0 0 1 1
use contact_8  contact_8_315
timestamp 1707688321
transform 1 0 6650 0 1 18943
box 0 0 1 1
use contact_8  contact_8_316
timestamp 1707688321
transform 1 0 7304 0 1 18957
box 0 0 1 1
use contact_8  contact_8_317
timestamp 1707688321
transform 1 0 7032 0 1 18957
box 0 0 1 1
use contact_8  contact_8_318
timestamp 1707688321
transform 1 0 6218 0 1 12623
box 0 0 1 1
use contact_8  contact_8_319
timestamp 1707688321
transform 1 0 6650 0 1 12623
box 0 0 1 1
use contact_8  contact_8_320
timestamp 1707688321
transform 1 0 7304 0 1 12637
box 0 0 1 1
use contact_8  contact_8_321
timestamp 1707688321
transform 1 0 7032 0 1 12637
box 0 0 1 1
use contact_8  contact_8_322
timestamp 1707688321
transform 1 0 7304 0 1 27647
box 0 0 1 1
use contact_8  contact_8_323
timestamp 1707688321
transform 1 0 7304 0 1 26067
box 0 0 1 1
use contact_8  contact_8_324
timestamp 1707688321
transform 1 0 7304 0 1 27252
box 0 0 1 1
use contact_8  contact_8_325
timestamp 1707688321
transform 1 0 7304 0 1 25672
box 0 0 1 1
use contact_8  contact_8_326
timestamp 1707688321
transform 1 0 7304 0 1 26462
box 0 0 1 1
use contact_8  contact_8_327
timestamp 1707688321
transform 1 0 7304 0 1 26857
box 0 0 1 1
use contact_8  contact_8_328
timestamp 1707688321
transform 1 0 7304 0 1 28042
box 0 0 1 1
use contact_8  contact_8_329
timestamp 1707688321
transform 1 0 6650 0 1 26053
box 0 0 1 1
use contact_8  contact_8_330
timestamp 1707688321
transform 1 0 6650 0 1 26485
box 0 0 1 1
use contact_8  contact_8_331
timestamp 1707688321
transform 1 0 6650 0 1 27633
box 0 0 1 1
use contact_8  contact_8_332
timestamp 1707688321
transform 1 0 6650 0 1 26843
box 0 0 1 1
use contact_8  contact_8_333
timestamp 1707688321
transform 1 0 6650 0 1 28065
box 0 0 1 1
use contact_8  contact_8_334
timestamp 1707688321
transform 1 0 6650 0 1 27275
box 0 0 1 1
use contact_8  contact_8_335
timestamp 1707688321
transform 1 0 6650 0 1 25695
box 0 0 1 1
use contact_8  contact_8_336
timestamp 1707688321
transform 1 0 7032 0 1 26462
box 0 0 1 1
use contact_8  contact_8_337
timestamp 1707688321
transform 1 0 7032 0 1 26067
box 0 0 1 1
use contact_8  contact_8_338
timestamp 1707688321
transform 1 0 7032 0 1 25672
box 0 0 1 1
use contact_8  contact_8_339
timestamp 1707688321
transform 1 0 7032 0 1 28042
box 0 0 1 1
use contact_8  contact_8_340
timestamp 1707688321
transform 1 0 7032 0 1 27647
box 0 0 1 1
use contact_8  contact_8_341
timestamp 1707688321
transform 1 0 7032 0 1 27252
box 0 0 1 1
use contact_8  contact_8_342
timestamp 1707688321
transform 1 0 7032 0 1 26857
box 0 0 1 1
use contact_8  contact_8_343
timestamp 1707688321
transform 1 0 6218 0 1 26485
box 0 0 1 1
use contact_8  contact_8_344
timestamp 1707688321
transform 1 0 6218 0 1 27633
box 0 0 1 1
use contact_8  contact_8_345
timestamp 1707688321
transform 1 0 6218 0 1 26053
box 0 0 1 1
use contact_8  contact_8_346
timestamp 1707688321
transform 1 0 6218 0 1 27275
box 0 0 1 1
use contact_8  contact_8_347
timestamp 1707688321
transform 1 0 6218 0 1 25695
box 0 0 1 1
use contact_8  contact_8_348
timestamp 1707688321
transform 1 0 6218 0 1 28065
box 0 0 1 1
use contact_8  contact_8_349
timestamp 1707688321
transform 1 0 6218 0 1 26843
box 0 0 1 1
use contact_8  contact_8_350
timestamp 1707688321
transform 1 0 5793 0 1 28065
box 0 0 1 1
use contact_8  contact_8_351
timestamp 1707688321
transform 1 0 5793 0 1 26111
box 0 0 1 1
use contact_8  contact_8_352
timestamp 1707688321
transform 1 0 5793 0 1 25695
box 0 0 1 1
use contact_8  contact_8_353
timestamp 1707688321
transform 1 0 5793 0 1 25321
box 0 0 1 1
use contact_8  contact_8_354
timestamp 1707688321
transform 1 0 5793 0 1 27691
box 0 0 1 1
use contact_8  contact_8_355
timestamp 1707688321
transform 1 0 5793 0 1 27275
box 0 0 1 1
use contact_8  contact_8_356
timestamp 1707688321
transform 1 0 5793 0 1 26901
box 0 0 1 1
use contact_8  contact_8_357
timestamp 1707688321
transform 1 0 5793 0 1 26485
box 0 0 1 1
use contact_8  contact_8_358
timestamp 1707688321
transform 1 0 6218 0 1 28855
box 0 0 1 1
use contact_8  contact_8_359
timestamp 1707688321
transform 1 0 5793 0 1 31225
box 0 0 1 1
use contact_8  contact_8_360
timestamp 1707688321
transform 1 0 5793 0 1 30851
box 0 0 1 1
use contact_8  contact_8_361
timestamp 1707688321
transform 1 0 5793 0 1 30435
box 0 0 1 1
use contact_8  contact_8_362
timestamp 1707688321
transform 1 0 5793 0 1 30061
box 0 0 1 1
use contact_8  contact_8_363
timestamp 1707688321
transform 1 0 5793 0 1 29645
box 0 0 1 1
use contact_8  contact_8_364
timestamp 1707688321
transform 1 0 5793 0 1 29271
box 0 0 1 1
use contact_8  contact_8_365
timestamp 1707688321
transform 1 0 5793 0 1 28855
box 0 0 1 1
use contact_8  contact_8_366
timestamp 1707688321
transform 1 0 5793 0 1 28481
box 0 0 1 1
use contact_8  contact_8_367
timestamp 1707688321
transform 1 0 6218 0 1 31225
box 0 0 1 1
use contact_8  contact_8_368
timestamp 1707688321
transform 1 0 6218 0 1 30793
box 0 0 1 1
use contact_8  contact_8_369
timestamp 1707688321
transform 1 0 6218 0 1 30435
box 0 0 1 1
use contact_8  contact_8_370
timestamp 1707688321
transform 1 0 6218 0 1 30003
box 0 0 1 1
use contact_8  contact_8_371
timestamp 1707688321
transform 1 0 6218 0 1 29645
box 0 0 1 1
use contact_8  contact_8_372
timestamp 1707688321
transform 1 0 6218 0 1 29213
box 0 0 1 1
use contact_8  contact_8_373
timestamp 1707688321
transform 1 0 6650 0 1 30003
box 0 0 1 1
use contact_8  contact_8_374
timestamp 1707688321
transform 1 0 6650 0 1 31225
box 0 0 1 1
use contact_8  contact_8_375
timestamp 1707688321
transform 1 0 6650 0 1 28855
box 0 0 1 1
use contact_8  contact_8_376
timestamp 1707688321
transform 1 0 6650 0 1 29213
box 0 0 1 1
use contact_8  contact_8_377
timestamp 1707688321
transform 1 0 6650 0 1 29645
box 0 0 1 1
use contact_8  contact_8_378
timestamp 1707688321
transform 1 0 6650 0 1 30435
box 0 0 1 1
use contact_8  contact_8_379
timestamp 1707688321
transform 1 0 6650 0 1 30793
box 0 0 1 1
use contact_8  contact_8_380
timestamp 1707688321
transform 1 0 7304 0 1 28832
box 0 0 1 1
use contact_8  contact_8_381
timestamp 1707688321
transform 1 0 7304 0 1 30807
box 0 0 1 1
use contact_8  contact_8_382
timestamp 1707688321
transform 1 0 7304 0 1 30017
box 0 0 1 1
use contact_8  contact_8_383
timestamp 1707688321
transform 1 0 7304 0 1 31202
box 0 0 1 1
use contact_8  contact_8_384
timestamp 1707688321
transform 1 0 7304 0 1 29622
box 0 0 1 1
use contact_8  contact_8_385
timestamp 1707688321
transform 1 0 7304 0 1 29227
box 0 0 1 1
use contact_8  contact_8_386
timestamp 1707688321
transform 1 0 7304 0 1 30412
box 0 0 1 1
use contact_8  contact_8_387
timestamp 1707688321
transform 1 0 7032 0 1 29227
box 0 0 1 1
use contact_8  contact_8_388
timestamp 1707688321
transform 1 0 7032 0 1 28832
box 0 0 1 1
use contact_8  contact_8_389
timestamp 1707688321
transform 1 0 7032 0 1 31202
box 0 0 1 1
use contact_8  contact_8_390
timestamp 1707688321
transform 1 0 7032 0 1 30807
box 0 0 1 1
use contact_8  contact_8_391
timestamp 1707688321
transform 1 0 7032 0 1 30412
box 0 0 1 1
use contact_8  contact_8_392
timestamp 1707688321
transform 1 0 7032 0 1 30017
box 0 0 1 1
use contact_8  contact_8_393
timestamp 1707688321
transform 1 0 7032 0 1 29622
box 0 0 1 1
use contact_8  contact_8_394
timestamp 1707688321
transform 1 0 6650 0 1 28423
box 0 0 1 1
use contact_8  contact_8_395
timestamp 1707688321
transform 1 0 7304 0 1 28437
box 0 0 1 1
use contact_8  contact_8_396
timestamp 1707688321
transform 1 0 7032 0 1 28437
box 0 0 1 1
use contact_8  contact_8_397
timestamp 1707688321
transform 1 0 6218 0 1 28423
box 0 0 1 1
use contact_8  contact_8_398
timestamp 1707688321
transform 1 0 7032 0 1 34362
box 0 0 1 1
use contact_8  contact_8_399
timestamp 1707688321
transform 1 0 7032 0 1 33967
box 0 0 1 1
use contact_8  contact_8_400
timestamp 1707688321
transform 1 0 7032 0 1 33572
box 0 0 1 1
use contact_8  contact_8_401
timestamp 1707688321
transform 1 0 7304 0 1 33177
box 0 0 1 1
use contact_8  contact_8_402
timestamp 1707688321
transform 1 0 7304 0 1 31992
box 0 0 1 1
use contact_8  contact_8_403
timestamp 1707688321
transform 1 0 7304 0 1 32387
box 0 0 1 1
use contact_8  contact_8_404
timestamp 1707688321
transform 1 0 7304 0 1 33572
box 0 0 1 1
use contact_8  contact_8_405
timestamp 1707688321
transform 1 0 7304 0 1 34362
box 0 0 1 1
use contact_8  contact_8_406
timestamp 1707688321
transform 1 0 7304 0 1 32782
box 0 0 1 1
use contact_8  contact_8_407
timestamp 1707688321
transform 1 0 7304 0 1 33967
box 0 0 1 1
use contact_8  contact_8_408
timestamp 1707688321
transform 1 0 6650 0 1 34743
box 0 0 1 1
use contact_8  contact_8_409
timestamp 1707688321
transform 1 0 6650 0 1 32373
box 0 0 1 1
use contact_8  contact_8_410
timestamp 1707688321
transform 1 0 6650 0 1 34385
box 0 0 1 1
use contact_8  contact_8_411
timestamp 1707688321
transform 1 0 6650 0 1 33953
box 0 0 1 1
use contact_8  contact_8_412
timestamp 1707688321
transform 1 0 6650 0 1 32015
box 0 0 1 1
use contact_8  contact_8_413
timestamp 1707688321
transform 1 0 6650 0 1 33595
box 0 0 1 1
use contact_8  contact_8_414
timestamp 1707688321
transform 1 0 6650 0 1 33163
box 0 0 1 1
use contact_8  contact_8_415
timestamp 1707688321
transform 1 0 6650 0 1 32805
box 0 0 1 1
use contact_8  contact_8_416
timestamp 1707688321
transform 1 0 7032 0 1 33177
box 0 0 1 1
use contact_8  contact_8_417
timestamp 1707688321
transform 1 0 7032 0 1 32782
box 0 0 1 1
use contact_8  contact_8_418
timestamp 1707688321
transform 1 0 7032 0 1 32387
box 0 0 1 1
use contact_8  contact_8_419
timestamp 1707688321
transform 1 0 7032 0 1 31992
box 0 0 1 1
use contact_8  contact_8_420
timestamp 1707688321
transform 1 0 6218 0 1 33163
box 0 0 1 1
use contact_8  contact_8_421
timestamp 1707688321
transform 1 0 6218 0 1 32805
box 0 0 1 1
use contact_8  contact_8_422
timestamp 1707688321
transform 1 0 6218 0 1 32373
box 0 0 1 1
use contact_8  contact_8_423
timestamp 1707688321
transform 1 0 6218 0 1 33595
box 0 0 1 1
use contact_8  contact_8_424
timestamp 1707688321
transform 1 0 6218 0 1 34743
box 0 0 1 1
use contact_8  contact_8_425
timestamp 1707688321
transform 1 0 6218 0 1 33953
box 0 0 1 1
use contact_8  contact_8_426
timestamp 1707688321
transform 1 0 6218 0 1 32015
box 0 0 1 1
use contact_8  contact_8_427
timestamp 1707688321
transform 1 0 6218 0 1 34385
box 0 0 1 1
use contact_8  contact_8_428
timestamp 1707688321
transform 1 0 5793 0 1 32805
box 0 0 1 1
use contact_8  contact_8_429
timestamp 1707688321
transform 1 0 5793 0 1 33221
box 0 0 1 1
use contact_8  contact_8_430
timestamp 1707688321
transform 1 0 5793 0 1 32431
box 0 0 1 1
use contact_8  contact_8_431
timestamp 1707688321
transform 1 0 5793 0 1 33595
box 0 0 1 1
use contact_8  contact_8_432
timestamp 1707688321
transform 1 0 5793 0 1 34011
box 0 0 1 1
use contact_8  contact_8_433
timestamp 1707688321
transform 1 0 5793 0 1 34385
box 0 0 1 1
use contact_8  contact_8_434
timestamp 1707688321
transform 1 0 5793 0 1 32015
box 0 0 1 1
use contact_8  contact_8_435
timestamp 1707688321
transform 1 0 5793 0 1 35175
box 0 0 1 1
use contact_8  contact_8_436
timestamp 1707688321
transform 1 0 5793 0 1 36381
box 0 0 1 1
use contact_8  contact_8_437
timestamp 1707688321
transform 1 0 5793 0 1 37545
box 0 0 1 1
use contact_8  contact_8_438
timestamp 1707688321
transform 1 0 5793 0 1 35591
box 0 0 1 1
use contact_8  contact_8_439
timestamp 1707688321
transform 1 0 5793 0 1 37171
box 0 0 1 1
use contact_8  contact_8_440
timestamp 1707688321
transform 1 0 5793 0 1 35965
box 0 0 1 1
use contact_8  contact_8_441
timestamp 1707688321
transform 1 0 5793 0 1 36755
box 0 0 1 1
use contact_8  contact_8_442
timestamp 1707688321
transform 1 0 6218 0 1 37903
box 0 0 1 1
use contact_8  contact_8_443
timestamp 1707688321
transform 1 0 6218 0 1 37545
box 0 0 1 1
use contact_8  contact_8_444
timestamp 1707688321
transform 1 0 6218 0 1 37113
box 0 0 1 1
use contact_8  contact_8_445
timestamp 1707688321
transform 1 0 6218 0 1 36755
box 0 0 1 1
use contact_8  contact_8_446
timestamp 1707688321
transform 1 0 6218 0 1 36323
box 0 0 1 1
use contact_8  contact_8_447
timestamp 1707688321
transform 1 0 6218 0 1 35965
box 0 0 1 1
use contact_8  contact_8_448
timestamp 1707688321
transform 1 0 6218 0 1 35533
box 0 0 1 1
use contact_8  contact_8_449
timestamp 1707688321
transform 1 0 6218 0 1 35175
box 0 0 1 1
use contact_8  contact_8_450
timestamp 1707688321
transform 1 0 7032 0 1 35942
box 0 0 1 1
use contact_8  contact_8_451
timestamp 1707688321
transform 1 0 6650 0 1 37903
box 0 0 1 1
use contact_8  contact_8_452
timestamp 1707688321
transform 1 0 6650 0 1 37545
box 0 0 1 1
use contact_8  contact_8_453
timestamp 1707688321
transform 1 0 6650 0 1 35533
box 0 0 1 1
use contact_8  contact_8_454
timestamp 1707688321
transform 1 0 6650 0 1 37113
box 0 0 1 1
use contact_8  contact_8_455
timestamp 1707688321
transform 1 0 6650 0 1 35965
box 0 0 1 1
use contact_8  contact_8_456
timestamp 1707688321
transform 1 0 6650 0 1 36755
box 0 0 1 1
use contact_8  contact_8_457
timestamp 1707688321
transform 1 0 6650 0 1 35175
box 0 0 1 1
use contact_8  contact_8_458
timestamp 1707688321
transform 1 0 6650 0 1 36323
box 0 0 1 1
use contact_8  contact_8_459
timestamp 1707688321
transform 1 0 7304 0 1 37522
box 0 0 1 1
use contact_8  contact_8_460
timestamp 1707688321
transform 1 0 7304 0 1 37127
box 0 0 1 1
use contact_8  contact_8_461
timestamp 1707688321
transform 1 0 7304 0 1 36732
box 0 0 1 1
use contact_8  contact_8_462
timestamp 1707688321
transform 1 0 7304 0 1 36337
box 0 0 1 1
use contact_8  contact_8_463
timestamp 1707688321
transform 1 0 7304 0 1 35942
box 0 0 1 1
use contact_8  contact_8_464
timestamp 1707688321
transform 1 0 7304 0 1 35547
box 0 0 1 1
use contact_8  contact_8_465
timestamp 1707688321
transform 1 0 7304 0 1 35152
box 0 0 1 1
use contact_8  contact_8_466
timestamp 1707688321
transform 1 0 7032 0 1 35547
box 0 0 1 1
use contact_8  contact_8_467
timestamp 1707688321
transform 1 0 7032 0 1 35152
box 0 0 1 1
use contact_8  contact_8_468
timestamp 1707688321
transform 1 0 7032 0 1 37522
box 0 0 1 1
use contact_8  contact_8_469
timestamp 1707688321
transform 1 0 7032 0 1 37127
box 0 0 1 1
use contact_8  contact_8_470
timestamp 1707688321
transform 1 0 7032 0 1 36732
box 0 0 1 1
use contact_8  contact_8_471
timestamp 1707688321
transform 1 0 7032 0 1 36337
box 0 0 1 1
use contact_8  contact_8_472
timestamp 1707688321
transform 1 0 5793 0 1 34801
box 0 0 1 1
use contact_8  contact_8_473
timestamp 1707688321
transform 1 0 7304 0 1 34757
box 0 0 1 1
use contact_8  contact_8_474
timestamp 1707688321
transform 1 0 7032 0 1 34757
box 0 0 1 1
use contact_8  contact_8_475
timestamp 1707688321
transform 1 0 5793 0 1 31641
box 0 0 1 1
use contact_8  contact_8_476
timestamp 1707688321
transform 1 0 7032 0 1 31597
box 0 0 1 1
use contact_8  contact_8_477
timestamp 1707688321
transform 1 0 6218 0 1 31583
box 0 0 1 1
use contact_8  contact_8_478
timestamp 1707688321
transform 1 0 6650 0 1 31583
box 0 0 1 1
use contact_8  contact_8_479
timestamp 1707688321
transform 1 0 7304 0 1 31597
box 0 0 1 1
use contact_8  contact_8_480
timestamp 1707688321
transform 1 0 6650 0 1 39915
box 0 0 1 1
use contact_8  contact_8_481
timestamp 1707688321
transform 1 0 6650 0 1 38693
box 0 0 1 1
use contact_8  contact_8_482
timestamp 1707688321
transform 1 0 6650 0 1 39483
box 0 0 1 1
use contact_8  contact_8_483
timestamp 1707688321
transform 1 0 6650 0 1 39125
box 0 0 1 1
use contact_8  contact_8_484
timestamp 1707688321
transform 1 0 6650 0 1 41063
box 0 0 1 1
use contact_8  contact_8_485
timestamp 1707688321
transform 1 0 6650 0 1 40705
box 0 0 1 1
use contact_8  contact_8_486
timestamp 1707688321
transform 1 0 6650 0 1 38335
box 0 0 1 1
use contact_8  contact_8_487
timestamp 1707688321
transform 1 0 6650 0 1 40273
box 0 0 1 1
use contact_8  contact_8_488
timestamp 1707688321
transform 1 0 7032 0 1 40682
box 0 0 1 1
use contact_8  contact_8_489
timestamp 1707688321
transform 1 0 7032 0 1 40287
box 0 0 1 1
use contact_8  contact_8_490
timestamp 1707688321
transform 1 0 7032 0 1 39892
box 0 0 1 1
use contact_8  contact_8_491
timestamp 1707688321
transform 1 0 7032 0 1 39497
box 0 0 1 1
use contact_8  contact_8_492
timestamp 1707688321
transform 1 0 7032 0 1 39102
box 0 0 1 1
use contact_8  contact_8_493
timestamp 1707688321
transform 1 0 7032 0 1 38707
box 0 0 1 1
use contact_8  contact_8_494
timestamp 1707688321
transform 1 0 7032 0 1 38312
box 0 0 1 1
use contact_8  contact_8_495
timestamp 1707688321
transform 1 0 7032 0 1 41077
box 0 0 1 1
use contact_8  contact_8_496
timestamp 1707688321
transform 1 0 7304 0 1 39892
box 0 0 1 1
use contact_8  contact_8_497
timestamp 1707688321
transform 1 0 7304 0 1 41077
box 0 0 1 1
use contact_8  contact_8_498
timestamp 1707688321
transform 1 0 7304 0 1 39102
box 0 0 1 1
use contact_8  contact_8_499
timestamp 1707688321
transform 1 0 7304 0 1 39497
box 0 0 1 1
use contact_8  contact_8_500
timestamp 1707688321
transform 1 0 7304 0 1 40287
box 0 0 1 1
use contact_8  contact_8_501
timestamp 1707688321
transform 1 0 7304 0 1 40682
box 0 0 1 1
use contact_8  contact_8_502
timestamp 1707688321
transform 1 0 7304 0 1 38707
box 0 0 1 1
use contact_8  contact_8_503
timestamp 1707688321
transform 1 0 7304 0 1 38312
box 0 0 1 1
use contact_8  contact_8_504
timestamp 1707688321
transform 1 0 6218 0 1 40705
box 0 0 1 1
use contact_8  contact_8_505
timestamp 1707688321
transform 1 0 5793 0 1 40705
box 0 0 1 1
use contact_8  contact_8_506
timestamp 1707688321
transform 1 0 5793 0 1 40331
box 0 0 1 1
use contact_8  contact_8_507
timestamp 1707688321
transform 1 0 5793 0 1 39915
box 0 0 1 1
use contact_8  contact_8_508
timestamp 1707688321
transform 1 0 5793 0 1 39541
box 0 0 1 1
use contact_8  contact_8_509
timestamp 1707688321
transform 1 0 5793 0 1 39125
box 0 0 1 1
use contact_8  contact_8_510
timestamp 1707688321
transform 1 0 5793 0 1 38751
box 0 0 1 1
use contact_8  contact_8_511
timestamp 1707688321
transform 1 0 5793 0 1 38335
box 0 0 1 1
use contact_8  contact_8_512
timestamp 1707688321
transform 1 0 6218 0 1 39915
box 0 0 1 1
use contact_8  contact_8_513
timestamp 1707688321
transform 1 0 6218 0 1 39125
box 0 0 1 1
use contact_8  contact_8_514
timestamp 1707688321
transform 1 0 6218 0 1 38693
box 0 0 1 1
use contact_8  contact_8_515
timestamp 1707688321
transform 1 0 6218 0 1 38335
box 0 0 1 1
use contact_8  contact_8_516
timestamp 1707688321
transform 1 0 6218 0 1 39483
box 0 0 1 1
use contact_8  contact_8_517
timestamp 1707688321
transform 1 0 6218 0 1 41063
box 0 0 1 1
use contact_8  contact_8_518
timestamp 1707688321
transform 1 0 6218 0 1 40273
box 0 0 1 1
use contact_8  contact_8_519
timestamp 1707688321
transform 1 0 5793 0 1 41495
box 0 0 1 1
use contact_8  contact_8_520
timestamp 1707688321
transform 1 0 5793 0 1 43865
box 0 0 1 1
use contact_8  contact_8_521
timestamp 1707688321
transform 1 0 5793 0 1 43491
box 0 0 1 1
use contact_8  contact_8_522
timestamp 1707688321
transform 1 0 5793 0 1 43075
box 0 0 1 1
use contact_8  contact_8_523
timestamp 1707688321
transform 1 0 5793 0 1 42701
box 0 0 1 1
use contact_8  contact_8_524
timestamp 1707688321
transform 1 0 5793 0 1 42285
box 0 0 1 1
use contact_8  contact_8_525
timestamp 1707688321
transform 1 0 5793 0 1 41911
box 0 0 1 1
use contact_8  contact_8_526
timestamp 1707688321
transform 1 0 6218 0 1 44223
box 0 0 1 1
use contact_8  contact_8_527
timestamp 1707688321
transform 1 0 6218 0 1 43865
box 0 0 1 1
use contact_8  contact_8_528
timestamp 1707688321
transform 1 0 6218 0 1 43433
box 0 0 1 1
use contact_8  contact_8_529
timestamp 1707688321
transform 1 0 6218 0 1 43075
box 0 0 1 1
use contact_8  contact_8_530
timestamp 1707688321
transform 1 0 6218 0 1 42643
box 0 0 1 1
use contact_8  contact_8_531
timestamp 1707688321
transform 1 0 6218 0 1 42285
box 0 0 1 1
use contact_8  contact_8_532
timestamp 1707688321
transform 1 0 6218 0 1 41853
box 0 0 1 1
use contact_8  contact_8_533
timestamp 1707688321
transform 1 0 6218 0 1 41495
box 0 0 1 1
use contact_8  contact_8_534
timestamp 1707688321
transform 1 0 7032 0 1 41472
box 0 0 1 1
use contact_8  contact_8_535
timestamp 1707688321
transform 1 0 6650 0 1 44223
box 0 0 1 1
use contact_8  contact_8_536
timestamp 1707688321
transform 1 0 6650 0 1 43075
box 0 0 1 1
use contact_8  contact_8_537
timestamp 1707688321
transform 1 0 6650 0 1 41495
box 0 0 1 1
use contact_8  contact_8_538
timestamp 1707688321
transform 1 0 6650 0 1 43865
box 0 0 1 1
use contact_8  contact_8_539
timestamp 1707688321
transform 1 0 6650 0 1 42285
box 0 0 1 1
use contact_8  contact_8_540
timestamp 1707688321
transform 1 0 6650 0 1 43433
box 0 0 1 1
use contact_8  contact_8_541
timestamp 1707688321
transform 1 0 6650 0 1 42643
box 0 0 1 1
use contact_8  contact_8_542
timestamp 1707688321
transform 1 0 6650 0 1 41853
box 0 0 1 1
use contact_8  contact_8_543
timestamp 1707688321
transform 1 0 7304 0 1 44237
box 0 0 1 1
use contact_8  contact_8_544
timestamp 1707688321
transform 1 0 7304 0 1 42262
box 0 0 1 1
use contact_8  contact_8_545
timestamp 1707688321
transform 1 0 7304 0 1 43052
box 0 0 1 1
use contact_8  contact_8_546
timestamp 1707688321
transform 1 0 7304 0 1 41867
box 0 0 1 1
use contact_8  contact_8_547
timestamp 1707688321
transform 1 0 7304 0 1 41472
box 0 0 1 1
use contact_8  contact_8_548
timestamp 1707688321
transform 1 0 7304 0 1 43447
box 0 0 1 1
use contact_8  contact_8_549
timestamp 1707688321
transform 1 0 7304 0 1 42657
box 0 0 1 1
use contact_8  contact_8_550
timestamp 1707688321
transform 1 0 7304 0 1 43842
box 0 0 1 1
use contact_8  contact_8_551
timestamp 1707688321
transform 1 0 7032 0 1 44237
box 0 0 1 1
use contact_8  contact_8_552
timestamp 1707688321
transform 1 0 7032 0 1 43842
box 0 0 1 1
use contact_8  contact_8_553
timestamp 1707688321
transform 1 0 7032 0 1 43447
box 0 0 1 1
use contact_8  contact_8_554
timestamp 1707688321
transform 1 0 7032 0 1 43052
box 0 0 1 1
use contact_8  contact_8_555
timestamp 1707688321
transform 1 0 7032 0 1 42657
box 0 0 1 1
use contact_8  contact_8_556
timestamp 1707688321
transform 1 0 7032 0 1 42262
box 0 0 1 1
use contact_8  contact_8_557
timestamp 1707688321
transform 1 0 7032 0 1 41867
box 0 0 1 1
use contact_8  contact_8_558
timestamp 1707688321
transform 1 0 5793 0 1 41121
box 0 0 1 1
use contact_8  contact_8_559
timestamp 1707688321
transform 1 0 7304 0 1 45422
box 0 0 1 1
use contact_8  contact_8_560
timestamp 1707688321
transform 1 0 7304 0 1 47002
box 0 0 1 1
use contact_8  contact_8_561
timestamp 1707688321
transform 1 0 7304 0 1 45817
box 0 0 1 1
use contact_8  contact_8_562
timestamp 1707688321
transform 1 0 7304 0 1 46607
box 0 0 1 1
use contact_8  contact_8_563
timestamp 1707688321
transform 1 0 7304 0 1 45027
box 0 0 1 1
use contact_8  contact_8_564
timestamp 1707688321
transform 1 0 7304 0 1 44632
box 0 0 1 1
use contact_8  contact_8_565
timestamp 1707688321
transform 1 0 6650 0 1 46235
box 0 0 1 1
use contact_8  contact_8_566
timestamp 1707688321
transform 1 0 6650 0 1 45803
box 0 0 1 1
use contact_8  contact_8_567
timestamp 1707688321
transform 1 0 6650 0 1 45445
box 0 0 1 1
use contact_8  contact_8_568
timestamp 1707688321
transform 1 0 6650 0 1 45013
box 0 0 1 1
use contact_8  contact_8_569
timestamp 1707688321
transform 1 0 6650 0 1 44655
box 0 0 1 1
use contact_8  contact_8_570
timestamp 1707688321
transform 1 0 6650 0 1 47383
box 0 0 1 1
use contact_8  contact_8_571
timestamp 1707688321
transform 1 0 6650 0 1 47025
box 0 0 1 1
use contact_8  contact_8_572
timestamp 1707688321
transform 1 0 6650 0 1 46593
box 0 0 1 1
use contact_8  contact_8_573
timestamp 1707688321
transform 1 0 7032 0 1 46212
box 0 0 1 1
use contact_8  contact_8_574
timestamp 1707688321
transform 1 0 7032 0 1 45817
box 0 0 1 1
use contact_8  contact_8_575
timestamp 1707688321
transform 1 0 7032 0 1 45422
box 0 0 1 1
use contact_8  contact_8_576
timestamp 1707688321
transform 1 0 7032 0 1 45027
box 0 0 1 1
use contact_8  contact_8_577
timestamp 1707688321
transform 1 0 7032 0 1 44632
box 0 0 1 1
use contact_8  contact_8_578
timestamp 1707688321
transform 1 0 7032 0 1 47397
box 0 0 1 1
use contact_8  contact_8_579
timestamp 1707688321
transform 1 0 7032 0 1 47002
box 0 0 1 1
use contact_8  contact_8_580
timestamp 1707688321
transform 1 0 7032 0 1 46607
box 0 0 1 1
use contact_8  contact_8_581
timestamp 1707688321
transform 1 0 7304 0 1 46212
box 0 0 1 1
use contact_8  contact_8_582
timestamp 1707688321
transform 1 0 7304 0 1 47397
box 0 0 1 1
use contact_8  contact_8_583
timestamp 1707688321
transform 1 0 6218 0 1 46235
box 0 0 1 1
use contact_8  contact_8_584
timestamp 1707688321
transform 1 0 6218 0 1 45445
box 0 0 1 1
use contact_8  contact_8_585
timestamp 1707688321
transform 1 0 6218 0 1 45803
box 0 0 1 1
use contact_8  contact_8_586
timestamp 1707688321
transform 1 0 6218 0 1 45013
box 0 0 1 1
use contact_8  contact_8_587
timestamp 1707688321
transform 1 0 6218 0 1 47025
box 0 0 1 1
use contact_8  contact_8_588
timestamp 1707688321
transform 1 0 6218 0 1 44655
box 0 0 1 1
use contact_8  contact_8_589
timestamp 1707688321
transform 1 0 6218 0 1 47383
box 0 0 1 1
use contact_8  contact_8_590
timestamp 1707688321
transform 1 0 6218 0 1 46593
box 0 0 1 1
use contact_8  contact_8_591
timestamp 1707688321
transform 1 0 5793 0 1 46651
box 0 0 1 1
use contact_8  contact_8_592
timestamp 1707688321
transform 1 0 5793 0 1 46235
box 0 0 1 1
use contact_8  contact_8_593
timestamp 1707688321
transform 1 0 5793 0 1 45861
box 0 0 1 1
use contact_8  contact_8_594
timestamp 1707688321
transform 1 0 5793 0 1 45445
box 0 0 1 1
use contact_8  contact_8_595
timestamp 1707688321
transform 1 0 5793 0 1 45071
box 0 0 1 1
use contact_8  contact_8_596
timestamp 1707688321
transform 1 0 5793 0 1 44655
box 0 0 1 1
use contact_8  contact_8_597
timestamp 1707688321
transform 1 0 5793 0 1 47025
box 0 0 1 1
use contact_8  contact_8_598
timestamp 1707688321
transform 1 0 5793 0 1 50185
box 0 0 1 1
use contact_8  contact_8_599
timestamp 1707688321
transform 1 0 5793 0 1 49811
box 0 0 1 1
use contact_8  contact_8_600
timestamp 1707688321
transform 1 0 5793 0 1 49395
box 0 0 1 1
use contact_8  contact_8_601
timestamp 1707688321
transform 1 0 5793 0 1 49021
box 0 0 1 1
use contact_8  contact_8_602
timestamp 1707688321
transform 1 0 5793 0 1 48605
box 0 0 1 1
use contact_8  contact_8_603
timestamp 1707688321
transform 1 0 5793 0 1 48231
box 0 0 1 1
use contact_8  contact_8_604
timestamp 1707688321
transform 1 0 5793 0 1 47815
box 0 0 1 1
use contact_8  contact_8_605
timestamp 1707688321
transform 1 0 6218 0 1 48173
box 0 0 1 1
use contact_8  contact_8_606
timestamp 1707688321
transform 1 0 6218 0 1 47815
box 0 0 1 1
use contact_8  contact_8_607
timestamp 1707688321
transform 1 0 6218 0 1 48605
box 0 0 1 1
use contact_8  contact_8_608
timestamp 1707688321
transform 1 0 6218 0 1 50185
box 0 0 1 1
use contact_8  contact_8_609
timestamp 1707688321
transform 1 0 6218 0 1 49753
box 0 0 1 1
use contact_8  contact_8_610
timestamp 1707688321
transform 1 0 6218 0 1 49395
box 0 0 1 1
use contact_8  contact_8_611
timestamp 1707688321
transform 1 0 6218 0 1 48963
box 0 0 1 1
use contact_8  contact_8_612
timestamp 1707688321
transform 1 0 7032 0 1 47792
box 0 0 1 1
use contact_8  contact_8_613
timestamp 1707688321
transform 1 0 6650 0 1 48963
box 0 0 1 1
use contact_8  contact_8_614
timestamp 1707688321
transform 1 0 6650 0 1 50185
box 0 0 1 1
use contact_8  contact_8_615
timestamp 1707688321
transform 1 0 6650 0 1 48173
box 0 0 1 1
use contact_8  contact_8_616
timestamp 1707688321
transform 1 0 6650 0 1 49753
box 0 0 1 1
use contact_8  contact_8_617
timestamp 1707688321
transform 1 0 6650 0 1 48605
box 0 0 1 1
use contact_8  contact_8_618
timestamp 1707688321
transform 1 0 6650 0 1 49395
box 0 0 1 1
use contact_8  contact_8_619
timestamp 1707688321
transform 1 0 6650 0 1 47815
box 0 0 1 1
use contact_8  contact_8_620
timestamp 1707688321
transform 1 0 7304 0 1 47792
box 0 0 1 1
use contact_8  contact_8_621
timestamp 1707688321
transform 1 0 7304 0 1 50162
box 0 0 1 1
use contact_8  contact_8_622
timestamp 1707688321
transform 1 0 7304 0 1 49767
box 0 0 1 1
use contact_8  contact_8_623
timestamp 1707688321
transform 1 0 7304 0 1 49372
box 0 0 1 1
use contact_8  contact_8_624
timestamp 1707688321
transform 1 0 7304 0 1 48977
box 0 0 1 1
use contact_8  contact_8_625
timestamp 1707688321
transform 1 0 7304 0 1 48582
box 0 0 1 1
use contact_8  contact_8_626
timestamp 1707688321
transform 1 0 7304 0 1 48187
box 0 0 1 1
use contact_8  contact_8_627
timestamp 1707688321
transform 1 0 7032 0 1 50162
box 0 0 1 1
use contact_8  contact_8_628
timestamp 1707688321
transform 1 0 7032 0 1 49767
box 0 0 1 1
use contact_8  contact_8_629
timestamp 1707688321
transform 1 0 7032 0 1 49372
box 0 0 1 1
use contact_8  contact_8_630
timestamp 1707688321
transform 1 0 7032 0 1 48977
box 0 0 1 1
use contact_8  contact_8_631
timestamp 1707688321
transform 1 0 7032 0 1 48582
box 0 0 1 1
use contact_8  contact_8_632
timestamp 1707688321
transform 1 0 7032 0 1 48187
box 0 0 1 1
use contact_8  contact_8_633
timestamp 1707688321
transform 1 0 5793 0 1 47441
box 0 0 1 1
use contact_8  contact_8_634
timestamp 1707688321
transform 1 0 5793 0 1 44281
box 0 0 1 1
use contact_8  contact_8_635
timestamp 1707688321
transform 1 0 5793 0 1 37961
box 0 0 1 1
use contact_8  contact_8_636
timestamp 1707688321
transform 1 0 7032 0 1 37917
box 0 0 1 1
use contact_8  contact_8_637
timestamp 1707688321
transform 1 0 7304 0 1 37917
box 0 0 1 1
use contact_8  contact_8_638
timestamp 1707688321
transform 1 0 7032 0 1 25277
box 0 0 1 1
use contact_8  contact_8_639
timestamp 1707688321
transform 1 0 6218 0 1 25263
box 0 0 1 1
use contact_8  contact_8_640
timestamp 1707688321
transform 1 0 6650 0 1 25263
box 0 0 1 1
use contact_8  contact_8_641
timestamp 1707688321
transform 1 0 7304 0 1 25277
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1707688321
transform 1 0 7303 0 1 2362
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1707688321
transform 1 0 7303 0 1 1572
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1707688321
transform 1 0 7303 0 1 2757
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1707688321
transform 1 0 7303 0 1 782
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1707688321
transform 1 0 7303 0 1 1177
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1707688321
transform 1 0 7303 0 1 1967
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1707688321
transform 1 0 7303 0 1 387
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1707688321
transform 1 0 6649 0 1 2348
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1707688321
transform 1 0 6649 0 1 768
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1707688321
transform 1 0 6649 0 1 2780
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1707688321
transform 1 0 6649 0 1 410
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1707688321
transform 1 0 6649 0 1 1990
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1707688321
transform 1 0 6649 0 1 1558
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1707688321
transform 1 0 6649 0 1 1200
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1707688321
transform 1 0 7031 0 1 2362
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1707688321
transform 1 0 7031 0 1 1967
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1707688321
transform 1 0 7031 0 1 1572
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1707688321
transform 1 0 7031 0 1 1177
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1707688321
transform 1 0 7031 0 1 782
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1707688321
transform 1 0 7031 0 1 387
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1707688321
transform 1 0 7031 0 1 2757
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1707688321
transform 1 0 5792 0 1 2780
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1707688321
transform 1 0 6217 0 1 1558
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1707688321
transform 1 0 6217 0 1 1200
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1707688321
transform 1 0 6217 0 1 768
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1707688321
transform 1 0 6217 0 1 410
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1707688321
transform 1 0 6217 0 1 1990
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1707688321
transform 1 0 6217 0 1 2780
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1707688321
transform 1 0 6217 0 1 2348
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1707688321
transform 1 0 5792 0 1 2406
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1707688321
transform 1 0 5792 0 1 1990
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1707688321
transform 1 0 5792 0 1 1616
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1707688321
transform 1 0 5792 0 1 1200
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1707688321
transform 1 0 5792 0 1 826
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1707688321
transform 1 0 5792 0 1 410
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1707688321
transform 1 0 5792 0 1 5940
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1707688321
transform 1 0 5792 0 1 5566
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1707688321
transform 1 0 5792 0 1 5150
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1707688321
transform 1 0 5792 0 1 4776
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1707688321
transform 1 0 5792 0 1 4360
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1707688321
transform 1 0 5792 0 1 3986
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1707688321
transform 1 0 5792 0 1 3570
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1707688321
transform 1 0 5792 0 1 3196
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1707688321
transform 1 0 6217 0 1 5940
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1707688321
transform 1 0 6217 0 1 5508
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1707688321
transform 1 0 6217 0 1 5150
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1707688321
transform 1 0 6217 0 1 4718
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1707688321
transform 1 0 6217 0 1 4360
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1707688321
transform 1 0 6217 0 1 3928
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1707688321
transform 1 0 6217 0 1 3570
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1707688321
transform 1 0 6217 0 1 3138
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1707688321
transform 1 0 6649 0 1 5150
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1707688321
transform 1 0 6649 0 1 3570
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1707688321
transform 1 0 6649 0 1 3928
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1707688321
transform 1 0 6649 0 1 4360
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1707688321
transform 1 0 6649 0 1 5940
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1707688321
transform 1 0 6649 0 1 4718
box 0 0 1 1
use contact_9  contact_9_57
timestamp 1707688321
transform 1 0 6649 0 1 3138
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1707688321
transform 1 0 6649 0 1 5508
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1707688321
transform 1 0 7303 0 1 3942
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1707688321
transform 1 0 7303 0 1 5127
box 0 0 1 1
use contact_9  contact_9_61
timestamp 1707688321
transform 1 0 7303 0 1 4337
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1707688321
transform 1 0 7303 0 1 3547
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1707688321
transform 1 0 7303 0 1 3152
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1707688321
transform 1 0 7303 0 1 4732
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1707688321
transform 1 0 7303 0 1 5917
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1707688321
transform 1 0 7303 0 1 5522
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1707688321
transform 1 0 7031 0 1 4337
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1707688321
transform 1 0 7031 0 1 3942
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1707688321
transform 1 0 7031 0 1 3547
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1707688321
transform 1 0 7031 0 1 3152
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1707688321
transform 1 0 7031 0 1 5917
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1707688321
transform 1 0 7031 0 1 5522
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1707688321
transform 1 0 7031 0 1 5127
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1707688321
transform 1 0 7031 0 1 4732
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1707688321
transform 1 0 7031 0 1 9077
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1707688321
transform 1 0 7303 0 1 6312
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1707688321
transform 1 0 7303 0 1 9077
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1707688321
transform 1 0 7303 0 1 7497
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1707688321
transform 1 0 7303 0 1 8682
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1707688321
transform 1 0 7303 0 1 6707
box 0 0 1 1
use contact_9  contact_9_81
timestamp 1707688321
transform 1 0 7303 0 1 8287
box 0 0 1 1
use contact_9  contact_9_82
timestamp 1707688321
transform 1 0 7303 0 1 7102
box 0 0 1 1
use contact_9  contact_9_83
timestamp 1707688321
transform 1 0 7303 0 1 7892
box 0 0 1 1
use contact_9  contact_9_84
timestamp 1707688321
transform 1 0 6649 0 1 7878
box 0 0 1 1
use contact_9  contact_9_85
timestamp 1707688321
transform 1 0 6649 0 1 7520
box 0 0 1 1
use contact_9  contact_9_86
timestamp 1707688321
transform 1 0 6649 0 1 7088
box 0 0 1 1
use contact_9  contact_9_87
timestamp 1707688321
transform 1 0 6649 0 1 6730
box 0 0 1 1
use contact_9  contact_9_88
timestamp 1707688321
transform 1 0 6649 0 1 9100
box 0 0 1 1
use contact_9  contact_9_89
timestamp 1707688321
transform 1 0 6649 0 1 8668
box 0 0 1 1
use contact_9  contact_9_90
timestamp 1707688321
transform 1 0 6649 0 1 8310
box 0 0 1 1
use contact_9  contact_9_91
timestamp 1707688321
transform 1 0 7031 0 1 8682
box 0 0 1 1
use contact_9  contact_9_92
timestamp 1707688321
transform 1 0 7031 0 1 8287
box 0 0 1 1
use contact_9  contact_9_93
timestamp 1707688321
transform 1 0 7031 0 1 7892
box 0 0 1 1
use contact_9  contact_9_94
timestamp 1707688321
transform 1 0 7031 0 1 7497
box 0 0 1 1
use contact_9  contact_9_95
timestamp 1707688321
transform 1 0 7031 0 1 7102
box 0 0 1 1
use contact_9  contact_9_96
timestamp 1707688321
transform 1 0 7031 0 1 6707
box 0 0 1 1
use contact_9  contact_9_97
timestamp 1707688321
transform 1 0 7031 0 1 6312
box 0 0 1 1
use contact_9  contact_9_98
timestamp 1707688321
transform 1 0 6217 0 1 6730
box 0 0 1 1
use contact_9  contact_9_99
timestamp 1707688321
transform 1 0 6217 0 1 8310
box 0 0 1 1
use contact_9  contact_9_100
timestamp 1707688321
transform 1 0 6217 0 1 7520
box 0 0 1 1
use contact_9  contact_9_101
timestamp 1707688321
transform 1 0 6217 0 1 9100
box 0 0 1 1
use contact_9  contact_9_102
timestamp 1707688321
transform 1 0 6217 0 1 7088
box 0 0 1 1
use contact_9  contact_9_103
timestamp 1707688321
transform 1 0 6217 0 1 7878
box 0 0 1 1
use contact_9  contact_9_104
timestamp 1707688321
transform 1 0 6217 0 1 8668
box 0 0 1 1
use contact_9  contact_9_105
timestamp 1707688321
transform 1 0 5792 0 1 9100
box 0 0 1 1
use contact_9  contact_9_106
timestamp 1707688321
transform 1 0 5792 0 1 8726
box 0 0 1 1
use contact_9  contact_9_107
timestamp 1707688321
transform 1 0 5792 0 1 8310
box 0 0 1 1
use contact_9  contact_9_108
timestamp 1707688321
transform 1 0 5792 0 1 7936
box 0 0 1 1
use contact_9  contact_9_109
timestamp 1707688321
transform 1 0 5792 0 1 7520
box 0 0 1 1
use contact_9  contact_9_110
timestamp 1707688321
transform 1 0 5792 0 1 7146
box 0 0 1 1
use contact_9  contact_9_111
timestamp 1707688321
transform 1 0 5792 0 1 6730
box 0 0 1 1
use contact_9  contact_9_112
timestamp 1707688321
transform 1 0 5792 0 1 6356
box 0 0 1 1
use contact_9  contact_9_113
timestamp 1707688321
transform 1 0 5792 0 1 12260
box 0 0 1 1
use contact_9  contact_9_114
timestamp 1707688321
transform 1 0 5792 0 1 11886
box 0 0 1 1
use contact_9  contact_9_115
timestamp 1707688321
transform 1 0 5792 0 1 11470
box 0 0 1 1
use contact_9  contact_9_116
timestamp 1707688321
transform 1 0 5792 0 1 11096
box 0 0 1 1
use contact_9  contact_9_117
timestamp 1707688321
transform 1 0 5792 0 1 10680
box 0 0 1 1
use contact_9  contact_9_118
timestamp 1707688321
transform 1 0 5792 0 1 10306
box 0 0 1 1
use contact_9  contact_9_119
timestamp 1707688321
transform 1 0 5792 0 1 9890
box 0 0 1 1
use contact_9  contact_9_120
timestamp 1707688321
transform 1 0 5792 0 1 9516
box 0 0 1 1
use contact_9  contact_9_121
timestamp 1707688321
transform 1 0 6217 0 1 10248
box 0 0 1 1
use contact_9  contact_9_122
timestamp 1707688321
transform 1 0 6217 0 1 9890
box 0 0 1 1
use contact_9  contact_9_123
timestamp 1707688321
transform 1 0 6217 0 1 10680
box 0 0 1 1
use contact_9  contact_9_124
timestamp 1707688321
transform 1 0 6217 0 1 12260
box 0 0 1 1
use contact_9  contact_9_125
timestamp 1707688321
transform 1 0 6217 0 1 11828
box 0 0 1 1
use contact_9  contact_9_126
timestamp 1707688321
transform 1 0 6217 0 1 11470
box 0 0 1 1
use contact_9  contact_9_127
timestamp 1707688321
transform 1 0 6217 0 1 11038
box 0 0 1 1
use contact_9  contact_9_128
timestamp 1707688321
transform 1 0 7031 0 1 9472
box 0 0 1 1
use contact_9  contact_9_129
timestamp 1707688321
transform 1 0 6649 0 1 9890
box 0 0 1 1
use contact_9  contact_9_130
timestamp 1707688321
transform 1 0 6649 0 1 11038
box 0 0 1 1
use contact_9  contact_9_131
timestamp 1707688321
transform 1 0 6649 0 1 12260
box 0 0 1 1
use contact_9  contact_9_132
timestamp 1707688321
transform 1 0 6649 0 1 10248
box 0 0 1 1
use contact_9  contact_9_133
timestamp 1707688321
transform 1 0 6649 0 1 11828
box 0 0 1 1
use contact_9  contact_9_134
timestamp 1707688321
transform 1 0 6649 0 1 10680
box 0 0 1 1
use contact_9  contact_9_135
timestamp 1707688321
transform 1 0 6649 0 1 11470
box 0 0 1 1
use contact_9  contact_9_136
timestamp 1707688321
transform 1 0 7303 0 1 12237
box 0 0 1 1
use contact_9  contact_9_137
timestamp 1707688321
transform 1 0 7303 0 1 11842
box 0 0 1 1
use contact_9  contact_9_138
timestamp 1707688321
transform 1 0 7303 0 1 11447
box 0 0 1 1
use contact_9  contact_9_139
timestamp 1707688321
transform 1 0 7303 0 1 11052
box 0 0 1 1
use contact_9  contact_9_140
timestamp 1707688321
transform 1 0 7303 0 1 10657
box 0 0 1 1
use contact_9  contact_9_141
timestamp 1707688321
transform 1 0 7303 0 1 10262
box 0 0 1 1
use contact_9  contact_9_142
timestamp 1707688321
transform 1 0 7303 0 1 9867
box 0 0 1 1
use contact_9  contact_9_143
timestamp 1707688321
transform 1 0 7303 0 1 9472
box 0 0 1 1
use contact_9  contact_9_144
timestamp 1707688321
transform 1 0 7031 0 1 12237
box 0 0 1 1
use contact_9  contact_9_145
timestamp 1707688321
transform 1 0 7031 0 1 11842
box 0 0 1 1
use contact_9  contact_9_146
timestamp 1707688321
transform 1 0 7031 0 1 11447
box 0 0 1 1
use contact_9  contact_9_147
timestamp 1707688321
transform 1 0 7031 0 1 11052
box 0 0 1 1
use contact_9  contact_9_148
timestamp 1707688321
transform 1 0 7031 0 1 10657
box 0 0 1 1
use contact_9  contact_9_149
timestamp 1707688321
transform 1 0 7031 0 1 10262
box 0 0 1 1
use contact_9  contact_9_150
timestamp 1707688321
transform 1 0 7031 0 1 9867
box 0 0 1 1
use contact_9  contact_9_151
timestamp 1707688321
transform 1 0 6217 0 1 9458
box 0 0 1 1
use contact_9  contact_9_152
timestamp 1707688321
transform 1 0 6649 0 1 9458
box 0 0 1 1
use contact_9  contact_9_153
timestamp 1707688321
transform 1 0 6217 0 1 6298
box 0 0 1 1
use contact_9  contact_9_154
timestamp 1707688321
transform 1 0 6649 0 1 6298
box 0 0 1 1
use contact_9  contact_9_155
timestamp 1707688321
transform 1 0 7303 0 1 14607
box 0 0 1 1
use contact_9  contact_9_156
timestamp 1707688321
transform 1 0 7303 0 1 15002
box 0 0 1 1
use contact_9  contact_9_157
timestamp 1707688321
transform 1 0 7303 0 1 14212
box 0 0 1 1
use contact_9  contact_9_158
timestamp 1707688321
transform 1 0 7303 0 1 13027
box 0 0 1 1
use contact_9  contact_9_159
timestamp 1707688321
transform 1 0 6649 0 1 13408
box 0 0 1 1
use contact_9  contact_9_160
timestamp 1707688321
transform 1 0 6649 0 1 14630
box 0 0 1 1
use contact_9  contact_9_161
timestamp 1707688321
transform 1 0 6649 0 1 15420
box 0 0 1 1
use contact_9  contact_9_162
timestamp 1707688321
transform 1 0 6649 0 1 14198
box 0 0 1 1
use contact_9  contact_9_163
timestamp 1707688321
transform 1 0 6649 0 1 13050
box 0 0 1 1
use contact_9  contact_9_164
timestamp 1707688321
transform 1 0 6649 0 1 13840
box 0 0 1 1
use contact_9  contact_9_165
timestamp 1707688321
transform 1 0 6649 0 1 14988
box 0 0 1 1
use contact_9  contact_9_166
timestamp 1707688321
transform 1 0 7031 0 1 14607
box 0 0 1 1
use contact_9  contact_9_167
timestamp 1707688321
transform 1 0 7031 0 1 13422
box 0 0 1 1
use contact_9  contact_9_168
timestamp 1707688321
transform 1 0 7031 0 1 15397
box 0 0 1 1
use contact_9  contact_9_169
timestamp 1707688321
transform 1 0 7031 0 1 15002
box 0 0 1 1
use contact_9  contact_9_170
timestamp 1707688321
transform 1 0 7031 0 1 13027
box 0 0 1 1
use contact_9  contact_9_171
timestamp 1707688321
transform 1 0 7031 0 1 13817
box 0 0 1 1
use contact_9  contact_9_172
timestamp 1707688321
transform 1 0 7031 0 1 14212
box 0 0 1 1
use contact_9  contact_9_173
timestamp 1707688321
transform 1 0 7303 0 1 13422
box 0 0 1 1
use contact_9  contact_9_174
timestamp 1707688321
transform 1 0 7303 0 1 15397
box 0 0 1 1
use contact_9  contact_9_175
timestamp 1707688321
transform 1 0 7303 0 1 13817
box 0 0 1 1
use contact_9  contact_9_176
timestamp 1707688321
transform 1 0 5792 0 1 13050
box 0 0 1 1
use contact_9  contact_9_177
timestamp 1707688321
transform 1 0 5792 0 1 12676
box 0 0 1 1
use contact_9  contact_9_178
timestamp 1707688321
transform 1 0 5792 0 1 13466
box 0 0 1 1
use contact_9  contact_9_179
timestamp 1707688321
transform 1 0 5792 0 1 15420
box 0 0 1 1
use contact_9  contact_9_180
timestamp 1707688321
transform 1 0 5792 0 1 15046
box 0 0 1 1
use contact_9  contact_9_181
timestamp 1707688321
transform 1 0 5792 0 1 14630
box 0 0 1 1
use contact_9  contact_9_182
timestamp 1707688321
transform 1 0 5792 0 1 14256
box 0 0 1 1
use contact_9  contact_9_183
timestamp 1707688321
transform 1 0 5792 0 1 13840
box 0 0 1 1
use contact_9  contact_9_184
timestamp 1707688321
transform 1 0 6217 0 1 13050
box 0 0 1 1
use contact_9  contact_9_185
timestamp 1707688321
transform 1 0 6217 0 1 15420
box 0 0 1 1
use contact_9  contact_9_186
timestamp 1707688321
transform 1 0 6217 0 1 14988
box 0 0 1 1
use contact_9  contact_9_187
timestamp 1707688321
transform 1 0 6217 0 1 14630
box 0 0 1 1
use contact_9  contact_9_188
timestamp 1707688321
transform 1 0 6217 0 1 14198
box 0 0 1 1
use contact_9  contact_9_189
timestamp 1707688321
transform 1 0 6217 0 1 13840
box 0 0 1 1
use contact_9  contact_9_190
timestamp 1707688321
transform 1 0 6217 0 1 13408
box 0 0 1 1
use contact_9  contact_9_191
timestamp 1707688321
transform 1 0 5792 0 1 18580
box 0 0 1 1
use contact_9  contact_9_192
timestamp 1707688321
transform 1 0 5792 0 1 18206
box 0 0 1 1
use contact_9  contact_9_193
timestamp 1707688321
transform 1 0 5792 0 1 17790
box 0 0 1 1
use contact_9  contact_9_194
timestamp 1707688321
transform 1 0 5792 0 1 17416
box 0 0 1 1
use contact_9  contact_9_195
timestamp 1707688321
transform 1 0 5792 0 1 17000
box 0 0 1 1
use contact_9  contact_9_196
timestamp 1707688321
transform 1 0 5792 0 1 16626
box 0 0 1 1
use contact_9  contact_9_197
timestamp 1707688321
transform 1 0 5792 0 1 16210
box 0 0 1 1
use contact_9  contact_9_198
timestamp 1707688321
transform 1 0 5792 0 1 15836
box 0 0 1 1
use contact_9  contact_9_199
timestamp 1707688321
transform 1 0 6217 0 1 18580
box 0 0 1 1
use contact_9  contact_9_200
timestamp 1707688321
transform 1 0 6217 0 1 18148
box 0 0 1 1
use contact_9  contact_9_201
timestamp 1707688321
transform 1 0 6217 0 1 17790
box 0 0 1 1
use contact_9  contact_9_202
timestamp 1707688321
transform 1 0 6217 0 1 17358
box 0 0 1 1
use contact_9  contact_9_203
timestamp 1707688321
transform 1 0 6217 0 1 17000
box 0 0 1 1
use contact_9  contact_9_204
timestamp 1707688321
transform 1 0 6217 0 1 16568
box 0 0 1 1
use contact_9  contact_9_205
timestamp 1707688321
transform 1 0 6217 0 1 16210
box 0 0 1 1
use contact_9  contact_9_206
timestamp 1707688321
transform 1 0 7031 0 1 18557
box 0 0 1 1
use contact_9  contact_9_207
timestamp 1707688321
transform 1 0 6649 0 1 16210
box 0 0 1 1
use contact_9  contact_9_208
timestamp 1707688321
transform 1 0 6649 0 1 17000
box 0 0 1 1
use contact_9  contact_9_209
timestamp 1707688321
transform 1 0 6649 0 1 18148
box 0 0 1 1
use contact_9  contact_9_210
timestamp 1707688321
transform 1 0 6649 0 1 17358
box 0 0 1 1
use contact_9  contact_9_211
timestamp 1707688321
transform 1 0 6649 0 1 16568
box 0 0 1 1
use contact_9  contact_9_212
timestamp 1707688321
transform 1 0 6649 0 1 17790
box 0 0 1 1
use contact_9  contact_9_213
timestamp 1707688321
transform 1 0 6649 0 1 18580
box 0 0 1 1
use contact_9  contact_9_214
timestamp 1707688321
transform 1 0 7303 0 1 16582
box 0 0 1 1
use contact_9  contact_9_215
timestamp 1707688321
transform 1 0 7303 0 1 18162
box 0 0 1 1
use contact_9  contact_9_216
timestamp 1707688321
transform 1 0 7303 0 1 16977
box 0 0 1 1
use contact_9  contact_9_217
timestamp 1707688321
transform 1 0 7303 0 1 17767
box 0 0 1 1
use contact_9  contact_9_218
timestamp 1707688321
transform 1 0 7303 0 1 16187
box 0 0 1 1
use contact_9  contact_9_219
timestamp 1707688321
transform 1 0 7303 0 1 17372
box 0 0 1 1
use contact_9  contact_9_220
timestamp 1707688321
transform 1 0 7303 0 1 18557
box 0 0 1 1
use contact_9  contact_9_221
timestamp 1707688321
transform 1 0 7031 0 1 17767
box 0 0 1 1
use contact_9  contact_9_222
timestamp 1707688321
transform 1 0 7031 0 1 17372
box 0 0 1 1
use contact_9  contact_9_223
timestamp 1707688321
transform 1 0 7031 0 1 16977
box 0 0 1 1
use contact_9  contact_9_224
timestamp 1707688321
transform 1 0 7031 0 1 16582
box 0 0 1 1
use contact_9  contact_9_225
timestamp 1707688321
transform 1 0 7031 0 1 16187
box 0 0 1 1
use contact_9  contact_9_226
timestamp 1707688321
transform 1 0 7031 0 1 18162
box 0 0 1 1
use contact_9  contact_9_227
timestamp 1707688321
transform 1 0 6217 0 1 15778
box 0 0 1 1
use contact_9  contact_9_228
timestamp 1707688321
transform 1 0 7031 0 1 15792
box 0 0 1 1
use contact_9  contact_9_229
timestamp 1707688321
transform 1 0 6649 0 1 15778
box 0 0 1 1
use contact_9  contact_9_230
timestamp 1707688321
transform 1 0 7303 0 1 15792
box 0 0 1 1
use contact_9  contact_9_231
timestamp 1707688321
transform 1 0 7031 0 1 21322
box 0 0 1 1
use contact_9  contact_9_232
timestamp 1707688321
transform 1 0 7031 0 1 20927
box 0 0 1 1
use contact_9  contact_9_233
timestamp 1707688321
transform 1 0 7031 0 1 20532
box 0 0 1 1
use contact_9  contact_9_234
timestamp 1707688321
transform 1 0 7031 0 1 20137
box 0 0 1 1
use contact_9  contact_9_235
timestamp 1707688321
transform 1 0 7031 0 1 19742
box 0 0 1 1
use contact_9  contact_9_236
timestamp 1707688321
transform 1 0 7303 0 1 19347
box 0 0 1 1
use contact_9  contact_9_237
timestamp 1707688321
transform 1 0 7303 0 1 20532
box 0 0 1 1
use contact_9  contact_9_238
timestamp 1707688321
transform 1 0 7303 0 1 21322
box 0 0 1 1
use contact_9  contact_9_239
timestamp 1707688321
transform 1 0 7303 0 1 20137
box 0 0 1 1
use contact_9  contact_9_240
timestamp 1707688321
transform 1 0 7303 0 1 21717
box 0 0 1 1
use contact_9  contact_9_241
timestamp 1707688321
transform 1 0 7303 0 1 19742
box 0 0 1 1
use contact_9  contact_9_242
timestamp 1707688321
transform 1 0 7303 0 1 20927
box 0 0 1 1
use contact_9  contact_9_243
timestamp 1707688321
transform 1 0 6649 0 1 20518
box 0 0 1 1
use contact_9  contact_9_244
timestamp 1707688321
transform 1 0 6649 0 1 20160
box 0 0 1 1
use contact_9  contact_9_245
timestamp 1707688321
transform 1 0 6649 0 1 19728
box 0 0 1 1
use contact_9  contact_9_246
timestamp 1707688321
transform 1 0 6649 0 1 19370
box 0 0 1 1
use contact_9  contact_9_247
timestamp 1707688321
transform 1 0 6649 0 1 21740
box 0 0 1 1
use contact_9  contact_9_248
timestamp 1707688321
transform 1 0 6649 0 1 21308
box 0 0 1 1
use contact_9  contact_9_249
timestamp 1707688321
transform 1 0 6649 0 1 20950
box 0 0 1 1
use contact_9  contact_9_250
timestamp 1707688321
transform 1 0 7031 0 1 19347
box 0 0 1 1
use contact_9  contact_9_251
timestamp 1707688321
transform 1 0 7031 0 1 21717
box 0 0 1 1
use contact_9  contact_9_252
timestamp 1707688321
transform 1 0 6217 0 1 20518
box 0 0 1 1
use contact_9  contact_9_253
timestamp 1707688321
transform 1 0 6217 0 1 21740
box 0 0 1 1
use contact_9  contact_9_254
timestamp 1707688321
transform 1 0 6217 0 1 20950
box 0 0 1 1
use contact_9  contact_9_255
timestamp 1707688321
transform 1 0 6217 0 1 20160
box 0 0 1 1
use contact_9  contact_9_256
timestamp 1707688321
transform 1 0 6217 0 1 19370
box 0 0 1 1
use contact_9  contact_9_257
timestamp 1707688321
transform 1 0 6217 0 1 21308
box 0 0 1 1
use contact_9  contact_9_258
timestamp 1707688321
transform 1 0 6217 0 1 19728
box 0 0 1 1
use contact_9  contact_9_259
timestamp 1707688321
transform 1 0 5792 0 1 18996
box 0 0 1 1
use contact_9  contact_9_260
timestamp 1707688321
transform 1 0 5792 0 1 19370
box 0 0 1 1
use contact_9  contact_9_261
timestamp 1707688321
transform 1 0 5792 0 1 20950
box 0 0 1 1
use contact_9  contact_9_262
timestamp 1707688321
transform 1 0 5792 0 1 19786
box 0 0 1 1
use contact_9  contact_9_263
timestamp 1707688321
transform 1 0 5792 0 1 20576
box 0 0 1 1
use contact_9  contact_9_264
timestamp 1707688321
transform 1 0 5792 0 1 21740
box 0 0 1 1
use contact_9  contact_9_265
timestamp 1707688321
transform 1 0 5792 0 1 20160
box 0 0 1 1
use contact_9  contact_9_266
timestamp 1707688321
transform 1 0 5792 0 1 21366
box 0 0 1 1
use contact_9  contact_9_267
timestamp 1707688321
transform 1 0 5792 0 1 22530
box 0 0 1 1
use contact_9  contact_9_268
timestamp 1707688321
transform 1 0 5792 0 1 24900
box 0 0 1 1
use contact_9  contact_9_269
timestamp 1707688321
transform 1 0 5792 0 1 24526
box 0 0 1 1
use contact_9  contact_9_270
timestamp 1707688321
transform 1 0 5792 0 1 24110
box 0 0 1 1
use contact_9  contact_9_271
timestamp 1707688321
transform 1 0 5792 0 1 22156
box 0 0 1 1
use contact_9  contact_9_272
timestamp 1707688321
transform 1 0 5792 0 1 23736
box 0 0 1 1
use contact_9  contact_9_273
timestamp 1707688321
transform 1 0 5792 0 1 23320
box 0 0 1 1
use contact_9  contact_9_274
timestamp 1707688321
transform 1 0 5792 0 1 22946
box 0 0 1 1
use contact_9  contact_9_275
timestamp 1707688321
transform 1 0 6217 0 1 22530
box 0 0 1 1
use contact_9  contact_9_276
timestamp 1707688321
transform 1 0 6217 0 1 22888
box 0 0 1 1
use contact_9  contact_9_277
timestamp 1707688321
transform 1 0 6217 0 1 23678
box 0 0 1 1
use contact_9  contact_9_278
timestamp 1707688321
transform 1 0 6217 0 1 24900
box 0 0 1 1
use contact_9  contact_9_279
timestamp 1707688321
transform 1 0 6217 0 1 23320
box 0 0 1 1
use contact_9  contact_9_280
timestamp 1707688321
transform 1 0 6217 0 1 24110
box 0 0 1 1
use contact_9  contact_9_281
timestamp 1707688321
transform 1 0 6217 0 1 24468
box 0 0 1 1
use contact_9  contact_9_282
timestamp 1707688321
transform 1 0 7031 0 1 22507
box 0 0 1 1
use contact_9  contact_9_283
timestamp 1707688321
transform 1 0 6649 0 1 24110
box 0 0 1 1
use contact_9  contact_9_284
timestamp 1707688321
transform 1 0 6649 0 1 22530
box 0 0 1 1
use contact_9  contact_9_285
timestamp 1707688321
transform 1 0 6649 0 1 23678
box 0 0 1 1
use contact_9  contact_9_286
timestamp 1707688321
transform 1 0 6649 0 1 23320
box 0 0 1 1
use contact_9  contact_9_287
timestamp 1707688321
transform 1 0 6649 0 1 24468
box 0 0 1 1
use contact_9  contact_9_288
timestamp 1707688321
transform 1 0 6649 0 1 22888
box 0 0 1 1
use contact_9  contact_9_289
timestamp 1707688321
transform 1 0 6649 0 1 24900
box 0 0 1 1
use contact_9  contact_9_290
timestamp 1707688321
transform 1 0 7303 0 1 24087
box 0 0 1 1
use contact_9  contact_9_291
timestamp 1707688321
transform 1 0 7303 0 1 23297
box 0 0 1 1
use contact_9  contact_9_292
timestamp 1707688321
transform 1 0 7303 0 1 23692
box 0 0 1 1
use contact_9  contact_9_293
timestamp 1707688321
transform 1 0 7303 0 1 22902
box 0 0 1 1
use contact_9  contact_9_294
timestamp 1707688321
transform 1 0 7303 0 1 22507
box 0 0 1 1
use contact_9  contact_9_295
timestamp 1707688321
transform 1 0 7303 0 1 24877
box 0 0 1 1
use contact_9  contact_9_296
timestamp 1707688321
transform 1 0 7303 0 1 24482
box 0 0 1 1
use contact_9  contact_9_297
timestamp 1707688321
transform 1 0 7031 0 1 24877
box 0 0 1 1
use contact_9  contact_9_298
timestamp 1707688321
transform 1 0 7031 0 1 24482
box 0 0 1 1
use contact_9  contact_9_299
timestamp 1707688321
transform 1 0 7031 0 1 24087
box 0 0 1 1
use contact_9  contact_9_300
timestamp 1707688321
transform 1 0 7031 0 1 23692
box 0 0 1 1
use contact_9  contact_9_301
timestamp 1707688321
transform 1 0 7031 0 1 23297
box 0 0 1 1
use contact_9  contact_9_302
timestamp 1707688321
transform 1 0 7031 0 1 22902
box 0 0 1 1
use contact_9  contact_9_303
timestamp 1707688321
transform 1 0 6217 0 1 22098
box 0 0 1 1
use contact_9  contact_9_304
timestamp 1707688321
transform 1 0 7031 0 1 22112
box 0 0 1 1
use contact_9  contact_9_305
timestamp 1707688321
transform 1 0 6649 0 1 22098
box 0 0 1 1
use contact_9  contact_9_306
timestamp 1707688321
transform 1 0 7303 0 1 22112
box 0 0 1 1
use contact_9  contact_9_307
timestamp 1707688321
transform 1 0 6217 0 1 18938
box 0 0 1 1
use contact_9  contact_9_308
timestamp 1707688321
transform 1 0 6649 0 1 18938
box 0 0 1 1
use contact_9  contact_9_309
timestamp 1707688321
transform 1 0 7303 0 1 18952
box 0 0 1 1
use contact_9  contact_9_310
timestamp 1707688321
transform 1 0 7031 0 1 18952
box 0 0 1 1
use contact_9  contact_9_311
timestamp 1707688321
transform 1 0 6217 0 1 12618
box 0 0 1 1
use contact_9  contact_9_312
timestamp 1707688321
transform 1 0 6649 0 1 12618
box 0 0 1 1
use contact_9  contact_9_313
timestamp 1707688321
transform 1 0 7303 0 1 12632
box 0 0 1 1
use contact_9  contact_9_314
timestamp 1707688321
transform 1 0 7031 0 1 12632
box 0 0 1 1
use contact_9  contact_9_315
timestamp 1707688321
transform 1 0 7303 0 1 27642
box 0 0 1 1
use contact_9  contact_9_316
timestamp 1707688321
transform 1 0 7303 0 1 26062
box 0 0 1 1
use contact_9  contact_9_317
timestamp 1707688321
transform 1 0 7303 0 1 27247
box 0 0 1 1
use contact_9  contact_9_318
timestamp 1707688321
transform 1 0 7303 0 1 25667
box 0 0 1 1
use contact_9  contact_9_319
timestamp 1707688321
transform 1 0 7303 0 1 26457
box 0 0 1 1
use contact_9  contact_9_320
timestamp 1707688321
transform 1 0 7303 0 1 26852
box 0 0 1 1
use contact_9  contact_9_321
timestamp 1707688321
transform 1 0 7303 0 1 28037
box 0 0 1 1
use contact_9  contact_9_322
timestamp 1707688321
transform 1 0 6649 0 1 26048
box 0 0 1 1
use contact_9  contact_9_323
timestamp 1707688321
transform 1 0 6649 0 1 26480
box 0 0 1 1
use contact_9  contact_9_324
timestamp 1707688321
transform 1 0 6649 0 1 27628
box 0 0 1 1
use contact_9  contact_9_325
timestamp 1707688321
transform 1 0 6649 0 1 26838
box 0 0 1 1
use contact_9  contact_9_326
timestamp 1707688321
transform 1 0 6649 0 1 28060
box 0 0 1 1
use contact_9  contact_9_327
timestamp 1707688321
transform 1 0 6649 0 1 27270
box 0 0 1 1
use contact_9  contact_9_328
timestamp 1707688321
transform 1 0 6649 0 1 25690
box 0 0 1 1
use contact_9  contact_9_329
timestamp 1707688321
transform 1 0 7031 0 1 26457
box 0 0 1 1
use contact_9  contact_9_330
timestamp 1707688321
transform 1 0 7031 0 1 26062
box 0 0 1 1
use contact_9  contact_9_331
timestamp 1707688321
transform 1 0 7031 0 1 25667
box 0 0 1 1
use contact_9  contact_9_332
timestamp 1707688321
transform 1 0 7031 0 1 28037
box 0 0 1 1
use contact_9  contact_9_333
timestamp 1707688321
transform 1 0 7031 0 1 27642
box 0 0 1 1
use contact_9  contact_9_334
timestamp 1707688321
transform 1 0 7031 0 1 27247
box 0 0 1 1
use contact_9  contact_9_335
timestamp 1707688321
transform 1 0 7031 0 1 26852
box 0 0 1 1
use contact_9  contact_9_336
timestamp 1707688321
transform 1 0 5792 0 1 28060
box 0 0 1 1
use contact_9  contact_9_337
timestamp 1707688321
transform 1 0 6217 0 1 26480
box 0 0 1 1
use contact_9  contact_9_338
timestamp 1707688321
transform 1 0 6217 0 1 27628
box 0 0 1 1
use contact_9  contact_9_339
timestamp 1707688321
transform 1 0 6217 0 1 26048
box 0 0 1 1
use contact_9  contact_9_340
timestamp 1707688321
transform 1 0 6217 0 1 27270
box 0 0 1 1
use contact_9  contact_9_341
timestamp 1707688321
transform 1 0 6217 0 1 25690
box 0 0 1 1
use contact_9  contact_9_342
timestamp 1707688321
transform 1 0 6217 0 1 28060
box 0 0 1 1
use contact_9  contact_9_343
timestamp 1707688321
transform 1 0 6217 0 1 26838
box 0 0 1 1
use contact_9  contact_9_344
timestamp 1707688321
transform 1 0 5792 0 1 26106
box 0 0 1 1
use contact_9  contact_9_345
timestamp 1707688321
transform 1 0 5792 0 1 25690
box 0 0 1 1
use contact_9  contact_9_346
timestamp 1707688321
transform 1 0 5792 0 1 25316
box 0 0 1 1
use contact_9  contact_9_347
timestamp 1707688321
transform 1 0 5792 0 1 27686
box 0 0 1 1
use contact_9  contact_9_348
timestamp 1707688321
transform 1 0 5792 0 1 27270
box 0 0 1 1
use contact_9  contact_9_349
timestamp 1707688321
transform 1 0 5792 0 1 26896
box 0 0 1 1
use contact_9  contact_9_350
timestamp 1707688321
transform 1 0 5792 0 1 26480
box 0 0 1 1
use contact_9  contact_9_351
timestamp 1707688321
transform 1 0 6217 0 1 28850
box 0 0 1 1
use contact_9  contact_9_352
timestamp 1707688321
transform 1 0 5792 0 1 31220
box 0 0 1 1
use contact_9  contact_9_353
timestamp 1707688321
transform 1 0 5792 0 1 30846
box 0 0 1 1
use contact_9  contact_9_354
timestamp 1707688321
transform 1 0 5792 0 1 30430
box 0 0 1 1
use contact_9  contact_9_355
timestamp 1707688321
transform 1 0 5792 0 1 30056
box 0 0 1 1
use contact_9  contact_9_356
timestamp 1707688321
transform 1 0 5792 0 1 29640
box 0 0 1 1
use contact_9  contact_9_357
timestamp 1707688321
transform 1 0 5792 0 1 29266
box 0 0 1 1
use contact_9  contact_9_358
timestamp 1707688321
transform 1 0 5792 0 1 28850
box 0 0 1 1
use contact_9  contact_9_359
timestamp 1707688321
transform 1 0 6217 0 1 31220
box 0 0 1 1
use contact_9  contact_9_360
timestamp 1707688321
transform 1 0 6217 0 1 30788
box 0 0 1 1
use contact_9  contact_9_361
timestamp 1707688321
transform 1 0 6217 0 1 30430
box 0 0 1 1
use contact_9  contact_9_362
timestamp 1707688321
transform 1 0 6217 0 1 29998
box 0 0 1 1
use contact_9  contact_9_363
timestamp 1707688321
transform 1 0 6217 0 1 29640
box 0 0 1 1
use contact_9  contact_9_364
timestamp 1707688321
transform 1 0 6217 0 1 29208
box 0 0 1 1
use contact_9  contact_9_365
timestamp 1707688321
transform 1 0 6649 0 1 29998
box 0 0 1 1
use contact_9  contact_9_366
timestamp 1707688321
transform 1 0 6649 0 1 31220
box 0 0 1 1
use contact_9  contact_9_367
timestamp 1707688321
transform 1 0 6649 0 1 28850
box 0 0 1 1
use contact_9  contact_9_368
timestamp 1707688321
transform 1 0 6649 0 1 29208
box 0 0 1 1
use contact_9  contact_9_369
timestamp 1707688321
transform 1 0 6649 0 1 29640
box 0 0 1 1
use contact_9  contact_9_370
timestamp 1707688321
transform 1 0 6649 0 1 30430
box 0 0 1 1
use contact_9  contact_9_371
timestamp 1707688321
transform 1 0 6649 0 1 30788
box 0 0 1 1
use contact_9  contact_9_372
timestamp 1707688321
transform 1 0 7303 0 1 28827
box 0 0 1 1
use contact_9  contact_9_373
timestamp 1707688321
transform 1 0 7303 0 1 30802
box 0 0 1 1
use contact_9  contact_9_374
timestamp 1707688321
transform 1 0 7303 0 1 30012
box 0 0 1 1
use contact_9  contact_9_375
timestamp 1707688321
transform 1 0 7303 0 1 31197
box 0 0 1 1
use contact_9  contact_9_376
timestamp 1707688321
transform 1 0 7303 0 1 29617
box 0 0 1 1
use contact_9  contact_9_377
timestamp 1707688321
transform 1 0 7303 0 1 29222
box 0 0 1 1
use contact_9  contact_9_378
timestamp 1707688321
transform 1 0 7303 0 1 30407
box 0 0 1 1
use contact_9  contact_9_379
timestamp 1707688321
transform 1 0 7031 0 1 29222
box 0 0 1 1
use contact_9  contact_9_380
timestamp 1707688321
transform 1 0 7031 0 1 28827
box 0 0 1 1
use contact_9  contact_9_381
timestamp 1707688321
transform 1 0 7031 0 1 31197
box 0 0 1 1
use contact_9  contact_9_382
timestamp 1707688321
transform 1 0 7031 0 1 30802
box 0 0 1 1
use contact_9  contact_9_383
timestamp 1707688321
transform 1 0 7031 0 1 30407
box 0 0 1 1
use contact_9  contact_9_384
timestamp 1707688321
transform 1 0 7031 0 1 30012
box 0 0 1 1
use contact_9  contact_9_385
timestamp 1707688321
transform 1 0 7031 0 1 29617
box 0 0 1 1
use contact_9  contact_9_386
timestamp 1707688321
transform 1 0 6649 0 1 28418
box 0 0 1 1
use contact_9  contact_9_387
timestamp 1707688321
transform 1 0 7303 0 1 28432
box 0 0 1 1
use contact_9  contact_9_388
timestamp 1707688321
transform 1 0 7031 0 1 28432
box 0 0 1 1
use contact_9  contact_9_389
timestamp 1707688321
transform 1 0 6217 0 1 28418
box 0 0 1 1
use contact_9  contact_9_390
timestamp 1707688321
transform 1 0 5792 0 1 28476
box 0 0 1 1
use contact_9  contact_9_391
timestamp 1707688321
transform 1 0 7031 0 1 34357
box 0 0 1 1
use contact_9  contact_9_392
timestamp 1707688321
transform 1 0 7031 0 1 33962
box 0 0 1 1
use contact_9  contact_9_393
timestamp 1707688321
transform 1 0 7031 0 1 33567
box 0 0 1 1
use contact_9  contact_9_394
timestamp 1707688321
transform 1 0 7303 0 1 33172
box 0 0 1 1
use contact_9  contact_9_395
timestamp 1707688321
transform 1 0 7303 0 1 31987
box 0 0 1 1
use contact_9  contact_9_396
timestamp 1707688321
transform 1 0 7303 0 1 32382
box 0 0 1 1
use contact_9  contact_9_397
timestamp 1707688321
transform 1 0 7303 0 1 33567
box 0 0 1 1
use contact_9  contact_9_398
timestamp 1707688321
transform 1 0 7303 0 1 34357
box 0 0 1 1
use contact_9  contact_9_399
timestamp 1707688321
transform 1 0 7303 0 1 32777
box 0 0 1 1
use contact_9  contact_9_400
timestamp 1707688321
transform 1 0 7303 0 1 33962
box 0 0 1 1
use contact_9  contact_9_401
timestamp 1707688321
transform 1 0 6649 0 1 32368
box 0 0 1 1
use contact_9  contact_9_402
timestamp 1707688321
transform 1 0 6649 0 1 34380
box 0 0 1 1
use contact_9  contact_9_403
timestamp 1707688321
transform 1 0 6649 0 1 33948
box 0 0 1 1
use contact_9  contact_9_404
timestamp 1707688321
transform 1 0 6649 0 1 32010
box 0 0 1 1
use contact_9  contact_9_405
timestamp 1707688321
transform 1 0 6649 0 1 33590
box 0 0 1 1
use contact_9  contact_9_406
timestamp 1707688321
transform 1 0 6649 0 1 33158
box 0 0 1 1
use contact_9  contact_9_407
timestamp 1707688321
transform 1 0 6649 0 1 32800
box 0 0 1 1
use contact_9  contact_9_408
timestamp 1707688321
transform 1 0 7031 0 1 33172
box 0 0 1 1
use contact_9  contact_9_409
timestamp 1707688321
transform 1 0 7031 0 1 32777
box 0 0 1 1
use contact_9  contact_9_410
timestamp 1707688321
transform 1 0 7031 0 1 32382
box 0 0 1 1
use contact_9  contact_9_411
timestamp 1707688321
transform 1 0 7031 0 1 31987
box 0 0 1 1
use contact_9  contact_9_412
timestamp 1707688321
transform 1 0 6217 0 1 33158
box 0 0 1 1
use contact_9  contact_9_413
timestamp 1707688321
transform 1 0 6217 0 1 32800
box 0 0 1 1
use contact_9  contact_9_414
timestamp 1707688321
transform 1 0 6217 0 1 32368
box 0 0 1 1
use contact_9  contact_9_415
timestamp 1707688321
transform 1 0 6217 0 1 33590
box 0 0 1 1
use contact_9  contact_9_416
timestamp 1707688321
transform 1 0 6217 0 1 33948
box 0 0 1 1
use contact_9  contact_9_417
timestamp 1707688321
transform 1 0 6217 0 1 32010
box 0 0 1 1
use contact_9  contact_9_418
timestamp 1707688321
transform 1 0 6217 0 1 34380
box 0 0 1 1
use contact_9  contact_9_419
timestamp 1707688321
transform 1 0 5792 0 1 32800
box 0 0 1 1
use contact_9  contact_9_420
timestamp 1707688321
transform 1 0 5792 0 1 33216
box 0 0 1 1
use contact_9  contact_9_421
timestamp 1707688321
transform 1 0 5792 0 1 32426
box 0 0 1 1
use contact_9  contact_9_422
timestamp 1707688321
transform 1 0 5792 0 1 33590
box 0 0 1 1
use contact_9  contact_9_423
timestamp 1707688321
transform 1 0 5792 0 1 34006
box 0 0 1 1
use contact_9  contact_9_424
timestamp 1707688321
transform 1 0 5792 0 1 34380
box 0 0 1 1
use contact_9  contact_9_425
timestamp 1707688321
transform 1 0 5792 0 1 32010
box 0 0 1 1
use contact_9  contact_9_426
timestamp 1707688321
transform 1 0 5792 0 1 35170
box 0 0 1 1
use contact_9  contact_9_427
timestamp 1707688321
transform 1 0 5792 0 1 36376
box 0 0 1 1
use contact_9  contact_9_428
timestamp 1707688321
transform 1 0 5792 0 1 37540
box 0 0 1 1
use contact_9  contact_9_429
timestamp 1707688321
transform 1 0 5792 0 1 35586
box 0 0 1 1
use contact_9  contact_9_430
timestamp 1707688321
transform 1 0 5792 0 1 37166
box 0 0 1 1
use contact_9  contact_9_431
timestamp 1707688321
transform 1 0 5792 0 1 35960
box 0 0 1 1
use contact_9  contact_9_432
timestamp 1707688321
transform 1 0 5792 0 1 36750
box 0 0 1 1
use contact_9  contact_9_433
timestamp 1707688321
transform 1 0 6217 0 1 37898
box 0 0 1 1
use contact_9  contact_9_434
timestamp 1707688321
transform 1 0 6217 0 1 37540
box 0 0 1 1
use contact_9  contact_9_435
timestamp 1707688321
transform 1 0 6217 0 1 37108
box 0 0 1 1
use contact_9  contact_9_436
timestamp 1707688321
transform 1 0 6217 0 1 36750
box 0 0 1 1
use contact_9  contact_9_437
timestamp 1707688321
transform 1 0 6217 0 1 36318
box 0 0 1 1
use contact_9  contact_9_438
timestamp 1707688321
transform 1 0 6217 0 1 35960
box 0 0 1 1
use contact_9  contact_9_439
timestamp 1707688321
transform 1 0 6217 0 1 35528
box 0 0 1 1
use contact_9  contact_9_440
timestamp 1707688321
transform 1 0 6217 0 1 35170
box 0 0 1 1
use contact_9  contact_9_441
timestamp 1707688321
transform 1 0 7031 0 1 35937
box 0 0 1 1
use contact_9  contact_9_442
timestamp 1707688321
transform 1 0 6649 0 1 37898
box 0 0 1 1
use contact_9  contact_9_443
timestamp 1707688321
transform 1 0 6649 0 1 37540
box 0 0 1 1
use contact_9  contact_9_444
timestamp 1707688321
transform 1 0 6649 0 1 35528
box 0 0 1 1
use contact_9  contact_9_445
timestamp 1707688321
transform 1 0 6649 0 1 37108
box 0 0 1 1
use contact_9  contact_9_446
timestamp 1707688321
transform 1 0 6649 0 1 35960
box 0 0 1 1
use contact_9  contact_9_447
timestamp 1707688321
transform 1 0 6649 0 1 36750
box 0 0 1 1
use contact_9  contact_9_448
timestamp 1707688321
transform 1 0 6649 0 1 35170
box 0 0 1 1
use contact_9  contact_9_449
timestamp 1707688321
transform 1 0 6649 0 1 36318
box 0 0 1 1
use contact_9  contact_9_450
timestamp 1707688321
transform 1 0 7303 0 1 37517
box 0 0 1 1
use contact_9  contact_9_451
timestamp 1707688321
transform 1 0 7303 0 1 37122
box 0 0 1 1
use contact_9  contact_9_452
timestamp 1707688321
transform 1 0 7303 0 1 36727
box 0 0 1 1
use contact_9  contact_9_453
timestamp 1707688321
transform 1 0 7303 0 1 36332
box 0 0 1 1
use contact_9  contact_9_454
timestamp 1707688321
transform 1 0 7303 0 1 35937
box 0 0 1 1
use contact_9  contact_9_455
timestamp 1707688321
transform 1 0 7303 0 1 35542
box 0 0 1 1
use contact_9  contact_9_456
timestamp 1707688321
transform 1 0 7303 0 1 35147
box 0 0 1 1
use contact_9  contact_9_457
timestamp 1707688321
transform 1 0 7031 0 1 35542
box 0 0 1 1
use contact_9  contact_9_458
timestamp 1707688321
transform 1 0 7031 0 1 35147
box 0 0 1 1
use contact_9  contact_9_459
timestamp 1707688321
transform 1 0 7031 0 1 37517
box 0 0 1 1
use contact_9  contact_9_460
timestamp 1707688321
transform 1 0 7031 0 1 37122
box 0 0 1 1
use contact_9  contact_9_461
timestamp 1707688321
transform 1 0 7031 0 1 36727
box 0 0 1 1
use contact_9  contact_9_462
timestamp 1707688321
transform 1 0 7031 0 1 36332
box 0 0 1 1
use contact_9  contact_9_463
timestamp 1707688321
transform 1 0 6217 0 1 34738
box 0 0 1 1
use contact_9  contact_9_464
timestamp 1707688321
transform 1 0 5792 0 1 34796
box 0 0 1 1
use contact_9  contact_9_465
timestamp 1707688321
transform 1 0 6649 0 1 34738
box 0 0 1 1
use contact_9  contact_9_466
timestamp 1707688321
transform 1 0 7303 0 1 34752
box 0 0 1 1
use contact_9  contact_9_467
timestamp 1707688321
transform 1 0 7031 0 1 34752
box 0 0 1 1
use contact_9  contact_9_468
timestamp 1707688321
transform 1 0 5792 0 1 31636
box 0 0 1 1
use contact_9  contact_9_469
timestamp 1707688321
transform 1 0 7031 0 1 31592
box 0 0 1 1
use contact_9  contact_9_470
timestamp 1707688321
transform 1 0 6217 0 1 31578
box 0 0 1 1
use contact_9  contact_9_471
timestamp 1707688321
transform 1 0 6649 0 1 31578
box 0 0 1 1
use contact_9  contact_9_472
timestamp 1707688321
transform 1 0 7303 0 1 31592
box 0 0 1 1
use contact_9  contact_9_473
timestamp 1707688321
transform 1 0 6649 0 1 39910
box 0 0 1 1
use contact_9  contact_9_474
timestamp 1707688321
transform 1 0 6649 0 1 38688
box 0 0 1 1
use contact_9  contact_9_475
timestamp 1707688321
transform 1 0 6649 0 1 39478
box 0 0 1 1
use contact_9  contact_9_476
timestamp 1707688321
transform 1 0 6649 0 1 39120
box 0 0 1 1
use contact_9  contact_9_477
timestamp 1707688321
transform 1 0 6649 0 1 41058
box 0 0 1 1
use contact_9  contact_9_478
timestamp 1707688321
transform 1 0 6649 0 1 40700
box 0 0 1 1
use contact_9  contact_9_479
timestamp 1707688321
transform 1 0 6649 0 1 38330
box 0 0 1 1
use contact_9  contact_9_480
timestamp 1707688321
transform 1 0 6649 0 1 40268
box 0 0 1 1
use contact_9  contact_9_481
timestamp 1707688321
transform 1 0 7031 0 1 40677
box 0 0 1 1
use contact_9  contact_9_482
timestamp 1707688321
transform 1 0 7031 0 1 40282
box 0 0 1 1
use contact_9  contact_9_483
timestamp 1707688321
transform 1 0 7031 0 1 39887
box 0 0 1 1
use contact_9  contact_9_484
timestamp 1707688321
transform 1 0 7031 0 1 39492
box 0 0 1 1
use contact_9  contact_9_485
timestamp 1707688321
transform 1 0 7031 0 1 39097
box 0 0 1 1
use contact_9  contact_9_486
timestamp 1707688321
transform 1 0 7031 0 1 38702
box 0 0 1 1
use contact_9  contact_9_487
timestamp 1707688321
transform 1 0 7031 0 1 38307
box 0 0 1 1
use contact_9  contact_9_488
timestamp 1707688321
transform 1 0 7031 0 1 41072
box 0 0 1 1
use contact_9  contact_9_489
timestamp 1707688321
transform 1 0 7303 0 1 39887
box 0 0 1 1
use contact_9  contact_9_490
timestamp 1707688321
transform 1 0 7303 0 1 41072
box 0 0 1 1
use contact_9  contact_9_491
timestamp 1707688321
transform 1 0 7303 0 1 39097
box 0 0 1 1
use contact_9  contact_9_492
timestamp 1707688321
transform 1 0 7303 0 1 39492
box 0 0 1 1
use contact_9  contact_9_493
timestamp 1707688321
transform 1 0 7303 0 1 40282
box 0 0 1 1
use contact_9  contact_9_494
timestamp 1707688321
transform 1 0 7303 0 1 40677
box 0 0 1 1
use contact_9  contact_9_495
timestamp 1707688321
transform 1 0 7303 0 1 38702
box 0 0 1 1
use contact_9  contact_9_496
timestamp 1707688321
transform 1 0 7303 0 1 38307
box 0 0 1 1
use contact_9  contact_9_497
timestamp 1707688321
transform 1 0 6217 0 1 40700
box 0 0 1 1
use contact_9  contact_9_498
timestamp 1707688321
transform 1 0 5792 0 1 40700
box 0 0 1 1
use contact_9  contact_9_499
timestamp 1707688321
transform 1 0 5792 0 1 40326
box 0 0 1 1
use contact_9  contact_9_500
timestamp 1707688321
transform 1 0 5792 0 1 39910
box 0 0 1 1
use contact_9  contact_9_501
timestamp 1707688321
transform 1 0 5792 0 1 39536
box 0 0 1 1
use contact_9  contact_9_502
timestamp 1707688321
transform 1 0 5792 0 1 39120
box 0 0 1 1
use contact_9  contact_9_503
timestamp 1707688321
transform 1 0 5792 0 1 38746
box 0 0 1 1
use contact_9  contact_9_504
timestamp 1707688321
transform 1 0 5792 0 1 38330
box 0 0 1 1
use contact_9  contact_9_505
timestamp 1707688321
transform 1 0 6217 0 1 39910
box 0 0 1 1
use contact_9  contact_9_506
timestamp 1707688321
transform 1 0 6217 0 1 39120
box 0 0 1 1
use contact_9  contact_9_507
timestamp 1707688321
transform 1 0 6217 0 1 38688
box 0 0 1 1
use contact_9  contact_9_508
timestamp 1707688321
transform 1 0 6217 0 1 38330
box 0 0 1 1
use contact_9  contact_9_509
timestamp 1707688321
transform 1 0 6217 0 1 39478
box 0 0 1 1
use contact_9  contact_9_510
timestamp 1707688321
transform 1 0 6217 0 1 41058
box 0 0 1 1
use contact_9  contact_9_511
timestamp 1707688321
transform 1 0 6217 0 1 40268
box 0 0 1 1
use contact_9  contact_9_512
timestamp 1707688321
transform 1 0 5792 0 1 41490
box 0 0 1 1
use contact_9  contact_9_513
timestamp 1707688321
transform 1 0 5792 0 1 43860
box 0 0 1 1
use contact_9  contact_9_514
timestamp 1707688321
transform 1 0 5792 0 1 43486
box 0 0 1 1
use contact_9  contact_9_515
timestamp 1707688321
transform 1 0 5792 0 1 43070
box 0 0 1 1
use contact_9  contact_9_516
timestamp 1707688321
transform 1 0 5792 0 1 42696
box 0 0 1 1
use contact_9  contact_9_517
timestamp 1707688321
transform 1 0 5792 0 1 42280
box 0 0 1 1
use contact_9  contact_9_518
timestamp 1707688321
transform 1 0 5792 0 1 41906
box 0 0 1 1
use contact_9  contact_9_519
timestamp 1707688321
transform 1 0 6217 0 1 44218
box 0 0 1 1
use contact_9  contact_9_520
timestamp 1707688321
transform 1 0 6217 0 1 43860
box 0 0 1 1
use contact_9  contact_9_521
timestamp 1707688321
transform 1 0 6217 0 1 43428
box 0 0 1 1
use contact_9  contact_9_522
timestamp 1707688321
transform 1 0 6217 0 1 43070
box 0 0 1 1
use contact_9  contact_9_523
timestamp 1707688321
transform 1 0 6217 0 1 42638
box 0 0 1 1
use contact_9  contact_9_524
timestamp 1707688321
transform 1 0 6217 0 1 42280
box 0 0 1 1
use contact_9  contact_9_525
timestamp 1707688321
transform 1 0 6217 0 1 41848
box 0 0 1 1
use contact_9  contact_9_526
timestamp 1707688321
transform 1 0 6217 0 1 41490
box 0 0 1 1
use contact_9  contact_9_527
timestamp 1707688321
transform 1 0 7031 0 1 41467
box 0 0 1 1
use contact_9  contact_9_528
timestamp 1707688321
transform 1 0 6649 0 1 44218
box 0 0 1 1
use contact_9  contact_9_529
timestamp 1707688321
transform 1 0 6649 0 1 43070
box 0 0 1 1
use contact_9  contact_9_530
timestamp 1707688321
transform 1 0 6649 0 1 41490
box 0 0 1 1
use contact_9  contact_9_531
timestamp 1707688321
transform 1 0 6649 0 1 43860
box 0 0 1 1
use contact_9  contact_9_532
timestamp 1707688321
transform 1 0 6649 0 1 42280
box 0 0 1 1
use contact_9  contact_9_533
timestamp 1707688321
transform 1 0 6649 0 1 43428
box 0 0 1 1
use contact_9  contact_9_534
timestamp 1707688321
transform 1 0 6649 0 1 42638
box 0 0 1 1
use contact_9  contact_9_535
timestamp 1707688321
transform 1 0 6649 0 1 41848
box 0 0 1 1
use contact_9  contact_9_536
timestamp 1707688321
transform 1 0 7303 0 1 44232
box 0 0 1 1
use contact_9  contact_9_537
timestamp 1707688321
transform 1 0 7303 0 1 42257
box 0 0 1 1
use contact_9  contact_9_538
timestamp 1707688321
transform 1 0 7303 0 1 43047
box 0 0 1 1
use contact_9  contact_9_539
timestamp 1707688321
transform 1 0 7303 0 1 41862
box 0 0 1 1
use contact_9  contact_9_540
timestamp 1707688321
transform 1 0 7303 0 1 41467
box 0 0 1 1
use contact_9  contact_9_541
timestamp 1707688321
transform 1 0 7303 0 1 43442
box 0 0 1 1
use contact_9  contact_9_542
timestamp 1707688321
transform 1 0 7303 0 1 42652
box 0 0 1 1
use contact_9  contact_9_543
timestamp 1707688321
transform 1 0 7303 0 1 43837
box 0 0 1 1
use contact_9  contact_9_544
timestamp 1707688321
transform 1 0 7031 0 1 44232
box 0 0 1 1
use contact_9  contact_9_545
timestamp 1707688321
transform 1 0 7031 0 1 43837
box 0 0 1 1
use contact_9  contact_9_546
timestamp 1707688321
transform 1 0 7031 0 1 43442
box 0 0 1 1
use contact_9  contact_9_547
timestamp 1707688321
transform 1 0 7031 0 1 43047
box 0 0 1 1
use contact_9  contact_9_548
timestamp 1707688321
transform 1 0 7031 0 1 42652
box 0 0 1 1
use contact_9  contact_9_549
timestamp 1707688321
transform 1 0 7031 0 1 42257
box 0 0 1 1
use contact_9  contact_9_550
timestamp 1707688321
transform 1 0 7031 0 1 41862
box 0 0 1 1
use contact_9  contact_9_551
timestamp 1707688321
transform 1 0 5792 0 1 41116
box 0 0 1 1
use contact_9  contact_9_552
timestamp 1707688321
transform 1 0 7303 0 1 45417
box 0 0 1 1
use contact_9  contact_9_553
timestamp 1707688321
transform 1 0 7303 0 1 46997
box 0 0 1 1
use contact_9  contact_9_554
timestamp 1707688321
transform 1 0 7303 0 1 45812
box 0 0 1 1
use contact_9  contact_9_555
timestamp 1707688321
transform 1 0 7303 0 1 46602
box 0 0 1 1
use contact_9  contact_9_556
timestamp 1707688321
transform 1 0 7303 0 1 45022
box 0 0 1 1
use contact_9  contact_9_557
timestamp 1707688321
transform 1 0 7303 0 1 44627
box 0 0 1 1
use contact_9  contact_9_558
timestamp 1707688321
transform 1 0 6649 0 1 46230
box 0 0 1 1
use contact_9  contact_9_559
timestamp 1707688321
transform 1 0 6649 0 1 45798
box 0 0 1 1
use contact_9  contact_9_560
timestamp 1707688321
transform 1 0 6649 0 1 45440
box 0 0 1 1
use contact_9  contact_9_561
timestamp 1707688321
transform 1 0 6649 0 1 45008
box 0 0 1 1
use contact_9  contact_9_562
timestamp 1707688321
transform 1 0 6649 0 1 44650
box 0 0 1 1
use contact_9  contact_9_563
timestamp 1707688321
transform 1 0 6649 0 1 47378
box 0 0 1 1
use contact_9  contact_9_564
timestamp 1707688321
transform 1 0 6649 0 1 47020
box 0 0 1 1
use contact_9  contact_9_565
timestamp 1707688321
transform 1 0 6649 0 1 46588
box 0 0 1 1
use contact_9  contact_9_566
timestamp 1707688321
transform 1 0 7031 0 1 46207
box 0 0 1 1
use contact_9  contact_9_567
timestamp 1707688321
transform 1 0 7031 0 1 45812
box 0 0 1 1
use contact_9  contact_9_568
timestamp 1707688321
transform 1 0 7031 0 1 45417
box 0 0 1 1
use contact_9  contact_9_569
timestamp 1707688321
transform 1 0 7031 0 1 45022
box 0 0 1 1
use contact_9  contact_9_570
timestamp 1707688321
transform 1 0 7031 0 1 44627
box 0 0 1 1
use contact_9  contact_9_571
timestamp 1707688321
transform 1 0 7031 0 1 47392
box 0 0 1 1
use contact_9  contact_9_572
timestamp 1707688321
transform 1 0 7031 0 1 46997
box 0 0 1 1
use contact_9  contact_9_573
timestamp 1707688321
transform 1 0 7031 0 1 46602
box 0 0 1 1
use contact_9  contact_9_574
timestamp 1707688321
transform 1 0 7303 0 1 46207
box 0 0 1 1
use contact_9  contact_9_575
timestamp 1707688321
transform 1 0 7303 0 1 47392
box 0 0 1 1
use contact_9  contact_9_576
timestamp 1707688321
transform 1 0 6217 0 1 46230
box 0 0 1 1
use contact_9  contact_9_577
timestamp 1707688321
transform 1 0 6217 0 1 45440
box 0 0 1 1
use contact_9  contact_9_578
timestamp 1707688321
transform 1 0 6217 0 1 45798
box 0 0 1 1
use contact_9  contact_9_579
timestamp 1707688321
transform 1 0 6217 0 1 45008
box 0 0 1 1
use contact_9  contact_9_580
timestamp 1707688321
transform 1 0 6217 0 1 47020
box 0 0 1 1
use contact_9  contact_9_581
timestamp 1707688321
transform 1 0 6217 0 1 44650
box 0 0 1 1
use contact_9  contact_9_582
timestamp 1707688321
transform 1 0 6217 0 1 47378
box 0 0 1 1
use contact_9  contact_9_583
timestamp 1707688321
transform 1 0 6217 0 1 46588
box 0 0 1 1
use contact_9  contact_9_584
timestamp 1707688321
transform 1 0 5792 0 1 46646
box 0 0 1 1
use contact_9  contact_9_585
timestamp 1707688321
transform 1 0 5792 0 1 46230
box 0 0 1 1
use contact_9  contact_9_586
timestamp 1707688321
transform 1 0 5792 0 1 45856
box 0 0 1 1
use contact_9  contact_9_587
timestamp 1707688321
transform 1 0 5792 0 1 45440
box 0 0 1 1
use contact_9  contact_9_588
timestamp 1707688321
transform 1 0 5792 0 1 45066
box 0 0 1 1
use contact_9  contact_9_589
timestamp 1707688321
transform 1 0 5792 0 1 44650
box 0 0 1 1
use contact_9  contact_9_590
timestamp 1707688321
transform 1 0 5792 0 1 47020
box 0 0 1 1
use contact_9  contact_9_591
timestamp 1707688321
transform 1 0 5792 0 1 50180
box 0 0 1 1
use contact_9  contact_9_592
timestamp 1707688321
transform 1 0 5792 0 1 49806
box 0 0 1 1
use contact_9  contact_9_593
timestamp 1707688321
transform 1 0 5792 0 1 49390
box 0 0 1 1
use contact_9  contact_9_594
timestamp 1707688321
transform 1 0 5792 0 1 49016
box 0 0 1 1
use contact_9  contact_9_595
timestamp 1707688321
transform 1 0 5792 0 1 48600
box 0 0 1 1
use contact_9  contact_9_596
timestamp 1707688321
transform 1 0 5792 0 1 48226
box 0 0 1 1
use contact_9  contact_9_597
timestamp 1707688321
transform 1 0 5792 0 1 47810
box 0 0 1 1
use contact_9  contact_9_598
timestamp 1707688321
transform 1 0 6217 0 1 48168
box 0 0 1 1
use contact_9  contact_9_599
timestamp 1707688321
transform 1 0 6217 0 1 47810
box 0 0 1 1
use contact_9  contact_9_600
timestamp 1707688321
transform 1 0 6217 0 1 48600
box 0 0 1 1
use contact_9  contact_9_601
timestamp 1707688321
transform 1 0 6217 0 1 50180
box 0 0 1 1
use contact_9  contact_9_602
timestamp 1707688321
transform 1 0 6217 0 1 49748
box 0 0 1 1
use contact_9  contact_9_603
timestamp 1707688321
transform 1 0 6217 0 1 49390
box 0 0 1 1
use contact_9  contact_9_604
timestamp 1707688321
transform 1 0 6217 0 1 48958
box 0 0 1 1
use contact_9  contact_9_605
timestamp 1707688321
transform 1 0 7031 0 1 47787
box 0 0 1 1
use contact_9  contact_9_606
timestamp 1707688321
transform 1 0 6649 0 1 48958
box 0 0 1 1
use contact_9  contact_9_607
timestamp 1707688321
transform 1 0 6649 0 1 50180
box 0 0 1 1
use contact_9  contact_9_608
timestamp 1707688321
transform 1 0 6649 0 1 48168
box 0 0 1 1
use contact_9  contact_9_609
timestamp 1707688321
transform 1 0 6649 0 1 49748
box 0 0 1 1
use contact_9  contact_9_610
timestamp 1707688321
transform 1 0 6649 0 1 48600
box 0 0 1 1
use contact_9  contact_9_611
timestamp 1707688321
transform 1 0 6649 0 1 49390
box 0 0 1 1
use contact_9  contact_9_612
timestamp 1707688321
transform 1 0 6649 0 1 47810
box 0 0 1 1
use contact_9  contact_9_613
timestamp 1707688321
transform 1 0 7303 0 1 47787
box 0 0 1 1
use contact_9  contact_9_614
timestamp 1707688321
transform 1 0 7303 0 1 50157
box 0 0 1 1
use contact_9  contact_9_615
timestamp 1707688321
transform 1 0 7303 0 1 49762
box 0 0 1 1
use contact_9  contact_9_616
timestamp 1707688321
transform 1 0 7303 0 1 49367
box 0 0 1 1
use contact_9  contact_9_617
timestamp 1707688321
transform 1 0 7303 0 1 48972
box 0 0 1 1
use contact_9  contact_9_618
timestamp 1707688321
transform 1 0 7303 0 1 48577
box 0 0 1 1
use contact_9  contact_9_619
timestamp 1707688321
transform 1 0 7303 0 1 48182
box 0 0 1 1
use contact_9  contact_9_620
timestamp 1707688321
transform 1 0 7031 0 1 50157
box 0 0 1 1
use contact_9  contact_9_621
timestamp 1707688321
transform 1 0 7031 0 1 49762
box 0 0 1 1
use contact_9  contact_9_622
timestamp 1707688321
transform 1 0 7031 0 1 49367
box 0 0 1 1
use contact_9  contact_9_623
timestamp 1707688321
transform 1 0 7031 0 1 48972
box 0 0 1 1
use contact_9  contact_9_624
timestamp 1707688321
transform 1 0 7031 0 1 48577
box 0 0 1 1
use contact_9  contact_9_625
timestamp 1707688321
transform 1 0 7031 0 1 48182
box 0 0 1 1
use contact_9  contact_9_626
timestamp 1707688321
transform 1 0 5792 0 1 47436
box 0 0 1 1
use contact_9  contact_9_627
timestamp 1707688321
transform 1 0 5792 0 1 44276
box 0 0 1 1
use contact_9  contact_9_628
timestamp 1707688321
transform 1 0 5792 0 1 37956
box 0 0 1 1
use contact_9  contact_9_629
timestamp 1707688321
transform 1 0 7031 0 1 37912
box 0 0 1 1
use contact_9  contact_9_630
timestamp 1707688321
transform 1 0 7303 0 1 37912
box 0 0 1 1
use contact_9  contact_9_631
timestamp 1707688321
transform 1 0 7031 0 1 25272
box 0 0 1 1
use contact_9  contact_9_632
timestamp 1707688321
transform 1 0 6217 0 1 25258
box 0 0 1 1
use contact_9  contact_9_633
timestamp 1707688321
transform 1 0 6649 0 1 25258
box 0 0 1 1
use contact_9  contact_9_634
timestamp 1707688321
transform 1 0 7303 0 1 25272
box 0 0 1 1
use contact_26  contact_26_0
timestamp 1707688321
transform 1 0 4655 0 1 2765
box 0 0 1 1
use contact_26  contact_26_1
timestamp 1707688321
transform 1 0 5135 0 1 5925
box 0 0 1 1
use contact_26  contact_26_2
timestamp 1707688321
transform 1 0 5055 0 1 5530
box 0 0 1 1
use contact_26  contact_26_3
timestamp 1707688321
transform 1 0 4975 0 1 5135
box 0 0 1 1
use contact_26  contact_26_4
timestamp 1707688321
transform 1 0 4895 0 1 4740
box 0 0 1 1
use contact_26  contact_26_5
timestamp 1707688321
transform 1 0 4815 0 1 3555
box 0 0 1 1
use contact_26  contact_26_6
timestamp 1707688321
transform 1 0 4735 0 1 3160
box 0 0 1 1
use contact_26  contact_26_7
timestamp 1707688321
transform 1 0 4575 0 1 2370
box 0 0 1 1
use contact_26  contact_26_8
timestamp 1707688321
transform 1 0 4495 0 1 1185
box 0 0 1 1
use contact_26  contact_26_9
timestamp 1707688321
transform 1 0 4415 0 1 790
box 0 0 1 1
use contact_26  contact_26_10
timestamp 1707688321
transform 1 0 4335 0 1 395
box 0 0 1 1
use contact_26  contact_26_11
timestamp 1707688321
transform 1 0 4255 0 1 0
box 0 0 1 1
use contact_26  contact_26_12
timestamp 1707688321
transform 1 0 5455 0 1 7505
box 0 0 1 1
use contact_26  contact_26_13
timestamp 1707688321
transform 1 0 5375 0 1 7110
box 0 0 1 1
use contact_26  contact_26_14
timestamp 1707688321
transform 1 0 5295 0 1 6715
box 0 0 1 1
use contact_26  contact_26_15
timestamp 1707688321
transform 1 0 5215 0 1 6320
box 0 0 1 1
use contact_27  contact_27_0
timestamp 1707688321
transform 1 0 4336 0 1 3866
box 0 0 1 1
use contact_27  contact_27_1
timestamp 1707688321
transform 1 0 4256 0 1 3238
box 0 0 1 1
use contact_27  contact_27_2
timestamp 1707688321
transform 1 0 4576 0 1 594
box 0 0 1 1
use contact_27  contact_27_3
timestamp 1707688321
transform 1 0 4496 0 1 3076
box 0 0 1 1
use contact_27  contact_27_4
timestamp 1707688321
transform 1 0 4336 0 1 706
box 0 0 1 1
use contact_27  contact_27_5
timestamp 1707688321
transform 1 0 4416 0 1 2448
box 0 0 1 1
use contact_27  contact_27_6
timestamp 1707688321
transform 1 0 4576 0 1 190
box 0 0 1 1
use contact_27  contact_27_7
timestamp 1707688321
transform 1 0 4336 0 1 2286
box 0 0 1 1
use contact_27  contact_27_8
timestamp 1707688321
transform 1 0 4256 0 1 78
box 0 0 1 1
use contact_27  contact_27_9
timestamp 1707688321
transform 1 0 4256 0 1 1658
box 0 0 1 1
use contact_27  contact_27_10
timestamp 1707688321
transform 1 0 4576 0 1 1384
box 0 0 1 1
use contact_27  contact_27_11
timestamp 1707688321
transform 1 0 4656 0 1 2964
box 0 0 1 1
use contact_27  contact_27_12
timestamp 1707688321
transform 1 0 4656 0 1 2560
box 0 0 1 1
use contact_27  contact_27_13
timestamp 1707688321
transform 1 0 4656 0 1 2174
box 0 0 1 1
use contact_27  contact_27_14
timestamp 1707688321
transform 1 0 4656 0 1 1770
box 0 0 1 1
use contact_27  contact_27_15
timestamp 1707688321
transform 1 0 4896 0 1 1294
box 0 0 1 1
use contact_27  contact_27_16
timestamp 1707688321
transform 1 0 4896 0 1 4230
box 0 0 1 1
use contact_27  contact_27_17
timestamp 1707688321
transform 1 0 4736 0 1 4140
box 0 0 1 1
use contact_27  contact_27_18
timestamp 1707688321
transform 1 0 4896 0 1 3664
box 0 0 1 1
use contact_27  contact_27_19
timestamp 1707688321
transform 1 0 4736 0 1 3754
box 0 0 1 1
use contact_27  contact_27_20
timestamp 1707688321
transform 1 0 4896 0 1 3440
box 0 0 1 1
use contact_27  contact_27_21
timestamp 1707688321
transform 1 0 4736 0 1 3350
box 0 0 1 1
use contact_27  contact_27_22
timestamp 1707688321
transform 1 0 4896 0 1 2874
box 0 0 1 1
use contact_27  contact_27_23
timestamp 1707688321
transform 1 0 4896 0 1 1070
box 0 0 1 1
use contact_27  contact_27_24
timestamp 1707688321
transform 1 0 4896 0 1 2650
box 0 0 1 1
use contact_27  contact_27_25
timestamp 1707688321
transform 1 0 4896 0 1 2084
box 0 0 1 1
use contact_27  contact_27_26
timestamp 1707688321
transform 1 0 4896 0 1 280
box 0 0 1 1
use contact_27  contact_27_27
timestamp 1707688321
transform 1 0 4896 0 1 1860
box 0 0 1 1
use contact_27  contact_27_28
timestamp 1707688321
transform 1 0 4896 0 1 6034
box 0 0 1 1
use contact_27  contact_27_29
timestamp 1707688321
transform 1 0 4816 0 1 6124
box 0 0 1 1
use contact_27  contact_27_30
timestamp 1707688321
transform 1 0 4896 0 1 5810
box 0 0 1 1
use contact_27  contact_27_31
timestamp 1707688321
transform 1 0 4816 0 1 5720
box 0 0 1 1
use contact_27  contact_27_32
timestamp 1707688321
transform 1 0 4896 0 1 5244
box 0 0 1 1
use contact_27  contact_27_33
timestamp 1707688321
transform 1 0 4816 0 1 5334
box 0 0 1 1
use contact_27  contact_27_34
timestamp 1707688321
transform 1 0 4896 0 1 504
box 0 0 1 1
use contact_27  contact_27_35
timestamp 1707688321
transform 1 0 4896 0 1 5020
box 0 0 1 1
use contact_27  contact_27_36
timestamp 1707688321
transform 1 0 4816 0 1 4930
box 0 0 1 1
use contact_27  contact_27_37
timestamp 1707688321
transform 1 0 4896 0 1 4454
box 0 0 1 1
use contact_27  contact_27_38
timestamp 1707688321
transform 1 0 4736 0 1 4544
box 0 0 1 1
use contact_27  contact_27_39
timestamp 1707688321
transform 1 0 4496 0 1 1496
box 0 0 1 1
use contact_27  contact_27_40
timestamp 1707688321
transform 1 0 4576 0 1 980
box 0 0 1 1
use contact_27  contact_27_41
timestamp 1707688321
transform 1 0 4416 0 1 868
box 0 0 1 1
use contact_27  contact_27_42
timestamp 1707688321
transform 1 0 4496 0 1 6236
box 0 0 1 1
use contact_27  contact_27_43
timestamp 1707688321
transform 1 0 4416 0 1 5608
box 0 0 1 1
use contact_27  contact_27_44
timestamp 1707688321
transform 1 0 4336 0 1 5446
box 0 0 1 1
use contact_27  contact_27_45
timestamp 1707688321
transform 1 0 4256 0 1 4818
box 0 0 1 1
use contact_27  contact_27_46
timestamp 1707688321
transform 1 0 4496 0 1 4656
box 0 0 1 1
use contact_27  contact_27_47
timestamp 1707688321
transform 1 0 4416 0 1 4028
box 0 0 1 1
use contact_27  contact_27_48
timestamp 1707688321
transform 1 0 4816 0 1 11250
box 0 0 1 1
use contact_27  contact_27_49
timestamp 1707688321
transform 1 0 4976 0 1 10774
box 0 0 1 1
use contact_27  contact_27_50
timestamp 1707688321
transform 1 0 4736 0 1 10864
box 0 0 1 1
use contact_27  contact_27_51
timestamp 1707688321
transform 1 0 4976 0 1 10550
box 0 0 1 1
use contact_27  contact_27_52
timestamp 1707688321
transform 1 0 4736 0 1 10460
box 0 0 1 1
use contact_27  contact_27_53
timestamp 1707688321
transform 1 0 4976 0 1 9984
box 0 0 1 1
use contact_27  contact_27_54
timestamp 1707688321
transform 1 0 4736 0 1 10074
box 0 0 1 1
use contact_27  contact_27_55
timestamp 1707688321
transform 1 0 4976 0 1 9760
box 0 0 1 1
use contact_27  contact_27_56
timestamp 1707688321
transform 1 0 4736 0 1 9670
box 0 0 1 1
use contact_27  contact_27_57
timestamp 1707688321
transform 1 0 4976 0 1 9194
box 0 0 1 1
use contact_27  contact_27_58
timestamp 1707688321
transform 1 0 4976 0 1 8970
box 0 0 1 1
use contact_27  contact_27_59
timestamp 1707688321
transform 1 0 4976 0 1 8404
box 0 0 1 1
use contact_27  contact_27_60
timestamp 1707688321
transform 1 0 4976 0 1 8180
box 0 0 1 1
use contact_27  contact_27_61
timestamp 1707688321
transform 1 0 4976 0 1 7614
box 0 0 1 1
use contact_27  contact_27_62
timestamp 1707688321
transform 1 0 4976 0 1 7390
box 0 0 1 1
use contact_27  contact_27_63
timestamp 1707688321
transform 1 0 4976 0 1 6824
box 0 0 1 1
use contact_27  contact_27_64
timestamp 1707688321
transform 1 0 4656 0 1 9284
box 0 0 1 1
use contact_27  contact_27_65
timestamp 1707688321
transform 1 0 4656 0 1 8880
box 0 0 1 1
use contact_27  contact_27_66
timestamp 1707688321
transform 1 0 4656 0 1 8494
box 0 0 1 1
use contact_27  contact_27_67
timestamp 1707688321
transform 1 0 4656 0 1 8090
box 0 0 1 1
use contact_27  contact_27_68
timestamp 1707688321
transform 1 0 4336 0 1 10186
box 0 0 1 1
use contact_27  contact_27_69
timestamp 1707688321
transform 1 0 4256 0 1 7978
box 0 0 1 1
use contact_27  contact_27_70
timestamp 1707688321
transform 1 0 4256 0 1 11138
box 0 0 1 1
use contact_27  contact_27_71
timestamp 1707688321
transform 1 0 4416 0 1 8768
box 0 0 1 1
use contact_27  contact_27_72
timestamp 1707688321
transform 1 0 4576 0 1 7300
box 0 0 1 1
use contact_27  contact_27_73
timestamp 1707688321
transform 1 0 4416 0 1 7188
box 0 0 1 1
use contact_27  contact_27_74
timestamp 1707688321
transform 1 0 4256 0 1 9558
box 0 0 1 1
use contact_27  contact_27_75
timestamp 1707688321
transform 1 0 4496 0 1 12556
box 0 0 1 1
use contact_27  contact_27_76
timestamp 1707688321
transform 1 0 4496 0 1 10976
box 0 0 1 1
use contact_27  contact_27_77
timestamp 1707688321
transform 1 0 4336 0 1 7026
box 0 0 1 1
use contact_27  contact_27_78
timestamp 1707688321
transform 1 0 4576 0 1 7704
box 0 0 1 1
use contact_27  contact_27_79
timestamp 1707688321
transform 1 0 4336 0 1 8606
box 0 0 1 1
use contact_27  contact_27_80
timestamp 1707688321
transform 1 0 4416 0 1 11928
box 0 0 1 1
use contact_27  contact_27_81
timestamp 1707688321
transform 1 0 4496 0 1 7816
box 0 0 1 1
use contact_27  contact_27_82
timestamp 1707688321
transform 1 0 4416 0 1 10348
box 0 0 1 1
use contact_27  contact_27_83
timestamp 1707688321
transform 1 0 4496 0 1 9396
box 0 0 1 1
use contact_27  contact_27_84
timestamp 1707688321
transform 1 0 4256 0 1 6398
box 0 0 1 1
use contact_27  contact_27_85
timestamp 1707688321
transform 1 0 4336 0 1 11766
box 0 0 1 1
use contact_27  contact_27_86
timestamp 1707688321
transform 1 0 4576 0 1 6510
box 0 0 1 1
use contact_27  contact_27_87
timestamp 1707688321
transform 1 0 4576 0 1 6914
box 0 0 1 1
use contact_27  contact_27_88
timestamp 1707688321
transform 1 0 4976 0 1 6600
box 0 0 1 1
use contact_27  contact_27_89
timestamp 1707688321
transform 1 0 4976 0 1 12354
box 0 0 1 1
use contact_27  contact_27_90
timestamp 1707688321
transform 1 0 4816 0 1 12444
box 0 0 1 1
use contact_27  contact_27_91
timestamp 1707688321
transform 1 0 4976 0 1 12130
box 0 0 1 1
use contact_27  contact_27_92
timestamp 1707688321
transform 1 0 4816 0 1 12040
box 0 0 1 1
use contact_27  contact_27_93
timestamp 1707688321
transform 1 0 4976 0 1 11564
box 0 0 1 1
use contact_27  contact_27_94
timestamp 1707688321
transform 1 0 4816 0 1 11654
box 0 0 1 1
use contact_27  contact_27_95
timestamp 1707688321
transform 1 0 4976 0 1 11340
box 0 0 1 1
use contact_27  contact_27_96
timestamp 1707688321
transform 1 0 0 0 1 194
box 0 0 1 1
use contact_27  contact_27_97
timestamp 1707688321
transform 1 0 480 0 1 5724
box 0 0 1 1
use contact_27  contact_27_98
timestamp 1707688321
transform 1 0 400 0 1 5330
box 0 0 1 1
use contact_27  contact_27_99
timestamp 1707688321
transform 1 0 320 0 1 4934
box 0 0 1 1
use contact_27  contact_27_100
timestamp 1707688321
transform 1 0 240 0 1 2960
box 0 0 1 1
use contact_27  contact_27_101
timestamp 1707688321
transform 1 0 160 0 1 2564
box 0 0 1 1
use contact_27  contact_27_102
timestamp 1707688321
transform 1 0 80 0 1 590
box 0 0 1 1
use contact_27  contact_27_103
timestamp 1707688321
transform 1 0 4736 0 1 15990
box 0 0 1 1
use contact_27  contact_27_104
timestamp 1707688321
transform 1 0 4816 0 1 18764
box 0 0 1 1
use contact_27  contact_27_105
timestamp 1707688321
transform 1 0 4736 0 1 16780
box 0 0 1 1
use contact_27  contact_27_106
timestamp 1707688321
transform 1 0 5056 0 1 17094
box 0 0 1 1
use contact_27  contact_27_107
timestamp 1707688321
transform 1 0 5056 0 1 15514
box 0 0 1 1
use contact_27  contact_27_108
timestamp 1707688321
transform 1 0 5056 0 1 13144
box 0 0 1 1
use contact_27  contact_27_109
timestamp 1707688321
transform 1 0 5056 0 1 13934
box 0 0 1 1
use contact_27  contact_27_110
timestamp 1707688321
transform 1 0 5056 0 1 18450
box 0 0 1 1
use contact_27  contact_27_111
timestamp 1707688321
transform 1 0 5056 0 1 15290
box 0 0 1 1
use contact_27  contact_27_112
timestamp 1707688321
transform 1 0 4816 0 1 18360
box 0 0 1 1
use contact_27  contact_27_113
timestamp 1707688321
transform 1 0 5056 0 1 14724
box 0 0 1 1
use contact_27  contact_27_114
timestamp 1707688321
transform 1 0 4736 0 1 17184
box 0 0 1 1
use contact_27  contact_27_115
timestamp 1707688321
transform 1 0 5056 0 1 16304
box 0 0 1 1
use contact_27  contact_27_116
timestamp 1707688321
transform 1 0 5056 0 1 17884
box 0 0 1 1
use contact_27  contact_27_117
timestamp 1707688321
transform 1 0 4816 0 1 17974
box 0 0 1 1
use contact_27  contact_27_118
timestamp 1707688321
transform 1 0 4736 0 1 16394
box 0 0 1 1
use contact_27  contact_27_119
timestamp 1707688321
transform 1 0 5056 0 1 16080
box 0 0 1 1
use contact_27  contact_27_120
timestamp 1707688321
transform 1 0 5056 0 1 13710
box 0 0 1 1
use contact_27  contact_27_121
timestamp 1707688321
transform 1 0 5056 0 1 16870
box 0 0 1 1
use contact_27  contact_27_122
timestamp 1707688321
transform 1 0 5056 0 1 14500
box 0 0 1 1
use contact_27  contact_27_123
timestamp 1707688321
transform 1 0 5056 0 1 12920
box 0 0 1 1
use contact_27  contact_27_124
timestamp 1707688321
transform 1 0 5056 0 1 17660
box 0 0 1 1
use contact_27  contact_27_125
timestamp 1707688321
transform 1 0 4816 0 1 17570
box 0 0 1 1
use contact_27  contact_27_126
timestamp 1707688321
transform 1 0 5056 0 1 18674
box 0 0 1 1
use contact_27  contact_27_127
timestamp 1707688321
transform 1 0 4416 0 1 16668
box 0 0 1 1
use contact_27  contact_27_128
timestamp 1707688321
transform 1 0 4336 0 1 16506
box 0 0 1 1
use contact_27  contact_27_129
timestamp 1707688321
transform 1 0 4256 0 1 15878
box 0 0 1 1
use contact_27  contact_27_130
timestamp 1707688321
transform 1 0 4336 0 1 13346
box 0 0 1 1
use contact_27  contact_27_131
timestamp 1707688321
transform 1 0 4576 0 1 13620
box 0 0 1 1
use contact_27  contact_27_132
timestamp 1707688321
transform 1 0 4256 0 1 14298
box 0 0 1 1
use contact_27  contact_27_133
timestamp 1707688321
transform 1 0 4336 0 1 14926
box 0 0 1 1
use contact_27  contact_27_134
timestamp 1707688321
transform 1 0 4256 0 1 12718
box 0 0 1 1
use contact_27  contact_27_135
timestamp 1707688321
transform 1 0 4496 0 1 15716
box 0 0 1 1
use contact_27  contact_27_136
timestamp 1707688321
transform 1 0 4496 0 1 14136
box 0 0 1 1
use contact_27  contact_27_137
timestamp 1707688321
transform 1 0 4336 0 1 18086
box 0 0 1 1
use contact_27  contact_27_138
timestamp 1707688321
transform 1 0 4496 0 1 17296
box 0 0 1 1
use contact_27  contact_27_139
timestamp 1707688321
transform 1 0 4416 0 1 13508
box 0 0 1 1
use contact_27  contact_27_140
timestamp 1707688321
transform 1 0 4256 0 1 17458
box 0 0 1 1
use contact_27  contact_27_141
timestamp 1707688321
transform 1 0 4416 0 1 15088
box 0 0 1 1
use contact_27  contact_27_142
timestamp 1707688321
transform 1 0 4576 0 1 12830
box 0 0 1 1
use contact_27  contact_27_143
timestamp 1707688321
transform 1 0 4496 0 1 18876
box 0 0 1 1
use contact_27  contact_27_144
timestamp 1707688321
transform 1 0 4576 0 1 14024
box 0 0 1 1
use contact_27  contact_27_145
timestamp 1707688321
transform 1 0 4576 0 1 13234
box 0 0 1 1
use contact_27  contact_27_146
timestamp 1707688321
transform 1 0 4416 0 1 18248
box 0 0 1 1
use contact_27  contact_27_147
timestamp 1707688321
transform 1 0 4656 0 1 15604
box 0 0 1 1
use contact_27  contact_27_148
timestamp 1707688321
transform 1 0 4656 0 1 15200
box 0 0 1 1
use contact_27  contact_27_149
timestamp 1707688321
transform 1 0 4656 0 1 14410
box 0 0 1 1
use contact_27  contact_27_150
timestamp 1707688321
transform 1 0 4656 0 1 14814
box 0 0 1 1
use contact_27  contact_27_151
timestamp 1707688321
transform 1 0 4256 0 1 23778
box 0 0 1 1
use contact_27  contact_27_152
timestamp 1707688321
transform 1 0 4576 0 1 19940
box 0 0 1 1
use contact_27  contact_27_153
timestamp 1707688321
transform 1 0 4256 0 1 22198
box 0 0 1 1
use contact_27  contact_27_154
timestamp 1707688321
transform 1 0 4496 0 1 25196
box 0 0 1 1
use contact_27  contact_27_155
timestamp 1707688321
transform 1 0 4256 0 1 20618
box 0 0 1 1
use contact_27  contact_27_156
timestamp 1707688321
transform 1 0 4416 0 1 21408
box 0 0 1 1
use contact_27  contact_27_157
timestamp 1707688321
transform 1 0 4336 0 1 24406
box 0 0 1 1
use contact_27  contact_27_158
timestamp 1707688321
transform 1 0 4336 0 1 19666
box 0 0 1 1
use contact_27  contact_27_159
timestamp 1707688321
transform 1 0 4336 0 1 22826
box 0 0 1 1
use contact_27  contact_27_160
timestamp 1707688321
transform 1 0 4416 0 1 19828
box 0 0 1 1
use contact_27  contact_27_161
timestamp 1707688321
transform 1 0 4256 0 1 19038
box 0 0 1 1
use contact_27  contact_27_162
timestamp 1707688321
transform 1 0 4496 0 1 23616
box 0 0 1 1
use contact_27  contact_27_163
timestamp 1707688321
transform 1 0 4416 0 1 22988
box 0 0 1 1
use contact_27  contact_27_164
timestamp 1707688321
transform 1 0 4336 0 1 21246
box 0 0 1 1
use contact_27  contact_27_165
timestamp 1707688321
transform 1 0 4576 0 1 20344
box 0 0 1 1
use contact_27  contact_27_166
timestamp 1707688321
transform 1 0 4496 0 1 22036
box 0 0 1 1
use contact_27  contact_27_167
timestamp 1707688321
transform 1 0 4496 0 1 20456
box 0 0 1 1
use contact_27  contact_27_168
timestamp 1707688321
transform 1 0 4416 0 1 24568
box 0 0 1 1
use contact_27  contact_27_169
timestamp 1707688321
transform 1 0 4576 0 1 19150
box 0 0 1 1
use contact_27  contact_27_170
timestamp 1707688321
transform 1 0 4576 0 1 19554
box 0 0 1 1
use contact_27  contact_27_171
timestamp 1707688321
transform 1 0 5136 0 1 23414
box 0 0 1 1
use contact_27  contact_27_172
timestamp 1707688321
transform 1 0 5136 0 1 22624
box 0 0 1 1
use contact_27  contact_27_173
timestamp 1707688321
transform 1 0 4736 0 1 23504
box 0 0 1 1
use contact_27  contact_27_174
timestamp 1707688321
transform 1 0 5136 0 1 23980
box 0 0 1 1
use contact_27  contact_27_175
timestamp 1707688321
transform 1 0 5136 0 1 24994
box 0 0 1 1
use contact_27  contact_27_176
timestamp 1707688321
transform 1 0 5136 0 1 21610
box 0 0 1 1
use contact_27  contact_27_177
timestamp 1707688321
transform 1 0 4816 0 1 25084
box 0 0 1 1
use contact_27  contact_27_178
timestamp 1707688321
transform 1 0 5136 0 1 22400
box 0 0 1 1
use contact_27  contact_27_179
timestamp 1707688321
transform 1 0 5136 0 1 21044
box 0 0 1 1
use contact_27  contact_27_180
timestamp 1707688321
transform 1 0 4816 0 1 23890
box 0 0 1 1
use contact_27  contact_27_181
timestamp 1707688321
transform 1 0 5136 0 1 23190
box 0 0 1 1
use contact_27  contact_27_182
timestamp 1707688321
transform 1 0 5136 0 1 20820
box 0 0 1 1
use contact_27  contact_27_183
timestamp 1707688321
transform 1 0 4736 0 1 22714
box 0 0 1 1
use contact_27  contact_27_184
timestamp 1707688321
transform 1 0 5136 0 1 20254
box 0 0 1 1
use contact_27  contact_27_185
timestamp 1707688321
transform 1 0 5136 0 1 20030
box 0 0 1 1
use contact_27  contact_27_186
timestamp 1707688321
transform 1 0 5136 0 1 24770
box 0 0 1 1
use contact_27  contact_27_187
timestamp 1707688321
transform 1 0 5136 0 1 19464
box 0 0 1 1
use contact_27  contact_27_188
timestamp 1707688321
transform 1 0 4816 0 1 24680
box 0 0 1 1
use contact_27  contact_27_189
timestamp 1707688321
transform 1 0 5136 0 1 19240
box 0 0 1 1
use contact_27  contact_27_190
timestamp 1707688321
transform 1 0 4736 0 1 23100
box 0 0 1 1
use contact_27  contact_27_191
timestamp 1707688321
transform 1 0 5136 0 1 24204
box 0 0 1 1
use contact_27  contact_27_192
timestamp 1707688321
transform 1 0 4816 0 1 24294
box 0 0 1 1
use contact_27  contact_27_193
timestamp 1707688321
transform 1 0 4736 0 1 22310
box 0 0 1 1
use contact_27  contact_27_194
timestamp 1707688321
transform 1 0 5136 0 1 21834
box 0 0 1 1
use contact_27  contact_27_195
timestamp 1707688321
transform 1 0 4656 0 1 21924
box 0 0 1 1
use contact_27  contact_27_196
timestamp 1707688321
transform 1 0 4656 0 1 21520
box 0 0 1 1
use contact_27  contact_27_197
timestamp 1707688321
transform 1 0 4656 0 1 21134
box 0 0 1 1
use contact_27  contact_27_198
timestamp 1707688321
transform 1 0 4656 0 1 20730
box 0 0 1 1
use contact_27  contact_27_199
timestamp 1707688321
transform 1 0 4816 0 1 31000
box 0 0 1 1
use contact_27  contact_27_200
timestamp 1707688321
transform 1 0 5216 0 1 30524
box 0 0 1 1
use contact_27  contact_27_201
timestamp 1707688321
transform 1 0 4816 0 1 30614
box 0 0 1 1
use contact_27  contact_27_202
timestamp 1707688321
transform 1 0 5216 0 1 25784
box 0 0 1 1
use contact_27  contact_27_203
timestamp 1707688321
transform 1 0 5216 0 1 30300
box 0 0 1 1
use contact_27  contact_27_204
timestamp 1707688321
transform 1 0 4816 0 1 30210
box 0 0 1 1
use contact_27  contact_27_205
timestamp 1707688321
transform 1 0 5216 0 1 29734
box 0 0 1 1
use contact_27  contact_27_206
timestamp 1707688321
transform 1 0 4736 0 1 29824
box 0 0 1 1
use contact_27  contact_27_207
timestamp 1707688321
transform 1 0 5216 0 1 26574
box 0 0 1 1
use contact_27  contact_27_208
timestamp 1707688321
transform 1 0 5216 0 1 29510
box 0 0 1 1
use contact_27  contact_27_209
timestamp 1707688321
transform 1 0 4736 0 1 29420
box 0 0 1 1
use contact_27  contact_27_210
timestamp 1707688321
transform 1 0 5216 0 1 28944
box 0 0 1 1
use contact_27  contact_27_211
timestamp 1707688321
transform 1 0 4736 0 1 29034
box 0 0 1 1
use contact_27  contact_27_212
timestamp 1707688321
transform 1 0 5216 0 1 28720
box 0 0 1 1
use contact_27  contact_27_213
timestamp 1707688321
transform 1 0 4736 0 1 28630
box 0 0 1 1
use contact_27  contact_27_214
timestamp 1707688321
transform 1 0 5216 0 1 28154
box 0 0 1 1
use contact_27  contact_27_215
timestamp 1707688321
transform 1 0 5216 0 1 26350
box 0 0 1 1
use contact_27  contact_27_216
timestamp 1707688321
transform 1 0 5216 0 1 27930
box 0 0 1 1
use contact_27  contact_27_217
timestamp 1707688321
transform 1 0 5216 0 1 27364
box 0 0 1 1
use contact_27  contact_27_218
timestamp 1707688321
transform 1 0 5216 0 1 25560
box 0 0 1 1
use contact_27  contact_27_219
timestamp 1707688321
transform 1 0 5216 0 1 27140
box 0 0 1 1
use contact_27  contact_27_220
timestamp 1707688321
transform 1 0 4496 0 1 29936
box 0 0 1 1
use contact_27  contact_27_221
timestamp 1707688321
transform 1 0 4416 0 1 29308
box 0 0 1 1
use contact_27  contact_27_222
timestamp 1707688321
transform 1 0 4336 0 1 29146
box 0 0 1 1
use contact_27  contact_27_223
timestamp 1707688321
transform 1 0 4256 0 1 28518
box 0 0 1 1
use contact_27  contact_27_224
timestamp 1707688321
transform 1 0 4576 0 1 25874
box 0 0 1 1
use contact_27  contact_27_225
timestamp 1707688321
transform 1 0 4496 0 1 28356
box 0 0 1 1
use contact_27  contact_27_226
timestamp 1707688321
transform 1 0 4336 0 1 25986
box 0 0 1 1
use contact_27  contact_27_227
timestamp 1707688321
transform 1 0 4416 0 1 27728
box 0 0 1 1
use contact_27  contact_27_228
timestamp 1707688321
transform 1 0 4576 0 1 25470
box 0 0 1 1
use contact_27  contact_27_229
timestamp 1707688321
transform 1 0 4336 0 1 27566
box 0 0 1 1
use contact_27  contact_27_230
timestamp 1707688321
transform 1 0 4256 0 1 25358
box 0 0 1 1
use contact_27  contact_27_231
timestamp 1707688321
transform 1 0 4256 0 1 26938
box 0 0 1 1
use contact_27  contact_27_232
timestamp 1707688321
transform 1 0 4576 0 1 26664
box 0 0 1 1
use contact_27  contact_27_233
timestamp 1707688321
transform 1 0 4496 0 1 26776
box 0 0 1 1
use contact_27  contact_27_234
timestamp 1707688321
transform 1 0 4576 0 1 26260
box 0 0 1 1
use contact_27  contact_27_235
timestamp 1707688321
transform 1 0 4416 0 1 26148
box 0 0 1 1
use contact_27  contact_27_236
timestamp 1707688321
transform 1 0 4496 0 1 31516
box 0 0 1 1
use contact_27  contact_27_237
timestamp 1707688321
transform 1 0 4416 0 1 30888
box 0 0 1 1
use contact_27  contact_27_238
timestamp 1707688321
transform 1 0 4336 0 1 30726
box 0 0 1 1
use contact_27  contact_27_239
timestamp 1707688321
transform 1 0 4256 0 1 30098
box 0 0 1 1
use contact_27  contact_27_240
timestamp 1707688321
transform 1 0 4656 0 1 28244
box 0 0 1 1
use contact_27  contact_27_241
timestamp 1707688321
transform 1 0 4656 0 1 27840
box 0 0 1 1
use contact_27  contact_27_242
timestamp 1707688321
transform 1 0 4656 0 1 27454
box 0 0 1 1
use contact_27  contact_27_243
timestamp 1707688321
transform 1 0 4656 0 1 27050
box 0 0 1 1
use contact_27  contact_27_244
timestamp 1707688321
transform 1 0 5216 0 1 31314
box 0 0 1 1
use contact_27  contact_27_245
timestamp 1707688321
transform 1 0 4816 0 1 31404
box 0 0 1 1
use contact_27  contact_27_246
timestamp 1707688321
transform 1 0 5216 0 1 31090
box 0 0 1 1
use contact_27  contact_27_247
timestamp 1707688321
transform 1 0 4496 0 1 33096
box 0 0 1 1
use contact_27  contact_27_248
timestamp 1707688321
transform 1 0 4256 0 1 36418
box 0 0 1 1
use contact_27  contact_27_249
timestamp 1707688321
transform 1 0 4336 0 1 35466
box 0 0 1 1
use contact_27  contact_27_250
timestamp 1707688321
transform 1 0 4416 0 1 37208
box 0 0 1 1
use contact_27  contact_27_251
timestamp 1707688321
transform 1 0 4336 0 1 37046
box 0 0 1 1
use contact_27  contact_27_252
timestamp 1707688321
transform 1 0 4336 0 1 33886
box 0 0 1 1
use contact_27  contact_27_253
timestamp 1707688321
transform 1 0 4576 0 1 32580
box 0 0 1 1
use contact_27  contact_27_254
timestamp 1707688321
transform 1 0 4256 0 1 34838
box 0 0 1 1
use contact_27  contact_27_255
timestamp 1707688321
transform 1 0 4416 0 1 32468
box 0 0 1 1
use contact_27  contact_27_256
timestamp 1707688321
transform 1 0 4576 0 1 31790
box 0 0 1 1
use contact_27  contact_27_257
timestamp 1707688321
transform 1 0 4256 0 1 31678
box 0 0 1 1
use contact_27  contact_27_258
timestamp 1707688321
transform 1 0 4256 0 1 33258
box 0 0 1 1
use contact_27  contact_27_259
timestamp 1707688321
transform 1 0 5296 0 1 35830
box 0 0 1 1
use contact_27  contact_27_260
timestamp 1707688321
transform 1 0 4736 0 1 35740
box 0 0 1 1
use contact_27  contact_27_261
timestamp 1707688321
transform 1 0 5296 0 1 35264
box 0 0 1 1
use contact_27  contact_27_262
timestamp 1707688321
transform 1 0 4736 0 1 35354
box 0 0 1 1
use contact_27  contact_27_263
timestamp 1707688321
transform 1 0 5296 0 1 35040
box 0 0 1 1
use contact_27  contact_27_264
timestamp 1707688321
transform 1 0 4736 0 1 34950
box 0 0 1 1
use contact_27  contact_27_265
timestamp 1707688321
transform 1 0 5296 0 1 34474
box 0 0 1 1
use contact_27  contact_27_266
timestamp 1707688321
transform 1 0 5296 0 1 36620
box 0 0 1 1
use contact_27  contact_27_267
timestamp 1707688321
transform 1 0 5296 0 1 34250
box 0 0 1 1
use contact_27  contact_27_268
timestamp 1707688321
transform 1 0 5296 0 1 33684
box 0 0 1 1
use contact_27  contact_27_269
timestamp 1707688321
transform 1 0 5296 0 1 33460
box 0 0 1 1
use contact_27  contact_27_270
timestamp 1707688321
transform 1 0 4816 0 1 36530
box 0 0 1 1
use contact_27  contact_27_271
timestamp 1707688321
transform 1 0 5296 0 1 32894
box 0 0 1 1
use contact_27  contact_27_272
timestamp 1707688321
transform 1 0 5296 0 1 32670
box 0 0 1 1
use contact_27  contact_27_273
timestamp 1707688321
transform 1 0 5296 0 1 32104
box 0 0 1 1
use contact_27  contact_27_274
timestamp 1707688321
transform 1 0 5296 0 1 31880
box 0 0 1 1
use contact_27  contact_27_275
timestamp 1707688321
transform 1 0 5296 0 1 36054
box 0 0 1 1
use contact_27  contact_27_276
timestamp 1707688321
transform 1 0 4736 0 1 36144
box 0 0 1 1
use contact_27  contact_27_277
timestamp 1707688321
transform 1 0 5296 0 1 37634
box 0 0 1 1
use contact_27  contact_27_278
timestamp 1707688321
transform 1 0 4816 0 1 37724
box 0 0 1 1
use contact_27  contact_27_279
timestamp 1707688321
transform 1 0 5296 0 1 37410
box 0 0 1 1
use contact_27  contact_27_280
timestamp 1707688321
transform 1 0 4816 0 1 37320
box 0 0 1 1
use contact_27  contact_27_281
timestamp 1707688321
transform 1 0 5296 0 1 36844
box 0 0 1 1
use contact_27  contact_27_282
timestamp 1707688321
transform 1 0 4816 0 1 36934
box 0 0 1 1
use contact_27  contact_27_283
timestamp 1707688321
transform 1 0 4656 0 1 34564
box 0 0 1 1
use contact_27  contact_27_284
timestamp 1707688321
transform 1 0 4656 0 1 34160
box 0 0 1 1
use contact_27  contact_27_285
timestamp 1707688321
transform 1 0 4656 0 1 33774
box 0 0 1 1
use contact_27  contact_27_286
timestamp 1707688321
transform 1 0 4656 0 1 33370
box 0 0 1 1
use contact_27  contact_27_287
timestamp 1707688321
transform 1 0 4496 0 1 36256
box 0 0 1 1
use contact_27  contact_27_288
timestamp 1707688321
transform 1 0 4496 0 1 34676
box 0 0 1 1
use contact_27  contact_27_289
timestamp 1707688321
transform 1 0 4496 0 1 37836
box 0 0 1 1
use contact_27  contact_27_290
timestamp 1707688321
transform 1 0 4576 0 1 32194
box 0 0 1 1
use contact_27  contact_27_291
timestamp 1707688321
transform 1 0 4336 0 1 32306
box 0 0 1 1
use contact_27  contact_27_292
timestamp 1707688321
transform 1 0 4416 0 1 35628
box 0 0 1 1
use contact_27  contact_27_293
timestamp 1707688321
transform 1 0 4576 0 1 32984
box 0 0 1 1
use contact_27  contact_27_294
timestamp 1707688321
transform 1 0 4416 0 1 34048
box 0 0 1 1
use contact_27  contact_27_295
timestamp 1707688321
transform 1 0 4816 0 1 44044
box 0 0 1 1
use contact_27  contact_27_296
timestamp 1707688321
transform 1 0 5376 0 1 43730
box 0 0 1 1
use contact_27  contact_27_297
timestamp 1707688321
transform 1 0 4816 0 1 43640
box 0 0 1 1
use contact_27  contact_27_298
timestamp 1707688321
transform 1 0 5376 0 1 41360
box 0 0 1 1
use contact_27  contact_27_299
timestamp 1707688321
transform 1 0 5376 0 1 42374
box 0 0 1 1
use contact_27  contact_27_300
timestamp 1707688321
transform 1 0 5376 0 1 38990
box 0 0 1 1
use contact_27  contact_27_301
timestamp 1707688321
transform 1 0 4736 0 1 42464
box 0 0 1 1
use contact_27  contact_27_302
timestamp 1707688321
transform 1 0 5376 0 1 43164
box 0 0 1 1
use contact_27  contact_27_303
timestamp 1707688321
transform 1 0 5376 0 1 40570
box 0 0 1 1
use contact_27  contact_27_304
timestamp 1707688321
transform 1 0 5376 0 1 43954
box 0 0 1 1
use contact_27  contact_27_305
timestamp 1707688321
transform 1 0 5376 0 1 41584
box 0 0 1 1
use contact_27  contact_27_306
timestamp 1707688321
transform 1 0 4816 0 1 43254
box 0 0 1 1
use contact_27  contact_27_307
timestamp 1707688321
transform 1 0 4736 0 1 41270
box 0 0 1 1
use contact_27  contact_27_308
timestamp 1707688321
transform 1 0 4736 0 1 41674
box 0 0 1 1
use contact_27  contact_27_309
timestamp 1707688321
transform 1 0 5376 0 1 40004
box 0 0 1 1
use contact_27  contact_27_310
timestamp 1707688321
transform 1 0 5376 0 1 39214
box 0 0 1 1
use contact_27  contact_27_311
timestamp 1707688321
transform 1 0 5376 0 1 42940
box 0 0 1 1
use contact_27  contact_27_312
timestamp 1707688321
transform 1 0 5376 0 1 38200
box 0 0 1 1
use contact_27  contact_27_313
timestamp 1707688321
transform 1 0 5376 0 1 39780
box 0 0 1 1
use contact_27  contact_27_314
timestamp 1707688321
transform 1 0 5376 0 1 42150
box 0 0 1 1
use contact_27  contact_27_315
timestamp 1707688321
transform 1 0 4816 0 1 42850
box 0 0 1 1
use contact_27  contact_27_316
timestamp 1707688321
transform 1 0 5376 0 1 40794
box 0 0 1 1
use contact_27  contact_27_317
timestamp 1707688321
transform 1 0 4736 0 1 42060
box 0 0 1 1
use contact_27  contact_27_318
timestamp 1707688321
transform 1 0 5376 0 1 38424
box 0 0 1 1
use contact_27  contact_27_319
timestamp 1707688321
transform 1 0 4496 0 1 44156
box 0 0 1 1
use contact_27  contact_27_320
timestamp 1707688321
transform 1 0 4416 0 1 41948
box 0 0 1 1
use contact_27  contact_27_321
timestamp 1707688321
transform 1 0 4416 0 1 43528
box 0 0 1 1
use contact_27  contact_27_322
timestamp 1707688321
transform 1 0 4496 0 1 40996
box 0 0 1 1
use contact_27  contact_27_323
timestamp 1707688321
transform 1 0 4576 0 1 38514
box 0 0 1 1
use contact_27  contact_27_324
timestamp 1707688321
transform 1 0 4336 0 1 41786
box 0 0 1 1
use contact_27  contact_27_325
timestamp 1707688321
transform 1 0 4256 0 1 41158
box 0 0 1 1
use contact_27  contact_27_326
timestamp 1707688321
transform 1 0 4416 0 1 40368
box 0 0 1 1
use contact_27  contact_27_327
timestamp 1707688321
transform 1 0 4256 0 1 39578
box 0 0 1 1
use contact_27  contact_27_328
timestamp 1707688321
transform 1 0 4256 0 1 37998
box 0 0 1 1
use contact_27  contact_27_329
timestamp 1707688321
transform 1 0 4336 0 1 40206
box 0 0 1 1
use contact_27  contact_27_330
timestamp 1707688321
transform 1 0 4576 0 1 38110
box 0 0 1 1
use contact_27  contact_27_331
timestamp 1707688321
transform 1 0 4496 0 1 39416
box 0 0 1 1
use contact_27  contact_27_332
timestamp 1707688321
transform 1 0 4256 0 1 42738
box 0 0 1 1
use contact_27  contact_27_333
timestamp 1707688321
transform 1 0 4496 0 1 42576
box 0 0 1 1
use contact_27  contact_27_334
timestamp 1707688321
transform 1 0 4576 0 1 38900
box 0 0 1 1
use contact_27  contact_27_335
timestamp 1707688321
transform 1 0 4336 0 1 38626
box 0 0 1 1
use contact_27  contact_27_336
timestamp 1707688321
transform 1 0 4416 0 1 38788
box 0 0 1 1
use contact_27  contact_27_337
timestamp 1707688321
transform 1 0 4336 0 1 43366
box 0 0 1 1
use contact_27  contact_27_338
timestamp 1707688321
transform 1 0 4576 0 1 39304
box 0 0 1 1
use contact_27  contact_27_339
timestamp 1707688321
transform 1 0 4656 0 1 40480
box 0 0 1 1
use contact_27  contact_27_340
timestamp 1707688321
transform 1 0 4656 0 1 40094
box 0 0 1 1
use contact_27  contact_27_341
timestamp 1707688321
transform 1 0 4656 0 1 39690
box 0 0 1 1
use contact_27  contact_27_342
timestamp 1707688321
transform 1 0 4656 0 1 40884
box 0 0 1 1
use contact_27  contact_27_343
timestamp 1707688321
transform 1 0 4256 0 1 49058
box 0 0 1 1
use contact_27  contact_27_344
timestamp 1707688321
transform 1 0 4576 0 1 44834
box 0 0 1 1
use contact_27  contact_27_345
timestamp 1707688321
transform 1 0 4256 0 1 45898
box 0 0 1 1
use contact_27  contact_27_346
timestamp 1707688321
transform 1 0 4416 0 1 46688
box 0 0 1 1
use contact_27  contact_27_347
timestamp 1707688321
transform 1 0 4576 0 1 45220
box 0 0 1 1
use contact_27  contact_27_348
timestamp 1707688321
transform 1 0 4496 0 1 50476
box 0 0 1 1
use contact_27  contact_27_349
timestamp 1707688321
transform 1 0 4256 0 1 47478
box 0 0 1 1
use contact_27  contact_27_350
timestamp 1707688321
transform 1 0 4496 0 1 48896
box 0 0 1 1
use contact_27  contact_27_351
timestamp 1707688321
transform 1 0 4416 0 1 45108
box 0 0 1 1
use contact_27  contact_27_352
timestamp 1707688321
transform 1 0 4336 0 1 44946
box 0 0 1 1
use contact_27  contact_27_353
timestamp 1707688321
transform 1 0 4416 0 1 49848
box 0 0 1 1
use contact_27  contact_27_354
timestamp 1707688321
transform 1 0 4576 0 1 45624
box 0 0 1 1
use contact_27  contact_27_355
timestamp 1707688321
transform 1 0 4336 0 1 46526
box 0 0 1 1
use contact_27  contact_27_356
timestamp 1707688321
transform 1 0 4416 0 1 48268
box 0 0 1 1
use contact_27  contact_27_357
timestamp 1707688321
transform 1 0 4496 0 1 47316
box 0 0 1 1
use contact_27  contact_27_358
timestamp 1707688321
transform 1 0 4336 0 1 49686
box 0 0 1 1
use contact_27  contact_27_359
timestamp 1707688321
transform 1 0 4496 0 1 45736
box 0 0 1 1
use contact_27  contact_27_360
timestamp 1707688321
transform 1 0 4576 0 1 44430
box 0 0 1 1
use contact_27  contact_27_361
timestamp 1707688321
transform 1 0 4256 0 1 44318
box 0 0 1 1
use contact_27  contact_27_362
timestamp 1707688321
transform 1 0 4336 0 1 48106
box 0 0 1 1
use contact_27  contact_27_363
timestamp 1707688321
transform 1 0 5456 0 1 50274
box 0 0 1 1
use contact_27  contact_27_364
timestamp 1707688321
transform 1 0 4816 0 1 50364
box 0 0 1 1
use contact_27  contact_27_365
timestamp 1707688321
transform 1 0 5456 0 1 50050
box 0 0 1 1
use contact_27  contact_27_366
timestamp 1707688321
transform 1 0 4816 0 1 49960
box 0 0 1 1
use contact_27  contact_27_367
timestamp 1707688321
transform 1 0 5456 0 1 49484
box 0 0 1 1
use contact_27  contact_27_368
timestamp 1707688321
transform 1 0 4816 0 1 49574
box 0 0 1 1
use contact_27  contact_27_369
timestamp 1707688321
transform 1 0 5456 0 1 49260
box 0 0 1 1
use contact_27  contact_27_370
timestamp 1707688321
transform 1 0 4816 0 1 49170
box 0 0 1 1
use contact_27  contact_27_371
timestamp 1707688321
transform 1 0 5456 0 1 48694
box 0 0 1 1
use contact_27  contact_27_372
timestamp 1707688321
transform 1 0 4736 0 1 48784
box 0 0 1 1
use contact_27  contact_27_373
timestamp 1707688321
transform 1 0 5456 0 1 44744
box 0 0 1 1
use contact_27  contact_27_374
timestamp 1707688321
transform 1 0 5456 0 1 48470
box 0 0 1 1
use contact_27  contact_27_375
timestamp 1707688321
transform 1 0 4736 0 1 48380
box 0 0 1 1
use contact_27  contact_27_376
timestamp 1707688321
transform 1 0 5456 0 1 47904
box 0 0 1 1
use contact_27  contact_27_377
timestamp 1707688321
transform 1 0 4736 0 1 47994
box 0 0 1 1
use contact_27  contact_27_378
timestamp 1707688321
transform 1 0 5456 0 1 47680
box 0 0 1 1
use contact_27  contact_27_379
timestamp 1707688321
transform 1 0 4736 0 1 47590
box 0 0 1 1
use contact_27  contact_27_380
timestamp 1707688321
transform 1 0 5456 0 1 47114
box 0 0 1 1
use contact_27  contact_27_381
timestamp 1707688321
transform 1 0 5456 0 1 46890
box 0 0 1 1
use contact_27  contact_27_382
timestamp 1707688321
transform 1 0 5456 0 1 46324
box 0 0 1 1
use contact_27  contact_27_383
timestamp 1707688321
transform 1 0 5456 0 1 44520
box 0 0 1 1
use contact_27  contact_27_384
timestamp 1707688321
transform 1 0 5456 0 1 46100
box 0 0 1 1
use contact_27  contact_27_385
timestamp 1707688321
transform 1 0 5456 0 1 45534
box 0 0 1 1
use contact_27  contact_27_386
timestamp 1707688321
transform 1 0 5456 0 1 45310
box 0 0 1 1
use contact_27  contact_27_387
timestamp 1707688321
transform 1 0 4656 0 1 47204
box 0 0 1 1
use contact_27  contact_27_388
timestamp 1707688321
transform 1 0 4656 0 1 46800
box 0 0 1 1
use contact_27  contact_27_389
timestamp 1707688321
transform 1 0 4656 0 1 46414
box 0 0 1 1
use contact_27  contact_27_390
timestamp 1707688321
transform 1 0 4656 0 1 46010
box 0 0 1 1
use contact_28  contact_28_0
timestamp 1707688321
transform 1 0 5664 0 1 877
box 0 0 1 1
use contact_28  contact_28_1
timestamp 1707688321
transform 1 0 5664 0 1 513
box 0 0 1 1
use contact_28  contact_28_2
timestamp 1707688321
transform 1 0 5664 0 1 1079
box 0 0 1 1
use contact_28  contact_28_3
timestamp 1707688321
transform 1 0 5664 0 1 3085
box 0 0 1 1
use contact_28  contact_28_4
timestamp 1707688321
transform 1 0 5664 0 1 1869
box 0 0 1 1
use contact_28  contact_28_5
timestamp 1707688321
transform 1 0 5664 0 1 289
box 0 0 1 1
use contact_28  contact_28_6
timestamp 1707688321
transform 1 0 5664 0 1 2659
box 0 0 1 1
use contact_28  contact_28_7
timestamp 1707688321
transform 1 0 5664 0 1 87
box 0 0 1 1
use contact_28  contact_28_8
timestamp 1707688321
transform 1 0 5664 0 1 715
box 0 0 1 1
use contact_28  contact_28_9
timestamp 1707688321
transform 1 0 5664 0 1 2093
box 0 0 1 1
use contact_28  contact_28_10
timestamp 1707688321
transform 1 0 5664 0 1 2883
box 0 0 1 1
use contact_28  contact_28_11
timestamp 1707688321
transform 1 0 5664 0 1 1505
box 0 0 1 1
use contact_28  contact_28_12
timestamp 1707688321
transform 1 0 5664 0 1 1303
box 0 0 1 1
use contact_28  contact_28_13
timestamp 1707688321
transform 1 0 5664 0 1 2295
box 0 0 1 1
use contact_28  contact_28_14
timestamp 1707688321
transform 1 0 5664 0 1 1667
box 0 0 1 1
use contact_28  contact_28_15
timestamp 1707688321
transform 1 0 5664 0 1 2457
box 0 0 1 1
use contact_28  contact_28_16
timestamp 1707688321
transform 1 0 5664 0 1 6043
box 0 0 1 1
use contact_28  contact_28_17
timestamp 1707688321
transform 1 0 5664 0 1 3449
box 0 0 1 1
use contact_28  contact_28_18
timestamp 1707688321
transform 1 0 5664 0 1 6245
box 0 0 1 1
use contact_28  contact_28_19
timestamp 1707688321
transform 1 0 5664 0 1 5819
box 0 0 1 1
use contact_28  contact_28_20
timestamp 1707688321
transform 1 0 5664 0 1 3247
box 0 0 1 1
use contact_28  contact_28_21
timestamp 1707688321
transform 1 0 5664 0 1 5617
box 0 0 1 1
use contact_28  contact_28_22
timestamp 1707688321
transform 1 0 5664 0 1 4665
box 0 0 1 1
use contact_28  contact_28_23
timestamp 1707688321
transform 1 0 5664 0 1 5253
box 0 0 1 1
use contact_28  contact_28_24
timestamp 1707688321
transform 1 0 5664 0 1 3875
box 0 0 1 1
use contact_28  contact_28_25
timestamp 1707688321
transform 1 0 5664 0 1 4239
box 0 0 1 1
use contact_28  contact_28_26
timestamp 1707688321
transform 1 0 5664 0 1 5455
box 0 0 1 1
use contact_28  contact_28_27
timestamp 1707688321
transform 1 0 5664 0 1 5029
box 0 0 1 1
use contact_28  contact_28_28
timestamp 1707688321
transform 1 0 5664 0 1 3673
box 0 0 1 1
use contact_28  contact_28_29
timestamp 1707688321
transform 1 0 5664 0 1 4827
box 0 0 1 1
use contact_28  contact_28_30
timestamp 1707688321
transform 1 0 5664 0 1 4463
box 0 0 1 1
use contact_28  contact_28_31
timestamp 1707688321
transform 1 0 5664 0 1 4037
box 0 0 1 1
use contact_28  contact_28_32
timestamp 1707688321
transform 1 0 5554 0 1 4149
box 0 0 1 1
use contact_28  contact_28_33
timestamp 1707688321
transform 1 0 5554 0 1 3763
box 0 0 1 1
use contact_28  contact_28_34
timestamp 1707688321
transform 1 0 5554 0 1 1393
box 0 0 1 1
use contact_28  contact_28_35
timestamp 1707688321
transform 1 0 5554 0 1 3359
box 0 0 1 1
use contact_28  contact_28_36
timestamp 1707688321
transform 1 0 5554 0 1 603
box 0 0 1 1
use contact_28  contact_28_37
timestamp 1707688321
transform 1 0 5554 0 1 2973
box 0 0 1 1
use contact_28  contact_28_38
timestamp 1707688321
transform 1 0 5554 0 1 2569
box 0 0 1 1
use contact_28  contact_28_39
timestamp 1707688321
transform 1 0 5554 0 1 989
box 0 0 1 1
use contact_28  contact_28_40
timestamp 1707688321
transform 1 0 5554 0 1 2183
box 0 0 1 1
use contact_28  contact_28_41
timestamp 1707688321
transform 1 0 5554 0 1 199
box 0 0 1 1
use contact_28  contact_28_42
timestamp 1707688321
transform 1 0 5554 0 1 6133
box 0 0 1 1
use contact_28  contact_28_43
timestamp 1707688321
transform 1 0 5554 0 1 5729
box 0 0 1 1
use contact_28  contact_28_44
timestamp 1707688321
transform 1 0 5554 0 1 1779
box 0 0 1 1
use contact_28  contact_28_45
timestamp 1707688321
transform 1 0 5554 0 1 5343
box 0 0 1 1
use contact_28  contact_28_46
timestamp 1707688321
transform 1 0 5554 0 1 4939
box 0 0 1 1
use contact_28  contact_28_47
timestamp 1707688321
transform 1 0 5554 0 1 4553
box 0 0 1 1
use contact_28  contact_28_48
timestamp 1707688321
transform 1 0 5554 0 1 11259
box 0 0 1 1
use contact_28  contact_28_49
timestamp 1707688321
transform 1 0 5554 0 1 10873
box 0 0 1 1
use contact_28  contact_28_50
timestamp 1707688321
transform 1 0 5554 0 1 10469
box 0 0 1 1
use contact_28  contact_28_51
timestamp 1707688321
transform 1 0 5554 0 1 10083
box 0 0 1 1
use contact_28  contact_28_52
timestamp 1707688321
transform 1 0 5554 0 1 9679
box 0 0 1 1
use contact_28  contact_28_53
timestamp 1707688321
transform 1 0 5554 0 1 9293
box 0 0 1 1
use contact_28  contact_28_54
timestamp 1707688321
transform 1 0 5554 0 1 8889
box 0 0 1 1
use contact_28  contact_28_55
timestamp 1707688321
transform 1 0 5554 0 1 6519
box 0 0 1 1
use contact_28  contact_28_56
timestamp 1707688321
transform 1 0 5554 0 1 8503
box 0 0 1 1
use contact_28  contact_28_57
timestamp 1707688321
transform 1 0 5554 0 1 8099
box 0 0 1 1
use contact_28  contact_28_58
timestamp 1707688321
transform 1 0 5554 0 1 7713
box 0 0 1 1
use contact_28  contact_28_59
timestamp 1707688321
transform 1 0 5554 0 1 7309
box 0 0 1 1
use contact_28  contact_28_60
timestamp 1707688321
transform 1 0 5554 0 1 6923
box 0 0 1 1
use contact_28  contact_28_61
timestamp 1707688321
transform 1 0 5554 0 1 12453
box 0 0 1 1
use contact_28  contact_28_62
timestamp 1707688321
transform 1 0 5554 0 1 12049
box 0 0 1 1
use contact_28  contact_28_63
timestamp 1707688321
transform 1 0 5554 0 1 11663
box 0 0 1 1
use contact_28  contact_28_64
timestamp 1707688321
transform 1 0 5664 0 1 7399
box 0 0 1 1
use contact_28  contact_28_65
timestamp 1707688321
transform 1 0 5664 0 1 7197
box 0 0 1 1
use contact_28  contact_28_66
timestamp 1707688321
transform 1 0 5664 0 1 9405
box 0 0 1 1
use contact_28  contact_28_67
timestamp 1707688321
transform 1 0 5664 0 1 8413
box 0 0 1 1
use contact_28  contact_28_68
timestamp 1707688321
transform 1 0 5664 0 1 8615
box 0 0 1 1
use contact_28  contact_28_69
timestamp 1707688321
transform 1 0 5664 0 1 6833
box 0 0 1 1
use contact_28  contact_28_70
timestamp 1707688321
transform 1 0 5664 0 1 9203
box 0 0 1 1
use contact_28  contact_28_71
timestamp 1707688321
transform 1 0 5664 0 1 8189
box 0 0 1 1
use contact_28  contact_28_72
timestamp 1707688321
transform 1 0 5664 0 1 8979
box 0 0 1 1
use contact_28  contact_28_73
timestamp 1707688321
transform 1 0 5664 0 1 7987
box 0 0 1 1
use contact_28  contact_28_74
timestamp 1707688321
transform 1 0 5664 0 1 7623
box 0 0 1 1
use contact_28  contact_28_75
timestamp 1707688321
transform 1 0 5664 0 1 7035
box 0 0 1 1
use contact_28  contact_28_76
timestamp 1707688321
transform 1 0 5664 0 1 6609
box 0 0 1 1
use contact_28  contact_28_77
timestamp 1707688321
transform 1 0 5664 0 1 7825
box 0 0 1 1
use contact_28  contact_28_78
timestamp 1707688321
transform 1 0 5664 0 1 8777
box 0 0 1 1
use contact_28  contact_28_79
timestamp 1707688321
transform 1 0 5664 0 1 6407
box 0 0 1 1
use contact_28  contact_28_80
timestamp 1707688321
transform 1 0 5664 0 1 11349
box 0 0 1 1
use contact_28  contact_28_81
timestamp 1707688321
transform 1 0 5664 0 1 11147
box 0 0 1 1
use contact_28  contact_28_82
timestamp 1707688321
transform 1 0 5664 0 1 10783
box 0 0 1 1
use contact_28  contact_28_83
timestamp 1707688321
transform 1 0 5664 0 1 10985
box 0 0 1 1
use contact_28  contact_28_84
timestamp 1707688321
transform 1 0 5664 0 1 10559
box 0 0 1 1
use contact_28  contact_28_85
timestamp 1707688321
transform 1 0 5664 0 1 11573
box 0 0 1 1
use contact_28  contact_28_86
timestamp 1707688321
transform 1 0 5664 0 1 9993
box 0 0 1 1
use contact_28  contact_28_87
timestamp 1707688321
transform 1 0 5664 0 1 10195
box 0 0 1 1
use contact_28  contact_28_88
timestamp 1707688321
transform 1 0 5664 0 1 11775
box 0 0 1 1
use contact_28  contact_28_89
timestamp 1707688321
transform 1 0 5664 0 1 10357
box 0 0 1 1
use contact_28  contact_28_90
timestamp 1707688321
transform 1 0 5664 0 1 9769
box 0 0 1 1
use contact_28  contact_28_91
timestamp 1707688321
transform 1 0 5664 0 1 9567
box 0 0 1 1
use contact_28  contact_28_92
timestamp 1707688321
transform 1 0 5664 0 1 12363
box 0 0 1 1
use contact_28  contact_28_93
timestamp 1707688321
transform 1 0 5664 0 1 12565
box 0 0 1 1
use contact_28  contact_28_94
timestamp 1707688321
transform 1 0 5664 0 1 12139
box 0 0 1 1
use contact_28  contact_28_95
timestamp 1707688321
transform 1 0 5664 0 1 11937
box 0 0 1 1
use contact_28  contact_28_96
timestamp 1707688321
transform 1 0 5664 0 1 15523
box 0 0 1 1
use contact_28  contact_28_97
timestamp 1707688321
transform 1 0 5664 0 1 15725
box 0 0 1 1
use contact_28  contact_28_98
timestamp 1707688321
transform 1 0 5664 0 1 15299
box 0 0 1 1
use contact_28  contact_28_99
timestamp 1707688321
transform 1 0 5664 0 1 15097
box 0 0 1 1
use contact_28  contact_28_100
timestamp 1707688321
transform 1 0 5664 0 1 14733
box 0 0 1 1
use contact_28  contact_28_101
timestamp 1707688321
transform 1 0 5664 0 1 14935
box 0 0 1 1
use contact_28  contact_28_102
timestamp 1707688321
transform 1 0 5664 0 1 14509
box 0 0 1 1
use contact_28  contact_28_103
timestamp 1707688321
transform 1 0 5664 0 1 14307
box 0 0 1 1
use contact_28  contact_28_104
timestamp 1707688321
transform 1 0 5664 0 1 13943
box 0 0 1 1
use contact_28  contact_28_105
timestamp 1707688321
transform 1 0 5664 0 1 14145
box 0 0 1 1
use contact_28  contact_28_106
timestamp 1707688321
transform 1 0 5664 0 1 13719
box 0 0 1 1
use contact_28  contact_28_107
timestamp 1707688321
transform 1 0 5664 0 1 13517
box 0 0 1 1
use contact_28  contact_28_108
timestamp 1707688321
transform 1 0 5664 0 1 13153
box 0 0 1 1
use contact_28  contact_28_109
timestamp 1707688321
transform 1 0 5664 0 1 13355
box 0 0 1 1
use contact_28  contact_28_110
timestamp 1707688321
transform 1 0 5664 0 1 12929
box 0 0 1 1
use contact_28  contact_28_111
timestamp 1707688321
transform 1 0 5664 0 1 12727
box 0 0 1 1
use contact_28  contact_28_112
timestamp 1707688321
transform 1 0 5664 0 1 15887
box 0 0 1 1
use contact_28  contact_28_113
timestamp 1707688321
transform 1 0 5664 0 1 18683
box 0 0 1 1
use contact_28  contact_28_114
timestamp 1707688321
transform 1 0 5664 0 1 18885
box 0 0 1 1
use contact_28  contact_28_115
timestamp 1707688321
transform 1 0 5664 0 1 18459
box 0 0 1 1
use contact_28  contact_28_116
timestamp 1707688321
transform 1 0 5664 0 1 18257
box 0 0 1 1
use contact_28  contact_28_117
timestamp 1707688321
transform 1 0 5664 0 1 17893
box 0 0 1 1
use contact_28  contact_28_118
timestamp 1707688321
transform 1 0 5664 0 1 18095
box 0 0 1 1
use contact_28  contact_28_119
timestamp 1707688321
transform 1 0 5664 0 1 17669
box 0 0 1 1
use contact_28  contact_28_120
timestamp 1707688321
transform 1 0 5664 0 1 17467
box 0 0 1 1
use contact_28  contact_28_121
timestamp 1707688321
transform 1 0 5664 0 1 17103
box 0 0 1 1
use contact_28  contact_28_122
timestamp 1707688321
transform 1 0 5664 0 1 17305
box 0 0 1 1
use contact_28  contact_28_123
timestamp 1707688321
transform 1 0 5664 0 1 16879
box 0 0 1 1
use contact_28  contact_28_124
timestamp 1707688321
transform 1 0 5664 0 1 16677
box 0 0 1 1
use contact_28  contact_28_125
timestamp 1707688321
transform 1 0 5664 0 1 16313
box 0 0 1 1
use contact_28  contact_28_126
timestamp 1707688321
transform 1 0 5664 0 1 16515
box 0 0 1 1
use contact_28  contact_28_127
timestamp 1707688321
transform 1 0 5664 0 1 16089
box 0 0 1 1
use contact_28  contact_28_128
timestamp 1707688321
transform 1 0 5554 0 1 15999
box 0 0 1 1
use contact_28  contact_28_129
timestamp 1707688321
transform 1 0 5554 0 1 18773
box 0 0 1 1
use contact_28  contact_28_130
timestamp 1707688321
transform 1 0 5554 0 1 15613
box 0 0 1 1
use contact_28  contact_28_131
timestamp 1707688321
transform 1 0 5554 0 1 15209
box 0 0 1 1
use contact_28  contact_28_132
timestamp 1707688321
transform 1 0 5554 0 1 14033
box 0 0 1 1
use contact_28  contact_28_133
timestamp 1707688321
transform 1 0 5554 0 1 18369
box 0 0 1 1
use contact_28  contact_28_134
timestamp 1707688321
transform 1 0 5554 0 1 13243
box 0 0 1 1
use contact_28  contact_28_135
timestamp 1707688321
transform 1 0 5554 0 1 17193
box 0 0 1 1
use contact_28  contact_28_136
timestamp 1707688321
transform 1 0 5554 0 1 14823
box 0 0 1 1
use contact_28  contact_28_137
timestamp 1707688321
transform 1 0 5554 0 1 17983
box 0 0 1 1
use contact_28  contact_28_138
timestamp 1707688321
transform 1 0 5554 0 1 16403
box 0 0 1 1
use contact_28  contact_28_139
timestamp 1707688321
transform 1 0 5554 0 1 13629
box 0 0 1 1
use contact_28  contact_28_140
timestamp 1707688321
transform 1 0 5554 0 1 14419
box 0 0 1 1
use contact_28  contact_28_141
timestamp 1707688321
transform 1 0 5554 0 1 17579
box 0 0 1 1
use contact_28  contact_28_142
timestamp 1707688321
transform 1 0 5554 0 1 12839
box 0 0 1 1
use contact_28  contact_28_143
timestamp 1707688321
transform 1 0 5554 0 1 16789
box 0 0 1 1
use contact_28  contact_28_144
timestamp 1707688321
transform 1 0 5554 0 1 23513
box 0 0 1 1
use contact_28  contact_28_145
timestamp 1707688321
transform 1 0 5554 0 1 21933
box 0 0 1 1
use contact_28  contact_28_146
timestamp 1707688321
transform 1 0 5554 0 1 25093
box 0 0 1 1
use contact_28  contact_28_147
timestamp 1707688321
transform 1 0 5554 0 1 21529
box 0 0 1 1
use contact_28  contact_28_148
timestamp 1707688321
transform 1 0 5554 0 1 23899
box 0 0 1 1
use contact_28  contact_28_149
timestamp 1707688321
transform 1 0 5554 0 1 21143
box 0 0 1 1
use contact_28  contact_28_150
timestamp 1707688321
transform 1 0 5554 0 1 22723
box 0 0 1 1
use contact_28  contact_28_151
timestamp 1707688321
transform 1 0 5554 0 1 20739
box 0 0 1 1
use contact_28  contact_28_152
timestamp 1707688321
transform 1 0 5554 0 1 23109
box 0 0 1 1
use contact_28  contact_28_153
timestamp 1707688321
transform 1 0 5554 0 1 20353
box 0 0 1 1
use contact_28  contact_28_154
timestamp 1707688321
transform 1 0 5554 0 1 19949
box 0 0 1 1
use contact_28  contact_28_155
timestamp 1707688321
transform 1 0 5554 0 1 24689
box 0 0 1 1
use contact_28  contact_28_156
timestamp 1707688321
transform 1 0 5554 0 1 19563
box 0 0 1 1
use contact_28  contact_28_157
timestamp 1707688321
transform 1 0 5554 0 1 19159
box 0 0 1 1
use contact_28  contact_28_158
timestamp 1707688321
transform 1 0 5554 0 1 22319
box 0 0 1 1
use contact_28  contact_28_159
timestamp 1707688321
transform 1 0 5554 0 1 24303
box 0 0 1 1
use contact_28  contact_28_160
timestamp 1707688321
transform 1 0 5664 0 1 22045
box 0 0 1 1
use contact_28  contact_28_161
timestamp 1707688321
transform 1 0 5664 0 1 21619
box 0 0 1 1
use contact_28  contact_28_162
timestamp 1707688321
transform 1 0 5664 0 1 21417
box 0 0 1 1
use contact_28  contact_28_163
timestamp 1707688321
transform 1 0 5664 0 1 21053
box 0 0 1 1
use contact_28  contact_28_164
timestamp 1707688321
transform 1 0 5664 0 1 21255
box 0 0 1 1
use contact_28  contact_28_165
timestamp 1707688321
transform 1 0 5664 0 1 20829
box 0 0 1 1
use contact_28  contact_28_166
timestamp 1707688321
transform 1 0 5664 0 1 20627
box 0 0 1 1
use contact_28  contact_28_167
timestamp 1707688321
transform 1 0 5664 0 1 20263
box 0 0 1 1
use contact_28  contact_28_168
timestamp 1707688321
transform 1 0 5664 0 1 20465
box 0 0 1 1
use contact_28  contact_28_169
timestamp 1707688321
transform 1 0 5664 0 1 20039
box 0 0 1 1
use contact_28  contact_28_170
timestamp 1707688321
transform 1 0 5664 0 1 19837
box 0 0 1 1
use contact_28  contact_28_171
timestamp 1707688321
transform 1 0 5664 0 1 19473
box 0 0 1 1
use contact_28  contact_28_172
timestamp 1707688321
transform 1 0 5664 0 1 19675
box 0 0 1 1
use contact_28  contact_28_173
timestamp 1707688321
transform 1 0 5664 0 1 19249
box 0 0 1 1
use contact_28  contact_28_174
timestamp 1707688321
transform 1 0 5664 0 1 19047
box 0 0 1 1
use contact_28  contact_28_175
timestamp 1707688321
transform 1 0 5664 0 1 21843
box 0 0 1 1
use contact_28  contact_28_176
timestamp 1707688321
transform 1 0 5664 0 1 25003
box 0 0 1 1
use contact_28  contact_28_177
timestamp 1707688321
transform 1 0 5664 0 1 25205
box 0 0 1 1
use contact_28  contact_28_178
timestamp 1707688321
transform 1 0 5664 0 1 24779
box 0 0 1 1
use contact_28  contact_28_179
timestamp 1707688321
transform 1 0 5664 0 1 24577
box 0 0 1 1
use contact_28  contact_28_180
timestamp 1707688321
transform 1 0 5664 0 1 24213
box 0 0 1 1
use contact_28  contact_28_181
timestamp 1707688321
transform 1 0 5664 0 1 24415
box 0 0 1 1
use contact_28  contact_28_182
timestamp 1707688321
transform 1 0 5664 0 1 23989
box 0 0 1 1
use contact_28  contact_28_183
timestamp 1707688321
transform 1 0 5664 0 1 23787
box 0 0 1 1
use contact_28  contact_28_184
timestamp 1707688321
transform 1 0 5664 0 1 22207
box 0 0 1 1
use contact_28  contact_28_185
timestamp 1707688321
transform 1 0 5664 0 1 23423
box 0 0 1 1
use contact_28  contact_28_186
timestamp 1707688321
transform 1 0 5664 0 1 23625
box 0 0 1 1
use contact_28  contact_28_187
timestamp 1707688321
transform 1 0 5664 0 1 23199
box 0 0 1 1
use contact_28  contact_28_188
timestamp 1707688321
transform 1 0 5664 0 1 22997
box 0 0 1 1
use contact_28  contact_28_189
timestamp 1707688321
transform 1 0 5664 0 1 22633
box 0 0 1 1
use contact_28  contact_28_190
timestamp 1707688321
transform 1 0 5664 0 1 22835
box 0 0 1 1
use contact_28  contact_28_191
timestamp 1707688321
transform 1 0 5664 0 1 22409
box 0 0 1 1
use contact_28  contact_28_192
timestamp 1707688321
transform 1 0 5664 0 1 27939
box 0 0 1 1
use contact_28  contact_28_193
timestamp 1707688321
transform 1 0 5664 0 1 26583
box 0 0 1 1
use contact_28  contact_28_194
timestamp 1707688321
transform 1 0 5664 0 1 26157
box 0 0 1 1
use contact_28  contact_28_195
timestamp 1707688321
transform 1 0 5664 0 1 25995
box 0 0 1 1
use contact_28  contact_28_196
timestamp 1707688321
transform 1 0 5664 0 1 26947
box 0 0 1 1
use contact_28  contact_28_197
timestamp 1707688321
transform 1 0 5664 0 1 27737
box 0 0 1 1
use contact_28  contact_28_198
timestamp 1707688321
transform 1 0 5664 0 1 27149
box 0 0 1 1
use contact_28  contact_28_199
timestamp 1707688321
transform 1 0 5664 0 1 25793
box 0 0 1 1
use contact_28  contact_28_200
timestamp 1707688321
transform 1 0 5664 0 1 27373
box 0 0 1 1
use contact_28  contact_28_201
timestamp 1707688321
transform 1 0 5664 0 1 26785
box 0 0 1 1
use contact_28  contact_28_202
timestamp 1707688321
transform 1 0 5664 0 1 25367
box 0 0 1 1
use contact_28  contact_28_203
timestamp 1707688321
transform 1 0 5664 0 1 25569
box 0 0 1 1
use contact_28  contact_28_204
timestamp 1707688321
transform 1 0 5664 0 1 28365
box 0 0 1 1
use contact_28  contact_28_205
timestamp 1707688321
transform 1 0 5664 0 1 27575
box 0 0 1 1
use contact_28  contact_28_206
timestamp 1707688321
transform 1 0 5664 0 1 26359
box 0 0 1 1
use contact_28  contact_28_207
timestamp 1707688321
transform 1 0 5664 0 1 28163
box 0 0 1 1
use contact_28  contact_28_208
timestamp 1707688321
transform 1 0 5664 0 1 30107
box 0 0 1 1
use contact_28  contact_28_209
timestamp 1707688321
transform 1 0 5664 0 1 29743
box 0 0 1 1
use contact_28  contact_28_210
timestamp 1707688321
transform 1 0 5664 0 1 29945
box 0 0 1 1
use contact_28  contact_28_211
timestamp 1707688321
transform 1 0 5664 0 1 29519
box 0 0 1 1
use contact_28  contact_28_212
timestamp 1707688321
transform 1 0 5664 0 1 29317
box 0 0 1 1
use contact_28  contact_28_213
timestamp 1707688321
transform 1 0 5664 0 1 28953
box 0 0 1 1
use contact_28  contact_28_214
timestamp 1707688321
transform 1 0 5664 0 1 30309
box 0 0 1 1
use contact_28  contact_28_215
timestamp 1707688321
transform 1 0 5664 0 1 29155
box 0 0 1 1
use contact_28  contact_28_216
timestamp 1707688321
transform 1 0 5664 0 1 31323
box 0 0 1 1
use contact_28  contact_28_217
timestamp 1707688321
transform 1 0 5664 0 1 28729
box 0 0 1 1
use contact_28  contact_28_218
timestamp 1707688321
transform 1 0 5664 0 1 31525
box 0 0 1 1
use contact_28  contact_28_219
timestamp 1707688321
transform 1 0 5664 0 1 31099
box 0 0 1 1
use contact_28  contact_28_220
timestamp 1707688321
transform 1 0 5664 0 1 28527
box 0 0 1 1
use contact_28  contact_28_221
timestamp 1707688321
transform 1 0 5664 0 1 30897
box 0 0 1 1
use contact_28  contact_28_222
timestamp 1707688321
transform 1 0 5664 0 1 30533
box 0 0 1 1
use contact_28  contact_28_223
timestamp 1707688321
transform 1 0 5664 0 1 30735
box 0 0 1 1
use contact_28  contact_28_224
timestamp 1707688321
transform 1 0 5554 0 1 27059
box 0 0 1 1
use contact_28  contact_28_225
timestamp 1707688321
transform 1 0 5554 0 1 30623
box 0 0 1 1
use contact_28  contact_28_226
timestamp 1707688321
transform 1 0 5554 0 1 30219
box 0 0 1 1
use contact_28  contact_28_227
timestamp 1707688321
transform 1 0 5554 0 1 29833
box 0 0 1 1
use contact_28  contact_28_228
timestamp 1707688321
transform 1 0 5554 0 1 29429
box 0 0 1 1
use contact_28  contact_28_229
timestamp 1707688321
transform 1 0 5554 0 1 29043
box 0 0 1 1
use contact_28  contact_28_230
timestamp 1707688321
transform 1 0 5554 0 1 26673
box 0 0 1 1
use contact_28  contact_28_231
timestamp 1707688321
transform 1 0 5554 0 1 28639
box 0 0 1 1
use contact_28  contact_28_232
timestamp 1707688321
transform 1 0 5554 0 1 25883
box 0 0 1 1
use contact_28  contact_28_233
timestamp 1707688321
transform 1 0 5554 0 1 28253
box 0 0 1 1
use contact_28  contact_28_234
timestamp 1707688321
transform 1 0 5554 0 1 27849
box 0 0 1 1
use contact_28  contact_28_235
timestamp 1707688321
transform 1 0 5554 0 1 26269
box 0 0 1 1
use contact_28  contact_28_236
timestamp 1707688321
transform 1 0 5554 0 1 27463
box 0 0 1 1
use contact_28  contact_28_237
timestamp 1707688321
transform 1 0 5554 0 1 25479
box 0 0 1 1
use contact_28  contact_28_238
timestamp 1707688321
transform 1 0 5554 0 1 31413
box 0 0 1 1
use contact_28  contact_28_239
timestamp 1707688321
transform 1 0 5554 0 1 31009
box 0 0 1 1
use contact_28  contact_28_240
timestamp 1707688321
transform 1 0 5554 0 1 35749
box 0 0 1 1
use contact_28  contact_28_241
timestamp 1707688321
transform 1 0 5554 0 1 35363
box 0 0 1 1
use contact_28  contact_28_242
timestamp 1707688321
transform 1 0 5554 0 1 34959
box 0 0 1 1
use contact_28  contact_28_243
timestamp 1707688321
transform 1 0 5554 0 1 34573
box 0 0 1 1
use contact_28  contact_28_244
timestamp 1707688321
transform 1 0 5554 0 1 34169
box 0 0 1 1
use contact_28  contact_28_245
timestamp 1707688321
transform 1 0 5554 0 1 33783
box 0 0 1 1
use contact_28  contact_28_246
timestamp 1707688321
transform 1 0 5554 0 1 36539
box 0 0 1 1
use contact_28  contact_28_247
timestamp 1707688321
transform 1 0 5554 0 1 33379
box 0 0 1 1
use contact_28  contact_28_248
timestamp 1707688321
transform 1 0 5554 0 1 32993
box 0 0 1 1
use contact_28  contact_28_249
timestamp 1707688321
transform 1 0 5554 0 1 32589
box 0 0 1 1
use contact_28  contact_28_250
timestamp 1707688321
transform 1 0 5554 0 1 32203
box 0 0 1 1
use contact_28  contact_28_251
timestamp 1707688321
transform 1 0 5554 0 1 31799
box 0 0 1 1
use contact_28  contact_28_252
timestamp 1707688321
transform 1 0 5554 0 1 36153
box 0 0 1 1
use contact_28  contact_28_253
timestamp 1707688321
transform 1 0 5554 0 1 37733
box 0 0 1 1
use contact_28  contact_28_254
timestamp 1707688321
transform 1 0 5554 0 1 37329
box 0 0 1 1
use contact_28  contact_28_255
timestamp 1707688321
transform 1 0 5554 0 1 36943
box 0 0 1 1
use contact_28  contact_28_256
timestamp 1707688321
transform 1 0 5664 0 1 34057
box 0 0 1 1
use contact_28  contact_28_257
timestamp 1707688321
transform 1 0 5664 0 1 33693
box 0 0 1 1
use contact_28  contact_28_258
timestamp 1707688321
transform 1 0 5664 0 1 33895
box 0 0 1 1
use contact_28  contact_28_259
timestamp 1707688321
transform 1 0 5664 0 1 33469
box 0 0 1 1
use contact_28  contact_28_260
timestamp 1707688321
transform 1 0 5664 0 1 33267
box 0 0 1 1
use contact_28  contact_28_261
timestamp 1707688321
transform 1 0 5664 0 1 32903
box 0 0 1 1
use contact_28  contact_28_262
timestamp 1707688321
transform 1 0 5664 0 1 33105
box 0 0 1 1
use contact_28  contact_28_263
timestamp 1707688321
transform 1 0 5664 0 1 32679
box 0 0 1 1
use contact_28  contact_28_264
timestamp 1707688321
transform 1 0 5664 0 1 32477
box 0 0 1 1
use contact_28  contact_28_265
timestamp 1707688321
transform 1 0 5664 0 1 32113
box 0 0 1 1
use contact_28  contact_28_266
timestamp 1707688321
transform 1 0 5664 0 1 34685
box 0 0 1 1
use contact_28  contact_28_267
timestamp 1707688321
transform 1 0 5664 0 1 32315
box 0 0 1 1
use contact_28  contact_28_268
timestamp 1707688321
transform 1 0 5664 0 1 31889
box 0 0 1 1
use contact_28  contact_28_269
timestamp 1707688321
transform 1 0 5664 0 1 34259
box 0 0 1 1
use contact_28  contact_28_270
timestamp 1707688321
transform 1 0 5664 0 1 31687
box 0 0 1 1
use contact_28  contact_28_271
timestamp 1707688321
transform 1 0 5664 0 1 34483
box 0 0 1 1
use contact_28  contact_28_272
timestamp 1707688321
transform 1 0 5664 0 1 37643
box 0 0 1 1
use contact_28  contact_28_273
timestamp 1707688321
transform 1 0 5664 0 1 37845
box 0 0 1 1
use contact_28  contact_28_274
timestamp 1707688321
transform 1 0 5664 0 1 37419
box 0 0 1 1
use contact_28  contact_28_275
timestamp 1707688321
transform 1 0 5664 0 1 37217
box 0 0 1 1
use contact_28  contact_28_276
timestamp 1707688321
transform 1 0 5664 0 1 36853
box 0 0 1 1
use contact_28  contact_28_277
timestamp 1707688321
transform 1 0 5664 0 1 37055
box 0 0 1 1
use contact_28  contact_28_278
timestamp 1707688321
transform 1 0 5664 0 1 36629
box 0 0 1 1
use contact_28  contact_28_279
timestamp 1707688321
transform 1 0 5664 0 1 36427
box 0 0 1 1
use contact_28  contact_28_280
timestamp 1707688321
transform 1 0 5664 0 1 36063
box 0 0 1 1
use contact_28  contact_28_281
timestamp 1707688321
transform 1 0 5664 0 1 36265
box 0 0 1 1
use contact_28  contact_28_282
timestamp 1707688321
transform 1 0 5664 0 1 35839
box 0 0 1 1
use contact_28  contact_28_283
timestamp 1707688321
transform 1 0 5664 0 1 35637
box 0 0 1 1
use contact_28  contact_28_284
timestamp 1707688321
transform 1 0 5664 0 1 35273
box 0 0 1 1
use contact_28  contact_28_285
timestamp 1707688321
transform 1 0 5664 0 1 35475
box 0 0 1 1
use contact_28  contact_28_286
timestamp 1707688321
transform 1 0 5664 0 1 35049
box 0 0 1 1
use contact_28  contact_28_287
timestamp 1707688321
transform 1 0 5664 0 1 34847
box 0 0 1 1
use contact_28  contact_28_288
timestamp 1707688321
transform 1 0 5664 0 1 40013
box 0 0 1 1
use contact_28  contact_28_289
timestamp 1707688321
transform 1 0 5664 0 1 40215
box 0 0 1 1
use contact_28  contact_28_290
timestamp 1707688321
transform 1 0 5664 0 1 39789
box 0 0 1 1
use contact_28  contact_28_291
timestamp 1707688321
transform 1 0 5664 0 1 39587
box 0 0 1 1
use contact_28  contact_28_292
timestamp 1707688321
transform 1 0 5664 0 1 39223
box 0 0 1 1
use contact_28  contact_28_293
timestamp 1707688321
transform 1 0 5664 0 1 39425
box 0 0 1 1
use contact_28  contact_28_294
timestamp 1707688321
transform 1 0 5664 0 1 38999
box 0 0 1 1
use contact_28  contact_28_295
timestamp 1707688321
transform 1 0 5664 0 1 38797
box 0 0 1 1
use contact_28  contact_28_296
timestamp 1707688321
transform 1 0 5664 0 1 38433
box 0 0 1 1
use contact_28  contact_28_297
timestamp 1707688321
transform 1 0 5664 0 1 38635
box 0 0 1 1
use contact_28  contact_28_298
timestamp 1707688321
transform 1 0 5664 0 1 38209
box 0 0 1 1
use contact_28  contact_28_299
timestamp 1707688321
transform 1 0 5664 0 1 38007
box 0 0 1 1
use contact_28  contact_28_300
timestamp 1707688321
transform 1 0 5664 0 1 40803
box 0 0 1 1
use contact_28  contact_28_301
timestamp 1707688321
transform 1 0 5664 0 1 41005
box 0 0 1 1
use contact_28  contact_28_302
timestamp 1707688321
transform 1 0 5664 0 1 40579
box 0 0 1 1
use contact_28  contact_28_303
timestamp 1707688321
transform 1 0 5664 0 1 40377
box 0 0 1 1
use contact_28  contact_28_304
timestamp 1707688321
transform 1 0 5664 0 1 43173
box 0 0 1 1
use contact_28  contact_28_305
timestamp 1707688321
transform 1 0 5664 0 1 43375
box 0 0 1 1
use contact_28  contact_28_306
timestamp 1707688321
transform 1 0 5664 0 1 42949
box 0 0 1 1
use contact_28  contact_28_307
timestamp 1707688321
transform 1 0 5664 0 1 42747
box 0 0 1 1
use contact_28  contact_28_308
timestamp 1707688321
transform 1 0 5664 0 1 42383
box 0 0 1 1
use contact_28  contact_28_309
timestamp 1707688321
transform 1 0 5664 0 1 42585
box 0 0 1 1
use contact_28  contact_28_310
timestamp 1707688321
transform 1 0 5664 0 1 42159
box 0 0 1 1
use contact_28  contact_28_311
timestamp 1707688321
transform 1 0 5664 0 1 41957
box 0 0 1 1
use contact_28  contact_28_312
timestamp 1707688321
transform 1 0 5664 0 1 41593
box 0 0 1 1
use contact_28  contact_28_313
timestamp 1707688321
transform 1 0 5664 0 1 41795
box 0 0 1 1
use contact_28  contact_28_314
timestamp 1707688321
transform 1 0 5664 0 1 41369
box 0 0 1 1
use contact_28  contact_28_315
timestamp 1707688321
transform 1 0 5664 0 1 41167
box 0 0 1 1
use contact_28  contact_28_316
timestamp 1707688321
transform 1 0 5664 0 1 43963
box 0 0 1 1
use contact_28  contact_28_317
timestamp 1707688321
transform 1 0 5664 0 1 44165
box 0 0 1 1
use contact_28  contact_28_318
timestamp 1707688321
transform 1 0 5664 0 1 43739
box 0 0 1 1
use contact_28  contact_28_319
timestamp 1707688321
transform 1 0 5664 0 1 43537
box 0 0 1 1
use contact_28  contact_28_320
timestamp 1707688321
transform 1 0 5554 0 1 40489
box 0 0 1 1
use contact_28  contact_28_321
timestamp 1707688321
transform 1 0 5554 0 1 43649
box 0 0 1 1
use contact_28  contact_28_322
timestamp 1707688321
transform 1 0 5554 0 1 38119
box 0 0 1 1
use contact_28  contact_28_323
timestamp 1707688321
transform 1 0 5554 0 1 39313
box 0 0 1 1
use contact_28  contact_28_324
timestamp 1707688321
transform 1 0 5554 0 1 42473
box 0 0 1 1
use contact_28  contact_28_325
timestamp 1707688321
transform 1 0 5554 0 1 43263
box 0 0 1 1
use contact_28  contact_28_326
timestamp 1707688321
transform 1 0 5554 0 1 38909
box 0 0 1 1
use contact_28  contact_28_327
timestamp 1707688321
transform 1 0 5554 0 1 41279
box 0 0 1 1
use contact_28  contact_28_328
timestamp 1707688321
transform 1 0 5554 0 1 41683
box 0 0 1 1
use contact_28  contact_28_329
timestamp 1707688321
transform 1 0 5554 0 1 38523
box 0 0 1 1
use contact_28  contact_28_330
timestamp 1707688321
transform 1 0 5554 0 1 42859
box 0 0 1 1
use contact_28  contact_28_331
timestamp 1707688321
transform 1 0 5554 0 1 40103
box 0 0 1 1
use contact_28  contact_28_332
timestamp 1707688321
transform 1 0 5554 0 1 42069
box 0 0 1 1
use contact_28  contact_28_333
timestamp 1707688321
transform 1 0 5554 0 1 44053
box 0 0 1 1
use contact_28  contact_28_334
timestamp 1707688321
transform 1 0 5554 0 1 40893
box 0 0 1 1
use contact_28  contact_28_335
timestamp 1707688321
transform 1 0 5554 0 1 39699
box 0 0 1 1
use contact_28  contact_28_336
timestamp 1707688321
transform 1 0 5554 0 1 45229
box 0 0 1 1
use contact_28  contact_28_337
timestamp 1707688321
transform 1 0 5554 0 1 50373
box 0 0 1 1
use contact_28  contact_28_338
timestamp 1707688321
transform 1 0 5554 0 1 49969
box 0 0 1 1
use contact_28  contact_28_339
timestamp 1707688321
transform 1 0 5554 0 1 49583
box 0 0 1 1
use contact_28  contact_28_340
timestamp 1707688321
transform 1 0 5554 0 1 49179
box 0 0 1 1
use contact_28  contact_28_341
timestamp 1707688321
transform 1 0 5554 0 1 48793
box 0 0 1 1
use contact_28  contact_28_342
timestamp 1707688321
transform 1 0 5554 0 1 48389
box 0 0 1 1
use contact_28  contact_28_343
timestamp 1707688321
transform 1 0 5554 0 1 48003
box 0 0 1 1
use contact_28  contact_28_344
timestamp 1707688321
transform 1 0 5554 0 1 47599
box 0 0 1 1
use contact_28  contact_28_345
timestamp 1707688321
transform 1 0 5554 0 1 47213
box 0 0 1 1
use contact_28  contact_28_346
timestamp 1707688321
transform 1 0 5554 0 1 46809
box 0 0 1 1
use contact_28  contact_28_347
timestamp 1707688321
transform 1 0 5554 0 1 44843
box 0 0 1 1
use contact_28  contact_28_348
timestamp 1707688321
transform 1 0 5554 0 1 44439
box 0 0 1 1
use contact_28  contact_28_349
timestamp 1707688321
transform 1 0 5554 0 1 46423
box 0 0 1 1
use contact_28  contact_28_350
timestamp 1707688321
transform 1 0 5554 0 1 46019
box 0 0 1 1
use contact_28  contact_28_351
timestamp 1707688321
transform 1 0 5554 0 1 45633
box 0 0 1 1
use contact_28  contact_28_352
timestamp 1707688321
transform 1 0 5664 0 1 46109
box 0 0 1 1
use contact_28  contact_28_353
timestamp 1707688321
transform 1 0 5664 0 1 45907
box 0 0 1 1
use contact_28  contact_28_354
timestamp 1707688321
transform 1 0 5664 0 1 45319
box 0 0 1 1
use contact_28  contact_28_355
timestamp 1707688321
transform 1 0 5664 0 1 45117
box 0 0 1 1
use contact_28  contact_28_356
timestamp 1707688321
transform 1 0 5664 0 1 46899
box 0 0 1 1
use contact_28  contact_28_357
timestamp 1707688321
transform 1 0 5664 0 1 46697
box 0 0 1 1
use contact_28  contact_28_358
timestamp 1707688321
transform 1 0 5664 0 1 45543
box 0 0 1 1
use contact_28  contact_28_359
timestamp 1707688321
transform 1 0 5664 0 1 45745
box 0 0 1 1
use contact_28  contact_28_360
timestamp 1707688321
transform 1 0 5664 0 1 44753
box 0 0 1 1
use contact_28  contact_28_361
timestamp 1707688321
transform 1 0 5664 0 1 44955
box 0 0 1 1
use contact_28  contact_28_362
timestamp 1707688321
transform 1 0 5664 0 1 44529
box 0 0 1 1
use contact_28  contact_28_363
timestamp 1707688321
transform 1 0 5664 0 1 44327
box 0 0 1 1
use contact_28  contact_28_364
timestamp 1707688321
transform 1 0 5664 0 1 46333
box 0 0 1 1
use contact_28  contact_28_365
timestamp 1707688321
transform 1 0 5664 0 1 46535
box 0 0 1 1
use contact_28  contact_28_366
timestamp 1707688321
transform 1 0 5664 0 1 47123
box 0 0 1 1
use contact_28  contact_28_367
timestamp 1707688321
transform 1 0 5664 0 1 47325
box 0 0 1 1
use contact_28  contact_28_368
timestamp 1707688321
transform 1 0 5664 0 1 48479
box 0 0 1 1
use contact_28  contact_28_369
timestamp 1707688321
transform 1 0 5664 0 1 48277
box 0 0 1 1
use contact_28  contact_28_370
timestamp 1707688321
transform 1 0 5664 0 1 47689
box 0 0 1 1
use contact_28  contact_28_371
timestamp 1707688321
transform 1 0 5664 0 1 47487
box 0 0 1 1
use contact_28  contact_28_372
timestamp 1707688321
transform 1 0 5664 0 1 47913
box 0 0 1 1
use contact_28  contact_28_373
timestamp 1707688321
transform 1 0 5664 0 1 48115
box 0 0 1 1
use contact_28  contact_28_374
timestamp 1707688321
transform 1 0 5664 0 1 50283
box 0 0 1 1
use contact_28  contact_28_375
timestamp 1707688321
transform 1 0 5664 0 1 50485
box 0 0 1 1
use contact_28  contact_28_376
timestamp 1707688321
transform 1 0 5664 0 1 50059
box 0 0 1 1
use contact_28  contact_28_377
timestamp 1707688321
transform 1 0 5664 0 1 49857
box 0 0 1 1
use contact_28  contact_28_378
timestamp 1707688321
transform 1 0 5664 0 1 49493
box 0 0 1 1
use contact_28  contact_28_379
timestamp 1707688321
transform 1 0 5664 0 1 49695
box 0 0 1 1
use contact_28  contact_28_380
timestamp 1707688321
transform 1 0 5664 0 1 49269
box 0 0 1 1
use contact_28  contact_28_381
timestamp 1707688321
transform 1 0 5664 0 1 49067
box 0 0 1 1
use contact_28  contact_28_382
timestamp 1707688321
transform 1 0 5664 0 1 48703
box 0 0 1 1
use contact_28  contact_28_383
timestamp 1707688321
transform 1 0 5664 0 1 48905
box 0 0 1 1
use contact_29  contact_29_0
timestamp 1707688321
transform 1 0 5665 0 1 1076
box 0 0 1 1
use contact_29  contact_29_1
timestamp 1707688321
transform 1 0 5665 0 1 3082
box 0 0 1 1
use contact_29  contact_29_2
timestamp 1707688321
transform 1 0 5665 0 1 2090
box 0 0 1 1
use contact_29  contact_29_3
timestamp 1707688321
transform 1 0 5665 0 1 1866
box 0 0 1 1
use contact_29  contact_29_4
timestamp 1707688321
transform 1 0 5665 0 1 286
box 0 0 1 1
use contact_29  contact_29_5
timestamp 1707688321
transform 1 0 5665 0 1 1300
box 0 0 1 1
use contact_29  contact_29_6
timestamp 1707688321
transform 1 0 5665 0 1 2656
box 0 0 1 1
use contact_29  contact_29_7
timestamp 1707688321
transform 1 0 5665 0 1 510
box 0 0 1 1
use contact_29  contact_29_8
timestamp 1707688321
transform 1 0 5665 0 1 84
box 0 0 1 1
use contact_29  contact_29_9
timestamp 1707688321
transform 1 0 5665 0 1 2454
box 0 0 1 1
use contact_29  contact_29_10
timestamp 1707688321
transform 1 0 5665 0 1 2880
box 0 0 1 1
use contact_29  contact_29_11
timestamp 1707688321
transform 1 0 5665 0 1 1502
box 0 0 1 1
use contact_29  contact_29_12
timestamp 1707688321
transform 1 0 5665 0 1 2292
box 0 0 1 1
use contact_29  contact_29_13
timestamp 1707688321
transform 1 0 5665 0 1 712
box 0 0 1 1
use contact_29  contact_29_14
timestamp 1707688321
transform 1 0 5665 0 1 1664
box 0 0 1 1
use contact_29  contact_29_15
timestamp 1707688321
transform 1 0 5665 0 1 874
box 0 0 1 1
use contact_29  contact_29_16
timestamp 1707688321
transform 1 0 5665 0 1 3446
box 0 0 1 1
use contact_29  contact_29_17
timestamp 1707688321
transform 1 0 5665 0 1 6040
box 0 0 1 1
use contact_29  contact_29_18
timestamp 1707688321
transform 1 0 5665 0 1 6242
box 0 0 1 1
use contact_29  contact_29_19
timestamp 1707688321
transform 1 0 5665 0 1 5816
box 0 0 1 1
use contact_29  contact_29_20
timestamp 1707688321
transform 1 0 5665 0 1 3244
box 0 0 1 1
use contact_29  contact_29_21
timestamp 1707688321
transform 1 0 5665 0 1 4662
box 0 0 1 1
use contact_29  contact_29_22
timestamp 1707688321
transform 1 0 5665 0 1 5614
box 0 0 1 1
use contact_29  contact_29_23
timestamp 1707688321
transform 1 0 5665 0 1 5250
box 0 0 1 1
use contact_29  contact_29_24
timestamp 1707688321
transform 1 0 5665 0 1 4236
box 0 0 1 1
use contact_29  contact_29_25
timestamp 1707688321
transform 1 0 5665 0 1 5452
box 0 0 1 1
use contact_29  contact_29_26
timestamp 1707688321
transform 1 0 5665 0 1 5026
box 0 0 1 1
use contact_29  contact_29_27
timestamp 1707688321
transform 1 0 5665 0 1 3670
box 0 0 1 1
use contact_29  contact_29_28
timestamp 1707688321
transform 1 0 5665 0 1 4824
box 0 0 1 1
use contact_29  contact_29_29
timestamp 1707688321
transform 1 0 5665 0 1 4460
box 0 0 1 1
use contact_29  contact_29_30
timestamp 1707688321
transform 1 0 5665 0 1 4034
box 0 0 1 1
use contact_29  contact_29_31
timestamp 1707688321
transform 1 0 5665 0 1 3872
box 0 0 1 1
use contact_29  contact_29_32
timestamp 1707688321
transform 1 0 5555 0 1 4146
box 0 0 1 1
use contact_29  contact_29_33
timestamp 1707688321
transform 1 0 5555 0 1 1390
box 0 0 1 1
use contact_29  contact_29_34
timestamp 1707688321
transform 1 0 5555 0 1 3760
box 0 0 1 1
use contact_29  contact_29_35
timestamp 1707688321
transform 1 0 5555 0 1 3356
box 0 0 1 1
use contact_29  contact_29_36
timestamp 1707688321
transform 1 0 5555 0 1 2970
box 0 0 1 1
use contact_29  contact_29_37
timestamp 1707688321
transform 1 0 5555 0 1 196
box 0 0 1 1
use contact_29  contact_29_38
timestamp 1707688321
transform 1 0 5555 0 1 2566
box 0 0 1 1
use contact_29  contact_29_39
timestamp 1707688321
transform 1 0 5555 0 1 986
box 0 0 1 1
use contact_29  contact_29_40
timestamp 1707688321
transform 1 0 5555 0 1 2180
box 0 0 1 1
use contact_29  contact_29_41
timestamp 1707688321
transform 1 0 5555 0 1 6130
box 0 0 1 1
use contact_29  contact_29_42
timestamp 1707688321
transform 1 0 5555 0 1 1776
box 0 0 1 1
use contact_29  contact_29_43
timestamp 1707688321
transform 1 0 5555 0 1 5726
box 0 0 1 1
use contact_29  contact_29_44
timestamp 1707688321
transform 1 0 5555 0 1 5340
box 0 0 1 1
use contact_29  contact_29_45
timestamp 1707688321
transform 1 0 5555 0 1 4936
box 0 0 1 1
use contact_29  contact_29_46
timestamp 1707688321
transform 1 0 5555 0 1 600
box 0 0 1 1
use contact_29  contact_29_47
timestamp 1707688321
transform 1 0 5555 0 1 4550
box 0 0 1 1
use contact_29  contact_29_48
timestamp 1707688321
transform 1 0 5555 0 1 11256
box 0 0 1 1
use contact_29  contact_29_49
timestamp 1707688321
transform 1 0 5555 0 1 10870
box 0 0 1 1
use contact_29  contact_29_50
timestamp 1707688321
transform 1 0 5555 0 1 10466
box 0 0 1 1
use contact_29  contact_29_51
timestamp 1707688321
transform 1 0 5555 0 1 10080
box 0 0 1 1
use contact_29  contact_29_52
timestamp 1707688321
transform 1 0 5555 0 1 9676
box 0 0 1 1
use contact_29  contact_29_53
timestamp 1707688321
transform 1 0 5555 0 1 9290
box 0 0 1 1
use contact_29  contact_29_54
timestamp 1707688321
transform 1 0 5555 0 1 6516
box 0 0 1 1
use contact_29  contact_29_55
timestamp 1707688321
transform 1 0 5555 0 1 8886
box 0 0 1 1
use contact_29  contact_29_56
timestamp 1707688321
transform 1 0 5555 0 1 8500
box 0 0 1 1
use contact_29  contact_29_57
timestamp 1707688321
transform 1 0 5555 0 1 8096
box 0 0 1 1
use contact_29  contact_29_58
timestamp 1707688321
transform 1 0 5555 0 1 7710
box 0 0 1 1
use contact_29  contact_29_59
timestamp 1707688321
transform 1 0 5555 0 1 7306
box 0 0 1 1
use contact_29  contact_29_60
timestamp 1707688321
transform 1 0 5555 0 1 6920
box 0 0 1 1
use contact_29  contact_29_61
timestamp 1707688321
transform 1 0 5555 0 1 12450
box 0 0 1 1
use contact_29  contact_29_62
timestamp 1707688321
transform 1 0 5555 0 1 12046
box 0 0 1 1
use contact_29  contact_29_63
timestamp 1707688321
transform 1 0 5555 0 1 11660
box 0 0 1 1
use contact_29  contact_29_64
timestamp 1707688321
transform 1 0 5665 0 1 7396
box 0 0 1 1
use contact_29  contact_29_65
timestamp 1707688321
transform 1 0 5665 0 1 7194
box 0 0 1 1
use contact_29  contact_29_66
timestamp 1707688321
transform 1 0 5665 0 1 9402
box 0 0 1 1
use contact_29  contact_29_67
timestamp 1707688321
transform 1 0 5665 0 1 8410
box 0 0 1 1
use contact_29  contact_29_68
timestamp 1707688321
transform 1 0 5665 0 1 8612
box 0 0 1 1
use contact_29  contact_29_69
timestamp 1707688321
transform 1 0 5665 0 1 6830
box 0 0 1 1
use contact_29  contact_29_70
timestamp 1707688321
transform 1 0 5665 0 1 9200
box 0 0 1 1
use contact_29  contact_29_71
timestamp 1707688321
transform 1 0 5665 0 1 8186
box 0 0 1 1
use contact_29  contact_29_72
timestamp 1707688321
transform 1 0 5665 0 1 8976
box 0 0 1 1
use contact_29  contact_29_73
timestamp 1707688321
transform 1 0 5665 0 1 7984
box 0 0 1 1
use contact_29  contact_29_74
timestamp 1707688321
transform 1 0 5665 0 1 7032
box 0 0 1 1
use contact_29  contact_29_75
timestamp 1707688321
transform 1 0 5665 0 1 6404
box 0 0 1 1
use contact_29  contact_29_76
timestamp 1707688321
transform 1 0 5665 0 1 7620
box 0 0 1 1
use contact_29  contact_29_77
timestamp 1707688321
transform 1 0 5665 0 1 8774
box 0 0 1 1
use contact_29  contact_29_78
timestamp 1707688321
transform 1 0 5665 0 1 6606
box 0 0 1 1
use contact_29  contact_29_79
timestamp 1707688321
transform 1 0 5665 0 1 7822
box 0 0 1 1
use contact_29  contact_29_80
timestamp 1707688321
transform 1 0 5665 0 1 11346
box 0 0 1 1
use contact_29  contact_29_81
timestamp 1707688321
transform 1 0 5665 0 1 11144
box 0 0 1 1
use contact_29  contact_29_82
timestamp 1707688321
transform 1 0 5665 0 1 10780
box 0 0 1 1
use contact_29  contact_29_83
timestamp 1707688321
transform 1 0 5665 0 1 10982
box 0 0 1 1
use contact_29  contact_29_84
timestamp 1707688321
transform 1 0 5665 0 1 10556
box 0 0 1 1
use contact_29  contact_29_85
timestamp 1707688321
transform 1 0 5665 0 1 11570
box 0 0 1 1
use contact_29  contact_29_86
timestamp 1707688321
transform 1 0 5665 0 1 9990
box 0 0 1 1
use contact_29  contact_29_87
timestamp 1707688321
transform 1 0 5665 0 1 10192
box 0 0 1 1
use contact_29  contact_29_88
timestamp 1707688321
transform 1 0 5665 0 1 11772
box 0 0 1 1
use contact_29  contact_29_89
timestamp 1707688321
transform 1 0 5665 0 1 10354
box 0 0 1 1
use contact_29  contact_29_90
timestamp 1707688321
transform 1 0 5665 0 1 9766
box 0 0 1 1
use contact_29  contact_29_91
timestamp 1707688321
transform 1 0 5665 0 1 9564
box 0 0 1 1
use contact_29  contact_29_92
timestamp 1707688321
transform 1 0 5665 0 1 12360
box 0 0 1 1
use contact_29  contact_29_93
timestamp 1707688321
transform 1 0 5665 0 1 12562
box 0 0 1 1
use contact_29  contact_29_94
timestamp 1707688321
transform 1 0 5665 0 1 12136
box 0 0 1 1
use contact_29  contact_29_95
timestamp 1707688321
transform 1 0 5665 0 1 11934
box 0 0 1 1
use contact_29  contact_29_96
timestamp 1707688321
transform 1 0 5665 0 1 15520
box 0 0 1 1
use contact_29  contact_29_97
timestamp 1707688321
transform 1 0 5665 0 1 15722
box 0 0 1 1
use contact_29  contact_29_98
timestamp 1707688321
transform 1 0 5665 0 1 15296
box 0 0 1 1
use contact_29  contact_29_99
timestamp 1707688321
transform 1 0 5665 0 1 15094
box 0 0 1 1
use contact_29  contact_29_100
timestamp 1707688321
transform 1 0 5665 0 1 14730
box 0 0 1 1
use contact_29  contact_29_101
timestamp 1707688321
transform 1 0 5665 0 1 14932
box 0 0 1 1
use contact_29  contact_29_102
timestamp 1707688321
transform 1 0 5665 0 1 14506
box 0 0 1 1
use contact_29  contact_29_103
timestamp 1707688321
transform 1 0 5665 0 1 14304
box 0 0 1 1
use contact_29  contact_29_104
timestamp 1707688321
transform 1 0 5665 0 1 13940
box 0 0 1 1
use contact_29  contact_29_105
timestamp 1707688321
transform 1 0 5665 0 1 14142
box 0 0 1 1
use contact_29  contact_29_106
timestamp 1707688321
transform 1 0 5665 0 1 13716
box 0 0 1 1
use contact_29  contact_29_107
timestamp 1707688321
transform 1 0 5665 0 1 13514
box 0 0 1 1
use contact_29  contact_29_108
timestamp 1707688321
transform 1 0 5665 0 1 13150
box 0 0 1 1
use contact_29  contact_29_109
timestamp 1707688321
transform 1 0 5665 0 1 13352
box 0 0 1 1
use contact_29  contact_29_110
timestamp 1707688321
transform 1 0 5665 0 1 12926
box 0 0 1 1
use contact_29  contact_29_111
timestamp 1707688321
transform 1 0 5665 0 1 12724
box 0 0 1 1
use contact_29  contact_29_112
timestamp 1707688321
transform 1 0 5665 0 1 18680
box 0 0 1 1
use contact_29  contact_29_113
timestamp 1707688321
transform 1 0 5665 0 1 18882
box 0 0 1 1
use contact_29  contact_29_114
timestamp 1707688321
transform 1 0 5665 0 1 18456
box 0 0 1 1
use contact_29  contact_29_115
timestamp 1707688321
transform 1 0 5665 0 1 18254
box 0 0 1 1
use contact_29  contact_29_116
timestamp 1707688321
transform 1 0 5665 0 1 17890
box 0 0 1 1
use contact_29  contact_29_117
timestamp 1707688321
transform 1 0 5665 0 1 18092
box 0 0 1 1
use contact_29  contact_29_118
timestamp 1707688321
transform 1 0 5665 0 1 17666
box 0 0 1 1
use contact_29  contact_29_119
timestamp 1707688321
transform 1 0 5665 0 1 17464
box 0 0 1 1
use contact_29  contact_29_120
timestamp 1707688321
transform 1 0 5665 0 1 17100
box 0 0 1 1
use contact_29  contact_29_121
timestamp 1707688321
transform 1 0 5665 0 1 17302
box 0 0 1 1
use contact_29  contact_29_122
timestamp 1707688321
transform 1 0 5665 0 1 16876
box 0 0 1 1
use contact_29  contact_29_123
timestamp 1707688321
transform 1 0 5665 0 1 16674
box 0 0 1 1
use contact_29  contact_29_124
timestamp 1707688321
transform 1 0 5665 0 1 16310
box 0 0 1 1
use contact_29  contact_29_125
timestamp 1707688321
transform 1 0 5665 0 1 16512
box 0 0 1 1
use contact_29  contact_29_126
timestamp 1707688321
transform 1 0 5665 0 1 16086
box 0 0 1 1
use contact_29  contact_29_127
timestamp 1707688321
transform 1 0 5665 0 1 15884
box 0 0 1 1
use contact_29  contact_29_128
timestamp 1707688321
transform 1 0 5555 0 1 15996
box 0 0 1 1
use contact_29  contact_29_129
timestamp 1707688321
transform 1 0 5555 0 1 18770
box 0 0 1 1
use contact_29  contact_29_130
timestamp 1707688321
transform 1 0 5555 0 1 15610
box 0 0 1 1
use contact_29  contact_29_131
timestamp 1707688321
transform 1 0 5555 0 1 17190
box 0 0 1 1
use contact_29  contact_29_132
timestamp 1707688321
transform 1 0 5555 0 1 13240
box 0 0 1 1
use contact_29  contact_29_133
timestamp 1707688321
transform 1 0 5555 0 1 14030
box 0 0 1 1
use contact_29  contact_29_134
timestamp 1707688321
transform 1 0 5555 0 1 15206
box 0 0 1 1
use contact_29  contact_29_135
timestamp 1707688321
transform 1 0 5555 0 1 18366
box 0 0 1 1
use contact_29  contact_29_136
timestamp 1707688321
transform 1 0 5555 0 1 14820
box 0 0 1 1
use contact_29  contact_29_137
timestamp 1707688321
transform 1 0 5555 0 1 16400
box 0 0 1 1
use contact_29  contact_29_138
timestamp 1707688321
transform 1 0 5555 0 1 17980
box 0 0 1 1
use contact_29  contact_29_139
timestamp 1707688321
transform 1 0 5555 0 1 13626
box 0 0 1 1
use contact_29  contact_29_140
timestamp 1707688321
transform 1 0 5555 0 1 14416
box 0 0 1 1
use contact_29  contact_29_141
timestamp 1707688321
transform 1 0 5555 0 1 17576
box 0 0 1 1
use contact_29  contact_29_142
timestamp 1707688321
transform 1 0 5555 0 1 12836
box 0 0 1 1
use contact_29  contact_29_143
timestamp 1707688321
transform 1 0 5555 0 1 16786
box 0 0 1 1
use contact_29  contact_29_144
timestamp 1707688321
transform 1 0 5555 0 1 21930
box 0 0 1 1
use contact_29  contact_29_145
timestamp 1707688321
transform 1 0 5555 0 1 23510
box 0 0 1 1
use contact_29  contact_29_146
timestamp 1707688321
transform 1 0 5555 0 1 22720
box 0 0 1 1
use contact_29  contact_29_147
timestamp 1707688321
transform 1 0 5555 0 1 23896
box 0 0 1 1
use contact_29  contact_29_148
timestamp 1707688321
transform 1 0 5555 0 1 25090
box 0 0 1 1
use contact_29  contact_29_149
timestamp 1707688321
transform 1 0 5555 0 1 21526
box 0 0 1 1
use contact_29  contact_29_150
timestamp 1707688321
transform 1 0 5555 0 1 21140
box 0 0 1 1
use contact_29  contact_29_151
timestamp 1707688321
transform 1 0 5555 0 1 20736
box 0 0 1 1
use contact_29  contact_29_152
timestamp 1707688321
transform 1 0 5555 0 1 23106
box 0 0 1 1
use contact_29  contact_29_153
timestamp 1707688321
transform 1 0 5555 0 1 20350
box 0 0 1 1
use contact_29  contact_29_154
timestamp 1707688321
transform 1 0 5555 0 1 19946
box 0 0 1 1
use contact_29  contact_29_155
timestamp 1707688321
transform 1 0 5555 0 1 24686
box 0 0 1 1
use contact_29  contact_29_156
timestamp 1707688321
transform 1 0 5555 0 1 19560
box 0 0 1 1
use contact_29  contact_29_157
timestamp 1707688321
transform 1 0 5555 0 1 19156
box 0 0 1 1
use contact_29  contact_29_158
timestamp 1707688321
transform 1 0 5555 0 1 22316
box 0 0 1 1
use contact_29  contact_29_159
timestamp 1707688321
transform 1 0 5555 0 1 24300
box 0 0 1 1
use contact_29  contact_29_160
timestamp 1707688321
transform 1 0 5665 0 1 21616
box 0 0 1 1
use contact_29  contact_29_161
timestamp 1707688321
transform 1 0 5665 0 1 21414
box 0 0 1 1
use contact_29  contact_29_162
timestamp 1707688321
transform 1 0 5665 0 1 21050
box 0 0 1 1
use contact_29  contact_29_163
timestamp 1707688321
transform 1 0 5665 0 1 21252
box 0 0 1 1
use contact_29  contact_29_164
timestamp 1707688321
transform 1 0 5665 0 1 20826
box 0 0 1 1
use contact_29  contact_29_165
timestamp 1707688321
transform 1 0 5665 0 1 20624
box 0 0 1 1
use contact_29  contact_29_166
timestamp 1707688321
transform 1 0 5665 0 1 20260
box 0 0 1 1
use contact_29  contact_29_167
timestamp 1707688321
transform 1 0 5665 0 1 20462
box 0 0 1 1
use contact_29  contact_29_168
timestamp 1707688321
transform 1 0 5665 0 1 20036
box 0 0 1 1
use contact_29  contact_29_169
timestamp 1707688321
transform 1 0 5665 0 1 19834
box 0 0 1 1
use contact_29  contact_29_170
timestamp 1707688321
transform 1 0 5665 0 1 19470
box 0 0 1 1
use contact_29  contact_29_171
timestamp 1707688321
transform 1 0 5665 0 1 19672
box 0 0 1 1
use contact_29  contact_29_172
timestamp 1707688321
transform 1 0 5665 0 1 19246
box 0 0 1 1
use contact_29  contact_29_173
timestamp 1707688321
transform 1 0 5665 0 1 19044
box 0 0 1 1
use contact_29  contact_29_174
timestamp 1707688321
transform 1 0 5665 0 1 21840
box 0 0 1 1
use contact_29  contact_29_175
timestamp 1707688321
transform 1 0 5665 0 1 22042
box 0 0 1 1
use contact_29  contact_29_176
timestamp 1707688321
transform 1 0 5665 0 1 25000
box 0 0 1 1
use contact_29  contact_29_177
timestamp 1707688321
transform 1 0 5665 0 1 25202
box 0 0 1 1
use contact_29  contact_29_178
timestamp 1707688321
transform 1 0 5665 0 1 24776
box 0 0 1 1
use contact_29  contact_29_179
timestamp 1707688321
transform 1 0 5665 0 1 24574
box 0 0 1 1
use contact_29  contact_29_180
timestamp 1707688321
transform 1 0 5665 0 1 24210
box 0 0 1 1
use contact_29  contact_29_181
timestamp 1707688321
transform 1 0 5665 0 1 24412
box 0 0 1 1
use contact_29  contact_29_182
timestamp 1707688321
transform 1 0 5665 0 1 23986
box 0 0 1 1
use contact_29  contact_29_183
timestamp 1707688321
transform 1 0 5665 0 1 23784
box 0 0 1 1
use contact_29  contact_29_184
timestamp 1707688321
transform 1 0 5665 0 1 23420
box 0 0 1 1
use contact_29  contact_29_185
timestamp 1707688321
transform 1 0 5665 0 1 23622
box 0 0 1 1
use contact_29  contact_29_186
timestamp 1707688321
transform 1 0 5665 0 1 23196
box 0 0 1 1
use contact_29  contact_29_187
timestamp 1707688321
transform 1 0 5665 0 1 22994
box 0 0 1 1
use contact_29  contact_29_188
timestamp 1707688321
transform 1 0 5665 0 1 22630
box 0 0 1 1
use contact_29  contact_29_189
timestamp 1707688321
transform 1 0 5665 0 1 22832
box 0 0 1 1
use contact_29  contact_29_190
timestamp 1707688321
transform 1 0 5665 0 1 22406
box 0 0 1 1
use contact_29  contact_29_191
timestamp 1707688321
transform 1 0 5665 0 1 22204
box 0 0 1 1
use contact_29  contact_29_192
timestamp 1707688321
transform 1 0 5665 0 1 26580
box 0 0 1 1
use contact_29  contact_29_193
timestamp 1707688321
transform 1 0 5665 0 1 27936
box 0 0 1 1
use contact_29  contact_29_194
timestamp 1707688321
transform 1 0 5665 0 1 25992
box 0 0 1 1
use contact_29  contact_29_195
timestamp 1707688321
transform 1 0 5665 0 1 26944
box 0 0 1 1
use contact_29  contact_29_196
timestamp 1707688321
transform 1 0 5665 0 1 27146
box 0 0 1 1
use contact_29  contact_29_197
timestamp 1707688321
transform 1 0 5665 0 1 25790
box 0 0 1 1
use contact_29  contact_29_198
timestamp 1707688321
transform 1 0 5665 0 1 27734
box 0 0 1 1
use contact_29  contact_29_199
timestamp 1707688321
transform 1 0 5665 0 1 26154
box 0 0 1 1
use contact_29  contact_29_200
timestamp 1707688321
transform 1 0 5665 0 1 25566
box 0 0 1 1
use contact_29  contact_29_201
timestamp 1707688321
transform 1 0 5665 0 1 27370
box 0 0 1 1
use contact_29  contact_29_202
timestamp 1707688321
transform 1 0 5665 0 1 26782
box 0 0 1 1
use contact_29  contact_29_203
timestamp 1707688321
transform 1 0 5665 0 1 28362
box 0 0 1 1
use contact_29  contact_29_204
timestamp 1707688321
transform 1 0 5665 0 1 26356
box 0 0 1 1
use contact_29  contact_29_205
timestamp 1707688321
transform 1 0 5665 0 1 27572
box 0 0 1 1
use contact_29  contact_29_206
timestamp 1707688321
transform 1 0 5665 0 1 25364
box 0 0 1 1
use contact_29  contact_29_207
timestamp 1707688321
transform 1 0 5665 0 1 28160
box 0 0 1 1
use contact_29  contact_29_208
timestamp 1707688321
transform 1 0 5665 0 1 30104
box 0 0 1 1
use contact_29  contact_29_209
timestamp 1707688321
transform 1 0 5665 0 1 29740
box 0 0 1 1
use contact_29  contact_29_210
timestamp 1707688321
transform 1 0 5665 0 1 29942
box 0 0 1 1
use contact_29  contact_29_211
timestamp 1707688321
transform 1 0 5665 0 1 29516
box 0 0 1 1
use contact_29  contact_29_212
timestamp 1707688321
transform 1 0 5665 0 1 29314
box 0 0 1 1
use contact_29  contact_29_213
timestamp 1707688321
transform 1 0 5665 0 1 28950
box 0 0 1 1
use contact_29  contact_29_214
timestamp 1707688321
transform 1 0 5665 0 1 30306
box 0 0 1 1
use contact_29  contact_29_215
timestamp 1707688321
transform 1 0 5665 0 1 29152
box 0 0 1 1
use contact_29  contact_29_216
timestamp 1707688321
transform 1 0 5665 0 1 28726
box 0 0 1 1
use contact_29  contact_29_217
timestamp 1707688321
transform 1 0 5665 0 1 31320
box 0 0 1 1
use contact_29  contact_29_218
timestamp 1707688321
transform 1 0 5665 0 1 31522
box 0 0 1 1
use contact_29  contact_29_219
timestamp 1707688321
transform 1 0 5665 0 1 31096
box 0 0 1 1
use contact_29  contact_29_220
timestamp 1707688321
transform 1 0 5665 0 1 28524
box 0 0 1 1
use contact_29  contact_29_221
timestamp 1707688321
transform 1 0 5665 0 1 30894
box 0 0 1 1
use contact_29  contact_29_222
timestamp 1707688321
transform 1 0 5665 0 1 30530
box 0 0 1 1
use contact_29  contact_29_223
timestamp 1707688321
transform 1 0 5665 0 1 30732
box 0 0 1 1
use contact_29  contact_29_224
timestamp 1707688321
transform 1 0 5555 0 1 30620
box 0 0 1 1
use contact_29  contact_29_225
timestamp 1707688321
transform 1 0 5555 0 1 30216
box 0 0 1 1
use contact_29  contact_29_226
timestamp 1707688321
transform 1 0 5555 0 1 25880
box 0 0 1 1
use contact_29  contact_29_227
timestamp 1707688321
transform 1 0 5555 0 1 29830
box 0 0 1 1
use contact_29  contact_29_228
timestamp 1707688321
transform 1 0 5555 0 1 29426
box 0 0 1 1
use contact_29  contact_29_229
timestamp 1707688321
transform 1 0 5555 0 1 26670
box 0 0 1 1
use contact_29  contact_29_230
timestamp 1707688321
transform 1 0 5555 0 1 29040
box 0 0 1 1
use contact_29  contact_29_231
timestamp 1707688321
transform 1 0 5555 0 1 28636
box 0 0 1 1
use contact_29  contact_29_232
timestamp 1707688321
transform 1 0 5555 0 1 28250
box 0 0 1 1
use contact_29  contact_29_233
timestamp 1707688321
transform 1 0 5555 0 1 25476
box 0 0 1 1
use contact_29  contact_29_234
timestamp 1707688321
transform 1 0 5555 0 1 27846
box 0 0 1 1
use contact_29  contact_29_235
timestamp 1707688321
transform 1 0 5555 0 1 26266
box 0 0 1 1
use contact_29  contact_29_236
timestamp 1707688321
transform 1 0 5555 0 1 27460
box 0 0 1 1
use contact_29  contact_29_237
timestamp 1707688321
transform 1 0 5555 0 1 31410
box 0 0 1 1
use contact_29  contact_29_238
timestamp 1707688321
transform 1 0 5555 0 1 27056
box 0 0 1 1
use contact_29  contact_29_239
timestamp 1707688321
transform 1 0 5555 0 1 31006
box 0 0 1 1
use contact_29  contact_29_240
timestamp 1707688321
transform 1 0 5555 0 1 35746
box 0 0 1 1
use contact_29  contact_29_241
timestamp 1707688321
transform 1 0 5555 0 1 35360
box 0 0 1 1
use contact_29  contact_29_242
timestamp 1707688321
transform 1 0 5555 0 1 34956
box 0 0 1 1
use contact_29  contact_29_243
timestamp 1707688321
transform 1 0 5555 0 1 34570
box 0 0 1 1
use contact_29  contact_29_244
timestamp 1707688321
transform 1 0 5555 0 1 34166
box 0 0 1 1
use contact_29  contact_29_245
timestamp 1707688321
transform 1 0 5555 0 1 36536
box 0 0 1 1
use contact_29  contact_29_246
timestamp 1707688321
transform 1 0 5555 0 1 33780
box 0 0 1 1
use contact_29  contact_29_247
timestamp 1707688321
transform 1 0 5555 0 1 33376
box 0 0 1 1
use contact_29  contact_29_248
timestamp 1707688321
transform 1 0 5555 0 1 32990
box 0 0 1 1
use contact_29  contact_29_249
timestamp 1707688321
transform 1 0 5555 0 1 32586
box 0 0 1 1
use contact_29  contact_29_250
timestamp 1707688321
transform 1 0 5555 0 1 32200
box 0 0 1 1
use contact_29  contact_29_251
timestamp 1707688321
transform 1 0 5555 0 1 31796
box 0 0 1 1
use contact_29  contact_29_252
timestamp 1707688321
transform 1 0 5555 0 1 36150
box 0 0 1 1
use contact_29  contact_29_253
timestamp 1707688321
transform 1 0 5555 0 1 37730
box 0 0 1 1
use contact_29  contact_29_254
timestamp 1707688321
transform 1 0 5555 0 1 37326
box 0 0 1 1
use contact_29  contact_29_255
timestamp 1707688321
transform 1 0 5555 0 1 36940
box 0 0 1 1
use contact_29  contact_29_256
timestamp 1707688321
transform 1 0 5665 0 1 34054
box 0 0 1 1
use contact_29  contact_29_257
timestamp 1707688321
transform 1 0 5665 0 1 33690
box 0 0 1 1
use contact_29  contact_29_258
timestamp 1707688321
transform 1 0 5665 0 1 33892
box 0 0 1 1
use contact_29  contact_29_259
timestamp 1707688321
transform 1 0 5665 0 1 33466
box 0 0 1 1
use contact_29  contact_29_260
timestamp 1707688321
transform 1 0 5665 0 1 33264
box 0 0 1 1
use contact_29  contact_29_261
timestamp 1707688321
transform 1 0 5665 0 1 32900
box 0 0 1 1
use contact_29  contact_29_262
timestamp 1707688321
transform 1 0 5665 0 1 33102
box 0 0 1 1
use contact_29  contact_29_263
timestamp 1707688321
transform 1 0 5665 0 1 32676
box 0 0 1 1
use contact_29  contact_29_264
timestamp 1707688321
transform 1 0 5665 0 1 32474
box 0 0 1 1
use contact_29  contact_29_265
timestamp 1707688321
transform 1 0 5665 0 1 32110
box 0 0 1 1
use contact_29  contact_29_266
timestamp 1707688321
transform 1 0 5665 0 1 34682
box 0 0 1 1
use contact_29  contact_29_267
timestamp 1707688321
transform 1 0 5665 0 1 32312
box 0 0 1 1
use contact_29  contact_29_268
timestamp 1707688321
transform 1 0 5665 0 1 31886
box 0 0 1 1
use contact_29  contact_29_269
timestamp 1707688321
transform 1 0 5665 0 1 34256
box 0 0 1 1
use contact_29  contact_29_270
timestamp 1707688321
transform 1 0 5665 0 1 31684
box 0 0 1 1
use contact_29  contact_29_271
timestamp 1707688321
transform 1 0 5665 0 1 34480
box 0 0 1 1
use contact_29  contact_29_272
timestamp 1707688321
transform 1 0 5665 0 1 37640
box 0 0 1 1
use contact_29  contact_29_273
timestamp 1707688321
transform 1 0 5665 0 1 37842
box 0 0 1 1
use contact_29  contact_29_274
timestamp 1707688321
transform 1 0 5665 0 1 37416
box 0 0 1 1
use contact_29  contact_29_275
timestamp 1707688321
transform 1 0 5665 0 1 37214
box 0 0 1 1
use contact_29  contact_29_276
timestamp 1707688321
transform 1 0 5665 0 1 36850
box 0 0 1 1
use contact_29  contact_29_277
timestamp 1707688321
transform 1 0 5665 0 1 37052
box 0 0 1 1
use contact_29  contact_29_278
timestamp 1707688321
transform 1 0 5665 0 1 36626
box 0 0 1 1
use contact_29  contact_29_279
timestamp 1707688321
transform 1 0 5665 0 1 36424
box 0 0 1 1
use contact_29  contact_29_280
timestamp 1707688321
transform 1 0 5665 0 1 36060
box 0 0 1 1
use contact_29  contact_29_281
timestamp 1707688321
transform 1 0 5665 0 1 36262
box 0 0 1 1
use contact_29  contact_29_282
timestamp 1707688321
transform 1 0 5665 0 1 35836
box 0 0 1 1
use contact_29  contact_29_283
timestamp 1707688321
transform 1 0 5665 0 1 35634
box 0 0 1 1
use contact_29  contact_29_284
timestamp 1707688321
transform 1 0 5665 0 1 35270
box 0 0 1 1
use contact_29  contact_29_285
timestamp 1707688321
transform 1 0 5665 0 1 35472
box 0 0 1 1
use contact_29  contact_29_286
timestamp 1707688321
transform 1 0 5665 0 1 35046
box 0 0 1 1
use contact_29  contact_29_287
timestamp 1707688321
transform 1 0 5665 0 1 34844
box 0 0 1 1
use contact_29  contact_29_288
timestamp 1707688321
transform 1 0 5665 0 1 40010
box 0 0 1 1
use contact_29  contact_29_289
timestamp 1707688321
transform 1 0 5665 0 1 40212
box 0 0 1 1
use contact_29  contact_29_290
timestamp 1707688321
transform 1 0 5665 0 1 39786
box 0 0 1 1
use contact_29  contact_29_291
timestamp 1707688321
transform 1 0 5665 0 1 39584
box 0 0 1 1
use contact_29  contact_29_292
timestamp 1707688321
transform 1 0 5665 0 1 39220
box 0 0 1 1
use contact_29  contact_29_293
timestamp 1707688321
transform 1 0 5665 0 1 39422
box 0 0 1 1
use contact_29  contact_29_294
timestamp 1707688321
transform 1 0 5665 0 1 38996
box 0 0 1 1
use contact_29  contact_29_295
timestamp 1707688321
transform 1 0 5665 0 1 38794
box 0 0 1 1
use contact_29  contact_29_296
timestamp 1707688321
transform 1 0 5665 0 1 38430
box 0 0 1 1
use contact_29  contact_29_297
timestamp 1707688321
transform 1 0 5665 0 1 38632
box 0 0 1 1
use contact_29  contact_29_298
timestamp 1707688321
transform 1 0 5665 0 1 38206
box 0 0 1 1
use contact_29  contact_29_299
timestamp 1707688321
transform 1 0 5665 0 1 38004
box 0 0 1 1
use contact_29  contact_29_300
timestamp 1707688321
transform 1 0 5665 0 1 40800
box 0 0 1 1
use contact_29  contact_29_301
timestamp 1707688321
transform 1 0 5665 0 1 41002
box 0 0 1 1
use contact_29  contact_29_302
timestamp 1707688321
transform 1 0 5665 0 1 40576
box 0 0 1 1
use contact_29  contact_29_303
timestamp 1707688321
transform 1 0 5665 0 1 40374
box 0 0 1 1
use contact_29  contact_29_304
timestamp 1707688321
transform 1 0 5665 0 1 43170
box 0 0 1 1
use contact_29  contact_29_305
timestamp 1707688321
transform 1 0 5665 0 1 43372
box 0 0 1 1
use contact_29  contact_29_306
timestamp 1707688321
transform 1 0 5665 0 1 42946
box 0 0 1 1
use contact_29  contact_29_307
timestamp 1707688321
transform 1 0 5665 0 1 42744
box 0 0 1 1
use contact_29  contact_29_308
timestamp 1707688321
transform 1 0 5665 0 1 42380
box 0 0 1 1
use contact_29  contact_29_309
timestamp 1707688321
transform 1 0 5665 0 1 42582
box 0 0 1 1
use contact_29  contact_29_310
timestamp 1707688321
transform 1 0 5665 0 1 42156
box 0 0 1 1
use contact_29  contact_29_311
timestamp 1707688321
transform 1 0 5665 0 1 41954
box 0 0 1 1
use contact_29  contact_29_312
timestamp 1707688321
transform 1 0 5665 0 1 41590
box 0 0 1 1
use contact_29  contact_29_313
timestamp 1707688321
transform 1 0 5665 0 1 41792
box 0 0 1 1
use contact_29  contact_29_314
timestamp 1707688321
transform 1 0 5665 0 1 41366
box 0 0 1 1
use contact_29  contact_29_315
timestamp 1707688321
transform 1 0 5665 0 1 41164
box 0 0 1 1
use contact_29  contact_29_316
timestamp 1707688321
transform 1 0 5665 0 1 43960
box 0 0 1 1
use contact_29  contact_29_317
timestamp 1707688321
transform 1 0 5665 0 1 44162
box 0 0 1 1
use contact_29  contact_29_318
timestamp 1707688321
transform 1 0 5665 0 1 43736
box 0 0 1 1
use contact_29  contact_29_319
timestamp 1707688321
transform 1 0 5665 0 1 43534
box 0 0 1 1
use contact_29  contact_29_320
timestamp 1707688321
transform 1 0 5555 0 1 40486
box 0 0 1 1
use contact_29  contact_29_321
timestamp 1707688321
transform 1 0 5555 0 1 43646
box 0 0 1 1
use contact_29  contact_29_322
timestamp 1707688321
transform 1 0 5555 0 1 38520
box 0 0 1 1
use contact_29  contact_29_323
timestamp 1707688321
transform 1 0 5555 0 1 42470
box 0 0 1 1
use contact_29  contact_29_324
timestamp 1707688321
transform 1 0 5555 0 1 38116
box 0 0 1 1
use contact_29  contact_29_325
timestamp 1707688321
transform 1 0 5555 0 1 43260
box 0 0 1 1
use contact_29  contact_29_326
timestamp 1707688321
transform 1 0 5555 0 1 41680
box 0 0 1 1
use contact_29  contact_29_327
timestamp 1707688321
transform 1 0 5555 0 1 41276
box 0 0 1 1
use contact_29  contact_29_328
timestamp 1707688321
transform 1 0 5555 0 1 38906
box 0 0 1 1
use contact_29  contact_29_329
timestamp 1707688321
transform 1 0 5555 0 1 44050
box 0 0 1 1
use contact_29  contact_29_330
timestamp 1707688321
transform 1 0 5555 0 1 40100
box 0 0 1 1
use contact_29  contact_29_331
timestamp 1707688321
transform 1 0 5555 0 1 42856
box 0 0 1 1
use contact_29  contact_29_332
timestamp 1707688321
transform 1 0 5555 0 1 42066
box 0 0 1 1
use contact_29  contact_29_333
timestamp 1707688321
transform 1 0 5555 0 1 40890
box 0 0 1 1
use contact_29  contact_29_334
timestamp 1707688321
transform 1 0 5555 0 1 39310
box 0 0 1 1
use contact_29  contact_29_335
timestamp 1707688321
transform 1 0 5555 0 1 39696
box 0 0 1 1
use contact_29  contact_29_336
timestamp 1707688321
transform 1 0 5555 0 1 50370
box 0 0 1 1
use contact_29  contact_29_337
timestamp 1707688321
transform 1 0 5555 0 1 49966
box 0 0 1 1
use contact_29  contact_29_338
timestamp 1707688321
transform 1 0 5555 0 1 49580
box 0 0 1 1
use contact_29  contact_29_339
timestamp 1707688321
transform 1 0 5555 0 1 49176
box 0 0 1 1
use contact_29  contact_29_340
timestamp 1707688321
transform 1 0 5555 0 1 48790
box 0 0 1 1
use contact_29  contact_29_341
timestamp 1707688321
transform 1 0 5555 0 1 48386
box 0 0 1 1
use contact_29  contact_29_342
timestamp 1707688321
transform 1 0 5555 0 1 48000
box 0 0 1 1
use contact_29  contact_29_343
timestamp 1707688321
transform 1 0 5555 0 1 47596
box 0 0 1 1
use contact_29  contact_29_344
timestamp 1707688321
transform 1 0 5555 0 1 47210
box 0 0 1 1
use contact_29  contact_29_345
timestamp 1707688321
transform 1 0 5555 0 1 44840
box 0 0 1 1
use contact_29  contact_29_346
timestamp 1707688321
transform 1 0 5555 0 1 46806
box 0 0 1 1
use contact_29  contact_29_347
timestamp 1707688321
transform 1 0 5555 0 1 46420
box 0 0 1 1
use contact_29  contact_29_348
timestamp 1707688321
transform 1 0 5555 0 1 46016
box 0 0 1 1
use contact_29  contact_29_349
timestamp 1707688321
transform 1 0 5555 0 1 44436
box 0 0 1 1
use contact_29  contact_29_350
timestamp 1707688321
transform 1 0 5555 0 1 45630
box 0 0 1 1
use contact_29  contact_29_351
timestamp 1707688321
transform 1 0 5555 0 1 45226
box 0 0 1 1
use contact_29  contact_29_352
timestamp 1707688321
transform 1 0 5665 0 1 46106
box 0 0 1 1
use contact_29  contact_29_353
timestamp 1707688321
transform 1 0 5665 0 1 45904
box 0 0 1 1
use contact_29  contact_29_354
timestamp 1707688321
transform 1 0 5665 0 1 45316
box 0 0 1 1
use contact_29  contact_29_355
timestamp 1707688321
transform 1 0 5665 0 1 45114
box 0 0 1 1
use contact_29  contact_29_356
timestamp 1707688321
transform 1 0 5665 0 1 46896
box 0 0 1 1
use contact_29  contact_29_357
timestamp 1707688321
transform 1 0 5665 0 1 46694
box 0 0 1 1
use contact_29  contact_29_358
timestamp 1707688321
transform 1 0 5665 0 1 45540
box 0 0 1 1
use contact_29  contact_29_359
timestamp 1707688321
transform 1 0 5665 0 1 45742
box 0 0 1 1
use contact_29  contact_29_360
timestamp 1707688321
transform 1 0 5665 0 1 44750
box 0 0 1 1
use contact_29  contact_29_361
timestamp 1707688321
transform 1 0 5665 0 1 44952
box 0 0 1 1
use contact_29  contact_29_362
timestamp 1707688321
transform 1 0 5665 0 1 44526
box 0 0 1 1
use contact_29  contact_29_363
timestamp 1707688321
transform 1 0 5665 0 1 44324
box 0 0 1 1
use contact_29  contact_29_364
timestamp 1707688321
transform 1 0 5665 0 1 46330
box 0 0 1 1
use contact_29  contact_29_365
timestamp 1707688321
transform 1 0 5665 0 1 46532
box 0 0 1 1
use contact_29  contact_29_366
timestamp 1707688321
transform 1 0 5665 0 1 47120
box 0 0 1 1
use contact_29  contact_29_367
timestamp 1707688321
transform 1 0 5665 0 1 47322
box 0 0 1 1
use contact_29  contact_29_368
timestamp 1707688321
transform 1 0 5665 0 1 48476
box 0 0 1 1
use contact_29  contact_29_369
timestamp 1707688321
transform 1 0 5665 0 1 48274
box 0 0 1 1
use contact_29  contact_29_370
timestamp 1707688321
transform 1 0 5665 0 1 47686
box 0 0 1 1
use contact_29  contact_29_371
timestamp 1707688321
transform 1 0 5665 0 1 47484
box 0 0 1 1
use contact_29  contact_29_372
timestamp 1707688321
transform 1 0 5665 0 1 47910
box 0 0 1 1
use contact_29  contact_29_373
timestamp 1707688321
transform 1 0 5665 0 1 48112
box 0 0 1 1
use contact_29  contact_29_374
timestamp 1707688321
transform 1 0 5665 0 1 50280
box 0 0 1 1
use contact_29  contact_29_375
timestamp 1707688321
transform 1 0 5665 0 1 50482
box 0 0 1 1
use contact_29  contact_29_376
timestamp 1707688321
transform 1 0 5665 0 1 50056
box 0 0 1 1
use contact_29  contact_29_377
timestamp 1707688321
transform 1 0 5665 0 1 49854
box 0 0 1 1
use contact_29  contact_29_378
timestamp 1707688321
transform 1 0 5665 0 1 49490
box 0 0 1 1
use contact_29  contact_29_379
timestamp 1707688321
transform 1 0 5665 0 1 49692
box 0 0 1 1
use contact_29  contact_29_380
timestamp 1707688321
transform 1 0 5665 0 1 49266
box 0 0 1 1
use contact_29  contact_29_381
timestamp 1707688321
transform 1 0 5665 0 1 49064
box 0 0 1 1
use contact_29  contact_29_382
timestamp 1707688321
transform 1 0 5665 0 1 48700
box 0 0 1 1
use contact_29  contact_29_383
timestamp 1707688321
transform 1 0 5665 0 1 48902
box 0 0 1 1
use hierarchical_predecode2x4  hierarchical_predecode2x4_0
timestamp 1707688321
transform 1 0 1282 0 1 29
box 62 -56 2930 1636
use hierarchical_predecode2x4  hierarchical_predecode2x4_1
timestamp 1707688321
transform 1 0 1282 0 1 2399
box 62 -56 2930 1636
use hierarchical_predecode3x8  hierarchical_predecode3x8_0
timestamp 1707688321
transform 1 0 606 0 1 4769
box 62 -60 3606 3220
<< labels >>
rlabel locali s 7257 31776 7257 31776 4 decode_80
port 88 nsew
rlabel locali s 7257 38096 7257 38096 4 decode_96
port 104 nsew
rlabel locali s 7257 49946 7257 49946 4 decode_126
port 134 nsew
rlabel locali s 7257 34146 7257 34146 4 decode_86
port 94 nsew
rlabel locali s 7257 41256 7257 41256 4 decode_104
port 112 nsew
rlabel locali s 7257 27036 7257 27036 4 decode_68
port 76 nsew
rlabel locali s 7257 48862 7257 48862 4 decode_123
port 131 nsew
rlabel locali s 7257 25456 7257 25456 4 decode_64
port 72 nsew
rlabel locali s 7257 30196 7257 30196 4 decode_76
port 84 nsew
rlabel locali s 7257 40962 7257 40962 4 decode_103
port 111 nsew
rlabel locali s 7257 26246 7257 26246 4 decode_66
port 74 nsew
rlabel locali s 7257 36516 7257 36516 4 decode_92
port 100 nsew
rlabel locali s 7257 48072 7257 48072 4 decode_121
port 129 nsew
rlabel locali s 7257 35432 7257 35432 4 decode_89
port 97 nsew
rlabel locali s 7257 25952 7257 25952 4 decode_65
port 73 nsew
rlabel locali s 7257 38592 7257 38592 4 decode_97
port 105 nsew
rlabel locali s 7257 31482 7257 31482 4 decode_79
port 87 nsew
rlabel locali s 7257 38886 7257 38886 4 decode_98
port 106 nsew
rlabel locali s 7257 36222 7257 36222 4 decode_91
port 99 nsew
rlabel locali s 7257 35726 7257 35726 4 decode_90
port 98 nsew
rlabel locali s 7257 49156 7257 49156 4 decode_124
port 132 nsew
rlabel locali s 7257 46492 7257 46492 4 decode_117
port 125 nsew
rlabel locali s 7257 44912 7257 44912 4 decode_113
port 121 nsew
rlabel locali s 7257 29112 7257 29112 4 decode_73
port 81 nsew
rlabel locali s 7257 50442 7257 50442 4 decode_127
port 135 nsew
rlabel locali s 7257 30986 7257 30986 4 decode_78
port 86 nsew
rlabel locali s 7257 32272 7257 32272 4 decode_81
port 89 nsew
rlabel locali s 7257 39676 7257 39676 4 decode_100
port 108 nsew
rlabel locali s 7257 29406 7257 29406 4 decode_74
port 82 nsew
rlabel locali s 7257 40466 7257 40466 4 decode_102
port 110 nsew
rlabel locali s 7257 42542 7257 42542 4 decode_107
port 115 nsew
rlabel locali s 7257 43626 7257 43626 4 decode_110
port 118 nsew
rlabel locali s 7257 45702 7257 45702 4 decode_115
port 123 nsew
rlabel locali s 7257 27532 7257 27532 4 decode_69
port 77 nsew
rlabel locali s 7257 29902 7257 29902 4 decode_75
port 83 nsew
rlabel locali s 7257 48366 7257 48366 4 decode_122
port 130 nsew
rlabel locali s 7257 45206 7257 45206 4 decode_114
port 122 nsew
rlabel locali s 7257 32566 7257 32566 4 decode_82
port 90 nsew
rlabel locali s 7257 42046 7257 42046 4 decode_106
port 114 nsew
rlabel locali s 7257 34936 7257 34936 4 decode_88
port 96 nsew
rlabel locali s 7257 41752 7257 41752 4 decode_105
port 113 nsew
rlabel locali s 7257 47576 7257 47576 4 decode_120
port 128 nsew
rlabel locali s 7257 33356 7257 33356 4 decode_84
port 92 nsew
rlabel locali s 7257 30692 7257 30692 4 decode_77
port 85 nsew
rlabel locali s 7257 33852 7257 33852 4 decode_85
port 93 nsew
rlabel locali s 7257 42836 7257 42836 4 decode_108
port 116 nsew
rlabel locali s 7257 44122 7257 44122 4 decode_111
port 119 nsew
rlabel locali s 7257 39382 7257 39382 4 decode_99
port 107 nsew
rlabel locali s 7257 34642 7257 34642 4 decode_87
port 95 nsew
rlabel locali s 7257 28322 7257 28322 4 decode_71
port 79 nsew
rlabel locali s 7257 37306 7257 37306 4 decode_94
port 102 nsew
rlabel locali s 7257 33062 7257 33062 4 decode_83
port 91 nsew
rlabel locali s 7257 40172 7257 40172 4 decode_101
port 109 nsew
rlabel locali s 7257 27826 7257 27826 4 decode_70
port 78 nsew
rlabel locali s 7257 37012 7257 37012 4 decode_93
port 101 nsew
rlabel locali s 7257 46786 7257 46786 4 decode_118
port 126 nsew
rlabel locali s 7257 26742 7257 26742 4 decode_67
port 75 nsew
rlabel locali s 7257 49652 7257 49652 4 decode_125
port 133 nsew
rlabel locali s 7257 45996 7257 45996 4 decode_116
port 124 nsew
rlabel locali s 7257 44416 7257 44416 4 decode_112
port 120 nsew
rlabel locali s 7257 28616 7257 28616 4 decode_72
port 80 nsew
rlabel locali s 7257 43332 7257 43332 4 decode_109
port 117 nsew
rlabel locali s 7257 47282 7257 47282 4 decode_119
port 127 nsew
rlabel locali s 7257 37802 7257 37802 4 decode_95
port 103 nsew
rlabel locali s 7257 14102 7257 14102 4 decode_35
port 43 nsew
rlabel locali s 7257 16472 7257 16472 4 decode_41
port 49 nsew
rlabel locali s 7257 2546 7257 2546 4 decode_6
port 14 nsew
rlabel locali s 7257 10446 7257 10446 4 decode_26
port 34 nsew
rlabel locali s 7257 966 7257 966 4 decode_2
port 10 nsew
rlabel locali s 7257 3042 7257 3042 4 decode_7
port 15 nsew
rlabel locali s 7257 12816 7257 12816 4 decode_32
port 40 nsew
rlabel locali s 7257 19926 7257 19926 4 decode_50
port 58 nsew
rlabel locali s 7257 18842 7257 18842 4 decode_47
port 55 nsew
rlabel locali s 7257 15186 7257 15186 4 decode_38
port 46 nsew
rlabel locali s 7257 13606 7257 13606 4 decode_34
port 42 nsew
rlabel locali s 7257 14892 7257 14892 4 decode_37
port 45 nsew
rlabel locali s 7257 4916 7257 4916 4 decode_12
port 20 nsew
rlabel locali s 7257 17556 7257 17556 4 decode_44
port 52 nsew
rlabel locali s 7257 1462 7257 1462 4 decode_3
port 11 nsew
rlabel locali s 7257 22296 7257 22296 4 decode_56
port 64 nsew
rlabel locali s 7257 9656 7257 9656 4 decode_24
port 32 nsew
rlabel locali s 7257 20422 7257 20422 4 decode_51
port 59 nsew
rlabel locali s 7257 9362 7257 9362 4 decode_23
port 31 nsew
rlabel locali s 7257 8572 7257 8572 4 decode_21
port 29 nsew
rlabel locali s 7257 2252 7257 2252 4 decode_5
port 13 nsew
rlabel locali s 7257 15976 7257 15976 4 decode_40
port 48 nsew
rlabel locali s 7257 14396 7257 14396 4 decode_36
port 44 nsew
rlabel locali s 7257 13312 7257 13312 4 decode_33
port 41 nsew
rlabel locali s 7257 25162 7257 25162 4 decode_63
port 71 nsew
rlabel locali s 7257 23876 7257 23876 4 decode_60
port 68 nsew
rlabel locali s 7257 8076 7257 8076 4 decode_20
port 28 nsew
rlabel locali s 7257 24372 7257 24372 4 decode_61
port 69 nsew
rlabel locali s 7257 11732 7257 11732 4 decode_29
port 37 nsew
rlabel locali s 7257 3832 7257 3832 4 decode_9
port 17 nsew
rlabel locali s 7257 5706 7257 5706 4 decode_14
port 22 nsew
rlabel locali s 7257 19136 7257 19136 4 decode_48
port 56 nsew
rlabel locali s 7257 21506 7257 21506 4 decode_54
port 62 nsew
rlabel locali s 7257 6992 7257 6992 4 decode_17
port 25 nsew
rlabel locali s 7257 672 7257 672 4 decode_1
port 9 nsew
rlabel locali s 7257 23086 7257 23086 4 decode_58
port 66 nsew
rlabel locali s 7257 4126 7257 4126 4 decode_10
port 18 nsew
rlabel locali s 7257 22002 7257 22002 4 decode_55
port 63 nsew
rlabel locali s 7257 176 7257 176 4 decode_0
port 8 nsew
rlabel locali s 7257 22792 7257 22792 4 decode_57
port 65 nsew
rlabel locali s 7257 8866 7257 8866 4 decode_22
port 30 nsew
rlabel locali s 7257 19632 7257 19632 4 decode_49
port 57 nsew
rlabel locali s 7257 24666 7257 24666 4 decode_62
port 70 nsew
rlabel locali s 7257 6202 7257 6202 4 decode_15
port 23 nsew
rlabel locali s 7257 7782 7257 7782 4 decode_19
port 27 nsew
rlabel locali s 7257 15682 7257 15682 4 decode_39
port 47 nsew
rlabel locali s 7257 10942 7257 10942 4 decode_27
port 35 nsew
rlabel locali s 7257 12522 7257 12522 4 decode_31
port 39 nsew
rlabel locali s 7257 4622 7257 4622 4 decode_11
port 19 nsew
rlabel locali s 7257 1756 7257 1756 4 decode_4
port 12 nsew
rlabel locali s 7257 10152 7257 10152 4 decode_25
port 33 nsew
rlabel locali s 7257 16766 7257 16766 4 decode_42
port 50 nsew
rlabel locali s 7257 11236 7257 11236 4 decode_28
port 36 nsew
rlabel locali s 7257 7286 7257 7286 4 decode_18
port 26 nsew
rlabel locali s 7257 17262 7257 17262 4 decode_43
port 51 nsew
rlabel locali s 7257 20716 7257 20716 4 decode_52
port 60 nsew
rlabel locali s 7257 21212 7257 21212 4 decode_53
port 61 nsew
rlabel locali s 7257 12026 7257 12026 4 decode_30
port 38 nsew
rlabel locali s 7257 18052 7257 18052 4 decode_45
port 53 nsew
rlabel locali s 7257 23582 7257 23582 4 decode_59
port 67 nsew
rlabel locali s 7257 5412 7257 5412 4 decode_13
port 21 nsew
rlabel locali s 7257 18346 7257 18346 4 decode_46
port 54 nsew
rlabel locali s 7257 6496 7257 6496 4 decode_16
port 24 nsew
rlabel locali s 7257 3336 7257 3336 4 decode_8
port 16 nsew
rlabel metal1 s 4608 25323 4608 25323 4 predecode_4
port 744 nsew
rlabel metal1 s 4688 25323 4688 25323 4 predecode_5
port 745 nsew
rlabel metal1 s 432 3979 432 3979 4 addr_5
port 6 nsew
rlabel metal1 s 4768 25323 4768 25323 4 predecode_6
port 746 nsew
rlabel metal1 s 5008 25323 5008 25323 4 predecode_9
port 747 nsew
rlabel metal1 s 5328 25323 5328 25323 4 predecode_13
port 748 nsew
rlabel metal1 s 4448 25323 4448 25323 4 predecode_2
port 749 nsew
rlabel metal1 s 4288 25323 4288 25323 4 predecode_0
port 750 nsew
rlabel metal1 s 5488 25323 5488 25323 4 predecode_15
port 751 nsew
rlabel metal1 s 4528 25323 4528 25323 4 predecode_3
port 752 nsew
rlabel metal1 s 5088 25323 5088 25323 4 predecode_10
port 753 nsew
rlabel metal1 s 272 3979 272 3979 4 addr_3
port 4 nsew
rlabel metal1 s 4928 25323 4928 25323 4 predecode_8
port 754 nsew
rlabel metal1 s 192 3979 192 3979 4 addr_2
port 3 nsew
rlabel metal1 s 112 3979 112 3979 4 addr_1
port 2 nsew
rlabel metal1 s 352 3979 352 3979 4 addr_4
port 5 nsew
rlabel metal1 s 512 3979 512 3979 4 addr_6
port 7 nsew
rlabel metal1 s 5248 25323 5248 25323 4 predecode_12
port 755 nsew
rlabel metal1 s 5168 25323 5168 25323 4 predecode_11
port 756 nsew
rlabel metal1 s 5408 25323 5408 25323 4 predecode_14
port 757 nsew
rlabel metal1 s 4368 25323 4368 25323 4 predecode_1
port 758 nsew
rlabel metal1 s 32 3979 32 3979 4 addr_0
port 1 nsew
rlabel metal1 s 4848 25323 4848 25323 4 predecode_7
port 743 nsew
rlabel metal3 s 7336 45059 7336 45059 4 vdd
port 136 nsew
rlabel metal3 s 7336 49009 7336 49009 4 vdd
port 136 nsew
rlabel metal3 s 6682 45045 6682 45045 4 vdd
port 136 nsew
rlabel metal3 s 6682 44687 6682 44687 4 vdd
port 136 nsew
rlabel metal3 s 7336 47429 7336 47429 4 vdd
port 136 nsew
rlabel metal3 s 7336 45454 7336 45454 4 vdd
port 136 nsew
rlabel metal3 s 6682 44255 6682 44255 4 vdd
port 136 nsew
rlabel metal3 s 7336 44269 7336 44269 4 vdd
port 136 nsew
rlabel metal3 s 6682 46267 6682 46267 4 vdd
port 136 nsew
rlabel metal3 s 7336 49799 7336 49799 4 vdd
port 136 nsew
rlabel metal3 s 6682 49785 6682 49785 4 vdd
port 136 nsew
rlabel metal3 s 7336 46639 7336 46639 4 vdd
port 136 nsew
rlabel metal3 s 6682 47415 6682 47415 4 vdd
port 136 nsew
rlabel metal3 s 6682 47847 6682 47847 4 vdd
port 136 nsew
rlabel metal3 s 7336 47824 7336 47824 4 vdd
port 136 nsew
rlabel metal3 s 6682 50217 6682 50217 4 vdd
port 136 nsew
rlabel metal3 s 7336 47034 7336 47034 4 vdd
port 136 nsew
rlabel metal3 s 6682 46625 6682 46625 4 vdd
port 136 nsew
rlabel metal3 s 6682 48205 6682 48205 4 vdd
port 136 nsew
rlabel metal3 s 6682 45835 6682 45835 4 vdd
port 136 nsew
rlabel metal3 s 7336 44664 7336 44664 4 vdd
port 136 nsew
rlabel metal3 s 6682 49427 6682 49427 4 vdd
port 136 nsew
rlabel metal3 s 7336 49404 7336 49404 4 vdd
port 136 nsew
rlabel metal3 s 7336 46244 7336 46244 4 vdd
port 136 nsew
rlabel metal3 s 7336 48219 7336 48219 4 vdd
port 136 nsew
rlabel metal3 s 7336 45849 7336 45849 4 vdd
port 136 nsew
rlabel metal3 s 6682 48995 6682 48995 4 vdd
port 136 nsew
rlabel metal3 s 6682 45477 6682 45477 4 vdd
port 136 nsew
rlabel metal3 s 6682 48637 6682 48637 4 vdd
port 136 nsew
rlabel metal3 s 6682 47057 6682 47057 4 vdd
port 136 nsew
rlabel metal3 s 7336 48614 7336 48614 4 vdd
port 136 nsew
rlabel metal3 s 7336 50194 7336 50194 4 vdd
port 136 nsew
rlabel metal3 s 7064 48614 7064 48614 4 gnd
port 137 nsew
rlabel metal3 s 7064 49009 7064 49009 4 gnd
port 137 nsew
rlabel metal3 s 7064 46244 7064 46244 4 gnd
port 137 nsew
rlabel metal3 s 7064 44664 7064 44664 4 gnd
port 137 nsew
rlabel metal3 s 7064 49404 7064 49404 4 gnd
port 137 nsew
rlabel metal3 s 7064 46639 7064 46639 4 gnd
port 137 nsew
rlabel metal3 s 7064 45059 7064 45059 4 gnd
port 137 nsew
rlabel metal3 s 7064 45454 7064 45454 4 gnd
port 137 nsew
rlabel metal3 s 7064 47824 7064 47824 4 gnd
port 137 nsew
rlabel metal3 s 7064 48219 7064 48219 4 gnd
port 137 nsew
rlabel metal3 s 7064 47429 7064 47429 4 gnd
port 137 nsew
rlabel metal3 s 7064 45849 7064 45849 4 gnd
port 137 nsew
rlabel metal3 s 7064 49799 7064 49799 4 gnd
port 137 nsew
rlabel metal3 s 7064 47034 7064 47034 4 gnd
port 137 nsew
rlabel metal3 s 7064 44269 7064 44269 4 gnd
port 137 nsew
rlabel metal3 s 7064 50194 7064 50194 4 gnd
port 137 nsew
rlabel metal3 s 6250 45477 6250 45477 4 vdd
port 136 nsew
rlabel metal3 s 6250 46267 6250 46267 4 vdd
port 136 nsew
rlabel metal3 s 6250 44687 6250 44687 4 vdd
port 136 nsew
rlabel metal3 s 6250 47057 6250 47057 4 vdd
port 136 nsew
rlabel metal3 s 5825 50217 5825 50217 4 gnd
port 137 nsew
rlabel metal3 s 5825 46267 5825 46267 4 gnd
port 137 nsew
rlabel metal3 s 5825 48263 5825 48263 4 gnd
port 137 nsew
rlabel metal3 s 5825 47473 5825 47473 4 gnd
port 137 nsew
rlabel metal3 s 5825 48637 5825 48637 4 gnd
port 137 nsew
rlabel metal3 s 5825 45103 5825 45103 4 gnd
port 137 nsew
rlabel metal3 s 6250 44255 6250 44255 4 vdd
port 136 nsew
rlabel metal3 s 5825 49053 5825 49053 4 gnd
port 137 nsew
rlabel metal3 s 6250 48995 6250 48995 4 vdd
port 136 nsew
rlabel metal3 s 6250 46625 6250 46625 4 vdd
port 136 nsew
rlabel metal3 s 6250 49785 6250 49785 4 vdd
port 136 nsew
rlabel metal3 s 5825 45477 5825 45477 4 gnd
port 137 nsew
rlabel metal3 s 5825 49843 5825 49843 4 gnd
port 137 nsew
rlabel metal3 s 6250 48205 6250 48205 4 vdd
port 136 nsew
rlabel metal3 s 5825 46683 5825 46683 4 gnd
port 137 nsew
rlabel metal3 s 5825 44687 5825 44687 4 gnd
port 137 nsew
rlabel metal3 s 5825 49427 5825 49427 4 gnd
port 137 nsew
rlabel metal3 s 6250 50217 6250 50217 4 vdd
port 136 nsew
rlabel metal3 s 5825 47847 5825 47847 4 gnd
port 137 nsew
rlabel metal3 s 5825 45893 5825 45893 4 gnd
port 137 nsew
rlabel metal3 s 6250 49427 6250 49427 4 vdd
port 136 nsew
rlabel metal3 s 6250 48637 6250 48637 4 vdd
port 136 nsew
rlabel metal3 s 5825 47057 5825 47057 4 gnd
port 137 nsew
rlabel metal3 s 6250 45835 6250 45835 4 vdd
port 136 nsew
rlabel metal3 s 6250 45045 6250 45045 4 vdd
port 136 nsew
rlabel metal3 s 5825 44313 5825 44313 4 gnd
port 137 nsew
rlabel metal3 s 6250 47415 6250 47415 4 vdd
port 136 nsew
rlabel metal3 s 6250 47847 6250 47847 4 vdd
port 136 nsew
rlabel metal3 s 6250 41885 6250 41885 4 vdd
port 136 nsew
rlabel metal3 s 6250 40737 6250 40737 4 vdd
port 136 nsew
rlabel metal3 s 6250 38367 6250 38367 4 vdd
port 136 nsew
rlabel metal3 s 6250 37935 6250 37935 4 vdd
port 136 nsew
rlabel metal3 s 5825 42733 5825 42733 4 gnd
port 137 nsew
rlabel metal3 s 6250 40305 6250 40305 4 vdd
port 136 nsew
rlabel metal3 s 6250 39515 6250 39515 4 vdd
port 136 nsew
rlabel metal3 s 6250 38725 6250 38725 4 vdd
port 136 nsew
rlabel metal3 s 6250 43465 6250 43465 4 vdd
port 136 nsew
rlabel metal3 s 6250 42317 6250 42317 4 vdd
port 136 nsew
rlabel metal3 s 5825 39947 5825 39947 4 gnd
port 137 nsew
rlabel metal3 s 5825 39573 5825 39573 4 gnd
port 137 nsew
rlabel metal3 s 5825 42317 5825 42317 4 gnd
port 137 nsew
rlabel metal3 s 5825 43107 5825 43107 4 gnd
port 137 nsew
rlabel metal3 s 5825 39157 5825 39157 4 gnd
port 137 nsew
rlabel metal3 s 6250 41527 6250 41527 4 vdd
port 136 nsew
rlabel metal3 s 5825 41527 5825 41527 4 gnd
port 137 nsew
rlabel metal3 s 5825 43897 5825 43897 4 gnd
port 137 nsew
rlabel metal3 s 5825 38783 5825 38783 4 gnd
port 137 nsew
rlabel metal3 s 5825 38367 5825 38367 4 gnd
port 137 nsew
rlabel metal3 s 5825 43523 5825 43523 4 gnd
port 137 nsew
rlabel metal3 s 6250 42675 6250 42675 4 vdd
port 136 nsew
rlabel metal3 s 5825 37993 5825 37993 4 gnd
port 137 nsew
rlabel metal3 s 5825 41153 5825 41153 4 gnd
port 137 nsew
rlabel metal3 s 6250 39157 6250 39157 4 vdd
port 136 nsew
rlabel metal3 s 5825 41943 5825 41943 4 gnd
port 137 nsew
rlabel metal3 s 5825 40363 5825 40363 4 gnd
port 137 nsew
rlabel metal3 s 6250 39947 6250 39947 4 vdd
port 136 nsew
rlabel metal3 s 6250 41095 6250 41095 4 vdd
port 136 nsew
rlabel metal3 s 6250 43107 6250 43107 4 vdd
port 136 nsew
rlabel metal3 s 5825 40737 5825 40737 4 gnd
port 137 nsew
rlabel metal3 s 6250 43897 6250 43897 4 vdd
port 136 nsew
rlabel metal3 s 7336 42689 7336 42689 4 vdd
port 136 nsew
rlabel metal3 s 7336 43874 7336 43874 4 vdd
port 136 nsew
rlabel metal3 s 6682 38725 6682 38725 4 vdd
port 136 nsew
rlabel metal3 s 7064 38344 7064 38344 4 gnd
port 137 nsew
rlabel metal3 s 6682 43465 6682 43465 4 vdd
port 136 nsew
rlabel metal3 s 6682 39947 6682 39947 4 vdd
port 136 nsew
rlabel metal3 s 7064 43874 7064 43874 4 gnd
port 137 nsew
rlabel metal3 s 7336 40714 7336 40714 4 vdd
port 136 nsew
rlabel metal3 s 7064 39134 7064 39134 4 gnd
port 137 nsew
rlabel metal3 s 7064 42689 7064 42689 4 gnd
port 137 nsew
rlabel metal3 s 7336 40319 7336 40319 4 vdd
port 136 nsew
rlabel metal3 s 6682 42317 6682 42317 4 vdd
port 136 nsew
rlabel metal3 s 7336 41899 7336 41899 4 vdd
port 136 nsew
rlabel metal3 s 6682 43107 6682 43107 4 vdd
port 136 nsew
rlabel metal3 s 7336 41109 7336 41109 4 vdd
port 136 nsew
rlabel metal3 s 7064 40319 7064 40319 4 gnd
port 137 nsew
rlabel metal3 s 7064 41504 7064 41504 4 gnd
port 137 nsew
rlabel metal3 s 6682 43897 6682 43897 4 vdd
port 136 nsew
rlabel metal3 s 7336 39924 7336 39924 4 vdd
port 136 nsew
rlabel metal3 s 6682 37935 6682 37935 4 vdd
port 136 nsew
rlabel metal3 s 6682 41885 6682 41885 4 vdd
port 136 nsew
rlabel metal3 s 7064 41899 7064 41899 4 gnd
port 137 nsew
rlabel metal3 s 6682 41095 6682 41095 4 vdd
port 136 nsew
rlabel metal3 s 6682 42675 6682 42675 4 vdd
port 136 nsew
rlabel metal3 s 7336 39529 7336 39529 4 vdd
port 136 nsew
rlabel metal3 s 6682 39515 6682 39515 4 vdd
port 136 nsew
rlabel metal3 s 7336 38344 7336 38344 4 vdd
port 136 nsew
rlabel metal3 s 7064 37949 7064 37949 4 gnd
port 137 nsew
rlabel metal3 s 7336 43084 7336 43084 4 vdd
port 136 nsew
rlabel metal3 s 7336 37949 7336 37949 4 vdd
port 136 nsew
rlabel metal3 s 6682 41527 6682 41527 4 vdd
port 136 nsew
rlabel metal3 s 6682 40737 6682 40737 4 vdd
port 136 nsew
rlabel metal3 s 6682 38367 6682 38367 4 vdd
port 136 nsew
rlabel metal3 s 7064 42294 7064 42294 4 gnd
port 137 nsew
rlabel metal3 s 7336 41504 7336 41504 4 vdd
port 136 nsew
rlabel metal3 s 7064 43479 7064 43479 4 gnd
port 137 nsew
rlabel metal3 s 7336 43479 7336 43479 4 vdd
port 136 nsew
rlabel metal3 s 7064 41109 7064 41109 4 gnd
port 137 nsew
rlabel metal3 s 7064 39924 7064 39924 4 gnd
port 137 nsew
rlabel metal3 s 7336 39134 7336 39134 4 vdd
port 136 nsew
rlabel metal3 s 6682 40305 6682 40305 4 vdd
port 136 nsew
rlabel metal3 s 7064 39529 7064 39529 4 gnd
port 137 nsew
rlabel metal3 s 6682 39157 6682 39157 4 vdd
port 136 nsew
rlabel metal3 s 7064 38739 7064 38739 4 gnd
port 137 nsew
rlabel metal3 s 7064 40714 7064 40714 4 gnd
port 137 nsew
rlabel metal3 s 7336 42294 7336 42294 4 vdd
port 136 nsew
rlabel metal3 s 7336 38739 7336 38739 4 vdd
port 136 nsew
rlabel metal3 s 7064 43084 7064 43084 4 gnd
port 137 nsew
rlabel metal3 s 6682 37145 6682 37145 4 vdd
port 136 nsew
rlabel metal3 s 6682 36355 6682 36355 4 vdd
port 136 nsew
rlabel metal3 s 6682 37577 6682 37577 4 vdd
port 136 nsew
rlabel metal3 s 7336 32814 7336 32814 4 vdd
port 136 nsew
rlabel metal3 s 7336 31629 7336 31629 4 vdd
port 136 nsew
rlabel metal3 s 7336 36764 7336 36764 4 vdd
port 136 nsew
rlabel metal3 s 7336 32024 7336 32024 4 vdd
port 136 nsew
rlabel metal3 s 6682 34417 6682 34417 4 vdd
port 136 nsew
rlabel metal3 s 6682 35207 6682 35207 4 vdd
port 136 nsew
rlabel metal3 s 7336 32419 7336 32419 4 vdd
port 136 nsew
rlabel metal3 s 7336 33604 7336 33604 4 vdd
port 136 nsew
rlabel metal3 s 6682 35565 6682 35565 4 vdd
port 136 nsew
rlabel metal3 s 6682 32837 6682 32837 4 vdd
port 136 nsew
rlabel metal3 s 7064 31629 7064 31629 4 gnd
port 137 nsew
rlabel metal3 s 7336 35184 7336 35184 4 vdd
port 136 nsew
rlabel metal3 s 7064 37554 7064 37554 4 gnd
port 137 nsew
rlabel metal3 s 6682 32047 6682 32047 4 vdd
port 136 nsew
rlabel metal3 s 7336 33209 7336 33209 4 vdd
port 136 nsew
rlabel metal3 s 7336 34789 7336 34789 4 vdd
port 136 nsew
rlabel metal3 s 6682 31615 6682 31615 4 vdd
port 136 nsew
rlabel metal3 s 6682 34775 6682 34775 4 vdd
port 136 nsew
rlabel metal3 s 7336 35579 7336 35579 4 vdd
port 136 nsew
rlabel metal3 s 7336 36369 7336 36369 4 vdd
port 136 nsew
rlabel metal3 s 7064 35974 7064 35974 4 gnd
port 137 nsew
rlabel metal3 s 7064 36369 7064 36369 4 gnd
port 137 nsew
rlabel metal3 s 7336 34394 7336 34394 4 vdd
port 136 nsew
rlabel metal3 s 7064 36764 7064 36764 4 gnd
port 137 nsew
rlabel metal3 s 7336 37159 7336 37159 4 vdd
port 136 nsew
rlabel metal3 s 6682 32405 6682 32405 4 vdd
port 136 nsew
rlabel metal3 s 6682 33195 6682 33195 4 vdd
port 136 nsew
rlabel metal3 s 6682 33627 6682 33627 4 vdd
port 136 nsew
rlabel metal3 s 7064 37159 7064 37159 4 gnd
port 137 nsew
rlabel metal3 s 7064 34394 7064 34394 4 gnd
port 137 nsew
rlabel metal3 s 7064 35579 7064 35579 4 gnd
port 137 nsew
rlabel metal3 s 7064 35184 7064 35184 4 gnd
port 137 nsew
rlabel metal3 s 7064 33999 7064 33999 4 gnd
port 137 nsew
rlabel metal3 s 7064 32024 7064 32024 4 gnd
port 137 nsew
rlabel metal3 s 7064 32814 7064 32814 4 gnd
port 137 nsew
rlabel metal3 s 6682 33985 6682 33985 4 vdd
port 136 nsew
rlabel metal3 s 7336 37554 7336 37554 4 vdd
port 136 nsew
rlabel metal3 s 7336 33999 7336 33999 4 vdd
port 136 nsew
rlabel metal3 s 6682 35997 6682 35997 4 vdd
port 136 nsew
rlabel metal3 s 7064 32419 7064 32419 4 gnd
port 137 nsew
rlabel metal3 s 7064 33209 7064 33209 4 gnd
port 137 nsew
rlabel metal3 s 6682 36787 6682 36787 4 vdd
port 136 nsew
rlabel metal3 s 7064 34789 7064 34789 4 gnd
port 137 nsew
rlabel metal3 s 7064 33604 7064 33604 4 gnd
port 137 nsew
rlabel metal3 s 7336 35974 7336 35974 4 vdd
port 136 nsew
rlabel metal3 s 5825 37577 5825 37577 4 gnd
port 137 nsew
rlabel metal3 s 5825 33627 5825 33627 4 gnd
port 137 nsew
rlabel metal3 s 5825 35623 5825 35623 4 gnd
port 137 nsew
rlabel metal3 s 6250 36787 6250 36787 4 vdd
port 136 nsew
rlabel metal3 s 5825 34417 5825 34417 4 gnd
port 137 nsew
rlabel metal3 s 6250 32047 6250 32047 4 vdd
port 136 nsew
rlabel metal3 s 6250 33627 6250 33627 4 vdd
port 136 nsew
rlabel metal3 s 5825 37203 5825 37203 4 gnd
port 137 nsew
rlabel metal3 s 5825 34833 5825 34833 4 gnd
port 137 nsew
rlabel metal3 s 6250 31615 6250 31615 4 vdd
port 136 nsew
rlabel metal3 s 5825 31673 5825 31673 4 gnd
port 137 nsew
rlabel metal3 s 6250 33985 6250 33985 4 vdd
port 136 nsew
rlabel metal3 s 6250 33195 6250 33195 4 vdd
port 136 nsew
rlabel metal3 s 5825 32463 5825 32463 4 gnd
port 137 nsew
rlabel metal3 s 6250 32405 6250 32405 4 vdd
port 136 nsew
rlabel metal3 s 5825 33253 5825 33253 4 gnd
port 137 nsew
rlabel metal3 s 6250 32837 6250 32837 4 vdd
port 136 nsew
rlabel metal3 s 5825 36787 5825 36787 4 gnd
port 137 nsew
rlabel metal3 s 5825 32837 5825 32837 4 gnd
port 137 nsew
rlabel metal3 s 5825 36413 5825 36413 4 gnd
port 137 nsew
rlabel metal3 s 6250 35565 6250 35565 4 vdd
port 136 nsew
rlabel metal3 s 6250 37577 6250 37577 4 vdd
port 136 nsew
rlabel metal3 s 5825 32047 5825 32047 4 gnd
port 137 nsew
rlabel metal3 s 5825 35997 5825 35997 4 gnd
port 137 nsew
rlabel metal3 s 6250 34417 6250 34417 4 vdd
port 136 nsew
rlabel metal3 s 6250 37145 6250 37145 4 vdd
port 136 nsew
rlabel metal3 s 5825 35207 5825 35207 4 gnd
port 137 nsew
rlabel metal3 s 6250 36355 6250 36355 4 vdd
port 136 nsew
rlabel metal3 s 5825 34043 5825 34043 4 gnd
port 137 nsew
rlabel metal3 s 6250 34775 6250 34775 4 vdd
port 136 nsew
rlabel metal3 s 6250 35997 6250 35997 4 vdd
port 136 nsew
rlabel metal3 s 6250 35207 6250 35207 4 vdd
port 136 nsew
rlabel metal3 s 6250 26085 6250 26085 4 vdd
port 136 nsew
rlabel metal3 s 5825 31257 5825 31257 4 gnd
port 137 nsew
rlabel metal3 s 5825 26517 5825 26517 4 gnd
port 137 nsew
rlabel metal3 s 6250 30035 6250 30035 4 vdd
port 136 nsew
rlabel metal3 s 6250 30825 6250 30825 4 vdd
port 136 nsew
rlabel metal3 s 5825 26143 5825 26143 4 gnd
port 137 nsew
rlabel metal3 s 5825 30467 5825 30467 4 gnd
port 137 nsew
rlabel metal3 s 6250 28455 6250 28455 4 vdd
port 136 nsew
rlabel metal3 s 5825 27723 5825 27723 4 gnd
port 137 nsew
rlabel metal3 s 5825 27307 5825 27307 4 gnd
port 137 nsew
rlabel metal3 s 6250 28887 6250 28887 4 vdd
port 136 nsew
rlabel metal3 s 5825 29677 5825 29677 4 gnd
port 137 nsew
rlabel metal3 s 5825 25727 5825 25727 4 gnd
port 137 nsew
rlabel metal3 s 6250 27307 6250 27307 4 vdd
port 136 nsew
rlabel metal3 s 5825 25353 5825 25353 4 gnd
port 137 nsew
rlabel metal3 s 5825 28887 5825 28887 4 gnd
port 137 nsew
rlabel metal3 s 6250 25727 6250 25727 4 vdd
port 136 nsew
rlabel metal3 s 6250 29245 6250 29245 4 vdd
port 136 nsew
rlabel metal3 s 6250 26517 6250 26517 4 vdd
port 136 nsew
rlabel metal3 s 5825 28513 5825 28513 4 gnd
port 137 nsew
rlabel metal3 s 6250 31257 6250 31257 4 vdd
port 136 nsew
rlabel metal3 s 5825 30093 5825 30093 4 gnd
port 137 nsew
rlabel metal3 s 6250 27665 6250 27665 4 vdd
port 136 nsew
rlabel metal3 s 5825 29303 5825 29303 4 gnd
port 137 nsew
rlabel metal3 s 6250 26875 6250 26875 4 vdd
port 136 nsew
rlabel metal3 s 6250 30467 6250 30467 4 vdd
port 136 nsew
rlabel metal3 s 5825 26933 5825 26933 4 gnd
port 137 nsew
rlabel metal3 s 6250 29677 6250 29677 4 vdd
port 136 nsew
rlabel metal3 s 5825 28097 5825 28097 4 gnd
port 137 nsew
rlabel metal3 s 6250 28097 6250 28097 4 vdd
port 136 nsew
rlabel metal3 s 5825 30883 5825 30883 4 gnd
port 137 nsew
rlabel metal3 s 7336 27284 7336 27284 4 vdd
port 136 nsew
rlabel metal3 s 7336 26099 7336 26099 4 vdd
port 136 nsew
rlabel metal3 s 7064 26494 7064 26494 4 gnd
port 137 nsew
rlabel metal3 s 6682 27307 6682 27307 4 vdd
port 136 nsew
rlabel metal3 s 6682 28455 6682 28455 4 vdd
port 136 nsew
rlabel metal3 s 7336 30839 7336 30839 4 vdd
port 136 nsew
rlabel metal3 s 7336 26494 7336 26494 4 vdd
port 136 nsew
rlabel metal3 s 7064 28864 7064 28864 4 gnd
port 137 nsew
rlabel metal3 s 7336 26889 7336 26889 4 vdd
port 136 nsew
rlabel metal3 s 7336 29654 7336 29654 4 vdd
port 136 nsew
rlabel metal3 s 6682 26875 6682 26875 4 vdd
port 136 nsew
rlabel metal3 s 6682 28097 6682 28097 4 vdd
port 136 nsew
rlabel metal3 s 7064 30839 7064 30839 4 gnd
port 137 nsew
rlabel metal3 s 7336 28469 7336 28469 4 vdd
port 136 nsew
rlabel metal3 s 7336 27679 7336 27679 4 vdd
port 136 nsew
rlabel metal3 s 6682 30035 6682 30035 4 vdd
port 136 nsew
rlabel metal3 s 6682 26517 6682 26517 4 vdd
port 136 nsew
rlabel metal3 s 6682 28887 6682 28887 4 vdd
port 136 nsew
rlabel metal3 s 7064 30444 7064 30444 4 gnd
port 137 nsew
rlabel metal3 s 7336 25704 7336 25704 4 vdd
port 136 nsew
rlabel metal3 s 7064 30049 7064 30049 4 gnd
port 137 nsew
rlabel metal3 s 6682 31257 6682 31257 4 vdd
port 136 nsew
rlabel metal3 s 6682 30467 6682 30467 4 vdd
port 136 nsew
rlabel metal3 s 7336 31234 7336 31234 4 vdd
port 136 nsew
rlabel metal3 s 6682 27665 6682 27665 4 vdd
port 136 nsew
rlabel metal3 s 7064 28469 7064 28469 4 gnd
port 137 nsew
rlabel metal3 s 7064 25704 7064 25704 4 gnd
port 137 nsew
rlabel metal3 s 7064 26889 7064 26889 4 gnd
port 137 nsew
rlabel metal3 s 7064 27284 7064 27284 4 gnd
port 137 nsew
rlabel metal3 s 6682 29245 6682 29245 4 vdd
port 136 nsew
rlabel metal3 s 7064 29259 7064 29259 4 gnd
port 137 nsew
rlabel metal3 s 7336 28074 7336 28074 4 vdd
port 136 nsew
rlabel metal3 s 7336 28864 7336 28864 4 vdd
port 136 nsew
rlabel metal3 s 7064 28074 7064 28074 4 gnd
port 137 nsew
rlabel metal3 s 7064 29654 7064 29654 4 gnd
port 137 nsew
rlabel metal3 s 6682 25727 6682 25727 4 vdd
port 136 nsew
rlabel metal3 s 7336 29259 7336 29259 4 vdd
port 136 nsew
rlabel metal3 s 6682 26085 6682 26085 4 vdd
port 136 nsew
rlabel metal3 s 6682 29677 6682 29677 4 vdd
port 136 nsew
rlabel metal3 s 7336 30444 7336 30444 4 vdd
port 136 nsew
rlabel metal3 s 7064 31234 7064 31234 4 gnd
port 137 nsew
rlabel metal3 s 7064 27679 7064 27679 4 gnd
port 137 nsew
rlabel metal3 s 7336 30049 7336 30049 4 vdd
port 136 nsew
rlabel metal3 s 6682 30825 6682 30825 4 vdd
port 136 nsew
rlabel metal3 s 7064 26099 7064 26099 4 gnd
port 137 nsew
rlabel metal3 s 1204 5164 1204 5164 4 gnd
port 137 nsew
rlabel metal3 s 6682 21345 6682 21345 4 vdd
port 136 nsew
rlabel metal3 s 6682 20987 6682 20987 4 vdd
port 136 nsew
rlabel metal3 s 6682 24937 6682 24937 4 vdd
port 136 nsew
rlabel metal3 s 7336 20174 7336 20174 4 vdd
port 136 nsew
rlabel metal3 s 6682 19765 6682 19765 4 vdd
port 136 nsew
rlabel metal3 s 6682 24147 6682 24147 4 vdd
port 136 nsew
rlabel metal3 s 6682 22567 6682 22567 4 vdd
port 136 nsew
rlabel metal3 s 6682 23715 6682 23715 4 vdd
port 136 nsew
rlabel metal3 s 7064 25309 7064 25309 4 gnd
port 137 nsew
rlabel metal3 s 6682 24505 6682 24505 4 vdd
port 136 nsew
rlabel metal3 s 7336 22939 7336 22939 4 vdd
port 136 nsew
rlabel metal3 s 6682 21777 6682 21777 4 vdd
port 136 nsew
rlabel metal3 s 7336 20569 7336 20569 4 vdd
port 136 nsew
rlabel metal3 s 6682 20555 6682 20555 4 vdd
port 136 nsew
rlabel metal3 s 7064 21754 7064 21754 4 gnd
port 137 nsew
rlabel metal3 s 7336 21754 7336 21754 4 vdd
port 136 nsew
rlabel metal3 s 7336 20964 7336 20964 4 vdd
port 136 nsew
rlabel metal3 s 7336 22544 7336 22544 4 vdd
port 136 nsew
rlabel metal3 s 6682 22135 6682 22135 4 vdd
port 136 nsew
rlabel metal3 s 7336 24914 7336 24914 4 vdd
port 136 nsew
rlabel metal3 s 7064 22544 7064 22544 4 gnd
port 137 nsew
rlabel metal3 s 7336 24124 7336 24124 4 vdd
port 136 nsew
rlabel metal3 s 6682 19407 6682 19407 4 vdd
port 136 nsew
rlabel metal3 s 6682 23357 6682 23357 4 vdd
port 136 nsew
rlabel metal3 s 7336 19384 7336 19384 4 vdd
port 136 nsew
rlabel metal3 s 7336 23729 7336 23729 4 vdd
port 136 nsew
rlabel metal3 s 7064 19384 7064 19384 4 gnd
port 137 nsew
rlabel metal3 s 6682 25295 6682 25295 4 vdd
port 136 nsew
rlabel metal3 s 7064 20569 7064 20569 4 gnd
port 137 nsew
rlabel metal3 s 7064 23334 7064 23334 4 gnd
port 137 nsew
rlabel metal3 s 7064 24914 7064 24914 4 gnd
port 137 nsew
rlabel metal3 s 7336 22149 7336 22149 4 vdd
port 136 nsew
rlabel metal3 s 7064 23729 7064 23729 4 gnd
port 137 nsew
rlabel metal3 s 7336 21359 7336 21359 4 vdd
port 136 nsew
rlabel metal3 s 7064 24519 7064 24519 4 gnd
port 137 nsew
rlabel metal3 s 7064 20964 7064 20964 4 gnd
port 137 nsew
rlabel metal3 s 7064 21359 7064 21359 4 gnd
port 137 nsew
rlabel metal3 s 7064 22939 7064 22939 4 gnd
port 137 nsew
rlabel metal3 s 7064 20174 7064 20174 4 gnd
port 137 nsew
rlabel metal3 s 7336 24519 7336 24519 4 vdd
port 136 nsew
rlabel metal3 s 6682 20197 6682 20197 4 vdd
port 136 nsew
rlabel metal3 s 7336 19779 7336 19779 4 vdd
port 136 nsew
rlabel metal3 s 7064 19779 7064 19779 4 gnd
port 137 nsew
rlabel metal3 s 7064 24124 7064 24124 4 gnd
port 137 nsew
rlabel metal3 s 7336 25309 7336 25309 4 vdd
port 136 nsew
rlabel metal3 s 6682 22925 6682 22925 4 vdd
port 136 nsew
rlabel metal3 s 7064 22149 7064 22149 4 gnd
port 137 nsew
rlabel metal3 s 7336 23334 7336 23334 4 vdd
port 136 nsew
rlabel metal3 s 6250 22567 6250 22567 4 vdd
port 136 nsew
rlabel metal3 s 5825 24147 5825 24147 4 gnd
port 137 nsew
rlabel metal3 s 5825 19823 5825 19823 4 gnd
port 137 nsew
rlabel metal3 s 5825 24937 5825 24937 4 gnd
port 137 nsew
rlabel metal3 s 6250 24505 6250 24505 4 vdd
port 136 nsew
rlabel metal3 s 6250 20555 6250 20555 4 vdd
port 136 nsew
rlabel metal3 s 6250 21777 6250 21777 4 vdd
port 136 nsew
rlabel metal3 s 6250 22135 6250 22135 4 vdd
port 136 nsew
rlabel metal3 s 5825 24563 5825 24563 4 gnd
port 137 nsew
rlabel metal3 s 5825 22983 5825 22983 4 gnd
port 137 nsew
rlabel metal3 s 6250 19765 6250 19765 4 vdd
port 136 nsew
rlabel metal3 s 6250 19407 6250 19407 4 vdd
port 136 nsew
rlabel metal3 s 6250 24937 6250 24937 4 vdd
port 136 nsew
rlabel metal3 s 5825 21403 5825 21403 4 gnd
port 137 nsew
rlabel metal3 s 6250 21345 6250 21345 4 vdd
port 136 nsew
rlabel metal3 s 5825 23773 5825 23773 4 gnd
port 137 nsew
rlabel metal3 s 6250 20197 6250 20197 4 vdd
port 136 nsew
rlabel metal3 s 5825 22567 5825 22567 4 gnd
port 137 nsew
rlabel metal3 s 6250 25295 6250 25295 4 vdd
port 136 nsew
rlabel metal3 s 5825 23357 5825 23357 4 gnd
port 137 nsew
rlabel metal3 s 6250 22925 6250 22925 4 vdd
port 136 nsew
rlabel metal3 s 6250 23715 6250 23715 4 vdd
port 136 nsew
rlabel metal3 s 5825 22193 5825 22193 4 gnd
port 137 nsew
rlabel metal3 s 6250 23357 6250 23357 4 vdd
port 136 nsew
rlabel metal3 s 5825 20613 5825 20613 4 gnd
port 137 nsew
rlabel metal3 s 6250 20987 6250 20987 4 vdd
port 136 nsew
rlabel metal3 s 5825 20987 5825 20987 4 gnd
port 137 nsew
rlabel metal3 s 5825 20197 5825 20197 4 gnd
port 137 nsew
rlabel metal3 s 6250 24147 6250 24147 4 vdd
port 136 nsew
rlabel metal3 s 5825 19407 5825 19407 4 gnd
port 137 nsew
rlabel metal3 s 5825 21777 5825 21777 4 gnd
port 137 nsew
rlabel metal3 s 6250 18617 6250 18617 4 vdd
port 136 nsew
rlabel metal3 s 6250 15025 6250 15025 4 vdd
port 136 nsew
rlabel metal3 s 5825 15457 5825 15457 4 gnd
port 137 nsew
rlabel metal3 s 5825 14667 5825 14667 4 gnd
port 137 nsew
rlabel metal3 s 6250 16605 6250 16605 4 vdd
port 136 nsew
rlabel metal3 s 6250 13445 6250 13445 4 vdd
port 136 nsew
rlabel metal3 s 6250 13087 6250 13087 4 vdd
port 136 nsew
rlabel metal3 s 6250 17037 6250 17037 4 vdd
port 136 nsew
rlabel metal3 s 6250 15457 6250 15457 4 vdd
port 136 nsew
rlabel metal3 s 5825 18617 5825 18617 4 gnd
port 137 nsew
rlabel metal3 s 5825 14293 5825 14293 4 gnd
port 137 nsew
rlabel metal3 s 6250 17395 6250 17395 4 vdd
port 136 nsew
rlabel metal3 s 5825 16247 5825 16247 4 gnd
port 137 nsew
rlabel metal3 s 5825 17827 5825 17827 4 gnd
port 137 nsew
rlabel metal3 s 6250 14235 6250 14235 4 vdd
port 136 nsew
rlabel metal3 s 5825 13087 5825 13087 4 gnd
port 137 nsew
rlabel metal3 s 6250 15815 6250 15815 4 vdd
port 136 nsew
rlabel metal3 s 5825 18243 5825 18243 4 gnd
port 137 nsew
rlabel metal3 s 5825 16663 5825 16663 4 gnd
port 137 nsew
rlabel metal3 s 6250 14667 6250 14667 4 vdd
port 136 nsew
rlabel metal3 s 6250 13877 6250 13877 4 vdd
port 136 nsew
rlabel metal3 s 5825 13877 5825 13877 4 gnd
port 137 nsew
rlabel metal3 s 5825 19033 5825 19033 4 gnd
port 137 nsew
rlabel metal3 s 6250 18185 6250 18185 4 vdd
port 136 nsew
rlabel metal3 s 6250 18975 6250 18975 4 vdd
port 136 nsew
rlabel metal3 s 5825 17037 5825 17037 4 gnd
port 137 nsew
rlabel metal3 s 6250 17827 6250 17827 4 vdd
port 136 nsew
rlabel metal3 s 6250 16247 6250 16247 4 vdd
port 136 nsew
rlabel metal3 s 5825 15873 5825 15873 4 gnd
port 137 nsew
rlabel metal3 s 5825 13503 5825 13503 4 gnd
port 137 nsew
rlabel metal3 s 5825 15083 5825 15083 4 gnd
port 137 nsew
rlabel metal3 s 5825 17453 5825 17453 4 gnd
port 137 nsew
rlabel metal3 s 7336 18989 7336 18989 4 vdd
port 136 nsew
rlabel metal3 s 7064 16619 7064 16619 4 gnd
port 137 nsew
rlabel metal3 s 7336 17014 7336 17014 4 vdd
port 136 nsew
rlabel metal3 s 6682 16605 6682 16605 4 vdd
port 136 nsew
rlabel metal3 s 7336 13459 7336 13459 4 vdd
port 136 nsew
rlabel metal3 s 7064 14644 7064 14644 4 gnd
port 137 nsew
rlabel metal3 s 6682 17037 6682 17037 4 vdd
port 136 nsew
rlabel metal3 s 7064 15039 7064 15039 4 gnd
port 137 nsew
rlabel metal3 s 7064 15829 7064 15829 4 gnd
port 137 nsew
rlabel metal3 s 7336 17804 7336 17804 4 vdd
port 136 nsew
rlabel metal3 s 7064 17014 7064 17014 4 gnd
port 137 nsew
rlabel metal3 s 7336 13854 7336 13854 4 vdd
port 136 nsew
rlabel metal3 s 6682 13087 6682 13087 4 vdd
port 136 nsew
rlabel metal3 s 7336 18594 7336 18594 4 vdd
port 136 nsew
rlabel metal3 s 7336 15829 7336 15829 4 vdd
port 136 nsew
rlabel metal3 s 7064 14249 7064 14249 4 gnd
port 137 nsew
rlabel metal3 s 6682 13445 6682 13445 4 vdd
port 136 nsew
rlabel metal3 s 6682 14667 6682 14667 4 vdd
port 136 nsew
rlabel metal3 s 7064 16224 7064 16224 4 gnd
port 137 nsew
rlabel metal3 s 7064 13064 7064 13064 4 gnd
port 137 nsew
rlabel metal3 s 7064 18199 7064 18199 4 gnd
port 137 nsew
rlabel metal3 s 6682 18185 6682 18185 4 vdd
port 136 nsew
rlabel metal3 s 7336 13064 7336 13064 4 vdd
port 136 nsew
rlabel metal3 s 6682 17827 6682 17827 4 vdd
port 136 nsew
rlabel metal3 s 6682 13877 6682 13877 4 vdd
port 136 nsew
rlabel metal3 s 7064 18594 7064 18594 4 gnd
port 137 nsew
rlabel metal3 s 6682 15457 6682 15457 4 vdd
port 136 nsew
rlabel metal3 s 7336 15434 7336 15434 4 vdd
port 136 nsew
rlabel metal3 s 7336 15039 7336 15039 4 vdd
port 136 nsew
rlabel metal3 s 6682 17395 6682 17395 4 vdd
port 136 nsew
rlabel metal3 s 7336 16619 7336 16619 4 vdd
port 136 nsew
rlabel metal3 s 7336 16224 7336 16224 4 vdd
port 136 nsew
rlabel metal3 s 6682 16247 6682 16247 4 vdd
port 136 nsew
rlabel metal3 s 7336 14644 7336 14644 4 vdd
port 136 nsew
rlabel metal3 s 7336 18199 7336 18199 4 vdd
port 136 nsew
rlabel metal3 s 6682 15815 6682 15815 4 vdd
port 136 nsew
rlabel metal3 s 6682 18975 6682 18975 4 vdd
port 136 nsew
rlabel metal3 s 6682 18617 6682 18617 4 vdd
port 136 nsew
rlabel metal3 s 7064 13854 7064 13854 4 gnd
port 137 nsew
rlabel metal3 s 6682 14235 6682 14235 4 vdd
port 136 nsew
rlabel metal3 s 7336 14249 7336 14249 4 vdd
port 136 nsew
rlabel metal3 s 7064 17409 7064 17409 4 gnd
port 137 nsew
rlabel metal3 s 7336 17409 7336 17409 4 vdd
port 136 nsew
rlabel metal3 s 7064 13459 7064 13459 4 gnd
port 137 nsew
rlabel metal3 s 7064 17804 7064 17804 4 gnd
port 137 nsew
rlabel metal3 s 7064 18989 7064 18989 4 gnd
port 137 nsew
rlabel metal3 s 7064 15434 7064 15434 4 gnd
port 137 nsew
rlabel metal3 s 6682 15025 6682 15025 4 vdd
port 136 nsew
rlabel metal3 s 6682 11075 6682 11075 4 vdd
port 136 nsew
rlabel metal3 s 6682 9495 6682 9495 4 vdd
port 136 nsew
rlabel metal3 s 7336 7139 7336 7139 4 vdd
port 136 nsew
rlabel metal3 s 7064 7139 7064 7139 4 gnd
port 137 nsew
rlabel metal3 s 7336 9509 7336 9509 4 vdd
port 136 nsew
rlabel metal3 s 7064 11879 7064 11879 4 gnd
port 137 nsew
rlabel metal3 s 7064 8719 7064 8719 4 gnd
port 137 nsew
rlabel metal3 s 6682 11507 6682 11507 4 vdd
port 136 nsew
rlabel metal3 s 6682 10717 6682 10717 4 vdd
port 136 nsew
rlabel metal3 s 7336 9904 7336 9904 4 vdd
port 136 nsew
rlabel metal3 s 6682 8347 6682 8347 4 vdd
port 136 nsew
rlabel metal3 s 6682 7557 6682 7557 4 vdd
port 136 nsew
rlabel metal3 s 7064 7534 7064 7534 4 gnd
port 137 nsew
rlabel metal3 s 7336 6744 7336 6744 4 vdd
port 136 nsew
rlabel metal3 s 6682 8705 6682 8705 4 vdd
port 136 nsew
rlabel metal3 s 6682 10285 6682 10285 4 vdd
port 136 nsew
rlabel metal3 s 7336 10299 7336 10299 4 vdd
port 136 nsew
rlabel metal3 s 6682 11865 6682 11865 4 vdd
port 136 nsew
rlabel metal3 s 7336 10694 7336 10694 4 vdd
port 136 nsew
rlabel metal3 s 7064 9114 7064 9114 4 gnd
port 137 nsew
rlabel metal3 s 7336 7534 7336 7534 4 vdd
port 136 nsew
rlabel metal3 s 7064 12669 7064 12669 4 gnd
port 137 nsew
rlabel metal3 s 6682 9137 6682 9137 4 vdd
port 136 nsew
rlabel metal3 s 7336 11089 7336 11089 4 vdd
port 136 nsew
rlabel metal3 s 7336 8719 7336 8719 4 vdd
port 136 nsew
rlabel metal3 s 7336 8324 7336 8324 4 vdd
port 136 nsew
rlabel metal3 s 7064 9509 7064 9509 4 gnd
port 137 nsew
rlabel metal3 s 7064 7929 7064 7929 4 gnd
port 137 nsew
rlabel metal3 s 7336 12274 7336 12274 4 vdd
port 136 nsew
rlabel metal3 s 7336 7929 7336 7929 4 vdd
port 136 nsew
rlabel metal3 s 6682 9927 6682 9927 4 vdd
port 136 nsew
rlabel metal3 s 7336 12669 7336 12669 4 vdd
port 136 nsew
rlabel metal3 s 7064 8324 7064 8324 4 gnd
port 137 nsew
rlabel metal3 s 6682 12655 6682 12655 4 vdd
port 136 nsew
rlabel metal3 s 6682 12297 6682 12297 4 vdd
port 136 nsew
rlabel metal3 s 6682 7915 6682 7915 4 vdd
port 136 nsew
rlabel metal3 s 7336 9114 7336 9114 4 vdd
port 136 nsew
rlabel metal3 s 6682 7125 6682 7125 4 vdd
port 136 nsew
rlabel metal3 s 7336 11484 7336 11484 4 vdd
port 136 nsew
rlabel metal3 s 6682 6767 6682 6767 4 vdd
port 136 nsew
rlabel metal3 s 7064 11484 7064 11484 4 gnd
port 137 nsew
rlabel metal3 s 7064 12274 7064 12274 4 gnd
port 137 nsew
rlabel metal3 s 7064 9904 7064 9904 4 gnd
port 137 nsew
rlabel metal3 s 7064 10694 7064 10694 4 gnd
port 137 nsew
rlabel metal3 s 7064 11089 7064 11089 4 gnd
port 137 nsew
rlabel metal3 s 7064 6744 7064 6744 4 gnd
port 137 nsew
rlabel metal3 s 7336 11879 7336 11879 4 vdd
port 136 nsew
rlabel metal3 s 7064 10299 7064 10299 4 gnd
port 137 nsew
rlabel metal3 s 5825 8347 5825 8347 4 gnd
port 137 nsew
rlabel metal3 s 6250 10717 6250 10717 4 vdd
port 136 nsew
rlabel metal3 s 5825 6767 5825 6767 4 gnd
port 137 nsew
rlabel metal3 s 5825 10717 5825 10717 4 gnd
port 137 nsew
rlabel metal3 s 5825 12713 5825 12713 4 gnd
port 137 nsew
rlabel metal3 s 5825 9553 5825 9553 4 gnd
port 137 nsew
rlabel metal3 s 6250 9495 6250 9495 4 vdd
port 136 nsew
rlabel metal3 s 5825 10343 5825 10343 4 gnd
port 137 nsew
rlabel metal3 s 5825 8763 5825 8763 4 gnd
port 137 nsew
rlabel metal3 s 6250 9137 6250 9137 4 vdd
port 136 nsew
rlabel metal3 s 5825 7183 5825 7183 4 gnd
port 137 nsew
rlabel metal3 s 5825 11507 5825 11507 4 gnd
port 137 nsew
rlabel metal3 s 6250 11507 6250 11507 4 vdd
port 136 nsew
rlabel metal3 s 6250 11865 6250 11865 4 vdd
port 136 nsew
rlabel metal3 s 6250 12297 6250 12297 4 vdd
port 136 nsew
rlabel metal3 s 6250 11075 6250 11075 4 vdd
port 136 nsew
rlabel metal3 s 5825 11133 5825 11133 4 gnd
port 137 nsew
rlabel metal3 s 5825 7557 5825 7557 4 gnd
port 137 nsew
rlabel metal3 s 6250 7915 6250 7915 4 vdd
port 136 nsew
rlabel metal3 s 5825 12297 5825 12297 4 gnd
port 137 nsew
rlabel metal3 s 5825 11923 5825 11923 4 gnd
port 137 nsew
rlabel metal3 s 6250 7557 6250 7557 4 vdd
port 136 nsew
rlabel metal3 s 6250 8347 6250 8347 4 vdd
port 136 nsew
rlabel metal3 s 5825 9927 5825 9927 4 gnd
port 137 nsew
rlabel metal3 s 6250 10285 6250 10285 4 vdd
port 136 nsew
rlabel metal3 s 6250 7125 6250 7125 4 vdd
port 136 nsew
rlabel metal3 s 6250 6767 6250 6767 4 vdd
port 136 nsew
rlabel metal3 s 5825 9137 5825 9137 4 gnd
port 137 nsew
rlabel metal3 s 6250 8705 6250 8705 4 vdd
port 136 nsew
rlabel metal3 s 5825 7973 5825 7973 4 gnd
port 137 nsew
rlabel metal3 s 6250 12655 6250 12655 4 vdd
port 136 nsew
rlabel metal3 s 6250 9927 6250 9927 4 vdd
port 136 nsew
rlabel metal3 s 4046 7534 4046 7534 4 vdd
port 136 nsew
rlabel metal3 s 3392 7557 3392 7557 4 vdd
port 136 nsew
rlabel metal3 s 2960 7557 2960 7557 4 vdd
port 136 nsew
rlabel metal3 s 4046 6744 4046 6744 4 vdd
port 136 nsew
rlabel metal3 s 3392 6767 3392 6767 4 vdd
port 136 nsew
rlabel metal3 s 3774 6744 3774 6744 4 gnd
port 137 nsew
rlabel metal3 s 2960 6767 2960 6767 4 vdd
port 136 nsew
rlabel metal3 s 2535 6767 2535 6767 4 gnd
port 137 nsew
rlabel metal3 s 2535 7557 2535 7557 4 gnd
port 137 nsew
rlabel metal3 s 3774 7534 3774 7534 4 gnd
port 137 nsew
rlabel metal3 s 4046 2794 4046 2794 4 vdd
port 136 nsew
rlabel metal3 s 2960 5187 2960 5187 4 vdd
port 136 nsew
rlabel metal3 s 3774 424 3774 424 4 gnd
port 137 nsew
rlabel metal3 s 2970 2801 2970 2801 4 gnd
port 137 nsew
rlabel metal3 s 3774 1214 3774 1214 4 gnd
port 137 nsew
rlabel metal3 s 3774 3584 3774 3584 4 gnd
port 137 nsew
rlabel metal3 s 2072 2794 2072 2794 4 vdd
port 136 nsew
rlabel metal3 s 4046 1214 4046 1214 4 vdd
port 136 nsew
rlabel metal3 s 2960 5977 2960 5977 4 vdd
port 136 nsew
rlabel metal3 s 3392 5977 3392 5977 4 vdd
port 136 nsew
rlabel metal3 s 3395 3591 3395 3591 4 vdd
port 136 nsew
rlabel metal3 s 3395 1221 3395 1221 4 vdd
port 136 nsew
rlabel metal3 s 3774 2794 3774 2794 4 gnd
port 137 nsew
rlabel metal3 s 1476 5164 1476 5164 4 vdd
port 136 nsew
rlabel metal3 s 3395 2801 3395 2801 4 vdd
port 136 nsew
rlabel metal3 s 1800 424 1800 424 4 gnd
port 137 nsew
rlabel metal3 s 3395 431 3395 431 4 vdd
port 136 nsew
rlabel metal3 s 3774 5954 3774 5954 4 gnd
port 137 nsew
rlabel metal3 s 4046 3584 4046 3584 4 vdd
port 136 nsew
rlabel metal3 s 2535 5187 2535 5187 4 gnd
port 137 nsew
rlabel metal3 s 2970 1221 2970 1221 4 gnd
port 137 nsew
rlabel metal3 s 2970 3591 2970 3591 4 gnd
port 137 nsew
rlabel metal3 s 2970 431 2970 431 4 gnd
port 137 nsew
rlabel metal3 s 2072 424 2072 424 4 vdd
port 136 nsew
rlabel metal3 s 4046 5954 4046 5954 4 vdd
port 136 nsew
rlabel metal3 s 3392 5187 3392 5187 4 vdd
port 136 nsew
rlabel metal3 s 1800 2794 1800 2794 4 gnd
port 137 nsew
rlabel metal3 s 2535 5977 2535 5977 4 gnd
port 137 nsew
rlabel metal3 s 3774 5164 3774 5164 4 gnd
port 137 nsew
rlabel metal3 s 4046 5164 4046 5164 4 vdd
port 136 nsew
rlabel metal3 s 4046 424 4046 424 4 vdd
port 136 nsew
rlabel metal3 s 5825 2817 5825 2817 4 gnd
port 137 nsew
rlabel metal3 s 6250 5545 6250 5545 4 vdd
port 136 nsew
rlabel metal3 s 5825 5187 5825 5187 4 gnd
port 137 nsew
rlabel metal3 s 6250 1237 6250 1237 4 vdd
port 136 nsew
rlabel metal3 s 5825 3607 5825 3607 4 gnd
port 137 nsew
rlabel metal3 s 6250 5187 6250 5187 4 vdd
port 136 nsew
rlabel metal3 s 6250 805 6250 805 4 vdd
port 136 nsew
rlabel metal3 s 5825 863 5825 863 4 gnd
port 137 nsew
rlabel metal3 s 6250 4755 6250 4755 4 vdd
port 136 nsew
rlabel metal3 s 6250 2027 6250 2027 4 vdd
port 136 nsew
rlabel metal3 s 6250 2385 6250 2385 4 vdd
port 136 nsew
rlabel metal3 s 6250 447 6250 447 4 vdd
port 136 nsew
rlabel metal3 s 6250 1595 6250 1595 4 vdd
port 136 nsew
rlabel metal3 s 6250 2817 6250 2817 4 vdd
port 136 nsew
rlabel metal3 s 5825 4023 5825 4023 4 gnd
port 137 nsew
rlabel metal3 s 5825 447 5825 447 4 gnd
port 137 nsew
rlabel metal3 s 6250 3965 6250 3965 4 vdd
port 136 nsew
rlabel metal3 s 5825 5977 5825 5977 4 gnd
port 137 nsew
rlabel metal3 s 6250 6335 6250 6335 4 vdd
port 136 nsew
rlabel metal3 s 6250 3607 6250 3607 4 vdd
port 136 nsew
rlabel metal3 s 5825 5603 5825 5603 4 gnd
port 137 nsew
rlabel metal3 s 5825 4397 5825 4397 4 gnd
port 137 nsew
rlabel metal3 s 5825 2027 5825 2027 4 gnd
port 137 nsew
rlabel metal3 s 5825 4813 5825 4813 4 gnd
port 137 nsew
rlabel metal3 s 5825 1237 5825 1237 4 gnd
port 137 nsew
rlabel metal3 s 5825 1653 5825 1653 4 gnd
port 137 nsew
rlabel metal3 s 6250 4397 6250 4397 4 vdd
port 136 nsew
rlabel metal3 s 5825 3233 5825 3233 4 gnd
port 137 nsew
rlabel metal3 s 6250 5977 6250 5977 4 vdd
port 136 nsew
rlabel metal3 s 5825 2443 5825 2443 4 gnd
port 137 nsew
rlabel metal3 s 5825 6393 5825 6393 4 gnd
port 137 nsew
rlabel metal3 s 6250 3175 6250 3175 4 vdd
port 136 nsew
rlabel metal3 s 7336 424 7336 424 4 vdd
port 136 nsew
rlabel metal3 s 6682 1595 6682 1595 4 vdd
port 136 nsew
rlabel metal3 s 6682 6335 6682 6335 4 vdd
port 136 nsew
rlabel metal3 s 7336 3584 7336 3584 4 vdd
port 136 nsew
rlabel metal3 s 7064 819 7064 819 4 gnd
port 137 nsew
rlabel metal3 s 6682 805 6682 805 4 vdd
port 136 nsew
rlabel metal3 s 7064 1214 7064 1214 4 gnd
port 137 nsew
rlabel metal3 s 7064 3189 7064 3189 4 gnd
port 137 nsew
rlabel metal3 s 7336 3189 7336 3189 4 vdd
port 136 nsew
rlabel metal3 s 6682 4397 6682 4397 4 vdd
port 136 nsew
rlabel metal3 s 7064 5164 7064 5164 4 gnd
port 137 nsew
rlabel metal3 s 7336 1214 7336 1214 4 vdd
port 136 nsew
rlabel metal3 s 6682 3965 6682 3965 4 vdd
port 136 nsew
rlabel metal3 s 7064 3979 7064 3979 4 gnd
port 137 nsew
rlabel metal3 s 6682 4755 6682 4755 4 vdd
port 136 nsew
rlabel metal3 s 7336 4769 7336 4769 4 vdd
port 136 nsew
rlabel metal3 s 7064 3584 7064 3584 4 gnd
port 137 nsew
rlabel metal3 s 7336 6349 7336 6349 4 vdd
port 136 nsew
rlabel metal3 s 6682 5977 6682 5977 4 vdd
port 136 nsew
rlabel metal3 s 7336 4374 7336 4374 4 vdd
port 136 nsew
rlabel metal3 s 7064 5559 7064 5559 4 gnd
port 137 nsew
rlabel metal3 s 7336 3979 7336 3979 4 vdd
port 136 nsew
rlabel metal3 s 6682 5187 6682 5187 4 vdd
port 136 nsew
rlabel metal3 s 7336 5559 7336 5559 4 vdd
port 136 nsew
rlabel metal3 s 6682 2385 6682 2385 4 vdd
port 136 nsew
rlabel metal3 s 7064 4374 7064 4374 4 gnd
port 137 nsew
rlabel metal3 s 7336 819 7336 819 4 vdd
port 136 nsew
rlabel metal3 s 7064 6349 7064 6349 4 gnd
port 137 nsew
rlabel metal3 s 6682 2817 6682 2817 4 vdd
port 136 nsew
rlabel metal3 s 7064 4769 7064 4769 4 gnd
port 137 nsew
rlabel metal3 s 7064 5954 7064 5954 4 gnd
port 137 nsew
rlabel metal3 s 7064 2004 7064 2004 4 gnd
port 137 nsew
rlabel metal3 s 7336 2004 7336 2004 4 vdd
port 136 nsew
rlabel metal3 s 7064 424 7064 424 4 gnd
port 137 nsew
rlabel metal3 s 7336 1609 7336 1609 4 vdd
port 136 nsew
rlabel metal3 s 7064 1609 7064 1609 4 gnd
port 137 nsew
rlabel metal3 s 7336 2399 7336 2399 4 vdd
port 136 nsew
rlabel metal3 s 6682 1237 6682 1237 4 vdd
port 136 nsew
rlabel metal3 s 7064 2399 7064 2399 4 gnd
port 137 nsew
rlabel metal3 s 6682 3175 6682 3175 4 vdd
port 136 nsew
rlabel metal3 s 6682 3607 6682 3607 4 vdd
port 136 nsew
rlabel metal3 s 7336 5954 7336 5954 4 vdd
port 136 nsew
rlabel metal3 s 6682 2027 6682 2027 4 vdd
port 136 nsew
rlabel metal3 s 6682 447 6682 447 4 vdd
port 136 nsew
rlabel metal3 s 7064 2794 7064 2794 4 gnd
port 137 nsew
rlabel metal3 s 7336 2794 7336 2794 4 vdd
port 136 nsew
rlabel metal3 s 7336 5164 7336 5164 4 vdd
port 136 nsew
rlabel metal3 s 6682 5545 6682 5545 4 vdd
port 136 nsew
<< properties >>
string FIXED_BBOX 0 0 7512 50588
string GDS_END 4076878
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3706318
<< end >>
