magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 125 0 128 90
<< via1 >>
rect 3 0 125 90
<< metal2 >>
rect 0 0 3 90
rect 125 0 128 90
<< properties >>
string GDS_END 78996986
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78996086
<< end >>
