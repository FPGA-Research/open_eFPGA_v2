magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 157 0 160 90
<< via1 >>
rect 3 0 157 90
<< metal2 >>
rect 0 0 3 90
rect 157 0 160 90
<< properties >>
string GDS_END 79750166
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79749074
<< end >>
