magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 90
rect 477 0 480 90
<< via1 >>
rect 3 0 477 90
<< metal2 >>
rect 0 0 3 90
rect 477 0 480 90
<< properties >>
string GDS_END 91747316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91744304
<< end >>
