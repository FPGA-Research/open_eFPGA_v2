magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 10 76 514 458
<< nmoslvt >>
rect 204 102 234 432
rect 290 102 320 432
<< ndiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 234 420 290 432
rect 234 386 245 420
rect 279 386 290 420
rect 234 352 290 386
rect 234 318 245 352
rect 279 318 290 352
rect 234 284 290 318
rect 234 250 245 284
rect 279 250 290 284
rect 234 216 290 250
rect 234 182 245 216
rect 279 182 290 216
rect 234 148 290 182
rect 234 114 245 148
rect 279 114 290 148
rect 234 102 290 114
rect 320 420 376 432
rect 320 386 331 420
rect 365 386 376 420
rect 320 352 376 386
rect 320 318 331 352
rect 365 318 376 352
rect 320 284 376 318
rect 320 250 331 284
rect 365 250 376 284
rect 320 216 376 250
rect 320 182 331 216
rect 365 182 376 216
rect 320 148 376 182
rect 320 114 331 148
rect 365 114 376 148
rect 320 102 376 114
<< ndiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 245 386 279 420
rect 245 318 279 352
rect 245 250 279 284
rect 245 182 279 216
rect 245 114 279 148
rect 331 386 365 420
rect 331 318 365 352
rect 331 250 365 284
rect 331 182 365 216
rect 331 114 365 148
<< psubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 430 386 488 432
rect 430 352 442 386
rect 476 352 488 386
rect 430 318 488 352
rect 430 284 442 318
rect 476 284 488 318
rect 430 250 488 284
rect 430 216 442 250
rect 476 216 488 250
rect 430 182 488 216
rect 430 148 442 182
rect 476 148 488 182
rect 430 102 488 148
<< psubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 442 352 476 386
rect 442 284 476 318
rect 442 216 476 250
rect 442 148 476 182
<< poly >>
rect 161 504 363 524
rect 161 470 177 504
rect 211 470 245 504
rect 279 470 313 504
rect 347 470 363 504
rect 161 454 363 470
rect 204 432 234 454
rect 290 432 320 454
rect 204 80 234 102
rect 290 80 320 102
rect 161 64 363 80
rect 161 30 177 64
rect 211 30 245 64
rect 279 30 313 64
rect 347 30 363 64
rect 161 10 363 30
<< polycont >>
rect 177 470 211 504
rect 245 470 279 504
rect 313 470 347 504
rect 177 30 211 64
rect 245 30 279 64
rect 313 30 347 64
<< locali >>
rect 161 470 173 504
rect 211 470 245 504
rect 279 470 313 504
rect 351 470 363 504
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 245 420 279 436
rect 245 352 279 358
rect 245 284 279 286
rect 245 248 279 250
rect 245 176 279 182
rect 245 98 279 114
rect 331 420 365 436
rect 331 352 365 358
rect 331 284 365 286
rect 331 248 365 250
rect 331 176 365 182
rect 442 392 476 402
rect 442 320 476 352
rect 442 250 476 284
rect 442 182 476 214
rect 442 132 476 142
rect 331 98 365 114
rect 161 30 173 64
rect 211 30 245 64
rect 279 30 313 64
rect 351 30 363 64
<< viali >>
rect 173 470 177 504
rect 177 470 207 504
rect 245 470 279 504
rect 317 470 347 504
rect 347 470 351 504
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 245 386 279 392
rect 245 358 279 386
rect 245 318 279 320
rect 245 286 279 318
rect 245 216 279 248
rect 245 214 279 216
rect 245 148 279 176
rect 245 142 279 148
rect 331 386 365 392
rect 331 358 365 386
rect 331 318 365 320
rect 331 286 365 318
rect 331 216 365 248
rect 331 214 365 216
rect 331 148 365 176
rect 331 142 365 148
rect 442 386 476 392
rect 442 358 476 386
rect 442 318 476 320
rect 442 286 476 318
rect 442 216 476 248
rect 442 214 476 216
rect 442 148 476 176
rect 442 142 476 148
rect 173 30 177 64
rect 177 30 207 64
rect 245 30 279 64
rect 317 30 347 64
rect 347 30 351 64
<< metal1 >>
rect 161 504 363 524
rect 161 470 173 504
rect 207 470 245 504
rect 279 470 317 504
rect 351 470 363 504
rect 161 458 363 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 236 414 288 420
rect 236 358 245 362
rect 279 358 288 362
rect 236 350 288 358
rect 236 286 245 298
rect 279 286 288 298
rect 236 248 288 286
rect 236 214 245 248
rect 279 214 288 248
rect 236 176 288 214
rect 236 142 245 176
rect 279 142 288 176
rect 236 114 288 142
rect 322 392 374 420
rect 322 358 331 392
rect 365 358 374 392
rect 322 320 374 358
rect 322 286 331 320
rect 365 286 374 320
rect 322 248 374 286
rect 322 236 331 248
rect 365 236 374 248
rect 322 176 374 184
rect 322 172 331 176
rect 365 172 374 176
rect 322 114 374 120
rect 430 392 488 420
rect 430 358 442 392
rect 476 358 488 392
rect 430 320 488 358
rect 430 286 442 320
rect 476 286 488 320
rect 430 248 488 286
rect 430 214 442 248
rect 476 214 488 248
rect 430 176 488 214
rect 430 142 442 176
rect 476 142 488 176
rect 430 114 488 142
rect 161 64 363 76
rect 161 30 173 64
rect 207 30 245 64
rect 279 30 317 64
rect 351 30 363 64
rect 161 10 363 30
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 236 392 288 414
rect 236 362 245 392
rect 245 362 279 392
rect 279 362 288 392
rect 236 320 288 350
rect 236 298 245 320
rect 245 298 279 320
rect 279 298 288 320
rect 322 214 331 236
rect 331 214 365 236
rect 365 214 374 236
rect 322 184 374 214
rect 322 142 331 172
rect 331 142 365 172
rect 365 142 374 172
rect 322 120 374 142
<< metal2 >>
rect 10 414 514 420
rect 10 362 236 414
rect 288 362 514 414
rect 10 350 514 362
rect 10 298 236 350
rect 288 298 514 350
rect 10 292 514 298
rect 10 236 514 242
rect 10 184 150 236
rect 202 184 322 236
rect 374 184 514 236
rect 10 172 514 184
rect 10 120 150 172
rect 202 120 322 172
rect 374 120 514 172
rect 10 114 514 120
<< labels >>
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 161 10 363 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 161 458 363 524 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 430 114 488 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 5936052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5928388
<< end >>
