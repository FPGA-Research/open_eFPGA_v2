magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 319 666
<< mvpmos >>
rect 0 0 200 600
<< mvpdiff >>
rect -50 0 0 600
rect 200 0 250 600
<< poly >>
rect 0 600 200 652
rect 0 -52 200 0
<< locali >>
rect -45 -4 -11 538
rect 211 -4 245 538
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 636
use DFL1sd_CDNS_5246887918534  DFL1sd_CDNS_5246887918534_1
timestamp 1707688321
transform 1 0 200 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 228 267 228 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 96466800
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96465786
<< end >>
