magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 2756 8032 7517 11445
rect 2756 4961 6830 8032
<< nwell >>
rect 6359 22018 6859 22186
rect 2676 11239 7597 11525
rect 2676 7987 2962 11239
rect 7311 8238 7597 11239
rect 6624 7987 7597 8238
rect 2676 7952 7597 7987
rect 2676 7819 6910 7952
rect 2676 5167 2962 7819
rect 6624 5167 6910 7819
rect 2676 3057 6910 5167
<< pwell >>
rect 348 39758 2616 39912
rect 348 168 502 39758
rect 2462 168 2616 39758
rect 7976 39758 10846 39912
rect 5338 39554 7510 39640
rect 5823 28364 7441 28450
rect 3056 7663 6550 7749
rect 3056 7311 5410 7663
rect 3056 5651 3142 7311
rect 5324 7216 5410 7311
rect 5324 5764 6050 7216
rect 5324 5651 5410 5764
rect 3056 5327 5410 5651
rect 6464 5327 6550 7663
rect 3056 5241 6550 5327
rect 7976 168 8062 39758
rect 9726 168 9812 39758
rect 10692 168 10846 39758
rect 348 14 2616 168
rect 7969 14 10846 168
<< mvndiff >>
rect 3208 7363 3808 7581
rect 3938 7363 4538 7581
rect 4668 7363 5268 7581
rect 5484 5790 5622 7190
rect 5886 5790 6024 7190
rect 3208 5381 3808 5599
rect 3938 5381 4538 5599
rect 4668 5381 5268 5599
<< mvpdiff >>
rect 2742 3291 2960 4691
rect 3686 3291 3907 4691
rect 3967 4491 4188 4691
rect 5946 4491 6167 4691
rect 3967 4161 4188 4361
rect 5946 4161 6167 4361
<< mvpsubdiff >>
rect 374 39852 448 39886
rect 482 39852 516 39886
rect 374 39818 516 39852
rect 476 39784 516 39818
rect 2522 39786 2590 39886
rect 2522 39784 2556 39786
rect 374 232 476 344
rect 408 198 442 232
rect 374 164 476 198
rect 408 142 476 164
rect 2488 39752 2556 39784
rect 2488 39718 2590 39752
rect 408 130 442 142
rect 374 40 442 130
rect 2448 108 2488 142
rect 8002 39784 8066 39886
rect 10752 39786 10820 39886
rect 10752 39784 10786 39786
rect 8002 39750 8036 39784
rect 8002 39682 8036 39716
rect 9752 39750 9786 39784
rect 9752 39682 9786 39716
rect 8002 39614 8036 39648
rect 5364 39580 5398 39614
rect 5432 39580 5468 39614
rect 5502 39580 5538 39614
rect 5572 39580 5608 39614
rect 5642 39580 5678 39614
rect 5712 39580 5748 39614
rect 5782 39580 5818 39614
rect 5852 39580 5888 39614
rect 5922 39580 5958 39614
rect 5992 39580 6028 39614
rect 6062 39580 6098 39614
rect 6132 39580 6168 39614
rect 6202 39580 6238 39614
rect 6272 39580 6308 39614
rect 6342 39580 6378 39614
rect 6412 39580 6448 39614
rect 6482 39580 6518 39614
rect 6552 39580 6588 39614
rect 6622 39580 6657 39614
rect 6691 39580 6726 39614
rect 6760 39580 6795 39614
rect 6829 39580 6864 39614
rect 6898 39580 6933 39614
rect 6967 39580 7002 39614
rect 7036 39580 7071 39614
rect 7105 39580 7140 39614
rect 7174 39580 7209 39614
rect 7243 39580 7278 39614
rect 7312 39580 7347 39614
rect 7381 39580 7416 39614
rect 7450 39580 7484 39614
rect 9752 39614 9786 39648
rect 8002 39546 8036 39580
rect 8002 39478 8036 39512
rect 8002 39410 8036 39444
rect 8002 39342 8036 39376
rect 8002 39274 8036 39308
rect 8002 39206 8036 39240
rect 8002 39138 8036 39172
rect 8002 39070 8036 39104
rect 8002 39002 8036 39036
rect 8002 38934 8036 38968
rect 8002 38866 8036 38900
rect 8002 38798 8036 38832
rect 8002 38730 8036 38764
rect 8002 38662 8036 38696
rect 8002 38594 8036 38628
rect 8002 38526 8036 38560
rect 8002 38458 8036 38492
rect 8002 38390 8036 38424
rect 8002 38322 8036 38356
rect 8002 38254 8036 38288
rect 8002 38186 8036 38220
rect 8002 38118 8036 38152
rect 8002 38050 8036 38084
rect 8002 37982 8036 38016
rect 8002 37914 8036 37948
rect 8002 37846 8036 37880
rect 8002 37778 8036 37812
rect 8002 37710 8036 37744
rect 8002 37642 8036 37676
rect 8002 37574 8036 37608
rect 8002 37506 8036 37540
rect 8002 37438 8036 37472
rect 8002 37370 8036 37404
rect 8002 37302 8036 37336
rect 8002 37234 8036 37268
rect 8002 37166 8036 37200
rect 8002 37098 8036 37132
rect 8002 37030 8036 37064
rect 8002 36962 8036 36996
rect 8002 36894 8036 36928
rect 8002 36826 8036 36860
rect 8002 36758 8036 36792
rect 8002 36690 8036 36724
rect 8002 36622 8036 36656
rect 8002 36554 8036 36588
rect 8002 36486 8036 36520
rect 8002 36418 8036 36452
rect 8002 36350 8036 36384
rect 8002 36282 8036 36316
rect 8002 36214 8036 36248
rect 8002 36146 8036 36180
rect 8002 36078 8036 36112
rect 8002 36010 8036 36044
rect 8002 35942 8036 35976
rect 8002 35874 8036 35908
rect 8002 35806 8036 35840
rect 8002 35738 8036 35772
rect 8002 35670 8036 35704
rect 8002 35602 8036 35636
rect 8002 35534 8036 35568
rect 8002 35466 8036 35500
rect 8002 35398 8036 35432
rect 8002 35330 8036 35364
rect 8002 35262 8036 35296
rect 8002 35194 8036 35228
rect 8002 35126 8036 35160
rect 8002 35058 8036 35092
rect 8002 34990 8036 35024
rect 8002 34922 8036 34956
rect 8002 34854 8036 34888
rect 8002 34786 8036 34820
rect 8002 34718 8036 34752
rect 8002 34650 8036 34684
rect 8002 34582 8036 34616
rect 8002 34514 8036 34548
rect 8002 34446 8036 34480
rect 8002 34378 8036 34412
rect 8002 34310 8036 34344
rect 8002 34242 8036 34276
rect 8002 34174 8036 34208
rect 8002 34106 8036 34140
rect 8002 34038 8036 34072
rect 8002 33970 8036 34004
rect 8002 33902 8036 33936
rect 8002 33834 8036 33868
rect 8002 33766 8036 33800
rect 8002 33698 8036 33732
rect 8002 33630 8036 33664
rect 8002 33562 8036 33596
rect 8002 33494 8036 33528
rect 8002 33426 8036 33460
rect 8002 33358 8036 33392
rect 8002 33290 8036 33324
rect 8002 33222 8036 33256
rect 8002 33154 8036 33188
rect 8002 33086 8036 33120
rect 8002 33018 8036 33052
rect 8002 32950 8036 32984
rect 8002 32882 8036 32916
rect 8002 32814 8036 32848
rect 8002 32746 8036 32780
rect 8002 32678 8036 32712
rect 8002 32610 8036 32644
rect 8002 32542 8036 32576
rect 8002 32474 8036 32508
rect 8002 32406 8036 32440
rect 8002 32338 8036 32372
rect 8002 32270 8036 32304
rect 8002 32202 8036 32236
rect 8002 32134 8036 32168
rect 8002 32066 8036 32100
rect 8002 31998 8036 32032
rect 8002 31930 8036 31964
rect 8002 31862 8036 31896
rect 8002 31794 8036 31828
rect 8002 31726 8036 31760
rect 8002 31658 8036 31692
rect 8002 31590 8036 31624
rect 8002 31522 8036 31556
rect 8002 31454 8036 31488
rect 8002 31386 8036 31420
rect 8002 31318 8036 31352
rect 8002 31250 8036 31284
rect 8002 31182 8036 31216
rect 8002 31114 8036 31148
rect 8002 31046 8036 31080
rect 8002 30978 8036 31012
rect 8002 30910 8036 30944
rect 8002 30842 8036 30876
rect 8002 30774 8036 30808
rect 8002 30706 8036 30740
rect 8002 30638 8036 30672
rect 8002 30570 8036 30604
rect 8002 30502 8036 30536
rect 8002 30434 8036 30468
rect 8002 30366 8036 30400
rect 8002 30298 8036 30332
rect 8002 30230 8036 30264
rect 8002 30162 8036 30196
rect 8002 30094 8036 30128
rect 8002 30026 8036 30060
rect 8002 29958 8036 29992
rect 8002 29890 8036 29924
rect 8002 29822 8036 29856
rect 8002 29754 8036 29788
rect 8002 29686 8036 29720
rect 8002 29618 8036 29652
rect 8002 29550 8036 29584
rect 8002 29482 8036 29516
rect 8002 29414 8036 29448
rect 8002 29346 8036 29380
rect 8002 29278 8036 29312
rect 8002 29210 8036 29244
rect 8002 29142 8036 29176
rect 8002 29074 8036 29108
rect 8002 29006 8036 29040
rect 8002 28938 8036 28972
rect 8002 28870 8036 28904
rect 8002 28802 8036 28836
rect 8002 28734 8036 28768
rect 8002 28666 8036 28700
rect 8002 28598 8036 28632
rect 8002 28530 8036 28564
rect 8002 28462 8036 28496
rect 5849 28390 5873 28424
rect 5907 28390 5944 28424
rect 5978 28390 6015 28424
rect 6049 28390 6086 28424
rect 6120 28390 6157 28424
rect 6191 28390 6228 28424
rect 6262 28390 6299 28424
rect 6333 28390 6370 28424
rect 6404 28390 6441 28424
rect 6475 28390 6512 28424
rect 6546 28390 6583 28424
rect 6617 28390 6654 28424
rect 6688 28390 6725 28424
rect 6759 28390 6796 28424
rect 6830 28390 6867 28424
rect 6901 28390 6937 28424
rect 6971 28390 7007 28424
rect 7041 28390 7077 28424
rect 7111 28390 7147 28424
rect 7181 28390 7217 28424
rect 7251 28390 7287 28424
rect 7321 28390 7357 28424
rect 7391 28390 7415 28424
rect 8002 28394 8036 28428
rect 8002 28326 8036 28360
rect 8002 28258 8036 28292
rect 8002 28190 8036 28224
rect 8002 28122 8036 28156
rect 8002 28054 8036 28088
rect 8002 27986 8036 28020
rect 8002 27918 8036 27952
rect 8002 27850 8036 27884
rect 8002 27782 8036 27816
rect 8002 27714 8036 27748
rect 8002 27646 8036 27680
rect 8002 27578 8036 27612
rect 8002 27510 8036 27544
rect 8002 27442 8036 27476
rect 8002 27374 8036 27408
rect 8002 27306 8036 27340
rect 8002 27238 8036 27272
rect 8002 27170 8036 27204
rect 8002 27102 8036 27136
rect 8002 27034 8036 27068
rect 8002 26966 8036 27000
rect 8002 26898 8036 26932
rect 8002 26830 8036 26864
rect 8002 26762 8036 26796
rect 8002 26694 8036 26728
rect 8002 26626 8036 26660
rect 8002 26558 8036 26592
rect 8002 26490 8036 26524
rect 8002 26422 8036 26456
rect 8002 26354 8036 26388
rect 8002 26286 8036 26320
rect 8002 26218 8036 26252
rect 8002 26150 8036 26184
rect 8002 26082 8036 26116
rect 8002 26014 8036 26048
rect 8002 25946 8036 25980
rect 8002 25878 8036 25912
rect 8002 25810 8036 25844
rect 8002 25742 8036 25776
rect 8002 25674 8036 25708
rect 8002 25606 8036 25640
rect 8002 25538 8036 25572
rect 8002 25470 8036 25504
rect 8002 25402 8036 25436
rect 8002 25334 8036 25368
rect 8002 25266 8036 25300
rect 8002 25198 8036 25232
rect 8002 25130 8036 25164
rect 8002 25062 8036 25096
rect 8002 24994 8036 25028
rect 8002 24926 8036 24960
rect 8002 24858 8036 24892
rect 8002 24790 8036 24824
rect 8002 24722 8036 24756
rect 8002 24654 8036 24688
rect 8002 24586 8036 24620
rect 8002 24518 8036 24552
rect 8002 24450 8036 24484
rect 8002 24382 8036 24416
rect 8002 24314 8036 24348
rect 8002 24246 8036 24280
rect 8002 24178 8036 24212
rect 8002 24110 8036 24144
rect 8002 24042 8036 24076
rect 8002 23974 8036 24008
rect 8002 23906 8036 23940
rect 8002 23838 8036 23872
rect 8002 23770 8036 23804
rect 8002 23702 8036 23736
rect 8002 23634 8036 23668
rect 8002 23566 8036 23600
rect 8002 23498 8036 23532
rect 8002 23430 8036 23464
rect 8002 23362 8036 23396
rect 8002 23294 8036 23328
rect 8002 23226 8036 23260
rect 8002 23158 8036 23192
rect 8002 23090 8036 23124
rect 8002 23022 8036 23056
rect 8002 22954 8036 22988
rect 8002 22886 8036 22920
rect 8002 22818 8036 22852
rect 8002 22750 8036 22784
rect 8002 22682 8036 22716
rect 8002 22614 8036 22648
rect 8002 22546 8036 22580
rect 8002 22478 8036 22512
rect 8002 22410 8036 22444
rect 8002 22342 8036 22376
rect 8002 22274 8036 22308
rect 8002 22206 8036 22240
rect 8002 22138 8036 22172
rect 8002 22070 8036 22104
rect 8002 22002 8036 22036
rect 8002 21934 8036 21968
rect 8002 21866 8036 21900
rect 8002 21798 8036 21832
rect 8002 21730 8036 21764
rect 8002 21662 8036 21696
rect 8002 21594 8036 21628
rect 8002 21526 8036 21560
rect 8002 21458 8036 21492
rect 8002 21390 8036 21424
rect 8002 21322 8036 21356
rect 8002 21254 8036 21288
rect 8002 21186 8036 21220
rect 8002 21118 8036 21152
rect 8002 21050 8036 21084
rect 8002 20982 8036 21016
rect 8002 20914 8036 20948
rect 8002 20846 8036 20880
rect 8002 20778 8036 20812
rect 8002 20710 8036 20744
rect 8002 20642 8036 20676
rect 8002 20574 8036 20608
rect 8002 20506 8036 20540
rect 8002 20438 8036 20472
rect 8002 20370 8036 20404
rect 8002 20302 8036 20336
rect 8002 20234 8036 20268
rect 8002 20166 8036 20200
rect 8002 20098 8036 20132
rect 8002 20030 8036 20064
rect 8002 19962 8036 19996
rect 8002 19894 8036 19928
rect 8002 19826 8036 19860
rect 8002 19758 8036 19792
rect 8002 19690 8036 19724
rect 8002 19622 8036 19656
rect 8002 19554 8036 19588
rect 8002 19486 8036 19520
rect 8002 19418 8036 19452
rect 8002 19350 8036 19384
rect 8002 19282 8036 19316
rect 8002 19214 8036 19248
rect 8002 19146 8036 19180
rect 8002 19078 8036 19112
rect 8002 19010 8036 19044
rect 8002 18942 8036 18976
rect 8002 18874 8036 18908
rect 8002 18806 8036 18840
rect 8002 18738 8036 18772
rect 8002 18670 8036 18704
rect 8002 18602 8036 18636
rect 8002 18534 8036 18568
rect 8002 18466 8036 18500
rect 8002 18398 8036 18432
rect 8002 18330 8036 18364
rect 8002 18262 8036 18296
rect 8002 18194 8036 18228
rect 8002 18126 8036 18160
rect 8002 18058 8036 18092
rect 8002 17990 8036 18024
rect 8002 17922 8036 17956
rect 8002 17854 8036 17888
rect 8002 17786 8036 17820
rect 8002 17718 8036 17752
rect 8002 17650 8036 17684
rect 8002 17582 8036 17616
rect 8002 17514 8036 17548
rect 8002 17446 8036 17480
rect 8002 17378 8036 17412
rect 8002 17310 8036 17344
rect 8002 17242 8036 17276
rect 8002 17174 8036 17208
rect 8002 17106 8036 17140
rect 8002 17038 8036 17072
rect 8002 16970 8036 17004
rect 8002 16902 8036 16936
rect 8002 16834 8036 16868
rect 8002 16766 8036 16800
rect 8002 16698 8036 16732
rect 8002 16630 8036 16664
rect 8002 16562 8036 16596
rect 8002 16494 8036 16528
rect 8002 16426 8036 16460
rect 8002 16358 8036 16392
rect 8002 16290 8036 16324
rect 8002 16222 8036 16256
rect 8002 16154 8036 16188
rect 8002 16086 8036 16120
rect 8002 16018 8036 16052
rect 8002 15950 8036 15984
rect 8002 15882 8036 15916
rect 8002 15814 8036 15848
rect 8002 15746 8036 15780
rect 8002 15678 8036 15712
rect 8002 15610 8036 15644
rect 8002 15542 8036 15576
rect 8002 15474 8036 15508
rect 8002 15406 8036 15440
rect 8002 15338 8036 15372
rect 8002 15270 8036 15304
rect 8002 15202 8036 15236
rect 8002 15134 8036 15168
rect 8002 15066 8036 15100
rect 8002 14998 8036 15032
rect 8002 14930 8036 14964
rect 8002 14862 8036 14896
rect 8002 14794 8036 14828
rect 8002 14726 8036 14760
rect 8002 14658 8036 14692
rect 8002 14590 8036 14624
rect 8002 14522 8036 14556
rect 8002 14454 8036 14488
rect 8002 14386 8036 14420
rect 8002 14318 8036 14352
rect 8002 14250 8036 14284
rect 8002 14182 8036 14216
rect 8002 14114 8036 14148
rect 8002 14046 8036 14080
rect 8002 13978 8036 14012
rect 8002 13910 8036 13944
rect 8002 13842 8036 13876
rect 8002 13774 8036 13808
rect 8002 13706 8036 13740
rect 8002 13638 8036 13672
rect 8002 13570 8036 13604
rect 8002 13502 8036 13536
rect 8002 13434 8036 13468
rect 8002 13366 8036 13400
rect 8002 13298 8036 13332
rect 8002 13230 8036 13264
rect 8002 13162 8036 13196
rect 8002 13094 8036 13128
rect 8002 13026 8036 13060
rect 8002 12958 8036 12992
rect 8002 12890 8036 12924
rect 8002 12822 8036 12856
rect 8002 12754 8036 12788
rect 8002 12686 8036 12720
rect 8002 12618 8036 12652
rect 8002 12550 8036 12584
rect 8002 12482 8036 12516
rect 8002 12414 8036 12448
rect 8002 12346 8036 12380
rect 8002 12278 8036 12312
rect 8002 12210 8036 12244
rect 8002 12142 8036 12176
rect 8002 12074 8036 12108
rect 8002 12006 8036 12040
rect 8002 11938 8036 11972
rect 8002 11870 8036 11904
rect 8002 11802 8036 11836
rect 8002 11734 8036 11768
rect 8002 11666 8036 11700
rect 8002 11598 8036 11632
rect 8002 11530 8036 11564
rect 8002 11462 8036 11496
rect 8002 11394 8036 11428
rect 8002 11326 8036 11360
rect 8002 11258 8036 11292
rect 8002 11190 8036 11224
rect 8002 11122 8036 11156
rect 8002 11054 8036 11088
rect 8002 10986 8036 11020
rect 8002 10918 8036 10952
rect 8002 10850 8036 10884
rect 8002 10782 8036 10816
rect 8002 10714 8036 10748
rect 8002 10646 8036 10680
rect 8002 10578 8036 10612
rect 8002 10510 8036 10544
rect 8002 10442 8036 10476
rect 8002 10374 8036 10408
rect 8002 10306 8036 10340
rect 8002 10238 8036 10272
rect 8002 10170 8036 10204
rect 8002 10102 8036 10136
rect 8002 10034 8036 10068
rect 8002 9966 8036 10000
rect 8002 9898 8036 9932
rect 8002 9830 8036 9864
rect 8002 9762 8036 9796
rect 8002 9694 8036 9728
rect 8002 9626 8036 9660
rect 8002 9558 8036 9592
rect 8002 9490 8036 9524
rect 8002 9422 8036 9456
rect 8002 9354 8036 9388
rect 8002 9286 8036 9320
rect 8002 9218 8036 9252
rect 8002 9150 8036 9184
rect 8002 9082 8036 9116
rect 8002 9014 8036 9048
rect 8002 8946 8036 8980
rect 8002 8878 8036 8912
rect 8002 8810 8036 8844
rect 8002 8742 8036 8776
rect 8002 8674 8036 8708
rect 8002 8606 8036 8640
rect 8002 8538 8036 8572
rect 8002 8470 8036 8504
rect 8002 8402 8036 8436
rect 8002 8334 8036 8368
rect 8002 8266 8036 8300
rect 8002 8198 8036 8232
rect 8002 8130 8036 8164
rect 3082 7689 3158 7723
rect 3192 7689 3226 7723
rect 3260 7689 3294 7723
rect 3328 7689 3362 7723
rect 3396 7689 3430 7723
rect 3464 7689 3498 7723
rect 3532 7689 3566 7723
rect 3600 7689 3634 7723
rect 3668 7689 3702 7723
rect 3736 7689 3770 7723
rect 3804 7689 3838 7723
rect 3872 7689 3906 7723
rect 3940 7689 3974 7723
rect 4008 7689 4042 7723
rect 4076 7689 4110 7723
rect 4144 7689 4178 7723
rect 4212 7689 4246 7723
rect 4280 7689 4314 7723
rect 4348 7689 4382 7723
rect 4416 7689 4450 7723
rect 4484 7689 4518 7723
rect 4552 7689 4586 7723
rect 4620 7689 4654 7723
rect 4688 7689 4722 7723
rect 4756 7689 4790 7723
rect 4824 7689 4858 7723
rect 4892 7689 4926 7723
rect 4960 7689 4994 7723
rect 5028 7689 5062 7723
rect 5096 7689 5130 7723
rect 5164 7689 5198 7723
rect 5232 7689 5266 7723
rect 5300 7689 5334 7723
rect 5368 7689 5402 7723
rect 5436 7689 5470 7723
rect 5504 7689 5538 7723
rect 5572 7689 5606 7723
rect 5640 7689 5674 7723
rect 5708 7689 5742 7723
rect 5776 7689 5810 7723
rect 5844 7689 5878 7723
rect 5912 7689 5946 7723
rect 5980 7689 6014 7723
rect 6048 7689 6082 7723
rect 6116 7689 6150 7723
rect 6184 7689 6218 7723
rect 6252 7689 6286 7723
rect 6320 7689 6354 7723
rect 6388 7689 6422 7723
rect 6456 7689 6524 7723
rect 3082 7655 3116 7689
rect 3082 7587 3116 7621
rect 5350 7655 5384 7689
rect 5350 7586 5384 7621
rect 3082 7519 3116 7553
rect 3082 7451 3116 7485
rect 3082 7383 3116 7417
rect 5350 7517 5384 7552
rect 5350 7448 5384 7483
rect 5350 7379 5384 7414
rect 3082 7315 3116 7349
rect 5350 7310 5384 7345
rect 3082 7247 3116 7281
rect 3082 7179 3116 7213
rect 3082 7111 3116 7145
rect 3082 7043 3116 7077
rect 3082 6975 3116 7009
rect 3082 6907 3116 6941
rect 3082 6839 3116 6873
rect 3082 6771 3116 6805
rect 3082 6703 3116 6737
rect 3082 6635 3116 6669
rect 3082 6567 3116 6601
rect 3082 6499 3116 6533
rect 3082 6431 3116 6465
rect 3082 6363 3116 6397
rect 3082 6295 3116 6329
rect 3082 6227 3116 6261
rect 3082 6159 3116 6193
rect 3082 6091 3116 6125
rect 3082 6023 3116 6057
rect 3082 5955 3116 5989
rect 3082 5887 3116 5921
rect 3082 5819 3116 5853
rect 3082 5751 3116 5785
rect 3082 5683 3116 5717
rect 5350 7241 5384 7276
rect 5350 7172 5384 7207
rect 6490 7613 6524 7689
rect 6490 7545 6524 7579
rect 6490 7477 6524 7511
rect 6490 7409 6524 7443
rect 6490 7341 6524 7375
rect 6490 7273 6524 7307
rect 6490 7205 6524 7239
rect 5350 7103 5384 7138
rect 5350 7034 5384 7069
rect 5350 6965 5384 7000
rect 5350 6896 5384 6931
rect 5350 6827 5384 6862
rect 5350 6758 5384 6793
rect 5350 6689 5384 6724
rect 5350 6620 5384 6655
rect 5350 6551 5384 6586
rect 5350 6482 5384 6517
rect 5350 6413 5384 6448
rect 5350 6344 5384 6379
rect 5350 6275 5384 6310
rect 5350 6206 5384 6241
rect 5350 6137 5384 6172
rect 5350 6068 5384 6103
rect 5350 5999 5384 6034
rect 5350 5929 5384 5965
rect 5350 5859 5384 5895
rect 5350 5789 5384 5825
rect 6490 7137 6524 7171
rect 6490 7069 6524 7103
rect 6490 7001 6524 7035
rect 6490 6933 6524 6967
rect 6490 6865 6524 6899
rect 6490 6797 6524 6831
rect 6490 6729 6524 6763
rect 6490 6661 6524 6695
rect 6490 6593 6524 6627
rect 5350 5719 5384 5755
rect 6490 6525 6524 6559
rect 6490 6457 6524 6491
rect 6490 6389 6524 6423
rect 6490 6321 6524 6355
rect 6490 6253 6524 6287
rect 6490 6185 6524 6219
rect 6490 6117 6524 6151
rect 6490 6049 6524 6083
rect 6490 5981 6524 6015
rect 6490 5913 6524 5947
rect 6490 5845 6524 5879
rect 6490 5777 6524 5811
rect 6490 5709 6524 5743
rect 3082 5615 3116 5649
rect 5350 5649 5384 5685
rect 3082 5547 3116 5581
rect 3082 5479 3116 5513
rect 3082 5411 3116 5445
rect 5350 5579 5384 5615
rect 5350 5509 5384 5545
rect 5350 5439 5384 5475
rect 3082 5301 3116 5377
rect 5350 5369 5384 5405
rect 5350 5301 5384 5335
rect 6490 5641 6524 5675
rect 6490 5573 6524 5607
rect 6490 5505 6524 5539
rect 6490 5437 6524 5471
rect 6490 5369 6524 5403
rect 6490 5301 6524 5335
rect 3082 5267 3150 5301
rect 3184 5267 3218 5301
rect 3252 5267 3286 5301
rect 3320 5267 3354 5301
rect 3388 5267 3422 5301
rect 3456 5267 3490 5301
rect 3524 5267 3558 5301
rect 3592 5267 3626 5301
rect 3660 5267 3694 5301
rect 3728 5267 3762 5301
rect 3796 5267 3830 5301
rect 3864 5267 3898 5301
rect 3932 5267 3966 5301
rect 4000 5267 4034 5301
rect 4068 5267 4102 5301
rect 4136 5267 4170 5301
rect 4204 5267 4238 5301
rect 4272 5267 4306 5301
rect 4340 5267 4374 5301
rect 4408 5267 4442 5301
rect 4476 5267 4510 5301
rect 4544 5267 4578 5301
rect 4612 5267 4646 5301
rect 4680 5267 4714 5301
rect 4748 5267 4782 5301
rect 4816 5267 4850 5301
rect 4884 5267 4918 5301
rect 4952 5267 4986 5301
rect 5020 5267 5054 5301
rect 5088 5267 5122 5301
rect 5156 5267 5190 5301
rect 5224 5267 5258 5301
rect 5292 5267 5326 5301
rect 5360 5267 5394 5301
rect 5428 5267 5462 5301
rect 5496 5267 5530 5301
rect 5564 5267 5598 5301
rect 5632 5267 5666 5301
rect 5700 5267 5734 5301
rect 5768 5267 5802 5301
rect 5836 5267 5870 5301
rect 5904 5267 5938 5301
rect 5972 5267 6006 5301
rect 6040 5267 6074 5301
rect 6108 5267 6142 5301
rect 6176 5267 6210 5301
rect 6244 5267 6278 5301
rect 6312 5267 6346 5301
rect 6380 5267 6414 5301
rect 6448 5267 6524 5301
rect 8002 8062 8036 8096
rect 8002 7994 8036 8028
rect 8002 7926 8036 7960
rect 8002 7858 8036 7892
rect 8002 7790 8036 7824
rect 8002 7722 8036 7756
rect 8002 7654 8036 7688
rect 8002 7586 8036 7620
rect 8002 7518 8036 7552
rect 8002 7450 8036 7484
rect 8002 7382 8036 7416
rect 8002 7314 8036 7348
rect 8002 7246 8036 7280
rect 8002 7178 8036 7212
rect 8002 7110 8036 7144
rect 8002 7042 8036 7076
rect 8002 6974 8036 7008
rect 8002 6906 8036 6940
rect 8002 6838 8036 6872
rect 8002 6770 8036 6804
rect 8002 6702 8036 6736
rect 8002 6634 8036 6668
rect 8002 6566 8036 6600
rect 8002 6498 8036 6532
rect 8002 6430 8036 6464
rect 8002 6362 8036 6396
rect 8002 6294 8036 6328
rect 8002 6226 8036 6260
rect 8002 6158 8036 6192
rect 8002 6090 8036 6124
rect 8002 6022 8036 6056
rect 8002 5954 8036 5988
rect 8002 5886 8036 5920
rect 8002 5818 8036 5852
rect 8002 5750 8036 5784
rect 8002 5682 8036 5716
rect 8002 5614 8036 5648
rect 8002 5546 8036 5580
rect 8002 5478 8036 5512
rect 8002 5410 8036 5444
rect 8002 5342 8036 5376
rect 8002 5274 8036 5308
rect 8002 5206 8036 5240
rect 8002 5138 8036 5172
rect 8002 5070 8036 5104
rect 8002 5002 8036 5036
rect 8002 4934 8036 4968
rect 8002 4866 8036 4900
rect 8002 4798 8036 4832
rect 8002 4730 8036 4764
rect 8002 4662 8036 4696
rect 8002 4593 8036 4628
rect 8002 4524 8036 4559
rect 8002 4455 8036 4490
rect 8002 4386 8036 4421
rect 8002 4317 8036 4352
rect 8002 4248 8036 4283
rect 8002 4179 8036 4214
rect 8002 4110 8036 4145
rect 8002 4041 8036 4076
rect 8002 3972 8036 4007
rect 8002 3903 8036 3938
rect 8002 3834 8036 3869
rect 8002 3765 8036 3800
rect 8002 3696 8036 3731
rect 8002 3627 8036 3662
rect 8002 3558 8036 3593
rect 8002 3489 8036 3524
rect 8002 3420 8036 3455
rect 8002 3351 8036 3386
rect 8002 3282 8036 3317
rect 8002 3213 8036 3248
rect 8002 3144 8036 3179
rect 8002 3075 8036 3110
rect 8002 3006 8036 3041
rect 8002 2937 8036 2972
rect 8002 2868 8036 2903
rect 8002 2799 8036 2834
rect 8002 2730 8036 2765
rect 8002 2661 8036 2696
rect 8002 2592 8036 2627
rect 8002 2523 8036 2558
rect 8002 2454 8036 2489
rect 8002 2385 8036 2420
rect 8002 2316 8036 2351
rect 8002 2247 8036 2282
rect 8002 2178 8036 2213
rect 8002 2109 8036 2144
rect 8002 2040 8036 2075
rect 8002 1971 8036 2006
rect 8002 1902 8036 1937
rect 8002 1833 8036 1868
rect 8002 1764 8036 1799
rect 8002 1695 8036 1730
rect 8002 1626 8036 1661
rect 8002 1557 8036 1592
rect 8002 1488 8036 1523
rect 8002 1419 8036 1454
rect 8002 1350 8036 1385
rect 8002 1281 8036 1316
rect 8002 1212 8036 1247
rect 8002 1143 8036 1178
rect 8002 1074 8036 1109
rect 8002 1005 8036 1040
rect 8002 936 8036 971
rect 8002 867 8036 902
rect 8002 798 8036 833
rect 8002 729 8036 764
rect 8002 660 8036 695
rect 8002 591 8036 626
rect 8002 522 8036 557
rect 8002 453 8036 488
rect 8002 384 8036 419
rect 8002 315 8036 350
rect 8002 246 8036 281
rect 8002 177 8036 212
rect 8002 142 8036 143
rect 9752 39546 9786 39580
rect 9752 39478 9786 39512
rect 9752 39410 9786 39444
rect 9752 39342 9786 39376
rect 9752 39274 9786 39308
rect 9752 39206 9786 39240
rect 9752 39138 9786 39172
rect 9752 39070 9786 39104
rect 9752 39002 9786 39036
rect 9752 38934 9786 38968
rect 9752 38866 9786 38900
rect 9752 38798 9786 38832
rect 9752 38730 9786 38764
rect 9752 38662 9786 38696
rect 9752 38594 9786 38628
rect 9752 38526 9786 38560
rect 9752 38458 9786 38492
rect 9752 38390 9786 38424
rect 9752 38322 9786 38356
rect 9752 38254 9786 38288
rect 9752 38186 9786 38220
rect 9752 38118 9786 38152
rect 9752 38050 9786 38084
rect 9752 37982 9786 38016
rect 9752 37914 9786 37948
rect 9752 37846 9786 37880
rect 9752 37778 9786 37812
rect 9752 37710 9786 37744
rect 9752 37642 9786 37676
rect 9752 37574 9786 37608
rect 9752 37506 9786 37540
rect 9752 37438 9786 37472
rect 9752 37370 9786 37404
rect 9752 37302 9786 37336
rect 9752 37234 9786 37268
rect 9752 37166 9786 37200
rect 9752 37098 9786 37132
rect 9752 37030 9786 37064
rect 9752 36962 9786 36996
rect 9752 36894 9786 36928
rect 9752 36826 9786 36860
rect 9752 36758 9786 36792
rect 9752 36690 9786 36724
rect 9752 36622 9786 36656
rect 9752 36554 9786 36588
rect 9752 36486 9786 36520
rect 9752 36418 9786 36452
rect 9752 36350 9786 36384
rect 9752 36282 9786 36316
rect 9752 36214 9786 36248
rect 9752 36146 9786 36180
rect 9752 36078 9786 36112
rect 9752 36010 9786 36044
rect 9752 35942 9786 35976
rect 9752 35874 9786 35908
rect 9752 35806 9786 35840
rect 9752 35738 9786 35772
rect 9752 35670 9786 35704
rect 9752 35602 9786 35636
rect 9752 35534 9786 35568
rect 9752 35466 9786 35500
rect 9752 35398 9786 35432
rect 9752 35330 9786 35364
rect 9752 35262 9786 35296
rect 9752 35194 9786 35228
rect 9752 35126 9786 35160
rect 9752 35058 9786 35092
rect 9752 34990 9786 35024
rect 9752 34922 9786 34956
rect 9752 34854 9786 34888
rect 9752 34786 9786 34820
rect 9752 34718 9786 34752
rect 9752 34650 9786 34684
rect 9752 34582 9786 34616
rect 9752 34514 9786 34548
rect 9752 34446 9786 34480
rect 9752 34378 9786 34412
rect 9752 34310 9786 34344
rect 9752 34242 9786 34276
rect 9752 34174 9786 34208
rect 9752 34106 9786 34140
rect 9752 34038 9786 34072
rect 9752 33970 9786 34004
rect 9752 33902 9786 33936
rect 9752 33834 9786 33868
rect 9752 33766 9786 33800
rect 9752 33698 9786 33732
rect 9752 33630 9786 33664
rect 9752 33562 9786 33596
rect 9752 33494 9786 33528
rect 9752 33426 9786 33460
rect 9752 33358 9786 33392
rect 9752 33290 9786 33324
rect 9752 33222 9786 33256
rect 9752 33154 9786 33188
rect 9752 33086 9786 33120
rect 9752 33018 9786 33052
rect 9752 32950 9786 32984
rect 9752 32882 9786 32916
rect 9752 32814 9786 32848
rect 9752 32746 9786 32780
rect 9752 32678 9786 32712
rect 9752 32610 9786 32644
rect 9752 32542 9786 32576
rect 9752 32474 9786 32508
rect 9752 32406 9786 32440
rect 9752 32338 9786 32372
rect 9752 32270 9786 32304
rect 9752 32202 9786 32236
rect 9752 32134 9786 32168
rect 9752 32066 9786 32100
rect 9752 31998 9786 32032
rect 9752 31930 9786 31964
rect 9752 31862 9786 31896
rect 9752 31794 9786 31828
rect 9752 31726 9786 31760
rect 9752 31658 9786 31692
rect 9752 31590 9786 31624
rect 9752 31522 9786 31556
rect 9752 31454 9786 31488
rect 9752 31386 9786 31420
rect 9752 31318 9786 31352
rect 9752 31250 9786 31284
rect 9752 31182 9786 31216
rect 9752 31114 9786 31148
rect 9752 31046 9786 31080
rect 9752 30978 9786 31012
rect 9752 30910 9786 30944
rect 9752 30842 9786 30876
rect 9752 30774 9786 30808
rect 9752 30706 9786 30740
rect 9752 30638 9786 30672
rect 9752 30570 9786 30604
rect 9752 30502 9786 30536
rect 9752 30434 9786 30468
rect 9752 30366 9786 30400
rect 9752 30298 9786 30332
rect 9752 30230 9786 30264
rect 9752 30162 9786 30196
rect 9752 30094 9786 30128
rect 9752 30026 9786 30060
rect 9752 29958 9786 29992
rect 9752 29890 9786 29924
rect 9752 29822 9786 29856
rect 9752 29754 9786 29788
rect 9752 29686 9786 29720
rect 9752 29618 9786 29652
rect 9752 29550 9786 29584
rect 9752 29482 9786 29516
rect 9752 29414 9786 29448
rect 9752 29346 9786 29380
rect 9752 29278 9786 29312
rect 9752 29210 9786 29244
rect 9752 29142 9786 29176
rect 9752 29074 9786 29108
rect 9752 29006 9786 29040
rect 9752 28938 9786 28972
rect 9752 28870 9786 28904
rect 9752 28802 9786 28836
rect 9752 28734 9786 28768
rect 9752 28666 9786 28700
rect 9752 28598 9786 28632
rect 9752 28530 9786 28564
rect 9752 28462 9786 28496
rect 9752 28394 9786 28428
rect 9752 28326 9786 28360
rect 9752 28258 9786 28292
rect 9752 28190 9786 28224
rect 9752 28122 9786 28156
rect 9752 28054 9786 28088
rect 9752 27986 9786 28020
rect 9752 27918 9786 27952
rect 9752 27850 9786 27884
rect 9752 27782 9786 27816
rect 9752 27714 9786 27748
rect 9752 27646 9786 27680
rect 9752 27578 9786 27612
rect 9752 27510 9786 27544
rect 9752 27442 9786 27476
rect 9752 27374 9786 27408
rect 9752 27306 9786 27340
rect 9752 27238 9786 27272
rect 9752 27170 9786 27204
rect 9752 27102 9786 27136
rect 9752 27034 9786 27068
rect 9752 26966 9786 27000
rect 9752 26898 9786 26932
rect 9752 26830 9786 26864
rect 9752 26762 9786 26796
rect 9752 26694 9786 26728
rect 9752 26626 9786 26660
rect 9752 26558 9786 26592
rect 9752 26490 9786 26524
rect 9752 26422 9786 26456
rect 9752 26354 9786 26388
rect 9752 26286 9786 26320
rect 9752 26218 9786 26252
rect 9752 26150 9786 26184
rect 9752 26082 9786 26116
rect 9752 26014 9786 26048
rect 9752 25946 9786 25980
rect 9752 25878 9786 25912
rect 9752 25810 9786 25844
rect 9752 25742 9786 25776
rect 9752 25674 9786 25708
rect 9752 25606 9786 25640
rect 9752 25538 9786 25572
rect 9752 25470 9786 25504
rect 9752 25402 9786 25436
rect 9752 25334 9786 25368
rect 9752 25266 9786 25300
rect 9752 25198 9786 25232
rect 9752 25130 9786 25164
rect 9752 25062 9786 25096
rect 9752 24994 9786 25028
rect 9752 24926 9786 24960
rect 9752 24858 9786 24892
rect 9752 24790 9786 24824
rect 9752 24722 9786 24756
rect 9752 24654 9786 24688
rect 9752 24586 9786 24620
rect 9752 24518 9786 24552
rect 9752 24450 9786 24484
rect 9752 24382 9786 24416
rect 9752 24314 9786 24348
rect 9752 24246 9786 24280
rect 9752 24178 9786 24212
rect 9752 24110 9786 24144
rect 9752 24042 9786 24076
rect 9752 23974 9786 24008
rect 9752 23906 9786 23940
rect 9752 23838 9786 23872
rect 9752 23770 9786 23804
rect 9752 23702 9786 23736
rect 9752 23634 9786 23668
rect 9752 23566 9786 23600
rect 9752 23498 9786 23532
rect 9752 23430 9786 23464
rect 9752 23362 9786 23396
rect 9752 23294 9786 23328
rect 9752 23226 9786 23260
rect 9752 23158 9786 23192
rect 9752 23090 9786 23124
rect 9752 23022 9786 23056
rect 9752 22954 9786 22988
rect 9752 22886 9786 22920
rect 9752 22818 9786 22852
rect 9752 22750 9786 22784
rect 9752 22682 9786 22716
rect 9752 22614 9786 22648
rect 9752 22546 9786 22580
rect 9752 22478 9786 22512
rect 9752 22410 9786 22444
rect 9752 22342 9786 22376
rect 9752 22274 9786 22308
rect 9752 22206 9786 22240
rect 9752 22138 9786 22172
rect 9752 22070 9786 22104
rect 9752 22002 9786 22036
rect 9752 21934 9786 21968
rect 9752 21866 9786 21900
rect 9752 21798 9786 21832
rect 9752 21730 9786 21764
rect 9752 21662 9786 21696
rect 9752 21594 9786 21628
rect 9752 21526 9786 21560
rect 9752 21458 9786 21492
rect 9752 21390 9786 21424
rect 9752 21322 9786 21356
rect 9752 21254 9786 21288
rect 9752 21186 9786 21220
rect 9752 21118 9786 21152
rect 9752 21050 9786 21084
rect 9752 20982 9786 21016
rect 9752 20914 9786 20948
rect 9752 20846 9786 20880
rect 9752 20778 9786 20812
rect 9752 20710 9786 20744
rect 9752 20642 9786 20676
rect 9752 20574 9786 20608
rect 9752 20506 9786 20540
rect 9752 20438 9786 20472
rect 9752 20370 9786 20404
rect 9752 20302 9786 20336
rect 9752 20234 9786 20268
rect 9752 20166 9786 20200
rect 9752 20098 9786 20132
rect 9752 20030 9786 20064
rect 9752 19962 9786 19996
rect 9752 19894 9786 19928
rect 9752 19826 9786 19860
rect 9752 19758 9786 19792
rect 9752 19690 9786 19724
rect 9752 19622 9786 19656
rect 9752 19554 9786 19588
rect 9752 19486 9786 19520
rect 9752 19418 9786 19452
rect 9752 19350 9786 19384
rect 9752 19282 9786 19316
rect 9752 19214 9786 19248
rect 9752 19146 9786 19180
rect 9752 19078 9786 19112
rect 9752 19010 9786 19044
rect 9752 18942 9786 18976
rect 9752 18874 9786 18908
rect 9752 18806 9786 18840
rect 9752 18738 9786 18772
rect 9752 18670 9786 18704
rect 9752 18602 9786 18636
rect 9752 18534 9786 18568
rect 9752 18466 9786 18500
rect 9752 18398 9786 18432
rect 9752 18330 9786 18364
rect 9752 18262 9786 18296
rect 9752 18194 9786 18228
rect 9752 18126 9786 18160
rect 9752 18058 9786 18092
rect 9752 17990 9786 18024
rect 9752 17922 9786 17956
rect 9752 17854 9786 17888
rect 9752 17786 9786 17820
rect 9752 17718 9786 17752
rect 9752 17650 9786 17684
rect 9752 17582 9786 17616
rect 9752 17514 9786 17548
rect 9752 17446 9786 17480
rect 9752 17378 9786 17412
rect 9752 17310 9786 17344
rect 9752 17242 9786 17276
rect 9752 17174 9786 17208
rect 9752 17106 9786 17140
rect 9752 17038 9786 17072
rect 9752 16970 9786 17004
rect 9752 16902 9786 16936
rect 9752 16834 9786 16868
rect 9752 16766 9786 16800
rect 9752 16698 9786 16732
rect 9752 16630 9786 16664
rect 9752 16562 9786 16596
rect 9752 16494 9786 16528
rect 9752 16426 9786 16460
rect 9752 16358 9786 16392
rect 9752 16290 9786 16324
rect 9752 16222 9786 16256
rect 9752 16154 9786 16188
rect 9752 16086 9786 16120
rect 9752 16018 9786 16052
rect 9752 15950 9786 15984
rect 9752 15882 9786 15916
rect 9752 15814 9786 15848
rect 9752 15746 9786 15780
rect 9752 15678 9786 15712
rect 9752 15610 9786 15644
rect 9752 15542 9786 15576
rect 9752 15474 9786 15508
rect 9752 15406 9786 15440
rect 9752 15338 9786 15372
rect 9752 15270 9786 15304
rect 9752 15202 9786 15236
rect 9752 15134 9786 15168
rect 9752 15066 9786 15100
rect 9752 14998 9786 15032
rect 9752 14930 9786 14964
rect 9752 14862 9786 14896
rect 9752 14794 9786 14828
rect 9752 14726 9786 14760
rect 9752 14658 9786 14692
rect 9752 14590 9786 14624
rect 9752 14522 9786 14556
rect 9752 14454 9786 14488
rect 9752 14386 9786 14420
rect 9752 14318 9786 14352
rect 9752 14250 9786 14284
rect 9752 14182 9786 14216
rect 9752 14114 9786 14148
rect 9752 14046 9786 14080
rect 9752 13978 9786 14012
rect 9752 13910 9786 13944
rect 9752 13842 9786 13876
rect 9752 13774 9786 13808
rect 9752 13706 9786 13740
rect 9752 13638 9786 13672
rect 9752 13570 9786 13604
rect 9752 13502 9786 13536
rect 9752 13434 9786 13468
rect 9752 13366 9786 13400
rect 9752 13298 9786 13332
rect 9752 13230 9786 13264
rect 9752 13162 9786 13196
rect 9752 13094 9786 13128
rect 9752 13026 9786 13060
rect 9752 12958 9786 12992
rect 9752 12890 9786 12924
rect 9752 12822 9786 12856
rect 9752 12754 9786 12788
rect 9752 12686 9786 12720
rect 9752 12618 9786 12652
rect 9752 12550 9786 12584
rect 9752 12482 9786 12516
rect 9752 12414 9786 12448
rect 9752 12346 9786 12380
rect 9752 12278 9786 12312
rect 9752 12210 9786 12244
rect 9752 12142 9786 12176
rect 9752 12074 9786 12108
rect 9752 12006 9786 12040
rect 9752 11938 9786 11972
rect 9752 11870 9786 11904
rect 9752 11802 9786 11836
rect 9752 11734 9786 11768
rect 9752 11666 9786 11700
rect 9752 11598 9786 11632
rect 9752 11530 9786 11564
rect 9752 11462 9786 11496
rect 9752 11394 9786 11428
rect 9752 11326 9786 11360
rect 9752 11258 9786 11292
rect 9752 11190 9786 11224
rect 9752 11122 9786 11156
rect 9752 11054 9786 11088
rect 9752 10986 9786 11020
rect 9752 10918 9786 10952
rect 9752 10850 9786 10884
rect 9752 10782 9786 10816
rect 9752 10714 9786 10748
rect 9752 10646 9786 10680
rect 9752 10578 9786 10612
rect 9752 10510 9786 10544
rect 9752 10442 9786 10476
rect 9752 10374 9786 10408
rect 9752 10306 9786 10340
rect 9752 10238 9786 10272
rect 9752 10170 9786 10204
rect 9752 10102 9786 10136
rect 9752 10034 9786 10068
rect 9752 9966 9786 10000
rect 9752 9898 9786 9932
rect 9752 9830 9786 9864
rect 9752 9762 9786 9796
rect 9752 9694 9786 9728
rect 9752 9626 9786 9660
rect 9752 9558 9786 9592
rect 9752 9490 9786 9524
rect 9752 9422 9786 9456
rect 9752 9354 9786 9388
rect 9752 9286 9786 9320
rect 9752 9218 9786 9252
rect 9752 9150 9786 9184
rect 9752 9082 9786 9116
rect 9752 9014 9786 9048
rect 9752 8946 9786 8980
rect 9752 8878 9786 8912
rect 9752 8810 9786 8844
rect 9752 8742 9786 8776
rect 9752 8674 9786 8708
rect 9752 8606 9786 8640
rect 9752 8538 9786 8572
rect 9752 8470 9786 8504
rect 9752 8402 9786 8436
rect 9752 8334 9786 8368
rect 9752 8266 9786 8300
rect 9752 8198 9786 8232
rect 9752 8130 9786 8164
rect 9752 8062 9786 8096
rect 9752 7994 9786 8028
rect 9752 7926 9786 7960
rect 9752 7858 9786 7892
rect 9752 7790 9786 7824
rect 9752 7722 9786 7756
rect 9752 7654 9786 7688
rect 9752 7586 9786 7620
rect 9752 7518 9786 7552
rect 9752 7450 9786 7484
rect 9752 7382 9786 7416
rect 9752 7314 9786 7348
rect 9752 7246 9786 7280
rect 9752 7178 9786 7212
rect 9752 7110 9786 7144
rect 9752 7042 9786 7076
rect 9752 6974 9786 7008
rect 9752 6906 9786 6940
rect 9752 6838 9786 6872
rect 9752 6770 9786 6804
rect 9752 6702 9786 6736
rect 9752 6634 9786 6668
rect 9752 6566 9786 6600
rect 9752 6498 9786 6532
rect 9752 6430 9786 6464
rect 9752 6362 9786 6396
rect 9752 6294 9786 6328
rect 9752 6226 9786 6260
rect 9752 6158 9786 6192
rect 9752 6090 9786 6124
rect 9752 6022 9786 6056
rect 9752 5954 9786 5988
rect 9752 5886 9786 5920
rect 9752 5818 9786 5852
rect 9752 5750 9786 5784
rect 9752 5682 9786 5716
rect 9752 5614 9786 5648
rect 9752 5546 9786 5580
rect 9752 5478 9786 5512
rect 9752 5410 9786 5444
rect 9752 5342 9786 5376
rect 9752 5274 9786 5308
rect 9752 5206 9786 5240
rect 9752 5138 9786 5172
rect 9752 5070 9786 5104
rect 9752 5002 9786 5036
rect 9752 4934 9786 4968
rect 9752 4866 9786 4900
rect 9752 4798 9786 4832
rect 9752 4730 9786 4764
rect 9752 4662 9786 4696
rect 9752 4594 9786 4628
rect 9752 4526 9786 4560
rect 9752 4458 9786 4492
rect 9752 4390 9786 4424
rect 9752 4322 9786 4356
rect 9752 4254 9786 4288
rect 9752 4186 9786 4220
rect 9752 4118 9786 4152
rect 9752 4050 9786 4084
rect 9752 3982 9786 4016
rect 9752 3914 9786 3948
rect 9752 3846 9786 3880
rect 9752 3778 9786 3812
rect 9752 3710 9786 3744
rect 9752 3642 9786 3676
rect 9752 3574 9786 3608
rect 9752 3506 9786 3540
rect 9752 3438 9786 3472
rect 9752 3370 9786 3404
rect 9752 3302 9786 3336
rect 9752 3234 9786 3268
rect 9752 3166 9786 3200
rect 9752 3098 9786 3132
rect 9752 3030 9786 3064
rect 9752 2962 9786 2996
rect 9752 2894 9786 2928
rect 9752 2826 9786 2860
rect 9752 2758 9786 2792
rect 9752 2690 9786 2724
rect 9752 2622 9786 2656
rect 9752 2554 9786 2588
rect 9752 2486 9786 2520
rect 9752 2418 9786 2452
rect 9752 2349 9786 2384
rect 9752 2280 9786 2315
rect 9752 2211 9786 2246
rect 9752 2142 9786 2177
rect 9752 2073 9786 2108
rect 9752 2004 9786 2039
rect 9752 1935 9786 1970
rect 9752 1866 9786 1901
rect 9752 1797 9786 1832
rect 9752 1728 9786 1763
rect 9752 1659 9786 1694
rect 9752 1590 9786 1625
rect 9752 1521 9786 1556
rect 9752 1452 9786 1487
rect 9752 1383 9786 1418
rect 9752 1314 9786 1349
rect 9752 1245 9786 1280
rect 9752 1176 9786 1211
rect 9752 1107 9786 1142
rect 9752 1038 9786 1073
rect 9752 969 9786 1004
rect 9752 900 9786 935
rect 9752 831 9786 866
rect 9752 762 9786 797
rect 9752 693 9786 728
rect 9752 624 9786 659
rect 9752 555 9786 590
rect 9752 486 9786 521
rect 9752 417 9786 452
rect 9752 348 9786 383
rect 9752 279 9786 314
rect 9752 210 9786 245
rect 9752 142 9786 176
rect 10718 39752 10786 39784
rect 10718 39718 10820 39752
rect 2448 74 2590 108
rect 2448 40 2482 74
rect 2516 40 2590 74
rect 7995 108 8096 142
rect 7995 74 8002 108
rect 8036 74 8096 108
rect 7995 40 8096 74
rect 10646 108 10718 142
rect 10646 74 10820 108
rect 10646 40 10680 74
rect 10714 40 10820 74
<< mvnsubdiff >>
rect 6426 22085 6520 22119
rect 6554 22085 6588 22119
rect 6622 22085 6656 22119
rect 6690 22085 6724 22119
rect 6758 22085 6792 22119
rect 2802 11365 2926 11399
rect 2960 11365 2994 11399
rect 3028 11365 3062 11399
rect 3096 11365 3130 11399
rect 3164 11365 3198 11399
rect 3232 11365 3266 11399
rect 3300 11365 3334 11399
rect 3368 11365 3402 11399
rect 3436 11365 3470 11399
rect 3504 11365 3538 11399
rect 3572 11365 3606 11399
rect 3640 11365 3674 11399
rect 3708 11365 3742 11399
rect 3776 11365 3810 11399
rect 3844 11365 3878 11399
rect 3912 11365 3946 11399
rect 3980 11365 4014 11399
rect 4048 11365 4082 11399
rect 4116 11365 4150 11399
rect 4184 11365 4218 11399
rect 4252 11365 4286 11399
rect 4320 11365 4354 11399
rect 4388 11365 4422 11399
rect 4456 11365 4490 11399
rect 4524 11365 4558 11399
rect 4592 11365 4626 11399
rect 4660 11365 4694 11399
rect 4728 11365 4762 11399
rect 4796 11365 4830 11399
rect 4864 11365 4898 11399
rect 4932 11365 4966 11399
rect 5000 11365 5034 11399
rect 5068 11365 5102 11399
rect 5136 11365 5170 11399
rect 5204 11365 5238 11399
rect 5272 11365 5306 11399
rect 5340 11365 5374 11399
rect 5408 11365 5442 11399
rect 5476 11365 5510 11399
rect 5544 11365 5578 11399
rect 5612 11365 5646 11399
rect 5680 11365 5714 11399
rect 5748 11365 5782 11399
rect 5816 11365 5850 11399
rect 5884 11365 5918 11399
rect 5952 11365 5986 11399
rect 6020 11365 6054 11399
rect 6088 11365 6122 11399
rect 6156 11365 6190 11399
rect 6224 11365 6258 11399
rect 6292 11365 6326 11399
rect 6360 11365 6394 11399
rect 6428 11365 6553 11399
rect 6587 11365 6621 11399
rect 6655 11365 6689 11399
rect 6723 11365 6757 11399
rect 6791 11365 6825 11399
rect 6859 11365 6893 11399
rect 6927 11365 6961 11399
rect 6995 11365 7029 11399
rect 7063 11365 7097 11399
rect 7131 11365 7165 11399
rect 7199 11365 7233 11399
rect 7267 11365 7301 11399
rect 7335 11365 7369 11399
rect 7403 11365 7471 11399
rect 2802 11331 2836 11365
rect 2802 11263 2836 11297
rect 2802 11195 2836 11229
rect 2802 11127 2836 11161
rect 2802 11059 2836 11093
rect 2802 10991 2836 11025
rect 2802 10923 2836 10957
rect 2802 10855 2836 10889
rect 2802 10787 2836 10821
rect 2802 10719 2836 10753
rect 2802 10651 2836 10685
rect 2802 10583 2836 10617
rect 2802 10515 2836 10549
rect 2802 10447 2836 10481
rect 2802 10379 2836 10413
rect 2802 10311 2836 10345
rect 2802 10243 2836 10277
rect 2802 10175 2836 10209
rect 2802 10107 2836 10141
rect 2802 10039 2836 10073
rect 2802 9971 2836 10005
rect 2802 9903 2836 9937
rect 2802 9835 2836 9869
rect 2802 9767 2836 9801
rect 2802 9699 2836 9733
rect 2802 9631 2836 9665
rect 2802 9563 2836 9597
rect 2802 9495 2836 9529
rect 2802 9427 2836 9461
rect 2802 9359 2836 9393
rect 2802 9291 2836 9325
rect 2802 9223 2836 9257
rect 2802 9155 2836 9189
rect 2802 9087 2836 9121
rect 2802 9019 2836 9053
rect 2802 8951 2836 8985
rect 2802 8883 2836 8917
rect 2802 8815 2836 8849
rect 2802 8747 2836 8781
rect 2802 8679 2836 8713
rect 2802 8611 2836 8645
rect 2802 8543 2836 8577
rect 2802 8475 2836 8509
rect 2802 8407 2836 8441
rect 2802 8339 2836 8373
rect 2802 8271 2836 8305
rect 2802 8203 2836 8237
rect 2802 8135 2836 8169
rect 7437 11318 7471 11365
rect 7437 11250 7471 11284
rect 7437 11182 7471 11216
rect 7437 11114 7471 11148
rect 7437 11046 7471 11080
rect 7437 10978 7471 11012
rect 7437 10910 7471 10944
rect 7437 10842 7471 10876
rect 7437 10774 7471 10808
rect 7437 10706 7471 10740
rect 7437 10638 7471 10672
rect 7437 10570 7471 10604
rect 7437 10502 7471 10536
rect 7437 10434 7471 10468
rect 7437 10366 7471 10400
rect 7437 10298 7471 10332
rect 7437 10230 7471 10264
rect 7437 10162 7471 10196
rect 7437 10094 7471 10128
rect 7437 10026 7471 10060
rect 7437 9958 7471 9992
rect 7437 9890 7471 9924
rect 7437 9822 7471 9856
rect 7437 9754 7471 9788
rect 7437 9686 7471 9720
rect 7437 9618 7471 9652
rect 7437 9472 7471 9584
rect 7437 9404 7471 9438
rect 7437 9336 7471 9370
rect 7437 9268 7471 9302
rect 7437 9200 7471 9234
rect 7437 9132 7471 9166
rect 7437 9064 7471 9098
rect 7437 8996 7471 9030
rect 7437 8928 7471 8962
rect 7437 8860 7471 8894
rect 7437 8792 7471 8826
rect 7437 8724 7471 8758
rect 7437 8656 7471 8690
rect 7437 8588 7471 8622
rect 7437 8520 7471 8554
rect 7437 8452 7471 8486
rect 7437 8384 7471 8418
rect 7437 8316 7471 8350
rect 7437 8248 7471 8282
rect 7437 8180 7471 8214
rect 7437 8112 7471 8146
rect 2802 8067 2836 8101
rect 2802 7999 2836 8033
rect 2802 7931 2836 7965
rect 6750 8078 6862 8112
rect 6896 8078 6930 8112
rect 6964 8078 6998 8112
rect 7032 8078 7100 8112
rect 7134 8078 7168 8112
rect 7202 8078 7236 8112
rect 7270 8078 7304 8112
rect 7338 8078 7471 8112
rect 6750 8044 6784 8078
rect 6750 7920 6784 8010
rect 2836 7897 2870 7920
rect 2802 7886 2870 7897
rect 2904 7886 2938 7920
rect 2972 7886 3006 7920
rect 3040 7886 3074 7920
rect 3108 7886 3142 7920
rect 3176 7886 3210 7920
rect 3244 7886 3278 7920
rect 3312 7886 3346 7920
rect 3380 7886 3414 7920
rect 3448 7886 3482 7920
rect 3516 7886 3550 7920
rect 3584 7886 3618 7920
rect 3652 7886 3686 7920
rect 3720 7886 3754 7920
rect 3788 7886 3822 7920
rect 3856 7886 3890 7920
rect 3924 7886 3958 7920
rect 3992 7886 4026 7920
rect 4060 7886 4094 7920
rect 4128 7886 4162 7920
rect 4196 7886 4230 7920
rect 4264 7886 4298 7920
rect 4332 7886 4366 7920
rect 4400 7886 4434 7920
rect 4468 7886 4502 7920
rect 4536 7886 4570 7920
rect 4604 7886 4638 7920
rect 4672 7886 4706 7920
rect 4740 7886 4774 7920
rect 4808 7886 4842 7920
rect 4876 7886 4910 7920
rect 4944 7886 4978 7920
rect 5012 7886 5046 7920
rect 5080 7886 5114 7920
rect 5148 7886 5182 7920
rect 5216 7886 5250 7920
rect 5284 7886 5318 7920
rect 5352 7886 5386 7920
rect 5420 7886 5454 7920
rect 5488 7886 5522 7920
rect 5556 7886 5590 7920
rect 5624 7886 5658 7920
rect 5692 7886 5726 7920
rect 5760 7886 5794 7920
rect 5828 7886 5862 7920
rect 5896 7886 5930 7920
rect 5964 7886 5998 7920
rect 6032 7886 6066 7920
rect 6100 7886 6134 7920
rect 6168 7886 6202 7920
rect 6236 7886 6270 7920
rect 6304 7886 6338 7920
rect 6372 7886 6406 7920
rect 6440 7886 6474 7920
rect 6508 7886 6542 7920
rect 6576 7886 6610 7920
rect 6644 7886 6678 7920
rect 6712 7897 6784 7920
rect 6712 7886 6750 7897
rect 2802 7863 2836 7886
rect 2802 7795 2836 7829
rect 2802 7727 2836 7761
rect 6750 7829 6784 7863
rect 6750 7761 6784 7795
rect 2802 7659 2836 7693
rect 2802 7591 2836 7625
rect 2802 7523 2836 7557
rect 2802 7455 2836 7489
rect 2802 7387 2836 7421
rect 2802 7319 2836 7353
rect 2802 7251 2836 7285
rect 2802 7183 2836 7217
rect 2802 7115 2836 7149
rect 2802 7047 2836 7081
rect 2802 6979 2836 7013
rect 2802 6911 2836 6945
rect 2802 6843 2836 6877
rect 2802 6775 2836 6809
rect 2802 6707 2836 6741
rect 2802 6639 2836 6673
rect 2802 6571 2836 6605
rect 2802 6503 2836 6537
rect 2802 6435 2836 6469
rect 2802 6367 2836 6401
rect 2802 6299 2836 6333
rect 2802 6231 2836 6265
rect 2802 6163 2836 6197
rect 2802 6095 2836 6129
rect 2802 6027 2836 6061
rect 2802 5959 2836 5993
rect 2802 5891 2836 5925
rect 2802 5823 2836 5857
rect 2802 5755 2836 5789
rect 2802 5687 2836 5721
rect 2802 5619 2836 5653
rect 2802 5551 2836 5585
rect 2802 5483 2836 5517
rect 2802 5415 2836 5449
rect 2802 5347 2836 5381
rect 2802 5279 2836 5313
rect 6750 7693 6784 7727
rect 6750 7625 6784 7659
rect 6750 7557 6784 7591
rect 6750 7489 6784 7523
rect 6750 7421 6784 7455
rect 6750 7353 6784 7387
rect 6750 7285 6784 7319
rect 6750 7217 6784 7251
rect 6750 7149 6784 7183
rect 6750 7081 6784 7115
rect 6750 7013 6784 7047
rect 6750 6945 6784 6979
rect 6750 6877 6784 6911
rect 6750 6809 6784 6843
rect 6750 6741 6784 6775
rect 6750 6673 6784 6707
rect 6750 6605 6784 6639
rect 6750 6537 6784 6571
rect 6750 6469 6784 6503
rect 6750 6401 6784 6435
rect 6750 6333 6784 6367
rect 6750 6265 6784 6299
rect 6750 6197 6784 6231
rect 6750 6129 6784 6163
rect 6750 6061 6784 6095
rect 6750 5993 6784 6027
rect 6750 5925 6784 5959
rect 6750 5857 6784 5891
rect 6750 5789 6784 5823
rect 6750 5721 6784 5755
rect 6750 5653 6784 5687
rect 6750 5585 6784 5619
rect 6750 5517 6784 5551
rect 6750 5449 6784 5483
rect 6750 5381 6784 5415
rect 6750 5313 6784 5347
rect 2802 5143 2836 5245
rect 2802 5041 2836 5109
rect 6750 5245 6784 5279
rect 6750 5177 6784 5211
rect 6750 5109 6784 5143
rect 6750 5041 6784 5075
rect 2802 5007 2870 5041
rect 2904 5007 2938 5041
rect 2972 5007 3006 5041
rect 3040 5007 3074 5041
rect 3108 5007 3142 5041
rect 3176 5007 3210 5041
rect 3244 5007 3278 5041
rect 3312 5007 3346 5041
rect 3380 5007 3414 5041
rect 3448 5007 3482 5041
rect 3516 5007 3550 5041
rect 3584 5007 3618 5041
rect 3652 5007 3686 5041
rect 3720 5007 3754 5041
rect 3788 5007 3822 5041
rect 3856 5007 3890 5041
rect 3924 5007 3958 5041
rect 3992 5007 4026 5041
rect 4060 5007 4094 5041
rect 4128 5007 4162 5041
rect 4196 5007 4230 5041
rect 4264 5007 4298 5041
rect 4332 5007 4366 5041
rect 4400 5007 4434 5041
rect 4468 5007 4502 5041
rect 4536 5007 4570 5041
rect 4604 5007 4638 5041
rect 4672 5007 4706 5041
rect 4740 5007 4774 5041
rect 4808 5007 4842 5041
rect 4876 5007 4910 5041
rect 4944 5007 4978 5041
rect 5012 5007 5046 5041
rect 5080 5007 5114 5041
rect 5148 5007 5182 5041
rect 5216 5007 5250 5041
rect 5284 5007 5318 5041
rect 5352 5007 5386 5041
rect 5420 5007 5454 5041
rect 5488 5007 5522 5041
rect 5556 5007 5590 5041
rect 5624 5007 5658 5041
rect 5692 5007 5726 5041
rect 5760 5007 5794 5041
rect 5828 5007 5862 5041
rect 5896 5007 5930 5041
rect 5964 5007 5998 5041
rect 6032 5007 6066 5041
rect 6100 5007 6134 5041
rect 6168 5007 6202 5041
rect 6236 5007 6270 5041
rect 6304 5007 6338 5041
rect 6372 5007 6406 5041
rect 6440 5007 6474 5041
rect 6508 5007 6542 5041
rect 6576 5007 6610 5041
rect 6644 5007 6678 5041
rect 6712 5007 6784 5041
rect 2802 4860 2887 4894
rect 2921 4860 2955 4894
rect 2989 4860 3023 4894
rect 3057 4860 3091 4894
rect 3125 4860 3159 4894
rect 3193 4860 3227 4894
rect 3261 4860 3295 4894
rect 3329 4860 3363 4894
rect 3397 4860 3431 4894
rect 3465 4860 3499 4894
rect 3533 4860 3567 4894
rect 3601 4860 3635 4894
rect 3669 4860 3703 4894
rect 3737 4860 3771 4894
rect 3805 4860 3839 4894
rect 3873 4860 3907 4894
rect 3941 4860 3975 4894
rect 4009 4860 4043 4894
rect 4077 4860 4111 4894
rect 4145 4860 4179 4894
rect 4213 4860 4247 4894
rect 4281 4860 4315 4894
rect 4349 4860 4383 4894
rect 4417 4860 4451 4894
rect 4485 4860 4519 4894
rect 4553 4860 4587 4894
rect 4621 4860 4655 4894
rect 4689 4860 4723 4894
rect 4757 4860 4791 4894
rect 4825 4860 4859 4894
rect 4893 4860 4927 4894
rect 4961 4860 4995 4894
rect 5029 4860 5063 4894
rect 5097 4860 5131 4894
rect 5165 4860 5199 4894
rect 5233 4860 5267 4894
rect 5301 4860 5335 4894
rect 5369 4860 5403 4894
rect 5437 4860 5471 4894
rect 5505 4860 5539 4894
rect 5573 4860 5607 4894
rect 5641 4860 5675 4894
rect 5709 4860 5743 4894
rect 5777 4860 5811 4894
rect 5845 4860 5879 4894
rect 5913 4860 5947 4894
rect 5981 4860 6015 4894
rect 6049 4860 6083 4894
rect 6117 4860 6151 4894
rect 6185 4860 6219 4894
rect 6253 4860 6287 4894
rect 6321 4860 6355 4894
rect 6389 4860 6423 4894
rect 6457 4860 6491 4894
rect 6525 4860 6559 4894
rect 6593 4860 6627 4894
rect 6661 4860 6695 4894
rect 6729 4860 6763 4894
rect 2743 3124 2778 3158
rect 2812 3124 2846 3158
rect 2880 3124 2914 3158
rect 2948 3124 2982 3158
rect 3016 3124 3050 3158
rect 3084 3124 3118 3158
rect 3152 3124 3186 3158
rect 3220 3124 3254 3158
rect 3288 3124 3322 3158
rect 3356 3124 3390 3158
rect 3424 3124 3458 3158
rect 3492 3124 3526 3158
rect 3560 3124 3594 3158
rect 3628 3124 3662 3158
rect 3696 3124 3730 3158
rect 3764 3124 3798 3158
rect 3832 3124 3866 3158
<< mvpsubdiffcont >>
rect 448 39852 482 39886
rect 374 344 476 39818
rect 516 39784 2522 39886
rect 374 198 408 232
rect 442 198 476 232
rect 374 130 408 164
rect 2556 39752 2590 39786
rect 442 40 2448 142
rect 2488 108 2590 39718
rect 8066 39784 10752 39886
rect 8002 39716 8036 39750
rect 8002 39648 8036 39682
rect 9752 39716 9786 39750
rect 5398 39580 5432 39614
rect 5468 39580 5502 39614
rect 5538 39580 5572 39614
rect 5608 39580 5642 39614
rect 5678 39580 5712 39614
rect 5748 39580 5782 39614
rect 5818 39580 5852 39614
rect 5888 39580 5922 39614
rect 5958 39580 5992 39614
rect 6028 39580 6062 39614
rect 6098 39580 6132 39614
rect 6168 39580 6202 39614
rect 6238 39580 6272 39614
rect 6308 39580 6342 39614
rect 6378 39580 6412 39614
rect 6448 39580 6482 39614
rect 6518 39580 6552 39614
rect 6588 39580 6622 39614
rect 6657 39580 6691 39614
rect 6726 39580 6760 39614
rect 6795 39580 6829 39614
rect 6864 39580 6898 39614
rect 6933 39580 6967 39614
rect 7002 39580 7036 39614
rect 7071 39580 7105 39614
rect 7140 39580 7174 39614
rect 7209 39580 7243 39614
rect 7278 39580 7312 39614
rect 7347 39580 7381 39614
rect 7416 39580 7450 39614
rect 8002 39580 8036 39614
rect 9752 39648 9786 39682
rect 8002 39512 8036 39546
rect 8002 39444 8036 39478
rect 8002 39376 8036 39410
rect 8002 39308 8036 39342
rect 8002 39240 8036 39274
rect 8002 39172 8036 39206
rect 8002 39104 8036 39138
rect 8002 39036 8036 39070
rect 8002 38968 8036 39002
rect 8002 38900 8036 38934
rect 8002 38832 8036 38866
rect 8002 38764 8036 38798
rect 8002 38696 8036 38730
rect 8002 38628 8036 38662
rect 8002 38560 8036 38594
rect 8002 38492 8036 38526
rect 8002 38424 8036 38458
rect 8002 38356 8036 38390
rect 8002 38288 8036 38322
rect 8002 38220 8036 38254
rect 8002 38152 8036 38186
rect 8002 38084 8036 38118
rect 8002 38016 8036 38050
rect 8002 37948 8036 37982
rect 8002 37880 8036 37914
rect 8002 37812 8036 37846
rect 8002 37744 8036 37778
rect 8002 37676 8036 37710
rect 8002 37608 8036 37642
rect 8002 37540 8036 37574
rect 8002 37472 8036 37506
rect 8002 37404 8036 37438
rect 8002 37336 8036 37370
rect 8002 37268 8036 37302
rect 8002 37200 8036 37234
rect 8002 37132 8036 37166
rect 8002 37064 8036 37098
rect 8002 36996 8036 37030
rect 8002 36928 8036 36962
rect 8002 36860 8036 36894
rect 8002 36792 8036 36826
rect 8002 36724 8036 36758
rect 8002 36656 8036 36690
rect 8002 36588 8036 36622
rect 8002 36520 8036 36554
rect 8002 36452 8036 36486
rect 8002 36384 8036 36418
rect 8002 36316 8036 36350
rect 8002 36248 8036 36282
rect 8002 36180 8036 36214
rect 8002 36112 8036 36146
rect 8002 36044 8036 36078
rect 8002 35976 8036 36010
rect 8002 35908 8036 35942
rect 8002 35840 8036 35874
rect 8002 35772 8036 35806
rect 8002 35704 8036 35738
rect 8002 35636 8036 35670
rect 8002 35568 8036 35602
rect 8002 35500 8036 35534
rect 8002 35432 8036 35466
rect 8002 35364 8036 35398
rect 8002 35296 8036 35330
rect 8002 35228 8036 35262
rect 8002 35160 8036 35194
rect 8002 35092 8036 35126
rect 8002 35024 8036 35058
rect 8002 34956 8036 34990
rect 8002 34888 8036 34922
rect 8002 34820 8036 34854
rect 8002 34752 8036 34786
rect 8002 34684 8036 34718
rect 8002 34616 8036 34650
rect 8002 34548 8036 34582
rect 8002 34480 8036 34514
rect 8002 34412 8036 34446
rect 8002 34344 8036 34378
rect 8002 34276 8036 34310
rect 8002 34208 8036 34242
rect 8002 34140 8036 34174
rect 8002 34072 8036 34106
rect 8002 34004 8036 34038
rect 8002 33936 8036 33970
rect 8002 33868 8036 33902
rect 8002 33800 8036 33834
rect 8002 33732 8036 33766
rect 8002 33664 8036 33698
rect 8002 33596 8036 33630
rect 8002 33528 8036 33562
rect 8002 33460 8036 33494
rect 8002 33392 8036 33426
rect 8002 33324 8036 33358
rect 8002 33256 8036 33290
rect 8002 33188 8036 33222
rect 8002 33120 8036 33154
rect 8002 33052 8036 33086
rect 8002 32984 8036 33018
rect 8002 32916 8036 32950
rect 8002 32848 8036 32882
rect 8002 32780 8036 32814
rect 8002 32712 8036 32746
rect 8002 32644 8036 32678
rect 8002 32576 8036 32610
rect 8002 32508 8036 32542
rect 8002 32440 8036 32474
rect 8002 32372 8036 32406
rect 8002 32304 8036 32338
rect 8002 32236 8036 32270
rect 8002 32168 8036 32202
rect 8002 32100 8036 32134
rect 8002 32032 8036 32066
rect 8002 31964 8036 31998
rect 8002 31896 8036 31930
rect 8002 31828 8036 31862
rect 8002 31760 8036 31794
rect 8002 31692 8036 31726
rect 8002 31624 8036 31658
rect 8002 31556 8036 31590
rect 8002 31488 8036 31522
rect 8002 31420 8036 31454
rect 8002 31352 8036 31386
rect 8002 31284 8036 31318
rect 8002 31216 8036 31250
rect 8002 31148 8036 31182
rect 8002 31080 8036 31114
rect 8002 31012 8036 31046
rect 8002 30944 8036 30978
rect 8002 30876 8036 30910
rect 8002 30808 8036 30842
rect 8002 30740 8036 30774
rect 8002 30672 8036 30706
rect 8002 30604 8036 30638
rect 8002 30536 8036 30570
rect 8002 30468 8036 30502
rect 8002 30400 8036 30434
rect 8002 30332 8036 30366
rect 8002 30264 8036 30298
rect 8002 30196 8036 30230
rect 8002 30128 8036 30162
rect 8002 30060 8036 30094
rect 8002 29992 8036 30026
rect 8002 29924 8036 29958
rect 8002 29856 8036 29890
rect 8002 29788 8036 29822
rect 8002 29720 8036 29754
rect 8002 29652 8036 29686
rect 8002 29584 8036 29618
rect 8002 29516 8036 29550
rect 8002 29448 8036 29482
rect 8002 29380 8036 29414
rect 8002 29312 8036 29346
rect 8002 29244 8036 29278
rect 8002 29176 8036 29210
rect 8002 29108 8036 29142
rect 8002 29040 8036 29074
rect 8002 28972 8036 29006
rect 8002 28904 8036 28938
rect 8002 28836 8036 28870
rect 8002 28768 8036 28802
rect 8002 28700 8036 28734
rect 8002 28632 8036 28666
rect 8002 28564 8036 28598
rect 8002 28496 8036 28530
rect 8002 28428 8036 28462
rect 5873 28390 5907 28424
rect 5944 28390 5978 28424
rect 6015 28390 6049 28424
rect 6086 28390 6120 28424
rect 6157 28390 6191 28424
rect 6228 28390 6262 28424
rect 6299 28390 6333 28424
rect 6370 28390 6404 28424
rect 6441 28390 6475 28424
rect 6512 28390 6546 28424
rect 6583 28390 6617 28424
rect 6654 28390 6688 28424
rect 6725 28390 6759 28424
rect 6796 28390 6830 28424
rect 6867 28390 6901 28424
rect 6937 28390 6971 28424
rect 7007 28390 7041 28424
rect 7077 28390 7111 28424
rect 7147 28390 7181 28424
rect 7217 28390 7251 28424
rect 7287 28390 7321 28424
rect 7357 28390 7391 28424
rect 8002 28360 8036 28394
rect 8002 28292 8036 28326
rect 8002 28224 8036 28258
rect 8002 28156 8036 28190
rect 8002 28088 8036 28122
rect 8002 28020 8036 28054
rect 8002 27952 8036 27986
rect 8002 27884 8036 27918
rect 8002 27816 8036 27850
rect 8002 27748 8036 27782
rect 8002 27680 8036 27714
rect 8002 27612 8036 27646
rect 8002 27544 8036 27578
rect 8002 27476 8036 27510
rect 8002 27408 8036 27442
rect 8002 27340 8036 27374
rect 8002 27272 8036 27306
rect 8002 27204 8036 27238
rect 8002 27136 8036 27170
rect 8002 27068 8036 27102
rect 8002 27000 8036 27034
rect 8002 26932 8036 26966
rect 8002 26864 8036 26898
rect 8002 26796 8036 26830
rect 8002 26728 8036 26762
rect 8002 26660 8036 26694
rect 8002 26592 8036 26626
rect 8002 26524 8036 26558
rect 8002 26456 8036 26490
rect 8002 26388 8036 26422
rect 8002 26320 8036 26354
rect 8002 26252 8036 26286
rect 8002 26184 8036 26218
rect 8002 26116 8036 26150
rect 8002 26048 8036 26082
rect 8002 25980 8036 26014
rect 8002 25912 8036 25946
rect 8002 25844 8036 25878
rect 8002 25776 8036 25810
rect 8002 25708 8036 25742
rect 8002 25640 8036 25674
rect 8002 25572 8036 25606
rect 8002 25504 8036 25538
rect 8002 25436 8036 25470
rect 8002 25368 8036 25402
rect 8002 25300 8036 25334
rect 8002 25232 8036 25266
rect 8002 25164 8036 25198
rect 8002 25096 8036 25130
rect 8002 25028 8036 25062
rect 8002 24960 8036 24994
rect 8002 24892 8036 24926
rect 8002 24824 8036 24858
rect 8002 24756 8036 24790
rect 8002 24688 8036 24722
rect 8002 24620 8036 24654
rect 8002 24552 8036 24586
rect 8002 24484 8036 24518
rect 8002 24416 8036 24450
rect 8002 24348 8036 24382
rect 8002 24280 8036 24314
rect 8002 24212 8036 24246
rect 8002 24144 8036 24178
rect 8002 24076 8036 24110
rect 8002 24008 8036 24042
rect 8002 23940 8036 23974
rect 8002 23872 8036 23906
rect 8002 23804 8036 23838
rect 8002 23736 8036 23770
rect 8002 23668 8036 23702
rect 8002 23600 8036 23634
rect 8002 23532 8036 23566
rect 8002 23464 8036 23498
rect 8002 23396 8036 23430
rect 8002 23328 8036 23362
rect 8002 23260 8036 23294
rect 8002 23192 8036 23226
rect 8002 23124 8036 23158
rect 8002 23056 8036 23090
rect 8002 22988 8036 23022
rect 8002 22920 8036 22954
rect 8002 22852 8036 22886
rect 8002 22784 8036 22818
rect 8002 22716 8036 22750
rect 8002 22648 8036 22682
rect 8002 22580 8036 22614
rect 8002 22512 8036 22546
rect 8002 22444 8036 22478
rect 8002 22376 8036 22410
rect 8002 22308 8036 22342
rect 8002 22240 8036 22274
rect 8002 22172 8036 22206
rect 8002 22104 8036 22138
rect 8002 22036 8036 22070
rect 8002 21968 8036 22002
rect 8002 21900 8036 21934
rect 8002 21832 8036 21866
rect 8002 21764 8036 21798
rect 8002 21696 8036 21730
rect 8002 21628 8036 21662
rect 8002 21560 8036 21594
rect 8002 21492 8036 21526
rect 8002 21424 8036 21458
rect 8002 21356 8036 21390
rect 8002 21288 8036 21322
rect 8002 21220 8036 21254
rect 8002 21152 8036 21186
rect 8002 21084 8036 21118
rect 8002 21016 8036 21050
rect 8002 20948 8036 20982
rect 8002 20880 8036 20914
rect 8002 20812 8036 20846
rect 8002 20744 8036 20778
rect 8002 20676 8036 20710
rect 8002 20608 8036 20642
rect 8002 20540 8036 20574
rect 8002 20472 8036 20506
rect 8002 20404 8036 20438
rect 8002 20336 8036 20370
rect 8002 20268 8036 20302
rect 8002 20200 8036 20234
rect 8002 20132 8036 20166
rect 8002 20064 8036 20098
rect 8002 19996 8036 20030
rect 8002 19928 8036 19962
rect 8002 19860 8036 19894
rect 8002 19792 8036 19826
rect 8002 19724 8036 19758
rect 8002 19656 8036 19690
rect 8002 19588 8036 19622
rect 8002 19520 8036 19554
rect 8002 19452 8036 19486
rect 8002 19384 8036 19418
rect 8002 19316 8036 19350
rect 8002 19248 8036 19282
rect 8002 19180 8036 19214
rect 8002 19112 8036 19146
rect 8002 19044 8036 19078
rect 8002 18976 8036 19010
rect 8002 18908 8036 18942
rect 8002 18840 8036 18874
rect 8002 18772 8036 18806
rect 8002 18704 8036 18738
rect 8002 18636 8036 18670
rect 8002 18568 8036 18602
rect 8002 18500 8036 18534
rect 8002 18432 8036 18466
rect 8002 18364 8036 18398
rect 8002 18296 8036 18330
rect 8002 18228 8036 18262
rect 8002 18160 8036 18194
rect 8002 18092 8036 18126
rect 8002 18024 8036 18058
rect 8002 17956 8036 17990
rect 8002 17888 8036 17922
rect 8002 17820 8036 17854
rect 8002 17752 8036 17786
rect 8002 17684 8036 17718
rect 8002 17616 8036 17650
rect 8002 17548 8036 17582
rect 8002 17480 8036 17514
rect 8002 17412 8036 17446
rect 8002 17344 8036 17378
rect 8002 17276 8036 17310
rect 8002 17208 8036 17242
rect 8002 17140 8036 17174
rect 8002 17072 8036 17106
rect 8002 17004 8036 17038
rect 8002 16936 8036 16970
rect 8002 16868 8036 16902
rect 8002 16800 8036 16834
rect 8002 16732 8036 16766
rect 8002 16664 8036 16698
rect 8002 16596 8036 16630
rect 8002 16528 8036 16562
rect 8002 16460 8036 16494
rect 8002 16392 8036 16426
rect 8002 16324 8036 16358
rect 8002 16256 8036 16290
rect 8002 16188 8036 16222
rect 8002 16120 8036 16154
rect 8002 16052 8036 16086
rect 8002 15984 8036 16018
rect 8002 15916 8036 15950
rect 8002 15848 8036 15882
rect 8002 15780 8036 15814
rect 8002 15712 8036 15746
rect 8002 15644 8036 15678
rect 8002 15576 8036 15610
rect 8002 15508 8036 15542
rect 8002 15440 8036 15474
rect 8002 15372 8036 15406
rect 8002 15304 8036 15338
rect 8002 15236 8036 15270
rect 8002 15168 8036 15202
rect 8002 15100 8036 15134
rect 8002 15032 8036 15066
rect 8002 14964 8036 14998
rect 8002 14896 8036 14930
rect 8002 14828 8036 14862
rect 8002 14760 8036 14794
rect 8002 14692 8036 14726
rect 8002 14624 8036 14658
rect 8002 14556 8036 14590
rect 8002 14488 8036 14522
rect 8002 14420 8036 14454
rect 8002 14352 8036 14386
rect 8002 14284 8036 14318
rect 8002 14216 8036 14250
rect 8002 14148 8036 14182
rect 8002 14080 8036 14114
rect 8002 14012 8036 14046
rect 8002 13944 8036 13978
rect 8002 13876 8036 13910
rect 8002 13808 8036 13842
rect 8002 13740 8036 13774
rect 8002 13672 8036 13706
rect 8002 13604 8036 13638
rect 8002 13536 8036 13570
rect 8002 13468 8036 13502
rect 8002 13400 8036 13434
rect 8002 13332 8036 13366
rect 8002 13264 8036 13298
rect 8002 13196 8036 13230
rect 8002 13128 8036 13162
rect 8002 13060 8036 13094
rect 8002 12992 8036 13026
rect 8002 12924 8036 12958
rect 8002 12856 8036 12890
rect 8002 12788 8036 12822
rect 8002 12720 8036 12754
rect 8002 12652 8036 12686
rect 8002 12584 8036 12618
rect 8002 12516 8036 12550
rect 8002 12448 8036 12482
rect 8002 12380 8036 12414
rect 8002 12312 8036 12346
rect 8002 12244 8036 12278
rect 8002 12176 8036 12210
rect 8002 12108 8036 12142
rect 8002 12040 8036 12074
rect 8002 11972 8036 12006
rect 8002 11904 8036 11938
rect 8002 11836 8036 11870
rect 8002 11768 8036 11802
rect 8002 11700 8036 11734
rect 8002 11632 8036 11666
rect 8002 11564 8036 11598
rect 8002 11496 8036 11530
rect 8002 11428 8036 11462
rect 8002 11360 8036 11394
rect 8002 11292 8036 11326
rect 8002 11224 8036 11258
rect 8002 11156 8036 11190
rect 8002 11088 8036 11122
rect 8002 11020 8036 11054
rect 8002 10952 8036 10986
rect 8002 10884 8036 10918
rect 8002 10816 8036 10850
rect 8002 10748 8036 10782
rect 8002 10680 8036 10714
rect 8002 10612 8036 10646
rect 8002 10544 8036 10578
rect 8002 10476 8036 10510
rect 8002 10408 8036 10442
rect 8002 10340 8036 10374
rect 8002 10272 8036 10306
rect 8002 10204 8036 10238
rect 8002 10136 8036 10170
rect 8002 10068 8036 10102
rect 8002 10000 8036 10034
rect 8002 9932 8036 9966
rect 8002 9864 8036 9898
rect 8002 9796 8036 9830
rect 8002 9728 8036 9762
rect 8002 9660 8036 9694
rect 8002 9592 8036 9626
rect 8002 9524 8036 9558
rect 8002 9456 8036 9490
rect 8002 9388 8036 9422
rect 8002 9320 8036 9354
rect 8002 9252 8036 9286
rect 8002 9184 8036 9218
rect 8002 9116 8036 9150
rect 8002 9048 8036 9082
rect 8002 8980 8036 9014
rect 8002 8912 8036 8946
rect 8002 8844 8036 8878
rect 8002 8776 8036 8810
rect 8002 8708 8036 8742
rect 8002 8640 8036 8674
rect 8002 8572 8036 8606
rect 8002 8504 8036 8538
rect 8002 8436 8036 8470
rect 8002 8368 8036 8402
rect 8002 8300 8036 8334
rect 8002 8232 8036 8266
rect 8002 8164 8036 8198
rect 8002 8096 8036 8130
rect 3158 7689 3192 7723
rect 3226 7689 3260 7723
rect 3294 7689 3328 7723
rect 3362 7689 3396 7723
rect 3430 7689 3464 7723
rect 3498 7689 3532 7723
rect 3566 7689 3600 7723
rect 3634 7689 3668 7723
rect 3702 7689 3736 7723
rect 3770 7689 3804 7723
rect 3838 7689 3872 7723
rect 3906 7689 3940 7723
rect 3974 7689 4008 7723
rect 4042 7689 4076 7723
rect 4110 7689 4144 7723
rect 4178 7689 4212 7723
rect 4246 7689 4280 7723
rect 4314 7689 4348 7723
rect 4382 7689 4416 7723
rect 4450 7689 4484 7723
rect 4518 7689 4552 7723
rect 4586 7689 4620 7723
rect 4654 7689 4688 7723
rect 4722 7689 4756 7723
rect 4790 7689 4824 7723
rect 4858 7689 4892 7723
rect 4926 7689 4960 7723
rect 4994 7689 5028 7723
rect 5062 7689 5096 7723
rect 5130 7689 5164 7723
rect 5198 7689 5232 7723
rect 5266 7689 5300 7723
rect 5334 7689 5368 7723
rect 5402 7689 5436 7723
rect 5470 7689 5504 7723
rect 5538 7689 5572 7723
rect 5606 7689 5640 7723
rect 5674 7689 5708 7723
rect 5742 7689 5776 7723
rect 5810 7689 5844 7723
rect 5878 7689 5912 7723
rect 5946 7689 5980 7723
rect 6014 7689 6048 7723
rect 6082 7689 6116 7723
rect 6150 7689 6184 7723
rect 6218 7689 6252 7723
rect 6286 7689 6320 7723
rect 6354 7689 6388 7723
rect 6422 7689 6456 7723
rect 3082 7621 3116 7655
rect 3082 7553 3116 7587
rect 5350 7621 5384 7655
rect 3082 7485 3116 7519
rect 3082 7417 3116 7451
rect 3082 7349 3116 7383
rect 5350 7552 5384 7586
rect 5350 7483 5384 7517
rect 5350 7414 5384 7448
rect 3082 7281 3116 7315
rect 5350 7345 5384 7379
rect 3082 7213 3116 7247
rect 3082 7145 3116 7179
rect 3082 7077 3116 7111
rect 3082 7009 3116 7043
rect 3082 6941 3116 6975
rect 3082 6873 3116 6907
rect 3082 6805 3116 6839
rect 3082 6737 3116 6771
rect 3082 6669 3116 6703
rect 3082 6601 3116 6635
rect 3082 6533 3116 6567
rect 3082 6465 3116 6499
rect 3082 6397 3116 6431
rect 3082 6329 3116 6363
rect 3082 6261 3116 6295
rect 3082 6193 3116 6227
rect 3082 6125 3116 6159
rect 3082 6057 3116 6091
rect 3082 5989 3116 6023
rect 3082 5921 3116 5955
rect 3082 5853 3116 5887
rect 3082 5785 3116 5819
rect 3082 5717 3116 5751
rect 3082 5649 3116 5683
rect 5350 7276 5384 7310
rect 5350 7207 5384 7241
rect 6490 7579 6524 7613
rect 6490 7511 6524 7545
rect 6490 7443 6524 7477
rect 6490 7375 6524 7409
rect 6490 7307 6524 7341
rect 6490 7239 6524 7273
rect 5350 7138 5384 7172
rect 5350 7069 5384 7103
rect 5350 7000 5384 7034
rect 5350 6931 5384 6965
rect 5350 6862 5384 6896
rect 5350 6793 5384 6827
rect 5350 6724 5384 6758
rect 5350 6655 5384 6689
rect 5350 6586 5384 6620
rect 5350 6517 5384 6551
rect 5350 6448 5384 6482
rect 5350 6379 5384 6413
rect 5350 6310 5384 6344
rect 5350 6241 5384 6275
rect 5350 6172 5384 6206
rect 5350 6103 5384 6137
rect 5350 6034 5384 6068
rect 5350 5965 5384 5999
rect 5350 5895 5384 5929
rect 5350 5825 5384 5859
rect 6490 7171 6524 7205
rect 6490 7103 6524 7137
rect 6490 7035 6524 7069
rect 6490 6967 6524 7001
rect 6490 6899 6524 6933
rect 6490 6831 6524 6865
rect 6490 6763 6524 6797
rect 6490 6695 6524 6729
rect 6490 6627 6524 6661
rect 6490 6559 6524 6593
rect 5350 5755 5384 5789
rect 5350 5685 5384 5719
rect 6490 6491 6524 6525
rect 6490 6423 6524 6457
rect 6490 6355 6524 6389
rect 6490 6287 6524 6321
rect 6490 6219 6524 6253
rect 6490 6151 6524 6185
rect 6490 6083 6524 6117
rect 6490 6015 6524 6049
rect 6490 5947 6524 5981
rect 6490 5879 6524 5913
rect 6490 5811 6524 5845
rect 6490 5743 6524 5777
rect 3082 5581 3116 5615
rect 5350 5615 5384 5649
rect 3082 5513 3116 5547
rect 3082 5445 3116 5479
rect 3082 5377 3116 5411
rect 5350 5545 5384 5579
rect 5350 5475 5384 5509
rect 5350 5405 5384 5439
rect 5350 5335 5384 5369
rect 6490 5675 6524 5709
rect 6490 5607 6524 5641
rect 6490 5539 6524 5573
rect 6490 5471 6524 5505
rect 6490 5403 6524 5437
rect 6490 5335 6524 5369
rect 3150 5267 3184 5301
rect 3218 5267 3252 5301
rect 3286 5267 3320 5301
rect 3354 5267 3388 5301
rect 3422 5267 3456 5301
rect 3490 5267 3524 5301
rect 3558 5267 3592 5301
rect 3626 5267 3660 5301
rect 3694 5267 3728 5301
rect 3762 5267 3796 5301
rect 3830 5267 3864 5301
rect 3898 5267 3932 5301
rect 3966 5267 4000 5301
rect 4034 5267 4068 5301
rect 4102 5267 4136 5301
rect 4170 5267 4204 5301
rect 4238 5267 4272 5301
rect 4306 5267 4340 5301
rect 4374 5267 4408 5301
rect 4442 5267 4476 5301
rect 4510 5267 4544 5301
rect 4578 5267 4612 5301
rect 4646 5267 4680 5301
rect 4714 5267 4748 5301
rect 4782 5267 4816 5301
rect 4850 5267 4884 5301
rect 4918 5267 4952 5301
rect 4986 5267 5020 5301
rect 5054 5267 5088 5301
rect 5122 5267 5156 5301
rect 5190 5267 5224 5301
rect 5258 5267 5292 5301
rect 5326 5267 5360 5301
rect 5394 5267 5428 5301
rect 5462 5267 5496 5301
rect 5530 5267 5564 5301
rect 5598 5267 5632 5301
rect 5666 5267 5700 5301
rect 5734 5267 5768 5301
rect 5802 5267 5836 5301
rect 5870 5267 5904 5301
rect 5938 5267 5972 5301
rect 6006 5267 6040 5301
rect 6074 5267 6108 5301
rect 6142 5267 6176 5301
rect 6210 5267 6244 5301
rect 6278 5267 6312 5301
rect 6346 5267 6380 5301
rect 6414 5267 6448 5301
rect 8002 8028 8036 8062
rect 8002 7960 8036 7994
rect 8002 7892 8036 7926
rect 8002 7824 8036 7858
rect 8002 7756 8036 7790
rect 8002 7688 8036 7722
rect 8002 7620 8036 7654
rect 8002 7552 8036 7586
rect 8002 7484 8036 7518
rect 8002 7416 8036 7450
rect 8002 7348 8036 7382
rect 8002 7280 8036 7314
rect 8002 7212 8036 7246
rect 8002 7144 8036 7178
rect 8002 7076 8036 7110
rect 8002 7008 8036 7042
rect 8002 6940 8036 6974
rect 8002 6872 8036 6906
rect 8002 6804 8036 6838
rect 8002 6736 8036 6770
rect 8002 6668 8036 6702
rect 8002 6600 8036 6634
rect 8002 6532 8036 6566
rect 8002 6464 8036 6498
rect 8002 6396 8036 6430
rect 8002 6328 8036 6362
rect 8002 6260 8036 6294
rect 8002 6192 8036 6226
rect 8002 6124 8036 6158
rect 8002 6056 8036 6090
rect 8002 5988 8036 6022
rect 8002 5920 8036 5954
rect 8002 5852 8036 5886
rect 8002 5784 8036 5818
rect 8002 5716 8036 5750
rect 8002 5648 8036 5682
rect 8002 5580 8036 5614
rect 8002 5512 8036 5546
rect 8002 5444 8036 5478
rect 8002 5376 8036 5410
rect 8002 5308 8036 5342
rect 8002 5240 8036 5274
rect 8002 5172 8036 5206
rect 8002 5104 8036 5138
rect 8002 5036 8036 5070
rect 8002 4968 8036 5002
rect 8002 4900 8036 4934
rect 8002 4832 8036 4866
rect 8002 4764 8036 4798
rect 8002 4696 8036 4730
rect 8002 4628 8036 4662
rect 8002 4559 8036 4593
rect 8002 4490 8036 4524
rect 8002 4421 8036 4455
rect 8002 4352 8036 4386
rect 8002 4283 8036 4317
rect 8002 4214 8036 4248
rect 8002 4145 8036 4179
rect 8002 4076 8036 4110
rect 8002 4007 8036 4041
rect 8002 3938 8036 3972
rect 8002 3869 8036 3903
rect 8002 3800 8036 3834
rect 8002 3731 8036 3765
rect 8002 3662 8036 3696
rect 8002 3593 8036 3627
rect 8002 3524 8036 3558
rect 8002 3455 8036 3489
rect 8002 3386 8036 3420
rect 8002 3317 8036 3351
rect 8002 3248 8036 3282
rect 8002 3179 8036 3213
rect 8002 3110 8036 3144
rect 8002 3041 8036 3075
rect 8002 2972 8036 3006
rect 8002 2903 8036 2937
rect 8002 2834 8036 2868
rect 8002 2765 8036 2799
rect 8002 2696 8036 2730
rect 8002 2627 8036 2661
rect 8002 2558 8036 2592
rect 8002 2489 8036 2523
rect 8002 2420 8036 2454
rect 8002 2351 8036 2385
rect 8002 2282 8036 2316
rect 8002 2213 8036 2247
rect 8002 2144 8036 2178
rect 8002 2075 8036 2109
rect 8002 2006 8036 2040
rect 8002 1937 8036 1971
rect 8002 1868 8036 1902
rect 8002 1799 8036 1833
rect 8002 1730 8036 1764
rect 8002 1661 8036 1695
rect 8002 1592 8036 1626
rect 8002 1523 8036 1557
rect 8002 1454 8036 1488
rect 8002 1385 8036 1419
rect 8002 1316 8036 1350
rect 8002 1247 8036 1281
rect 8002 1178 8036 1212
rect 8002 1109 8036 1143
rect 8002 1040 8036 1074
rect 8002 971 8036 1005
rect 8002 902 8036 936
rect 8002 833 8036 867
rect 8002 764 8036 798
rect 8002 695 8036 729
rect 8002 626 8036 660
rect 8002 557 8036 591
rect 8002 488 8036 522
rect 8002 419 8036 453
rect 8002 350 8036 384
rect 8002 281 8036 315
rect 8002 212 8036 246
rect 8002 143 8036 177
rect 9752 39580 9786 39614
rect 9752 39512 9786 39546
rect 9752 39444 9786 39478
rect 9752 39376 9786 39410
rect 9752 39308 9786 39342
rect 9752 39240 9786 39274
rect 9752 39172 9786 39206
rect 9752 39104 9786 39138
rect 9752 39036 9786 39070
rect 9752 38968 9786 39002
rect 9752 38900 9786 38934
rect 9752 38832 9786 38866
rect 9752 38764 9786 38798
rect 9752 38696 9786 38730
rect 9752 38628 9786 38662
rect 9752 38560 9786 38594
rect 9752 38492 9786 38526
rect 9752 38424 9786 38458
rect 9752 38356 9786 38390
rect 9752 38288 9786 38322
rect 9752 38220 9786 38254
rect 9752 38152 9786 38186
rect 9752 38084 9786 38118
rect 9752 38016 9786 38050
rect 9752 37948 9786 37982
rect 9752 37880 9786 37914
rect 9752 37812 9786 37846
rect 9752 37744 9786 37778
rect 9752 37676 9786 37710
rect 9752 37608 9786 37642
rect 9752 37540 9786 37574
rect 9752 37472 9786 37506
rect 9752 37404 9786 37438
rect 9752 37336 9786 37370
rect 9752 37268 9786 37302
rect 9752 37200 9786 37234
rect 9752 37132 9786 37166
rect 9752 37064 9786 37098
rect 9752 36996 9786 37030
rect 9752 36928 9786 36962
rect 9752 36860 9786 36894
rect 9752 36792 9786 36826
rect 9752 36724 9786 36758
rect 9752 36656 9786 36690
rect 9752 36588 9786 36622
rect 9752 36520 9786 36554
rect 9752 36452 9786 36486
rect 9752 36384 9786 36418
rect 9752 36316 9786 36350
rect 9752 36248 9786 36282
rect 9752 36180 9786 36214
rect 9752 36112 9786 36146
rect 9752 36044 9786 36078
rect 9752 35976 9786 36010
rect 9752 35908 9786 35942
rect 9752 35840 9786 35874
rect 9752 35772 9786 35806
rect 9752 35704 9786 35738
rect 9752 35636 9786 35670
rect 9752 35568 9786 35602
rect 9752 35500 9786 35534
rect 9752 35432 9786 35466
rect 9752 35364 9786 35398
rect 9752 35296 9786 35330
rect 9752 35228 9786 35262
rect 9752 35160 9786 35194
rect 9752 35092 9786 35126
rect 9752 35024 9786 35058
rect 9752 34956 9786 34990
rect 9752 34888 9786 34922
rect 9752 34820 9786 34854
rect 9752 34752 9786 34786
rect 9752 34684 9786 34718
rect 9752 34616 9786 34650
rect 9752 34548 9786 34582
rect 9752 34480 9786 34514
rect 9752 34412 9786 34446
rect 9752 34344 9786 34378
rect 9752 34276 9786 34310
rect 9752 34208 9786 34242
rect 9752 34140 9786 34174
rect 9752 34072 9786 34106
rect 9752 34004 9786 34038
rect 9752 33936 9786 33970
rect 9752 33868 9786 33902
rect 9752 33800 9786 33834
rect 9752 33732 9786 33766
rect 9752 33664 9786 33698
rect 9752 33596 9786 33630
rect 9752 33528 9786 33562
rect 9752 33460 9786 33494
rect 9752 33392 9786 33426
rect 9752 33324 9786 33358
rect 9752 33256 9786 33290
rect 9752 33188 9786 33222
rect 9752 33120 9786 33154
rect 9752 33052 9786 33086
rect 9752 32984 9786 33018
rect 9752 32916 9786 32950
rect 9752 32848 9786 32882
rect 9752 32780 9786 32814
rect 9752 32712 9786 32746
rect 9752 32644 9786 32678
rect 9752 32576 9786 32610
rect 9752 32508 9786 32542
rect 9752 32440 9786 32474
rect 9752 32372 9786 32406
rect 9752 32304 9786 32338
rect 9752 32236 9786 32270
rect 9752 32168 9786 32202
rect 9752 32100 9786 32134
rect 9752 32032 9786 32066
rect 9752 31964 9786 31998
rect 9752 31896 9786 31930
rect 9752 31828 9786 31862
rect 9752 31760 9786 31794
rect 9752 31692 9786 31726
rect 9752 31624 9786 31658
rect 9752 31556 9786 31590
rect 9752 31488 9786 31522
rect 9752 31420 9786 31454
rect 9752 31352 9786 31386
rect 9752 31284 9786 31318
rect 9752 31216 9786 31250
rect 9752 31148 9786 31182
rect 9752 31080 9786 31114
rect 9752 31012 9786 31046
rect 9752 30944 9786 30978
rect 9752 30876 9786 30910
rect 9752 30808 9786 30842
rect 9752 30740 9786 30774
rect 9752 30672 9786 30706
rect 9752 30604 9786 30638
rect 9752 30536 9786 30570
rect 9752 30468 9786 30502
rect 9752 30400 9786 30434
rect 9752 30332 9786 30366
rect 9752 30264 9786 30298
rect 9752 30196 9786 30230
rect 9752 30128 9786 30162
rect 9752 30060 9786 30094
rect 9752 29992 9786 30026
rect 9752 29924 9786 29958
rect 9752 29856 9786 29890
rect 9752 29788 9786 29822
rect 9752 29720 9786 29754
rect 9752 29652 9786 29686
rect 9752 29584 9786 29618
rect 9752 29516 9786 29550
rect 9752 29448 9786 29482
rect 9752 29380 9786 29414
rect 9752 29312 9786 29346
rect 9752 29244 9786 29278
rect 9752 29176 9786 29210
rect 9752 29108 9786 29142
rect 9752 29040 9786 29074
rect 9752 28972 9786 29006
rect 9752 28904 9786 28938
rect 9752 28836 9786 28870
rect 9752 28768 9786 28802
rect 9752 28700 9786 28734
rect 9752 28632 9786 28666
rect 9752 28564 9786 28598
rect 9752 28496 9786 28530
rect 9752 28428 9786 28462
rect 9752 28360 9786 28394
rect 9752 28292 9786 28326
rect 9752 28224 9786 28258
rect 9752 28156 9786 28190
rect 9752 28088 9786 28122
rect 9752 28020 9786 28054
rect 9752 27952 9786 27986
rect 9752 27884 9786 27918
rect 9752 27816 9786 27850
rect 9752 27748 9786 27782
rect 9752 27680 9786 27714
rect 9752 27612 9786 27646
rect 9752 27544 9786 27578
rect 9752 27476 9786 27510
rect 9752 27408 9786 27442
rect 9752 27340 9786 27374
rect 9752 27272 9786 27306
rect 9752 27204 9786 27238
rect 9752 27136 9786 27170
rect 9752 27068 9786 27102
rect 9752 27000 9786 27034
rect 9752 26932 9786 26966
rect 9752 26864 9786 26898
rect 9752 26796 9786 26830
rect 9752 26728 9786 26762
rect 9752 26660 9786 26694
rect 9752 26592 9786 26626
rect 9752 26524 9786 26558
rect 9752 26456 9786 26490
rect 9752 26388 9786 26422
rect 9752 26320 9786 26354
rect 9752 26252 9786 26286
rect 9752 26184 9786 26218
rect 9752 26116 9786 26150
rect 9752 26048 9786 26082
rect 9752 25980 9786 26014
rect 9752 25912 9786 25946
rect 9752 25844 9786 25878
rect 9752 25776 9786 25810
rect 9752 25708 9786 25742
rect 9752 25640 9786 25674
rect 9752 25572 9786 25606
rect 9752 25504 9786 25538
rect 9752 25436 9786 25470
rect 9752 25368 9786 25402
rect 9752 25300 9786 25334
rect 9752 25232 9786 25266
rect 9752 25164 9786 25198
rect 9752 25096 9786 25130
rect 9752 25028 9786 25062
rect 9752 24960 9786 24994
rect 9752 24892 9786 24926
rect 9752 24824 9786 24858
rect 9752 24756 9786 24790
rect 9752 24688 9786 24722
rect 9752 24620 9786 24654
rect 9752 24552 9786 24586
rect 9752 24484 9786 24518
rect 9752 24416 9786 24450
rect 9752 24348 9786 24382
rect 9752 24280 9786 24314
rect 9752 24212 9786 24246
rect 9752 24144 9786 24178
rect 9752 24076 9786 24110
rect 9752 24008 9786 24042
rect 9752 23940 9786 23974
rect 9752 23872 9786 23906
rect 9752 23804 9786 23838
rect 9752 23736 9786 23770
rect 9752 23668 9786 23702
rect 9752 23600 9786 23634
rect 9752 23532 9786 23566
rect 9752 23464 9786 23498
rect 9752 23396 9786 23430
rect 9752 23328 9786 23362
rect 9752 23260 9786 23294
rect 9752 23192 9786 23226
rect 9752 23124 9786 23158
rect 9752 23056 9786 23090
rect 9752 22988 9786 23022
rect 9752 22920 9786 22954
rect 9752 22852 9786 22886
rect 9752 22784 9786 22818
rect 9752 22716 9786 22750
rect 9752 22648 9786 22682
rect 9752 22580 9786 22614
rect 9752 22512 9786 22546
rect 9752 22444 9786 22478
rect 9752 22376 9786 22410
rect 9752 22308 9786 22342
rect 9752 22240 9786 22274
rect 9752 22172 9786 22206
rect 9752 22104 9786 22138
rect 9752 22036 9786 22070
rect 9752 21968 9786 22002
rect 9752 21900 9786 21934
rect 9752 21832 9786 21866
rect 9752 21764 9786 21798
rect 9752 21696 9786 21730
rect 9752 21628 9786 21662
rect 9752 21560 9786 21594
rect 9752 21492 9786 21526
rect 9752 21424 9786 21458
rect 9752 21356 9786 21390
rect 9752 21288 9786 21322
rect 9752 21220 9786 21254
rect 9752 21152 9786 21186
rect 9752 21084 9786 21118
rect 9752 21016 9786 21050
rect 9752 20948 9786 20982
rect 9752 20880 9786 20914
rect 9752 20812 9786 20846
rect 9752 20744 9786 20778
rect 9752 20676 9786 20710
rect 9752 20608 9786 20642
rect 9752 20540 9786 20574
rect 9752 20472 9786 20506
rect 9752 20404 9786 20438
rect 9752 20336 9786 20370
rect 9752 20268 9786 20302
rect 9752 20200 9786 20234
rect 9752 20132 9786 20166
rect 9752 20064 9786 20098
rect 9752 19996 9786 20030
rect 9752 19928 9786 19962
rect 9752 19860 9786 19894
rect 9752 19792 9786 19826
rect 9752 19724 9786 19758
rect 9752 19656 9786 19690
rect 9752 19588 9786 19622
rect 9752 19520 9786 19554
rect 9752 19452 9786 19486
rect 9752 19384 9786 19418
rect 9752 19316 9786 19350
rect 9752 19248 9786 19282
rect 9752 19180 9786 19214
rect 9752 19112 9786 19146
rect 9752 19044 9786 19078
rect 9752 18976 9786 19010
rect 9752 18908 9786 18942
rect 9752 18840 9786 18874
rect 9752 18772 9786 18806
rect 9752 18704 9786 18738
rect 9752 18636 9786 18670
rect 9752 18568 9786 18602
rect 9752 18500 9786 18534
rect 9752 18432 9786 18466
rect 9752 18364 9786 18398
rect 9752 18296 9786 18330
rect 9752 18228 9786 18262
rect 9752 18160 9786 18194
rect 9752 18092 9786 18126
rect 9752 18024 9786 18058
rect 9752 17956 9786 17990
rect 9752 17888 9786 17922
rect 9752 17820 9786 17854
rect 9752 17752 9786 17786
rect 9752 17684 9786 17718
rect 9752 17616 9786 17650
rect 9752 17548 9786 17582
rect 9752 17480 9786 17514
rect 9752 17412 9786 17446
rect 9752 17344 9786 17378
rect 9752 17276 9786 17310
rect 9752 17208 9786 17242
rect 9752 17140 9786 17174
rect 9752 17072 9786 17106
rect 9752 17004 9786 17038
rect 9752 16936 9786 16970
rect 9752 16868 9786 16902
rect 9752 16800 9786 16834
rect 9752 16732 9786 16766
rect 9752 16664 9786 16698
rect 9752 16596 9786 16630
rect 9752 16528 9786 16562
rect 9752 16460 9786 16494
rect 9752 16392 9786 16426
rect 9752 16324 9786 16358
rect 9752 16256 9786 16290
rect 9752 16188 9786 16222
rect 9752 16120 9786 16154
rect 9752 16052 9786 16086
rect 9752 15984 9786 16018
rect 9752 15916 9786 15950
rect 9752 15848 9786 15882
rect 9752 15780 9786 15814
rect 9752 15712 9786 15746
rect 9752 15644 9786 15678
rect 9752 15576 9786 15610
rect 9752 15508 9786 15542
rect 9752 15440 9786 15474
rect 9752 15372 9786 15406
rect 9752 15304 9786 15338
rect 9752 15236 9786 15270
rect 9752 15168 9786 15202
rect 9752 15100 9786 15134
rect 9752 15032 9786 15066
rect 9752 14964 9786 14998
rect 9752 14896 9786 14930
rect 9752 14828 9786 14862
rect 9752 14760 9786 14794
rect 9752 14692 9786 14726
rect 9752 14624 9786 14658
rect 9752 14556 9786 14590
rect 9752 14488 9786 14522
rect 9752 14420 9786 14454
rect 9752 14352 9786 14386
rect 9752 14284 9786 14318
rect 9752 14216 9786 14250
rect 9752 14148 9786 14182
rect 9752 14080 9786 14114
rect 9752 14012 9786 14046
rect 9752 13944 9786 13978
rect 9752 13876 9786 13910
rect 9752 13808 9786 13842
rect 9752 13740 9786 13774
rect 9752 13672 9786 13706
rect 9752 13604 9786 13638
rect 9752 13536 9786 13570
rect 9752 13468 9786 13502
rect 9752 13400 9786 13434
rect 9752 13332 9786 13366
rect 9752 13264 9786 13298
rect 9752 13196 9786 13230
rect 9752 13128 9786 13162
rect 9752 13060 9786 13094
rect 9752 12992 9786 13026
rect 9752 12924 9786 12958
rect 9752 12856 9786 12890
rect 9752 12788 9786 12822
rect 9752 12720 9786 12754
rect 9752 12652 9786 12686
rect 9752 12584 9786 12618
rect 9752 12516 9786 12550
rect 9752 12448 9786 12482
rect 9752 12380 9786 12414
rect 9752 12312 9786 12346
rect 9752 12244 9786 12278
rect 9752 12176 9786 12210
rect 9752 12108 9786 12142
rect 9752 12040 9786 12074
rect 9752 11972 9786 12006
rect 9752 11904 9786 11938
rect 9752 11836 9786 11870
rect 9752 11768 9786 11802
rect 9752 11700 9786 11734
rect 9752 11632 9786 11666
rect 9752 11564 9786 11598
rect 9752 11496 9786 11530
rect 9752 11428 9786 11462
rect 9752 11360 9786 11394
rect 9752 11292 9786 11326
rect 9752 11224 9786 11258
rect 9752 11156 9786 11190
rect 9752 11088 9786 11122
rect 9752 11020 9786 11054
rect 9752 10952 9786 10986
rect 9752 10884 9786 10918
rect 9752 10816 9786 10850
rect 9752 10748 9786 10782
rect 9752 10680 9786 10714
rect 9752 10612 9786 10646
rect 9752 10544 9786 10578
rect 9752 10476 9786 10510
rect 9752 10408 9786 10442
rect 9752 10340 9786 10374
rect 9752 10272 9786 10306
rect 9752 10204 9786 10238
rect 9752 10136 9786 10170
rect 9752 10068 9786 10102
rect 9752 10000 9786 10034
rect 9752 9932 9786 9966
rect 9752 9864 9786 9898
rect 9752 9796 9786 9830
rect 9752 9728 9786 9762
rect 9752 9660 9786 9694
rect 9752 9592 9786 9626
rect 9752 9524 9786 9558
rect 9752 9456 9786 9490
rect 9752 9388 9786 9422
rect 9752 9320 9786 9354
rect 9752 9252 9786 9286
rect 9752 9184 9786 9218
rect 9752 9116 9786 9150
rect 9752 9048 9786 9082
rect 9752 8980 9786 9014
rect 9752 8912 9786 8946
rect 9752 8844 9786 8878
rect 9752 8776 9786 8810
rect 9752 8708 9786 8742
rect 9752 8640 9786 8674
rect 9752 8572 9786 8606
rect 9752 8504 9786 8538
rect 9752 8436 9786 8470
rect 9752 8368 9786 8402
rect 9752 8300 9786 8334
rect 9752 8232 9786 8266
rect 9752 8164 9786 8198
rect 9752 8096 9786 8130
rect 9752 8028 9786 8062
rect 9752 7960 9786 7994
rect 9752 7892 9786 7926
rect 9752 7824 9786 7858
rect 9752 7756 9786 7790
rect 9752 7688 9786 7722
rect 9752 7620 9786 7654
rect 9752 7552 9786 7586
rect 9752 7484 9786 7518
rect 9752 7416 9786 7450
rect 9752 7348 9786 7382
rect 9752 7280 9786 7314
rect 9752 7212 9786 7246
rect 9752 7144 9786 7178
rect 9752 7076 9786 7110
rect 9752 7008 9786 7042
rect 9752 6940 9786 6974
rect 9752 6872 9786 6906
rect 9752 6804 9786 6838
rect 9752 6736 9786 6770
rect 9752 6668 9786 6702
rect 9752 6600 9786 6634
rect 9752 6532 9786 6566
rect 9752 6464 9786 6498
rect 9752 6396 9786 6430
rect 9752 6328 9786 6362
rect 9752 6260 9786 6294
rect 9752 6192 9786 6226
rect 9752 6124 9786 6158
rect 9752 6056 9786 6090
rect 9752 5988 9786 6022
rect 9752 5920 9786 5954
rect 9752 5852 9786 5886
rect 9752 5784 9786 5818
rect 9752 5716 9786 5750
rect 9752 5648 9786 5682
rect 9752 5580 9786 5614
rect 9752 5512 9786 5546
rect 9752 5444 9786 5478
rect 9752 5376 9786 5410
rect 9752 5308 9786 5342
rect 9752 5240 9786 5274
rect 9752 5172 9786 5206
rect 9752 5104 9786 5138
rect 9752 5036 9786 5070
rect 9752 4968 9786 5002
rect 9752 4900 9786 4934
rect 9752 4832 9786 4866
rect 9752 4764 9786 4798
rect 9752 4696 9786 4730
rect 9752 4628 9786 4662
rect 9752 4560 9786 4594
rect 9752 4492 9786 4526
rect 9752 4424 9786 4458
rect 9752 4356 9786 4390
rect 9752 4288 9786 4322
rect 9752 4220 9786 4254
rect 9752 4152 9786 4186
rect 9752 4084 9786 4118
rect 9752 4016 9786 4050
rect 9752 3948 9786 3982
rect 9752 3880 9786 3914
rect 9752 3812 9786 3846
rect 9752 3744 9786 3778
rect 9752 3676 9786 3710
rect 9752 3608 9786 3642
rect 9752 3540 9786 3574
rect 9752 3472 9786 3506
rect 9752 3404 9786 3438
rect 9752 3336 9786 3370
rect 9752 3268 9786 3302
rect 9752 3200 9786 3234
rect 9752 3132 9786 3166
rect 9752 3064 9786 3098
rect 9752 2996 9786 3030
rect 9752 2928 9786 2962
rect 9752 2860 9786 2894
rect 9752 2792 9786 2826
rect 9752 2724 9786 2758
rect 9752 2656 9786 2690
rect 9752 2588 9786 2622
rect 9752 2520 9786 2554
rect 9752 2452 9786 2486
rect 9752 2384 9786 2418
rect 9752 2315 9786 2349
rect 9752 2246 9786 2280
rect 9752 2177 9786 2211
rect 9752 2108 9786 2142
rect 9752 2039 9786 2073
rect 9752 1970 9786 2004
rect 9752 1901 9786 1935
rect 9752 1832 9786 1866
rect 9752 1763 9786 1797
rect 9752 1694 9786 1728
rect 9752 1625 9786 1659
rect 9752 1556 9786 1590
rect 9752 1487 9786 1521
rect 9752 1418 9786 1452
rect 9752 1349 9786 1383
rect 9752 1280 9786 1314
rect 9752 1211 9786 1245
rect 9752 1142 9786 1176
rect 9752 1073 9786 1107
rect 9752 1004 9786 1038
rect 9752 935 9786 969
rect 9752 866 9786 900
rect 9752 797 9786 831
rect 9752 728 9786 762
rect 9752 659 9786 693
rect 9752 590 9786 624
rect 9752 521 9786 555
rect 9752 452 9786 486
rect 9752 383 9786 417
rect 9752 314 9786 348
rect 9752 245 9786 279
rect 9752 176 9786 210
rect 10786 39752 10820 39786
rect 2482 40 2516 74
rect 8002 74 8036 108
rect 8096 40 10646 142
rect 10718 108 10820 39718
rect 10680 40 10714 74
<< mvnsubdiffcont >>
rect 6520 22085 6554 22119
rect 6588 22085 6622 22119
rect 6656 22085 6690 22119
rect 6724 22085 6758 22119
rect 2926 11365 2960 11399
rect 2994 11365 3028 11399
rect 3062 11365 3096 11399
rect 3130 11365 3164 11399
rect 3198 11365 3232 11399
rect 3266 11365 3300 11399
rect 3334 11365 3368 11399
rect 3402 11365 3436 11399
rect 3470 11365 3504 11399
rect 3538 11365 3572 11399
rect 3606 11365 3640 11399
rect 3674 11365 3708 11399
rect 3742 11365 3776 11399
rect 3810 11365 3844 11399
rect 3878 11365 3912 11399
rect 3946 11365 3980 11399
rect 4014 11365 4048 11399
rect 4082 11365 4116 11399
rect 4150 11365 4184 11399
rect 4218 11365 4252 11399
rect 4286 11365 4320 11399
rect 4354 11365 4388 11399
rect 4422 11365 4456 11399
rect 4490 11365 4524 11399
rect 4558 11365 4592 11399
rect 4626 11365 4660 11399
rect 4694 11365 4728 11399
rect 4762 11365 4796 11399
rect 4830 11365 4864 11399
rect 4898 11365 4932 11399
rect 4966 11365 5000 11399
rect 5034 11365 5068 11399
rect 5102 11365 5136 11399
rect 5170 11365 5204 11399
rect 5238 11365 5272 11399
rect 5306 11365 5340 11399
rect 5374 11365 5408 11399
rect 5442 11365 5476 11399
rect 5510 11365 5544 11399
rect 5578 11365 5612 11399
rect 5646 11365 5680 11399
rect 5714 11365 5748 11399
rect 5782 11365 5816 11399
rect 5850 11365 5884 11399
rect 5918 11365 5952 11399
rect 5986 11365 6020 11399
rect 6054 11365 6088 11399
rect 6122 11365 6156 11399
rect 6190 11365 6224 11399
rect 6258 11365 6292 11399
rect 6326 11365 6360 11399
rect 6394 11365 6428 11399
rect 6553 11365 6587 11399
rect 6621 11365 6655 11399
rect 6689 11365 6723 11399
rect 6757 11365 6791 11399
rect 6825 11365 6859 11399
rect 6893 11365 6927 11399
rect 6961 11365 6995 11399
rect 7029 11365 7063 11399
rect 7097 11365 7131 11399
rect 7165 11365 7199 11399
rect 7233 11365 7267 11399
rect 7301 11365 7335 11399
rect 7369 11365 7403 11399
rect 2802 11297 2836 11331
rect 2802 11229 2836 11263
rect 2802 11161 2836 11195
rect 2802 11093 2836 11127
rect 2802 11025 2836 11059
rect 2802 10957 2836 10991
rect 2802 10889 2836 10923
rect 2802 10821 2836 10855
rect 2802 10753 2836 10787
rect 2802 10685 2836 10719
rect 2802 10617 2836 10651
rect 2802 10549 2836 10583
rect 2802 10481 2836 10515
rect 2802 10413 2836 10447
rect 2802 10345 2836 10379
rect 2802 10277 2836 10311
rect 2802 10209 2836 10243
rect 2802 10141 2836 10175
rect 2802 10073 2836 10107
rect 2802 10005 2836 10039
rect 2802 9937 2836 9971
rect 2802 9869 2836 9903
rect 2802 9801 2836 9835
rect 2802 9733 2836 9767
rect 2802 9665 2836 9699
rect 2802 9597 2836 9631
rect 2802 9529 2836 9563
rect 2802 9461 2836 9495
rect 2802 9393 2836 9427
rect 2802 9325 2836 9359
rect 2802 9257 2836 9291
rect 2802 9189 2836 9223
rect 2802 9121 2836 9155
rect 2802 9053 2836 9087
rect 2802 8985 2836 9019
rect 2802 8917 2836 8951
rect 2802 8849 2836 8883
rect 2802 8781 2836 8815
rect 2802 8713 2836 8747
rect 2802 8645 2836 8679
rect 2802 8577 2836 8611
rect 2802 8509 2836 8543
rect 2802 8441 2836 8475
rect 2802 8373 2836 8407
rect 2802 8305 2836 8339
rect 2802 8237 2836 8271
rect 2802 8169 2836 8203
rect 2802 8101 2836 8135
rect 7437 11284 7471 11318
rect 7437 11216 7471 11250
rect 7437 11148 7471 11182
rect 7437 11080 7471 11114
rect 7437 11012 7471 11046
rect 7437 10944 7471 10978
rect 7437 10876 7471 10910
rect 7437 10808 7471 10842
rect 7437 10740 7471 10774
rect 7437 10672 7471 10706
rect 7437 10604 7471 10638
rect 7437 10536 7471 10570
rect 7437 10468 7471 10502
rect 7437 10400 7471 10434
rect 7437 10332 7471 10366
rect 7437 10264 7471 10298
rect 7437 10196 7471 10230
rect 7437 10128 7471 10162
rect 7437 10060 7471 10094
rect 7437 9992 7471 10026
rect 7437 9924 7471 9958
rect 7437 9856 7471 9890
rect 7437 9788 7471 9822
rect 7437 9720 7471 9754
rect 7437 9652 7471 9686
rect 7437 9584 7471 9618
rect 7437 9438 7471 9472
rect 7437 9370 7471 9404
rect 7437 9302 7471 9336
rect 7437 9234 7471 9268
rect 7437 9166 7471 9200
rect 7437 9098 7471 9132
rect 7437 9030 7471 9064
rect 7437 8962 7471 8996
rect 7437 8894 7471 8928
rect 7437 8826 7471 8860
rect 7437 8758 7471 8792
rect 7437 8690 7471 8724
rect 7437 8622 7471 8656
rect 7437 8554 7471 8588
rect 7437 8486 7471 8520
rect 7437 8418 7471 8452
rect 7437 8350 7471 8384
rect 7437 8282 7471 8316
rect 7437 8214 7471 8248
rect 7437 8146 7471 8180
rect 2802 8033 2836 8067
rect 2802 7965 2836 7999
rect 2802 7897 2836 7931
rect 6862 8078 6896 8112
rect 6930 8078 6964 8112
rect 6998 8078 7032 8112
rect 7100 8078 7134 8112
rect 7168 8078 7202 8112
rect 7236 8078 7270 8112
rect 7304 8078 7338 8112
rect 6750 8010 6784 8044
rect 2870 7886 2904 7920
rect 2938 7886 2972 7920
rect 3006 7886 3040 7920
rect 3074 7886 3108 7920
rect 3142 7886 3176 7920
rect 3210 7886 3244 7920
rect 3278 7886 3312 7920
rect 3346 7886 3380 7920
rect 3414 7886 3448 7920
rect 3482 7886 3516 7920
rect 3550 7886 3584 7920
rect 3618 7886 3652 7920
rect 3686 7886 3720 7920
rect 3754 7886 3788 7920
rect 3822 7886 3856 7920
rect 3890 7886 3924 7920
rect 3958 7886 3992 7920
rect 4026 7886 4060 7920
rect 4094 7886 4128 7920
rect 4162 7886 4196 7920
rect 4230 7886 4264 7920
rect 4298 7886 4332 7920
rect 4366 7886 4400 7920
rect 4434 7886 4468 7920
rect 4502 7886 4536 7920
rect 4570 7886 4604 7920
rect 4638 7886 4672 7920
rect 4706 7886 4740 7920
rect 4774 7886 4808 7920
rect 4842 7886 4876 7920
rect 4910 7886 4944 7920
rect 4978 7886 5012 7920
rect 5046 7886 5080 7920
rect 5114 7886 5148 7920
rect 5182 7886 5216 7920
rect 5250 7886 5284 7920
rect 5318 7886 5352 7920
rect 5386 7886 5420 7920
rect 5454 7886 5488 7920
rect 5522 7886 5556 7920
rect 5590 7886 5624 7920
rect 5658 7886 5692 7920
rect 5726 7886 5760 7920
rect 5794 7886 5828 7920
rect 5862 7886 5896 7920
rect 5930 7886 5964 7920
rect 5998 7886 6032 7920
rect 6066 7886 6100 7920
rect 6134 7886 6168 7920
rect 6202 7886 6236 7920
rect 6270 7886 6304 7920
rect 6338 7886 6372 7920
rect 6406 7886 6440 7920
rect 6474 7886 6508 7920
rect 6542 7886 6576 7920
rect 6610 7886 6644 7920
rect 6678 7886 6712 7920
rect 2802 7829 2836 7863
rect 2802 7761 2836 7795
rect 2802 7693 2836 7727
rect 6750 7863 6784 7897
rect 6750 7795 6784 7829
rect 6750 7727 6784 7761
rect 2802 7625 2836 7659
rect 2802 7557 2836 7591
rect 2802 7489 2836 7523
rect 2802 7421 2836 7455
rect 2802 7353 2836 7387
rect 2802 7285 2836 7319
rect 2802 7217 2836 7251
rect 2802 7149 2836 7183
rect 2802 7081 2836 7115
rect 2802 7013 2836 7047
rect 2802 6945 2836 6979
rect 2802 6877 2836 6911
rect 2802 6809 2836 6843
rect 2802 6741 2836 6775
rect 2802 6673 2836 6707
rect 2802 6605 2836 6639
rect 2802 6537 2836 6571
rect 2802 6469 2836 6503
rect 2802 6401 2836 6435
rect 2802 6333 2836 6367
rect 2802 6265 2836 6299
rect 2802 6197 2836 6231
rect 2802 6129 2836 6163
rect 2802 6061 2836 6095
rect 2802 5993 2836 6027
rect 2802 5925 2836 5959
rect 2802 5857 2836 5891
rect 2802 5789 2836 5823
rect 2802 5721 2836 5755
rect 2802 5653 2836 5687
rect 2802 5585 2836 5619
rect 2802 5517 2836 5551
rect 2802 5449 2836 5483
rect 2802 5381 2836 5415
rect 2802 5313 2836 5347
rect 2802 5245 2836 5279
rect 6750 7659 6784 7693
rect 6750 7591 6784 7625
rect 6750 7523 6784 7557
rect 6750 7455 6784 7489
rect 6750 7387 6784 7421
rect 6750 7319 6784 7353
rect 6750 7251 6784 7285
rect 6750 7183 6784 7217
rect 6750 7115 6784 7149
rect 6750 7047 6784 7081
rect 6750 6979 6784 7013
rect 6750 6911 6784 6945
rect 6750 6843 6784 6877
rect 6750 6775 6784 6809
rect 6750 6707 6784 6741
rect 6750 6639 6784 6673
rect 6750 6571 6784 6605
rect 6750 6503 6784 6537
rect 6750 6435 6784 6469
rect 6750 6367 6784 6401
rect 6750 6299 6784 6333
rect 6750 6231 6784 6265
rect 6750 6163 6784 6197
rect 6750 6095 6784 6129
rect 6750 6027 6784 6061
rect 6750 5959 6784 5993
rect 6750 5891 6784 5925
rect 6750 5823 6784 5857
rect 6750 5755 6784 5789
rect 6750 5687 6784 5721
rect 6750 5619 6784 5653
rect 6750 5551 6784 5585
rect 6750 5483 6784 5517
rect 6750 5415 6784 5449
rect 6750 5347 6784 5381
rect 6750 5279 6784 5313
rect 2802 5109 2836 5143
rect 6750 5211 6784 5245
rect 6750 5143 6784 5177
rect 6750 5075 6784 5109
rect 2870 5007 2904 5041
rect 2938 5007 2972 5041
rect 3006 5007 3040 5041
rect 3074 5007 3108 5041
rect 3142 5007 3176 5041
rect 3210 5007 3244 5041
rect 3278 5007 3312 5041
rect 3346 5007 3380 5041
rect 3414 5007 3448 5041
rect 3482 5007 3516 5041
rect 3550 5007 3584 5041
rect 3618 5007 3652 5041
rect 3686 5007 3720 5041
rect 3754 5007 3788 5041
rect 3822 5007 3856 5041
rect 3890 5007 3924 5041
rect 3958 5007 3992 5041
rect 4026 5007 4060 5041
rect 4094 5007 4128 5041
rect 4162 5007 4196 5041
rect 4230 5007 4264 5041
rect 4298 5007 4332 5041
rect 4366 5007 4400 5041
rect 4434 5007 4468 5041
rect 4502 5007 4536 5041
rect 4570 5007 4604 5041
rect 4638 5007 4672 5041
rect 4706 5007 4740 5041
rect 4774 5007 4808 5041
rect 4842 5007 4876 5041
rect 4910 5007 4944 5041
rect 4978 5007 5012 5041
rect 5046 5007 5080 5041
rect 5114 5007 5148 5041
rect 5182 5007 5216 5041
rect 5250 5007 5284 5041
rect 5318 5007 5352 5041
rect 5386 5007 5420 5041
rect 5454 5007 5488 5041
rect 5522 5007 5556 5041
rect 5590 5007 5624 5041
rect 5658 5007 5692 5041
rect 5726 5007 5760 5041
rect 5794 5007 5828 5041
rect 5862 5007 5896 5041
rect 5930 5007 5964 5041
rect 5998 5007 6032 5041
rect 6066 5007 6100 5041
rect 6134 5007 6168 5041
rect 6202 5007 6236 5041
rect 6270 5007 6304 5041
rect 6338 5007 6372 5041
rect 6406 5007 6440 5041
rect 6474 5007 6508 5041
rect 6542 5007 6576 5041
rect 6610 5007 6644 5041
rect 6678 5007 6712 5041
rect 2887 4860 2921 4894
rect 2955 4860 2989 4894
rect 3023 4860 3057 4894
rect 3091 4860 3125 4894
rect 3159 4860 3193 4894
rect 3227 4860 3261 4894
rect 3295 4860 3329 4894
rect 3363 4860 3397 4894
rect 3431 4860 3465 4894
rect 3499 4860 3533 4894
rect 3567 4860 3601 4894
rect 3635 4860 3669 4894
rect 3703 4860 3737 4894
rect 3771 4860 3805 4894
rect 3839 4860 3873 4894
rect 3907 4860 3941 4894
rect 3975 4860 4009 4894
rect 4043 4860 4077 4894
rect 4111 4860 4145 4894
rect 4179 4860 4213 4894
rect 4247 4860 4281 4894
rect 4315 4860 4349 4894
rect 4383 4860 4417 4894
rect 4451 4860 4485 4894
rect 4519 4860 4553 4894
rect 4587 4860 4621 4894
rect 4655 4860 4689 4894
rect 4723 4860 4757 4894
rect 4791 4860 4825 4894
rect 4859 4860 4893 4894
rect 4927 4860 4961 4894
rect 4995 4860 5029 4894
rect 5063 4860 5097 4894
rect 5131 4860 5165 4894
rect 5199 4860 5233 4894
rect 5267 4860 5301 4894
rect 5335 4860 5369 4894
rect 5403 4860 5437 4894
rect 5471 4860 5505 4894
rect 5539 4860 5573 4894
rect 5607 4860 5641 4894
rect 5675 4860 5709 4894
rect 5743 4860 5777 4894
rect 5811 4860 5845 4894
rect 5879 4860 5913 4894
rect 5947 4860 5981 4894
rect 6015 4860 6049 4894
rect 6083 4860 6117 4894
rect 6151 4860 6185 4894
rect 6219 4860 6253 4894
rect 6287 4860 6321 4894
rect 6355 4860 6389 4894
rect 6423 4860 6457 4894
rect 6491 4860 6525 4894
rect 6559 4860 6593 4894
rect 6627 4860 6661 4894
rect 6695 4860 6729 4894
rect 2778 3124 2812 3158
rect 2846 3124 2880 3158
rect 2914 3124 2948 3158
rect 2982 3124 3016 3158
rect 3050 3124 3084 3158
rect 3118 3124 3152 3158
rect 3186 3124 3220 3158
rect 3254 3124 3288 3158
rect 3322 3124 3356 3158
rect 3390 3124 3424 3158
rect 3458 3124 3492 3158
rect 3526 3124 3560 3158
rect 3594 3124 3628 3158
rect 3662 3124 3696 3158
rect 3730 3124 3764 3158
rect 3798 3124 3832 3158
<< poly >>
rect 8132 39651 8198 39667
rect 8132 39617 8148 39651
rect 8182 39617 8198 39651
rect 8132 39595 8198 39617
rect 9590 39651 9656 39667
rect 9590 39617 9606 39651
rect 9640 39617 9656 39651
rect 9590 39595 9656 39617
rect 7516 39431 7582 39447
rect 7516 39397 7532 39431
rect 7566 39397 7582 39431
rect 7516 39363 7582 39397
rect 7516 39329 7532 39363
rect 7566 39329 7582 39363
rect 7516 39295 7582 39329
rect 7516 39261 7532 39295
rect 7566 39261 7582 39295
rect 7516 39227 7582 39261
rect 7516 39193 7532 39227
rect 7566 39193 7582 39227
rect 7516 39159 7582 39193
rect 7516 39125 7532 39159
rect 7566 39125 7582 39159
rect 7516 39091 7582 39125
rect 7516 39057 7532 39091
rect 7566 39057 7582 39091
rect 7516 39023 7582 39057
rect 7516 38989 7532 39023
rect 7566 38989 7582 39023
rect 7516 38955 7582 38989
rect 7516 38921 7532 38955
rect 7566 38921 7582 38955
rect 7516 38887 7582 38921
rect 7516 38853 7532 38887
rect 7566 38853 7582 38887
rect 7516 38819 7582 38853
rect 7516 38785 7532 38819
rect 7566 38785 7582 38819
rect 7516 38751 7582 38785
rect 7516 38717 7532 38751
rect 7566 38717 7582 38751
rect 7516 38683 7582 38717
rect 7516 38649 7532 38683
rect 7566 38649 7582 38683
rect 7516 38615 7582 38649
rect 7516 38581 7532 38615
rect 7566 38581 7582 38615
rect 7516 38547 7582 38581
rect 7516 38513 7532 38547
rect 7566 38513 7582 38547
rect 7516 38479 7582 38513
rect 7516 38445 7532 38479
rect 7566 38445 7582 38479
rect 7516 38411 7582 38445
rect 7516 38377 7532 38411
rect 7566 38377 7582 38411
rect 7516 38343 7582 38377
rect 7516 38309 7532 38343
rect 7566 38309 7582 38343
rect 7516 38275 7582 38309
rect 7516 38241 7532 38275
rect 7566 38241 7582 38275
rect 7516 38207 7582 38241
rect 7516 38173 7532 38207
rect 7566 38173 7582 38207
rect 7516 38139 7582 38173
rect 7516 38105 7532 38139
rect 7566 38105 7582 38139
rect 7516 38071 7582 38105
rect 7516 38037 7532 38071
rect 7566 38037 7582 38071
rect 7516 38003 7582 38037
rect 7516 37969 7532 38003
rect 7566 37969 7582 38003
rect 7516 37935 7582 37969
rect 7516 37901 7532 37935
rect 7566 37901 7582 37935
rect 7516 37867 7582 37901
rect 7516 37833 7532 37867
rect 7566 37833 7582 37867
rect 7516 37799 7582 37833
rect 7516 37765 7532 37799
rect 7566 37765 7582 37799
rect 7516 37731 7582 37765
rect 7516 37697 7532 37731
rect 7566 37697 7582 37731
rect 7516 37663 7582 37697
rect 7516 37629 7532 37663
rect 7566 37629 7582 37663
rect 7516 37595 7582 37629
rect 7516 37561 7532 37595
rect 7566 37561 7582 37595
rect 7516 37527 7582 37561
rect 7516 37493 7532 37527
rect 7566 37493 7582 37527
rect 7516 37459 7582 37493
rect 7516 37425 7532 37459
rect 7566 37425 7582 37459
rect 7516 37391 7582 37425
rect 7516 37357 7532 37391
rect 7566 37357 7582 37391
rect 7516 37323 7582 37357
rect 7516 37289 7532 37323
rect 7566 37289 7582 37323
rect 7516 37255 7582 37289
rect 7516 37221 7532 37255
rect 7566 37221 7582 37255
rect 7516 37187 7582 37221
rect 7516 37153 7532 37187
rect 7566 37153 7582 37187
rect 7516 37119 7582 37153
rect 7516 37085 7532 37119
rect 7566 37085 7582 37119
rect 7516 37051 7582 37085
rect 7516 37017 7532 37051
rect 7566 37017 7582 37051
rect 7516 36983 7582 37017
rect 7516 36949 7532 36983
rect 7566 36949 7582 36983
rect 7516 36915 7582 36949
rect 7516 36881 7532 36915
rect 7566 36881 7582 36915
rect 7516 36847 7582 36881
rect 7516 36813 7532 36847
rect 7566 36813 7582 36847
rect 7516 36779 7582 36813
rect 7516 36745 7532 36779
rect 7566 36745 7582 36779
rect 7516 36711 7582 36745
rect 7516 36677 7532 36711
rect 7566 36677 7582 36711
rect 7516 36643 7582 36677
rect 7516 36609 7532 36643
rect 7566 36609 7582 36643
rect 7516 36575 7582 36609
rect 7516 36541 7532 36575
rect 7566 36541 7582 36575
rect 7516 36507 7582 36541
rect 7516 36473 7532 36507
rect 7566 36473 7582 36507
rect 7516 36439 7582 36473
rect 7516 36405 7532 36439
rect 7566 36405 7582 36439
rect 7516 36370 7582 36405
rect 7516 36336 7532 36370
rect 7566 36336 7582 36370
rect 7516 36301 7582 36336
rect 7516 36267 7532 36301
rect 7566 36267 7582 36301
rect 7516 36232 7582 36267
rect 7516 36198 7532 36232
rect 7566 36198 7582 36232
rect 7516 36163 7582 36198
rect 7516 36129 7532 36163
rect 7566 36129 7582 36163
rect 7516 36094 7582 36129
rect 7516 36060 7532 36094
rect 7566 36060 7582 36094
rect 7516 36025 7582 36060
rect 7516 35991 7532 36025
rect 7566 35991 7582 36025
rect 7516 35956 7582 35991
rect 7516 35922 7532 35956
rect 7566 35922 7582 35956
rect 7516 35887 7582 35922
rect 7516 35853 7532 35887
rect 7566 35853 7582 35887
rect 7516 35818 7582 35853
rect 7516 35784 7532 35818
rect 7566 35784 7582 35818
rect 7516 35749 7582 35784
rect 7516 35715 7532 35749
rect 7566 35715 7582 35749
rect 7516 35680 7582 35715
rect 7516 35646 7532 35680
rect 7566 35646 7582 35680
rect 7516 35611 7582 35646
rect 7516 35577 7532 35611
rect 7566 35577 7582 35611
rect 7516 35542 7582 35577
rect 7516 35508 7532 35542
rect 7566 35508 7582 35542
rect 7516 35473 7582 35508
rect 7516 35439 7532 35473
rect 7566 35439 7582 35473
rect 7516 35404 7582 35439
rect 7516 35370 7532 35404
rect 7566 35370 7582 35404
rect 7516 35335 7582 35370
rect 7516 35301 7532 35335
rect 7566 35301 7582 35335
rect 7516 35266 7582 35301
rect 7516 35232 7532 35266
rect 7566 35232 7582 35266
rect 7516 35197 7582 35232
rect 7516 35163 7532 35197
rect 7566 35163 7582 35197
rect 7516 35128 7582 35163
rect 7516 35094 7532 35128
rect 7566 35094 7582 35128
rect 7516 35059 7582 35094
rect 7516 35025 7532 35059
rect 7566 35025 7582 35059
rect 7516 34990 7582 35025
rect 7516 34956 7532 34990
rect 7566 34956 7582 34990
rect 7516 34921 7582 34956
rect 7516 34887 7532 34921
rect 7566 34887 7582 34921
rect 7516 34852 7582 34887
rect 7516 34818 7532 34852
rect 7566 34818 7582 34852
rect 7516 34783 7582 34818
rect 7516 34749 7532 34783
rect 7566 34749 7582 34783
rect 7516 34714 7582 34749
rect 7516 34680 7532 34714
rect 7566 34680 7582 34714
rect 7516 34645 7582 34680
rect 7516 34611 7532 34645
rect 7566 34611 7582 34645
rect 7516 34576 7582 34611
rect 7516 34542 7532 34576
rect 7566 34542 7582 34576
rect 7516 34507 7582 34542
rect 7516 34473 7532 34507
rect 7566 34473 7582 34507
rect 7516 34438 7582 34473
rect 7516 34404 7532 34438
rect 7566 34404 7582 34438
rect 7516 34369 7582 34404
rect 7516 34335 7532 34369
rect 7566 34335 7582 34369
rect 7516 34300 7582 34335
rect 7516 34266 7532 34300
rect 7566 34266 7582 34300
rect 7516 34231 7582 34266
rect 7516 34197 7532 34231
rect 7566 34197 7582 34231
rect 7516 34162 7582 34197
rect 7516 34128 7532 34162
rect 7566 34128 7582 34162
rect 7516 34093 7582 34128
rect 7516 34059 7532 34093
rect 7566 34059 7582 34093
rect 7516 34024 7582 34059
rect 7516 33990 7532 34024
rect 7566 33990 7582 34024
rect 7516 33955 7582 33990
rect 7516 33921 7532 33955
rect 7566 33921 7582 33955
rect 7516 33886 7582 33921
rect 7516 33852 7532 33886
rect 7566 33852 7582 33886
rect 7516 33817 7582 33852
rect 7516 33783 7532 33817
rect 7566 33783 7582 33817
rect 7516 33748 7582 33783
rect 7516 33714 7532 33748
rect 7566 33714 7582 33748
rect 7516 33679 7582 33714
rect 7516 33645 7532 33679
rect 7566 33645 7582 33679
rect 7516 33610 7582 33645
rect 7516 33576 7532 33610
rect 7566 33576 7582 33610
rect 7516 33541 7582 33576
rect 7516 33507 7532 33541
rect 7566 33507 7582 33541
rect 7516 33472 7582 33507
rect 7516 33438 7532 33472
rect 7566 33438 7582 33472
rect 7516 33403 7582 33438
rect 7516 33369 7532 33403
rect 7566 33369 7582 33403
rect 7516 33334 7582 33369
rect 7516 33300 7532 33334
rect 7566 33300 7582 33334
rect 7516 33265 7582 33300
rect 7516 33231 7532 33265
rect 7566 33231 7582 33265
rect 7516 33196 7582 33231
rect 7516 33162 7532 33196
rect 7566 33162 7582 33196
rect 7516 33127 7582 33162
rect 7516 33093 7532 33127
rect 7566 33093 7582 33127
rect 7516 33058 7582 33093
rect 7516 33024 7532 33058
rect 7566 33024 7582 33058
rect 7516 32989 7582 33024
rect 7516 32955 7532 32989
rect 7566 32955 7582 32989
rect 7516 32920 7582 32955
rect 7516 32886 7532 32920
rect 7566 32886 7582 32920
rect 7516 32851 7582 32886
rect 7516 32817 7532 32851
rect 7566 32817 7582 32851
rect 7516 32782 7582 32817
rect 7516 32748 7532 32782
rect 7566 32748 7582 32782
rect 7516 32713 7582 32748
rect 7516 32679 7532 32713
rect 7566 32679 7582 32713
rect 7516 32663 7582 32679
rect 7516 32591 7582 32607
rect 7516 32557 7532 32591
rect 7566 32557 7582 32591
rect 7516 32522 7582 32557
rect 7516 32488 7532 32522
rect 7566 32488 7582 32522
rect 7516 32453 7582 32488
rect 7516 32419 7532 32453
rect 7566 32419 7582 32453
rect 7516 32384 7582 32419
rect 7516 32350 7532 32384
rect 7566 32350 7582 32384
rect 7516 32315 7582 32350
rect 7516 32281 7532 32315
rect 7566 32281 7582 32315
rect 7516 32246 7582 32281
rect 7516 32212 7532 32246
rect 7566 32212 7582 32246
rect 7516 32177 7582 32212
rect 7516 32143 7532 32177
rect 7566 32143 7582 32177
rect 7516 32108 7582 32143
rect 7516 32074 7532 32108
rect 7566 32074 7582 32108
rect 7516 32039 7582 32074
rect 7516 32005 7532 32039
rect 7566 32005 7582 32039
rect 7516 31970 7582 32005
rect 7516 31936 7532 31970
rect 7566 31936 7582 31970
rect 7516 31901 7582 31936
rect 7516 31867 7532 31901
rect 7566 31867 7582 31901
rect 7516 31832 7582 31867
rect 7516 31798 7532 31832
rect 7566 31798 7582 31832
rect 7516 31763 7582 31798
rect 7516 31729 7532 31763
rect 7566 31729 7582 31763
rect 7516 31693 7582 31729
rect 7516 31659 7532 31693
rect 7566 31659 7582 31693
rect 7516 31623 7582 31659
rect 7516 31589 7532 31623
rect 7566 31589 7582 31623
rect 7516 31553 7582 31589
rect 7516 31519 7532 31553
rect 7566 31519 7582 31553
rect 7516 31483 7582 31519
rect 7516 31449 7532 31483
rect 7566 31449 7582 31483
rect 7516 31413 7582 31449
rect 7516 31379 7532 31413
rect 7566 31379 7582 31413
rect 7516 31343 7582 31379
rect 7516 31309 7532 31343
rect 7566 31309 7582 31343
rect 7516 31273 7582 31309
rect 7516 31239 7532 31273
rect 7566 31239 7582 31273
rect 7516 31203 7582 31239
rect 7516 31169 7532 31203
rect 7566 31169 7582 31203
rect 7516 31133 7582 31169
rect 7516 31099 7532 31133
rect 7566 31099 7582 31133
rect 7516 31063 7582 31099
rect 7516 31029 7532 31063
rect 7566 31029 7582 31063
rect 7516 30993 7582 31029
rect 7516 30959 7532 30993
rect 7566 30959 7582 30993
rect 7516 30923 7582 30959
rect 7516 30889 7532 30923
rect 7566 30889 7582 30923
rect 7516 30853 7582 30889
rect 7516 30819 7532 30853
rect 7566 30819 7582 30853
rect 7516 30783 7582 30819
rect 7516 30749 7532 30783
rect 7566 30749 7582 30783
rect 7516 30713 7582 30749
rect 7516 30679 7532 30713
rect 7566 30679 7582 30713
rect 7516 30643 7582 30679
rect 7516 30609 7532 30643
rect 7566 30609 7582 30643
rect 7516 30573 7582 30609
rect 7516 30539 7532 30573
rect 7566 30539 7582 30573
rect 7516 30503 7582 30539
rect 7516 30469 7532 30503
rect 7566 30469 7582 30503
rect 7516 30433 7582 30469
rect 7516 30399 7532 30433
rect 7566 30399 7582 30433
rect 7516 30383 7582 30399
rect 6788 29888 6922 29904
rect 6788 29854 6804 29888
rect 6838 29854 6872 29888
rect 6906 29854 6922 29888
rect 6788 29838 6922 29854
rect 6978 29888 7112 29904
rect 6978 29854 6994 29888
rect 7028 29854 7062 29888
rect 7096 29854 7112 29888
rect 6978 29838 7112 29854
rect 5838 29566 7438 29582
rect 5838 29532 5854 29566
rect 5888 29532 5924 29566
rect 5958 29532 5994 29566
rect 6028 29532 6064 29566
rect 6098 29532 6134 29566
rect 6168 29532 6204 29566
rect 6238 29532 6274 29566
rect 6308 29532 6344 29566
rect 6378 29532 6414 29566
rect 6448 29532 6484 29566
rect 6518 29532 6554 29566
rect 6588 29532 6624 29566
rect 6658 29532 6694 29566
rect 6728 29532 6764 29566
rect 6798 29532 6834 29566
rect 6868 29532 6904 29566
rect 6938 29532 6974 29566
rect 7008 29532 7043 29566
rect 7077 29532 7112 29566
rect 7146 29532 7181 29566
rect 7215 29532 7250 29566
rect 7284 29532 7319 29566
rect 7353 29532 7388 29566
rect 7422 29532 7438 29566
rect 5838 29516 7438 29532
rect 5864 29194 6664 29210
rect 5864 29160 5880 29194
rect 5914 29160 5954 29194
rect 5988 29160 6028 29194
rect 6062 29160 6102 29194
rect 6136 29160 6176 29194
rect 6210 29160 6249 29194
rect 6283 29160 6322 29194
rect 6356 29160 6395 29194
rect 6429 29160 6468 29194
rect 6502 29160 6541 29194
rect 6575 29160 6614 29194
rect 6648 29160 6664 29194
rect 5864 29144 6664 29160
rect 6934 29194 7068 29210
rect 6934 29160 6950 29194
rect 6984 29160 7018 29194
rect 7052 29160 7068 29194
rect 6934 29144 7068 29160
rect 7300 29194 7434 29210
rect 7300 29160 7316 29194
rect 7350 29160 7384 29194
rect 7418 29160 7434 29194
rect 7300 29144 7434 29160
rect 5864 28822 6664 28838
rect 5864 28788 5880 28822
rect 5914 28788 5954 28822
rect 5988 28788 6028 28822
rect 6062 28788 6102 28822
rect 6136 28788 6176 28822
rect 6210 28788 6249 28822
rect 6283 28788 6322 28822
rect 6356 28788 6395 28822
rect 6429 28788 6468 28822
rect 6502 28788 6541 28822
rect 6575 28788 6614 28822
rect 6648 28788 6664 28822
rect 5864 28772 6664 28788
rect 6934 28822 7068 28838
rect 6934 28788 6950 28822
rect 6984 28788 7018 28822
rect 7052 28788 7068 28822
rect 6934 28772 7068 28788
rect 2757 27094 2827 27110
rect 2757 27060 2773 27094
rect 2807 27060 2827 27094
rect 2757 27044 2827 27060
rect 6050 27094 6120 27110
rect 6050 27060 6070 27094
rect 6104 27060 6120 27094
rect 6050 27044 6120 27060
rect 6447 21604 6581 21620
rect 6447 21570 6463 21604
rect 6497 21570 6531 21604
rect 6565 21570 6581 21604
rect 6447 21554 6581 21570
rect 6637 21604 6771 21620
rect 6637 21570 6653 21604
rect 6687 21570 6721 21604
rect 6755 21570 6771 21604
rect 6637 21554 6771 21570
rect 3840 7265 3906 7281
rect 3840 7231 3856 7265
rect 3890 7231 3906 7265
rect 3840 7196 3906 7231
rect 3840 7162 3856 7196
rect 3890 7162 3906 7196
rect 3840 7127 3906 7162
rect 3840 7093 3856 7127
rect 3890 7093 3906 7127
rect 3840 7058 3906 7093
rect 3840 7024 3856 7058
rect 3890 7024 3906 7058
rect 3840 6989 3906 7024
rect 3840 6955 3856 6989
rect 3890 6955 3906 6989
rect 3840 6920 3906 6955
rect 3840 6886 3856 6920
rect 3890 6886 3906 6920
rect 3840 6851 3906 6886
rect 3840 6817 3856 6851
rect 3890 6817 3906 6851
rect 3840 6781 3906 6817
rect 3840 6747 3856 6781
rect 3890 6747 3906 6781
rect 3840 6711 3906 6747
rect 3840 6677 3856 6711
rect 3890 6677 3906 6711
rect 3840 6641 3906 6677
rect 3840 6607 3856 6641
rect 3890 6607 3906 6641
rect 3840 6571 3906 6607
rect 3840 6537 3856 6571
rect 3890 6537 3906 6571
rect 3840 6501 3906 6537
rect 3840 6467 3856 6501
rect 3890 6467 3906 6501
rect 3840 6431 3906 6467
rect 3840 6397 3856 6431
rect 3890 6397 3906 6431
rect 3840 6361 3906 6397
rect 3840 6327 3856 6361
rect 3890 6327 3906 6361
rect 3840 6291 3906 6327
rect 3840 6257 3856 6291
rect 3890 6257 3906 6291
rect 3840 6221 3906 6257
rect 3840 6187 3856 6221
rect 3890 6187 3906 6221
rect 3840 6151 3906 6187
rect 3840 6117 3856 6151
rect 3890 6117 3906 6151
rect 3840 6081 3906 6117
rect 3840 6047 3856 6081
rect 3890 6047 3906 6081
rect 3840 6011 3906 6047
rect 3840 5977 3856 6011
rect 3890 5977 3906 6011
rect 3840 5941 3906 5977
rect 3840 5907 3856 5941
rect 3890 5907 3906 5941
rect 3840 5871 3906 5907
rect 3840 5837 3856 5871
rect 3890 5837 3906 5871
rect 3840 5801 3906 5837
rect 3840 5767 3856 5801
rect 3890 5767 3906 5801
rect 3840 5731 3906 5767
rect 3840 5697 3856 5731
rect 3890 5697 3906 5731
rect 3840 5681 3906 5697
rect 4570 7265 4636 7281
rect 4570 7231 4586 7265
rect 4620 7231 4636 7265
rect 4570 7196 4636 7231
rect 4570 7162 4586 7196
rect 4620 7162 4636 7196
rect 4570 7127 4636 7162
rect 4570 7093 4586 7127
rect 4620 7093 4636 7127
rect 4570 7058 4636 7093
rect 4570 7024 4586 7058
rect 4620 7024 4636 7058
rect 4570 6989 4636 7024
rect 4570 6955 4586 6989
rect 4620 6955 4636 6989
rect 4570 6920 4636 6955
rect 4570 6886 4586 6920
rect 4620 6886 4636 6920
rect 4570 6851 4636 6886
rect 4570 6817 4586 6851
rect 4620 6817 4636 6851
rect 4570 6781 4636 6817
rect 4570 6747 4586 6781
rect 4620 6747 4636 6781
rect 4570 6711 4636 6747
rect 4570 6677 4586 6711
rect 4620 6677 4636 6711
rect 4570 6641 4636 6677
rect 4570 6607 4586 6641
rect 4620 6607 4636 6641
rect 4570 6571 4636 6607
rect 4570 6537 4586 6571
rect 4620 6537 4636 6571
rect 4570 6501 4636 6537
rect 4570 6467 4586 6501
rect 4620 6467 4636 6501
rect 4570 6431 4636 6467
rect 4570 6397 4586 6431
rect 4620 6397 4636 6431
rect 4570 6361 4636 6397
rect 4570 6327 4586 6361
rect 4620 6327 4636 6361
rect 4570 6291 4636 6327
rect 4570 6257 4586 6291
rect 4620 6257 4636 6291
rect 4570 6221 4636 6257
rect 4570 6187 4586 6221
rect 4620 6187 4636 6221
rect 4570 6151 4636 6187
rect 4570 6117 4586 6151
rect 4620 6117 4636 6151
rect 4570 6081 4636 6117
rect 4570 6047 4586 6081
rect 4620 6047 4636 6081
rect 4570 6011 4636 6047
rect 4570 5977 4586 6011
rect 4620 5977 4636 6011
rect 4570 5941 4636 5977
rect 4570 5907 4586 5941
rect 4620 5907 4636 5941
rect 4570 5871 4636 5907
rect 4570 5837 4586 5871
rect 4620 5837 4636 5871
rect 4570 5801 4636 5837
rect 4570 5767 4586 5801
rect 4620 5767 4636 5801
rect 4570 5731 4636 5767
rect 4570 5697 4586 5731
rect 4620 5697 4636 5731
rect 4570 5681 4636 5697
rect 6084 7108 6150 7124
rect 6084 7074 6100 7108
rect 6134 7074 6150 7108
rect 6084 7025 6150 7074
rect 6084 6991 6100 7025
rect 6134 6991 6150 7025
rect 6084 6942 6150 6991
rect 6084 6908 6100 6942
rect 6134 6908 6150 6942
rect 6084 6858 6150 6908
rect 6084 6824 6100 6858
rect 6134 6824 6150 6858
rect 6084 6774 6150 6824
rect 6084 6740 6100 6774
rect 6134 6740 6150 6774
rect 6084 6724 6150 6740
rect 6084 6536 6150 6552
rect 6084 6502 6100 6536
rect 6134 6502 6150 6536
rect 6084 6463 6150 6502
rect 6084 6429 6100 6463
rect 6134 6429 6150 6463
rect 6084 6390 6150 6429
rect 6084 6356 6100 6390
rect 6134 6356 6150 6390
rect 6084 6317 6150 6356
rect 6084 6283 6100 6317
rect 6134 6283 6150 6317
rect 6084 6244 6150 6283
rect 6084 6210 6100 6244
rect 6134 6210 6150 6244
rect 6084 6171 6150 6210
rect 6084 6137 6100 6171
rect 6134 6137 6150 6171
rect 6084 6098 6150 6137
rect 6084 6064 6100 6098
rect 6134 6064 6150 6098
rect 6084 6024 6150 6064
rect 6084 5990 6100 6024
rect 6134 5990 6150 6024
rect 6084 5950 6150 5990
rect 6084 5916 6100 5950
rect 6134 5916 6150 5950
rect 6084 5876 6150 5916
rect 6084 5842 6100 5876
rect 6134 5842 6150 5876
rect 6084 5802 6150 5842
rect 6084 5768 6100 5802
rect 6134 5768 6150 5802
rect 5670 5742 5804 5758
rect 6084 5752 6150 5768
rect 5670 5708 5686 5742
rect 5720 5708 5754 5742
rect 5788 5708 5804 5742
rect 5670 5692 5804 5708
rect 3039 4773 3607 4789
rect 3039 4739 3055 4773
rect 3089 4739 3127 4773
rect 3161 4739 3199 4773
rect 3233 4739 3271 4773
rect 3305 4739 3343 4773
rect 3377 4739 3415 4773
rect 3449 4739 3486 4773
rect 3520 4739 3557 4773
rect 3591 4739 3607 4773
rect 3039 4723 3607 4739
rect 6320 4660 6386 4676
rect 6320 4626 6336 4660
rect 6370 4626 6386 4660
rect 6320 4589 6386 4626
rect 6320 4555 6336 4589
rect 6370 4555 6386 4589
rect 6320 4518 6386 4555
rect 6320 4484 6336 4518
rect 6370 4484 6386 4518
rect 4267 4443 5867 4459
rect 4267 4409 4283 4443
rect 4317 4409 4353 4443
rect 4387 4409 4423 4443
rect 4457 4409 4493 4443
rect 4527 4409 4563 4443
rect 4597 4409 4633 4443
rect 4667 4409 4703 4443
rect 4737 4409 4773 4443
rect 4807 4409 4843 4443
rect 4877 4409 4913 4443
rect 4947 4409 4983 4443
rect 5017 4409 5053 4443
rect 5087 4409 5123 4443
rect 5157 4409 5193 4443
rect 5227 4409 5263 4443
rect 5297 4409 5333 4443
rect 5367 4409 5403 4443
rect 5437 4409 5472 4443
rect 5506 4409 5541 4443
rect 5575 4409 5610 4443
rect 5644 4409 5679 4443
rect 5713 4409 5748 4443
rect 5782 4409 5817 4443
rect 5851 4409 5867 4443
rect 4267 4393 5867 4409
rect 6320 4446 6386 4484
rect 6320 4412 6336 4446
rect 6370 4412 6386 4446
rect 6320 4374 6386 4412
rect 6320 4340 6336 4374
rect 6370 4340 6386 4374
rect 6320 4302 6386 4340
rect 6320 4268 6336 4302
rect 6370 4268 6386 4302
rect 6320 4230 6386 4268
rect 6320 4196 6336 4230
rect 6370 4196 6386 4230
rect 6320 4158 6386 4196
rect 6320 4124 6336 4158
rect 6370 4124 6386 4158
rect 6320 4086 6386 4124
rect 4211 4049 5867 4065
rect 4211 4015 4227 4049
rect 4261 4015 4297 4049
rect 4331 4015 4367 4049
rect 4401 4015 4437 4049
rect 4471 4015 4506 4049
rect 4540 4015 4575 4049
rect 4609 4015 4644 4049
rect 4678 4015 4713 4049
rect 4747 4015 4782 4049
rect 4816 4015 4851 4049
rect 4885 4015 4920 4049
rect 4954 4015 4989 4049
rect 5023 4015 5058 4049
rect 5092 4015 5127 4049
rect 5161 4015 5196 4049
rect 5230 4015 5265 4049
rect 5299 4015 5334 4049
rect 5368 4015 5403 4049
rect 5437 4015 5472 4049
rect 5506 4015 5541 4049
rect 5575 4015 5610 4049
rect 5644 4015 5679 4049
rect 5713 4015 5748 4049
rect 5782 4015 5817 4049
rect 5851 4015 5867 4049
rect 4211 3999 5867 4015
rect 6320 4052 6336 4086
rect 6370 4052 6386 4086
rect 6320 4014 6386 4052
rect 6320 3980 6336 4014
rect 6370 3980 6386 4014
rect 6320 3942 6386 3980
rect 6320 3908 6336 3942
rect 6370 3908 6386 3942
rect 6320 3870 6386 3908
rect 6320 3836 6336 3870
rect 6370 3836 6386 3870
rect 6320 3820 6386 3836
<< polycont >>
rect 8148 39617 8182 39651
rect 9606 39617 9640 39651
rect 7532 39397 7566 39431
rect 7532 39329 7566 39363
rect 7532 39261 7566 39295
rect 7532 39193 7566 39227
rect 7532 39125 7566 39159
rect 7532 39057 7566 39091
rect 7532 38989 7566 39023
rect 7532 38921 7566 38955
rect 7532 38853 7566 38887
rect 7532 38785 7566 38819
rect 7532 38717 7566 38751
rect 7532 38649 7566 38683
rect 7532 38581 7566 38615
rect 7532 38513 7566 38547
rect 7532 38445 7566 38479
rect 7532 38377 7566 38411
rect 7532 38309 7566 38343
rect 7532 38241 7566 38275
rect 7532 38173 7566 38207
rect 7532 38105 7566 38139
rect 7532 38037 7566 38071
rect 7532 37969 7566 38003
rect 7532 37901 7566 37935
rect 7532 37833 7566 37867
rect 7532 37765 7566 37799
rect 7532 37697 7566 37731
rect 7532 37629 7566 37663
rect 7532 37561 7566 37595
rect 7532 37493 7566 37527
rect 7532 37425 7566 37459
rect 7532 37357 7566 37391
rect 7532 37289 7566 37323
rect 7532 37221 7566 37255
rect 7532 37153 7566 37187
rect 7532 37085 7566 37119
rect 7532 37017 7566 37051
rect 7532 36949 7566 36983
rect 7532 36881 7566 36915
rect 7532 36813 7566 36847
rect 7532 36745 7566 36779
rect 7532 36677 7566 36711
rect 7532 36609 7566 36643
rect 7532 36541 7566 36575
rect 7532 36473 7566 36507
rect 7532 36405 7566 36439
rect 7532 36336 7566 36370
rect 7532 36267 7566 36301
rect 7532 36198 7566 36232
rect 7532 36129 7566 36163
rect 7532 36060 7566 36094
rect 7532 35991 7566 36025
rect 7532 35922 7566 35956
rect 7532 35853 7566 35887
rect 7532 35784 7566 35818
rect 7532 35715 7566 35749
rect 7532 35646 7566 35680
rect 7532 35577 7566 35611
rect 7532 35508 7566 35542
rect 7532 35439 7566 35473
rect 7532 35370 7566 35404
rect 7532 35301 7566 35335
rect 7532 35232 7566 35266
rect 7532 35163 7566 35197
rect 7532 35094 7566 35128
rect 7532 35025 7566 35059
rect 7532 34956 7566 34990
rect 7532 34887 7566 34921
rect 7532 34818 7566 34852
rect 7532 34749 7566 34783
rect 7532 34680 7566 34714
rect 7532 34611 7566 34645
rect 7532 34542 7566 34576
rect 7532 34473 7566 34507
rect 7532 34404 7566 34438
rect 7532 34335 7566 34369
rect 7532 34266 7566 34300
rect 7532 34197 7566 34231
rect 7532 34128 7566 34162
rect 7532 34059 7566 34093
rect 7532 33990 7566 34024
rect 7532 33921 7566 33955
rect 7532 33852 7566 33886
rect 7532 33783 7566 33817
rect 7532 33714 7566 33748
rect 7532 33645 7566 33679
rect 7532 33576 7566 33610
rect 7532 33507 7566 33541
rect 7532 33438 7566 33472
rect 7532 33369 7566 33403
rect 7532 33300 7566 33334
rect 7532 33231 7566 33265
rect 7532 33162 7566 33196
rect 7532 33093 7566 33127
rect 7532 33024 7566 33058
rect 7532 32955 7566 32989
rect 7532 32886 7566 32920
rect 7532 32817 7566 32851
rect 7532 32748 7566 32782
rect 7532 32679 7566 32713
rect 7532 32557 7566 32591
rect 7532 32488 7566 32522
rect 7532 32419 7566 32453
rect 7532 32350 7566 32384
rect 7532 32281 7566 32315
rect 7532 32212 7566 32246
rect 7532 32143 7566 32177
rect 7532 32074 7566 32108
rect 7532 32005 7566 32039
rect 7532 31936 7566 31970
rect 7532 31867 7566 31901
rect 7532 31798 7566 31832
rect 7532 31729 7566 31763
rect 7532 31659 7566 31693
rect 7532 31589 7566 31623
rect 7532 31519 7566 31553
rect 7532 31449 7566 31483
rect 7532 31379 7566 31413
rect 7532 31309 7566 31343
rect 7532 31239 7566 31273
rect 7532 31169 7566 31203
rect 7532 31099 7566 31133
rect 7532 31029 7566 31063
rect 7532 30959 7566 30993
rect 7532 30889 7566 30923
rect 7532 30819 7566 30853
rect 7532 30749 7566 30783
rect 7532 30679 7566 30713
rect 7532 30609 7566 30643
rect 7532 30539 7566 30573
rect 7532 30469 7566 30503
rect 7532 30399 7566 30433
rect 6804 29854 6838 29888
rect 6872 29854 6906 29888
rect 6994 29854 7028 29888
rect 7062 29854 7096 29888
rect 5854 29532 5888 29566
rect 5924 29532 5958 29566
rect 5994 29532 6028 29566
rect 6064 29532 6098 29566
rect 6134 29532 6168 29566
rect 6204 29532 6238 29566
rect 6274 29532 6308 29566
rect 6344 29532 6378 29566
rect 6414 29532 6448 29566
rect 6484 29532 6518 29566
rect 6554 29532 6588 29566
rect 6624 29532 6658 29566
rect 6694 29532 6728 29566
rect 6764 29532 6798 29566
rect 6834 29532 6868 29566
rect 6904 29532 6938 29566
rect 6974 29532 7008 29566
rect 7043 29532 7077 29566
rect 7112 29532 7146 29566
rect 7181 29532 7215 29566
rect 7250 29532 7284 29566
rect 7319 29532 7353 29566
rect 7388 29532 7422 29566
rect 5880 29160 5914 29194
rect 5954 29160 5988 29194
rect 6028 29160 6062 29194
rect 6102 29160 6136 29194
rect 6176 29160 6210 29194
rect 6249 29160 6283 29194
rect 6322 29160 6356 29194
rect 6395 29160 6429 29194
rect 6468 29160 6502 29194
rect 6541 29160 6575 29194
rect 6614 29160 6648 29194
rect 6950 29160 6984 29194
rect 7018 29160 7052 29194
rect 7316 29160 7350 29194
rect 7384 29160 7418 29194
rect 5880 28788 5914 28822
rect 5954 28788 5988 28822
rect 6028 28788 6062 28822
rect 6102 28788 6136 28822
rect 6176 28788 6210 28822
rect 6249 28788 6283 28822
rect 6322 28788 6356 28822
rect 6395 28788 6429 28822
rect 6468 28788 6502 28822
rect 6541 28788 6575 28822
rect 6614 28788 6648 28822
rect 6950 28788 6984 28822
rect 7018 28788 7052 28822
rect 2773 27060 2807 27094
rect 6070 27060 6104 27094
rect 6463 21570 6497 21604
rect 6531 21570 6565 21604
rect 6653 21570 6687 21604
rect 6721 21570 6755 21604
rect 3856 7231 3890 7265
rect 3856 7162 3890 7196
rect 3856 7093 3890 7127
rect 3856 7024 3890 7058
rect 3856 6955 3890 6989
rect 3856 6886 3890 6920
rect 3856 6817 3890 6851
rect 3856 6747 3890 6781
rect 3856 6677 3890 6711
rect 3856 6607 3890 6641
rect 3856 6537 3890 6571
rect 3856 6467 3890 6501
rect 3856 6397 3890 6431
rect 3856 6327 3890 6361
rect 3856 6257 3890 6291
rect 3856 6187 3890 6221
rect 3856 6117 3890 6151
rect 3856 6047 3890 6081
rect 3856 5977 3890 6011
rect 3856 5907 3890 5941
rect 3856 5837 3890 5871
rect 3856 5767 3890 5801
rect 3856 5697 3890 5731
rect 4586 7231 4620 7265
rect 4586 7162 4620 7196
rect 4586 7093 4620 7127
rect 4586 7024 4620 7058
rect 4586 6955 4620 6989
rect 4586 6886 4620 6920
rect 4586 6817 4620 6851
rect 4586 6747 4620 6781
rect 4586 6677 4620 6711
rect 4586 6607 4620 6641
rect 4586 6537 4620 6571
rect 4586 6467 4620 6501
rect 4586 6397 4620 6431
rect 4586 6327 4620 6361
rect 4586 6257 4620 6291
rect 4586 6187 4620 6221
rect 4586 6117 4620 6151
rect 4586 6047 4620 6081
rect 4586 5977 4620 6011
rect 4586 5907 4620 5941
rect 4586 5837 4620 5871
rect 4586 5767 4620 5801
rect 4586 5697 4620 5731
rect 6100 7074 6134 7108
rect 6100 6991 6134 7025
rect 6100 6908 6134 6942
rect 6100 6824 6134 6858
rect 6100 6740 6134 6774
rect 6100 6502 6134 6536
rect 6100 6429 6134 6463
rect 6100 6356 6134 6390
rect 6100 6283 6134 6317
rect 6100 6210 6134 6244
rect 6100 6137 6134 6171
rect 6100 6064 6134 6098
rect 6100 5990 6134 6024
rect 6100 5916 6134 5950
rect 6100 5842 6134 5876
rect 6100 5768 6134 5802
rect 5686 5708 5720 5742
rect 5754 5708 5788 5742
rect 3055 4739 3089 4773
rect 3127 4739 3161 4773
rect 3199 4739 3233 4773
rect 3271 4739 3305 4773
rect 3343 4739 3377 4773
rect 3415 4739 3449 4773
rect 3486 4739 3520 4773
rect 3557 4739 3591 4773
rect 6336 4626 6370 4660
rect 6336 4555 6370 4589
rect 6336 4484 6370 4518
rect 4283 4409 4317 4443
rect 4353 4409 4387 4443
rect 4423 4409 4457 4443
rect 4493 4409 4527 4443
rect 4563 4409 4597 4443
rect 4633 4409 4667 4443
rect 4703 4409 4737 4443
rect 4773 4409 4807 4443
rect 4843 4409 4877 4443
rect 4913 4409 4947 4443
rect 4983 4409 5017 4443
rect 5053 4409 5087 4443
rect 5123 4409 5157 4443
rect 5193 4409 5227 4443
rect 5263 4409 5297 4443
rect 5333 4409 5367 4443
rect 5403 4409 5437 4443
rect 5472 4409 5506 4443
rect 5541 4409 5575 4443
rect 5610 4409 5644 4443
rect 5679 4409 5713 4443
rect 5748 4409 5782 4443
rect 5817 4409 5851 4443
rect 6336 4412 6370 4446
rect 6336 4340 6370 4374
rect 6336 4268 6370 4302
rect 6336 4196 6370 4230
rect 6336 4124 6370 4158
rect 4227 4015 4261 4049
rect 4297 4015 4331 4049
rect 4367 4015 4401 4049
rect 4437 4015 4471 4049
rect 4506 4015 4540 4049
rect 4575 4015 4609 4049
rect 4644 4015 4678 4049
rect 4713 4015 4747 4049
rect 4782 4015 4816 4049
rect 4851 4015 4885 4049
rect 4920 4015 4954 4049
rect 4989 4015 5023 4049
rect 5058 4015 5092 4049
rect 5127 4015 5161 4049
rect 5196 4015 5230 4049
rect 5265 4015 5299 4049
rect 5334 4015 5368 4049
rect 5403 4015 5437 4049
rect 5472 4015 5506 4049
rect 5541 4015 5575 4049
rect 5610 4015 5644 4049
rect 5679 4015 5713 4049
rect 5748 4015 5782 4049
rect 5817 4015 5851 4049
rect 6336 4052 6370 4086
rect 6336 3980 6370 4014
rect 6336 3908 6370 3942
rect 6336 3836 6370 3870
<< locali >>
rect 366 39888 2599 39894
rect 366 39854 445 39888
rect 479 39886 518 39888
rect 552 39886 591 39888
rect 625 39886 664 39888
rect 698 39886 737 39888
rect 771 39886 810 39888
rect 844 39886 884 39888
rect 918 39886 958 39888
rect 992 39886 1032 39888
rect 1066 39886 1106 39888
rect 1140 39886 1216 39888
rect 1250 39886 1290 39888
rect 1324 39886 1364 39888
rect 1398 39886 1438 39888
rect 1472 39886 1512 39888
rect 1546 39886 1587 39888
rect 1621 39886 1662 39888
rect 1696 39886 1737 39888
rect 1771 39886 1812 39888
rect 1846 39886 1887 39888
rect 1921 39886 1962 39888
rect 1996 39886 2037 39888
rect 2071 39886 2112 39888
rect 2146 39886 2187 39888
rect 2221 39886 2262 39888
rect 2296 39886 2337 39888
rect 2371 39886 2412 39888
rect 2446 39886 2487 39888
rect 2521 39886 2599 39888
rect 366 39852 448 39854
rect 482 39852 516 39886
rect 366 39818 516 39852
rect 366 39816 374 39818
rect 476 39816 516 39818
rect 2522 39816 2599 39886
rect 366 39782 372 39816
rect 478 39784 516 39816
rect 478 39782 518 39784
rect 552 39782 591 39784
rect 625 39782 664 39784
rect 698 39782 737 39784
rect 771 39782 810 39784
rect 844 39782 884 39784
rect 918 39782 958 39784
rect 992 39782 1032 39784
rect 1066 39782 1106 39784
rect 1140 39782 1216 39784
rect 1250 39782 1290 39784
rect 1324 39782 1364 39784
rect 1398 39782 1438 39784
rect 1472 39782 1512 39784
rect 1546 39782 1587 39784
rect 1621 39782 1662 39784
rect 1696 39782 1737 39784
rect 1771 39782 1812 39784
rect 1846 39782 1887 39784
rect 1921 39782 1962 39784
rect 1996 39782 2037 39784
rect 2071 39782 2112 39784
rect 2146 39782 2187 39784
rect 2221 39782 2262 39784
rect 2296 39782 2337 39784
rect 2371 39782 2412 39784
rect 2446 39782 2487 39784
rect 366 39743 374 39782
rect 476 39776 2487 39782
rect 476 39743 484 39776
rect 366 39709 372 39743
rect 478 39709 484 39743
rect 366 39670 374 39709
rect 476 39670 484 39709
rect 366 39636 372 39670
rect 478 39636 484 39670
rect 366 39597 374 39636
rect 476 39597 484 39636
rect 366 39563 372 39597
rect 478 39563 484 39597
rect 366 39524 374 39563
rect 476 39524 484 39563
rect 366 39490 372 39524
rect 478 39490 484 39524
rect 366 39451 374 39490
rect 476 39451 484 39490
rect 548 39667 566 39701
rect 600 39667 638 39701
rect 548 39628 672 39667
rect 548 39594 566 39628
rect 600 39594 638 39628
rect 548 39555 672 39594
rect 548 39521 566 39555
rect 600 39521 638 39555
rect 548 39489 672 39521
rect 2344 39679 2382 39713
rect 2310 39640 2416 39679
rect 2344 39606 2382 39640
rect 2310 39567 2416 39606
rect 2344 39533 2382 39567
rect 2310 39490 2416 39533
rect 366 39417 372 39451
rect 478 39417 484 39451
rect 366 39378 374 39417
rect 476 39378 484 39417
rect 366 39344 372 39378
rect 478 39344 484 39378
rect 366 39305 374 39344
rect 476 39305 484 39344
rect 366 39271 372 39305
rect 478 39271 484 39305
rect 366 39232 374 39271
rect 476 39232 484 39271
rect 366 39198 372 39232
rect 478 39198 484 39232
rect 366 39159 374 39198
rect 476 39159 484 39198
rect 366 39125 372 39159
rect 478 39125 484 39159
rect 366 39086 374 39125
rect 476 39086 484 39125
rect 366 39052 372 39086
rect 478 39052 484 39086
rect 366 39013 374 39052
rect 476 39013 484 39052
rect 366 38979 372 39013
rect 478 38979 484 39013
rect 366 38940 374 38979
rect 476 38940 484 38979
rect 366 38906 372 38940
rect 478 38906 484 38940
rect 366 38867 374 38906
rect 476 38867 484 38906
rect 366 38833 372 38867
rect 478 38833 484 38867
rect 366 38794 374 38833
rect 476 38794 484 38833
rect 366 38760 372 38794
rect 478 38760 484 38794
rect 366 38721 374 38760
rect 476 38721 484 38760
rect 366 38687 372 38721
rect 478 38687 484 38721
rect 366 38648 374 38687
rect 476 38648 484 38687
rect 366 38614 372 38648
rect 478 38614 484 38648
rect 366 38575 374 38614
rect 476 38575 484 38614
rect 366 38541 372 38575
rect 478 38541 484 38575
rect 366 38502 374 38541
rect 476 38502 484 38541
rect 366 38468 372 38502
rect 478 38468 484 38502
rect 366 38429 374 38468
rect 476 38429 484 38468
rect 366 38395 372 38429
rect 478 38395 484 38429
rect 366 38356 374 38395
rect 476 38356 484 38395
rect 366 38322 372 38356
rect 478 38322 484 38356
rect 366 38283 374 38322
rect 476 38283 484 38322
rect 366 38249 372 38283
rect 478 38249 484 38283
rect 366 38210 374 38249
rect 476 38210 484 38249
rect 366 38176 372 38210
rect 478 38176 484 38210
rect 366 38137 374 38176
rect 476 38137 484 38176
rect 366 38103 372 38137
rect 478 38103 484 38137
rect 366 38064 374 38103
rect 476 38064 484 38103
rect 366 38030 372 38064
rect 478 38030 484 38064
rect 366 37991 374 38030
rect 476 37991 484 38030
rect 366 37957 372 37991
rect 478 37957 484 37991
rect 366 37918 374 37957
rect 476 37918 484 37957
rect 366 37884 372 37918
rect 478 37884 484 37918
rect 366 37845 374 37884
rect 476 37845 484 37884
rect 366 37811 372 37845
rect 478 37811 484 37845
rect 366 37772 374 37811
rect 476 37772 484 37811
rect 366 37738 372 37772
rect 478 37738 484 37772
rect 366 37699 374 37738
rect 476 37699 484 37738
rect 366 37665 372 37699
rect 478 37665 484 37699
rect 366 37626 374 37665
rect 476 37626 484 37665
rect 366 37592 372 37626
rect 478 37592 484 37626
rect 366 37553 374 37592
rect 476 37553 484 37592
rect 366 37519 372 37553
rect 478 37519 484 37553
rect 366 37480 374 37519
rect 476 37480 484 37519
rect 366 37446 372 37480
rect 478 37446 484 37480
rect 366 37407 374 37446
rect 476 37407 484 37446
rect 366 37373 372 37407
rect 478 37373 484 37407
rect 366 37334 374 37373
rect 476 37334 484 37373
rect 366 436 372 37334
rect 478 436 484 37334
rect 366 398 374 436
rect 476 398 484 436
rect 2481 2918 2487 39776
rect 2593 2918 2599 39816
rect 8002 39889 10828 39895
rect 8002 39855 8040 39889
rect 8074 39886 8116 39889
rect 8150 39886 8192 39889
rect 8226 39886 8268 39889
rect 8302 39886 8345 39889
rect 8379 39886 8422 39889
rect 8456 39886 8499 39889
rect 8533 39886 8576 39889
rect 8610 39886 8653 39889
rect 8687 39886 8730 39889
rect 8764 39886 8840 39889
rect 10458 39886 10497 39889
rect 10531 39886 10570 39889
rect 10604 39886 10643 39889
rect 10677 39886 10716 39889
rect 10750 39886 10828 39889
rect 8002 39817 8066 39855
rect 8002 39783 8040 39817
rect 10752 39817 10828 39886
rect 8074 39783 8116 39784
rect 8150 39783 8192 39784
rect 8226 39783 8268 39784
rect 8302 39783 8345 39784
rect 8379 39783 8422 39784
rect 8456 39783 8499 39784
rect 8533 39783 8576 39784
rect 8610 39783 8653 39784
rect 8687 39783 8730 39784
rect 8764 39783 8840 39784
rect 10458 39783 10497 39784
rect 10531 39783 10570 39784
rect 10604 39783 10643 39784
rect 10677 39783 10716 39784
rect 8002 39777 10716 39783
rect 8002 39750 8036 39777
rect 8034 39708 8036 39716
rect 9746 39750 9792 39777
rect 8000 39682 8036 39708
rect 8000 39670 8002 39682
rect 8034 39636 8036 39648
rect 5370 39614 7536 39620
rect 5364 39580 5398 39614
rect 5436 39580 5468 39614
rect 5510 39580 5538 39614
rect 5584 39580 5608 39614
rect 5658 39580 5678 39614
rect 5732 39580 5748 39614
rect 5806 39580 5818 39614
rect 5880 39580 5888 39614
rect 5954 39580 5958 39614
rect 5992 39580 5994 39614
rect 6062 39580 6068 39614
rect 6132 39580 6142 39614
rect 6202 39580 6216 39614
rect 6272 39580 6290 39614
rect 6342 39580 6364 39614
rect 6412 39580 6438 39614
rect 6482 39580 6512 39614
rect 6552 39580 6586 39614
rect 6622 39580 6657 39614
rect 6694 39580 6726 39614
rect 6768 39580 6795 39614
rect 6842 39580 6864 39614
rect 6916 39580 6933 39614
rect 6990 39580 7002 39614
rect 7064 39580 7071 39614
rect 7138 39580 7140 39614
rect 7174 39580 7178 39614
rect 7243 39580 7251 39614
rect 7312 39580 7324 39614
rect 7381 39580 7397 39614
rect 7450 39580 7470 39614
rect 7504 39580 7536 39614
rect 5370 39574 7536 39580
rect 8000 39614 8036 39636
rect 8000 39598 8002 39614
rect 8034 39564 8036 39580
rect 8000 39546 8036 39564
rect 8000 39526 8002 39546
rect 8146 39679 8184 39713
rect 8112 39651 8218 39679
rect 8112 39640 8148 39651
rect 8146 39617 8148 39640
rect 8182 39640 8218 39651
rect 8182 39617 8184 39640
rect 8146 39606 8184 39617
rect 8112 39567 8218 39606
rect 8146 39533 8184 39567
rect 9598 39679 9636 39713
rect 9564 39651 9670 39679
rect 9564 39640 9606 39651
rect 9640 39640 9670 39651
rect 9598 39617 9606 39640
rect 9598 39606 9636 39617
rect 9564 39567 9670 39606
rect 9598 39533 9636 39567
rect 9746 39711 9752 39750
rect 9786 39711 9792 39750
rect 9746 39682 9792 39711
rect 9746 39639 9752 39682
rect 9786 39639 9792 39682
rect 9746 39614 9792 39639
rect 9746 39567 9752 39614
rect 9786 39567 9792 39614
rect 9746 39546 9792 39567
rect 8034 39492 8036 39512
rect 8000 39478 8036 39492
rect 8000 39454 8002 39478
rect 7532 39431 7566 39447
rect 7532 39363 7566 39397
rect 7532 39295 7566 39322
rect 7532 39227 7566 39250
rect 7532 39159 7566 39178
rect 7532 39091 7566 39106
rect 7532 39023 7566 39034
rect 7532 38955 7566 38962
rect 7532 38887 7566 38890
rect 7532 38852 7566 38853
rect 7532 38780 7566 38785
rect 7532 38708 7566 38717
rect 7532 38636 7566 38649
rect 7532 38564 7566 38581
rect 7532 38492 7566 38513
rect 7532 38420 7566 38445
rect 7532 38348 7566 38377
rect 7532 38276 7566 38309
rect 7532 38207 7566 38241
rect 7532 38139 7566 38170
rect 7532 38071 7566 38098
rect 7532 38003 7566 38026
rect 7532 37935 7566 37954
rect 7532 37867 7566 37882
rect 7532 37799 7566 37810
rect 7532 37731 7566 37738
rect 7532 37663 7566 37666
rect 7532 37628 7566 37629
rect 7532 37556 7566 37561
rect 7532 37484 7566 37493
rect 7532 37412 7566 37425
rect 7532 37340 7566 37357
rect 7532 37267 7566 37289
rect 7532 37194 7566 37221
rect 7532 37121 7566 37153
rect 7532 37051 7566 37085
rect 7532 36983 7566 37014
rect 7532 36915 7566 36941
rect 7532 36847 7566 36868
rect 7532 36779 7566 36795
rect 7532 36711 7566 36722
rect 7532 36643 7566 36649
rect 7532 36575 7566 36576
rect 7532 36537 7566 36541
rect 7532 36464 7566 36473
rect 7532 36391 7566 36405
rect 7532 36318 7566 36336
rect 7532 36245 7566 36267
rect 7532 36172 7566 36198
rect 7532 36099 7566 36129
rect 7532 36026 7566 36060
rect 7532 35956 7566 35991
rect 7532 35887 7566 35919
rect 7532 35818 7566 35846
rect 7532 35749 7566 35773
rect 7532 35680 7566 35700
rect 7532 35611 7566 35627
rect 7532 35542 7566 35554
rect 7532 35473 7566 35481
rect 7532 35404 7566 35408
rect 7532 35369 7566 35370
rect 7532 35296 7566 35301
rect 7532 35223 7566 35232
rect 7532 35150 7566 35163
rect 7532 35077 7566 35094
rect 7532 35004 7566 35025
rect 7532 34931 7566 34956
rect 7532 34858 7566 34887
rect 7532 34785 7566 34818
rect 7532 34714 7566 34749
rect 7532 34645 7566 34678
rect 7532 34576 7566 34605
rect 7532 34507 7566 34532
rect 7532 34438 7566 34459
rect 7532 34369 7566 34386
rect 7532 34300 7566 34313
rect 7532 34231 7566 34240
rect 7532 34162 7566 34167
rect 7532 34093 7566 34094
rect 7532 34055 7566 34059
rect 7532 33982 7566 33990
rect 7532 33909 7566 33921
rect 7532 33836 7566 33852
rect 7532 33763 7566 33783
rect 7532 33690 7566 33714
rect 7532 33617 7566 33645
rect 7532 33544 7566 33576
rect 7532 33472 7566 33507
rect 7532 33403 7566 33437
rect 7532 33334 7566 33364
rect 7532 33265 7566 33291
rect 7532 33196 7566 33218
rect 7532 33127 7566 33145
rect 7532 33058 7566 33072
rect 7532 32989 7566 32999
rect 7532 32920 7566 32926
rect 7532 32851 7566 32853
rect 7532 32814 7566 32817
rect 7532 32741 7566 32748
rect 7532 32663 7566 32679
rect 8034 39420 8036 39444
rect 8000 39410 8036 39420
rect 8000 39382 8002 39410
rect 8034 39348 8036 39376
rect 8000 39342 8036 39348
rect 8000 39310 8002 39342
rect 8034 39276 8036 39308
rect 8000 39274 8036 39276
rect 8000 39240 8002 39274
rect 8000 39238 8036 39240
rect 8034 39206 8036 39238
rect 8000 39172 8002 39204
rect 8000 39166 8036 39172
rect 8034 39138 8036 39166
rect 8000 39104 8002 39132
rect 8000 39094 8036 39104
rect 8034 39070 8036 39094
rect 8000 39036 8002 39060
rect 8000 39022 8036 39036
rect 8034 39002 8036 39022
rect 8000 38968 8002 38988
rect 8000 38950 8036 38968
rect 8034 38934 8036 38950
rect 8000 38900 8002 38916
rect 8000 38878 8036 38900
rect 8034 38866 8036 38878
rect 8000 38832 8002 38844
rect 8000 38806 8036 38832
rect 8034 38798 8036 38806
rect 8000 38764 8002 38772
rect 8000 38734 8036 38764
rect 8034 38730 8036 38734
rect 8000 38696 8002 38700
rect 8000 38662 8036 38696
rect 8000 38594 8036 38628
rect 8000 38590 8002 38594
rect 8034 38556 8036 38560
rect 8000 38526 8036 38556
rect 8000 38518 8002 38526
rect 8034 38484 8036 38492
rect 8000 38458 8036 38484
rect 8000 38446 8002 38458
rect 8034 38412 8036 38424
rect 8000 38390 8036 38412
rect 8000 38374 8002 38390
rect 8034 38340 8036 38356
rect 8000 38322 8036 38340
rect 8000 38302 8002 38322
rect 8034 38268 8036 38288
rect 8000 38254 8036 38268
rect 8000 38230 8002 38254
rect 8034 38196 8036 38220
rect 8000 38186 8036 38196
rect 8000 38158 8002 38186
rect 8034 38124 8036 38152
rect 8000 38118 8036 38124
rect 8000 38086 8002 38118
rect 8034 38052 8036 38084
rect 8000 38050 8036 38052
rect 8000 38016 8002 38050
rect 8000 38014 8036 38016
rect 8034 37982 8036 38014
rect 8000 37948 8002 37980
rect 8000 37942 8036 37948
rect 8034 37914 8036 37942
rect 8000 37880 8002 37908
rect 8000 37870 8036 37880
rect 8034 37846 8036 37870
rect 8000 37812 8002 37836
rect 8000 37798 8036 37812
rect 8034 37778 8036 37798
rect 8000 37744 8002 37764
rect 8000 37726 8036 37744
rect 8034 37710 8036 37726
rect 8000 37676 8002 37692
rect 8000 37654 8036 37676
rect 8034 37642 8036 37654
rect 8000 37608 8002 37620
rect 8000 37582 8036 37608
rect 8034 37574 8036 37582
rect 8000 37540 8002 37548
rect 8000 37510 8036 37540
rect 8034 37506 8036 37510
rect 8000 37472 8002 37476
rect 8000 37438 8036 37472
rect 8000 37370 8036 37404
rect 8000 37366 8002 37370
rect 8034 37332 8036 37336
rect 8000 37302 8036 37332
rect 8000 37294 8002 37302
rect 8034 37260 8036 37268
rect 8000 37234 8036 37260
rect 8000 37222 8002 37234
rect 8034 37188 8036 37200
rect 8000 37166 8036 37188
rect 8000 37150 8002 37166
rect 8034 37116 8036 37132
rect 8000 37098 8036 37116
rect 8000 37078 8002 37098
rect 8034 37044 8036 37064
rect 8000 37030 8036 37044
rect 8000 37006 8002 37030
rect 8034 36972 8036 36996
rect 8000 36962 8036 36972
rect 8000 36934 8002 36962
rect 8034 36900 8036 36928
rect 8000 36894 8036 36900
rect 8000 36862 8002 36894
rect 8034 36828 8036 36860
rect 8000 36826 8036 36828
rect 8000 36792 8002 36826
rect 8000 36790 8036 36792
rect 8034 36758 8036 36790
rect 8000 36724 8002 36756
rect 8000 36718 8036 36724
rect 8034 36690 8036 36718
rect 8000 36656 8002 36684
rect 8000 36646 8036 36656
rect 8034 36622 8036 36646
rect 8000 36588 8002 36612
rect 8000 36574 8036 36588
rect 8034 36554 8036 36574
rect 8000 36520 8002 36540
rect 8000 36502 8036 36520
rect 8034 36486 8036 36502
rect 8000 36452 8002 36468
rect 8000 36430 8036 36452
rect 8034 36418 8036 36430
rect 8000 36384 8002 36396
rect 8000 36358 8036 36384
rect 8034 36350 8036 36358
rect 8000 36316 8002 36324
rect 8000 36286 8036 36316
rect 8034 36282 8036 36286
rect 8000 36248 8002 36252
rect 8000 36214 8036 36248
rect 8000 36146 8036 36180
rect 8000 36142 8002 36146
rect 8034 36108 8036 36112
rect 8000 36078 8036 36108
rect 8000 36070 8002 36078
rect 8034 36036 8036 36044
rect 8000 36010 8036 36036
rect 8000 35998 8002 36010
rect 8034 35964 8036 35976
rect 8000 35942 8036 35964
rect 8000 35926 8002 35942
rect 8034 35892 8036 35908
rect 8000 35874 8036 35892
rect 8000 35854 8002 35874
rect 8034 35820 8036 35840
rect 8000 35806 8036 35820
rect 8000 35782 8002 35806
rect 8034 35748 8036 35772
rect 8000 35738 8036 35748
rect 8000 35710 8002 35738
rect 8034 35676 8036 35704
rect 8000 35670 8036 35676
rect 8000 35638 8002 35670
rect 8034 35604 8036 35636
rect 8000 35602 8036 35604
rect 8000 35568 8002 35602
rect 8000 35566 8036 35568
rect 8034 35534 8036 35566
rect 8000 35500 8002 35532
rect 8000 35494 8036 35500
rect 8034 35466 8036 35494
rect 8000 35432 8002 35460
rect 8000 35422 8036 35432
rect 8034 35398 8036 35422
rect 8000 35364 8002 35388
rect 8000 35350 8036 35364
rect 8034 35330 8036 35350
rect 8000 35296 8002 35316
rect 8000 35278 8036 35296
rect 8034 35262 8036 35278
rect 8000 35228 8002 35244
rect 8000 35206 8036 35228
rect 8034 35194 8036 35206
rect 8000 35160 8002 35172
rect 8000 35134 8036 35160
rect 8034 35126 8036 35134
rect 8000 35092 8002 35100
rect 8000 35062 8036 35092
rect 8034 35058 8036 35062
rect 8000 35024 8002 35028
rect 8000 34990 8036 35024
rect 8000 34922 8036 34956
rect 8000 34918 8002 34922
rect 8034 34884 8036 34888
rect 8000 34854 8036 34884
rect 8000 34846 8002 34854
rect 8034 34812 8036 34820
rect 8000 34786 8036 34812
rect 8000 34774 8002 34786
rect 8034 34740 8036 34752
rect 8000 34718 8036 34740
rect 8000 34702 8002 34718
rect 8034 34668 8036 34684
rect 8000 34650 8036 34668
rect 8000 34630 8002 34650
rect 8034 34596 8036 34616
rect 8000 34582 8036 34596
rect 8000 34558 8002 34582
rect 8034 34524 8036 34548
rect 8000 34514 8036 34524
rect 8000 34486 8002 34514
rect 8034 34452 8036 34480
rect 8000 34446 8036 34452
rect 8000 34414 8002 34446
rect 8034 34380 8036 34412
rect 8000 34378 8036 34380
rect 8000 34344 8002 34378
rect 8000 34342 8036 34344
rect 8034 34310 8036 34342
rect 8000 34276 8002 34308
rect 8000 34270 8036 34276
rect 8034 34242 8036 34270
rect 8000 34208 8002 34236
rect 8000 34198 8036 34208
rect 8034 34174 8036 34198
rect 8000 34140 8002 34164
rect 8000 34126 8036 34140
rect 8034 34106 8036 34126
rect 8000 34072 8002 34092
rect 8000 34054 8036 34072
rect 8034 34038 8036 34054
rect 8000 34004 8002 34020
rect 8000 33982 8036 34004
rect 8034 33970 8036 33982
rect 8000 33936 8002 33948
rect 8000 33910 8036 33936
rect 8034 33902 8036 33910
rect 8000 33868 8002 33876
rect 8000 33838 8036 33868
rect 8034 33834 8036 33838
rect 8000 33800 8002 33804
rect 8000 33766 8036 33800
rect 8000 33698 8036 33732
rect 8000 33694 8002 33698
rect 8034 33660 8036 33664
rect 8000 33630 8036 33660
rect 8000 33622 8002 33630
rect 8034 33588 8036 33596
rect 8000 33562 8036 33588
rect 8000 33550 8002 33562
rect 8034 33516 8036 33528
rect 8000 33494 8036 33516
rect 8000 33478 8002 33494
rect 8034 33444 8036 33460
rect 8000 33426 8036 33444
rect 8000 33406 8002 33426
rect 8034 33372 8036 33392
rect 8000 33358 8036 33372
rect 8000 33334 8002 33358
rect 8034 33300 8036 33324
rect 8000 33290 8036 33300
rect 8000 33262 8002 33290
rect 8034 33228 8036 33256
rect 8000 33222 8036 33228
rect 8000 33190 8002 33222
rect 8034 33156 8036 33188
rect 8000 33154 8036 33156
rect 8000 33120 8002 33154
rect 8000 33118 8036 33120
rect 8034 33086 8036 33118
rect 8000 33052 8002 33084
rect 8000 33046 8036 33052
rect 8034 33018 8036 33046
rect 8000 32984 8002 33012
rect 8000 32974 8036 32984
rect 8034 32950 8036 32974
rect 8000 32916 8002 32940
rect 8000 32902 8036 32916
rect 8034 32882 8036 32902
rect 8000 32848 8002 32868
rect 8000 32830 8036 32848
rect 8034 32814 8036 32830
rect 8000 32780 8002 32796
rect 8000 32758 8036 32780
rect 8034 32746 8036 32758
rect 8000 32712 8002 32724
rect 8000 32686 8036 32712
rect 8034 32678 8036 32686
rect 8000 32644 8002 32652
rect 8000 32614 8036 32644
rect 8034 32610 8036 32614
rect 7532 32591 7566 32607
rect 7532 32539 7566 32557
rect 7532 32467 7566 32488
rect 7532 32395 7566 32419
rect 7532 32323 7566 32350
rect 7532 32251 7566 32281
rect 7532 32179 7566 32212
rect 7532 32108 7566 32143
rect 7532 32039 7566 32073
rect 7532 31970 7566 32001
rect 7532 31901 7566 31929
rect 7532 31832 7566 31857
rect 7532 31763 7566 31785
rect 7532 31693 7566 31713
rect 7532 31623 7566 31641
rect 7532 31553 7566 31569
rect 7532 31483 7566 31497
rect 7532 31413 7566 31425
rect 7532 31343 7566 31353
rect 7532 31273 7566 31281
rect 7532 31203 7566 31209
rect 7532 31133 7566 31137
rect 7532 31063 7566 31065
rect 7532 31026 7566 31029
rect 7532 30953 7566 30959
rect 7532 30880 7566 30889
rect 7532 30807 7566 30819
rect 7532 30734 7566 30749
rect 7532 30661 7566 30679
rect 7532 30588 7566 30609
rect 7532 30515 7566 30539
rect 7532 30442 7566 30469
rect 7532 30383 7566 30399
rect 8000 32576 8002 32580
rect 8000 32542 8036 32576
rect 8000 32474 8036 32508
rect 8000 32470 8002 32474
rect 8034 32436 8036 32440
rect 8000 32406 8036 32436
rect 8000 32398 8002 32406
rect 8034 32364 8036 32372
rect 8000 32338 8036 32364
rect 8000 32326 8002 32338
rect 8034 32292 8036 32304
rect 8000 32270 8036 32292
rect 8000 32254 8002 32270
rect 8034 32220 8036 32236
rect 8000 32202 8036 32220
rect 8000 32182 8002 32202
rect 8034 32148 8036 32168
rect 8000 32134 8036 32148
rect 8000 32110 8002 32134
rect 8034 32076 8036 32100
rect 8000 32066 8036 32076
rect 8000 32038 8002 32066
rect 8034 32004 8036 32032
rect 8000 31998 8036 32004
rect 8000 31966 8002 31998
rect 8034 31932 8036 31964
rect 8000 31930 8036 31932
rect 8000 31896 8002 31930
rect 8000 31894 8036 31896
rect 8034 31862 8036 31894
rect 8000 31828 8002 31860
rect 8000 31822 8036 31828
rect 8034 31794 8036 31822
rect 8000 31760 8002 31788
rect 8000 31750 8036 31760
rect 8034 31726 8036 31750
rect 8000 31692 8002 31716
rect 8000 31678 8036 31692
rect 8034 31658 8036 31678
rect 8000 31624 8002 31644
rect 8000 31606 8036 31624
rect 8034 31590 8036 31606
rect 8000 31556 8002 31572
rect 8000 31534 8036 31556
rect 8034 31522 8036 31534
rect 8000 31488 8002 31500
rect 8000 31462 8036 31488
rect 8034 31454 8036 31462
rect 8000 31420 8002 31428
rect 8000 31390 8036 31420
rect 8034 31386 8036 31390
rect 8000 31352 8002 31356
rect 8000 31318 8036 31352
rect 8000 31250 8036 31284
rect 8000 31246 8002 31250
rect 8034 31212 8036 31216
rect 8000 31182 8036 31212
rect 8000 31174 8002 31182
rect 8034 31140 8036 31148
rect 8000 31114 8036 31140
rect 8000 31102 8002 31114
rect 8034 31068 8036 31080
rect 8000 31046 8036 31068
rect 8000 31030 8002 31046
rect 8034 30996 8036 31012
rect 8000 30978 8036 30996
rect 8000 30958 8002 30978
rect 8034 30924 8036 30944
rect 8000 30910 8036 30924
rect 8000 30886 8002 30910
rect 8034 30852 8036 30876
rect 8000 30842 8036 30852
rect 8000 30814 8002 30842
rect 8034 30780 8036 30808
rect 8000 30774 8036 30780
rect 8000 30742 8002 30774
rect 8034 30708 8036 30740
rect 8000 30706 8036 30708
rect 8000 30672 8002 30706
rect 8000 30670 8036 30672
rect 8034 30638 8036 30670
rect 8000 30604 8002 30636
rect 8000 30598 8036 30604
rect 8034 30570 8036 30598
rect 8000 30536 8002 30564
rect 8000 30526 8036 30536
rect 8034 30502 8036 30526
rect 8000 30468 8002 30492
rect 8000 30454 8036 30468
rect 8034 30434 8036 30454
rect 8000 30400 8002 30420
rect 8000 30382 8036 30400
rect 8034 30366 8036 30382
rect 8000 30332 8002 30348
rect 8000 30310 8036 30332
rect 8034 30298 8036 30310
rect 8000 30264 8002 30276
rect 8000 30238 8036 30264
rect 8034 30230 8036 30238
rect 8000 30196 8002 30204
rect 8000 30166 8036 30196
rect 8034 30162 8036 30166
rect 8000 30128 8002 30132
rect 8000 30094 8036 30128
rect 8000 30026 8036 30060
rect 8000 30022 8002 30026
rect 8034 29988 8036 29992
rect 8000 29958 8036 29988
rect 8000 29950 8002 29958
rect 8034 29916 8036 29924
rect 8000 29890 8036 29916
rect 6838 29854 6853 29888
rect 6906 29854 6922 29888
rect 6978 29854 6994 29888
rect 7047 29854 7062 29888
rect 8000 29878 8002 29890
rect 8034 29844 8036 29856
rect 8000 29822 8036 29844
rect 8000 29806 8002 29822
rect 8034 29772 8036 29788
rect 8000 29754 8036 29772
rect 8000 29734 8002 29754
rect 8034 29700 8036 29720
rect 8000 29686 8036 29700
rect 8000 29662 8002 29686
rect 8034 29628 8036 29652
rect 8000 29618 8036 29628
rect 8000 29590 8002 29618
rect 5838 29565 5854 29566
rect 5888 29565 5924 29566
rect 5838 29532 5850 29565
rect 5888 29532 5923 29565
rect 5958 29532 5994 29566
rect 6028 29565 6064 29566
rect 6098 29565 6134 29566
rect 6168 29565 6204 29566
rect 6238 29565 6274 29566
rect 6308 29565 6344 29566
rect 6378 29565 6414 29566
rect 6448 29565 6484 29566
rect 6518 29565 6554 29566
rect 6588 29565 6624 29566
rect 6658 29565 6694 29566
rect 6728 29565 6764 29566
rect 6798 29565 6834 29566
rect 6868 29565 6904 29566
rect 6030 29532 6064 29565
rect 6103 29532 6134 29565
rect 6176 29532 6204 29565
rect 6249 29532 6274 29565
rect 6322 29532 6344 29565
rect 6395 29532 6414 29565
rect 6468 29532 6484 29565
rect 6541 29532 6554 29565
rect 6613 29532 6624 29565
rect 6685 29532 6694 29565
rect 6757 29532 6764 29565
rect 6829 29532 6834 29565
rect 6901 29532 6904 29565
rect 6938 29565 6974 29566
rect 6938 29532 6939 29565
rect 5884 29531 5923 29532
rect 5957 29531 5996 29532
rect 6030 29531 6069 29532
rect 6103 29531 6142 29532
rect 6176 29531 6215 29532
rect 6249 29531 6288 29532
rect 6322 29531 6361 29532
rect 6395 29531 6434 29532
rect 6468 29531 6507 29532
rect 6541 29531 6579 29532
rect 6613 29531 6651 29532
rect 6685 29531 6723 29532
rect 6757 29531 6795 29532
rect 6829 29531 6867 29532
rect 6901 29531 6939 29532
rect 6973 29532 6974 29565
rect 7008 29565 7043 29566
rect 7077 29565 7112 29566
rect 7146 29565 7181 29566
rect 7215 29565 7250 29566
rect 7284 29565 7319 29566
rect 7353 29565 7388 29566
rect 7422 29565 7438 29566
rect 7008 29532 7011 29565
rect 7077 29532 7083 29565
rect 7146 29532 7155 29565
rect 7215 29532 7227 29565
rect 7284 29532 7299 29565
rect 7353 29532 7371 29565
rect 7422 29532 7443 29565
rect 6973 29531 7011 29532
rect 7045 29531 7083 29532
rect 7117 29531 7155 29532
rect 7189 29531 7227 29532
rect 7261 29531 7299 29532
rect 7333 29531 7371 29532
rect 7405 29531 7443 29532
rect 8034 29556 8036 29584
rect 8000 29550 8036 29556
rect 8000 29518 8002 29550
rect 8034 29484 8036 29516
rect 8000 29482 8036 29484
rect 8000 29448 8002 29482
rect 8000 29446 8036 29448
rect 8034 29414 8036 29446
rect 8000 29380 8002 29412
rect 8000 29374 8036 29380
rect 8034 29346 8036 29374
rect 8000 29312 8002 29340
rect 8000 29302 8036 29312
rect 8034 29278 8036 29302
rect 8000 29244 8002 29268
rect 8000 29230 8036 29244
rect 8034 29210 8036 29230
rect 5864 29160 5880 29194
rect 5914 29160 5939 29194
rect 5988 29160 6020 29194
rect 6062 29160 6101 29194
rect 6136 29160 6176 29194
rect 6216 29160 6249 29194
rect 6297 29160 6322 29194
rect 6378 29160 6395 29194
rect 6459 29160 6468 29194
rect 6502 29160 6505 29194
rect 6539 29160 6541 29194
rect 6575 29160 6585 29194
rect 6648 29160 6664 29194
rect 6934 29160 6946 29194
rect 6984 29160 7018 29194
rect 7052 29160 7068 29194
rect 7300 29160 7314 29194
rect 7350 29160 7384 29194
rect 7420 29160 7434 29194
rect 8000 29176 8002 29196
rect 8000 29158 8036 29176
rect 8034 29142 8036 29158
rect 8000 29108 8002 29124
rect 8000 29086 8036 29108
rect 8034 29074 8036 29086
rect 8000 29040 8002 29052
rect 8000 29014 8036 29040
rect 8034 29006 8036 29014
rect 8000 28972 8002 28980
rect 8000 28942 8036 28972
rect 8034 28938 8036 28942
rect 8000 28904 8002 28908
rect 8000 28870 8036 28904
rect 5864 28788 5880 28822
rect 5914 28788 5939 28822
rect 5988 28788 6020 28822
rect 6062 28788 6101 28822
rect 6136 28788 6176 28822
rect 6216 28788 6249 28822
rect 6297 28788 6322 28822
rect 6378 28788 6395 28822
rect 6459 28788 6468 28822
rect 6502 28788 6505 28822
rect 6539 28788 6541 28822
rect 6575 28788 6585 28822
rect 6648 28788 6664 28822
rect 6934 28788 6946 28822
rect 6984 28788 7018 28822
rect 7052 28788 7068 28822
rect 8000 28802 8036 28836
rect 8000 28798 8002 28802
rect 8034 28764 8036 28768
rect 8000 28734 8036 28764
rect 8000 28726 8002 28734
rect 8034 28692 8036 28700
rect 8000 28666 8036 28692
rect 8000 28654 8002 28666
rect 8034 28620 8036 28632
rect 8000 28598 8036 28620
rect 8000 28582 8002 28598
rect 8034 28548 8036 28564
rect 8000 28530 8036 28548
rect 8000 28510 8002 28530
rect 8034 28476 8036 28496
rect 8000 28462 8036 28476
rect 8000 28438 8002 28462
rect 5849 28390 5867 28424
rect 5907 28390 5943 28424
rect 5978 28390 6015 28424
rect 6053 28390 6086 28424
rect 6129 28390 6157 28424
rect 6205 28390 6228 28424
rect 6280 28390 6299 28424
rect 6355 28390 6370 28424
rect 6430 28390 6441 28424
rect 6505 28390 6512 28424
rect 6580 28390 6583 28424
rect 6617 28390 6621 28424
rect 6688 28390 6696 28424
rect 6759 28390 6771 28424
rect 6830 28390 6846 28424
rect 6901 28390 6921 28424
rect 6971 28390 6996 28424
rect 7041 28390 7071 28424
rect 7111 28390 7146 28424
rect 7181 28390 7217 28424
rect 7255 28390 7287 28424
rect 7330 28390 7357 28424
rect 7405 28390 7415 28424
rect 8034 28404 8036 28428
rect 8000 28394 8036 28404
rect 8000 28366 8002 28394
rect 8034 28332 8036 28360
rect 8000 28326 8036 28332
rect 8000 28294 8002 28326
rect 8034 28260 8036 28292
rect 8000 28258 8036 28260
rect 8000 28224 8002 28258
rect 8000 28222 8036 28224
rect 8034 28190 8036 28222
rect 8000 28156 8002 28188
rect 8000 28150 8036 28156
rect 8034 28122 8036 28150
rect 8000 28088 8002 28116
rect 8000 28078 8036 28088
rect 8034 28054 8036 28078
rect 8000 28020 8002 28044
rect 8000 28006 8036 28020
rect 8034 27986 8036 28006
rect 8000 27952 8002 27972
rect 8000 27934 8036 27952
rect 8034 27918 8036 27934
rect 8000 27884 8002 27900
rect 8000 27862 8036 27884
rect 8034 27850 8036 27862
rect 8000 27816 8002 27828
rect 8000 27790 8036 27816
rect 8034 27782 8036 27790
rect 8000 27748 8002 27756
rect 8000 27718 8036 27748
rect 8034 27714 8036 27718
rect 8000 27680 8002 27684
rect 8000 27646 8036 27680
rect 8000 27578 8036 27612
rect 8000 27574 8002 27578
rect 8034 27540 8036 27544
rect 8000 27510 8036 27540
rect 8000 27502 8002 27510
rect 8034 27468 8036 27476
rect 8000 27442 8036 27468
rect 8000 27430 8002 27442
rect 8034 27396 8036 27408
rect 8000 27374 8036 27396
rect 8000 27358 8002 27374
rect 8034 27324 8036 27340
rect 8000 27306 8036 27324
rect 8000 27286 8002 27306
rect 8034 27252 8036 27272
rect 8000 27238 8036 27252
rect 8000 27214 8002 27238
rect 8034 27180 8036 27204
rect 8000 27170 8036 27180
rect 8000 27142 8002 27170
rect 2757 27094 2825 27126
rect 2757 27060 2773 27094
rect 2807 27092 2825 27094
rect 2859 27092 2875 27126
rect 2807 27060 2875 27092
rect 2757 27054 2875 27060
rect 2757 27020 2825 27054
rect 2859 27020 2875 27054
rect 5917 27094 6120 27111
rect 5917 27088 6070 27094
rect 6104 27088 6120 27094
rect 5917 27054 5929 27088
rect 5963 27060 6070 27088
rect 5963 27054 6071 27060
rect 6105 27054 6120 27088
rect 5917 27037 6120 27054
rect 5917 27032 6117 27037
rect 8034 27108 8036 27136
rect 8000 27102 8036 27108
rect 8000 27070 8002 27102
rect 8034 27036 8036 27068
rect 8000 27034 8036 27036
rect 8000 27000 8002 27034
rect 8000 26998 8036 27000
rect 8034 26966 8036 26998
rect 8000 26932 8002 26964
rect 8000 26926 8036 26932
rect 8034 26898 8036 26926
rect 8000 26864 8002 26892
rect 8000 26854 8036 26864
rect 8034 26830 8036 26854
rect 8000 26796 8002 26820
rect 8000 26782 8036 26796
rect 8034 26762 8036 26782
rect 8000 26728 8002 26748
rect 8000 26710 8036 26728
rect 8034 26694 8036 26710
rect 8000 26660 8002 26676
rect 8000 26638 8036 26660
rect 8034 26626 8036 26638
rect 8000 26592 8002 26604
rect 8000 26566 8036 26592
rect 8034 26558 8036 26566
rect 8000 26524 8002 26532
rect 8000 26494 8036 26524
rect 8034 26490 8036 26494
rect 8000 26456 8002 26460
rect 8000 26422 8036 26456
rect 8000 26354 8036 26388
rect 8000 26350 8002 26354
rect 8034 26316 8036 26320
rect 8000 26286 8036 26316
rect 8000 26278 8002 26286
rect 8034 26244 8036 26252
rect 8000 26218 8036 26244
rect 8000 26206 8002 26218
rect 8034 26172 8036 26184
rect 8000 26150 8036 26172
rect 8000 26134 8002 26150
rect 8034 26100 8036 26116
rect 8000 26082 8036 26100
rect 8000 26062 8002 26082
rect 8034 26028 8036 26048
rect 8000 26014 8036 26028
rect 8000 25990 8002 26014
rect 8034 25956 8036 25980
rect 8000 25946 8036 25956
rect 8000 25918 8002 25946
rect 8034 25884 8036 25912
rect 8000 25878 8036 25884
rect 8000 25846 8002 25878
rect 8034 25812 8036 25844
rect 8000 25810 8036 25812
rect 8000 25776 8002 25810
rect 8000 25774 8036 25776
rect 8034 25742 8036 25774
rect 8000 25708 8002 25740
rect 8000 25702 8036 25708
rect 8034 25674 8036 25702
rect 8000 25640 8002 25668
rect 8000 25630 8036 25640
rect 8034 25606 8036 25630
rect 8000 25572 8002 25596
rect 8000 25558 8036 25572
rect 8034 25538 8036 25558
rect 8000 25504 8002 25524
rect 8000 25486 8036 25504
rect 8034 25470 8036 25486
rect 8000 25436 8002 25452
rect 8000 25414 8036 25436
rect 8034 25402 8036 25414
rect 8000 25368 8002 25380
rect 8000 25342 8036 25368
rect 8034 25334 8036 25342
rect 8000 25300 8002 25308
rect 8000 25270 8036 25300
rect 8034 25266 8036 25270
rect 8000 25232 8002 25236
rect 8000 25198 8036 25232
rect 8000 25130 8036 25164
rect 8000 25126 8002 25130
rect 8034 25092 8036 25096
rect 8000 25062 8036 25092
rect 8000 25054 8002 25062
rect 8034 25020 8036 25028
rect 8000 24994 8036 25020
rect 8000 24982 8002 24994
rect 8034 24948 8036 24960
rect 8000 24926 8036 24948
rect 8000 24910 8002 24926
rect 8034 24876 8036 24892
rect 8000 24858 8036 24876
rect 8000 24838 8002 24858
rect 8034 24804 8036 24824
rect 8000 24790 8036 24804
rect 8000 24766 8002 24790
rect 8034 24732 8036 24756
rect 8000 24722 8036 24732
rect 8000 24694 8002 24722
rect 8034 24660 8036 24688
rect 8000 24654 8036 24660
rect 8000 24622 8002 24654
rect 8034 24588 8036 24620
rect 8000 24586 8036 24588
rect 8000 24552 8002 24586
rect 8000 24550 8036 24552
rect 8034 24518 8036 24550
rect 8000 24484 8002 24516
rect 8000 24478 8036 24484
rect 8034 24450 8036 24478
rect 8000 24416 8002 24444
rect 8000 24406 8036 24416
rect 8034 24382 8036 24406
rect 8000 24348 8002 24372
rect 8000 24334 8036 24348
rect 8034 24314 8036 24334
rect 8000 24280 8002 24300
rect 8000 24262 8036 24280
rect 8034 24246 8036 24262
rect 8000 24212 8002 24228
rect 8000 24190 8036 24212
rect 8034 24178 8036 24190
rect 8000 24144 8002 24156
rect 8000 24118 8036 24144
rect 8034 24110 8036 24118
rect 8000 24076 8002 24084
rect 8000 24046 8036 24076
rect 8034 24042 8036 24046
rect 8000 24008 8002 24012
rect 8000 23974 8036 24008
rect 8000 23906 8036 23940
rect 8000 23902 8002 23906
rect 8034 23868 8036 23872
rect 8000 23838 8036 23868
rect 8000 23830 8002 23838
rect 8034 23796 8036 23804
rect 8000 23770 8036 23796
rect 8000 23758 8002 23770
rect 8034 23724 8036 23736
rect 8000 23702 8036 23724
rect 8000 23686 8002 23702
rect 8034 23652 8036 23668
rect 8000 23634 8036 23652
rect 8000 23614 8002 23634
rect 8034 23580 8036 23600
rect 8000 23566 8036 23580
rect 8000 23542 8002 23566
rect 8034 23508 8036 23532
rect 8000 23498 8036 23508
rect 8000 23470 8002 23498
rect 8034 23436 8036 23464
rect 8000 23430 8036 23436
rect 8000 23398 8002 23430
rect 8034 23364 8036 23396
rect 8000 23362 8036 23364
rect 8000 23328 8002 23362
rect 8000 23326 8036 23328
rect 8034 23294 8036 23326
rect 8000 23260 8002 23292
rect 8000 23254 8036 23260
rect 8034 23226 8036 23254
rect 8000 23192 8002 23220
rect 8000 23182 8036 23192
rect 8034 23158 8036 23182
rect 8000 23124 8002 23148
rect 8000 23110 8036 23124
rect 8034 23090 8036 23110
rect 8000 23056 8002 23076
rect 8000 23038 8036 23056
rect 8034 23022 8036 23038
rect 8000 22988 8002 23004
rect 8000 22966 8036 22988
rect 8034 22954 8036 22966
rect 8000 22920 8002 22932
rect 8000 22894 8036 22920
rect 8034 22886 8036 22894
rect 8000 22852 8002 22860
rect 8000 22822 8036 22852
rect 8034 22818 8036 22822
rect 8000 22784 8002 22788
rect 8000 22750 8036 22784
rect 8000 22682 8036 22716
rect 8000 22678 8002 22682
rect 8034 22644 8036 22648
rect 8000 22614 8036 22644
rect 8000 22606 8002 22614
rect 8034 22572 8036 22580
rect 8000 22546 8036 22572
rect 8000 22534 8002 22546
rect 8034 22500 8036 22512
rect 8000 22478 8036 22500
rect 8000 22462 8002 22478
rect 8034 22428 8036 22444
rect 8000 22410 8036 22428
rect 8000 22390 8002 22410
rect 8034 22356 8036 22376
rect 8000 22342 8036 22356
rect 8000 22318 8002 22342
rect 8034 22284 8036 22308
rect 8000 22274 8036 22284
rect 8000 22246 8002 22274
rect 8034 22212 8036 22240
rect 8000 22206 8036 22212
rect 8000 22174 8002 22206
rect 8034 22140 8036 22172
rect 8000 22138 8036 22140
rect 6426 22085 6442 22119
rect 6476 22085 6517 22119
rect 6554 22085 6588 22119
rect 6626 22085 6656 22119
rect 6701 22085 6724 22119
rect 6776 22085 6792 22119
rect 8000 22104 8002 22138
rect 8000 22102 8036 22104
rect 8034 22070 8036 22102
rect 8000 22036 8002 22068
rect 8000 22030 8036 22036
rect 8034 22002 8036 22030
rect 8000 21968 8002 21996
rect 8000 21958 8036 21968
rect 8034 21934 8036 21958
rect 8000 21900 8002 21924
rect 8000 21886 8036 21900
rect 8034 21866 8036 21886
rect 8000 21832 8002 21852
rect 8000 21814 8036 21832
rect 8034 21798 8036 21814
rect 8000 21764 8002 21780
rect 8000 21742 8036 21764
rect 8034 21730 8036 21742
rect 8000 21696 8002 21708
rect 8000 21670 8036 21696
rect 8034 21662 8036 21670
rect 8000 21628 8002 21636
rect 6497 21570 6514 21604
rect 6565 21570 6581 21604
rect 6637 21570 6653 21604
rect 6706 21570 6721 21604
rect 8000 21598 8036 21628
rect 8034 21594 8036 21598
rect 8000 21560 8002 21564
rect 8000 21526 8036 21560
rect 8000 21458 8036 21492
rect 8000 21454 8002 21458
rect 8034 21420 8036 21424
rect 8000 21390 8036 21420
rect 8000 21382 8002 21390
rect 8034 21348 8036 21356
rect 8000 21322 8036 21348
rect 8000 21310 8002 21322
rect 8034 21276 8036 21288
rect 8000 21254 8036 21276
rect 8000 21238 8002 21254
rect 8034 21204 8036 21220
rect 8000 21186 8036 21204
rect 8000 21166 8002 21186
rect 8034 21132 8036 21152
rect 8000 21118 8036 21132
rect 8000 21094 8002 21118
rect 8034 21060 8036 21084
rect 8000 21050 8036 21060
rect 8000 21022 8002 21050
rect 8034 20988 8036 21016
rect 8000 20982 8036 20988
rect 8000 20950 8002 20982
rect 8034 20916 8036 20948
rect 8000 20914 8036 20916
rect 8000 20880 8002 20914
rect 8000 20878 8036 20880
rect 8034 20846 8036 20878
rect 8000 20812 8002 20844
rect 8000 20806 8036 20812
rect 8034 20778 8036 20806
rect 8000 20744 8002 20772
rect 8000 20734 8036 20744
rect 8034 20710 8036 20734
rect 8000 20676 8002 20700
rect 8000 20662 8036 20676
rect 8034 20642 8036 20662
rect 8000 20608 8002 20628
rect 8000 20590 8036 20608
rect 8034 20574 8036 20590
rect 8000 20540 8002 20556
rect 8000 20518 8036 20540
rect 8034 20506 8036 20518
rect 8000 20472 8002 20484
rect 8000 20446 8036 20472
rect 8034 20438 8036 20446
rect 8000 20404 8002 20412
rect 8000 20374 8036 20404
rect 8034 20370 8036 20374
rect 8000 20336 8002 20340
rect 8000 20302 8036 20336
rect 8000 20234 8036 20268
rect 8000 20230 8002 20234
rect 8034 20196 8036 20200
rect 8000 20166 8036 20196
rect 8000 20158 8002 20166
rect 8034 20124 8036 20132
rect 8000 20098 8036 20124
rect 8000 20086 8002 20098
rect 8034 20052 8036 20064
rect 8000 20030 8036 20052
rect 8000 20014 8002 20030
rect 8034 19980 8036 19996
rect 8000 19962 8036 19980
rect 8000 19942 8002 19962
rect 8034 19908 8036 19928
rect 8000 19894 8036 19908
rect 8000 19870 8002 19894
rect 8034 19836 8036 19860
rect 8000 19826 8036 19836
rect 8000 19798 8002 19826
rect 8034 19764 8036 19792
rect 8000 19758 8036 19764
rect 8000 19726 8002 19758
rect 8034 19692 8036 19724
rect 8000 19690 8036 19692
rect 8000 19656 8002 19690
rect 8000 19654 8036 19656
rect 8034 19622 8036 19654
rect 8000 19588 8002 19620
rect 8000 19582 8036 19588
rect 8034 19554 8036 19582
rect 8000 19520 8002 19548
rect 8000 19510 8036 19520
rect 8034 19486 8036 19510
rect 8000 19452 8002 19476
rect 8000 19438 8036 19452
rect 8034 19418 8036 19438
rect 8000 19384 8002 19404
rect 8000 19366 8036 19384
rect 8034 19350 8036 19366
rect 8000 19316 8002 19332
rect 8000 19294 8036 19316
rect 8034 19282 8036 19294
rect 8000 19248 8002 19260
rect 8000 19222 8036 19248
rect 8034 19214 8036 19222
rect 8000 19180 8002 19188
rect 8000 19150 8036 19180
rect 8034 19146 8036 19150
rect 8000 19112 8002 19116
rect 8000 19078 8036 19112
rect 8000 19010 8036 19044
rect 8000 19006 8002 19010
rect 8034 18972 8036 18976
rect 8000 18942 8036 18972
rect 8000 18934 8002 18942
rect 8034 18900 8036 18908
rect 8000 18874 8036 18900
rect 8000 18862 8002 18874
rect 8034 18828 8036 18840
rect 8000 18806 8036 18828
rect 8000 18790 8002 18806
rect 8034 18756 8036 18772
rect 8000 18738 8036 18756
rect 8000 18718 8002 18738
rect 8034 18684 8036 18704
rect 8000 18670 8036 18684
rect 8000 18646 8002 18670
rect 8034 18612 8036 18636
rect 8000 18602 8036 18612
rect 8000 18574 8002 18602
rect 8034 18540 8036 18568
rect 8000 18534 8036 18540
rect 8000 18502 8002 18534
rect 8034 18468 8036 18500
rect 8000 18466 8036 18468
rect 8000 18432 8002 18466
rect 8000 18430 8036 18432
rect 8034 18398 8036 18430
rect 8000 18364 8002 18396
rect 8000 18358 8036 18364
rect 8034 18330 8036 18358
rect 8000 18296 8002 18324
rect 8000 18286 8036 18296
rect 8034 18262 8036 18286
rect 8000 18228 8002 18252
rect 8000 18214 8036 18228
rect 8034 18194 8036 18214
rect 8000 18160 8002 18180
rect 8000 18142 8036 18160
rect 8034 18126 8036 18142
rect 8000 18092 8002 18108
rect 8000 18070 8036 18092
rect 8034 18058 8036 18070
rect 8000 18024 8002 18036
rect 8000 17998 8036 18024
rect 8034 17990 8036 17998
rect 8000 17956 8002 17964
rect 8000 17926 8036 17956
rect 8034 17922 8036 17926
rect 8000 17888 8002 17892
rect 8000 17854 8036 17888
rect 8000 17786 8036 17820
rect 8000 17782 8002 17786
rect 8034 17748 8036 17752
rect 8000 17718 8036 17748
rect 8000 17710 8002 17718
rect 8034 17676 8036 17684
rect 8000 17650 8036 17676
rect 8000 17638 8002 17650
rect 8034 17604 8036 17616
rect 8000 17582 8036 17604
rect 8000 17566 8002 17582
rect 8034 17532 8036 17548
rect 8000 17514 8036 17532
rect 8000 17494 8002 17514
rect 8034 17460 8036 17480
rect 8000 17446 8036 17460
rect 8000 17422 8002 17446
rect 8034 17388 8036 17412
rect 8000 17378 8036 17388
rect 8000 17350 8002 17378
rect 8034 17316 8036 17344
rect 8000 17310 8036 17316
rect 8000 17278 8002 17310
rect 8034 17244 8036 17276
rect 8000 17242 8036 17244
rect 8000 17208 8002 17242
rect 8000 17206 8036 17208
rect 8034 17174 8036 17206
rect 8000 17140 8002 17172
rect 8000 17134 8036 17140
rect 8034 17106 8036 17134
rect 8000 17072 8002 17100
rect 8000 17062 8036 17072
rect 8034 17038 8036 17062
rect 8000 17004 8002 17028
rect 8000 16990 8036 17004
rect 8034 16970 8036 16990
rect 8000 16936 8002 16956
rect 8000 16918 8036 16936
rect 8034 16902 8036 16918
rect 8000 16868 8002 16884
rect 8000 16846 8036 16868
rect 8034 16834 8036 16846
rect 8000 16800 8002 16812
rect 8000 16774 8036 16800
rect 8034 16766 8036 16774
rect 8000 16732 8002 16740
rect 8000 16702 8036 16732
rect 8034 16698 8036 16702
rect 8000 16664 8002 16668
rect 8000 16630 8036 16664
rect 8000 16562 8036 16596
rect 8000 16558 8002 16562
rect 8034 16524 8036 16528
rect 8000 16494 8036 16524
rect 8000 16486 8002 16494
rect 8034 16452 8036 16460
rect 8000 16426 8036 16452
rect 8000 16414 8002 16426
rect 8034 16380 8036 16392
rect 8000 16358 8036 16380
rect 8000 16342 8002 16358
rect 8034 16308 8036 16324
rect 8000 16290 8036 16308
rect 8000 16270 8002 16290
rect 8034 16236 8036 16256
rect 8000 16222 8036 16236
rect 8000 16198 8002 16222
rect 8034 16164 8036 16188
rect 8000 16154 8036 16164
rect 8000 16126 8002 16154
rect 8034 16092 8036 16120
rect 8000 16086 8036 16092
rect 8000 16054 8002 16086
rect 8034 16020 8036 16052
rect 8000 16018 8036 16020
rect 8000 15984 8002 16018
rect 8000 15982 8036 15984
rect 8034 15950 8036 15982
rect 8000 15916 8002 15948
rect 8000 15910 8036 15916
rect 8034 15882 8036 15910
rect 8000 15848 8002 15876
rect 8000 15838 8036 15848
rect 8034 15814 8036 15838
rect 8000 15780 8002 15804
rect 8000 15766 8036 15780
rect 8034 15746 8036 15766
rect 8000 15712 8002 15732
rect 8000 15694 8036 15712
rect 8034 15678 8036 15694
rect 8000 15644 8002 15660
rect 8000 15622 8036 15644
rect 8034 15610 8036 15622
rect 8000 15576 8002 15588
rect 8000 15550 8036 15576
rect 8034 15542 8036 15550
rect 8000 15508 8002 15516
rect 8000 15478 8036 15508
rect 8034 15474 8036 15478
rect 8000 15440 8002 15444
rect 8000 15406 8036 15440
rect 8000 15338 8036 15372
rect 8000 15334 8002 15338
rect 8034 15300 8036 15304
rect 8000 15270 8036 15300
rect 8000 15262 8002 15270
rect 8034 15228 8036 15236
rect 8000 15202 8036 15228
rect 8000 15190 8002 15202
rect 8034 15156 8036 15168
rect 8000 15134 8036 15156
rect 8000 15118 8002 15134
rect 8034 15084 8036 15100
rect 8000 15066 8036 15084
rect 8000 15046 8002 15066
rect 8034 15012 8036 15032
rect 8000 14998 8036 15012
rect 8000 14974 8002 14998
rect 8034 14940 8036 14964
rect 8000 14930 8036 14940
rect 8000 14902 8002 14930
rect 8034 14868 8036 14896
rect 8000 14862 8036 14868
rect 8000 14830 8002 14862
rect 8034 14796 8036 14828
rect 8000 14794 8036 14796
rect 8000 14760 8002 14794
rect 8000 14758 8036 14760
rect 8034 14726 8036 14758
rect 8000 14692 8002 14724
rect 8000 14686 8036 14692
rect 8034 14658 8036 14686
rect 8000 14624 8002 14652
rect 8000 14614 8036 14624
rect 8034 14590 8036 14614
rect 8000 14556 8002 14580
rect 8000 14542 8036 14556
rect 8034 14522 8036 14542
rect 8000 14488 8002 14508
rect 8000 14470 8036 14488
rect 8034 14454 8036 14470
rect 8000 14420 8002 14436
rect 8000 14398 8036 14420
rect 8034 14386 8036 14398
rect 8000 14352 8002 14364
rect 8000 14326 8036 14352
rect 8034 14318 8036 14326
rect 8000 14284 8002 14292
rect 8000 14254 8036 14284
rect 8034 14250 8036 14254
rect 8000 14216 8002 14220
rect 8000 14182 8036 14216
rect 8000 14114 8036 14148
rect 8000 14110 8002 14114
rect 8034 14076 8036 14080
rect 8000 14046 8036 14076
rect 8000 14038 8002 14046
rect 8034 14004 8036 14012
rect 8000 13978 8036 14004
rect 8000 13966 8002 13978
rect 8034 13932 8036 13944
rect 8000 13910 8036 13932
rect 8000 13894 8002 13910
rect 8034 13860 8036 13876
rect 8000 13842 8036 13860
rect 8000 13822 8002 13842
rect 8034 13788 8036 13808
rect 8000 13774 8036 13788
rect 8000 13750 8002 13774
rect 8034 13716 8036 13740
rect 8000 13706 8036 13716
rect 8000 13678 8002 13706
rect 8034 13644 8036 13672
rect 8000 13638 8036 13644
rect 8000 13606 8002 13638
rect 8034 13572 8036 13604
rect 8000 13570 8036 13572
rect 8000 13536 8002 13570
rect 8000 13534 8036 13536
rect 8034 13502 8036 13534
rect 8000 13468 8002 13500
rect 8000 13462 8036 13468
rect 8034 13434 8036 13462
rect 8000 13400 8002 13428
rect 8000 13390 8036 13400
rect 8034 13366 8036 13390
rect 8000 13332 8002 13356
rect 8000 13318 8036 13332
rect 8034 13298 8036 13318
rect 8000 13264 8002 13284
rect 8000 13246 8036 13264
rect 8034 13230 8036 13246
rect 8000 13196 8002 13212
rect 8000 13174 8036 13196
rect 8034 13162 8036 13174
rect 8000 13128 8002 13140
rect 8000 13102 8036 13128
rect 8034 13094 8036 13102
rect 8000 13060 8002 13068
rect 8000 13030 8036 13060
rect 8034 13026 8036 13030
rect 8000 12992 8002 12996
rect 8000 12958 8036 12992
rect 8000 12890 8036 12924
rect 8000 12886 8002 12890
rect 8034 12852 8036 12856
rect 8000 12822 8036 12852
rect 8000 12814 8002 12822
rect 8034 12780 8036 12788
rect 8000 12754 8036 12780
rect 8000 12742 8002 12754
rect 8034 12708 8036 12720
rect 8000 12686 8036 12708
rect 8000 12670 8002 12686
rect 8034 12636 8036 12652
rect 8000 12618 8036 12636
rect 8000 12598 8002 12618
rect 8034 12564 8036 12584
rect 8000 12550 8036 12564
rect 8000 12526 8002 12550
rect 8034 12492 8036 12516
rect 8000 12482 8036 12492
rect 8000 12454 8002 12482
rect 8034 12420 8036 12448
rect 8000 12414 8036 12420
rect 8000 12382 8002 12414
rect 8034 12348 8036 12380
rect 8000 12346 8036 12348
rect 8000 12312 8002 12346
rect 8000 12310 8036 12312
rect 8034 12278 8036 12310
rect 8000 12244 8002 12276
rect 8000 12238 8036 12244
rect 8034 12210 8036 12238
rect 8000 12176 8002 12204
rect 8000 12166 8036 12176
rect 8034 12142 8036 12166
rect 8000 12108 8002 12132
rect 8000 12094 8036 12108
rect 8034 12074 8036 12094
rect 8000 12040 8002 12060
rect 8000 12022 8036 12040
rect 8034 12006 8036 12022
rect 8000 11972 8002 11988
rect 8000 11950 8036 11972
rect 8034 11938 8036 11950
rect 8000 11904 8002 11916
rect 8000 11878 8036 11904
rect 8034 11870 8036 11878
rect 8000 11836 8002 11844
rect 8000 11806 8036 11836
rect 8034 11802 8036 11806
rect 8000 11768 8002 11772
rect 8000 11734 8036 11768
rect 8000 11666 8036 11700
rect 8000 11662 8002 11666
rect 8034 11628 8036 11632
rect 8000 11598 8036 11628
rect 8000 11590 8002 11598
rect 8034 11556 8036 11564
rect 8000 11530 8036 11556
rect 8000 11518 8002 11530
rect 8034 11484 8036 11496
rect 8000 11462 8036 11484
rect 8000 11446 8002 11462
rect 8034 11412 8036 11428
rect 2796 11399 7477 11405
rect 2796 11365 2879 11399
rect 2913 11365 2926 11399
rect 2990 11365 2994 11399
rect 3028 11365 3033 11399
rect 3096 11365 3110 11399
rect 3164 11365 3188 11399
rect 3232 11365 3266 11399
rect 3300 11365 3334 11399
rect 3378 11365 3402 11399
rect 3456 11365 3470 11399
rect 3534 11365 3538 11399
rect 3572 11365 3578 11399
rect 3640 11365 3656 11399
rect 3708 11365 3742 11399
rect 3800 11365 3810 11399
rect 3873 11365 3878 11399
rect 3980 11365 3985 11399
rect 4048 11365 4058 11399
rect 4116 11365 4131 11399
rect 4184 11365 4204 11399
rect 4252 11365 4277 11399
rect 4320 11365 4350 11399
rect 4388 11365 4422 11399
rect 4457 11365 4490 11399
rect 4530 11365 4558 11399
rect 4603 11365 4626 11399
rect 4676 11365 4694 11399
rect 4749 11365 4762 11399
rect 4822 11365 4830 11399
rect 4895 11365 4898 11399
rect 4932 11365 4934 11399
rect 5000 11365 5007 11399
rect 5068 11365 5080 11399
rect 5136 11365 5153 11399
rect 5204 11365 5226 11399
rect 5272 11365 5299 11399
rect 5340 11365 5372 11399
rect 5408 11365 5442 11399
rect 5479 11365 5510 11399
rect 5552 11365 5578 11399
rect 5625 11365 5646 11399
rect 5698 11365 5714 11399
rect 5771 11365 5782 11399
rect 5845 11365 5850 11399
rect 5884 11365 5885 11399
rect 5952 11365 5959 11399
rect 6020 11365 6033 11399
rect 6088 11365 6107 11399
rect 6156 11365 6181 11399
rect 6224 11365 6255 11399
rect 6292 11365 6326 11399
rect 6363 11365 6394 11399
rect 6437 11365 6477 11399
rect 6511 11365 6551 11399
rect 6587 11365 6621 11399
rect 6659 11365 6689 11399
rect 6733 11365 6757 11399
rect 6807 11365 6825 11399
rect 6881 11365 6893 11399
rect 6955 11365 6961 11399
rect 7063 11365 7069 11399
rect 7131 11365 7143 11399
rect 7199 11365 7217 11399
rect 7267 11365 7291 11399
rect 7335 11365 7365 11399
rect 7403 11365 7477 11399
rect 2796 11359 7477 11365
rect 2796 11331 2842 11359
rect 2796 11293 2802 11331
rect 2836 11293 2842 11331
rect 2796 11263 2842 11293
rect 2796 11220 2802 11263
rect 2836 11220 2842 11263
rect 2796 11195 2842 11220
rect 2796 11147 2802 11195
rect 2836 11147 2842 11195
rect 2796 11127 2842 11147
rect 2796 11074 2802 11127
rect 2836 11074 2842 11127
rect 2796 11059 2842 11074
rect 2796 11001 2802 11059
rect 2836 11001 2842 11059
rect 2796 10991 2842 11001
rect 2796 10928 2802 10991
rect 2836 10928 2842 10991
rect 2796 10923 2842 10928
rect 2796 10821 2802 10923
rect 2836 10821 2842 10923
rect 2796 10816 2842 10821
rect 2796 10753 2802 10816
rect 2836 10753 2842 10816
rect 2796 10743 2842 10753
rect 2796 10685 2802 10743
rect 2836 10685 2842 10743
rect 2796 10670 2842 10685
rect 2796 10617 2802 10670
rect 2836 10617 2842 10670
rect 2796 10597 2842 10617
rect 2796 10549 2802 10597
rect 2836 10549 2842 10597
rect 2796 10524 2842 10549
rect 2796 10481 2802 10524
rect 2836 10481 2842 10524
rect 2796 10451 2842 10481
rect 2796 10413 2802 10451
rect 2836 10413 2842 10451
rect 2796 10379 2842 10413
rect 2796 10344 2802 10379
rect 2836 10344 2842 10379
rect 2796 10311 2842 10344
rect 2796 10271 2802 10311
rect 2836 10271 2842 10311
rect 2796 10243 2842 10271
rect 2796 10198 2802 10243
rect 2836 10198 2842 10243
rect 2796 10175 2842 10198
rect 2796 10125 2802 10175
rect 2836 10125 2842 10175
rect 2796 10107 2842 10125
rect 2796 10052 2802 10107
rect 2836 10052 2842 10107
rect 2796 10039 2842 10052
rect 2796 9979 2802 10039
rect 2836 9979 2842 10039
rect 2796 9971 2842 9979
rect 2796 9906 2802 9971
rect 2836 9906 2842 9971
rect 2796 9903 2842 9906
rect 2796 9869 2802 9903
rect 2836 9869 2842 9903
rect 2796 9867 2842 9869
rect 2796 9801 2802 9867
rect 2836 9801 2842 9867
rect 2796 9794 2842 9801
rect 2796 9733 2802 9794
rect 2836 9733 2842 9794
rect 2796 9721 2842 9733
rect 2796 9665 2802 9721
rect 2836 9665 2842 9721
rect 2796 9648 2842 9665
rect 2796 9597 2802 9648
rect 2836 9597 2842 9648
rect 2796 9575 2842 9597
rect 2796 9529 2802 9575
rect 2836 9529 2842 9575
rect 2796 9502 2842 9529
rect 2796 9461 2802 9502
rect 2836 9461 2842 9502
rect 2796 9429 2842 9461
rect 2796 9393 2802 9429
rect 2836 9393 2842 9429
rect 2796 9359 2842 9393
rect 2796 9322 2802 9359
rect 2836 9322 2842 9359
rect 2796 9291 2842 9322
rect 2796 9249 2802 9291
rect 2836 9249 2842 9291
rect 2796 9223 2842 9249
rect 2796 9176 2802 9223
rect 2836 9176 2842 9223
rect 2796 9155 2842 9176
rect 2796 9103 2802 9155
rect 2836 9103 2842 9155
rect 2796 9087 2842 9103
rect 2796 9030 2802 9087
rect 2836 9030 2842 9087
rect 2796 9019 2842 9030
rect 2796 8957 2802 9019
rect 2836 8957 2842 9019
rect 2796 8951 2842 8957
rect 2796 8884 2802 8951
rect 2836 8884 2842 8951
rect 2796 8883 2842 8884
rect 2796 8849 2802 8883
rect 2836 8849 2842 8883
rect 2796 8845 2842 8849
rect 2796 8781 2802 8845
rect 2836 8781 2842 8845
rect 2796 8772 2842 8781
rect 2796 8713 2802 8772
rect 2836 8713 2842 8772
rect 2796 8699 2842 8713
rect 2796 8645 2802 8699
rect 2836 8645 2842 8699
rect 2796 8626 2842 8645
rect 2796 8577 2802 8626
rect 2836 8577 2842 8626
rect 2796 8553 2842 8577
rect 2796 8509 2802 8553
rect 2836 8509 2842 8553
rect 2796 8480 2842 8509
rect 2796 8441 2802 8480
rect 2836 8441 2842 8480
rect 2796 8407 2842 8441
rect 2796 8373 2802 8407
rect 2836 8373 2842 8407
rect 2796 8339 2842 8373
rect 2796 8300 2802 8339
rect 2836 8300 2842 8339
rect 2796 8271 2842 8300
rect 2796 8227 2802 8271
rect 2836 8227 2842 8271
rect 2796 8203 2842 8227
rect 2796 8154 2802 8203
rect 2836 8154 2842 8203
rect 2796 8135 2842 8154
rect 2796 8081 2802 8135
rect 2836 8081 2842 8135
rect 7431 11325 7477 11359
rect 7431 11284 7437 11325
rect 7471 11284 7477 11325
rect 7431 11251 7477 11284
rect 7431 11216 7437 11251
rect 7471 11216 7477 11251
rect 7431 11182 7477 11216
rect 7431 11143 7437 11182
rect 7471 11143 7477 11182
rect 7431 11114 7477 11143
rect 7431 11069 7437 11114
rect 7471 11069 7477 11114
rect 7431 11046 7477 11069
rect 7431 10995 7437 11046
rect 7471 10995 7477 11046
rect 7431 10978 7477 10995
rect 7431 10921 7437 10978
rect 7471 10921 7477 10978
rect 7431 10910 7477 10921
rect 7431 10846 7437 10910
rect 7471 10846 7477 10910
rect 7431 10842 7477 10846
rect 7431 10808 7437 10842
rect 7471 10808 7477 10842
rect 7431 10805 7477 10808
rect 7431 10740 7437 10805
rect 7471 10740 7477 10805
rect 7431 10730 7477 10740
rect 7431 10672 7437 10730
rect 7471 10672 7477 10730
rect 7431 10655 7477 10672
rect 7431 10604 7437 10655
rect 7471 10604 7477 10655
rect 7431 10580 7477 10604
rect 7431 10536 7437 10580
rect 7471 10536 7477 10580
rect 7431 10505 7477 10536
rect 7431 10468 7437 10505
rect 7471 10468 7477 10505
rect 7431 10434 7477 10468
rect 7431 10367 7437 10434
rect 7471 10367 7477 10434
rect 7431 10366 7477 10367
rect 7431 10332 7437 10366
rect 7471 10332 7477 10366
rect 7431 10328 7477 10332
rect 7431 10264 7437 10328
rect 7471 10264 7477 10328
rect 7431 10255 7477 10264
rect 7431 10196 7437 10255
rect 7471 10196 7477 10255
rect 7431 10182 7477 10196
rect 7431 10128 7437 10182
rect 7471 10128 7477 10182
rect 7431 10108 7477 10128
rect 7431 10060 7437 10108
rect 7471 10060 7477 10108
rect 7431 10034 7477 10060
rect 7431 9992 7437 10034
rect 7471 9992 7477 10034
rect 7431 9960 7477 9992
rect 7431 9924 7437 9960
rect 7471 9924 7477 9960
rect 7431 9890 7477 9924
rect 7431 9852 7437 9890
rect 7471 9852 7477 9890
rect 7431 9822 7477 9852
rect 7431 9778 7437 9822
rect 7471 9778 7477 9822
rect 7431 9754 7477 9778
rect 7431 9704 7437 9754
rect 7471 9704 7477 9754
rect 7431 9686 7477 9704
rect 7431 9630 7437 9686
rect 7471 9630 7477 9686
rect 7431 9618 7477 9630
rect 7431 9556 7437 9618
rect 7471 9556 7477 9618
rect 7431 9516 7477 9556
rect 7431 9482 7437 9516
rect 7471 9482 7477 9516
rect 7431 9472 7477 9482
rect 7431 9408 7437 9472
rect 7471 9408 7477 9472
rect 7431 9404 7477 9408
rect 7431 9370 7437 9404
rect 7471 9370 7477 9404
rect 7431 9368 7477 9370
rect 7431 9302 7437 9368
rect 7471 9302 7477 9368
rect 7431 9294 7477 9302
rect 7431 9234 7437 9294
rect 7471 9234 7477 9294
rect 7431 9220 7477 9234
rect 7431 9166 7437 9220
rect 7471 9166 7477 9220
rect 7431 9146 7477 9166
rect 7431 9098 7437 9146
rect 7471 9098 7477 9146
rect 7431 9072 7477 9098
rect 7431 9030 7437 9072
rect 7471 9030 7477 9072
rect 7431 8998 7477 9030
rect 7431 8962 7437 8998
rect 7471 8962 7477 8998
rect 7431 8928 7477 8962
rect 7431 8890 7437 8928
rect 7471 8890 7477 8928
rect 7431 8860 7477 8890
rect 7431 8816 7437 8860
rect 7471 8816 7477 8860
rect 7431 8792 7477 8816
rect 7431 8742 7437 8792
rect 7471 8742 7477 8792
rect 7431 8724 7477 8742
rect 7431 8668 7437 8724
rect 7471 8668 7477 8724
rect 7431 8656 7477 8668
rect 7431 8594 7437 8656
rect 7471 8594 7477 8656
rect 7431 8588 7477 8594
rect 7431 8486 7437 8588
rect 7471 8486 7477 8588
rect 7431 8480 7477 8486
rect 7431 8418 7437 8480
rect 7471 8418 7477 8480
rect 7431 8406 7477 8418
rect 7431 8350 7437 8406
rect 7471 8350 7477 8406
rect 7431 8332 7477 8350
rect 7431 8282 7437 8332
rect 7471 8282 7477 8332
rect 7431 8258 7477 8282
rect 7431 8214 7437 8258
rect 7471 8214 7477 8258
rect 7431 8184 7477 8214
rect 7431 8146 7437 8184
rect 7471 8146 7477 8184
rect 2796 8067 2842 8081
rect 2796 8008 2802 8067
rect 2836 8008 2842 8067
rect 2796 7999 2842 8008
rect 2796 7935 2802 7999
rect 2836 7935 2842 7999
rect 2796 7931 2842 7935
rect 2796 7897 2802 7931
rect 2836 7920 2842 7931
rect 6744 8112 6790 8126
rect 7431 8118 7477 8146
rect 7016 8112 7477 8118
rect 6744 8094 6862 8112
rect 6744 8060 6750 8094
rect 6784 8078 6862 8094
rect 6896 8078 6930 8112
rect 6964 8078 6998 8112
rect 7032 8078 7048 8112
rect 7082 8078 7100 8112
rect 7160 8078 7168 8112
rect 7202 8078 7204 8112
rect 7270 8078 7282 8112
rect 7338 8078 7360 8112
rect 7394 8078 7477 8112
rect 6784 8060 6790 8078
rect 7016 8072 7477 8078
rect 8000 11394 8036 11412
rect 8000 11374 8002 11394
rect 8034 11340 8036 11360
rect 8000 11326 8036 11340
rect 8000 11302 8002 11326
rect 8034 11268 8036 11292
rect 8000 11258 8036 11268
rect 8000 11230 8002 11258
rect 8034 11196 8036 11224
rect 8000 11190 8036 11196
rect 8000 11158 8002 11190
rect 8034 11124 8036 11156
rect 8000 11122 8036 11124
rect 8000 11088 8002 11122
rect 8000 11086 8036 11088
rect 8034 11054 8036 11086
rect 8000 11020 8002 11052
rect 8000 11014 8036 11020
rect 8034 10986 8036 11014
rect 8000 10952 8002 10980
rect 8000 10942 8036 10952
rect 8034 10918 8036 10942
rect 8000 10884 8002 10908
rect 8000 10870 8036 10884
rect 8034 10850 8036 10870
rect 8000 10816 8002 10836
rect 8000 10798 8036 10816
rect 8034 10782 8036 10798
rect 8000 10748 8002 10764
rect 8000 10726 8036 10748
rect 8034 10714 8036 10726
rect 8000 10680 8002 10692
rect 8000 10654 8036 10680
rect 8034 10646 8036 10654
rect 8000 10612 8002 10620
rect 8000 10582 8036 10612
rect 8034 10578 8036 10582
rect 8000 10544 8002 10548
rect 8000 10510 8036 10544
rect 8000 10442 8036 10476
rect 8000 10438 8002 10442
rect 8034 10404 8036 10408
rect 8000 10374 8036 10404
rect 8000 10366 8002 10374
rect 8034 10332 8036 10340
rect 8000 10306 8036 10332
rect 8000 10294 8002 10306
rect 8034 10260 8036 10272
rect 8000 10238 8036 10260
rect 8000 10222 8002 10238
rect 8034 10188 8036 10204
rect 8000 10170 8036 10188
rect 8000 10150 8002 10170
rect 8034 10116 8036 10136
rect 8000 10102 8036 10116
rect 8000 10078 8002 10102
rect 8034 10044 8036 10068
rect 8000 10034 8036 10044
rect 8000 10006 8002 10034
rect 8034 9972 8036 10000
rect 8000 9966 8036 9972
rect 8000 9934 8002 9966
rect 8034 9900 8036 9932
rect 8000 9898 8036 9900
rect 8000 9864 8002 9898
rect 8000 9862 8036 9864
rect 8034 9830 8036 9862
rect 8000 9796 8002 9828
rect 8000 9790 8036 9796
rect 8034 9762 8036 9790
rect 8000 9728 8002 9756
rect 8000 9718 8036 9728
rect 8034 9694 8036 9718
rect 8000 9660 8002 9684
rect 8000 9646 8036 9660
rect 8034 9626 8036 9646
rect 8000 9592 8002 9612
rect 8000 9574 8036 9592
rect 8034 9558 8036 9574
rect 8000 9524 8002 9540
rect 8000 9502 8036 9524
rect 8034 9490 8036 9502
rect 8000 9456 8002 9468
rect 8000 9430 8036 9456
rect 8034 9422 8036 9430
rect 8000 9388 8002 9396
rect 8000 9358 8036 9388
rect 8034 9354 8036 9358
rect 8000 9320 8002 9324
rect 8000 9286 8036 9320
rect 8000 9218 8036 9252
rect 8000 9214 8002 9218
rect 8034 9180 8036 9184
rect 8000 9150 8036 9180
rect 8000 9142 8002 9150
rect 8034 9108 8036 9116
rect 8000 9082 8036 9108
rect 8000 9070 8002 9082
rect 8034 9036 8036 9048
rect 8000 9014 8036 9036
rect 8000 8998 8002 9014
rect 8034 8964 8036 8980
rect 8000 8946 8036 8964
rect 8000 8926 8002 8946
rect 8034 8892 8036 8912
rect 8000 8878 8036 8892
rect 8000 8854 8002 8878
rect 8034 8820 8036 8844
rect 8000 8810 8036 8820
rect 8000 8782 8002 8810
rect 8034 8748 8036 8776
rect 8000 8742 8036 8748
rect 8000 8710 8002 8742
rect 8034 8676 8036 8708
rect 8000 8674 8036 8676
rect 8000 8640 8002 8674
rect 8000 8638 8036 8640
rect 8034 8606 8036 8638
rect 8000 8572 8002 8604
rect 8000 8566 8036 8572
rect 8034 8538 8036 8566
rect 8000 8504 8002 8532
rect 8000 8494 8036 8504
rect 8034 8470 8036 8494
rect 8000 8436 8002 8460
rect 8000 8422 8036 8436
rect 8034 8402 8036 8422
rect 8000 8368 8002 8388
rect 8000 8350 8036 8368
rect 8034 8334 8036 8350
rect 8000 8300 8002 8316
rect 8000 8278 8036 8300
rect 8034 8266 8036 8278
rect 8000 8232 8002 8244
rect 8000 8206 8036 8232
rect 8034 8198 8036 8206
rect 8000 8164 8002 8172
rect 8000 8134 8036 8164
rect 8034 8130 8036 8134
rect 8000 8096 8002 8100
rect 6744 8044 6790 8060
rect 6744 8010 6750 8044
rect 6784 8010 6790 8044
rect 6744 7992 6790 8010
rect 6744 7958 6750 7992
rect 6784 7958 6790 7992
rect 6744 7920 6790 7958
rect 2836 7897 2870 7920
rect 2796 7896 2870 7897
rect 2796 7829 2802 7896
rect 2836 7886 2870 7896
rect 2904 7886 2938 7920
rect 2972 7886 3006 7920
rect 3040 7886 3074 7920
rect 3108 7886 3142 7920
rect 3176 7886 3210 7920
rect 3244 7886 3278 7920
rect 3312 7886 3346 7920
rect 3380 7886 3414 7920
rect 3448 7886 3482 7920
rect 3516 7886 3550 7920
rect 3584 7886 3618 7920
rect 3652 7886 3686 7920
rect 3720 7886 3754 7920
rect 3788 7886 3822 7920
rect 3856 7886 3890 7920
rect 3924 7886 3958 7920
rect 3992 7886 4026 7920
rect 4060 7886 4094 7920
rect 4128 7886 4162 7920
rect 4196 7886 4230 7920
rect 4264 7886 4298 7920
rect 4332 7886 4366 7920
rect 4400 7886 4434 7920
rect 4468 7886 4502 7920
rect 4536 7886 4570 7920
rect 4604 7886 4638 7920
rect 4672 7886 4706 7920
rect 4740 7886 4774 7920
rect 4808 7886 4842 7920
rect 4876 7886 4910 7920
rect 4944 7886 4978 7920
rect 5012 7886 5046 7920
rect 5080 7886 5114 7920
rect 5148 7886 5182 7920
rect 5216 7886 5250 7920
rect 5284 7886 5318 7920
rect 5352 7886 5386 7920
rect 5420 7886 5454 7920
rect 5488 7886 5522 7920
rect 5556 7886 5590 7920
rect 5624 7886 5658 7920
rect 5692 7886 5726 7920
rect 5760 7886 5794 7920
rect 5828 7886 5862 7920
rect 5896 7886 5930 7920
rect 5964 7886 5998 7920
rect 6032 7886 6066 7920
rect 6100 7886 6134 7920
rect 6168 7886 6202 7920
rect 6236 7886 6270 7920
rect 6304 7886 6338 7920
rect 6372 7886 6406 7920
rect 6440 7886 6474 7920
rect 6508 7886 6542 7920
rect 6576 7886 6610 7920
rect 6644 7886 6678 7920
rect 6712 7897 6790 7920
rect 6712 7886 6750 7897
rect 2836 7829 2842 7886
rect 2796 7823 2842 7829
rect 2796 7761 2802 7823
rect 2836 7761 2842 7823
rect 2796 7750 2842 7761
rect 2796 7693 2802 7750
rect 2836 7693 2842 7750
rect 6744 7854 6750 7886
rect 6784 7854 6790 7897
rect 6744 7829 6790 7854
rect 6744 7781 6750 7829
rect 6784 7781 6790 7829
rect 6744 7761 6790 7781
rect 2796 7677 2842 7693
rect 2796 7625 2802 7677
rect 2836 7625 2842 7677
rect 2796 7604 2842 7625
rect 2796 7557 2802 7604
rect 2836 7557 2842 7604
rect 2796 7531 2842 7557
rect 2796 7489 2802 7531
rect 2836 7489 2842 7531
rect 2796 7458 2842 7489
rect 2796 7421 2802 7458
rect 2836 7421 2842 7458
rect 2796 7387 2842 7421
rect 2796 7351 2802 7387
rect 2836 7351 2842 7387
rect 2796 7319 2842 7351
rect 2796 7278 2802 7319
rect 2836 7278 2842 7319
rect 2796 7251 2842 7278
rect 2796 7205 2802 7251
rect 2836 7205 2842 7251
rect 2796 7183 2842 7205
rect 2796 7132 2802 7183
rect 2836 7132 2842 7183
rect 2796 7115 2842 7132
rect 2796 7059 2802 7115
rect 2836 7059 2842 7115
rect 2796 7047 2842 7059
rect 2796 6986 2802 7047
rect 2836 6986 2842 7047
rect 2796 6979 2842 6986
rect 2796 6913 2802 6979
rect 2836 6913 2842 6979
rect 2796 6911 2842 6913
rect 2796 6877 2802 6911
rect 2836 6877 2842 6911
rect 2796 6874 2842 6877
rect 2796 6809 2802 6874
rect 2836 6809 2842 6874
rect 2796 6801 2842 6809
rect 2796 6741 2802 6801
rect 2836 6741 2842 6801
rect 2796 6729 2842 6741
rect 2796 6673 2802 6729
rect 2836 6673 2842 6729
rect 2796 6657 2842 6673
rect 2796 6605 2802 6657
rect 2836 6605 2842 6657
rect 2796 6585 2842 6605
rect 2796 6537 2802 6585
rect 2836 6537 2842 6585
rect 2796 6513 2842 6537
rect 2796 6469 2802 6513
rect 2836 6469 2842 6513
rect 2796 6441 2842 6469
rect 2796 6401 2802 6441
rect 2836 6401 2842 6441
rect 2796 6369 2842 6401
rect 2796 6333 2802 6369
rect 2836 6333 2842 6369
rect 2796 6299 2842 6333
rect 2796 6263 2802 6299
rect 2836 6263 2842 6299
rect 2796 6231 2842 6263
rect 2796 6191 2802 6231
rect 2836 6191 2842 6231
rect 2796 6163 2842 6191
rect 2796 6119 2802 6163
rect 2836 6119 2842 6163
rect 2796 6095 2842 6119
rect 2796 6047 2802 6095
rect 2836 6047 2842 6095
rect 2796 6027 2842 6047
rect 2796 5975 2802 6027
rect 2836 5975 2842 6027
rect 2796 5959 2842 5975
rect 2796 5903 2802 5959
rect 2836 5903 2842 5959
rect 2796 5891 2842 5903
rect 2796 5831 2802 5891
rect 2836 5831 2842 5891
rect 2796 5823 2842 5831
rect 2796 5759 2802 5823
rect 2836 5759 2842 5823
rect 2796 5755 2842 5759
rect 2796 5653 2802 5755
rect 2836 5653 2842 5755
rect 2796 5649 2842 5653
rect 2796 5585 2802 5649
rect 2836 5585 2842 5649
rect 2796 5577 2842 5585
rect 2796 5517 2802 5577
rect 2836 5517 2842 5577
rect 2796 5505 2842 5517
rect 2796 5449 2802 5505
rect 2836 5449 2842 5505
rect 2796 5433 2842 5449
rect 2796 5381 2802 5433
rect 2836 5381 2842 5433
rect 2796 5361 2842 5381
rect 2796 5313 2802 5361
rect 2836 5313 2842 5361
rect 2796 5289 2842 5313
rect 2796 5245 2802 5289
rect 2836 5245 2842 5289
rect 3076 7723 6530 7729
rect 3076 7689 3158 7723
rect 3198 7689 3226 7723
rect 3280 7689 3294 7723
rect 3396 7689 3411 7723
rect 3464 7689 3494 7723
rect 3532 7689 3566 7723
rect 3600 7689 3604 7723
rect 3668 7689 3676 7723
rect 3736 7689 3748 7723
rect 3804 7689 3820 7723
rect 3872 7689 3892 7723
rect 3940 7689 3964 7723
rect 4008 7689 4036 7723
rect 4076 7689 4108 7723
rect 4144 7689 4178 7723
rect 4214 7689 4246 7723
rect 4286 7689 4314 7723
rect 4358 7689 4382 7723
rect 4430 7689 4450 7723
rect 4502 7689 4518 7723
rect 4574 7689 4586 7723
rect 4646 7689 4654 7723
rect 4718 7689 4722 7723
rect 4824 7689 4828 7723
rect 4892 7689 4900 7723
rect 4960 7689 4972 7723
rect 5028 7689 5044 7723
rect 5096 7689 5116 7723
rect 5164 7689 5188 7723
rect 5232 7689 5260 7723
rect 5300 7689 5332 7723
rect 5368 7689 5402 7723
rect 5438 7689 5470 7723
rect 5510 7689 5538 7723
rect 5582 7689 5606 7723
rect 5654 7689 5674 7723
rect 5726 7689 5742 7723
rect 5798 7689 5810 7723
rect 5870 7689 5878 7723
rect 5942 7689 5946 7723
rect 6048 7689 6053 7723
rect 6116 7689 6126 7723
rect 6184 7689 6199 7723
rect 6252 7689 6272 7723
rect 6320 7689 6345 7723
rect 6388 7689 6418 7723
rect 6456 7689 6530 7723
rect 3076 7683 6530 7689
rect 3076 7655 3122 7683
rect 3076 7617 3082 7655
rect 3116 7617 3122 7655
rect 3076 7587 3122 7617
rect 3076 7543 3082 7587
rect 3116 7543 3122 7587
rect 3076 7519 3122 7543
rect 3076 7469 3082 7519
rect 3116 7469 3122 7519
rect 3076 7451 3122 7469
rect 3076 7395 3082 7451
rect 3116 7395 3122 7451
rect 3076 7383 3122 7395
rect 3076 7321 3082 7383
rect 3116 7321 3122 7383
rect 3076 7315 3122 7321
rect 3076 7213 3082 7315
rect 3116 7213 3122 7315
rect 5344 7655 5390 7683
rect 5344 7617 5350 7655
rect 5384 7617 5390 7655
rect 5344 7586 5390 7617
rect 5344 7544 5350 7586
rect 5384 7544 5390 7586
rect 5344 7517 5390 7544
rect 5344 7471 5350 7517
rect 5384 7471 5390 7517
rect 5344 7448 5390 7471
rect 5344 7398 5350 7448
rect 5384 7398 5390 7448
rect 5344 7379 5390 7398
rect 5344 7325 5350 7379
rect 5384 7325 5390 7379
rect 5344 7310 5390 7325
rect 3076 7207 3122 7213
rect 3076 7145 3082 7207
rect 3116 7145 3122 7207
rect 3076 7133 3122 7145
rect 3076 7077 3082 7133
rect 3116 7077 3122 7133
rect 3076 7059 3122 7077
rect 3076 7009 3082 7059
rect 3116 7009 3122 7059
rect 3076 6985 3122 7009
rect 3076 6941 3082 6985
rect 3116 6941 3122 6985
rect 3076 6911 3122 6941
rect 3076 6873 3082 6911
rect 3116 6873 3122 6911
rect 3076 6839 3122 6873
rect 3076 6803 3082 6839
rect 3116 6803 3122 6839
rect 3076 6771 3122 6803
rect 3076 6729 3082 6771
rect 3116 6729 3122 6771
rect 3076 6703 3122 6729
rect 3076 6655 3082 6703
rect 3116 6655 3122 6703
rect 3076 6635 3122 6655
rect 3076 6581 3082 6635
rect 3116 6581 3122 6635
rect 3076 6567 3122 6581
rect 3076 6508 3082 6567
rect 3116 6508 3122 6567
rect 3076 6499 3122 6508
rect 3076 6435 3082 6499
rect 3116 6435 3122 6499
rect 3076 6431 3122 6435
rect 3076 6397 3082 6431
rect 3116 6397 3122 6431
rect 3076 6396 3122 6397
rect 3076 6329 3082 6396
rect 3116 6329 3122 6396
rect 3076 6323 3122 6329
rect 3076 6261 3082 6323
rect 3116 6261 3122 6323
rect 3076 6250 3122 6261
rect 3076 6193 3082 6250
rect 3116 6193 3122 6250
rect 3076 6177 3122 6193
rect 3076 6125 3082 6177
rect 3116 6125 3122 6177
rect 3076 6104 3122 6125
rect 3076 6057 3082 6104
rect 3116 6057 3122 6104
rect 3076 6031 3122 6057
rect 3076 5989 3082 6031
rect 3116 5989 3122 6031
rect 3076 5958 3122 5989
rect 3076 5921 3082 5958
rect 3116 5921 3122 5958
rect 3076 5887 3122 5921
rect 3076 5851 3082 5887
rect 3116 5851 3122 5887
rect 3076 5819 3122 5851
rect 3076 5778 3082 5819
rect 3116 5778 3122 5819
rect 3076 5751 3122 5778
rect 3076 5705 3082 5751
rect 3116 5705 3122 5751
rect 3076 5683 3122 5705
rect 3076 5632 3082 5683
rect 3116 5632 3122 5683
rect 3856 7265 3890 7281
rect 3856 7196 3890 7231
rect 3856 7127 3890 7159
rect 3856 7058 3890 7085
rect 3856 6989 3890 7011
rect 3856 6920 3890 6937
rect 3856 6851 3890 6863
rect 3856 6781 3890 6789
rect 3856 6711 3890 6715
rect 3856 6675 3890 6677
rect 3856 6601 3890 6607
rect 3856 6527 3890 6537
rect 3856 6452 3890 6467
rect 3856 6377 3890 6397
rect 3856 6302 3890 6327
rect 3856 6227 3890 6257
rect 3856 6152 3890 6187
rect 3856 6081 3890 6117
rect 3856 6011 3890 6043
rect 3856 5941 3890 5968
rect 3856 5871 3890 5893
rect 3856 5801 3890 5818
rect 3856 5731 3890 5743
rect 3856 5681 3890 5697
rect 4586 7265 4620 7281
rect 4586 7196 4620 7231
rect 4586 7127 4620 7159
rect 4586 7058 4620 7085
rect 4586 6989 4620 7011
rect 4586 6920 4620 6937
rect 4586 6851 4620 6863
rect 4586 6781 4620 6789
rect 4586 6711 4620 6715
rect 4586 6675 4620 6677
rect 4586 6601 4620 6607
rect 4586 6527 4620 6537
rect 4586 6452 4620 6467
rect 4586 6377 4620 6397
rect 4586 6302 4620 6327
rect 4586 6227 4620 6257
rect 4586 6152 4620 6187
rect 4586 6081 4620 6117
rect 4586 6011 4620 6043
rect 4586 5941 4620 5968
rect 4586 5871 4620 5893
rect 4586 5801 4620 5818
rect 4586 5731 4620 5743
rect 4586 5681 4620 5697
rect 5344 7252 5350 7310
rect 5384 7252 5390 7310
rect 5344 7241 5390 7252
rect 5344 7179 5350 7241
rect 5384 7179 5390 7241
rect 5344 7172 5390 7179
rect 5344 7106 5350 7172
rect 5384 7106 5390 7172
rect 6484 7650 6530 7683
rect 6484 7616 6490 7650
rect 6524 7616 6530 7650
rect 6484 7613 6530 7616
rect 6484 7579 6490 7613
rect 6524 7579 6530 7613
rect 6484 7577 6530 7579
rect 6484 7511 6490 7577
rect 6524 7511 6530 7577
rect 6484 7504 6530 7511
rect 6484 7443 6490 7504
rect 6524 7443 6530 7504
rect 6484 7431 6530 7443
rect 6484 7375 6490 7431
rect 6524 7375 6530 7431
rect 6484 7358 6530 7375
rect 6484 7307 6490 7358
rect 6524 7307 6530 7358
rect 6484 7285 6530 7307
rect 6484 7239 6490 7285
rect 6524 7239 6530 7285
rect 6484 7212 6530 7239
rect 6484 7171 6490 7212
rect 6524 7171 6530 7212
rect 6484 7139 6530 7171
rect 5344 7103 5390 7106
rect 5344 7069 5350 7103
rect 5384 7069 5390 7103
rect 5344 7067 5390 7069
rect 5344 7000 5350 7067
rect 5384 7000 5390 7067
rect 5344 6994 5390 7000
rect 5344 6931 5350 6994
rect 5384 6931 5390 6994
rect 5344 6921 5390 6931
rect 5344 6862 5350 6921
rect 5384 6862 5390 6921
rect 5344 6848 5390 6862
rect 5344 6793 5350 6848
rect 5384 6793 5390 6848
rect 5344 6775 5390 6793
rect 5344 6724 5350 6775
rect 5384 6724 5390 6775
rect 6100 7108 6134 7124
rect 6100 7046 6134 7074
rect 6100 6954 6134 6991
rect 6100 6862 6134 6908
rect 6100 6774 6134 6824
rect 6100 6724 6134 6736
rect 6484 7103 6490 7139
rect 6524 7103 6530 7139
rect 6484 7069 6530 7103
rect 6484 7032 6490 7069
rect 6524 7032 6530 7069
rect 6484 7001 6530 7032
rect 6484 6959 6490 7001
rect 6524 6959 6530 7001
rect 6484 6933 6530 6959
rect 6484 6886 6490 6933
rect 6524 6886 6530 6933
rect 6484 6865 6530 6886
rect 6484 6813 6490 6865
rect 6524 6813 6530 6865
rect 6484 6797 6530 6813
rect 6484 6740 6490 6797
rect 6524 6740 6530 6797
rect 6484 6729 6530 6740
rect 5344 6702 5390 6724
rect 5344 6655 5350 6702
rect 5384 6655 5390 6702
rect 5344 6629 5390 6655
rect 5344 6586 5350 6629
rect 5384 6586 5390 6629
rect 5344 6556 5390 6586
rect 5344 6517 5350 6556
rect 5384 6517 5390 6556
rect 6484 6667 6490 6729
rect 6524 6667 6530 6729
rect 6484 6661 6530 6667
rect 6484 6594 6490 6661
rect 6524 6594 6530 6661
rect 6484 6593 6530 6594
rect 6484 6559 6490 6593
rect 6524 6559 6530 6593
rect 6484 6555 6530 6559
rect 5344 6483 5390 6517
rect 5344 6448 5350 6483
rect 5384 6448 5390 6483
rect 5344 6413 5390 6448
rect 5344 6375 5350 6413
rect 5384 6375 5390 6413
rect 5344 6344 5390 6375
rect 5344 6301 5350 6344
rect 5384 6301 5390 6344
rect 5344 6275 5390 6301
rect 5344 6227 5350 6275
rect 5384 6227 5390 6275
rect 5344 6206 5390 6227
rect 5344 6153 5350 6206
rect 5384 6153 5390 6206
rect 5344 6137 5390 6153
rect 5344 6079 5350 6137
rect 5384 6079 5390 6137
rect 5344 6068 5390 6079
rect 5344 6005 5350 6068
rect 5384 6005 5390 6068
rect 5344 5999 5390 6005
rect 5344 5931 5350 5999
rect 5384 5931 5390 5999
rect 5344 5929 5390 5931
rect 5344 5895 5350 5929
rect 5384 5895 5390 5929
rect 5344 5891 5390 5895
rect 5344 5825 5350 5891
rect 5384 5825 5390 5891
rect 5344 5817 5390 5825
rect 5344 5755 5350 5817
rect 5384 5755 5390 5817
rect 5344 5743 5390 5755
rect 6100 6536 6134 6552
rect 6100 6463 6134 6472
rect 6100 6390 6134 6396
rect 6100 6354 6134 6356
rect 6100 6317 6134 6320
rect 6100 6278 6134 6283
rect 6100 6202 6134 6210
rect 6100 6126 6134 6137
rect 6100 6050 6134 6064
rect 6100 5973 6134 5990
rect 6100 5896 6134 5916
rect 6100 5819 6134 5842
rect 6100 5752 6134 5768
rect 6484 6491 6490 6555
rect 6524 6491 6530 6555
rect 6484 6482 6530 6491
rect 6484 6423 6490 6482
rect 6524 6423 6530 6482
rect 6484 6409 6530 6423
rect 6484 6355 6490 6409
rect 6524 6355 6530 6409
rect 6484 6335 6530 6355
rect 6484 6287 6490 6335
rect 6524 6287 6530 6335
rect 6484 6261 6530 6287
rect 6484 6219 6490 6261
rect 6524 6219 6530 6261
rect 6484 6187 6530 6219
rect 6484 6151 6490 6187
rect 6524 6151 6530 6187
rect 6484 6117 6530 6151
rect 6484 6079 6490 6117
rect 6524 6079 6530 6117
rect 6484 6049 6530 6079
rect 6484 6005 6490 6049
rect 6524 6005 6530 6049
rect 6484 5981 6530 6005
rect 6484 5931 6490 5981
rect 6524 5931 6530 5981
rect 6484 5913 6530 5931
rect 6484 5857 6490 5913
rect 6524 5857 6530 5913
rect 6484 5845 6530 5857
rect 6484 5783 6490 5845
rect 6524 5783 6530 5845
rect 6484 5777 6530 5783
rect 5344 5685 5350 5743
rect 5384 5685 5390 5743
rect 5720 5708 5729 5742
rect 5788 5708 5804 5742
rect 3076 5615 3122 5632
rect 3076 5559 3082 5615
rect 3116 5559 3122 5615
rect 3076 5547 3122 5559
rect 3076 5486 3082 5547
rect 3116 5486 3122 5547
rect 3076 5479 3122 5486
rect 3076 5413 3082 5479
rect 3116 5413 3122 5479
rect 3076 5411 3122 5413
rect 3076 5377 3082 5411
rect 3116 5377 3122 5411
rect 3076 5374 3122 5377
rect 3076 5340 3082 5374
rect 3116 5340 3122 5374
rect 3076 5307 3122 5340
rect 5344 5669 5390 5685
rect 5344 5615 5350 5669
rect 5384 5615 5390 5669
rect 5344 5595 5390 5615
rect 5344 5545 5350 5595
rect 5384 5545 5390 5595
rect 5344 5521 5390 5545
rect 5344 5475 5350 5521
rect 5384 5475 5390 5521
rect 5344 5447 5390 5475
rect 5344 5405 5350 5447
rect 5384 5405 5390 5447
rect 5344 5373 5390 5405
rect 5344 5335 5350 5373
rect 5384 5335 5390 5373
rect 5344 5307 5390 5335
rect 6484 5675 6490 5777
rect 6524 5675 6530 5777
rect 6484 5669 6530 5675
rect 6484 5607 6490 5669
rect 6524 5607 6530 5669
rect 6484 5595 6530 5607
rect 6484 5539 6490 5595
rect 6524 5539 6530 5595
rect 6484 5521 6530 5539
rect 6484 5471 6490 5521
rect 6524 5471 6530 5521
rect 6484 5447 6530 5471
rect 6484 5403 6490 5447
rect 6524 5403 6530 5447
rect 6484 5373 6530 5403
rect 6484 5335 6490 5373
rect 6524 5335 6530 5373
rect 6484 5307 6530 5335
rect 3076 5301 3655 5307
rect 3880 5301 6530 5307
rect 3076 5267 3150 5301
rect 3188 5267 3218 5301
rect 3274 5267 3286 5301
rect 3320 5267 3326 5301
rect 3388 5267 3412 5301
rect 3456 5267 3490 5301
rect 3532 5267 3558 5301
rect 3617 5267 3626 5301
rect 3660 5267 3694 5301
rect 3728 5267 3762 5301
rect 3796 5267 3830 5301
rect 3864 5267 3898 5301
rect 3952 5267 3966 5301
rect 4026 5267 4034 5301
rect 4100 5267 4102 5301
rect 4136 5267 4140 5301
rect 4204 5267 4214 5301
rect 4272 5267 4288 5301
rect 4340 5267 4362 5301
rect 4408 5267 4436 5301
rect 4476 5267 4510 5301
rect 4544 5267 4578 5301
rect 4618 5267 4646 5301
rect 4692 5267 4714 5301
rect 4766 5267 4782 5301
rect 4840 5267 4850 5301
rect 4914 5267 4918 5301
rect 4952 5267 4954 5301
rect 5020 5267 5028 5301
rect 5088 5267 5102 5301
rect 5156 5267 5176 5301
rect 5224 5267 5249 5301
rect 5292 5267 5322 5301
rect 5360 5267 5394 5301
rect 5429 5267 5462 5301
rect 5502 5267 5530 5301
rect 5575 5267 5598 5301
rect 5648 5267 5666 5301
rect 5721 5267 5734 5301
rect 5794 5267 5802 5301
rect 5867 5267 5870 5301
rect 5904 5267 5906 5301
rect 5972 5267 5979 5301
rect 6040 5267 6052 5301
rect 6108 5267 6125 5301
rect 6176 5267 6198 5301
rect 6244 5267 6271 5301
rect 6312 5267 6344 5301
rect 6380 5267 6414 5301
rect 6451 5267 6530 5301
rect 3076 5261 3655 5267
rect 3880 5261 6530 5267
rect 6744 7708 6750 7761
rect 6784 7708 6790 7761
rect 6744 7693 6790 7708
rect 6744 7635 6750 7693
rect 6784 7635 6790 7693
rect 6744 7625 6790 7635
rect 6744 7562 6750 7625
rect 6784 7562 6790 7625
rect 6744 7557 6790 7562
rect 6744 7455 6750 7557
rect 6784 7455 6790 7557
rect 6744 7450 6790 7455
rect 6744 7387 6750 7450
rect 6784 7387 6790 7450
rect 6744 7377 6790 7387
rect 6744 7319 6750 7377
rect 6784 7319 6790 7377
rect 6744 7304 6790 7319
rect 6744 7251 6750 7304
rect 6784 7251 6790 7304
rect 6744 7231 6790 7251
rect 6744 7183 6750 7231
rect 6784 7183 6790 7231
rect 6744 7158 6790 7183
rect 6744 7115 6750 7158
rect 6784 7115 6790 7158
rect 6744 7085 6790 7115
rect 6744 7047 6750 7085
rect 6784 7047 6790 7085
rect 6744 7013 6790 7047
rect 6744 6978 6750 7013
rect 6784 6978 6790 7013
rect 6744 6945 6790 6978
rect 6744 6905 6750 6945
rect 6784 6905 6790 6945
rect 6744 6877 6790 6905
rect 6744 6832 6750 6877
rect 6784 6832 6790 6877
rect 6744 6809 6790 6832
rect 6744 6759 6750 6809
rect 6784 6759 6790 6809
rect 6744 6741 6790 6759
rect 6744 6686 6750 6741
rect 6784 6686 6790 6741
rect 6744 6673 6790 6686
rect 6744 6613 6750 6673
rect 6784 6613 6790 6673
rect 6744 6605 6790 6613
rect 6744 6540 6750 6605
rect 6784 6540 6790 6605
rect 6744 6537 6790 6540
rect 6744 6503 6750 6537
rect 6784 6503 6790 6537
rect 6744 6501 6790 6503
rect 6744 6435 6750 6501
rect 6784 6435 6790 6501
rect 6744 6428 6790 6435
rect 6744 6367 6750 6428
rect 6784 6367 6790 6428
rect 6744 6355 6790 6367
rect 6744 6299 6750 6355
rect 6784 6299 6790 6355
rect 6744 6282 6790 6299
rect 6744 6231 6750 6282
rect 6784 6231 6790 6282
rect 6744 6209 6790 6231
rect 6744 6163 6750 6209
rect 6784 6163 6790 6209
rect 6744 6136 6790 6163
rect 6744 6095 6750 6136
rect 6784 6095 6790 6136
rect 6744 6063 6790 6095
rect 6744 6027 6750 6063
rect 6784 6027 6790 6063
rect 6744 5993 6790 6027
rect 6744 5956 6750 5993
rect 6784 5956 6790 5993
rect 6744 5925 6790 5956
rect 6744 5883 6750 5925
rect 6784 5883 6790 5925
rect 6744 5857 6790 5883
rect 6744 5810 6750 5857
rect 6784 5810 6790 5857
rect 6744 5789 6790 5810
rect 6744 5737 6750 5789
rect 6784 5737 6790 5789
rect 6744 5721 6790 5737
rect 6744 5664 6750 5721
rect 6784 5664 6790 5721
rect 6744 5653 6790 5664
rect 6744 5591 6750 5653
rect 6784 5591 6790 5653
rect 6744 5585 6790 5591
rect 6744 5518 6750 5585
rect 6784 5518 6790 5585
rect 6744 5517 6790 5518
rect 6744 5483 6750 5517
rect 6784 5483 6790 5517
rect 6744 5479 6790 5483
rect 6744 5415 6750 5479
rect 6784 5415 6790 5479
rect 6744 5406 6790 5415
rect 6744 5347 6750 5406
rect 6784 5347 6790 5406
rect 6744 5333 6790 5347
rect 6744 5279 6750 5333
rect 6784 5279 6790 5333
rect 2796 5217 2842 5245
rect 2796 5183 2802 5217
rect 2836 5183 2842 5217
rect 2796 5145 2842 5183
rect 2796 5109 2802 5145
rect 2836 5109 2842 5145
rect 2796 5073 2842 5109
rect 2796 5039 2802 5073
rect 2836 5041 2842 5073
rect 6744 5260 6790 5279
rect 6744 5211 6750 5260
rect 6784 5211 6790 5260
rect 6744 5187 6790 5211
rect 6744 5143 6750 5187
rect 6784 5143 6790 5187
rect 6744 5113 6790 5143
rect 6744 5075 6750 5113
rect 6784 5075 6790 5113
rect 6744 5047 6790 5075
rect 3880 5041 6790 5047
rect 2836 5039 2870 5041
rect 2796 5007 2870 5039
rect 2933 5007 2938 5041
rect 2972 5007 2977 5041
rect 3040 5007 3056 5041
rect 3108 5007 3135 5041
rect 3176 5007 3210 5041
rect 3248 5007 3278 5041
rect 3327 5007 3346 5041
rect 3406 5007 3414 5041
rect 3448 5007 3451 5041
rect 3516 5007 3530 5041
rect 3584 5007 3609 5041
rect 3652 5007 3686 5041
rect 3720 5007 3754 5041
rect 3788 5007 3822 5041
rect 3856 5007 3890 5041
rect 3952 5007 3958 5041
rect 4025 5007 4026 5041
rect 4060 5007 4064 5041
rect 4128 5007 4137 5041
rect 4196 5007 4210 5041
rect 4264 5007 4283 5041
rect 4332 5007 4356 5041
rect 4400 5007 4429 5041
rect 4468 5007 4502 5041
rect 4536 5007 4570 5041
rect 4609 5007 4638 5041
rect 4682 5007 4706 5041
rect 4755 5007 4774 5041
rect 4828 5007 4842 5041
rect 4901 5007 4910 5041
rect 4974 5007 4978 5041
rect 5012 5007 5013 5041
rect 5080 5007 5086 5041
rect 5148 5007 5159 5041
rect 5216 5007 5232 5041
rect 5284 5007 5305 5041
rect 5352 5007 5378 5041
rect 5420 5007 5451 5041
rect 5488 5007 5522 5041
rect 5558 5007 5590 5041
rect 5631 5007 5658 5041
rect 5704 5007 5726 5041
rect 5776 5007 5794 5041
rect 5848 5007 5862 5041
rect 5920 5007 5930 5041
rect 5992 5007 5998 5041
rect 6064 5007 6066 5041
rect 6100 5007 6102 5041
rect 6168 5007 6174 5041
rect 6236 5007 6246 5041
rect 6304 5007 6318 5041
rect 6372 5007 6390 5041
rect 6440 5007 6462 5041
rect 6508 5007 6534 5041
rect 6576 5007 6606 5041
rect 6644 5007 6678 5041
rect 6712 5007 6790 5041
rect 2796 5001 2842 5007
rect 3880 5001 6790 5007
rect 8000 8062 8036 8096
rect 8000 7994 8036 8028
rect 8000 7990 8002 7994
rect 8034 7956 8036 7960
rect 8000 7926 8036 7956
rect 8000 7918 8002 7926
rect 8034 7884 8036 7892
rect 8000 7858 8036 7884
rect 8000 7846 8002 7858
rect 8034 7812 8036 7824
rect 8000 7790 8036 7812
rect 8000 7774 8002 7790
rect 8034 7740 8036 7756
rect 8000 7722 8036 7740
rect 8000 7702 8002 7722
rect 8034 7668 8036 7688
rect 8000 7654 8036 7668
rect 8000 7630 8002 7654
rect 8034 7596 8036 7620
rect 8000 7586 8036 7596
rect 8000 7558 8002 7586
rect 8034 7524 8036 7552
rect 8000 7518 8036 7524
rect 8000 7486 8002 7518
rect 8034 7452 8036 7484
rect 8000 7450 8036 7452
rect 8000 7416 8002 7450
rect 8000 7414 8036 7416
rect 8034 7382 8036 7414
rect 8000 7348 8002 7380
rect 8000 7342 8036 7348
rect 8034 7314 8036 7342
rect 8000 7280 8002 7308
rect 8000 7270 8036 7280
rect 8034 7246 8036 7270
rect 8000 7212 8002 7236
rect 8000 7198 8036 7212
rect 8034 7178 8036 7198
rect 8000 7144 8002 7164
rect 8000 7126 8036 7144
rect 8034 7110 8036 7126
rect 8000 7076 8002 7092
rect 8000 7054 8036 7076
rect 8034 7042 8036 7054
rect 8000 7008 8002 7020
rect 8000 6982 8036 7008
rect 8034 6974 8036 6982
rect 8000 6940 8002 6948
rect 8000 6910 8036 6940
rect 8034 6906 8036 6910
rect 8000 6872 8002 6876
rect 8000 6838 8036 6872
rect 8000 6770 8036 6804
rect 8000 6766 8002 6770
rect 8034 6732 8036 6736
rect 8000 6702 8036 6732
rect 8000 6694 8002 6702
rect 8034 6660 8036 6668
rect 8000 6634 8036 6660
rect 8000 6622 8002 6634
rect 8034 6588 8036 6600
rect 8000 6566 8036 6588
rect 8000 6550 8002 6566
rect 8034 6516 8036 6532
rect 8000 6498 8036 6516
rect 8000 6478 8002 6498
rect 8034 6444 8036 6464
rect 8000 6430 8036 6444
rect 8000 6406 8002 6430
rect 8034 6372 8036 6396
rect 8000 6362 8036 6372
rect 8000 6334 8002 6362
rect 8034 6300 8036 6328
rect 8000 6294 8036 6300
rect 8000 6262 8002 6294
rect 8034 6228 8036 6260
rect 8000 6226 8036 6228
rect 8000 6192 8002 6226
rect 8000 6190 8036 6192
rect 8034 6158 8036 6190
rect 8000 6124 8002 6156
rect 8000 6118 8036 6124
rect 8034 6090 8036 6118
rect 8000 6056 8002 6084
rect 8000 6046 8036 6056
rect 8034 6022 8036 6046
rect 8000 5988 8002 6012
rect 8000 5974 8036 5988
rect 8034 5954 8036 5974
rect 8000 5920 8002 5940
rect 8000 5902 8036 5920
rect 8034 5886 8036 5902
rect 8000 5852 8002 5868
rect 8000 5830 8036 5852
rect 8034 5818 8036 5830
rect 8000 5784 8002 5796
rect 8000 5758 8036 5784
rect 8034 5750 8036 5758
rect 8000 5716 8002 5724
rect 8000 5686 8036 5716
rect 8034 5682 8036 5686
rect 8000 5648 8002 5652
rect 8000 5614 8036 5648
rect 8000 5546 8036 5580
rect 8000 5542 8002 5546
rect 8034 5508 8036 5512
rect 8000 5478 8036 5508
rect 8000 5470 8002 5478
rect 8034 5436 8036 5444
rect 8000 5410 8036 5436
rect 8000 5398 8002 5410
rect 8034 5364 8036 5376
rect 8000 5342 8036 5364
rect 8000 5326 8002 5342
rect 8034 5292 8036 5308
rect 8000 5274 8036 5292
rect 8000 5254 8002 5274
rect 8034 5220 8036 5240
rect 8000 5206 8036 5220
rect 8000 5182 8002 5206
rect 8034 5148 8036 5172
rect 8000 5138 8036 5148
rect 8000 5110 8002 5138
rect 8034 5076 8036 5104
rect 8000 5070 8036 5076
rect 8000 5038 8002 5070
rect 8034 5004 8036 5036
rect 8000 5002 8036 5004
rect 8000 4968 8002 5002
rect 8000 4966 8036 4968
rect 8034 4934 8036 4966
rect 8000 4900 8002 4932
rect 8000 4894 8036 4900
rect 2802 4860 2803 4894
rect 2837 4860 2876 4894
rect 2921 4860 2949 4894
rect 2989 4860 3022 4894
rect 3057 4860 3091 4894
rect 3129 4860 3159 4894
rect 3202 4860 3227 4894
rect 3275 4860 3295 4894
rect 3348 4860 3363 4894
rect 3421 4860 3431 4894
rect 3495 4860 3499 4894
rect 3533 4860 3535 4894
rect 3601 4860 3609 4894
rect 3669 4860 3703 4894
rect 3737 4860 3771 4894
rect 3805 4860 3839 4894
rect 3873 4860 3892 4894
rect 3941 4860 3965 4894
rect 4009 4860 4038 4894
rect 4077 4860 4111 4894
rect 4145 4860 4179 4894
rect 4218 4860 4247 4894
rect 4291 4860 4315 4894
rect 4364 4860 4383 4894
rect 4437 4860 4451 4894
rect 4510 4860 4519 4894
rect 4583 4860 4587 4894
rect 4621 4860 4622 4894
rect 4689 4860 4695 4894
rect 4757 4860 4768 4894
rect 4825 4860 4841 4894
rect 4893 4860 4914 4894
rect 4961 4860 4987 4894
rect 5029 4860 5060 4894
rect 5097 4860 5131 4894
rect 5167 4860 5199 4894
rect 5239 4860 5267 4894
rect 5311 4860 5335 4894
rect 5383 4860 5403 4894
rect 5455 4860 5471 4894
rect 5527 4860 5539 4894
rect 5599 4860 5607 4894
rect 5671 4860 5675 4894
rect 5777 4860 5781 4894
rect 5845 4860 5853 4894
rect 5913 4860 5925 4894
rect 5981 4860 5997 4894
rect 6049 4860 6069 4894
rect 6117 4860 6141 4894
rect 6185 4860 6213 4894
rect 6253 4860 6285 4894
rect 6321 4860 6355 4894
rect 6391 4860 6423 4894
rect 6463 4860 6491 4894
rect 6535 4860 6559 4894
rect 6607 4860 6627 4894
rect 6679 4860 6695 4894
rect 6751 4860 6763 4894
rect 8034 4866 8036 4894
rect 8000 4832 8002 4860
rect 8000 4822 8036 4832
rect 8034 4798 8036 4822
rect 3039 4739 3055 4773
rect 3089 4739 3127 4773
rect 3166 4739 3199 4773
rect 3249 4739 3271 4773
rect 3332 4739 3343 4773
rect 3377 4739 3381 4773
rect 3449 4739 3463 4773
rect 3520 4739 3545 4773
rect 3591 4739 3607 4773
rect 8000 4764 8002 4788
rect 8000 4750 8036 4764
rect 8034 4730 8036 4750
rect 6464 4687 6509 4721
rect 6543 4687 6588 4721
rect 8000 4696 8002 4716
rect 2994 4561 3028 4599
rect 2994 4489 3028 4527
rect 2994 4417 3028 4455
rect 2994 4345 3028 4383
rect 2994 4273 3028 4311
rect 2994 4201 3028 4239
rect 2994 4129 3028 4167
rect 2994 4057 3028 4095
rect 2994 3985 3028 4023
rect 2994 3913 3028 3951
rect 2994 3841 3028 3879
rect 2994 3769 3028 3807
rect 2994 3697 3028 3735
rect 2994 3625 3028 3663
rect 2994 3553 3028 3591
rect 2994 3481 3028 3519
rect 2994 3409 3028 3447
rect 2994 3337 3028 3375
rect 3150 4561 3184 4599
rect 3150 4489 3184 4527
rect 3150 4417 3184 4455
rect 3150 4345 3184 4383
rect 3150 4273 3184 4311
rect 3150 4201 3184 4239
rect 3150 4129 3184 4167
rect 3150 4057 3184 4095
rect 3150 3985 3184 4023
rect 3150 3913 3184 3951
rect 3150 3841 3184 3879
rect 3150 3769 3184 3807
rect 3150 3697 3184 3735
rect 3150 3625 3184 3663
rect 3150 3553 3184 3591
rect 3150 3481 3184 3519
rect 3150 3409 3184 3447
rect 3150 3337 3184 3375
rect 3306 4561 3340 4599
rect 3306 4489 3340 4527
rect 3306 4417 3340 4455
rect 3306 4345 3340 4383
rect 3306 4273 3340 4311
rect 3306 4201 3340 4239
rect 3306 4129 3340 4167
rect 3306 4057 3340 4095
rect 3306 3985 3340 4023
rect 3306 3913 3340 3951
rect 3306 3841 3340 3879
rect 3306 3769 3340 3807
rect 3306 3697 3340 3735
rect 3306 3625 3340 3663
rect 3306 3553 3340 3591
rect 3306 3481 3340 3519
rect 3306 3409 3340 3447
rect 3306 3337 3340 3375
rect 3462 4561 3496 4599
rect 3462 4489 3496 4527
rect 3462 4417 3496 4455
rect 3462 4345 3496 4383
rect 3462 4273 3496 4311
rect 3462 4201 3496 4239
rect 3462 4129 3496 4167
rect 3462 4057 3496 4095
rect 3462 3985 3496 4023
rect 3462 3913 3496 3951
rect 3462 3841 3496 3879
rect 3462 3769 3496 3807
rect 3462 3697 3496 3735
rect 3462 3625 3496 3663
rect 3462 3553 3496 3591
rect 3462 3481 3496 3519
rect 3462 3409 3496 3447
rect 3462 3337 3496 3375
rect 3618 4561 3652 4599
rect 3618 4489 3652 4527
rect 4222 4537 4256 4645
rect 8000 4678 8036 4696
rect 5878 4537 5912 4645
rect 6336 4660 6370 4676
rect 6336 4589 6370 4626
rect 6336 4518 6370 4555
rect 3618 4417 3652 4455
rect 6336 4452 6370 4484
rect 4267 4409 4283 4443
rect 4317 4409 4334 4443
rect 4387 4409 4407 4443
rect 4457 4409 4480 4443
rect 4527 4409 4553 4443
rect 4597 4409 4626 4443
rect 4667 4409 4699 4443
rect 4737 4409 4772 4443
rect 4807 4409 4843 4443
rect 4879 4409 4913 4443
rect 4952 4409 4983 4443
rect 5024 4409 5053 4443
rect 5096 4409 5123 4443
rect 5168 4409 5193 4443
rect 5240 4409 5263 4443
rect 5312 4409 5333 4443
rect 5384 4409 5403 4443
rect 5456 4409 5472 4443
rect 5528 4409 5541 4443
rect 5600 4409 5610 4443
rect 5672 4409 5679 4443
rect 5713 4409 5748 4443
rect 5782 4409 5817 4443
rect 5851 4409 5867 4443
rect 3618 4345 3652 4383
rect 6336 4377 6370 4412
rect 3618 4273 3652 4311
rect 3618 4201 3652 4239
rect 4222 4205 4256 4313
rect 5878 4205 5912 4313
rect 6336 4302 6370 4340
rect 6336 4230 6370 4268
rect 8034 4662 8036 4678
rect 8000 4628 8002 4644
rect 8000 4606 8036 4628
rect 8034 4593 8036 4606
rect 8000 4559 8002 4572
rect 8000 4534 8036 4559
rect 8034 4524 8036 4534
rect 8000 4490 8002 4500
rect 8000 4462 8036 4490
rect 8034 4455 8036 4462
rect 8000 4421 8002 4428
rect 8000 4390 8036 4421
rect 8034 4386 8036 4390
rect 8000 4352 8002 4356
rect 8000 4318 8036 4352
rect 8034 4317 8036 4318
rect 8000 4283 8002 4284
rect 6464 4231 6509 4265
rect 6543 4231 6588 4265
rect 8000 4248 8036 4283
rect 8000 4246 8002 4248
rect 3618 4129 3652 4167
rect 3618 4057 3652 4095
rect 6336 4158 6370 4193
rect 6336 4086 6370 4117
rect 3618 3985 3652 4023
rect 4211 4015 4227 4049
rect 4261 4015 4293 4049
rect 4331 4015 4367 4049
rect 4401 4015 4437 4049
rect 4475 4015 4506 4049
rect 4549 4015 4575 4049
rect 4622 4015 4644 4049
rect 4695 4015 4713 4049
rect 4768 4015 4782 4049
rect 4841 4015 4851 4049
rect 4914 4015 4920 4049
rect 4987 4015 4989 4049
rect 5023 4015 5026 4049
rect 5092 4015 5099 4049
rect 5161 4015 5172 4049
rect 5230 4015 5245 4049
rect 5299 4015 5318 4049
rect 5368 4015 5391 4049
rect 5437 4015 5464 4049
rect 5506 4015 5537 4049
rect 5575 4015 5610 4049
rect 5644 4015 5679 4049
rect 5717 4015 5748 4049
rect 5790 4015 5817 4049
rect 5851 4015 5867 4049
rect 6336 4014 6370 4041
rect 3618 3913 3652 3951
rect 3618 3841 3652 3879
rect 3618 3769 3652 3807
rect 4166 3809 4200 3915
rect 5022 3880 5056 3921
rect 5022 3805 5056 3846
rect 5878 3882 5912 3921
rect 5878 3809 5912 3848
rect 6336 3942 6370 3965
rect 6336 3870 6370 3889
rect 6336 3820 6370 3836
rect 8034 4212 8036 4214
rect 8000 4179 8036 4212
rect 8000 4174 8002 4179
rect 8034 4140 8036 4145
rect 8000 4110 8036 4140
rect 8000 4101 8002 4110
rect 8034 4067 8036 4076
rect 8000 4041 8036 4067
rect 8000 4028 8002 4041
rect 8034 3994 8036 4007
rect 8000 3972 8036 3994
rect 8000 3955 8002 3972
rect 8034 3921 8036 3938
rect 8000 3903 8036 3921
rect 8000 3882 8002 3903
rect 8034 3848 8036 3869
rect 8000 3834 8036 3848
rect 8000 3809 8002 3834
rect 6464 3775 6509 3809
rect 6543 3775 6588 3809
rect 8034 3775 8036 3800
rect 3618 3697 3652 3735
rect 3618 3625 3652 3663
rect 3618 3553 3652 3591
rect 3618 3481 3652 3519
rect 3618 3409 3652 3447
rect 3618 3337 3652 3375
rect 8000 3765 8036 3775
rect 8000 3736 8002 3765
rect 8034 3702 8036 3731
rect 8000 3696 8036 3702
rect 8000 3663 8002 3696
rect 8034 3629 8036 3662
rect 8000 3627 8036 3629
rect 8000 3593 8002 3627
rect 8000 3590 8036 3593
rect 8034 3558 8036 3590
rect 8000 3524 8002 3556
rect 8000 3517 8036 3524
rect 8034 3489 8036 3517
rect 8000 3455 8002 3483
rect 8000 3444 8036 3455
rect 8034 3420 8036 3444
rect 8000 3386 8002 3410
rect 8000 3371 8036 3386
rect 8034 3351 8036 3371
rect 8000 3317 8002 3337
rect 8000 3298 8036 3317
rect 8034 3282 8036 3298
rect 8000 3248 8002 3264
rect 8000 3225 8036 3248
rect 8034 3213 8036 3225
rect 8000 3179 8002 3191
rect 2718 3124 2760 3158
rect 2812 3124 2836 3158
rect 2880 3124 2912 3158
rect 2948 3124 2982 3158
rect 3022 3124 3050 3158
rect 3098 3124 3118 3158
rect 3174 3124 3186 3158
rect 3250 3124 3254 3158
rect 3288 3124 3292 3158
rect 3356 3124 3368 3158
rect 3424 3124 3444 3158
rect 3492 3124 3520 3158
rect 3560 3124 3594 3158
rect 3629 3124 3662 3158
rect 3704 3124 3730 3158
rect 3779 3124 3798 3158
rect 3854 3124 3866 3158
rect 8000 3152 8036 3179
rect 8034 3144 8036 3152
rect 2481 2879 2488 2918
rect 2590 2879 2599 2918
rect 2481 2845 2487 2879
rect 2593 2845 2599 2879
rect 2481 2806 2488 2845
rect 2590 2806 2599 2845
rect 2481 2772 2487 2806
rect 2593 2772 2599 2806
rect 2481 2733 2488 2772
rect 2590 2733 2599 2772
rect 2481 2699 2487 2733
rect 2593 2699 2599 2733
rect 2481 2660 2488 2699
rect 2590 2660 2599 2699
rect 2481 2626 2487 2660
rect 2593 2626 2599 2660
rect 2481 2587 2488 2626
rect 2590 2587 2599 2626
rect 2481 2553 2487 2587
rect 2593 2553 2599 2587
rect 2481 2514 2488 2553
rect 2590 2514 2599 2553
rect 2481 2480 2487 2514
rect 2593 2480 2599 2514
rect 2481 2441 2488 2480
rect 2590 2441 2599 2480
rect 2481 2407 2487 2441
rect 2593 2407 2599 2441
rect 2481 2368 2488 2407
rect 2590 2368 2599 2407
rect 2481 2334 2487 2368
rect 2593 2334 2599 2368
rect 2481 2295 2488 2334
rect 2590 2295 2599 2334
rect 2481 2261 2487 2295
rect 2593 2261 2599 2295
rect 2481 2222 2488 2261
rect 2590 2222 2599 2261
rect 2481 2188 2487 2222
rect 2593 2188 2599 2222
rect 2481 2149 2488 2188
rect 2590 2149 2599 2188
rect 2481 2115 2487 2149
rect 2593 2115 2599 2149
rect 2481 2076 2488 2115
rect 2590 2076 2599 2115
rect 2481 2042 2487 2076
rect 2593 2042 2599 2076
rect 2481 2003 2488 2042
rect 2590 2003 2599 2042
rect 2481 1969 2487 2003
rect 2593 1969 2599 2003
rect 2481 1930 2488 1969
rect 2590 1930 2599 1969
rect 2481 1896 2487 1930
rect 2593 1896 2599 1930
rect 2481 1857 2488 1896
rect 2590 1857 2599 1896
rect 2481 1823 2487 1857
rect 2593 1823 2599 1857
rect 2481 1784 2488 1823
rect 2590 1784 2599 1823
rect 2481 1750 2487 1784
rect 2593 1750 2599 1784
rect 2481 1711 2488 1750
rect 2590 1711 2599 1750
rect 2481 1677 2487 1711
rect 2593 1677 2599 1711
rect 2481 1638 2488 1677
rect 2590 1638 2599 1677
rect 2481 1604 2487 1638
rect 2593 1604 2599 1638
rect 2481 1565 2488 1604
rect 2590 1565 2599 1604
rect 2481 1531 2487 1565
rect 2593 1531 2599 1565
rect 2481 1492 2488 1531
rect 2590 1492 2599 1531
rect 2481 1458 2487 1492
rect 2593 1458 2599 1492
rect 2481 1419 2488 1458
rect 2590 1419 2599 1458
rect 2481 1385 2487 1419
rect 2593 1385 2599 1419
rect 2481 1346 2488 1385
rect 2590 1346 2599 1385
rect 2481 1312 2487 1346
rect 2593 1312 2599 1346
rect 2481 1273 2488 1312
rect 2590 1273 2599 1312
rect 2481 1239 2487 1273
rect 2593 1239 2599 1273
rect 2481 1200 2488 1239
rect 2590 1200 2599 1239
rect 2481 1166 2487 1200
rect 2593 1166 2599 1200
rect 2481 1127 2488 1166
rect 2590 1127 2599 1166
rect 2481 1093 2487 1127
rect 2593 1093 2599 1127
rect 2481 1054 2488 1093
rect 2590 1054 2599 1093
rect 2481 1020 2487 1054
rect 2593 1020 2599 1054
rect 2481 981 2488 1020
rect 2590 981 2599 1020
rect 2481 947 2487 981
rect 2593 947 2599 981
rect 2481 908 2488 947
rect 2590 908 2599 947
rect 2481 874 2487 908
rect 2593 874 2599 908
rect 2481 835 2488 874
rect 2590 835 2599 874
rect 2481 801 2487 835
rect 2593 801 2599 835
rect 2481 762 2488 801
rect 2590 762 2599 801
rect 2481 728 2487 762
rect 2593 728 2599 762
rect 2481 689 2488 728
rect 2590 689 2599 728
rect 2481 655 2487 689
rect 2593 655 2599 689
rect 2481 616 2488 655
rect 2590 616 2599 655
rect 2481 582 2487 616
rect 2593 582 2599 616
rect 2481 543 2488 582
rect 2590 543 2599 582
rect 2481 509 2487 543
rect 2593 509 2599 543
rect 2481 470 2488 509
rect 2590 470 2599 509
rect 2481 436 2487 470
rect 2593 436 2599 470
rect 2481 398 2488 436
rect 374 232 476 344
rect 408 198 442 232
rect 374 164 476 198
rect 408 142 476 164
rect 408 130 442 142
rect 374 40 442 130
rect 2448 108 2488 142
rect 2590 398 2599 436
rect 8000 3110 8002 3118
rect 8000 3079 8036 3110
rect 8034 3075 8036 3079
rect 8000 3041 8002 3045
rect 8000 3006 8036 3041
rect 8000 2937 8036 2972
rect 8000 2933 8002 2937
rect 8034 2899 8036 2903
rect 8000 2868 8036 2899
rect 8000 2860 8002 2868
rect 8034 2826 8036 2834
rect 8000 2799 8036 2826
rect 8000 2787 8002 2799
rect 8034 2753 8036 2765
rect 8000 2730 8036 2753
rect 8000 2714 8002 2730
rect 8034 2680 8036 2696
rect 8000 2661 8036 2680
rect 8000 2641 8002 2661
rect 8034 2607 8036 2627
rect 8000 2592 8036 2607
rect 8000 2568 8002 2592
rect 8034 2534 8036 2558
rect 8000 2523 8036 2534
rect 8000 2495 8002 2523
rect 8034 2461 8036 2489
rect 8000 2454 8036 2461
rect 8000 2422 8002 2454
rect 8034 2388 8036 2420
rect 8000 2385 8036 2388
rect 8000 2351 8002 2385
rect 8000 2349 8036 2351
rect 8034 2316 8036 2349
rect 8000 2282 8002 2315
rect 8000 2276 8036 2282
rect 8034 2247 8036 2276
rect 8000 2213 8002 2242
rect 8000 2203 8036 2213
rect 8034 2178 8036 2203
rect 8000 2144 8002 2169
rect 8000 2130 8036 2144
rect 8034 2109 8036 2130
rect 8000 2075 8002 2096
rect 8000 2057 8036 2075
rect 8034 2040 8036 2057
rect 8000 2006 8002 2023
rect 8000 1984 8036 2006
rect 8034 1971 8036 1984
rect 8000 1937 8002 1950
rect 8000 1911 8036 1937
rect 8034 1902 8036 1911
rect 8000 1868 8002 1877
rect 8000 1838 8036 1868
rect 8034 1833 8036 1838
rect 8000 1799 8002 1804
rect 8000 1765 8036 1799
rect 8034 1764 8036 1765
rect 8000 1730 8002 1731
rect 8000 1695 8036 1730
rect 8000 1692 8002 1695
rect 8034 1658 8036 1661
rect 8000 1626 8036 1658
rect 8000 1619 8002 1626
rect 8034 1585 8036 1592
rect 8000 1557 8036 1585
rect 8000 1546 8002 1557
rect 8034 1512 8036 1523
rect 8000 1488 8036 1512
rect 8000 1473 8002 1488
rect 8034 1439 8036 1454
rect 8000 1419 8036 1439
rect 8000 1400 8002 1419
rect 8034 1366 8036 1385
rect 8000 1350 8036 1366
rect 8000 1327 8002 1350
rect 8034 1293 8036 1316
rect 8000 1281 8036 1293
rect 8000 1254 8002 1281
rect 8034 1220 8036 1247
rect 8000 1212 8036 1220
rect 8000 1181 8002 1212
rect 8034 1147 8036 1178
rect 8000 1143 8036 1147
rect 8000 1109 8002 1143
rect 8000 1108 8036 1109
rect 8034 1074 8036 1108
rect 8000 1040 8002 1074
rect 8000 1035 8036 1040
rect 8034 1005 8036 1035
rect 8000 971 8002 1001
rect 8000 962 8036 971
rect 8034 936 8036 962
rect 8000 902 8002 928
rect 8000 889 8036 902
rect 8034 867 8036 889
rect 8000 833 8002 855
rect 8000 816 8036 833
rect 8034 798 8036 816
rect 8000 764 8002 782
rect 8000 743 8036 764
rect 8034 729 8036 743
rect 8000 695 8002 709
rect 8000 670 8036 695
rect 8034 660 8036 670
rect 8000 626 8002 636
rect 8000 597 8036 626
rect 8034 591 8036 597
rect 8000 557 8002 563
rect 8000 524 8036 557
rect 8034 522 8036 524
rect 8000 488 8002 490
rect 8000 453 8036 488
rect 8000 451 8002 453
rect 8034 417 8036 419
rect 8000 384 8036 417
rect 9746 39495 9752 39546
rect 9786 39495 9792 39546
rect 9746 39478 9792 39495
rect 10593 39679 10631 39713
rect 10559 39640 10665 39679
rect 10593 39606 10631 39640
rect 10559 39567 10665 39606
rect 10593 39533 10631 39567
rect 10559 39487 10665 39533
rect 9746 39423 9752 39478
rect 9786 39423 9792 39478
rect 9746 39410 9792 39423
rect 9746 39351 9752 39410
rect 9786 39351 9792 39410
rect 9746 39342 9792 39351
rect 9746 39279 9752 39342
rect 9786 39279 9792 39342
rect 9746 39274 9792 39279
rect 9746 39207 9752 39274
rect 9786 39207 9792 39274
rect 9746 39206 9792 39207
rect 9746 39172 9752 39206
rect 9786 39172 9792 39206
rect 9746 39169 9792 39172
rect 9746 39104 9752 39169
rect 9786 39104 9792 39169
rect 9746 39097 9792 39104
rect 9746 39036 9752 39097
rect 9786 39036 9792 39097
rect 9746 39025 9792 39036
rect 9746 38968 9752 39025
rect 9786 38968 9792 39025
rect 9746 38953 9792 38968
rect 9746 38900 9752 38953
rect 9786 38900 9792 38953
rect 9746 38881 9792 38900
rect 9746 38832 9752 38881
rect 9786 38832 9792 38881
rect 9746 38809 9792 38832
rect 9746 38764 9752 38809
rect 9786 38764 9792 38809
rect 9746 38737 9792 38764
rect 9746 38696 9752 38737
rect 9786 38696 9792 38737
rect 9746 38665 9792 38696
rect 9746 38628 9752 38665
rect 9786 38628 9792 38665
rect 9746 38594 9792 38628
rect 9746 38559 9752 38594
rect 9786 38559 9792 38594
rect 9746 38526 9792 38559
rect 9746 38487 9752 38526
rect 9786 38487 9792 38526
rect 9746 38458 9792 38487
rect 9746 38415 9752 38458
rect 9786 38415 9792 38458
rect 9746 38390 9792 38415
rect 9746 38343 9752 38390
rect 9786 38343 9792 38390
rect 9746 38322 9792 38343
rect 9746 38271 9752 38322
rect 9786 38271 9792 38322
rect 9746 38254 9792 38271
rect 9746 38199 9752 38254
rect 9786 38199 9792 38254
rect 9746 38186 9792 38199
rect 9746 38127 9752 38186
rect 9786 38127 9792 38186
rect 9746 38118 9792 38127
rect 9746 38055 9752 38118
rect 9786 38055 9792 38118
rect 9746 38050 9792 38055
rect 9746 37983 9752 38050
rect 9786 37983 9792 38050
rect 9746 37982 9792 37983
rect 9746 37948 9752 37982
rect 9786 37948 9792 37982
rect 9746 37945 9792 37948
rect 9746 37880 9752 37945
rect 9786 37880 9792 37945
rect 9746 37873 9792 37880
rect 9746 37812 9752 37873
rect 9786 37812 9792 37873
rect 9746 37801 9792 37812
rect 9746 37744 9752 37801
rect 9786 37744 9792 37801
rect 9746 37729 9792 37744
rect 9746 37676 9752 37729
rect 9786 37676 9792 37729
rect 9746 37657 9792 37676
rect 9746 37608 9752 37657
rect 9786 37608 9792 37657
rect 9746 37585 9792 37608
rect 9746 37540 9752 37585
rect 9786 37540 9792 37585
rect 9746 37513 9792 37540
rect 9746 37472 9752 37513
rect 9786 37472 9792 37513
rect 9746 37441 9792 37472
rect 9746 37404 9752 37441
rect 9786 37404 9792 37441
rect 9746 37370 9792 37404
rect 9746 37335 9752 37370
rect 9786 37335 9792 37370
rect 9746 37302 9792 37335
rect 9746 37263 9752 37302
rect 9786 37263 9792 37302
rect 9746 37234 9792 37263
rect 9746 37191 9752 37234
rect 9786 37191 9792 37234
rect 9746 37166 9792 37191
rect 9746 37119 9752 37166
rect 9786 37119 9792 37166
rect 9746 37098 9792 37119
rect 9746 37047 9752 37098
rect 9786 37047 9792 37098
rect 9746 37030 9792 37047
rect 9746 36975 9752 37030
rect 9786 36975 9792 37030
rect 9746 36962 9792 36975
rect 9746 36903 9752 36962
rect 9786 36903 9792 36962
rect 9746 36894 9792 36903
rect 9746 36831 9752 36894
rect 9786 36831 9792 36894
rect 9746 36826 9792 36831
rect 9746 36759 9752 36826
rect 9786 36759 9792 36826
rect 9746 36758 9792 36759
rect 9746 36724 9752 36758
rect 9786 36724 9792 36758
rect 9746 36721 9792 36724
rect 9746 36656 9752 36721
rect 9786 36656 9792 36721
rect 9746 36649 9792 36656
rect 9746 36588 9752 36649
rect 9786 36588 9792 36649
rect 9746 36577 9792 36588
rect 9746 36520 9752 36577
rect 9786 36520 9792 36577
rect 9746 36505 9792 36520
rect 9746 36452 9752 36505
rect 9786 36452 9792 36505
rect 9746 36433 9792 36452
rect 9746 36384 9752 36433
rect 9786 36384 9792 36433
rect 9746 36361 9792 36384
rect 9746 36316 9752 36361
rect 9786 36316 9792 36361
rect 9746 36289 9792 36316
rect 9746 36248 9752 36289
rect 9786 36248 9792 36289
rect 9746 36217 9792 36248
rect 9746 36180 9752 36217
rect 9786 36180 9792 36217
rect 9746 36146 9792 36180
rect 9746 36111 9752 36146
rect 9786 36111 9792 36146
rect 9746 36078 9792 36111
rect 9746 36039 9752 36078
rect 9786 36039 9792 36078
rect 9746 36010 9792 36039
rect 9746 35967 9752 36010
rect 9786 35967 9792 36010
rect 9746 35942 9792 35967
rect 9746 35895 9752 35942
rect 9786 35895 9792 35942
rect 9746 35874 9792 35895
rect 9746 35823 9752 35874
rect 9786 35823 9792 35874
rect 9746 35806 9792 35823
rect 9746 35751 9752 35806
rect 9786 35751 9792 35806
rect 9746 35738 9792 35751
rect 9746 35679 9752 35738
rect 9786 35679 9792 35738
rect 9746 35670 9792 35679
rect 9746 35607 9752 35670
rect 9786 35607 9792 35670
rect 9746 35602 9792 35607
rect 9746 35535 9752 35602
rect 9786 35535 9792 35602
rect 9746 35534 9792 35535
rect 9746 35500 9752 35534
rect 9786 35500 9792 35534
rect 9746 35497 9792 35500
rect 9746 35432 9752 35497
rect 9786 35432 9792 35497
rect 9746 35425 9792 35432
rect 9746 35364 9752 35425
rect 9786 35364 9792 35425
rect 9746 35353 9792 35364
rect 9746 35296 9752 35353
rect 9786 35296 9792 35353
rect 9746 35281 9792 35296
rect 9746 35228 9752 35281
rect 9786 35228 9792 35281
rect 9746 35209 9792 35228
rect 9746 35160 9752 35209
rect 9786 35160 9792 35209
rect 9746 35137 9792 35160
rect 9746 35092 9752 35137
rect 9786 35092 9792 35137
rect 9746 35065 9792 35092
rect 9746 35024 9752 35065
rect 9786 35024 9792 35065
rect 9746 34993 9792 35024
rect 9746 34956 9752 34993
rect 9786 34956 9792 34993
rect 9746 34922 9792 34956
rect 9746 34887 9752 34922
rect 9786 34887 9792 34922
rect 9746 34854 9792 34887
rect 9746 34815 9752 34854
rect 9786 34815 9792 34854
rect 9746 34786 9792 34815
rect 9746 34743 9752 34786
rect 9786 34743 9792 34786
rect 9746 34718 9792 34743
rect 9746 34671 9752 34718
rect 9786 34671 9792 34718
rect 9746 34650 9792 34671
rect 9746 34599 9752 34650
rect 9786 34599 9792 34650
rect 9746 34582 9792 34599
rect 9746 34527 9752 34582
rect 9786 34527 9792 34582
rect 9746 34514 9792 34527
rect 9746 34455 9752 34514
rect 9786 34455 9792 34514
rect 9746 34446 9792 34455
rect 9746 34383 9752 34446
rect 9786 34383 9792 34446
rect 9746 34378 9792 34383
rect 9746 34311 9752 34378
rect 9786 34311 9792 34378
rect 9746 34310 9792 34311
rect 9746 34276 9752 34310
rect 9786 34276 9792 34310
rect 9746 34273 9792 34276
rect 9746 34208 9752 34273
rect 9786 34208 9792 34273
rect 9746 34201 9792 34208
rect 9746 34140 9752 34201
rect 9786 34140 9792 34201
rect 9746 34129 9792 34140
rect 9746 34072 9752 34129
rect 9786 34072 9792 34129
rect 9746 34057 9792 34072
rect 9746 34004 9752 34057
rect 9786 34004 9792 34057
rect 9746 33985 9792 34004
rect 9746 33936 9752 33985
rect 9786 33936 9792 33985
rect 9746 33913 9792 33936
rect 9746 33868 9752 33913
rect 9786 33868 9792 33913
rect 9746 33841 9792 33868
rect 9746 33800 9752 33841
rect 9786 33800 9792 33841
rect 9746 33769 9792 33800
rect 9746 33732 9752 33769
rect 9786 33732 9792 33769
rect 9746 33698 9792 33732
rect 9746 33663 9752 33698
rect 9786 33663 9792 33698
rect 9746 33630 9792 33663
rect 9746 33591 9752 33630
rect 9786 33591 9792 33630
rect 9746 33562 9792 33591
rect 9746 33519 9752 33562
rect 9786 33519 9792 33562
rect 9746 33494 9792 33519
rect 9746 33447 9752 33494
rect 9786 33447 9792 33494
rect 9746 33426 9792 33447
rect 9746 33375 9752 33426
rect 9786 33375 9792 33426
rect 9746 33358 9792 33375
rect 9746 33303 9752 33358
rect 9786 33303 9792 33358
rect 9746 33290 9792 33303
rect 9746 33231 9752 33290
rect 9786 33231 9792 33290
rect 9746 33222 9792 33231
rect 9746 33159 9752 33222
rect 9786 33159 9792 33222
rect 9746 33154 9792 33159
rect 9746 33087 9752 33154
rect 9786 33087 9792 33154
rect 9746 33086 9792 33087
rect 9746 33052 9752 33086
rect 9786 33052 9792 33086
rect 9746 33049 9792 33052
rect 9746 32984 9752 33049
rect 9786 32984 9792 33049
rect 9746 32977 9792 32984
rect 9746 32916 9752 32977
rect 9786 32916 9792 32977
rect 9746 32905 9792 32916
rect 9746 32848 9752 32905
rect 9786 32848 9792 32905
rect 9746 32833 9792 32848
rect 9746 32780 9752 32833
rect 9786 32780 9792 32833
rect 9746 32761 9792 32780
rect 9746 32712 9752 32761
rect 9786 32712 9792 32761
rect 9746 32689 9792 32712
rect 9746 32644 9752 32689
rect 9786 32644 9792 32689
rect 9746 32617 9792 32644
rect 9746 32576 9752 32617
rect 9786 32576 9792 32617
rect 9746 32545 9792 32576
rect 9746 32508 9752 32545
rect 9786 32508 9792 32545
rect 9746 32474 9792 32508
rect 9746 32439 9752 32474
rect 9786 32439 9792 32474
rect 9746 32406 9792 32439
rect 9746 32367 9752 32406
rect 9786 32367 9792 32406
rect 9746 32338 9792 32367
rect 9746 32295 9752 32338
rect 9786 32295 9792 32338
rect 9746 32270 9792 32295
rect 9746 32223 9752 32270
rect 9786 32223 9792 32270
rect 9746 32202 9792 32223
rect 9746 32151 9752 32202
rect 9786 32151 9792 32202
rect 9746 32134 9792 32151
rect 9746 32079 9752 32134
rect 9786 32079 9792 32134
rect 9746 32066 9792 32079
rect 9746 32007 9752 32066
rect 9786 32007 9792 32066
rect 9746 31998 9792 32007
rect 9746 31935 9752 31998
rect 9786 31935 9792 31998
rect 9746 31930 9792 31935
rect 9746 31863 9752 31930
rect 9786 31863 9792 31930
rect 9746 31862 9792 31863
rect 9746 31828 9752 31862
rect 9786 31828 9792 31862
rect 9746 31825 9792 31828
rect 9746 31760 9752 31825
rect 9786 31760 9792 31825
rect 9746 31753 9792 31760
rect 9746 31692 9752 31753
rect 9786 31692 9792 31753
rect 9746 31681 9792 31692
rect 9746 31624 9752 31681
rect 9786 31624 9792 31681
rect 9746 31609 9792 31624
rect 9746 31556 9752 31609
rect 9786 31556 9792 31609
rect 9746 31537 9792 31556
rect 9746 31488 9752 31537
rect 9786 31488 9792 31537
rect 9746 31465 9792 31488
rect 9746 31420 9752 31465
rect 9786 31420 9792 31465
rect 9746 31393 9792 31420
rect 9746 31352 9752 31393
rect 9786 31352 9792 31393
rect 9746 31321 9792 31352
rect 9746 31284 9752 31321
rect 9786 31284 9792 31321
rect 9746 31250 9792 31284
rect 9746 31215 9752 31250
rect 9786 31215 9792 31250
rect 9746 31182 9792 31215
rect 9746 31143 9752 31182
rect 9786 31143 9792 31182
rect 9746 31114 9792 31143
rect 9746 31071 9752 31114
rect 9786 31071 9792 31114
rect 9746 31046 9792 31071
rect 9746 30999 9752 31046
rect 9786 30999 9792 31046
rect 9746 30978 9792 30999
rect 9746 30927 9752 30978
rect 9786 30927 9792 30978
rect 9746 30910 9792 30927
rect 9746 30855 9752 30910
rect 9786 30855 9792 30910
rect 9746 30842 9792 30855
rect 9746 30783 9752 30842
rect 9786 30783 9792 30842
rect 9746 30774 9792 30783
rect 9746 30711 9752 30774
rect 9786 30711 9792 30774
rect 9746 30706 9792 30711
rect 9746 30639 9752 30706
rect 9786 30639 9792 30706
rect 9746 30638 9792 30639
rect 9746 30604 9752 30638
rect 9786 30604 9792 30638
rect 9746 30601 9792 30604
rect 9746 30536 9752 30601
rect 9786 30536 9792 30601
rect 9746 30529 9792 30536
rect 9746 30468 9752 30529
rect 9786 30468 9792 30529
rect 9746 30457 9792 30468
rect 9746 30400 9752 30457
rect 9786 30400 9792 30457
rect 9746 30385 9792 30400
rect 9746 30332 9752 30385
rect 9786 30332 9792 30385
rect 9746 30313 9792 30332
rect 9746 30264 9752 30313
rect 9786 30264 9792 30313
rect 9746 30241 9792 30264
rect 9746 30196 9752 30241
rect 9786 30196 9792 30241
rect 9746 30169 9792 30196
rect 9746 30128 9752 30169
rect 9786 30128 9792 30169
rect 9746 30097 9792 30128
rect 9746 30060 9752 30097
rect 9786 30060 9792 30097
rect 9746 30026 9792 30060
rect 9746 29991 9752 30026
rect 9786 29991 9792 30026
rect 9746 29958 9792 29991
rect 9746 29919 9752 29958
rect 9786 29919 9792 29958
rect 9746 29890 9792 29919
rect 9746 29847 9752 29890
rect 9786 29847 9792 29890
rect 9746 29822 9792 29847
rect 9746 29775 9752 29822
rect 9786 29775 9792 29822
rect 9746 29754 9792 29775
rect 9746 29703 9752 29754
rect 9786 29703 9792 29754
rect 9746 29686 9792 29703
rect 9746 29631 9752 29686
rect 9786 29631 9792 29686
rect 9746 29618 9792 29631
rect 9746 29559 9752 29618
rect 9786 29559 9792 29618
rect 9746 29550 9792 29559
rect 9746 29487 9752 29550
rect 9786 29487 9792 29550
rect 9746 29482 9792 29487
rect 9746 29415 9752 29482
rect 9786 29415 9792 29482
rect 9746 29414 9792 29415
rect 9746 29380 9752 29414
rect 9786 29380 9792 29414
rect 9746 29377 9792 29380
rect 9746 29312 9752 29377
rect 9786 29312 9792 29377
rect 9746 29305 9792 29312
rect 9746 29244 9752 29305
rect 9786 29244 9792 29305
rect 9746 29233 9792 29244
rect 9746 29176 9752 29233
rect 9786 29176 9792 29233
rect 9746 29161 9792 29176
rect 9746 29108 9752 29161
rect 9786 29108 9792 29161
rect 9746 29089 9792 29108
rect 9746 29040 9752 29089
rect 9786 29040 9792 29089
rect 9746 29017 9792 29040
rect 9746 28972 9752 29017
rect 9786 28972 9792 29017
rect 9746 28945 9792 28972
rect 9746 28904 9752 28945
rect 9786 28904 9792 28945
rect 9746 28873 9792 28904
rect 9746 28836 9752 28873
rect 9786 28836 9792 28873
rect 9746 28802 9792 28836
rect 9746 28767 9752 28802
rect 9786 28767 9792 28802
rect 9746 28734 9792 28767
rect 9746 28695 9752 28734
rect 9786 28695 9792 28734
rect 9746 28666 9792 28695
rect 9746 28623 9752 28666
rect 9786 28623 9792 28666
rect 9746 28598 9792 28623
rect 9746 28551 9752 28598
rect 9786 28551 9792 28598
rect 9746 28530 9792 28551
rect 9746 28479 9752 28530
rect 9786 28479 9792 28530
rect 9746 28462 9792 28479
rect 9746 28407 9752 28462
rect 9786 28407 9792 28462
rect 9746 28394 9792 28407
rect 9746 28335 9752 28394
rect 9786 28335 9792 28394
rect 9746 28326 9792 28335
rect 9746 28263 9752 28326
rect 9786 28263 9792 28326
rect 9746 28258 9792 28263
rect 9746 28191 9752 28258
rect 9786 28191 9792 28258
rect 9746 28190 9792 28191
rect 9746 28156 9752 28190
rect 9786 28156 9792 28190
rect 9746 28153 9792 28156
rect 9746 28088 9752 28153
rect 9786 28088 9792 28153
rect 9746 28081 9792 28088
rect 9746 28020 9752 28081
rect 9786 28020 9792 28081
rect 9746 28009 9792 28020
rect 9746 27952 9752 28009
rect 9786 27952 9792 28009
rect 9746 27937 9792 27952
rect 9746 27884 9752 27937
rect 9786 27884 9792 27937
rect 9746 27865 9792 27884
rect 9746 27816 9752 27865
rect 9786 27816 9792 27865
rect 9746 27793 9792 27816
rect 9746 27748 9752 27793
rect 9786 27748 9792 27793
rect 9746 27721 9792 27748
rect 9746 27680 9752 27721
rect 9786 27680 9792 27721
rect 9746 27649 9792 27680
rect 9746 27612 9752 27649
rect 9786 27612 9792 27649
rect 9746 27578 9792 27612
rect 9746 27543 9752 27578
rect 9786 27543 9792 27578
rect 9746 27510 9792 27543
rect 9746 27471 9752 27510
rect 9786 27471 9792 27510
rect 9746 27442 9792 27471
rect 9746 27399 9752 27442
rect 9786 27399 9792 27442
rect 9746 27374 9792 27399
rect 9746 27327 9752 27374
rect 9786 27327 9792 27374
rect 9746 27306 9792 27327
rect 9746 27255 9752 27306
rect 9786 27255 9792 27306
rect 9746 27238 9792 27255
rect 9746 27183 9752 27238
rect 9786 27183 9792 27238
rect 9746 27170 9792 27183
rect 9746 27111 9752 27170
rect 9786 27111 9792 27170
rect 9746 27102 9792 27111
rect 9746 27039 9752 27102
rect 9786 27039 9792 27102
rect 9746 27034 9792 27039
rect 9746 26967 9752 27034
rect 9786 26967 9792 27034
rect 9746 26966 9792 26967
rect 9746 26932 9752 26966
rect 9786 26932 9792 26966
rect 9746 26929 9792 26932
rect 9746 26864 9752 26929
rect 9786 26864 9792 26929
rect 9746 26857 9792 26864
rect 9746 26796 9752 26857
rect 9786 26796 9792 26857
rect 9746 26785 9792 26796
rect 9746 26728 9752 26785
rect 9786 26728 9792 26785
rect 9746 26713 9792 26728
rect 9746 26660 9752 26713
rect 9786 26660 9792 26713
rect 9746 26641 9792 26660
rect 9746 26592 9752 26641
rect 9786 26592 9792 26641
rect 9746 26569 9792 26592
rect 9746 26524 9752 26569
rect 9786 26524 9792 26569
rect 9746 26497 9792 26524
rect 9746 26456 9752 26497
rect 9786 26456 9792 26497
rect 9746 26425 9792 26456
rect 9746 26388 9752 26425
rect 9786 26388 9792 26425
rect 9746 26354 9792 26388
rect 9746 26319 9752 26354
rect 9786 26319 9792 26354
rect 9746 26286 9792 26319
rect 9746 26247 9752 26286
rect 9786 26247 9792 26286
rect 9746 26218 9792 26247
rect 9746 26175 9752 26218
rect 9786 26175 9792 26218
rect 9746 26150 9792 26175
rect 9746 26103 9752 26150
rect 9786 26103 9792 26150
rect 9746 26082 9792 26103
rect 9746 26031 9752 26082
rect 9786 26031 9792 26082
rect 9746 26014 9792 26031
rect 9746 25959 9752 26014
rect 9786 25959 9792 26014
rect 9746 25946 9792 25959
rect 9746 25887 9752 25946
rect 9786 25887 9792 25946
rect 9746 25878 9792 25887
rect 9746 25815 9752 25878
rect 9786 25815 9792 25878
rect 9746 25810 9792 25815
rect 9746 25743 9752 25810
rect 9786 25743 9792 25810
rect 9746 25742 9792 25743
rect 9746 25708 9752 25742
rect 9786 25708 9792 25742
rect 9746 25705 9792 25708
rect 9746 25640 9752 25705
rect 9786 25640 9792 25705
rect 9746 25633 9792 25640
rect 9746 25572 9752 25633
rect 9786 25572 9792 25633
rect 9746 25561 9792 25572
rect 9746 25504 9752 25561
rect 9786 25504 9792 25561
rect 9746 25489 9792 25504
rect 9746 25436 9752 25489
rect 9786 25436 9792 25489
rect 9746 25417 9792 25436
rect 9746 25368 9752 25417
rect 9786 25368 9792 25417
rect 9746 25345 9792 25368
rect 9746 25300 9752 25345
rect 9786 25300 9792 25345
rect 9746 25273 9792 25300
rect 9746 25232 9752 25273
rect 9786 25232 9792 25273
rect 9746 25201 9792 25232
rect 9746 25164 9752 25201
rect 9786 25164 9792 25201
rect 9746 25130 9792 25164
rect 9746 25095 9752 25130
rect 9786 25095 9792 25130
rect 9746 25062 9792 25095
rect 9746 25023 9752 25062
rect 9786 25023 9792 25062
rect 9746 24994 9792 25023
rect 9746 24951 9752 24994
rect 9786 24951 9792 24994
rect 9746 24926 9792 24951
rect 9746 24879 9752 24926
rect 9786 24879 9792 24926
rect 9746 24858 9792 24879
rect 9746 24807 9752 24858
rect 9786 24807 9792 24858
rect 9746 24790 9792 24807
rect 9746 24735 9752 24790
rect 9786 24735 9792 24790
rect 9746 24722 9792 24735
rect 9746 24663 9752 24722
rect 9786 24663 9792 24722
rect 9746 24654 9792 24663
rect 9746 24591 9752 24654
rect 9786 24591 9792 24654
rect 9746 24586 9792 24591
rect 9746 24519 9752 24586
rect 9786 24519 9792 24586
rect 9746 24518 9792 24519
rect 9746 24484 9752 24518
rect 9786 24484 9792 24518
rect 9746 24481 9792 24484
rect 9746 24416 9752 24481
rect 9786 24416 9792 24481
rect 9746 24409 9792 24416
rect 9746 24348 9752 24409
rect 9786 24348 9792 24409
rect 9746 24337 9792 24348
rect 9746 24280 9752 24337
rect 9786 24280 9792 24337
rect 9746 24265 9792 24280
rect 9746 24212 9752 24265
rect 9786 24212 9792 24265
rect 9746 24193 9792 24212
rect 9746 24144 9752 24193
rect 9786 24144 9792 24193
rect 9746 24121 9792 24144
rect 9746 24076 9752 24121
rect 9786 24076 9792 24121
rect 9746 24049 9792 24076
rect 9746 24008 9752 24049
rect 9786 24008 9792 24049
rect 9746 23977 9792 24008
rect 9746 23940 9752 23977
rect 9786 23940 9792 23977
rect 9746 23906 9792 23940
rect 9746 23871 9752 23906
rect 9786 23871 9792 23906
rect 9746 23838 9792 23871
rect 9746 23799 9752 23838
rect 9786 23799 9792 23838
rect 9746 23770 9792 23799
rect 9746 23727 9752 23770
rect 9786 23727 9792 23770
rect 9746 23702 9792 23727
rect 9746 23655 9752 23702
rect 9786 23655 9792 23702
rect 9746 23634 9792 23655
rect 9746 23583 9752 23634
rect 9786 23583 9792 23634
rect 9746 23566 9792 23583
rect 9746 23511 9752 23566
rect 9786 23511 9792 23566
rect 9746 23498 9792 23511
rect 9746 23439 9752 23498
rect 9786 23439 9792 23498
rect 9746 23430 9792 23439
rect 9746 23367 9752 23430
rect 9786 23367 9792 23430
rect 9746 23362 9792 23367
rect 9746 23295 9752 23362
rect 9786 23295 9792 23362
rect 9746 23294 9792 23295
rect 9746 23260 9752 23294
rect 9786 23260 9792 23294
rect 9746 23257 9792 23260
rect 9746 23192 9752 23257
rect 9786 23192 9792 23257
rect 9746 23185 9792 23192
rect 9746 23124 9752 23185
rect 9786 23124 9792 23185
rect 9746 23113 9792 23124
rect 9746 23056 9752 23113
rect 9786 23056 9792 23113
rect 9746 23041 9792 23056
rect 9746 22988 9752 23041
rect 9786 22988 9792 23041
rect 9746 22969 9792 22988
rect 9746 22920 9752 22969
rect 9786 22920 9792 22969
rect 9746 22897 9792 22920
rect 9746 22852 9752 22897
rect 9786 22852 9792 22897
rect 9746 22825 9792 22852
rect 9746 22784 9752 22825
rect 9786 22784 9792 22825
rect 9746 22753 9792 22784
rect 9746 22716 9752 22753
rect 9786 22716 9792 22753
rect 9746 22682 9792 22716
rect 9746 22647 9752 22682
rect 9786 22647 9792 22682
rect 9746 22614 9792 22647
rect 9746 22575 9752 22614
rect 9786 22575 9792 22614
rect 9746 22546 9792 22575
rect 9746 22503 9752 22546
rect 9786 22503 9792 22546
rect 9746 22478 9792 22503
rect 9746 22431 9752 22478
rect 9786 22431 9792 22478
rect 9746 22410 9792 22431
rect 9746 22359 9752 22410
rect 9786 22359 9792 22410
rect 9746 22342 9792 22359
rect 9746 22287 9752 22342
rect 9786 22287 9792 22342
rect 9746 22274 9792 22287
rect 9746 22215 9752 22274
rect 9786 22215 9792 22274
rect 9746 22206 9792 22215
rect 9746 22143 9752 22206
rect 9786 22143 9792 22206
rect 9746 22138 9792 22143
rect 9746 22071 9752 22138
rect 9786 22071 9792 22138
rect 9746 22070 9792 22071
rect 9746 22036 9752 22070
rect 9786 22036 9792 22070
rect 9746 22033 9792 22036
rect 9746 21968 9752 22033
rect 9786 21968 9792 22033
rect 9746 21961 9792 21968
rect 9746 21900 9752 21961
rect 9786 21900 9792 21961
rect 9746 21889 9792 21900
rect 9746 21832 9752 21889
rect 9786 21832 9792 21889
rect 9746 21817 9792 21832
rect 9746 21764 9752 21817
rect 9786 21764 9792 21817
rect 9746 21745 9792 21764
rect 9746 21696 9752 21745
rect 9786 21696 9792 21745
rect 9746 21673 9792 21696
rect 9746 21628 9752 21673
rect 9786 21628 9792 21673
rect 9746 21601 9792 21628
rect 9746 21560 9752 21601
rect 9786 21560 9792 21601
rect 9746 21529 9792 21560
rect 9746 21492 9752 21529
rect 9786 21492 9792 21529
rect 9746 21458 9792 21492
rect 9746 21423 9752 21458
rect 9786 21423 9792 21458
rect 9746 21390 9792 21423
rect 9746 21351 9752 21390
rect 9786 21351 9792 21390
rect 9746 21322 9792 21351
rect 9746 21279 9752 21322
rect 9786 21279 9792 21322
rect 9746 21254 9792 21279
rect 9746 21207 9752 21254
rect 9786 21207 9792 21254
rect 9746 21186 9792 21207
rect 9746 21135 9752 21186
rect 9786 21135 9792 21186
rect 9746 21118 9792 21135
rect 9746 21063 9752 21118
rect 9786 21063 9792 21118
rect 9746 21050 9792 21063
rect 9746 20991 9752 21050
rect 9786 20991 9792 21050
rect 9746 20982 9792 20991
rect 9746 20919 9752 20982
rect 9786 20919 9792 20982
rect 9746 20914 9792 20919
rect 9746 20847 9752 20914
rect 9786 20847 9792 20914
rect 9746 20846 9792 20847
rect 9746 20812 9752 20846
rect 9786 20812 9792 20846
rect 9746 20809 9792 20812
rect 9746 20744 9752 20809
rect 9786 20744 9792 20809
rect 9746 20737 9792 20744
rect 9746 20676 9752 20737
rect 9786 20676 9792 20737
rect 9746 20665 9792 20676
rect 9746 20608 9752 20665
rect 9786 20608 9792 20665
rect 9746 20593 9792 20608
rect 9746 20540 9752 20593
rect 9786 20540 9792 20593
rect 9746 20521 9792 20540
rect 9746 20472 9752 20521
rect 9786 20472 9792 20521
rect 9746 20449 9792 20472
rect 9746 20404 9752 20449
rect 9786 20404 9792 20449
rect 9746 20377 9792 20404
rect 9746 20336 9752 20377
rect 9786 20336 9792 20377
rect 9746 20305 9792 20336
rect 9746 20268 9752 20305
rect 9786 20268 9792 20305
rect 9746 20234 9792 20268
rect 9746 20199 9752 20234
rect 9786 20199 9792 20234
rect 9746 20166 9792 20199
rect 9746 20127 9752 20166
rect 9786 20127 9792 20166
rect 9746 20098 9792 20127
rect 9746 20055 9752 20098
rect 9786 20055 9792 20098
rect 9746 20030 9792 20055
rect 9746 19983 9752 20030
rect 9786 19983 9792 20030
rect 9746 19962 9792 19983
rect 9746 19911 9752 19962
rect 9786 19911 9792 19962
rect 9746 19894 9792 19911
rect 9746 19839 9752 19894
rect 9786 19839 9792 19894
rect 9746 19826 9792 19839
rect 9746 19767 9752 19826
rect 9786 19767 9792 19826
rect 9746 19758 9792 19767
rect 9746 19695 9752 19758
rect 9786 19695 9792 19758
rect 9746 19690 9792 19695
rect 9746 19623 9752 19690
rect 9786 19623 9792 19690
rect 9746 19622 9792 19623
rect 9746 19588 9752 19622
rect 9786 19588 9792 19622
rect 9746 19585 9792 19588
rect 9746 19520 9752 19585
rect 9786 19520 9792 19585
rect 9746 19513 9792 19520
rect 9746 19452 9752 19513
rect 9786 19452 9792 19513
rect 9746 19441 9792 19452
rect 9746 19384 9752 19441
rect 9786 19384 9792 19441
rect 9746 19369 9792 19384
rect 9746 19316 9752 19369
rect 9786 19316 9792 19369
rect 9746 19297 9792 19316
rect 9746 19248 9752 19297
rect 9786 19248 9792 19297
rect 9746 19225 9792 19248
rect 9746 19180 9752 19225
rect 9786 19180 9792 19225
rect 9746 19153 9792 19180
rect 9746 19112 9752 19153
rect 9786 19112 9792 19153
rect 9746 19081 9792 19112
rect 9746 19044 9752 19081
rect 9786 19044 9792 19081
rect 9746 19010 9792 19044
rect 9746 18975 9752 19010
rect 9786 18975 9792 19010
rect 9746 18942 9792 18975
rect 9746 18903 9752 18942
rect 9786 18903 9792 18942
rect 9746 18874 9792 18903
rect 9746 18831 9752 18874
rect 9786 18831 9792 18874
rect 9746 18806 9792 18831
rect 9746 18759 9752 18806
rect 9786 18759 9792 18806
rect 9746 18738 9792 18759
rect 9746 18687 9752 18738
rect 9786 18687 9792 18738
rect 9746 18670 9792 18687
rect 9746 18615 9752 18670
rect 9786 18615 9792 18670
rect 9746 18602 9792 18615
rect 9746 18543 9752 18602
rect 9786 18543 9792 18602
rect 9746 18534 9792 18543
rect 9746 18471 9752 18534
rect 9786 18471 9792 18534
rect 9746 18466 9792 18471
rect 9746 18399 9752 18466
rect 9786 18399 9792 18466
rect 9746 18398 9792 18399
rect 9746 18364 9752 18398
rect 9786 18364 9792 18398
rect 9746 18361 9792 18364
rect 9746 18296 9752 18361
rect 9786 18296 9792 18361
rect 9746 18289 9792 18296
rect 9746 18228 9752 18289
rect 9786 18228 9792 18289
rect 9746 18217 9792 18228
rect 9746 18160 9752 18217
rect 9786 18160 9792 18217
rect 9746 18145 9792 18160
rect 9746 18092 9752 18145
rect 9786 18092 9792 18145
rect 9746 18073 9792 18092
rect 9746 18024 9752 18073
rect 9786 18024 9792 18073
rect 9746 18001 9792 18024
rect 9746 17956 9752 18001
rect 9786 17956 9792 18001
rect 9746 17929 9792 17956
rect 9746 17888 9752 17929
rect 9786 17888 9792 17929
rect 9746 17857 9792 17888
rect 9746 17820 9752 17857
rect 9786 17820 9792 17857
rect 9746 17786 9792 17820
rect 9746 17751 9752 17786
rect 9786 17751 9792 17786
rect 9746 17718 9792 17751
rect 9746 17679 9752 17718
rect 9786 17679 9792 17718
rect 9746 17650 9792 17679
rect 9746 17607 9752 17650
rect 9786 17607 9792 17650
rect 9746 17582 9792 17607
rect 9746 17535 9752 17582
rect 9786 17535 9792 17582
rect 9746 17514 9792 17535
rect 9746 17463 9752 17514
rect 9786 17463 9792 17514
rect 9746 17446 9792 17463
rect 9746 17391 9752 17446
rect 9786 17391 9792 17446
rect 9746 17378 9792 17391
rect 9746 17319 9752 17378
rect 9786 17319 9792 17378
rect 9746 17310 9792 17319
rect 9746 17247 9752 17310
rect 9786 17247 9792 17310
rect 9746 17242 9792 17247
rect 9746 17175 9752 17242
rect 9786 17175 9792 17242
rect 9746 17174 9792 17175
rect 9746 17140 9752 17174
rect 9786 17140 9792 17174
rect 9746 17137 9792 17140
rect 9746 17072 9752 17137
rect 9786 17072 9792 17137
rect 9746 17065 9792 17072
rect 9746 17004 9752 17065
rect 9786 17004 9792 17065
rect 9746 16993 9792 17004
rect 9746 16936 9752 16993
rect 9786 16936 9792 16993
rect 9746 16921 9792 16936
rect 9746 16868 9752 16921
rect 9786 16868 9792 16921
rect 9746 16849 9792 16868
rect 9746 16800 9752 16849
rect 9786 16800 9792 16849
rect 9746 16777 9792 16800
rect 9746 16732 9752 16777
rect 9786 16732 9792 16777
rect 9746 16705 9792 16732
rect 9746 16664 9752 16705
rect 9786 16664 9792 16705
rect 9746 16633 9792 16664
rect 9746 16596 9752 16633
rect 9786 16596 9792 16633
rect 9746 16562 9792 16596
rect 9746 16527 9752 16562
rect 9786 16527 9792 16562
rect 9746 16494 9792 16527
rect 9746 16455 9752 16494
rect 9786 16455 9792 16494
rect 9746 16426 9792 16455
rect 9746 16383 9752 16426
rect 9786 16383 9792 16426
rect 9746 16358 9792 16383
rect 9746 16311 9752 16358
rect 9786 16311 9792 16358
rect 9746 16290 9792 16311
rect 9746 16239 9752 16290
rect 9786 16239 9792 16290
rect 9746 16222 9792 16239
rect 9746 16167 9752 16222
rect 9786 16167 9792 16222
rect 9746 16154 9792 16167
rect 9746 16095 9752 16154
rect 9786 16095 9792 16154
rect 9746 16086 9792 16095
rect 9746 16023 9752 16086
rect 9786 16023 9792 16086
rect 9746 16018 9792 16023
rect 9746 15951 9752 16018
rect 9786 15951 9792 16018
rect 9746 15950 9792 15951
rect 9746 15916 9752 15950
rect 9786 15916 9792 15950
rect 9746 15913 9792 15916
rect 9746 15848 9752 15913
rect 9786 15848 9792 15913
rect 9746 15841 9792 15848
rect 9746 15780 9752 15841
rect 9786 15780 9792 15841
rect 9746 15769 9792 15780
rect 9746 15712 9752 15769
rect 9786 15712 9792 15769
rect 9746 15697 9792 15712
rect 9746 15644 9752 15697
rect 9786 15644 9792 15697
rect 9746 15625 9792 15644
rect 9746 15576 9752 15625
rect 9786 15576 9792 15625
rect 9746 15553 9792 15576
rect 9746 15508 9752 15553
rect 9786 15508 9792 15553
rect 9746 15481 9792 15508
rect 9746 15440 9752 15481
rect 9786 15440 9792 15481
rect 9746 15409 9792 15440
rect 9746 15372 9752 15409
rect 9786 15372 9792 15409
rect 9746 15338 9792 15372
rect 9746 15303 9752 15338
rect 9786 15303 9792 15338
rect 9746 15270 9792 15303
rect 9746 15231 9752 15270
rect 9786 15231 9792 15270
rect 9746 15202 9792 15231
rect 9746 15159 9752 15202
rect 9786 15159 9792 15202
rect 9746 15134 9792 15159
rect 9746 15087 9752 15134
rect 9786 15087 9792 15134
rect 9746 15066 9792 15087
rect 9746 15015 9752 15066
rect 9786 15015 9792 15066
rect 9746 14998 9792 15015
rect 9746 14943 9752 14998
rect 9786 14943 9792 14998
rect 9746 14930 9792 14943
rect 9746 14871 9752 14930
rect 9786 14871 9792 14930
rect 9746 14862 9792 14871
rect 9746 14799 9752 14862
rect 9786 14799 9792 14862
rect 9746 14794 9792 14799
rect 9746 14727 9752 14794
rect 9786 14727 9792 14794
rect 9746 14726 9792 14727
rect 9746 14692 9752 14726
rect 9786 14692 9792 14726
rect 9746 14689 9792 14692
rect 9746 14624 9752 14689
rect 9786 14624 9792 14689
rect 9746 14617 9792 14624
rect 9746 14556 9752 14617
rect 9786 14556 9792 14617
rect 9746 14545 9792 14556
rect 9746 14488 9752 14545
rect 9786 14488 9792 14545
rect 9746 14473 9792 14488
rect 9746 14420 9752 14473
rect 9786 14420 9792 14473
rect 9746 14401 9792 14420
rect 9746 14352 9752 14401
rect 9786 14352 9792 14401
rect 9746 14329 9792 14352
rect 9746 14284 9752 14329
rect 9786 14284 9792 14329
rect 9746 14257 9792 14284
rect 9746 14216 9752 14257
rect 9786 14216 9792 14257
rect 9746 14185 9792 14216
rect 9746 14148 9752 14185
rect 9786 14148 9792 14185
rect 9746 14114 9792 14148
rect 9746 14079 9752 14114
rect 9786 14079 9792 14114
rect 9746 14046 9792 14079
rect 9746 14007 9752 14046
rect 9786 14007 9792 14046
rect 9746 13978 9792 14007
rect 9746 13935 9752 13978
rect 9786 13935 9792 13978
rect 9746 13910 9792 13935
rect 9746 13863 9752 13910
rect 9786 13863 9792 13910
rect 9746 13842 9792 13863
rect 9746 13791 9752 13842
rect 9786 13791 9792 13842
rect 9746 13774 9792 13791
rect 9746 13719 9752 13774
rect 9786 13719 9792 13774
rect 9746 13706 9792 13719
rect 9746 13647 9752 13706
rect 9786 13647 9792 13706
rect 9746 13638 9792 13647
rect 9746 13575 9752 13638
rect 9786 13575 9792 13638
rect 9746 13570 9792 13575
rect 9746 13503 9752 13570
rect 9786 13503 9792 13570
rect 9746 13502 9792 13503
rect 9746 13468 9752 13502
rect 9786 13468 9792 13502
rect 9746 13465 9792 13468
rect 9746 13400 9752 13465
rect 9786 13400 9792 13465
rect 9746 13393 9792 13400
rect 9746 13332 9752 13393
rect 9786 13332 9792 13393
rect 9746 13321 9792 13332
rect 9746 13264 9752 13321
rect 9786 13264 9792 13321
rect 9746 13249 9792 13264
rect 9746 13196 9752 13249
rect 9786 13196 9792 13249
rect 9746 13177 9792 13196
rect 9746 13128 9752 13177
rect 9786 13128 9792 13177
rect 9746 13105 9792 13128
rect 9746 13060 9752 13105
rect 9786 13060 9792 13105
rect 9746 13033 9792 13060
rect 9746 12992 9752 13033
rect 9786 12992 9792 13033
rect 9746 12961 9792 12992
rect 9746 12924 9752 12961
rect 9786 12924 9792 12961
rect 9746 12890 9792 12924
rect 9746 12855 9752 12890
rect 9786 12855 9792 12890
rect 9746 12822 9792 12855
rect 9746 12783 9752 12822
rect 9786 12783 9792 12822
rect 9746 12754 9792 12783
rect 9746 12711 9752 12754
rect 9786 12711 9792 12754
rect 9746 12686 9792 12711
rect 9746 12639 9752 12686
rect 9786 12639 9792 12686
rect 9746 12618 9792 12639
rect 9746 12567 9752 12618
rect 9786 12567 9792 12618
rect 9746 12550 9792 12567
rect 9746 12495 9752 12550
rect 9786 12495 9792 12550
rect 9746 12482 9792 12495
rect 9746 12423 9752 12482
rect 9786 12423 9792 12482
rect 9746 12414 9792 12423
rect 9746 12351 9752 12414
rect 9786 12351 9792 12414
rect 9746 12346 9792 12351
rect 9746 12279 9752 12346
rect 9786 12279 9792 12346
rect 9746 12278 9792 12279
rect 9746 12244 9752 12278
rect 9786 12244 9792 12278
rect 9746 12241 9792 12244
rect 9746 12176 9752 12241
rect 9786 12176 9792 12241
rect 9746 12169 9792 12176
rect 9746 12108 9752 12169
rect 9786 12108 9792 12169
rect 9746 12097 9792 12108
rect 9746 12040 9752 12097
rect 9786 12040 9792 12097
rect 9746 12025 9792 12040
rect 9746 11972 9752 12025
rect 9786 11972 9792 12025
rect 9746 11953 9792 11972
rect 9746 11904 9752 11953
rect 9786 11904 9792 11953
rect 9746 11881 9792 11904
rect 9746 11836 9752 11881
rect 9786 11836 9792 11881
rect 9746 11809 9792 11836
rect 9746 11768 9752 11809
rect 9786 11768 9792 11809
rect 9746 11737 9792 11768
rect 9746 11700 9752 11737
rect 9786 11700 9792 11737
rect 9746 11666 9792 11700
rect 9746 11631 9752 11666
rect 9786 11631 9792 11666
rect 9746 11598 9792 11631
rect 9746 11559 9752 11598
rect 9786 11559 9792 11598
rect 9746 11530 9792 11559
rect 9746 11487 9752 11530
rect 9786 11487 9792 11530
rect 9746 11462 9792 11487
rect 9746 11415 9752 11462
rect 9786 11415 9792 11462
rect 9746 11394 9792 11415
rect 9746 11343 9752 11394
rect 9786 11343 9792 11394
rect 9746 11326 9792 11343
rect 9746 11271 9752 11326
rect 9786 11271 9792 11326
rect 9746 11258 9792 11271
rect 9746 11199 9752 11258
rect 9786 11199 9792 11258
rect 9746 11190 9792 11199
rect 9746 11127 9752 11190
rect 9786 11127 9792 11190
rect 9746 11122 9792 11127
rect 9746 11055 9752 11122
rect 9786 11055 9792 11122
rect 9746 11054 9792 11055
rect 9746 11020 9752 11054
rect 9786 11020 9792 11054
rect 9746 11017 9792 11020
rect 9746 10952 9752 11017
rect 9786 10952 9792 11017
rect 9746 10945 9792 10952
rect 9746 10884 9752 10945
rect 9786 10884 9792 10945
rect 9746 10873 9792 10884
rect 9746 10816 9752 10873
rect 9786 10816 9792 10873
rect 9746 10801 9792 10816
rect 9746 10748 9752 10801
rect 9786 10748 9792 10801
rect 9746 10729 9792 10748
rect 9746 10680 9752 10729
rect 9786 10680 9792 10729
rect 9746 10657 9792 10680
rect 9746 10612 9752 10657
rect 9786 10612 9792 10657
rect 9746 10585 9792 10612
rect 9746 10544 9752 10585
rect 9786 10544 9792 10585
rect 9746 10513 9792 10544
rect 9746 10476 9752 10513
rect 9786 10476 9792 10513
rect 9746 10442 9792 10476
rect 9746 10407 9752 10442
rect 9786 10407 9792 10442
rect 9746 10374 9792 10407
rect 9746 10335 9752 10374
rect 9786 10335 9792 10374
rect 9746 10306 9792 10335
rect 9746 10263 9752 10306
rect 9786 10263 9792 10306
rect 9746 10238 9792 10263
rect 9746 10191 9752 10238
rect 9786 10191 9792 10238
rect 9746 10170 9792 10191
rect 9746 10119 9752 10170
rect 9786 10119 9792 10170
rect 9746 10102 9792 10119
rect 9746 10047 9752 10102
rect 9786 10047 9792 10102
rect 9746 10034 9792 10047
rect 9746 9975 9752 10034
rect 9786 9975 9792 10034
rect 9746 9966 9792 9975
rect 9746 9903 9752 9966
rect 9786 9903 9792 9966
rect 9746 9898 9792 9903
rect 9746 9831 9752 9898
rect 9786 9831 9792 9898
rect 9746 9830 9792 9831
rect 9746 9796 9752 9830
rect 9786 9796 9792 9830
rect 9746 9793 9792 9796
rect 9746 9728 9752 9793
rect 9786 9728 9792 9793
rect 9746 9721 9792 9728
rect 9746 9660 9752 9721
rect 9786 9660 9792 9721
rect 9746 9649 9792 9660
rect 9746 9592 9752 9649
rect 9786 9592 9792 9649
rect 9746 9577 9792 9592
rect 9746 9524 9752 9577
rect 9786 9524 9792 9577
rect 9746 9505 9792 9524
rect 9746 9456 9752 9505
rect 9786 9456 9792 9505
rect 9746 9433 9792 9456
rect 9746 9388 9752 9433
rect 9786 9388 9792 9433
rect 9746 9361 9792 9388
rect 9746 9320 9752 9361
rect 9786 9320 9792 9361
rect 9746 9289 9792 9320
rect 9746 9252 9752 9289
rect 9786 9252 9792 9289
rect 9746 9218 9792 9252
rect 9746 9183 9752 9218
rect 9786 9183 9792 9218
rect 9746 9150 9792 9183
rect 9746 9111 9752 9150
rect 9786 9111 9792 9150
rect 9746 9082 9792 9111
rect 9746 9039 9752 9082
rect 9786 9039 9792 9082
rect 9746 9014 9792 9039
rect 9746 8967 9752 9014
rect 9786 8967 9792 9014
rect 9746 8946 9792 8967
rect 9746 8895 9752 8946
rect 9786 8895 9792 8946
rect 9746 8878 9792 8895
rect 9746 8823 9752 8878
rect 9786 8823 9792 8878
rect 9746 8810 9792 8823
rect 9746 8751 9752 8810
rect 9786 8751 9792 8810
rect 9746 8742 9792 8751
rect 9746 8679 9752 8742
rect 9786 8679 9792 8742
rect 9746 8674 9792 8679
rect 9746 8607 9752 8674
rect 9786 8607 9792 8674
rect 9746 8606 9792 8607
rect 9746 8572 9752 8606
rect 9786 8572 9792 8606
rect 9746 8569 9792 8572
rect 9746 8504 9752 8569
rect 9786 8504 9792 8569
rect 9746 8497 9792 8504
rect 9746 8436 9752 8497
rect 9786 8436 9792 8497
rect 9746 8425 9792 8436
rect 9746 8368 9752 8425
rect 9786 8368 9792 8425
rect 9746 8353 9792 8368
rect 9746 8300 9752 8353
rect 9786 8300 9792 8353
rect 9746 8281 9792 8300
rect 9746 8232 9752 8281
rect 9786 8232 9792 8281
rect 9746 8209 9792 8232
rect 9746 8164 9752 8209
rect 9786 8164 9792 8209
rect 9746 8137 9792 8164
rect 9746 8096 9752 8137
rect 9786 8096 9792 8137
rect 9746 8065 9792 8096
rect 9746 8028 9752 8065
rect 9786 8028 9792 8065
rect 9746 7994 9792 8028
rect 9746 7959 9752 7994
rect 9786 7959 9792 7994
rect 9746 7926 9792 7959
rect 9746 7887 9752 7926
rect 9786 7887 9792 7926
rect 9746 7858 9792 7887
rect 9746 7815 9752 7858
rect 9786 7815 9792 7858
rect 9746 7790 9792 7815
rect 9746 7743 9752 7790
rect 9786 7743 9792 7790
rect 9746 7722 9792 7743
rect 9746 7671 9752 7722
rect 9786 7671 9792 7722
rect 9746 7654 9792 7671
rect 9746 7599 9752 7654
rect 9786 7599 9792 7654
rect 9746 7586 9792 7599
rect 9746 7527 9752 7586
rect 9786 7527 9792 7586
rect 9746 7518 9792 7527
rect 9746 7455 9752 7518
rect 9786 7455 9792 7518
rect 9746 7450 9792 7455
rect 9746 7383 9752 7450
rect 9786 7383 9792 7450
rect 9746 7382 9792 7383
rect 9746 7348 9752 7382
rect 9786 7348 9792 7382
rect 9746 7345 9792 7348
rect 9746 7280 9752 7345
rect 9786 7280 9792 7345
rect 9746 7273 9792 7280
rect 9746 7212 9752 7273
rect 9786 7212 9792 7273
rect 9746 7201 9792 7212
rect 9746 7144 9752 7201
rect 9786 7144 9792 7201
rect 9746 7129 9792 7144
rect 9746 7076 9752 7129
rect 9786 7076 9792 7129
rect 9746 7057 9792 7076
rect 9746 7008 9752 7057
rect 9786 7008 9792 7057
rect 9746 6985 9792 7008
rect 9746 6940 9752 6985
rect 9786 6940 9792 6985
rect 9746 6913 9792 6940
rect 9746 6872 9752 6913
rect 9786 6872 9792 6913
rect 9746 6841 9792 6872
rect 9746 6804 9752 6841
rect 9786 6804 9792 6841
rect 9746 6770 9792 6804
rect 9746 6735 9752 6770
rect 9786 6735 9792 6770
rect 9746 6702 9792 6735
rect 9746 6663 9752 6702
rect 9786 6663 9792 6702
rect 9746 6634 9792 6663
rect 9746 6591 9752 6634
rect 9786 6591 9792 6634
rect 9746 6566 9792 6591
rect 9746 6519 9752 6566
rect 9786 6519 9792 6566
rect 9746 6498 9792 6519
rect 9746 6447 9752 6498
rect 9786 6447 9792 6498
rect 9746 6430 9792 6447
rect 9746 6375 9752 6430
rect 9786 6375 9792 6430
rect 9746 6362 9792 6375
rect 9746 6303 9752 6362
rect 9786 6303 9792 6362
rect 9746 6294 9792 6303
rect 9746 6231 9752 6294
rect 9786 6231 9792 6294
rect 9746 6226 9792 6231
rect 9746 6159 9752 6226
rect 9786 6159 9792 6226
rect 9746 6158 9792 6159
rect 9746 6124 9752 6158
rect 9786 6124 9792 6158
rect 9746 6121 9792 6124
rect 9746 6056 9752 6121
rect 9786 6056 9792 6121
rect 9746 6049 9792 6056
rect 9746 5988 9752 6049
rect 9786 5988 9792 6049
rect 9746 5977 9792 5988
rect 9746 5920 9752 5977
rect 9786 5920 9792 5977
rect 9746 5905 9792 5920
rect 9746 5852 9752 5905
rect 9786 5852 9792 5905
rect 9746 5833 9792 5852
rect 9746 5784 9752 5833
rect 9786 5784 9792 5833
rect 9746 5761 9792 5784
rect 9746 5716 9752 5761
rect 9786 5716 9792 5761
rect 9746 5689 9792 5716
rect 9746 5648 9752 5689
rect 9786 5648 9792 5689
rect 9746 5617 9792 5648
rect 9746 5580 9752 5617
rect 9786 5580 9792 5617
rect 9746 5546 9792 5580
rect 9746 5511 9752 5546
rect 9786 5511 9792 5546
rect 9746 5478 9792 5511
rect 9746 5439 9752 5478
rect 9786 5439 9792 5478
rect 9746 5410 9792 5439
rect 9746 5367 9752 5410
rect 9786 5367 9792 5410
rect 9746 5342 9792 5367
rect 9746 5295 9752 5342
rect 9786 5295 9792 5342
rect 9746 5274 9792 5295
rect 9746 5223 9752 5274
rect 9786 5223 9792 5274
rect 9746 5206 9792 5223
rect 9746 5151 9752 5206
rect 9786 5151 9792 5206
rect 9746 5138 9792 5151
rect 9746 5079 9752 5138
rect 9786 5079 9792 5138
rect 9746 5070 9792 5079
rect 9746 5007 9752 5070
rect 9786 5007 9792 5070
rect 9746 5002 9792 5007
rect 9746 4935 9752 5002
rect 9786 4935 9792 5002
rect 9746 4934 9792 4935
rect 9746 4900 9752 4934
rect 9786 4900 9792 4934
rect 9746 4897 9792 4900
rect 9746 4832 9752 4897
rect 9786 4832 9792 4897
rect 9746 4825 9792 4832
rect 9746 4764 9752 4825
rect 9786 4764 9792 4825
rect 9746 4753 9792 4764
rect 9746 4696 9752 4753
rect 9786 4696 9792 4753
rect 9746 4681 9792 4696
rect 9746 4628 9752 4681
rect 9786 4628 9792 4681
rect 9746 4609 9792 4628
rect 9746 4560 9752 4609
rect 9786 4560 9792 4609
rect 9746 4537 9792 4560
rect 9746 4492 9752 4537
rect 9786 4492 9792 4537
rect 9746 4465 9792 4492
rect 9746 4424 9752 4465
rect 9786 4424 9792 4465
rect 9746 4393 9792 4424
rect 9746 4356 9752 4393
rect 9786 4356 9792 4393
rect 9746 4322 9792 4356
rect 9746 4287 9752 4322
rect 9786 4287 9792 4322
rect 9746 4254 9792 4287
rect 9746 4215 9752 4254
rect 9786 4215 9792 4254
rect 9746 4186 9792 4215
rect 9746 4143 9752 4186
rect 9786 4143 9792 4186
rect 9746 4118 9792 4143
rect 9746 4071 9752 4118
rect 9786 4071 9792 4118
rect 9746 4050 9792 4071
rect 9746 3999 9752 4050
rect 9786 3999 9792 4050
rect 9746 3982 9792 3999
rect 9746 3927 9752 3982
rect 9786 3927 9792 3982
rect 9746 3914 9792 3927
rect 9746 3855 9752 3914
rect 9786 3855 9792 3914
rect 9746 3846 9792 3855
rect 9746 3783 9752 3846
rect 9786 3783 9792 3846
rect 9746 3778 9792 3783
rect 9746 3711 9752 3778
rect 9786 3711 9792 3778
rect 9746 3710 9792 3711
rect 9746 3676 9752 3710
rect 9786 3676 9792 3710
rect 9746 3673 9792 3676
rect 9746 3608 9752 3673
rect 9786 3608 9792 3673
rect 9746 3601 9792 3608
rect 9746 3540 9752 3601
rect 9786 3540 9792 3601
rect 9746 3529 9792 3540
rect 9746 3472 9752 3529
rect 9786 3472 9792 3529
rect 9746 3457 9792 3472
rect 9746 3404 9752 3457
rect 9786 3404 9792 3457
rect 9746 3385 9792 3404
rect 9746 3336 9752 3385
rect 9786 3336 9792 3385
rect 9746 3313 9792 3336
rect 9746 3268 9752 3313
rect 9786 3268 9792 3313
rect 9746 3241 9792 3268
rect 9746 3200 9752 3241
rect 9786 3200 9792 3241
rect 9746 3168 9792 3200
rect 9746 3132 9752 3168
rect 9786 3132 9792 3168
rect 9746 3098 9792 3132
rect 9746 3061 9752 3098
rect 9786 3061 9792 3098
rect 9746 3030 9792 3061
rect 9746 2988 9752 3030
rect 9786 2988 9792 3030
rect 9746 2962 9792 2988
rect 9746 2915 9752 2962
rect 9786 2915 9792 2962
rect 9746 2894 9792 2915
rect 9746 2842 9752 2894
rect 9786 2842 9792 2894
rect 9746 2826 9792 2842
rect 9746 2769 9752 2826
rect 9786 2769 9792 2826
rect 9746 2758 9792 2769
rect 9746 2696 9752 2758
rect 9786 2696 9792 2758
rect 9746 2690 9792 2696
rect 9746 2623 9752 2690
rect 9786 2623 9792 2690
rect 9746 2622 9792 2623
rect 9746 2588 9752 2622
rect 9786 2588 9792 2622
rect 9746 2584 9792 2588
rect 9746 2520 9752 2584
rect 9786 2520 9792 2584
rect 9746 2511 9792 2520
rect 9746 2452 9752 2511
rect 9786 2452 9792 2511
rect 9746 2438 9792 2452
rect 9746 2384 9752 2438
rect 9786 2384 9792 2438
rect 9746 2365 9792 2384
rect 9746 2315 9752 2365
rect 9786 2315 9792 2365
rect 9746 2292 9792 2315
rect 9746 2246 9752 2292
rect 9786 2246 9792 2292
rect 9746 2219 9792 2246
rect 9746 2177 9752 2219
rect 9786 2177 9792 2219
rect 9746 2146 9792 2177
rect 9746 2108 9752 2146
rect 9786 2108 9792 2146
rect 9746 2073 9792 2108
rect 9746 2039 9752 2073
rect 9786 2039 9792 2073
rect 9746 2004 9792 2039
rect 9746 1966 9752 2004
rect 9786 1966 9792 2004
rect 9746 1935 9792 1966
rect 9746 1893 9752 1935
rect 9786 1893 9792 1935
rect 9746 1866 9792 1893
rect 9746 1820 9752 1866
rect 9786 1820 9792 1866
rect 9746 1797 9792 1820
rect 9746 1747 9752 1797
rect 9786 1747 9792 1797
rect 9746 1728 9792 1747
rect 9746 1674 9752 1728
rect 9786 1674 9792 1728
rect 9746 1659 9792 1674
rect 9746 1601 9752 1659
rect 9786 1601 9792 1659
rect 9746 1590 9792 1601
rect 9746 1528 9752 1590
rect 9786 1528 9792 1590
rect 9746 1521 9792 1528
rect 9746 1455 9752 1521
rect 9786 1455 9792 1521
rect 9746 1452 9792 1455
rect 9746 1418 9752 1452
rect 9786 1418 9792 1452
rect 9746 1416 9792 1418
rect 9746 1349 9752 1416
rect 9786 1349 9792 1416
rect 10710 2487 10716 39777
rect 10822 2487 10828 39817
rect 10710 2448 10718 2487
rect 10820 2448 10828 2487
rect 10710 2414 10716 2448
rect 10822 2414 10828 2448
rect 10710 2375 10718 2414
rect 10820 2375 10828 2414
rect 10710 2341 10716 2375
rect 10822 2341 10828 2375
rect 10710 2302 10718 2341
rect 10820 2302 10828 2341
rect 10710 2268 10716 2302
rect 10822 2268 10828 2302
rect 10710 2229 10718 2268
rect 10820 2229 10828 2268
rect 10710 2195 10716 2229
rect 10822 2195 10828 2229
rect 10710 2156 10718 2195
rect 10820 2156 10828 2195
rect 10710 2122 10716 2156
rect 10822 2122 10828 2156
rect 10710 2083 10718 2122
rect 10820 2083 10828 2122
rect 10710 2049 10716 2083
rect 10822 2049 10828 2083
rect 10710 2010 10718 2049
rect 10820 2010 10828 2049
rect 10710 1976 10716 2010
rect 10822 1976 10828 2010
rect 10710 1937 10718 1976
rect 10820 1937 10828 1976
rect 10710 1903 10716 1937
rect 10822 1903 10828 1937
rect 10710 1864 10718 1903
rect 10820 1864 10828 1903
rect 10710 1830 10716 1864
rect 10822 1830 10828 1864
rect 10710 1791 10718 1830
rect 10820 1791 10828 1830
rect 10710 1757 10716 1791
rect 10822 1757 10828 1791
rect 10710 1718 10718 1757
rect 10820 1718 10828 1757
rect 10710 1684 10716 1718
rect 10822 1684 10828 1718
rect 10710 1645 10718 1684
rect 10820 1645 10828 1684
rect 10710 1611 10716 1645
rect 10822 1611 10828 1645
rect 10710 1572 10718 1611
rect 10820 1572 10828 1611
rect 10710 1538 10716 1572
rect 10822 1538 10828 1572
rect 10710 1499 10718 1538
rect 10820 1499 10828 1538
rect 10710 1465 10716 1499
rect 10822 1465 10828 1499
rect 10710 1426 10718 1465
rect 10820 1426 10828 1465
rect 9746 1343 9792 1349
rect 9746 1280 9752 1343
rect 9786 1280 9792 1343
rect 9859 1399 10243 1411
rect 9859 1293 10137 1399
rect 10710 1392 10716 1426
rect 10822 1392 10828 1426
rect 10710 1353 10718 1392
rect 10820 1353 10828 1392
rect 10710 1319 10716 1353
rect 10822 1319 10828 1353
rect 9746 1270 9792 1280
rect 9746 1211 9752 1270
rect 9786 1211 9792 1270
rect 9746 1197 9792 1211
rect 9746 1142 9752 1197
rect 9786 1142 9792 1197
rect 9746 1124 9792 1142
rect 9746 1073 9752 1124
rect 9786 1073 9792 1124
rect 9746 1051 9792 1073
rect 9746 1004 9752 1051
rect 9786 1004 9792 1051
rect 9746 978 9792 1004
rect 9746 935 9752 978
rect 9786 935 9792 978
rect 9746 905 9792 935
rect 9746 866 9752 905
rect 9786 866 9792 905
rect 9746 832 9792 866
rect 9746 797 9752 832
rect 9786 797 9792 832
rect 9746 762 9792 797
rect 9746 725 9752 762
rect 9786 725 9792 762
rect 9746 693 9792 725
rect 9746 652 9752 693
rect 9786 652 9792 693
rect 9746 624 9792 652
rect 9746 579 9752 624
rect 9786 579 9792 624
rect 9746 555 9792 579
rect 9746 506 9752 555
rect 9786 506 9792 555
rect 9746 486 9792 506
rect 9746 433 9752 486
rect 9786 433 9792 486
rect 9746 417 9792 433
rect 9746 401 9752 417
rect 8000 378 8002 384
rect 8034 344 8036 350
rect 8000 315 8036 344
rect 8000 305 8002 315
rect 8034 271 8036 281
rect 8000 246 8036 271
rect 8000 232 8002 246
rect 8034 198 8036 212
rect 8000 177 8036 198
rect 8000 159 8002 177
rect 2448 74 2590 108
rect 2448 40 2482 74
rect 2516 40 2590 74
rect 7977 125 8000 142
rect 8034 142 8036 143
rect 9786 401 9792 417
rect 10710 1280 10718 1319
rect 10820 1280 10828 1319
rect 10710 1246 10716 1280
rect 10822 1246 10828 1280
rect 10710 1207 10718 1246
rect 10820 1207 10828 1246
rect 10710 1173 10716 1207
rect 10822 1173 10828 1207
rect 10710 1134 10718 1173
rect 10820 1134 10828 1173
rect 10710 1100 10716 1134
rect 10822 1100 10828 1134
rect 10710 1061 10718 1100
rect 10820 1061 10828 1100
rect 10710 1027 10716 1061
rect 10822 1027 10828 1061
rect 10710 988 10718 1027
rect 10820 988 10828 1027
rect 10710 954 10716 988
rect 10822 954 10828 988
rect 10710 915 10718 954
rect 10820 915 10828 954
rect 10710 881 10716 915
rect 10822 881 10828 915
rect 10710 842 10718 881
rect 10820 842 10828 881
rect 10710 808 10716 842
rect 10822 808 10828 842
rect 10710 769 10718 808
rect 10820 769 10828 808
rect 10710 735 10716 769
rect 10822 735 10828 769
rect 10710 696 10718 735
rect 10820 696 10828 735
rect 10710 662 10716 696
rect 10822 662 10828 696
rect 10710 623 10718 662
rect 10820 623 10828 662
rect 10710 589 10716 623
rect 10822 589 10828 623
rect 10710 550 10718 589
rect 10820 550 10828 589
rect 10710 516 10716 550
rect 10822 516 10828 550
rect 10710 477 10718 516
rect 10820 477 10828 516
rect 10710 443 10716 477
rect 10822 443 10828 477
rect 10710 404 10718 443
rect 10820 404 10828 443
rect 9752 348 9786 383
rect 9752 279 9786 314
rect 9752 210 9786 245
rect 9752 142 9786 176
rect 10710 370 10716 404
rect 10822 370 10828 404
rect 10710 331 10718 370
rect 10820 331 10828 370
rect 10710 297 10716 331
rect 10822 297 10828 331
rect 10710 258 10718 297
rect 10820 258 10828 297
rect 10710 224 10716 258
rect 10822 224 10828 258
rect 10710 185 10718 224
rect 10820 185 10828 224
rect 10710 151 10716 185
rect 10822 151 10828 185
rect 10710 142 10718 151
rect 8034 125 8096 142
rect 7977 108 8096 125
rect 7977 86 8002 108
rect 7977 52 8000 86
rect 8036 74 8096 108
rect 8034 52 8096 74
rect 7977 40 8096 52
rect 10646 112 10718 142
rect 10820 112 10828 151
rect 10646 78 10716 112
rect 10750 78 10788 108
rect 10822 78 10828 112
rect 10646 74 10828 78
rect 10646 40 10680 74
rect 10714 40 10828 74
<< viali >>
rect 445 39886 479 39888
rect 518 39886 552 39888
rect 591 39886 625 39888
rect 664 39886 698 39888
rect 737 39886 771 39888
rect 810 39886 844 39888
rect 884 39886 918 39888
rect 958 39886 992 39888
rect 1032 39886 1066 39888
rect 1106 39886 1140 39888
rect 1216 39886 1250 39888
rect 1290 39886 1324 39888
rect 1364 39886 1398 39888
rect 1438 39886 1472 39888
rect 1512 39886 1546 39888
rect 1587 39886 1621 39888
rect 1662 39886 1696 39888
rect 1737 39886 1771 39888
rect 1812 39886 1846 39888
rect 1887 39886 1921 39888
rect 1962 39886 1996 39888
rect 2037 39886 2071 39888
rect 2112 39886 2146 39888
rect 2187 39886 2221 39888
rect 2262 39886 2296 39888
rect 2337 39886 2371 39888
rect 2412 39886 2446 39888
rect 2487 39886 2521 39888
rect 445 39854 448 39886
rect 448 39854 479 39886
rect 518 39854 552 39886
rect 591 39854 625 39886
rect 664 39854 698 39886
rect 737 39854 771 39886
rect 810 39854 844 39886
rect 884 39854 918 39886
rect 958 39854 992 39886
rect 1032 39854 1066 39886
rect 1106 39854 1140 39886
rect 1216 39854 1250 39886
rect 1290 39854 1324 39886
rect 1364 39854 1398 39886
rect 1438 39854 1472 39886
rect 1512 39854 1546 39886
rect 1587 39854 1621 39886
rect 1662 39854 1696 39886
rect 1737 39854 1771 39886
rect 1812 39854 1846 39886
rect 1887 39854 1921 39886
rect 1962 39854 1996 39886
rect 2037 39854 2071 39886
rect 2112 39854 2146 39886
rect 2187 39854 2221 39886
rect 2262 39854 2296 39886
rect 2337 39854 2371 39886
rect 2412 39854 2446 39886
rect 2487 39854 2521 39886
rect 372 39782 374 39816
rect 374 39782 406 39816
rect 444 39782 476 39816
rect 476 39782 478 39816
rect 518 39784 552 39816
rect 591 39784 625 39816
rect 664 39784 698 39816
rect 737 39784 771 39816
rect 810 39784 844 39816
rect 884 39784 918 39816
rect 958 39784 992 39816
rect 1032 39784 1066 39816
rect 1106 39784 1140 39816
rect 1216 39784 1250 39816
rect 1290 39784 1324 39816
rect 1364 39784 1398 39816
rect 1438 39784 1472 39816
rect 1512 39784 1546 39816
rect 1587 39784 1621 39816
rect 1662 39784 1696 39816
rect 1737 39784 1771 39816
rect 1812 39784 1846 39816
rect 1887 39784 1921 39816
rect 1962 39784 1996 39816
rect 2037 39784 2071 39816
rect 2112 39784 2146 39816
rect 2187 39784 2221 39816
rect 2262 39784 2296 39816
rect 2337 39784 2371 39816
rect 2412 39784 2446 39816
rect 2487 39784 2522 39816
rect 2522 39786 2593 39816
rect 2522 39784 2556 39786
rect 518 39782 552 39784
rect 591 39782 625 39784
rect 664 39782 698 39784
rect 737 39782 771 39784
rect 810 39782 844 39784
rect 884 39782 918 39784
rect 958 39782 992 39784
rect 1032 39782 1066 39784
rect 1106 39782 1140 39784
rect 1216 39782 1250 39784
rect 1290 39782 1324 39784
rect 1364 39782 1398 39784
rect 1438 39782 1472 39784
rect 1512 39782 1546 39784
rect 1587 39782 1621 39784
rect 1662 39782 1696 39784
rect 1737 39782 1771 39784
rect 1812 39782 1846 39784
rect 1887 39782 1921 39784
rect 1962 39782 1996 39784
rect 2037 39782 2071 39784
rect 2112 39782 2146 39784
rect 2187 39782 2221 39784
rect 2262 39782 2296 39784
rect 2337 39782 2371 39784
rect 2412 39782 2446 39784
rect 372 39709 374 39743
rect 374 39709 406 39743
rect 444 39709 476 39743
rect 476 39709 478 39743
rect 372 39636 374 39670
rect 374 39636 406 39670
rect 444 39636 476 39670
rect 476 39636 478 39670
rect 372 39563 374 39597
rect 374 39563 406 39597
rect 444 39563 476 39597
rect 476 39563 478 39597
rect 372 39490 374 39524
rect 374 39490 406 39524
rect 444 39490 476 39524
rect 476 39490 478 39524
rect 566 39667 600 39701
rect 638 39667 672 39701
rect 566 39594 600 39628
rect 638 39594 672 39628
rect 566 39521 600 39555
rect 638 39521 672 39555
rect 2310 39679 2344 39713
rect 2382 39679 2416 39713
rect 2310 39606 2344 39640
rect 2382 39606 2416 39640
rect 2310 39533 2344 39567
rect 2382 39533 2416 39567
rect 372 39417 374 39451
rect 374 39417 406 39451
rect 444 39417 476 39451
rect 476 39417 478 39451
rect 372 39344 374 39378
rect 374 39344 406 39378
rect 444 39344 476 39378
rect 476 39344 478 39378
rect 372 39271 374 39305
rect 374 39271 406 39305
rect 444 39271 476 39305
rect 476 39271 478 39305
rect 372 39198 374 39232
rect 374 39198 406 39232
rect 444 39198 476 39232
rect 476 39198 478 39232
rect 372 39125 374 39159
rect 374 39125 406 39159
rect 444 39125 476 39159
rect 476 39125 478 39159
rect 372 39052 374 39086
rect 374 39052 406 39086
rect 444 39052 476 39086
rect 476 39052 478 39086
rect 372 38979 374 39013
rect 374 38979 406 39013
rect 444 38979 476 39013
rect 476 38979 478 39013
rect 372 38906 374 38940
rect 374 38906 406 38940
rect 444 38906 476 38940
rect 476 38906 478 38940
rect 372 38833 374 38867
rect 374 38833 406 38867
rect 444 38833 476 38867
rect 476 38833 478 38867
rect 372 38760 374 38794
rect 374 38760 406 38794
rect 444 38760 476 38794
rect 476 38760 478 38794
rect 372 38687 374 38721
rect 374 38687 406 38721
rect 444 38687 476 38721
rect 476 38687 478 38721
rect 372 38614 374 38648
rect 374 38614 406 38648
rect 444 38614 476 38648
rect 476 38614 478 38648
rect 372 38541 374 38575
rect 374 38541 406 38575
rect 444 38541 476 38575
rect 476 38541 478 38575
rect 372 38468 374 38502
rect 374 38468 406 38502
rect 444 38468 476 38502
rect 476 38468 478 38502
rect 372 38395 374 38429
rect 374 38395 406 38429
rect 444 38395 476 38429
rect 476 38395 478 38429
rect 372 38322 374 38356
rect 374 38322 406 38356
rect 444 38322 476 38356
rect 476 38322 478 38356
rect 372 38249 374 38283
rect 374 38249 406 38283
rect 444 38249 476 38283
rect 476 38249 478 38283
rect 372 38176 374 38210
rect 374 38176 406 38210
rect 444 38176 476 38210
rect 476 38176 478 38210
rect 372 38103 374 38137
rect 374 38103 406 38137
rect 444 38103 476 38137
rect 476 38103 478 38137
rect 372 38030 374 38064
rect 374 38030 406 38064
rect 444 38030 476 38064
rect 476 38030 478 38064
rect 372 37957 374 37991
rect 374 37957 406 37991
rect 444 37957 476 37991
rect 476 37957 478 37991
rect 372 37884 374 37918
rect 374 37884 406 37918
rect 444 37884 476 37918
rect 476 37884 478 37918
rect 372 37811 374 37845
rect 374 37811 406 37845
rect 444 37811 476 37845
rect 476 37811 478 37845
rect 372 37738 374 37772
rect 374 37738 406 37772
rect 444 37738 476 37772
rect 476 37738 478 37772
rect 372 37665 374 37699
rect 374 37665 406 37699
rect 444 37665 476 37699
rect 476 37665 478 37699
rect 372 37592 374 37626
rect 374 37592 406 37626
rect 444 37592 476 37626
rect 476 37592 478 37626
rect 372 37519 374 37553
rect 374 37519 406 37553
rect 444 37519 476 37553
rect 476 37519 478 37553
rect 372 37446 374 37480
rect 374 37446 406 37480
rect 444 37446 476 37480
rect 476 37446 478 37480
rect 372 37373 374 37407
rect 374 37373 406 37407
rect 444 37373 476 37407
rect 476 37373 478 37407
rect 372 436 374 37334
rect 374 436 476 37334
rect 476 436 478 37334
rect 2487 39752 2556 39784
rect 2556 39752 2590 39786
rect 2590 39752 2593 39786
rect 2487 39718 2593 39752
rect 2487 2918 2488 39718
rect 2488 2918 2590 39718
rect 2590 2918 2593 39718
rect 8040 39886 8074 39889
rect 8116 39886 8150 39889
rect 8192 39886 8226 39889
rect 8268 39886 8302 39889
rect 8345 39886 8379 39889
rect 8422 39886 8456 39889
rect 8499 39886 8533 39889
rect 8576 39886 8610 39889
rect 8653 39886 8687 39889
rect 8730 39886 8764 39889
rect 8840 39886 10458 39889
rect 10497 39886 10531 39889
rect 10570 39886 10604 39889
rect 10643 39886 10677 39889
rect 10716 39886 10750 39889
rect 8040 39855 8066 39886
rect 8066 39855 8074 39886
rect 8116 39855 8150 39886
rect 8192 39855 8226 39886
rect 8268 39855 8302 39886
rect 8345 39855 8379 39886
rect 8422 39855 8456 39886
rect 8499 39855 8533 39886
rect 8576 39855 8610 39886
rect 8653 39855 8687 39886
rect 8730 39855 8764 39886
rect 8040 39784 8066 39817
rect 8066 39784 8074 39817
rect 8116 39784 8150 39817
rect 8192 39784 8226 39817
rect 8268 39784 8302 39817
rect 8345 39784 8379 39817
rect 8422 39784 8456 39817
rect 8499 39784 8533 39817
rect 8576 39784 8610 39817
rect 8653 39784 8687 39817
rect 8730 39784 8764 39817
rect 8840 39784 10458 39886
rect 10497 39855 10531 39886
rect 10570 39855 10604 39886
rect 10643 39855 10677 39886
rect 10716 39855 10750 39886
rect 10497 39784 10531 39817
rect 10570 39784 10604 39817
rect 10643 39784 10677 39817
rect 10716 39784 10752 39817
rect 10752 39786 10822 39817
rect 10752 39784 10786 39786
rect 8040 39783 8074 39784
rect 8116 39783 8150 39784
rect 8192 39783 8226 39784
rect 8268 39783 8302 39784
rect 8345 39783 8379 39784
rect 8422 39783 8456 39784
rect 8499 39783 8533 39784
rect 8576 39783 8610 39784
rect 8653 39783 8687 39784
rect 8730 39783 8764 39784
rect 8840 39783 10458 39784
rect 10497 39783 10531 39784
rect 10570 39783 10604 39784
rect 10643 39783 10677 39784
rect 8000 39716 8002 39742
rect 8002 39716 8034 39742
rect 8000 39708 8034 39716
rect 8000 39648 8002 39670
rect 8002 39648 8034 39670
rect 8000 39636 8034 39648
rect 5402 39580 5432 39614
rect 5432 39580 5436 39614
rect 5476 39580 5502 39614
rect 5502 39580 5510 39614
rect 5550 39580 5572 39614
rect 5572 39580 5584 39614
rect 5624 39580 5642 39614
rect 5642 39580 5658 39614
rect 5698 39580 5712 39614
rect 5712 39580 5732 39614
rect 5772 39580 5782 39614
rect 5782 39580 5806 39614
rect 5846 39580 5852 39614
rect 5852 39580 5880 39614
rect 5920 39580 5922 39614
rect 5922 39580 5954 39614
rect 5994 39580 6028 39614
rect 6068 39580 6098 39614
rect 6098 39580 6102 39614
rect 6142 39580 6168 39614
rect 6168 39580 6176 39614
rect 6216 39580 6238 39614
rect 6238 39580 6250 39614
rect 6290 39580 6308 39614
rect 6308 39580 6324 39614
rect 6364 39580 6378 39614
rect 6378 39580 6398 39614
rect 6438 39580 6448 39614
rect 6448 39580 6472 39614
rect 6512 39580 6518 39614
rect 6518 39580 6546 39614
rect 6586 39580 6588 39614
rect 6588 39580 6620 39614
rect 6660 39580 6691 39614
rect 6691 39580 6694 39614
rect 6734 39580 6760 39614
rect 6760 39580 6768 39614
rect 6808 39580 6829 39614
rect 6829 39580 6842 39614
rect 6882 39580 6898 39614
rect 6898 39580 6916 39614
rect 6956 39580 6967 39614
rect 6967 39580 6990 39614
rect 7030 39580 7036 39614
rect 7036 39580 7064 39614
rect 7104 39580 7105 39614
rect 7105 39580 7138 39614
rect 7178 39580 7209 39614
rect 7209 39580 7212 39614
rect 7251 39580 7278 39614
rect 7278 39580 7285 39614
rect 7324 39580 7347 39614
rect 7347 39580 7358 39614
rect 7397 39580 7416 39614
rect 7416 39580 7431 39614
rect 7470 39580 7504 39614
rect 8000 39580 8002 39598
rect 8002 39580 8034 39598
rect 8000 39564 8034 39580
rect 8112 39679 8146 39713
rect 8184 39679 8218 39713
rect 8112 39606 8146 39640
rect 8184 39606 8218 39640
rect 8112 39533 8146 39567
rect 8184 39533 8218 39567
rect 9564 39679 9598 39713
rect 9636 39679 9670 39713
rect 9564 39606 9598 39640
rect 9636 39617 9640 39640
rect 9640 39617 9670 39640
rect 9636 39606 9670 39617
rect 9564 39533 9598 39567
rect 9636 39533 9670 39567
rect 9752 39716 9786 39745
rect 9752 39711 9786 39716
rect 9752 39648 9786 39673
rect 9752 39639 9786 39648
rect 9752 39580 9786 39601
rect 9752 39567 9786 39580
rect 8000 39512 8002 39526
rect 8002 39512 8034 39526
rect 8000 39492 8034 39512
rect 7532 39329 7566 39356
rect 7532 39322 7566 39329
rect 7532 39261 7566 39284
rect 7532 39250 7566 39261
rect 7532 39193 7566 39212
rect 7532 39178 7566 39193
rect 7532 39125 7566 39140
rect 7532 39106 7566 39125
rect 7532 39057 7566 39068
rect 7532 39034 7566 39057
rect 7532 38989 7566 38996
rect 7532 38962 7566 38989
rect 7532 38921 7566 38924
rect 7532 38890 7566 38921
rect 7532 38819 7566 38852
rect 7532 38818 7566 38819
rect 7532 38751 7566 38780
rect 7532 38746 7566 38751
rect 7532 38683 7566 38708
rect 7532 38674 7566 38683
rect 7532 38615 7566 38636
rect 7532 38602 7566 38615
rect 7532 38547 7566 38564
rect 7532 38530 7566 38547
rect 7532 38479 7566 38492
rect 7532 38458 7566 38479
rect 7532 38411 7566 38420
rect 7532 38386 7566 38411
rect 7532 38343 7566 38348
rect 7532 38314 7566 38343
rect 7532 38275 7566 38276
rect 7532 38242 7566 38275
rect 7532 38173 7566 38204
rect 7532 38170 7566 38173
rect 7532 38105 7566 38132
rect 7532 38098 7566 38105
rect 7532 38037 7566 38060
rect 7532 38026 7566 38037
rect 7532 37969 7566 37988
rect 7532 37954 7566 37969
rect 7532 37901 7566 37916
rect 7532 37882 7566 37901
rect 7532 37833 7566 37844
rect 7532 37810 7566 37833
rect 7532 37765 7566 37772
rect 7532 37738 7566 37765
rect 7532 37697 7566 37700
rect 7532 37666 7566 37697
rect 7532 37595 7566 37628
rect 7532 37594 7566 37595
rect 7532 37527 7566 37556
rect 7532 37522 7566 37527
rect 7532 37459 7566 37484
rect 7532 37450 7566 37459
rect 7532 37391 7566 37412
rect 7532 37378 7566 37391
rect 7532 37323 7566 37340
rect 7532 37306 7566 37323
rect 7532 37255 7566 37267
rect 7532 37233 7566 37255
rect 7532 37187 7566 37194
rect 7532 37160 7566 37187
rect 7532 37119 7566 37121
rect 7532 37087 7566 37119
rect 7532 37017 7566 37048
rect 7532 37014 7566 37017
rect 7532 36949 7566 36975
rect 7532 36941 7566 36949
rect 7532 36881 7566 36902
rect 7532 36868 7566 36881
rect 7532 36813 7566 36829
rect 7532 36795 7566 36813
rect 7532 36745 7566 36756
rect 7532 36722 7566 36745
rect 7532 36677 7566 36683
rect 7532 36649 7566 36677
rect 7532 36609 7566 36610
rect 7532 36576 7566 36609
rect 7532 36507 7566 36537
rect 7532 36503 7566 36507
rect 7532 36439 7566 36464
rect 7532 36430 7566 36439
rect 7532 36370 7566 36391
rect 7532 36357 7566 36370
rect 7532 36301 7566 36318
rect 7532 36284 7566 36301
rect 7532 36232 7566 36245
rect 7532 36211 7566 36232
rect 7532 36163 7566 36172
rect 7532 36138 7566 36163
rect 7532 36094 7566 36099
rect 7532 36065 7566 36094
rect 7532 36025 7566 36026
rect 7532 35992 7566 36025
rect 7532 35922 7566 35953
rect 7532 35919 7566 35922
rect 7532 35853 7566 35880
rect 7532 35846 7566 35853
rect 7532 35784 7566 35807
rect 7532 35773 7566 35784
rect 7532 35715 7566 35734
rect 7532 35700 7566 35715
rect 7532 35646 7566 35661
rect 7532 35627 7566 35646
rect 7532 35577 7566 35588
rect 7532 35554 7566 35577
rect 7532 35508 7566 35515
rect 7532 35481 7566 35508
rect 7532 35439 7566 35442
rect 7532 35408 7566 35439
rect 7532 35335 7566 35369
rect 7532 35266 7566 35296
rect 7532 35262 7566 35266
rect 7532 35197 7566 35223
rect 7532 35189 7566 35197
rect 7532 35128 7566 35150
rect 7532 35116 7566 35128
rect 7532 35059 7566 35077
rect 7532 35043 7566 35059
rect 7532 34990 7566 35004
rect 7532 34970 7566 34990
rect 7532 34921 7566 34931
rect 7532 34897 7566 34921
rect 7532 34852 7566 34858
rect 7532 34824 7566 34852
rect 7532 34783 7566 34785
rect 7532 34751 7566 34783
rect 7532 34680 7566 34712
rect 7532 34678 7566 34680
rect 7532 34611 7566 34639
rect 7532 34605 7566 34611
rect 7532 34542 7566 34566
rect 7532 34532 7566 34542
rect 7532 34473 7566 34493
rect 7532 34459 7566 34473
rect 7532 34404 7566 34420
rect 7532 34386 7566 34404
rect 7532 34335 7566 34347
rect 7532 34313 7566 34335
rect 7532 34266 7566 34274
rect 7532 34240 7566 34266
rect 7532 34197 7566 34201
rect 7532 34167 7566 34197
rect 7532 34094 7566 34128
rect 7532 34024 7566 34055
rect 7532 34021 7566 34024
rect 7532 33955 7566 33982
rect 7532 33948 7566 33955
rect 7532 33886 7566 33909
rect 7532 33875 7566 33886
rect 7532 33817 7566 33836
rect 7532 33802 7566 33817
rect 7532 33748 7566 33763
rect 7532 33729 7566 33748
rect 7532 33679 7566 33690
rect 7532 33656 7566 33679
rect 7532 33610 7566 33617
rect 7532 33583 7566 33610
rect 7532 33541 7566 33544
rect 7532 33510 7566 33541
rect 7532 33438 7566 33471
rect 7532 33437 7566 33438
rect 7532 33369 7566 33398
rect 7532 33364 7566 33369
rect 7532 33300 7566 33325
rect 7532 33291 7566 33300
rect 7532 33231 7566 33252
rect 7532 33218 7566 33231
rect 7532 33162 7566 33179
rect 7532 33145 7566 33162
rect 7532 33093 7566 33106
rect 7532 33072 7566 33093
rect 7532 33024 7566 33033
rect 7532 32999 7566 33024
rect 7532 32955 7566 32960
rect 7532 32926 7566 32955
rect 7532 32886 7566 32887
rect 7532 32853 7566 32886
rect 7532 32782 7566 32814
rect 7532 32780 7566 32782
rect 7532 32713 7566 32741
rect 7532 32707 7566 32713
rect 8000 39444 8002 39454
rect 8002 39444 8034 39454
rect 8000 39420 8034 39444
rect 8000 39376 8002 39382
rect 8002 39376 8034 39382
rect 8000 39348 8034 39376
rect 8000 39308 8002 39310
rect 8002 39308 8034 39310
rect 8000 39276 8034 39308
rect 8000 39206 8034 39238
rect 8000 39204 8002 39206
rect 8002 39204 8034 39206
rect 8000 39138 8034 39166
rect 8000 39132 8002 39138
rect 8002 39132 8034 39138
rect 8000 39070 8034 39094
rect 8000 39060 8002 39070
rect 8002 39060 8034 39070
rect 8000 39002 8034 39022
rect 8000 38988 8002 39002
rect 8002 38988 8034 39002
rect 8000 38934 8034 38950
rect 8000 38916 8002 38934
rect 8002 38916 8034 38934
rect 8000 38866 8034 38878
rect 8000 38844 8002 38866
rect 8002 38844 8034 38866
rect 8000 38798 8034 38806
rect 8000 38772 8002 38798
rect 8002 38772 8034 38798
rect 8000 38730 8034 38734
rect 8000 38700 8002 38730
rect 8002 38700 8034 38730
rect 8000 38628 8002 38662
rect 8002 38628 8034 38662
rect 8000 38560 8002 38590
rect 8002 38560 8034 38590
rect 8000 38556 8034 38560
rect 8000 38492 8002 38518
rect 8002 38492 8034 38518
rect 8000 38484 8034 38492
rect 8000 38424 8002 38446
rect 8002 38424 8034 38446
rect 8000 38412 8034 38424
rect 8000 38356 8002 38374
rect 8002 38356 8034 38374
rect 8000 38340 8034 38356
rect 8000 38288 8002 38302
rect 8002 38288 8034 38302
rect 8000 38268 8034 38288
rect 8000 38220 8002 38230
rect 8002 38220 8034 38230
rect 8000 38196 8034 38220
rect 8000 38152 8002 38158
rect 8002 38152 8034 38158
rect 8000 38124 8034 38152
rect 8000 38084 8002 38086
rect 8002 38084 8034 38086
rect 8000 38052 8034 38084
rect 8000 37982 8034 38014
rect 8000 37980 8002 37982
rect 8002 37980 8034 37982
rect 8000 37914 8034 37942
rect 8000 37908 8002 37914
rect 8002 37908 8034 37914
rect 8000 37846 8034 37870
rect 8000 37836 8002 37846
rect 8002 37836 8034 37846
rect 8000 37778 8034 37798
rect 8000 37764 8002 37778
rect 8002 37764 8034 37778
rect 8000 37710 8034 37726
rect 8000 37692 8002 37710
rect 8002 37692 8034 37710
rect 8000 37642 8034 37654
rect 8000 37620 8002 37642
rect 8002 37620 8034 37642
rect 8000 37574 8034 37582
rect 8000 37548 8002 37574
rect 8002 37548 8034 37574
rect 8000 37506 8034 37510
rect 8000 37476 8002 37506
rect 8002 37476 8034 37506
rect 8000 37404 8002 37438
rect 8002 37404 8034 37438
rect 8000 37336 8002 37366
rect 8002 37336 8034 37366
rect 8000 37332 8034 37336
rect 8000 37268 8002 37294
rect 8002 37268 8034 37294
rect 8000 37260 8034 37268
rect 8000 37200 8002 37222
rect 8002 37200 8034 37222
rect 8000 37188 8034 37200
rect 8000 37132 8002 37150
rect 8002 37132 8034 37150
rect 8000 37116 8034 37132
rect 8000 37064 8002 37078
rect 8002 37064 8034 37078
rect 8000 37044 8034 37064
rect 8000 36996 8002 37006
rect 8002 36996 8034 37006
rect 8000 36972 8034 36996
rect 8000 36928 8002 36934
rect 8002 36928 8034 36934
rect 8000 36900 8034 36928
rect 8000 36860 8002 36862
rect 8002 36860 8034 36862
rect 8000 36828 8034 36860
rect 8000 36758 8034 36790
rect 8000 36756 8002 36758
rect 8002 36756 8034 36758
rect 8000 36690 8034 36718
rect 8000 36684 8002 36690
rect 8002 36684 8034 36690
rect 8000 36622 8034 36646
rect 8000 36612 8002 36622
rect 8002 36612 8034 36622
rect 8000 36554 8034 36574
rect 8000 36540 8002 36554
rect 8002 36540 8034 36554
rect 8000 36486 8034 36502
rect 8000 36468 8002 36486
rect 8002 36468 8034 36486
rect 8000 36418 8034 36430
rect 8000 36396 8002 36418
rect 8002 36396 8034 36418
rect 8000 36350 8034 36358
rect 8000 36324 8002 36350
rect 8002 36324 8034 36350
rect 8000 36282 8034 36286
rect 8000 36252 8002 36282
rect 8002 36252 8034 36282
rect 8000 36180 8002 36214
rect 8002 36180 8034 36214
rect 8000 36112 8002 36142
rect 8002 36112 8034 36142
rect 8000 36108 8034 36112
rect 8000 36044 8002 36070
rect 8002 36044 8034 36070
rect 8000 36036 8034 36044
rect 8000 35976 8002 35998
rect 8002 35976 8034 35998
rect 8000 35964 8034 35976
rect 8000 35908 8002 35926
rect 8002 35908 8034 35926
rect 8000 35892 8034 35908
rect 8000 35840 8002 35854
rect 8002 35840 8034 35854
rect 8000 35820 8034 35840
rect 8000 35772 8002 35782
rect 8002 35772 8034 35782
rect 8000 35748 8034 35772
rect 8000 35704 8002 35710
rect 8002 35704 8034 35710
rect 8000 35676 8034 35704
rect 8000 35636 8002 35638
rect 8002 35636 8034 35638
rect 8000 35604 8034 35636
rect 8000 35534 8034 35566
rect 8000 35532 8002 35534
rect 8002 35532 8034 35534
rect 8000 35466 8034 35494
rect 8000 35460 8002 35466
rect 8002 35460 8034 35466
rect 8000 35398 8034 35422
rect 8000 35388 8002 35398
rect 8002 35388 8034 35398
rect 8000 35330 8034 35350
rect 8000 35316 8002 35330
rect 8002 35316 8034 35330
rect 8000 35262 8034 35278
rect 8000 35244 8002 35262
rect 8002 35244 8034 35262
rect 8000 35194 8034 35206
rect 8000 35172 8002 35194
rect 8002 35172 8034 35194
rect 8000 35126 8034 35134
rect 8000 35100 8002 35126
rect 8002 35100 8034 35126
rect 8000 35058 8034 35062
rect 8000 35028 8002 35058
rect 8002 35028 8034 35058
rect 8000 34956 8002 34990
rect 8002 34956 8034 34990
rect 8000 34888 8002 34918
rect 8002 34888 8034 34918
rect 8000 34884 8034 34888
rect 8000 34820 8002 34846
rect 8002 34820 8034 34846
rect 8000 34812 8034 34820
rect 8000 34752 8002 34774
rect 8002 34752 8034 34774
rect 8000 34740 8034 34752
rect 8000 34684 8002 34702
rect 8002 34684 8034 34702
rect 8000 34668 8034 34684
rect 8000 34616 8002 34630
rect 8002 34616 8034 34630
rect 8000 34596 8034 34616
rect 8000 34548 8002 34558
rect 8002 34548 8034 34558
rect 8000 34524 8034 34548
rect 8000 34480 8002 34486
rect 8002 34480 8034 34486
rect 8000 34452 8034 34480
rect 8000 34412 8002 34414
rect 8002 34412 8034 34414
rect 8000 34380 8034 34412
rect 8000 34310 8034 34342
rect 8000 34308 8002 34310
rect 8002 34308 8034 34310
rect 8000 34242 8034 34270
rect 8000 34236 8002 34242
rect 8002 34236 8034 34242
rect 8000 34174 8034 34198
rect 8000 34164 8002 34174
rect 8002 34164 8034 34174
rect 8000 34106 8034 34126
rect 8000 34092 8002 34106
rect 8002 34092 8034 34106
rect 8000 34038 8034 34054
rect 8000 34020 8002 34038
rect 8002 34020 8034 34038
rect 8000 33970 8034 33982
rect 8000 33948 8002 33970
rect 8002 33948 8034 33970
rect 8000 33902 8034 33910
rect 8000 33876 8002 33902
rect 8002 33876 8034 33902
rect 8000 33834 8034 33838
rect 8000 33804 8002 33834
rect 8002 33804 8034 33834
rect 8000 33732 8002 33766
rect 8002 33732 8034 33766
rect 8000 33664 8002 33694
rect 8002 33664 8034 33694
rect 8000 33660 8034 33664
rect 8000 33596 8002 33622
rect 8002 33596 8034 33622
rect 8000 33588 8034 33596
rect 8000 33528 8002 33550
rect 8002 33528 8034 33550
rect 8000 33516 8034 33528
rect 8000 33460 8002 33478
rect 8002 33460 8034 33478
rect 8000 33444 8034 33460
rect 8000 33392 8002 33406
rect 8002 33392 8034 33406
rect 8000 33372 8034 33392
rect 8000 33324 8002 33334
rect 8002 33324 8034 33334
rect 8000 33300 8034 33324
rect 8000 33256 8002 33262
rect 8002 33256 8034 33262
rect 8000 33228 8034 33256
rect 8000 33188 8002 33190
rect 8002 33188 8034 33190
rect 8000 33156 8034 33188
rect 8000 33086 8034 33118
rect 8000 33084 8002 33086
rect 8002 33084 8034 33086
rect 8000 33018 8034 33046
rect 8000 33012 8002 33018
rect 8002 33012 8034 33018
rect 8000 32950 8034 32974
rect 8000 32940 8002 32950
rect 8002 32940 8034 32950
rect 8000 32882 8034 32902
rect 8000 32868 8002 32882
rect 8002 32868 8034 32882
rect 8000 32814 8034 32830
rect 8000 32796 8002 32814
rect 8002 32796 8034 32814
rect 8000 32746 8034 32758
rect 8000 32724 8002 32746
rect 8002 32724 8034 32746
rect 8000 32678 8034 32686
rect 8000 32652 8002 32678
rect 8002 32652 8034 32678
rect 8000 32610 8034 32614
rect 7532 32522 7566 32539
rect 7532 32505 7566 32522
rect 7532 32453 7566 32467
rect 7532 32433 7566 32453
rect 7532 32384 7566 32395
rect 7532 32361 7566 32384
rect 7532 32315 7566 32323
rect 7532 32289 7566 32315
rect 7532 32246 7566 32251
rect 7532 32217 7566 32246
rect 7532 32177 7566 32179
rect 7532 32145 7566 32177
rect 7532 32074 7566 32107
rect 7532 32073 7566 32074
rect 7532 32005 7566 32035
rect 7532 32001 7566 32005
rect 7532 31936 7566 31963
rect 7532 31929 7566 31936
rect 7532 31867 7566 31891
rect 7532 31857 7566 31867
rect 7532 31798 7566 31819
rect 7532 31785 7566 31798
rect 7532 31729 7566 31747
rect 7532 31713 7566 31729
rect 7532 31659 7566 31675
rect 7532 31641 7566 31659
rect 7532 31589 7566 31603
rect 7532 31569 7566 31589
rect 7532 31519 7566 31531
rect 7532 31497 7566 31519
rect 7532 31449 7566 31459
rect 7532 31425 7566 31449
rect 7532 31379 7566 31387
rect 7532 31353 7566 31379
rect 7532 31309 7566 31315
rect 7532 31281 7566 31309
rect 7532 31239 7566 31243
rect 7532 31209 7566 31239
rect 7532 31169 7566 31171
rect 7532 31137 7566 31169
rect 7532 31065 7566 31099
rect 7532 30993 7566 31026
rect 7532 30992 7566 30993
rect 7532 30923 7566 30953
rect 7532 30919 7566 30923
rect 7532 30853 7566 30880
rect 7532 30846 7566 30853
rect 7532 30783 7566 30807
rect 7532 30773 7566 30783
rect 7532 30713 7566 30734
rect 7532 30700 7566 30713
rect 7532 30643 7566 30661
rect 7532 30627 7566 30643
rect 7532 30573 7566 30588
rect 7532 30554 7566 30573
rect 7532 30503 7566 30515
rect 7532 30481 7566 30503
rect 7532 30433 7566 30442
rect 7532 30408 7566 30433
rect 8000 32580 8002 32610
rect 8002 32580 8034 32610
rect 8000 32508 8002 32542
rect 8002 32508 8034 32542
rect 8000 32440 8002 32470
rect 8002 32440 8034 32470
rect 8000 32436 8034 32440
rect 8000 32372 8002 32398
rect 8002 32372 8034 32398
rect 8000 32364 8034 32372
rect 8000 32304 8002 32326
rect 8002 32304 8034 32326
rect 8000 32292 8034 32304
rect 8000 32236 8002 32254
rect 8002 32236 8034 32254
rect 8000 32220 8034 32236
rect 8000 32168 8002 32182
rect 8002 32168 8034 32182
rect 8000 32148 8034 32168
rect 8000 32100 8002 32110
rect 8002 32100 8034 32110
rect 8000 32076 8034 32100
rect 8000 32032 8002 32038
rect 8002 32032 8034 32038
rect 8000 32004 8034 32032
rect 8000 31964 8002 31966
rect 8002 31964 8034 31966
rect 8000 31932 8034 31964
rect 8000 31862 8034 31894
rect 8000 31860 8002 31862
rect 8002 31860 8034 31862
rect 8000 31794 8034 31822
rect 8000 31788 8002 31794
rect 8002 31788 8034 31794
rect 8000 31726 8034 31750
rect 8000 31716 8002 31726
rect 8002 31716 8034 31726
rect 8000 31658 8034 31678
rect 8000 31644 8002 31658
rect 8002 31644 8034 31658
rect 8000 31590 8034 31606
rect 8000 31572 8002 31590
rect 8002 31572 8034 31590
rect 8000 31522 8034 31534
rect 8000 31500 8002 31522
rect 8002 31500 8034 31522
rect 8000 31454 8034 31462
rect 8000 31428 8002 31454
rect 8002 31428 8034 31454
rect 8000 31386 8034 31390
rect 8000 31356 8002 31386
rect 8002 31356 8034 31386
rect 8000 31284 8002 31318
rect 8002 31284 8034 31318
rect 8000 31216 8002 31246
rect 8002 31216 8034 31246
rect 8000 31212 8034 31216
rect 8000 31148 8002 31174
rect 8002 31148 8034 31174
rect 8000 31140 8034 31148
rect 8000 31080 8002 31102
rect 8002 31080 8034 31102
rect 8000 31068 8034 31080
rect 8000 31012 8002 31030
rect 8002 31012 8034 31030
rect 8000 30996 8034 31012
rect 8000 30944 8002 30958
rect 8002 30944 8034 30958
rect 8000 30924 8034 30944
rect 8000 30876 8002 30886
rect 8002 30876 8034 30886
rect 8000 30852 8034 30876
rect 8000 30808 8002 30814
rect 8002 30808 8034 30814
rect 8000 30780 8034 30808
rect 8000 30740 8002 30742
rect 8002 30740 8034 30742
rect 8000 30708 8034 30740
rect 8000 30638 8034 30670
rect 8000 30636 8002 30638
rect 8002 30636 8034 30638
rect 8000 30570 8034 30598
rect 8000 30564 8002 30570
rect 8002 30564 8034 30570
rect 8000 30502 8034 30526
rect 8000 30492 8002 30502
rect 8002 30492 8034 30502
rect 8000 30434 8034 30454
rect 8000 30420 8002 30434
rect 8002 30420 8034 30434
rect 8000 30366 8034 30382
rect 8000 30348 8002 30366
rect 8002 30348 8034 30366
rect 8000 30298 8034 30310
rect 8000 30276 8002 30298
rect 8002 30276 8034 30298
rect 8000 30230 8034 30238
rect 8000 30204 8002 30230
rect 8002 30204 8034 30230
rect 8000 30162 8034 30166
rect 8000 30132 8002 30162
rect 8002 30132 8034 30162
rect 8000 30060 8002 30094
rect 8002 30060 8034 30094
rect 8000 29992 8002 30022
rect 8002 29992 8034 30022
rect 8000 29988 8034 29992
rect 8000 29924 8002 29950
rect 8002 29924 8034 29950
rect 8000 29916 8034 29924
rect 6781 29854 6804 29888
rect 6804 29854 6815 29888
rect 6853 29854 6872 29888
rect 6872 29854 6887 29888
rect 7013 29854 7028 29888
rect 7028 29854 7047 29888
rect 7085 29854 7096 29888
rect 7096 29854 7119 29888
rect 8000 29856 8002 29878
rect 8002 29856 8034 29878
rect 8000 29844 8034 29856
rect 8000 29788 8002 29806
rect 8002 29788 8034 29806
rect 8000 29772 8034 29788
rect 8000 29720 8002 29734
rect 8002 29720 8034 29734
rect 8000 29700 8034 29720
rect 8000 29652 8002 29662
rect 8002 29652 8034 29662
rect 8000 29628 8034 29652
rect 8000 29584 8002 29590
rect 8002 29584 8034 29590
rect 5850 29532 5854 29565
rect 5854 29532 5884 29565
rect 5923 29532 5924 29565
rect 5924 29532 5957 29565
rect 5996 29532 6028 29565
rect 6028 29532 6030 29565
rect 6069 29532 6098 29565
rect 6098 29532 6103 29565
rect 6142 29532 6168 29565
rect 6168 29532 6176 29565
rect 6215 29532 6238 29565
rect 6238 29532 6249 29565
rect 6288 29532 6308 29565
rect 6308 29532 6322 29565
rect 6361 29532 6378 29565
rect 6378 29532 6395 29565
rect 6434 29532 6448 29565
rect 6448 29532 6468 29565
rect 6507 29532 6518 29565
rect 6518 29532 6541 29565
rect 6579 29532 6588 29565
rect 6588 29532 6613 29565
rect 6651 29532 6658 29565
rect 6658 29532 6685 29565
rect 6723 29532 6728 29565
rect 6728 29532 6757 29565
rect 6795 29532 6798 29565
rect 6798 29532 6829 29565
rect 6867 29532 6868 29565
rect 6868 29532 6901 29565
rect 5850 29531 5884 29532
rect 5923 29531 5957 29532
rect 5996 29531 6030 29532
rect 6069 29531 6103 29532
rect 6142 29531 6176 29532
rect 6215 29531 6249 29532
rect 6288 29531 6322 29532
rect 6361 29531 6395 29532
rect 6434 29531 6468 29532
rect 6507 29531 6541 29532
rect 6579 29531 6613 29532
rect 6651 29531 6685 29532
rect 6723 29531 6757 29532
rect 6795 29531 6829 29532
rect 6867 29531 6901 29532
rect 6939 29531 6973 29565
rect 7011 29532 7043 29565
rect 7043 29532 7045 29565
rect 7083 29532 7112 29565
rect 7112 29532 7117 29565
rect 7155 29532 7181 29565
rect 7181 29532 7189 29565
rect 7227 29532 7250 29565
rect 7250 29532 7261 29565
rect 7299 29532 7319 29565
rect 7319 29532 7333 29565
rect 7371 29532 7388 29565
rect 7388 29532 7405 29565
rect 7011 29531 7045 29532
rect 7083 29531 7117 29532
rect 7155 29531 7189 29532
rect 7227 29531 7261 29532
rect 7299 29531 7333 29532
rect 7371 29531 7405 29532
rect 7443 29531 7477 29565
rect 8000 29556 8034 29584
rect 8000 29516 8002 29518
rect 8002 29516 8034 29518
rect 8000 29484 8034 29516
rect 8000 29414 8034 29446
rect 8000 29412 8002 29414
rect 8002 29412 8034 29414
rect 8000 29346 8034 29374
rect 8000 29340 8002 29346
rect 8002 29340 8034 29346
rect 8000 29278 8034 29302
rect 8000 29268 8002 29278
rect 8002 29268 8034 29278
rect 8000 29210 8034 29230
rect 8000 29196 8002 29210
rect 8002 29196 8034 29210
rect 5939 29160 5954 29194
rect 5954 29160 5973 29194
rect 6020 29160 6028 29194
rect 6028 29160 6054 29194
rect 6101 29160 6102 29194
rect 6102 29160 6135 29194
rect 6182 29160 6210 29194
rect 6210 29160 6216 29194
rect 6263 29160 6283 29194
rect 6283 29160 6297 29194
rect 6344 29160 6356 29194
rect 6356 29160 6378 29194
rect 6425 29160 6429 29194
rect 6429 29160 6459 29194
rect 6505 29160 6539 29194
rect 6585 29160 6614 29194
rect 6614 29160 6619 29194
rect 6946 29160 6950 29194
rect 6950 29160 6980 29194
rect 7018 29160 7052 29194
rect 7314 29160 7316 29194
rect 7316 29160 7348 29194
rect 7386 29160 7418 29194
rect 7418 29160 7420 29194
rect 8000 29142 8034 29158
rect 8000 29124 8002 29142
rect 8002 29124 8034 29142
rect 8000 29074 8034 29086
rect 8000 29052 8002 29074
rect 8002 29052 8034 29074
rect 8000 29006 8034 29014
rect 8000 28980 8002 29006
rect 8002 28980 8034 29006
rect 8000 28938 8034 28942
rect 8000 28908 8002 28938
rect 8002 28908 8034 28938
rect 8000 28836 8002 28870
rect 8002 28836 8034 28870
rect 5939 28788 5954 28822
rect 5954 28788 5973 28822
rect 6020 28788 6028 28822
rect 6028 28788 6054 28822
rect 6101 28788 6102 28822
rect 6102 28788 6135 28822
rect 6182 28788 6210 28822
rect 6210 28788 6216 28822
rect 6263 28788 6283 28822
rect 6283 28788 6297 28822
rect 6344 28788 6356 28822
rect 6356 28788 6378 28822
rect 6425 28788 6429 28822
rect 6429 28788 6459 28822
rect 6505 28788 6539 28822
rect 6585 28788 6614 28822
rect 6614 28788 6619 28822
rect 6946 28788 6950 28822
rect 6950 28788 6980 28822
rect 7018 28788 7052 28822
rect 8000 28768 8002 28798
rect 8002 28768 8034 28798
rect 8000 28764 8034 28768
rect 8000 28700 8002 28726
rect 8002 28700 8034 28726
rect 8000 28692 8034 28700
rect 8000 28632 8002 28654
rect 8002 28632 8034 28654
rect 8000 28620 8034 28632
rect 8000 28564 8002 28582
rect 8002 28564 8034 28582
rect 8000 28548 8034 28564
rect 8000 28496 8002 28510
rect 8002 28496 8034 28510
rect 8000 28476 8034 28496
rect 8000 28428 8002 28438
rect 8002 28428 8034 28438
rect 5867 28390 5873 28424
rect 5873 28390 5901 28424
rect 5943 28390 5944 28424
rect 5944 28390 5977 28424
rect 6019 28390 6049 28424
rect 6049 28390 6053 28424
rect 6095 28390 6120 28424
rect 6120 28390 6129 28424
rect 6171 28390 6191 28424
rect 6191 28390 6205 28424
rect 6246 28390 6262 28424
rect 6262 28390 6280 28424
rect 6321 28390 6333 28424
rect 6333 28390 6355 28424
rect 6396 28390 6404 28424
rect 6404 28390 6430 28424
rect 6471 28390 6475 28424
rect 6475 28390 6505 28424
rect 6546 28390 6580 28424
rect 6621 28390 6654 28424
rect 6654 28390 6655 28424
rect 6696 28390 6725 28424
rect 6725 28390 6730 28424
rect 6771 28390 6796 28424
rect 6796 28390 6805 28424
rect 6846 28390 6867 28424
rect 6867 28390 6880 28424
rect 6921 28390 6937 28424
rect 6937 28390 6955 28424
rect 6996 28390 7007 28424
rect 7007 28390 7030 28424
rect 7071 28390 7077 28424
rect 7077 28390 7105 28424
rect 7146 28390 7147 28424
rect 7147 28390 7180 28424
rect 7221 28390 7251 28424
rect 7251 28390 7255 28424
rect 7296 28390 7321 28424
rect 7321 28390 7330 28424
rect 7371 28390 7391 28424
rect 7391 28390 7405 28424
rect 8000 28404 8034 28428
rect 8000 28360 8002 28366
rect 8002 28360 8034 28366
rect 8000 28332 8034 28360
rect 8000 28292 8002 28294
rect 8002 28292 8034 28294
rect 8000 28260 8034 28292
rect 8000 28190 8034 28222
rect 8000 28188 8002 28190
rect 8002 28188 8034 28190
rect 8000 28122 8034 28150
rect 8000 28116 8002 28122
rect 8002 28116 8034 28122
rect 8000 28054 8034 28078
rect 8000 28044 8002 28054
rect 8002 28044 8034 28054
rect 8000 27986 8034 28006
rect 8000 27972 8002 27986
rect 8002 27972 8034 27986
rect 8000 27918 8034 27934
rect 8000 27900 8002 27918
rect 8002 27900 8034 27918
rect 8000 27850 8034 27862
rect 8000 27828 8002 27850
rect 8002 27828 8034 27850
rect 8000 27782 8034 27790
rect 8000 27756 8002 27782
rect 8002 27756 8034 27782
rect 8000 27714 8034 27718
rect 8000 27684 8002 27714
rect 8002 27684 8034 27714
rect 8000 27612 8002 27646
rect 8002 27612 8034 27646
rect 8000 27544 8002 27574
rect 8002 27544 8034 27574
rect 8000 27540 8034 27544
rect 8000 27476 8002 27502
rect 8002 27476 8034 27502
rect 8000 27468 8034 27476
rect 8000 27408 8002 27430
rect 8002 27408 8034 27430
rect 8000 27396 8034 27408
rect 8000 27340 8002 27358
rect 8002 27340 8034 27358
rect 8000 27324 8034 27340
rect 8000 27272 8002 27286
rect 8002 27272 8034 27286
rect 8000 27252 8034 27272
rect 8000 27204 8002 27214
rect 8002 27204 8034 27214
rect 8000 27180 8034 27204
rect 8000 27136 8002 27142
rect 8002 27136 8034 27142
rect 2825 27092 2859 27126
rect 2825 27020 2859 27054
rect 5929 27054 5963 27088
rect 6071 27060 6104 27088
rect 6104 27060 6105 27088
rect 6071 27054 6105 27060
rect 6485 27012 6591 27118
rect 8000 27108 8034 27136
rect 6843 26985 6949 27091
rect 7318 26974 7424 27080
rect 7682 26974 7788 27080
rect 8000 27068 8002 27070
rect 8002 27068 8034 27070
rect 8000 27036 8034 27068
rect 8000 26966 8034 26998
rect 8000 26964 8002 26966
rect 8002 26964 8034 26966
rect 8000 26898 8034 26926
rect 8000 26892 8002 26898
rect 8002 26892 8034 26898
rect 8000 26830 8034 26854
rect 8000 26820 8002 26830
rect 8002 26820 8034 26830
rect 8000 26762 8034 26782
rect 8000 26748 8002 26762
rect 8002 26748 8034 26762
rect 8000 26694 8034 26710
rect 8000 26676 8002 26694
rect 8002 26676 8034 26694
rect 8000 26626 8034 26638
rect 8000 26604 8002 26626
rect 8002 26604 8034 26626
rect 8000 26558 8034 26566
rect 8000 26532 8002 26558
rect 8002 26532 8034 26558
rect 8000 26490 8034 26494
rect 8000 26460 8002 26490
rect 8002 26460 8034 26490
rect 8000 26388 8002 26422
rect 8002 26388 8034 26422
rect 8000 26320 8002 26350
rect 8002 26320 8034 26350
rect 8000 26316 8034 26320
rect 8000 26252 8002 26278
rect 8002 26252 8034 26278
rect 8000 26244 8034 26252
rect 8000 26184 8002 26206
rect 8002 26184 8034 26206
rect 8000 26172 8034 26184
rect 8000 26116 8002 26134
rect 8002 26116 8034 26134
rect 8000 26100 8034 26116
rect 8000 26048 8002 26062
rect 8002 26048 8034 26062
rect 8000 26028 8034 26048
rect 8000 25980 8002 25990
rect 8002 25980 8034 25990
rect 8000 25956 8034 25980
rect 8000 25912 8002 25918
rect 8002 25912 8034 25918
rect 8000 25884 8034 25912
rect 8000 25844 8002 25846
rect 8002 25844 8034 25846
rect 8000 25812 8034 25844
rect 8000 25742 8034 25774
rect 8000 25740 8002 25742
rect 8002 25740 8034 25742
rect 8000 25674 8034 25702
rect 8000 25668 8002 25674
rect 8002 25668 8034 25674
rect 8000 25606 8034 25630
rect 8000 25596 8002 25606
rect 8002 25596 8034 25606
rect 8000 25538 8034 25558
rect 8000 25524 8002 25538
rect 8002 25524 8034 25538
rect 8000 25470 8034 25486
rect 8000 25452 8002 25470
rect 8002 25452 8034 25470
rect 8000 25402 8034 25414
rect 8000 25380 8002 25402
rect 8002 25380 8034 25402
rect 8000 25334 8034 25342
rect 8000 25308 8002 25334
rect 8002 25308 8034 25334
rect 8000 25266 8034 25270
rect 8000 25236 8002 25266
rect 8002 25236 8034 25266
rect 8000 25164 8002 25198
rect 8002 25164 8034 25198
rect 8000 25096 8002 25126
rect 8002 25096 8034 25126
rect 8000 25092 8034 25096
rect 8000 25028 8002 25054
rect 8002 25028 8034 25054
rect 8000 25020 8034 25028
rect 8000 24960 8002 24982
rect 8002 24960 8034 24982
rect 8000 24948 8034 24960
rect 8000 24892 8002 24910
rect 8002 24892 8034 24910
rect 8000 24876 8034 24892
rect 8000 24824 8002 24838
rect 8002 24824 8034 24838
rect 8000 24804 8034 24824
rect 8000 24756 8002 24766
rect 8002 24756 8034 24766
rect 8000 24732 8034 24756
rect 8000 24688 8002 24694
rect 8002 24688 8034 24694
rect 8000 24660 8034 24688
rect 8000 24620 8002 24622
rect 8002 24620 8034 24622
rect 8000 24588 8034 24620
rect 8000 24518 8034 24550
rect 8000 24516 8002 24518
rect 8002 24516 8034 24518
rect 8000 24450 8034 24478
rect 8000 24444 8002 24450
rect 8002 24444 8034 24450
rect 8000 24382 8034 24406
rect 8000 24372 8002 24382
rect 8002 24372 8034 24382
rect 8000 24314 8034 24334
rect 8000 24300 8002 24314
rect 8002 24300 8034 24314
rect 8000 24246 8034 24262
rect 8000 24228 8002 24246
rect 8002 24228 8034 24246
rect 8000 24178 8034 24190
rect 8000 24156 8002 24178
rect 8002 24156 8034 24178
rect 8000 24110 8034 24118
rect 8000 24084 8002 24110
rect 8002 24084 8034 24110
rect 8000 24042 8034 24046
rect 8000 24012 8002 24042
rect 8002 24012 8034 24042
rect 8000 23940 8002 23974
rect 8002 23940 8034 23974
rect 8000 23872 8002 23902
rect 8002 23872 8034 23902
rect 8000 23868 8034 23872
rect 8000 23804 8002 23830
rect 8002 23804 8034 23830
rect 8000 23796 8034 23804
rect 8000 23736 8002 23758
rect 8002 23736 8034 23758
rect 8000 23724 8034 23736
rect 8000 23668 8002 23686
rect 8002 23668 8034 23686
rect 8000 23652 8034 23668
rect 8000 23600 8002 23614
rect 8002 23600 8034 23614
rect 8000 23580 8034 23600
rect 8000 23532 8002 23542
rect 8002 23532 8034 23542
rect 8000 23508 8034 23532
rect 8000 23464 8002 23470
rect 8002 23464 8034 23470
rect 8000 23436 8034 23464
rect 8000 23396 8002 23398
rect 8002 23396 8034 23398
rect 8000 23364 8034 23396
rect 8000 23294 8034 23326
rect 8000 23292 8002 23294
rect 8002 23292 8034 23294
rect 8000 23226 8034 23254
rect 8000 23220 8002 23226
rect 8002 23220 8034 23226
rect 8000 23158 8034 23182
rect 8000 23148 8002 23158
rect 8002 23148 8034 23158
rect 8000 23090 8034 23110
rect 8000 23076 8002 23090
rect 8002 23076 8034 23090
rect 8000 23022 8034 23038
rect 8000 23004 8002 23022
rect 8002 23004 8034 23022
rect 8000 22954 8034 22966
rect 8000 22932 8002 22954
rect 8002 22932 8034 22954
rect 8000 22886 8034 22894
rect 8000 22860 8002 22886
rect 8002 22860 8034 22886
rect 8000 22818 8034 22822
rect 8000 22788 8002 22818
rect 8002 22788 8034 22818
rect 8000 22716 8002 22750
rect 8002 22716 8034 22750
rect 8000 22648 8002 22678
rect 8002 22648 8034 22678
rect 8000 22644 8034 22648
rect 8000 22580 8002 22606
rect 8002 22580 8034 22606
rect 8000 22572 8034 22580
rect 8000 22512 8002 22534
rect 8002 22512 8034 22534
rect 8000 22500 8034 22512
rect 8000 22444 8002 22462
rect 8002 22444 8034 22462
rect 8000 22428 8034 22444
rect 8000 22376 8002 22390
rect 8002 22376 8034 22390
rect 8000 22356 8034 22376
rect 8000 22308 8002 22318
rect 8002 22308 8034 22318
rect 8000 22284 8034 22308
rect 8000 22240 8002 22246
rect 8002 22240 8034 22246
rect 8000 22212 8034 22240
rect 8000 22172 8002 22174
rect 8002 22172 8034 22174
rect 8000 22140 8034 22172
rect 6442 22085 6476 22119
rect 6517 22085 6520 22119
rect 6520 22085 6551 22119
rect 6592 22085 6622 22119
rect 6622 22085 6626 22119
rect 6667 22085 6690 22119
rect 6690 22085 6701 22119
rect 6742 22085 6758 22119
rect 6758 22085 6776 22119
rect 8000 22070 8034 22102
rect 8000 22068 8002 22070
rect 8002 22068 8034 22070
rect 8000 22002 8034 22030
rect 8000 21996 8002 22002
rect 8002 21996 8034 22002
rect 8000 21934 8034 21958
rect 8000 21924 8002 21934
rect 8002 21924 8034 21934
rect 8000 21866 8034 21886
rect 8000 21852 8002 21866
rect 8002 21852 8034 21866
rect 8000 21798 8034 21814
rect 8000 21780 8002 21798
rect 8002 21780 8034 21798
rect 8000 21730 8034 21742
rect 8000 21708 8002 21730
rect 8002 21708 8034 21730
rect 8000 21662 8034 21670
rect 8000 21636 8002 21662
rect 8002 21636 8034 21662
rect 6442 21570 6463 21604
rect 6463 21570 6476 21604
rect 6514 21570 6531 21604
rect 6531 21570 6548 21604
rect 6672 21570 6687 21604
rect 6687 21570 6706 21604
rect 6744 21570 6755 21604
rect 6755 21570 6778 21604
rect 8000 21594 8034 21598
rect 8000 21564 8002 21594
rect 8002 21564 8034 21594
rect 8000 21492 8002 21526
rect 8002 21492 8034 21526
rect 8000 21424 8002 21454
rect 8002 21424 8034 21454
rect 8000 21420 8034 21424
rect 8000 21356 8002 21382
rect 8002 21356 8034 21382
rect 8000 21348 8034 21356
rect 8000 21288 8002 21310
rect 8002 21288 8034 21310
rect 8000 21276 8034 21288
rect 8000 21220 8002 21238
rect 8002 21220 8034 21238
rect 8000 21204 8034 21220
rect 8000 21152 8002 21166
rect 8002 21152 8034 21166
rect 8000 21132 8034 21152
rect 8000 21084 8002 21094
rect 8002 21084 8034 21094
rect 8000 21060 8034 21084
rect 8000 21016 8002 21022
rect 8002 21016 8034 21022
rect 8000 20988 8034 21016
rect 8000 20948 8002 20950
rect 8002 20948 8034 20950
rect 8000 20916 8034 20948
rect 8000 20846 8034 20878
rect 8000 20844 8002 20846
rect 8002 20844 8034 20846
rect 8000 20778 8034 20806
rect 8000 20772 8002 20778
rect 8002 20772 8034 20778
rect 8000 20710 8034 20734
rect 8000 20700 8002 20710
rect 8002 20700 8034 20710
rect 8000 20642 8034 20662
rect 8000 20628 8002 20642
rect 8002 20628 8034 20642
rect 8000 20574 8034 20590
rect 8000 20556 8002 20574
rect 8002 20556 8034 20574
rect 8000 20506 8034 20518
rect 8000 20484 8002 20506
rect 8002 20484 8034 20506
rect 8000 20438 8034 20446
rect 8000 20412 8002 20438
rect 8002 20412 8034 20438
rect 8000 20370 8034 20374
rect 8000 20340 8002 20370
rect 8002 20340 8034 20370
rect 8000 20268 8002 20302
rect 8002 20268 8034 20302
rect 8000 20200 8002 20230
rect 8002 20200 8034 20230
rect 8000 20196 8034 20200
rect 8000 20132 8002 20158
rect 8002 20132 8034 20158
rect 8000 20124 8034 20132
rect 8000 20064 8002 20086
rect 8002 20064 8034 20086
rect 8000 20052 8034 20064
rect 8000 19996 8002 20014
rect 8002 19996 8034 20014
rect 8000 19980 8034 19996
rect 8000 19928 8002 19942
rect 8002 19928 8034 19942
rect 8000 19908 8034 19928
rect 8000 19860 8002 19870
rect 8002 19860 8034 19870
rect 8000 19836 8034 19860
rect 8000 19792 8002 19798
rect 8002 19792 8034 19798
rect 8000 19764 8034 19792
rect 8000 19724 8002 19726
rect 8002 19724 8034 19726
rect 8000 19692 8034 19724
rect 8000 19622 8034 19654
rect 8000 19620 8002 19622
rect 8002 19620 8034 19622
rect 8000 19554 8034 19582
rect 8000 19548 8002 19554
rect 8002 19548 8034 19554
rect 8000 19486 8034 19510
rect 8000 19476 8002 19486
rect 8002 19476 8034 19486
rect 8000 19418 8034 19438
rect 8000 19404 8002 19418
rect 8002 19404 8034 19418
rect 8000 19350 8034 19366
rect 8000 19332 8002 19350
rect 8002 19332 8034 19350
rect 8000 19282 8034 19294
rect 8000 19260 8002 19282
rect 8002 19260 8034 19282
rect 8000 19214 8034 19222
rect 8000 19188 8002 19214
rect 8002 19188 8034 19214
rect 8000 19146 8034 19150
rect 8000 19116 8002 19146
rect 8002 19116 8034 19146
rect 8000 19044 8002 19078
rect 8002 19044 8034 19078
rect 8000 18976 8002 19006
rect 8002 18976 8034 19006
rect 8000 18972 8034 18976
rect 8000 18908 8002 18934
rect 8002 18908 8034 18934
rect 8000 18900 8034 18908
rect 8000 18840 8002 18862
rect 8002 18840 8034 18862
rect 8000 18828 8034 18840
rect 8000 18772 8002 18790
rect 8002 18772 8034 18790
rect 8000 18756 8034 18772
rect 8000 18704 8002 18718
rect 8002 18704 8034 18718
rect 8000 18684 8034 18704
rect 8000 18636 8002 18646
rect 8002 18636 8034 18646
rect 8000 18612 8034 18636
rect 8000 18568 8002 18574
rect 8002 18568 8034 18574
rect 8000 18540 8034 18568
rect 8000 18500 8002 18502
rect 8002 18500 8034 18502
rect 8000 18468 8034 18500
rect 8000 18398 8034 18430
rect 8000 18396 8002 18398
rect 8002 18396 8034 18398
rect 8000 18330 8034 18358
rect 8000 18324 8002 18330
rect 8002 18324 8034 18330
rect 8000 18262 8034 18286
rect 8000 18252 8002 18262
rect 8002 18252 8034 18262
rect 8000 18194 8034 18214
rect 8000 18180 8002 18194
rect 8002 18180 8034 18194
rect 8000 18126 8034 18142
rect 8000 18108 8002 18126
rect 8002 18108 8034 18126
rect 8000 18058 8034 18070
rect 8000 18036 8002 18058
rect 8002 18036 8034 18058
rect 8000 17990 8034 17998
rect 8000 17964 8002 17990
rect 8002 17964 8034 17990
rect 8000 17922 8034 17926
rect 8000 17892 8002 17922
rect 8002 17892 8034 17922
rect 8000 17820 8002 17854
rect 8002 17820 8034 17854
rect 8000 17752 8002 17782
rect 8002 17752 8034 17782
rect 8000 17748 8034 17752
rect 8000 17684 8002 17710
rect 8002 17684 8034 17710
rect 8000 17676 8034 17684
rect 8000 17616 8002 17638
rect 8002 17616 8034 17638
rect 8000 17604 8034 17616
rect 8000 17548 8002 17566
rect 8002 17548 8034 17566
rect 8000 17532 8034 17548
rect 8000 17480 8002 17494
rect 8002 17480 8034 17494
rect 8000 17460 8034 17480
rect 8000 17412 8002 17422
rect 8002 17412 8034 17422
rect 8000 17388 8034 17412
rect 8000 17344 8002 17350
rect 8002 17344 8034 17350
rect 8000 17316 8034 17344
rect 8000 17276 8002 17278
rect 8002 17276 8034 17278
rect 8000 17244 8034 17276
rect 8000 17174 8034 17206
rect 8000 17172 8002 17174
rect 8002 17172 8034 17174
rect 8000 17106 8034 17134
rect 8000 17100 8002 17106
rect 8002 17100 8034 17106
rect 8000 17038 8034 17062
rect 8000 17028 8002 17038
rect 8002 17028 8034 17038
rect 8000 16970 8034 16990
rect 8000 16956 8002 16970
rect 8002 16956 8034 16970
rect 8000 16902 8034 16918
rect 8000 16884 8002 16902
rect 8002 16884 8034 16902
rect 8000 16834 8034 16846
rect 8000 16812 8002 16834
rect 8002 16812 8034 16834
rect 8000 16766 8034 16774
rect 8000 16740 8002 16766
rect 8002 16740 8034 16766
rect 8000 16698 8034 16702
rect 8000 16668 8002 16698
rect 8002 16668 8034 16698
rect 8000 16596 8002 16630
rect 8002 16596 8034 16630
rect 8000 16528 8002 16558
rect 8002 16528 8034 16558
rect 8000 16524 8034 16528
rect 8000 16460 8002 16486
rect 8002 16460 8034 16486
rect 8000 16452 8034 16460
rect 8000 16392 8002 16414
rect 8002 16392 8034 16414
rect 8000 16380 8034 16392
rect 8000 16324 8002 16342
rect 8002 16324 8034 16342
rect 8000 16308 8034 16324
rect 8000 16256 8002 16270
rect 8002 16256 8034 16270
rect 8000 16236 8034 16256
rect 8000 16188 8002 16198
rect 8002 16188 8034 16198
rect 8000 16164 8034 16188
rect 8000 16120 8002 16126
rect 8002 16120 8034 16126
rect 8000 16092 8034 16120
rect 8000 16052 8002 16054
rect 8002 16052 8034 16054
rect 8000 16020 8034 16052
rect 8000 15950 8034 15982
rect 8000 15948 8002 15950
rect 8002 15948 8034 15950
rect 8000 15882 8034 15910
rect 8000 15876 8002 15882
rect 8002 15876 8034 15882
rect 8000 15814 8034 15838
rect 8000 15804 8002 15814
rect 8002 15804 8034 15814
rect 8000 15746 8034 15766
rect 8000 15732 8002 15746
rect 8002 15732 8034 15746
rect 8000 15678 8034 15694
rect 8000 15660 8002 15678
rect 8002 15660 8034 15678
rect 8000 15610 8034 15622
rect 8000 15588 8002 15610
rect 8002 15588 8034 15610
rect 8000 15542 8034 15550
rect 8000 15516 8002 15542
rect 8002 15516 8034 15542
rect 8000 15474 8034 15478
rect 8000 15444 8002 15474
rect 8002 15444 8034 15474
rect 8000 15372 8002 15406
rect 8002 15372 8034 15406
rect 8000 15304 8002 15334
rect 8002 15304 8034 15334
rect 8000 15300 8034 15304
rect 8000 15236 8002 15262
rect 8002 15236 8034 15262
rect 8000 15228 8034 15236
rect 8000 15168 8002 15190
rect 8002 15168 8034 15190
rect 8000 15156 8034 15168
rect 8000 15100 8002 15118
rect 8002 15100 8034 15118
rect 8000 15084 8034 15100
rect 8000 15032 8002 15046
rect 8002 15032 8034 15046
rect 8000 15012 8034 15032
rect 8000 14964 8002 14974
rect 8002 14964 8034 14974
rect 8000 14940 8034 14964
rect 8000 14896 8002 14902
rect 8002 14896 8034 14902
rect 8000 14868 8034 14896
rect 8000 14828 8002 14830
rect 8002 14828 8034 14830
rect 8000 14796 8034 14828
rect 8000 14726 8034 14758
rect 8000 14724 8002 14726
rect 8002 14724 8034 14726
rect 8000 14658 8034 14686
rect 8000 14652 8002 14658
rect 8002 14652 8034 14658
rect 8000 14590 8034 14614
rect 8000 14580 8002 14590
rect 8002 14580 8034 14590
rect 8000 14522 8034 14542
rect 8000 14508 8002 14522
rect 8002 14508 8034 14522
rect 8000 14454 8034 14470
rect 8000 14436 8002 14454
rect 8002 14436 8034 14454
rect 8000 14386 8034 14398
rect 8000 14364 8002 14386
rect 8002 14364 8034 14386
rect 8000 14318 8034 14326
rect 8000 14292 8002 14318
rect 8002 14292 8034 14318
rect 8000 14250 8034 14254
rect 8000 14220 8002 14250
rect 8002 14220 8034 14250
rect 8000 14148 8002 14182
rect 8002 14148 8034 14182
rect 8000 14080 8002 14110
rect 8002 14080 8034 14110
rect 8000 14076 8034 14080
rect 8000 14012 8002 14038
rect 8002 14012 8034 14038
rect 8000 14004 8034 14012
rect 8000 13944 8002 13966
rect 8002 13944 8034 13966
rect 8000 13932 8034 13944
rect 8000 13876 8002 13894
rect 8002 13876 8034 13894
rect 8000 13860 8034 13876
rect 8000 13808 8002 13822
rect 8002 13808 8034 13822
rect 8000 13788 8034 13808
rect 8000 13740 8002 13750
rect 8002 13740 8034 13750
rect 8000 13716 8034 13740
rect 8000 13672 8002 13678
rect 8002 13672 8034 13678
rect 8000 13644 8034 13672
rect 8000 13604 8002 13606
rect 8002 13604 8034 13606
rect 8000 13572 8034 13604
rect 8000 13502 8034 13534
rect 8000 13500 8002 13502
rect 8002 13500 8034 13502
rect 8000 13434 8034 13462
rect 8000 13428 8002 13434
rect 8002 13428 8034 13434
rect 8000 13366 8034 13390
rect 8000 13356 8002 13366
rect 8002 13356 8034 13366
rect 8000 13298 8034 13318
rect 8000 13284 8002 13298
rect 8002 13284 8034 13298
rect 8000 13230 8034 13246
rect 8000 13212 8002 13230
rect 8002 13212 8034 13230
rect 8000 13162 8034 13174
rect 8000 13140 8002 13162
rect 8002 13140 8034 13162
rect 8000 13094 8034 13102
rect 8000 13068 8002 13094
rect 8002 13068 8034 13094
rect 8000 13026 8034 13030
rect 8000 12996 8002 13026
rect 8002 12996 8034 13026
rect 8000 12924 8002 12958
rect 8002 12924 8034 12958
rect 8000 12856 8002 12886
rect 8002 12856 8034 12886
rect 8000 12852 8034 12856
rect 8000 12788 8002 12814
rect 8002 12788 8034 12814
rect 8000 12780 8034 12788
rect 8000 12720 8002 12742
rect 8002 12720 8034 12742
rect 8000 12708 8034 12720
rect 8000 12652 8002 12670
rect 8002 12652 8034 12670
rect 8000 12636 8034 12652
rect 8000 12584 8002 12598
rect 8002 12584 8034 12598
rect 8000 12564 8034 12584
rect 8000 12516 8002 12526
rect 8002 12516 8034 12526
rect 8000 12492 8034 12516
rect 8000 12448 8002 12454
rect 8002 12448 8034 12454
rect 8000 12420 8034 12448
rect 8000 12380 8002 12382
rect 8002 12380 8034 12382
rect 8000 12348 8034 12380
rect 8000 12278 8034 12310
rect 8000 12276 8002 12278
rect 8002 12276 8034 12278
rect 8000 12210 8034 12238
rect 8000 12204 8002 12210
rect 8002 12204 8034 12210
rect 8000 12142 8034 12166
rect 8000 12132 8002 12142
rect 8002 12132 8034 12142
rect 8000 12074 8034 12094
rect 8000 12060 8002 12074
rect 8002 12060 8034 12074
rect 8000 12006 8034 12022
rect 8000 11988 8002 12006
rect 8002 11988 8034 12006
rect 8000 11938 8034 11950
rect 8000 11916 8002 11938
rect 8002 11916 8034 11938
rect 8000 11870 8034 11878
rect 8000 11844 8002 11870
rect 8002 11844 8034 11870
rect 8000 11802 8034 11806
rect 8000 11772 8002 11802
rect 8002 11772 8034 11802
rect 8000 11700 8002 11734
rect 8002 11700 8034 11734
rect 8000 11632 8002 11662
rect 8002 11632 8034 11662
rect 8000 11628 8034 11632
rect 8000 11564 8002 11590
rect 8002 11564 8034 11590
rect 8000 11556 8034 11564
rect 8000 11496 8002 11518
rect 8002 11496 8034 11518
rect 8000 11484 8034 11496
rect 8000 11428 8002 11446
rect 8002 11428 8034 11446
rect 8000 11412 8034 11428
rect 2879 11365 2913 11399
rect 2956 11365 2960 11399
rect 2960 11365 2990 11399
rect 3033 11365 3062 11399
rect 3062 11365 3067 11399
rect 3110 11365 3130 11399
rect 3130 11365 3144 11399
rect 3188 11365 3198 11399
rect 3198 11365 3222 11399
rect 3266 11365 3300 11399
rect 3344 11365 3368 11399
rect 3368 11365 3378 11399
rect 3422 11365 3436 11399
rect 3436 11365 3456 11399
rect 3500 11365 3504 11399
rect 3504 11365 3534 11399
rect 3578 11365 3606 11399
rect 3606 11365 3612 11399
rect 3656 11365 3674 11399
rect 3674 11365 3690 11399
rect 3766 11365 3776 11399
rect 3776 11365 3800 11399
rect 3839 11365 3844 11399
rect 3844 11365 3873 11399
rect 3912 11365 3946 11399
rect 3985 11365 4014 11399
rect 4014 11365 4019 11399
rect 4058 11365 4082 11399
rect 4082 11365 4092 11399
rect 4131 11365 4150 11399
rect 4150 11365 4165 11399
rect 4204 11365 4218 11399
rect 4218 11365 4238 11399
rect 4277 11365 4286 11399
rect 4286 11365 4311 11399
rect 4350 11365 4354 11399
rect 4354 11365 4384 11399
rect 4423 11365 4456 11399
rect 4456 11365 4457 11399
rect 4496 11365 4524 11399
rect 4524 11365 4530 11399
rect 4569 11365 4592 11399
rect 4592 11365 4603 11399
rect 4642 11365 4660 11399
rect 4660 11365 4676 11399
rect 4715 11365 4728 11399
rect 4728 11365 4749 11399
rect 4788 11365 4796 11399
rect 4796 11365 4822 11399
rect 4861 11365 4864 11399
rect 4864 11365 4895 11399
rect 4934 11365 4966 11399
rect 4966 11365 4968 11399
rect 5007 11365 5034 11399
rect 5034 11365 5041 11399
rect 5080 11365 5102 11399
rect 5102 11365 5114 11399
rect 5153 11365 5170 11399
rect 5170 11365 5187 11399
rect 5226 11365 5238 11399
rect 5238 11365 5260 11399
rect 5299 11365 5306 11399
rect 5306 11365 5333 11399
rect 5372 11365 5374 11399
rect 5374 11365 5406 11399
rect 5445 11365 5476 11399
rect 5476 11365 5479 11399
rect 5518 11365 5544 11399
rect 5544 11365 5552 11399
rect 5591 11365 5612 11399
rect 5612 11365 5625 11399
rect 5664 11365 5680 11399
rect 5680 11365 5698 11399
rect 5737 11365 5748 11399
rect 5748 11365 5771 11399
rect 5811 11365 5816 11399
rect 5816 11365 5845 11399
rect 5885 11365 5918 11399
rect 5918 11365 5919 11399
rect 5959 11365 5986 11399
rect 5986 11365 5993 11399
rect 6033 11365 6054 11399
rect 6054 11365 6067 11399
rect 6107 11365 6122 11399
rect 6122 11365 6141 11399
rect 6181 11365 6190 11399
rect 6190 11365 6215 11399
rect 6255 11365 6258 11399
rect 6258 11365 6289 11399
rect 6329 11365 6360 11399
rect 6360 11365 6363 11399
rect 6403 11365 6428 11399
rect 6428 11365 6437 11399
rect 6477 11365 6511 11399
rect 6551 11365 6553 11399
rect 6553 11365 6585 11399
rect 6625 11365 6655 11399
rect 6655 11365 6659 11399
rect 6699 11365 6723 11399
rect 6723 11365 6733 11399
rect 6773 11365 6791 11399
rect 6791 11365 6807 11399
rect 6847 11365 6859 11399
rect 6859 11365 6881 11399
rect 6921 11365 6927 11399
rect 6927 11365 6955 11399
rect 6995 11365 7029 11399
rect 7069 11365 7097 11399
rect 7097 11365 7103 11399
rect 7143 11365 7165 11399
rect 7165 11365 7177 11399
rect 7217 11365 7233 11399
rect 7233 11365 7251 11399
rect 7291 11365 7301 11399
rect 7301 11365 7325 11399
rect 7365 11365 7369 11399
rect 7369 11365 7399 11399
rect 2802 11297 2836 11327
rect 2802 11293 2836 11297
rect 2802 11229 2836 11254
rect 2802 11220 2836 11229
rect 2802 11161 2836 11181
rect 2802 11147 2836 11161
rect 2802 11093 2836 11108
rect 2802 11074 2836 11093
rect 2802 11025 2836 11035
rect 2802 11001 2836 11025
rect 2802 10957 2836 10962
rect 2802 10928 2836 10957
rect 2802 10855 2836 10889
rect 2802 10787 2836 10816
rect 2802 10782 2836 10787
rect 2802 10719 2836 10743
rect 2802 10709 2836 10719
rect 2802 10651 2836 10670
rect 2802 10636 2836 10651
rect 2802 10583 2836 10597
rect 2802 10563 2836 10583
rect 2802 10515 2836 10524
rect 2802 10490 2836 10515
rect 2802 10447 2836 10451
rect 2802 10417 2836 10447
rect 2802 10345 2836 10378
rect 2802 10344 2836 10345
rect 2802 10277 2836 10305
rect 2802 10271 2836 10277
rect 2802 10209 2836 10232
rect 2802 10198 2836 10209
rect 2802 10141 2836 10159
rect 2802 10125 2836 10141
rect 2802 10073 2836 10086
rect 2802 10052 2836 10073
rect 2802 10005 2836 10013
rect 2802 9979 2836 10005
rect 2802 9937 2836 9940
rect 2802 9906 2836 9937
rect 2802 9835 2836 9867
rect 2802 9833 2836 9835
rect 2802 9767 2836 9794
rect 2802 9760 2836 9767
rect 2802 9699 2836 9721
rect 2802 9687 2836 9699
rect 2802 9631 2836 9648
rect 2802 9614 2836 9631
rect 2802 9563 2836 9575
rect 2802 9541 2836 9563
rect 2802 9495 2836 9502
rect 2802 9468 2836 9495
rect 2802 9427 2836 9429
rect 2802 9395 2836 9427
rect 2802 9325 2836 9356
rect 2802 9322 2836 9325
rect 2802 9257 2836 9283
rect 2802 9249 2836 9257
rect 2802 9189 2836 9210
rect 2802 9176 2836 9189
rect 2802 9121 2836 9137
rect 2802 9103 2836 9121
rect 2802 9053 2836 9064
rect 2802 9030 2836 9053
rect 2802 8985 2836 8991
rect 2802 8957 2836 8985
rect 2802 8917 2836 8918
rect 2802 8884 2836 8917
rect 2802 8815 2836 8845
rect 2802 8811 2836 8815
rect 2802 8747 2836 8772
rect 2802 8738 2836 8747
rect 2802 8679 2836 8699
rect 2802 8665 2836 8679
rect 2802 8611 2836 8626
rect 2802 8592 2836 8611
rect 2802 8543 2836 8553
rect 2802 8519 2836 8543
rect 2802 8475 2836 8480
rect 2802 8446 2836 8475
rect 2802 8373 2836 8407
rect 2802 8305 2836 8334
rect 2802 8300 2836 8305
rect 2802 8237 2836 8261
rect 2802 8227 2836 8237
rect 2802 8169 2836 8188
rect 2802 8154 2836 8169
rect 2802 8101 2836 8115
rect 2802 8081 2836 8101
rect 7437 11318 7471 11325
rect 7437 11291 7471 11318
rect 7437 11250 7471 11251
rect 7437 11217 7471 11250
rect 7437 11148 7471 11177
rect 7437 11143 7471 11148
rect 7437 11080 7471 11103
rect 7437 11069 7471 11080
rect 7437 11012 7471 11029
rect 7437 10995 7471 11012
rect 7437 10944 7471 10955
rect 7437 10921 7471 10944
rect 7437 10876 7471 10880
rect 7437 10846 7471 10876
rect 7437 10774 7471 10805
rect 7437 10771 7471 10774
rect 7437 10706 7471 10730
rect 7437 10696 7471 10706
rect 7437 10638 7471 10655
rect 7437 10621 7471 10638
rect 7437 10570 7471 10580
rect 7437 10546 7471 10570
rect 7437 10502 7471 10505
rect 7437 10471 7471 10502
rect 7437 10400 7471 10401
rect 7437 10367 7471 10400
rect 7437 10298 7471 10328
rect 7437 10294 7471 10298
rect 7437 10230 7471 10255
rect 7437 10221 7471 10230
rect 7437 10162 7471 10182
rect 7437 10148 7471 10162
rect 7437 10094 7471 10108
rect 7437 10074 7471 10094
rect 7437 10026 7471 10034
rect 7437 10000 7471 10026
rect 7437 9958 7471 9960
rect 7437 9926 7471 9958
rect 7437 9856 7471 9886
rect 7437 9852 7471 9856
rect 7437 9788 7471 9812
rect 7437 9778 7471 9788
rect 7437 9720 7471 9738
rect 7437 9704 7471 9720
rect 7437 9652 7471 9664
rect 7437 9630 7471 9652
rect 7437 9584 7471 9590
rect 7437 9556 7471 9584
rect 7437 9482 7471 9516
rect 7437 9438 7471 9442
rect 7437 9408 7471 9438
rect 7437 9336 7471 9368
rect 7437 9334 7471 9336
rect 7437 9268 7471 9294
rect 7437 9260 7471 9268
rect 7437 9200 7471 9220
rect 7437 9186 7471 9200
rect 7437 9132 7471 9146
rect 7437 9112 7471 9132
rect 7437 9064 7471 9072
rect 7437 9038 7471 9064
rect 7437 8996 7471 8998
rect 7437 8964 7471 8996
rect 7437 8894 7471 8924
rect 7437 8890 7471 8894
rect 7437 8826 7471 8850
rect 7437 8816 7471 8826
rect 7437 8758 7471 8776
rect 7437 8742 7471 8758
rect 7437 8690 7471 8702
rect 7437 8668 7471 8690
rect 7437 8622 7471 8628
rect 7437 8594 7471 8622
rect 7437 8520 7471 8554
rect 7437 8452 7471 8480
rect 7437 8446 7471 8452
rect 7437 8384 7471 8406
rect 7437 8372 7471 8384
rect 7437 8316 7471 8332
rect 7437 8298 7471 8316
rect 7437 8248 7471 8258
rect 7437 8224 7471 8248
rect 7437 8180 7471 8184
rect 7437 8150 7471 8180
rect 2802 8033 2836 8042
rect 2802 8008 2836 8033
rect 2802 7965 2836 7969
rect 2802 7935 2836 7965
rect 6750 8060 6784 8094
rect 7048 8078 7082 8112
rect 7126 8078 7134 8112
rect 7134 8078 7160 8112
rect 7204 8078 7236 8112
rect 7236 8078 7238 8112
rect 7282 8078 7304 8112
rect 7304 8078 7316 8112
rect 7360 8078 7394 8112
rect 8000 11360 8002 11374
rect 8002 11360 8034 11374
rect 8000 11340 8034 11360
rect 8000 11292 8002 11302
rect 8002 11292 8034 11302
rect 8000 11268 8034 11292
rect 8000 11224 8002 11230
rect 8002 11224 8034 11230
rect 8000 11196 8034 11224
rect 8000 11156 8002 11158
rect 8002 11156 8034 11158
rect 8000 11124 8034 11156
rect 8000 11054 8034 11086
rect 8000 11052 8002 11054
rect 8002 11052 8034 11054
rect 8000 10986 8034 11014
rect 8000 10980 8002 10986
rect 8002 10980 8034 10986
rect 8000 10918 8034 10942
rect 8000 10908 8002 10918
rect 8002 10908 8034 10918
rect 8000 10850 8034 10870
rect 8000 10836 8002 10850
rect 8002 10836 8034 10850
rect 8000 10782 8034 10798
rect 8000 10764 8002 10782
rect 8002 10764 8034 10782
rect 8000 10714 8034 10726
rect 8000 10692 8002 10714
rect 8002 10692 8034 10714
rect 8000 10646 8034 10654
rect 8000 10620 8002 10646
rect 8002 10620 8034 10646
rect 8000 10578 8034 10582
rect 8000 10548 8002 10578
rect 8002 10548 8034 10578
rect 8000 10476 8002 10510
rect 8002 10476 8034 10510
rect 8000 10408 8002 10438
rect 8002 10408 8034 10438
rect 8000 10404 8034 10408
rect 8000 10340 8002 10366
rect 8002 10340 8034 10366
rect 8000 10332 8034 10340
rect 8000 10272 8002 10294
rect 8002 10272 8034 10294
rect 8000 10260 8034 10272
rect 8000 10204 8002 10222
rect 8002 10204 8034 10222
rect 8000 10188 8034 10204
rect 8000 10136 8002 10150
rect 8002 10136 8034 10150
rect 8000 10116 8034 10136
rect 8000 10068 8002 10078
rect 8002 10068 8034 10078
rect 8000 10044 8034 10068
rect 8000 10000 8002 10006
rect 8002 10000 8034 10006
rect 8000 9972 8034 10000
rect 8000 9932 8002 9934
rect 8002 9932 8034 9934
rect 8000 9900 8034 9932
rect 8000 9830 8034 9862
rect 8000 9828 8002 9830
rect 8002 9828 8034 9830
rect 8000 9762 8034 9790
rect 8000 9756 8002 9762
rect 8002 9756 8034 9762
rect 8000 9694 8034 9718
rect 8000 9684 8002 9694
rect 8002 9684 8034 9694
rect 8000 9626 8034 9646
rect 8000 9612 8002 9626
rect 8002 9612 8034 9626
rect 8000 9558 8034 9574
rect 8000 9540 8002 9558
rect 8002 9540 8034 9558
rect 8000 9490 8034 9502
rect 8000 9468 8002 9490
rect 8002 9468 8034 9490
rect 8000 9422 8034 9430
rect 8000 9396 8002 9422
rect 8002 9396 8034 9422
rect 8000 9354 8034 9358
rect 8000 9324 8002 9354
rect 8002 9324 8034 9354
rect 8000 9252 8002 9286
rect 8002 9252 8034 9286
rect 8000 9184 8002 9214
rect 8002 9184 8034 9214
rect 8000 9180 8034 9184
rect 8000 9116 8002 9142
rect 8002 9116 8034 9142
rect 8000 9108 8034 9116
rect 8000 9048 8002 9070
rect 8002 9048 8034 9070
rect 8000 9036 8034 9048
rect 8000 8980 8002 8998
rect 8002 8980 8034 8998
rect 8000 8964 8034 8980
rect 8000 8912 8002 8926
rect 8002 8912 8034 8926
rect 8000 8892 8034 8912
rect 8000 8844 8002 8854
rect 8002 8844 8034 8854
rect 8000 8820 8034 8844
rect 8000 8776 8002 8782
rect 8002 8776 8034 8782
rect 8000 8748 8034 8776
rect 8000 8708 8002 8710
rect 8002 8708 8034 8710
rect 8000 8676 8034 8708
rect 8000 8606 8034 8638
rect 8000 8604 8002 8606
rect 8002 8604 8034 8606
rect 8000 8538 8034 8566
rect 8000 8532 8002 8538
rect 8002 8532 8034 8538
rect 8000 8470 8034 8494
rect 8000 8460 8002 8470
rect 8002 8460 8034 8470
rect 8000 8402 8034 8422
rect 8000 8388 8002 8402
rect 8002 8388 8034 8402
rect 8000 8334 8034 8350
rect 8000 8316 8002 8334
rect 8002 8316 8034 8334
rect 8000 8266 8034 8278
rect 8000 8244 8002 8266
rect 8002 8244 8034 8266
rect 8000 8198 8034 8206
rect 8000 8172 8002 8198
rect 8002 8172 8034 8198
rect 8000 8130 8034 8134
rect 8000 8100 8002 8130
rect 8002 8100 8034 8130
rect 6750 7958 6784 7992
rect 2802 7863 2836 7896
rect 2802 7862 2836 7863
rect 2802 7795 2836 7823
rect 2802 7789 2836 7795
rect 2802 7727 2836 7750
rect 2802 7716 2836 7727
rect 6750 7863 6784 7888
rect 6750 7854 6784 7863
rect 6750 7795 6784 7815
rect 6750 7781 6784 7795
rect 2802 7659 2836 7677
rect 2802 7643 2836 7659
rect 2802 7591 2836 7604
rect 2802 7570 2836 7591
rect 2802 7523 2836 7531
rect 2802 7497 2836 7523
rect 2802 7455 2836 7458
rect 2802 7424 2836 7455
rect 2802 7353 2836 7385
rect 2802 7351 2836 7353
rect 2802 7285 2836 7312
rect 2802 7278 2836 7285
rect 2802 7217 2836 7239
rect 2802 7205 2836 7217
rect 2802 7149 2836 7166
rect 2802 7132 2836 7149
rect 2802 7081 2836 7093
rect 2802 7059 2836 7081
rect 2802 7013 2836 7020
rect 2802 6986 2836 7013
rect 2802 6945 2836 6947
rect 2802 6913 2836 6945
rect 2802 6843 2836 6874
rect 2802 6840 2836 6843
rect 2802 6775 2836 6801
rect 2802 6767 2836 6775
rect 2802 6707 2836 6729
rect 2802 6695 2836 6707
rect 2802 6639 2836 6657
rect 2802 6623 2836 6639
rect 2802 6571 2836 6585
rect 2802 6551 2836 6571
rect 2802 6503 2836 6513
rect 2802 6479 2836 6503
rect 2802 6435 2836 6441
rect 2802 6407 2836 6435
rect 2802 6367 2836 6369
rect 2802 6335 2836 6367
rect 2802 6265 2836 6297
rect 2802 6263 2836 6265
rect 2802 6197 2836 6225
rect 2802 6191 2836 6197
rect 2802 6129 2836 6153
rect 2802 6119 2836 6129
rect 2802 6061 2836 6081
rect 2802 6047 2836 6061
rect 2802 5993 2836 6009
rect 2802 5975 2836 5993
rect 2802 5925 2836 5937
rect 2802 5903 2836 5925
rect 2802 5857 2836 5865
rect 2802 5831 2836 5857
rect 2802 5789 2836 5793
rect 2802 5759 2836 5789
rect 2802 5687 2836 5721
rect 2802 5619 2836 5649
rect 2802 5615 2836 5619
rect 2802 5551 2836 5577
rect 2802 5543 2836 5551
rect 2802 5483 2836 5505
rect 2802 5471 2836 5483
rect 2802 5415 2836 5433
rect 2802 5399 2836 5415
rect 2802 5347 2836 5361
rect 2802 5327 2836 5347
rect 2802 5279 2836 5289
rect 2802 5255 2836 5279
rect 3164 7689 3192 7723
rect 3192 7689 3198 7723
rect 3246 7689 3260 7723
rect 3260 7689 3280 7723
rect 3328 7689 3362 7723
rect 3411 7689 3430 7723
rect 3430 7689 3445 7723
rect 3494 7689 3498 7723
rect 3498 7689 3528 7723
rect 3604 7689 3634 7723
rect 3634 7689 3638 7723
rect 3676 7689 3702 7723
rect 3702 7689 3710 7723
rect 3748 7689 3770 7723
rect 3770 7689 3782 7723
rect 3820 7689 3838 7723
rect 3838 7689 3854 7723
rect 3892 7689 3906 7723
rect 3906 7689 3926 7723
rect 3964 7689 3974 7723
rect 3974 7689 3998 7723
rect 4036 7689 4042 7723
rect 4042 7689 4070 7723
rect 4108 7689 4110 7723
rect 4110 7689 4142 7723
rect 4180 7689 4212 7723
rect 4212 7689 4214 7723
rect 4252 7689 4280 7723
rect 4280 7689 4286 7723
rect 4324 7689 4348 7723
rect 4348 7689 4358 7723
rect 4396 7689 4416 7723
rect 4416 7689 4430 7723
rect 4468 7689 4484 7723
rect 4484 7689 4502 7723
rect 4540 7689 4552 7723
rect 4552 7689 4574 7723
rect 4612 7689 4620 7723
rect 4620 7689 4646 7723
rect 4684 7689 4688 7723
rect 4688 7689 4718 7723
rect 4756 7689 4790 7723
rect 4828 7689 4858 7723
rect 4858 7689 4862 7723
rect 4900 7689 4926 7723
rect 4926 7689 4934 7723
rect 4972 7689 4994 7723
rect 4994 7689 5006 7723
rect 5044 7689 5062 7723
rect 5062 7689 5078 7723
rect 5116 7689 5130 7723
rect 5130 7689 5150 7723
rect 5188 7689 5198 7723
rect 5198 7689 5222 7723
rect 5260 7689 5266 7723
rect 5266 7689 5294 7723
rect 5332 7689 5334 7723
rect 5334 7689 5366 7723
rect 5404 7689 5436 7723
rect 5436 7689 5438 7723
rect 5476 7689 5504 7723
rect 5504 7689 5510 7723
rect 5548 7689 5572 7723
rect 5572 7689 5582 7723
rect 5620 7689 5640 7723
rect 5640 7689 5654 7723
rect 5692 7689 5708 7723
rect 5708 7689 5726 7723
rect 5764 7689 5776 7723
rect 5776 7689 5798 7723
rect 5836 7689 5844 7723
rect 5844 7689 5870 7723
rect 5908 7689 5912 7723
rect 5912 7689 5942 7723
rect 5980 7689 6014 7723
rect 6053 7689 6082 7723
rect 6082 7689 6087 7723
rect 6126 7689 6150 7723
rect 6150 7689 6160 7723
rect 6199 7689 6218 7723
rect 6218 7689 6233 7723
rect 6272 7689 6286 7723
rect 6286 7689 6306 7723
rect 6345 7689 6354 7723
rect 6354 7689 6379 7723
rect 6418 7689 6422 7723
rect 6422 7689 6452 7723
rect 3082 7621 3116 7651
rect 3082 7617 3116 7621
rect 3082 7553 3116 7577
rect 3082 7543 3116 7553
rect 3082 7485 3116 7503
rect 3082 7469 3116 7485
rect 3082 7417 3116 7429
rect 3082 7395 3116 7417
rect 3082 7349 3116 7355
rect 3082 7321 3116 7349
rect 3082 7247 3116 7281
rect 5350 7621 5384 7651
rect 5350 7617 5384 7621
rect 5350 7552 5384 7578
rect 5350 7544 5384 7552
rect 5350 7483 5384 7505
rect 5350 7471 5384 7483
rect 5350 7414 5384 7432
rect 5350 7398 5384 7414
rect 5350 7345 5384 7359
rect 5350 7325 5384 7345
rect 3082 7179 3116 7207
rect 3082 7173 3116 7179
rect 3082 7111 3116 7133
rect 3082 7099 3116 7111
rect 3082 7043 3116 7059
rect 3082 7025 3116 7043
rect 3082 6975 3116 6985
rect 3082 6951 3116 6975
rect 3082 6907 3116 6911
rect 3082 6877 3116 6907
rect 3082 6805 3116 6837
rect 3082 6803 3116 6805
rect 3082 6737 3116 6763
rect 3082 6729 3116 6737
rect 3082 6669 3116 6689
rect 3082 6655 3116 6669
rect 3082 6601 3116 6615
rect 3082 6581 3116 6601
rect 3082 6533 3116 6542
rect 3082 6508 3116 6533
rect 3082 6465 3116 6469
rect 3082 6435 3116 6465
rect 3082 6363 3116 6396
rect 3082 6362 3116 6363
rect 3082 6295 3116 6323
rect 3082 6289 3116 6295
rect 3082 6227 3116 6250
rect 3082 6216 3116 6227
rect 3082 6159 3116 6177
rect 3082 6143 3116 6159
rect 3082 6091 3116 6104
rect 3082 6070 3116 6091
rect 3082 6023 3116 6031
rect 3082 5997 3116 6023
rect 3082 5955 3116 5958
rect 3082 5924 3116 5955
rect 3082 5853 3116 5885
rect 3082 5851 3116 5853
rect 3082 5785 3116 5812
rect 3082 5778 3116 5785
rect 3082 5717 3116 5739
rect 3082 5705 3116 5717
rect 3082 5649 3116 5666
rect 3082 5632 3116 5649
rect 3856 7162 3890 7193
rect 3856 7159 3890 7162
rect 3856 7093 3890 7119
rect 3856 7085 3890 7093
rect 3856 7024 3890 7045
rect 3856 7011 3890 7024
rect 3856 6955 3890 6971
rect 3856 6937 3890 6955
rect 3856 6886 3890 6897
rect 3856 6863 3890 6886
rect 3856 6817 3890 6823
rect 3856 6789 3890 6817
rect 3856 6747 3890 6749
rect 3856 6715 3890 6747
rect 3856 6641 3890 6675
rect 3856 6571 3890 6601
rect 3856 6567 3890 6571
rect 3856 6501 3890 6527
rect 3856 6493 3890 6501
rect 3856 6431 3890 6452
rect 3856 6418 3890 6431
rect 3856 6361 3890 6377
rect 3856 6343 3890 6361
rect 3856 6291 3890 6302
rect 3856 6268 3890 6291
rect 3856 6221 3890 6227
rect 3856 6193 3890 6221
rect 3856 6151 3890 6152
rect 3856 6118 3890 6151
rect 3856 6047 3890 6077
rect 3856 6043 3890 6047
rect 3856 5977 3890 6002
rect 3856 5968 3890 5977
rect 3856 5907 3890 5927
rect 3856 5893 3890 5907
rect 3856 5837 3890 5852
rect 3856 5818 3890 5837
rect 3856 5767 3890 5777
rect 3856 5743 3890 5767
rect 4586 7162 4620 7193
rect 4586 7159 4620 7162
rect 4586 7093 4620 7119
rect 4586 7085 4620 7093
rect 4586 7024 4620 7045
rect 4586 7011 4620 7024
rect 4586 6955 4620 6971
rect 4586 6937 4620 6955
rect 4586 6886 4620 6897
rect 4586 6863 4620 6886
rect 4586 6817 4620 6823
rect 4586 6789 4620 6817
rect 4586 6747 4620 6749
rect 4586 6715 4620 6747
rect 4586 6641 4620 6675
rect 4586 6571 4620 6601
rect 4586 6567 4620 6571
rect 4586 6501 4620 6527
rect 4586 6493 4620 6501
rect 4586 6431 4620 6452
rect 4586 6418 4620 6431
rect 4586 6361 4620 6377
rect 4586 6343 4620 6361
rect 4586 6291 4620 6302
rect 4586 6268 4620 6291
rect 4586 6221 4620 6227
rect 4586 6193 4620 6221
rect 4586 6151 4620 6152
rect 4586 6118 4620 6151
rect 4586 6047 4620 6077
rect 4586 6043 4620 6047
rect 4586 5977 4620 6002
rect 4586 5968 4620 5977
rect 4586 5907 4620 5927
rect 4586 5893 4620 5907
rect 4586 5837 4620 5852
rect 4586 5818 4620 5837
rect 4586 5767 4620 5777
rect 4586 5743 4620 5767
rect 5350 7276 5384 7286
rect 5350 7252 5384 7276
rect 5350 7207 5384 7213
rect 5350 7179 5384 7207
rect 5350 7138 5384 7140
rect 5350 7106 5384 7138
rect 6490 7616 6524 7650
rect 6490 7545 6524 7577
rect 6490 7543 6524 7545
rect 6490 7477 6524 7504
rect 6490 7470 6524 7477
rect 6490 7409 6524 7431
rect 6490 7397 6524 7409
rect 6490 7341 6524 7358
rect 6490 7324 6524 7341
rect 6490 7273 6524 7285
rect 6490 7251 6524 7273
rect 6490 7205 6524 7212
rect 6490 7178 6524 7205
rect 5350 7034 5384 7067
rect 5350 7033 5384 7034
rect 5350 6965 5384 6994
rect 5350 6960 5384 6965
rect 5350 6896 5384 6921
rect 5350 6887 5384 6896
rect 5350 6827 5384 6848
rect 5350 6814 5384 6827
rect 5350 6758 5384 6775
rect 5350 6741 5384 6758
rect 6100 7025 6134 7046
rect 6100 7012 6134 7025
rect 6100 6942 6134 6954
rect 6100 6920 6134 6942
rect 6100 6858 6134 6862
rect 6100 6828 6134 6858
rect 6100 6740 6134 6770
rect 6100 6736 6134 6740
rect 6490 7137 6524 7139
rect 6490 7105 6524 7137
rect 6490 7035 6524 7066
rect 6490 7032 6524 7035
rect 6490 6967 6524 6993
rect 6490 6959 6524 6967
rect 6490 6899 6524 6920
rect 6490 6886 6524 6899
rect 6490 6831 6524 6847
rect 6490 6813 6524 6831
rect 6490 6763 6524 6774
rect 6490 6740 6524 6763
rect 5350 6689 5384 6702
rect 5350 6668 5384 6689
rect 5350 6620 5384 6629
rect 5350 6595 5384 6620
rect 5350 6551 5384 6556
rect 5350 6522 5384 6551
rect 6490 6695 6524 6701
rect 6490 6667 6524 6695
rect 6490 6627 6524 6628
rect 6490 6594 6524 6627
rect 5350 6482 5384 6483
rect 5350 6449 5384 6482
rect 5350 6379 5384 6409
rect 5350 6375 5384 6379
rect 5350 6310 5384 6335
rect 5350 6301 5384 6310
rect 5350 6241 5384 6261
rect 5350 6227 5384 6241
rect 5350 6172 5384 6187
rect 5350 6153 5384 6172
rect 5350 6103 5384 6113
rect 5350 6079 5384 6103
rect 5350 6034 5384 6039
rect 5350 6005 5384 6034
rect 5350 5931 5384 5965
rect 5350 5859 5384 5891
rect 5350 5857 5384 5859
rect 5350 5789 5384 5817
rect 5350 5783 5384 5789
rect 6100 6502 6134 6506
rect 6100 6472 6134 6502
rect 6100 6429 6134 6430
rect 6100 6396 6134 6429
rect 6100 6320 6134 6354
rect 6100 6244 6134 6278
rect 6100 6171 6134 6202
rect 6100 6168 6134 6171
rect 6100 6098 6134 6126
rect 6100 6092 6134 6098
rect 6100 6024 6134 6050
rect 6100 6016 6134 6024
rect 6100 5950 6134 5973
rect 6100 5939 6134 5950
rect 6100 5876 6134 5896
rect 6100 5862 6134 5876
rect 6100 5802 6134 5819
rect 6100 5785 6134 5802
rect 6490 6525 6524 6555
rect 6490 6521 6524 6525
rect 6490 6457 6524 6482
rect 6490 6448 6524 6457
rect 6490 6389 6524 6409
rect 6490 6375 6524 6389
rect 6490 6321 6524 6335
rect 6490 6301 6524 6321
rect 6490 6253 6524 6261
rect 6490 6227 6524 6253
rect 6490 6185 6524 6187
rect 6490 6153 6524 6185
rect 6490 6083 6524 6113
rect 6490 6079 6524 6083
rect 6490 6015 6524 6039
rect 6490 6005 6524 6015
rect 6490 5947 6524 5965
rect 6490 5931 6524 5947
rect 6490 5879 6524 5891
rect 6490 5857 6524 5879
rect 6490 5811 6524 5817
rect 6490 5783 6524 5811
rect 5350 5719 5384 5743
rect 5350 5709 5384 5719
rect 5657 5708 5686 5742
rect 5686 5708 5691 5742
rect 5729 5708 5754 5742
rect 5754 5708 5763 5742
rect 3082 5581 3116 5593
rect 3082 5559 3116 5581
rect 3082 5513 3116 5520
rect 3082 5486 3116 5513
rect 3082 5445 3116 5447
rect 3082 5413 3116 5445
rect 3082 5340 3116 5374
rect 5350 5649 5384 5669
rect 5350 5635 5384 5649
rect 5350 5579 5384 5595
rect 5350 5561 5384 5579
rect 5350 5509 5384 5521
rect 5350 5487 5384 5509
rect 5350 5439 5384 5447
rect 5350 5413 5384 5439
rect 5350 5369 5384 5373
rect 5350 5339 5384 5369
rect 6490 5709 6524 5743
rect 6490 5641 6524 5669
rect 6490 5635 6524 5641
rect 6490 5573 6524 5595
rect 6490 5561 6524 5573
rect 6490 5505 6524 5521
rect 6490 5487 6524 5505
rect 6490 5437 6524 5447
rect 6490 5413 6524 5437
rect 6490 5369 6524 5373
rect 6490 5339 6524 5369
rect 3154 5267 3184 5301
rect 3184 5267 3188 5301
rect 3240 5267 3252 5301
rect 3252 5267 3274 5301
rect 3326 5267 3354 5301
rect 3354 5267 3360 5301
rect 3412 5267 3422 5301
rect 3422 5267 3446 5301
rect 3498 5267 3524 5301
rect 3524 5267 3532 5301
rect 3583 5267 3592 5301
rect 3592 5267 3617 5301
rect 3918 5267 3932 5301
rect 3932 5267 3952 5301
rect 3992 5267 4000 5301
rect 4000 5267 4026 5301
rect 4066 5267 4068 5301
rect 4068 5267 4100 5301
rect 4140 5267 4170 5301
rect 4170 5267 4174 5301
rect 4214 5267 4238 5301
rect 4238 5267 4248 5301
rect 4288 5267 4306 5301
rect 4306 5267 4322 5301
rect 4362 5267 4374 5301
rect 4374 5267 4396 5301
rect 4436 5267 4442 5301
rect 4442 5267 4470 5301
rect 4510 5267 4544 5301
rect 4584 5267 4612 5301
rect 4612 5267 4618 5301
rect 4658 5267 4680 5301
rect 4680 5267 4692 5301
rect 4732 5267 4748 5301
rect 4748 5267 4766 5301
rect 4806 5267 4816 5301
rect 4816 5267 4840 5301
rect 4880 5267 4884 5301
rect 4884 5267 4914 5301
rect 4954 5267 4986 5301
rect 4986 5267 4988 5301
rect 5028 5267 5054 5301
rect 5054 5267 5062 5301
rect 5102 5267 5122 5301
rect 5122 5267 5136 5301
rect 5176 5267 5190 5301
rect 5190 5267 5210 5301
rect 5249 5267 5258 5301
rect 5258 5267 5283 5301
rect 5322 5267 5326 5301
rect 5326 5267 5356 5301
rect 5395 5267 5428 5301
rect 5428 5267 5429 5301
rect 5468 5267 5496 5301
rect 5496 5267 5502 5301
rect 5541 5267 5564 5301
rect 5564 5267 5575 5301
rect 5614 5267 5632 5301
rect 5632 5267 5648 5301
rect 5687 5267 5700 5301
rect 5700 5267 5721 5301
rect 5760 5267 5768 5301
rect 5768 5267 5794 5301
rect 5833 5267 5836 5301
rect 5836 5267 5867 5301
rect 5906 5267 5938 5301
rect 5938 5267 5940 5301
rect 5979 5267 6006 5301
rect 6006 5267 6013 5301
rect 6052 5267 6074 5301
rect 6074 5267 6086 5301
rect 6125 5267 6142 5301
rect 6142 5267 6159 5301
rect 6198 5267 6210 5301
rect 6210 5267 6232 5301
rect 6271 5267 6278 5301
rect 6278 5267 6305 5301
rect 6344 5267 6346 5301
rect 6346 5267 6378 5301
rect 6417 5267 6448 5301
rect 6448 5267 6451 5301
rect 6750 7727 6784 7742
rect 6750 7708 6784 7727
rect 6750 7659 6784 7669
rect 6750 7635 6784 7659
rect 6750 7591 6784 7596
rect 6750 7562 6784 7591
rect 6750 7489 6784 7523
rect 6750 7421 6784 7450
rect 6750 7416 6784 7421
rect 6750 7353 6784 7377
rect 6750 7343 6784 7353
rect 6750 7285 6784 7304
rect 6750 7270 6784 7285
rect 6750 7217 6784 7231
rect 6750 7197 6784 7217
rect 6750 7149 6784 7158
rect 6750 7124 6784 7149
rect 6750 7081 6784 7085
rect 6750 7051 6784 7081
rect 6750 6979 6784 7012
rect 6750 6978 6784 6979
rect 6750 6911 6784 6939
rect 6750 6905 6784 6911
rect 6750 6843 6784 6866
rect 6750 6832 6784 6843
rect 6750 6775 6784 6793
rect 6750 6759 6784 6775
rect 6750 6707 6784 6720
rect 6750 6686 6784 6707
rect 6750 6639 6784 6647
rect 6750 6613 6784 6639
rect 6750 6571 6784 6574
rect 6750 6540 6784 6571
rect 6750 6469 6784 6501
rect 6750 6467 6784 6469
rect 6750 6401 6784 6428
rect 6750 6394 6784 6401
rect 6750 6333 6784 6355
rect 6750 6321 6784 6333
rect 6750 6265 6784 6282
rect 6750 6248 6784 6265
rect 6750 6197 6784 6209
rect 6750 6175 6784 6197
rect 6750 6129 6784 6136
rect 6750 6102 6784 6129
rect 6750 6061 6784 6063
rect 6750 6029 6784 6061
rect 6750 5959 6784 5990
rect 6750 5956 6784 5959
rect 6750 5891 6784 5917
rect 6750 5883 6784 5891
rect 6750 5823 6784 5844
rect 6750 5810 6784 5823
rect 6750 5755 6784 5771
rect 6750 5737 6784 5755
rect 6750 5687 6784 5698
rect 6750 5664 6784 5687
rect 6750 5619 6784 5625
rect 6750 5591 6784 5619
rect 6750 5551 6784 5552
rect 6750 5518 6784 5551
rect 6750 5449 6784 5479
rect 6750 5445 6784 5449
rect 6750 5381 6784 5406
rect 6750 5372 6784 5381
rect 6750 5313 6784 5333
rect 6750 5299 6784 5313
rect 2802 5183 2836 5217
rect 2802 5143 2836 5145
rect 2802 5111 2836 5143
rect 2802 5039 2836 5073
rect 6750 5245 6784 5260
rect 6750 5226 6784 5245
rect 6750 5177 6784 5187
rect 6750 5153 6784 5177
rect 6750 5109 6784 5113
rect 6750 5079 6784 5109
rect 2899 5007 2904 5041
rect 2904 5007 2933 5041
rect 2977 5007 3006 5041
rect 3006 5007 3011 5041
rect 3056 5007 3074 5041
rect 3074 5007 3090 5041
rect 3135 5007 3142 5041
rect 3142 5007 3169 5041
rect 3214 5007 3244 5041
rect 3244 5007 3248 5041
rect 3293 5007 3312 5041
rect 3312 5007 3327 5041
rect 3372 5007 3380 5041
rect 3380 5007 3406 5041
rect 3451 5007 3482 5041
rect 3482 5007 3485 5041
rect 3530 5007 3550 5041
rect 3550 5007 3564 5041
rect 3609 5007 3618 5041
rect 3618 5007 3643 5041
rect 3918 5007 3924 5041
rect 3924 5007 3952 5041
rect 3991 5007 3992 5041
rect 3992 5007 4025 5041
rect 4064 5007 4094 5041
rect 4094 5007 4098 5041
rect 4137 5007 4162 5041
rect 4162 5007 4171 5041
rect 4210 5007 4230 5041
rect 4230 5007 4244 5041
rect 4283 5007 4298 5041
rect 4298 5007 4317 5041
rect 4356 5007 4366 5041
rect 4366 5007 4390 5041
rect 4429 5007 4434 5041
rect 4434 5007 4463 5041
rect 4502 5007 4536 5041
rect 4575 5007 4604 5041
rect 4604 5007 4609 5041
rect 4648 5007 4672 5041
rect 4672 5007 4682 5041
rect 4721 5007 4740 5041
rect 4740 5007 4755 5041
rect 4794 5007 4808 5041
rect 4808 5007 4828 5041
rect 4867 5007 4876 5041
rect 4876 5007 4901 5041
rect 4940 5007 4944 5041
rect 4944 5007 4974 5041
rect 5013 5007 5046 5041
rect 5046 5007 5047 5041
rect 5086 5007 5114 5041
rect 5114 5007 5120 5041
rect 5159 5007 5182 5041
rect 5182 5007 5193 5041
rect 5232 5007 5250 5041
rect 5250 5007 5266 5041
rect 5305 5007 5318 5041
rect 5318 5007 5339 5041
rect 5378 5007 5386 5041
rect 5386 5007 5412 5041
rect 5451 5007 5454 5041
rect 5454 5007 5485 5041
rect 5524 5007 5556 5041
rect 5556 5007 5558 5041
rect 5597 5007 5624 5041
rect 5624 5007 5631 5041
rect 5670 5007 5692 5041
rect 5692 5007 5704 5041
rect 5742 5007 5760 5041
rect 5760 5007 5776 5041
rect 5814 5007 5828 5041
rect 5828 5007 5848 5041
rect 5886 5007 5896 5041
rect 5896 5007 5920 5041
rect 5958 5007 5964 5041
rect 5964 5007 5992 5041
rect 6030 5007 6032 5041
rect 6032 5007 6064 5041
rect 6102 5007 6134 5041
rect 6134 5007 6136 5041
rect 6174 5007 6202 5041
rect 6202 5007 6208 5041
rect 6246 5007 6270 5041
rect 6270 5007 6280 5041
rect 6318 5007 6338 5041
rect 6338 5007 6352 5041
rect 6390 5007 6406 5041
rect 6406 5007 6424 5041
rect 6462 5007 6474 5041
rect 6474 5007 6496 5041
rect 6534 5007 6542 5041
rect 6542 5007 6568 5041
rect 6606 5007 6610 5041
rect 6610 5007 6640 5041
rect 6678 5007 6712 5041
rect 8000 8028 8002 8062
rect 8002 8028 8034 8062
rect 8000 7960 8002 7990
rect 8002 7960 8034 7990
rect 8000 7956 8034 7960
rect 8000 7892 8002 7918
rect 8002 7892 8034 7918
rect 8000 7884 8034 7892
rect 8000 7824 8002 7846
rect 8002 7824 8034 7846
rect 8000 7812 8034 7824
rect 8000 7756 8002 7774
rect 8002 7756 8034 7774
rect 8000 7740 8034 7756
rect 8000 7688 8002 7702
rect 8002 7688 8034 7702
rect 8000 7668 8034 7688
rect 8000 7620 8002 7630
rect 8002 7620 8034 7630
rect 8000 7596 8034 7620
rect 8000 7552 8002 7558
rect 8002 7552 8034 7558
rect 8000 7524 8034 7552
rect 8000 7484 8002 7486
rect 8002 7484 8034 7486
rect 8000 7452 8034 7484
rect 8000 7382 8034 7414
rect 8000 7380 8002 7382
rect 8002 7380 8034 7382
rect 8000 7314 8034 7342
rect 8000 7308 8002 7314
rect 8002 7308 8034 7314
rect 8000 7246 8034 7270
rect 8000 7236 8002 7246
rect 8002 7236 8034 7246
rect 8000 7178 8034 7198
rect 8000 7164 8002 7178
rect 8002 7164 8034 7178
rect 8000 7110 8034 7126
rect 8000 7092 8002 7110
rect 8002 7092 8034 7110
rect 8000 7042 8034 7054
rect 8000 7020 8002 7042
rect 8002 7020 8034 7042
rect 8000 6974 8034 6982
rect 8000 6948 8002 6974
rect 8002 6948 8034 6974
rect 8000 6906 8034 6910
rect 8000 6876 8002 6906
rect 8002 6876 8034 6906
rect 8000 6804 8002 6838
rect 8002 6804 8034 6838
rect 8000 6736 8002 6766
rect 8002 6736 8034 6766
rect 8000 6732 8034 6736
rect 8000 6668 8002 6694
rect 8002 6668 8034 6694
rect 8000 6660 8034 6668
rect 8000 6600 8002 6622
rect 8002 6600 8034 6622
rect 8000 6588 8034 6600
rect 8000 6532 8002 6550
rect 8002 6532 8034 6550
rect 8000 6516 8034 6532
rect 8000 6464 8002 6478
rect 8002 6464 8034 6478
rect 8000 6444 8034 6464
rect 8000 6396 8002 6406
rect 8002 6396 8034 6406
rect 8000 6372 8034 6396
rect 8000 6328 8002 6334
rect 8002 6328 8034 6334
rect 8000 6300 8034 6328
rect 8000 6260 8002 6262
rect 8002 6260 8034 6262
rect 8000 6228 8034 6260
rect 8000 6158 8034 6190
rect 8000 6156 8002 6158
rect 8002 6156 8034 6158
rect 8000 6090 8034 6118
rect 8000 6084 8002 6090
rect 8002 6084 8034 6090
rect 8000 6022 8034 6046
rect 8000 6012 8002 6022
rect 8002 6012 8034 6022
rect 8000 5954 8034 5974
rect 8000 5940 8002 5954
rect 8002 5940 8034 5954
rect 8000 5886 8034 5902
rect 8000 5868 8002 5886
rect 8002 5868 8034 5886
rect 8000 5818 8034 5830
rect 8000 5796 8002 5818
rect 8002 5796 8034 5818
rect 8000 5750 8034 5758
rect 8000 5724 8002 5750
rect 8002 5724 8034 5750
rect 8000 5682 8034 5686
rect 8000 5652 8002 5682
rect 8002 5652 8034 5682
rect 8000 5580 8002 5614
rect 8002 5580 8034 5614
rect 8000 5512 8002 5542
rect 8002 5512 8034 5542
rect 8000 5508 8034 5512
rect 8000 5444 8002 5470
rect 8002 5444 8034 5470
rect 8000 5436 8034 5444
rect 8000 5376 8002 5398
rect 8002 5376 8034 5398
rect 8000 5364 8034 5376
rect 8000 5308 8002 5326
rect 8002 5308 8034 5326
rect 8000 5292 8034 5308
rect 8000 5240 8002 5254
rect 8002 5240 8034 5254
rect 8000 5220 8034 5240
rect 8000 5172 8002 5182
rect 8002 5172 8034 5182
rect 8000 5148 8034 5172
rect 8000 5104 8002 5110
rect 8002 5104 8034 5110
rect 8000 5076 8034 5104
rect 8000 5036 8002 5038
rect 8002 5036 8034 5038
rect 8000 5004 8034 5036
rect 8000 4934 8034 4966
rect 8000 4932 8002 4934
rect 8002 4932 8034 4934
rect 2803 4860 2837 4894
rect 2876 4860 2887 4894
rect 2887 4860 2910 4894
rect 2949 4860 2955 4894
rect 2955 4860 2983 4894
rect 3022 4860 3023 4894
rect 3023 4860 3056 4894
rect 3095 4860 3125 4894
rect 3125 4860 3129 4894
rect 3168 4860 3193 4894
rect 3193 4860 3202 4894
rect 3241 4860 3261 4894
rect 3261 4860 3275 4894
rect 3314 4860 3329 4894
rect 3329 4860 3348 4894
rect 3387 4860 3397 4894
rect 3397 4860 3421 4894
rect 3461 4860 3465 4894
rect 3465 4860 3495 4894
rect 3535 4860 3567 4894
rect 3567 4860 3569 4894
rect 3609 4860 3635 4894
rect 3635 4860 3643 4894
rect 3892 4860 3907 4894
rect 3907 4860 3926 4894
rect 3965 4860 3975 4894
rect 3975 4860 3999 4894
rect 4038 4860 4043 4894
rect 4043 4860 4072 4894
rect 4111 4860 4145 4894
rect 4184 4860 4213 4894
rect 4213 4860 4218 4894
rect 4257 4860 4281 4894
rect 4281 4860 4291 4894
rect 4330 4860 4349 4894
rect 4349 4860 4364 4894
rect 4403 4860 4417 4894
rect 4417 4860 4437 4894
rect 4476 4860 4485 4894
rect 4485 4860 4510 4894
rect 4549 4860 4553 4894
rect 4553 4860 4583 4894
rect 4622 4860 4655 4894
rect 4655 4860 4656 4894
rect 4695 4860 4723 4894
rect 4723 4860 4729 4894
rect 4768 4860 4791 4894
rect 4791 4860 4802 4894
rect 4841 4860 4859 4894
rect 4859 4860 4875 4894
rect 4914 4860 4927 4894
rect 4927 4860 4948 4894
rect 4987 4860 4995 4894
rect 4995 4860 5021 4894
rect 5060 4860 5063 4894
rect 5063 4860 5094 4894
rect 5133 4860 5165 4894
rect 5165 4860 5167 4894
rect 5205 4860 5233 4894
rect 5233 4860 5239 4894
rect 5277 4860 5301 4894
rect 5301 4860 5311 4894
rect 5349 4860 5369 4894
rect 5369 4860 5383 4894
rect 5421 4860 5437 4894
rect 5437 4860 5455 4894
rect 5493 4860 5505 4894
rect 5505 4860 5527 4894
rect 5565 4860 5573 4894
rect 5573 4860 5599 4894
rect 5637 4860 5641 4894
rect 5641 4860 5671 4894
rect 5709 4860 5743 4894
rect 5781 4860 5811 4894
rect 5811 4860 5815 4894
rect 5853 4860 5879 4894
rect 5879 4860 5887 4894
rect 5925 4860 5947 4894
rect 5947 4860 5959 4894
rect 5997 4860 6015 4894
rect 6015 4860 6031 4894
rect 6069 4860 6083 4894
rect 6083 4860 6103 4894
rect 6141 4860 6151 4894
rect 6151 4860 6175 4894
rect 6213 4860 6219 4894
rect 6219 4860 6247 4894
rect 6285 4860 6287 4894
rect 6287 4860 6319 4894
rect 6357 4860 6389 4894
rect 6389 4860 6391 4894
rect 6429 4860 6457 4894
rect 6457 4860 6463 4894
rect 6501 4860 6525 4894
rect 6525 4860 6535 4894
rect 6573 4860 6593 4894
rect 6593 4860 6607 4894
rect 6645 4860 6661 4894
rect 6661 4860 6679 4894
rect 6717 4860 6729 4894
rect 6729 4860 6751 4894
rect 8000 4866 8034 4894
rect 8000 4860 8002 4866
rect 8002 4860 8034 4866
rect 8000 4798 8034 4822
rect 8000 4788 8002 4798
rect 8002 4788 8034 4798
rect 3132 4739 3161 4773
rect 3161 4739 3166 4773
rect 3215 4739 3233 4773
rect 3233 4739 3249 4773
rect 3298 4739 3305 4773
rect 3305 4739 3332 4773
rect 3381 4739 3415 4773
rect 3463 4739 3486 4773
rect 3486 4739 3497 4773
rect 3545 4739 3557 4773
rect 3557 4739 3579 4773
rect 8000 4730 8034 4750
rect 6430 4687 6464 4721
rect 6509 4687 6543 4721
rect 6588 4687 6622 4721
rect 8000 4716 8002 4730
rect 8002 4716 8034 4730
rect 4222 4645 4256 4679
rect 2994 4599 3028 4633
rect 2994 4527 3028 4561
rect 2994 4455 3028 4489
rect 2994 4383 3028 4417
rect 2994 4311 3028 4345
rect 2994 4239 3028 4273
rect 2994 4167 3028 4201
rect 2994 4095 3028 4129
rect 2994 4023 3028 4057
rect 2994 3951 3028 3985
rect 2994 3879 3028 3913
rect 2994 3807 3028 3841
rect 2994 3735 3028 3769
rect 2994 3663 3028 3697
rect 2994 3591 3028 3625
rect 2994 3519 3028 3553
rect 2994 3447 3028 3481
rect 2994 3375 3028 3409
rect 2994 3303 3028 3337
rect 3150 4599 3184 4633
rect 3150 4527 3184 4561
rect 3150 4455 3184 4489
rect 3150 4383 3184 4417
rect 3150 4311 3184 4345
rect 3150 4239 3184 4273
rect 3150 4167 3184 4201
rect 3150 4095 3184 4129
rect 3150 4023 3184 4057
rect 3150 3951 3184 3985
rect 3150 3879 3184 3913
rect 3150 3807 3184 3841
rect 3150 3735 3184 3769
rect 3150 3663 3184 3697
rect 3150 3591 3184 3625
rect 3150 3519 3184 3553
rect 3150 3447 3184 3481
rect 3150 3375 3184 3409
rect 3150 3303 3184 3337
rect 3306 4599 3340 4633
rect 3306 4527 3340 4561
rect 3306 4455 3340 4489
rect 3306 4383 3340 4417
rect 3306 4311 3340 4345
rect 3306 4239 3340 4273
rect 3306 4167 3340 4201
rect 3306 4095 3340 4129
rect 3306 4023 3340 4057
rect 3306 3951 3340 3985
rect 3306 3879 3340 3913
rect 3306 3807 3340 3841
rect 3306 3735 3340 3769
rect 3306 3663 3340 3697
rect 3306 3591 3340 3625
rect 3306 3519 3340 3553
rect 3306 3447 3340 3481
rect 3306 3375 3340 3409
rect 3306 3303 3340 3337
rect 3462 4599 3496 4633
rect 3462 4527 3496 4561
rect 3462 4455 3496 4489
rect 3462 4383 3496 4417
rect 3462 4311 3496 4345
rect 3462 4239 3496 4273
rect 3462 4167 3496 4201
rect 3462 4095 3496 4129
rect 3462 4023 3496 4057
rect 3462 3951 3496 3985
rect 3462 3879 3496 3913
rect 3462 3807 3496 3841
rect 3462 3735 3496 3769
rect 3462 3663 3496 3697
rect 3462 3591 3496 3625
rect 3462 3519 3496 3553
rect 3462 3447 3496 3481
rect 3462 3375 3496 3409
rect 3462 3303 3496 3337
rect 3618 4599 3652 4633
rect 3618 4527 3652 4561
rect 4222 4503 4256 4537
rect 5878 4645 5912 4679
rect 5878 4503 5912 4537
rect 3618 4455 3652 4489
rect 6336 4446 6370 4452
rect 3618 4383 3652 4417
rect 4334 4409 4353 4443
rect 4353 4409 4368 4443
rect 4407 4409 4423 4443
rect 4423 4409 4441 4443
rect 4480 4409 4493 4443
rect 4493 4409 4514 4443
rect 4553 4409 4563 4443
rect 4563 4409 4587 4443
rect 4626 4409 4633 4443
rect 4633 4409 4660 4443
rect 4699 4409 4703 4443
rect 4703 4409 4733 4443
rect 4772 4409 4773 4443
rect 4773 4409 4806 4443
rect 4845 4409 4877 4443
rect 4877 4409 4879 4443
rect 4918 4409 4947 4443
rect 4947 4409 4952 4443
rect 4990 4409 5017 4443
rect 5017 4409 5024 4443
rect 5062 4409 5087 4443
rect 5087 4409 5096 4443
rect 5134 4409 5157 4443
rect 5157 4409 5168 4443
rect 5206 4409 5227 4443
rect 5227 4409 5240 4443
rect 5278 4409 5297 4443
rect 5297 4409 5312 4443
rect 5350 4409 5367 4443
rect 5367 4409 5384 4443
rect 5422 4409 5437 4443
rect 5437 4409 5456 4443
rect 5494 4409 5506 4443
rect 5506 4409 5528 4443
rect 5566 4409 5575 4443
rect 5575 4409 5600 4443
rect 5638 4409 5644 4443
rect 5644 4409 5672 4443
rect 6336 4418 6370 4446
rect 6336 4374 6370 4377
rect 3618 4311 3652 4345
rect 3618 4239 3652 4273
rect 3618 4167 3652 4201
rect 4222 4313 4256 4347
rect 4222 4171 4256 4205
rect 5878 4313 5912 4347
rect 5878 4171 5912 4205
rect 6336 4343 6370 4374
rect 6336 4268 6370 4302
rect 8000 4662 8034 4678
rect 8000 4644 8002 4662
rect 8002 4644 8034 4662
rect 8000 4593 8034 4606
rect 8000 4572 8002 4593
rect 8002 4572 8034 4593
rect 8000 4524 8034 4534
rect 8000 4500 8002 4524
rect 8002 4500 8034 4524
rect 8000 4455 8034 4462
rect 8000 4428 8002 4455
rect 8002 4428 8034 4455
rect 8000 4386 8034 4390
rect 8000 4356 8002 4386
rect 8002 4356 8034 4386
rect 8000 4317 8034 4318
rect 8000 4284 8002 4317
rect 8002 4284 8034 4317
rect 6430 4231 6464 4265
rect 6509 4231 6543 4265
rect 6588 4231 6622 4265
rect 6336 4196 6370 4227
rect 6336 4193 6370 4196
rect 3618 4095 3652 4129
rect 3618 4023 3652 4057
rect 6336 4124 6370 4151
rect 6336 4117 6370 4124
rect 6336 4052 6370 4075
rect 4293 4015 4297 4049
rect 4297 4015 4327 4049
rect 4367 4015 4401 4049
rect 4441 4015 4471 4049
rect 4471 4015 4475 4049
rect 4515 4015 4540 4049
rect 4540 4015 4549 4049
rect 4588 4015 4609 4049
rect 4609 4015 4622 4049
rect 4661 4015 4678 4049
rect 4678 4015 4695 4049
rect 4734 4015 4747 4049
rect 4747 4015 4768 4049
rect 4807 4015 4816 4049
rect 4816 4015 4841 4049
rect 4880 4015 4885 4049
rect 4885 4015 4914 4049
rect 4953 4015 4954 4049
rect 4954 4015 4987 4049
rect 5026 4015 5058 4049
rect 5058 4015 5060 4049
rect 5099 4015 5127 4049
rect 5127 4015 5133 4049
rect 5172 4015 5196 4049
rect 5196 4015 5206 4049
rect 5245 4015 5265 4049
rect 5265 4015 5279 4049
rect 5318 4015 5334 4049
rect 5334 4015 5352 4049
rect 5391 4015 5403 4049
rect 5403 4015 5425 4049
rect 5464 4015 5472 4049
rect 5472 4015 5498 4049
rect 5537 4015 5541 4049
rect 5541 4015 5571 4049
rect 5610 4015 5644 4049
rect 5683 4015 5713 4049
rect 5713 4015 5717 4049
rect 5756 4015 5782 4049
rect 5782 4015 5790 4049
rect 6336 4041 6370 4052
rect 3618 3951 3652 3985
rect 6336 3980 6370 3999
rect 6336 3965 6370 3980
rect 3618 3879 3652 3913
rect 3618 3807 3652 3841
rect 4166 3915 4200 3949
rect 4166 3775 4200 3809
rect 5022 3921 5056 3955
rect 5022 3846 5056 3880
rect 5022 3771 5056 3805
rect 5878 3921 5912 3955
rect 5878 3848 5912 3882
rect 6336 3908 6370 3923
rect 6336 3889 6370 3908
rect 8000 4214 8002 4246
rect 8002 4214 8034 4246
rect 8000 4212 8034 4214
rect 8000 4145 8002 4174
rect 8002 4145 8034 4174
rect 8000 4140 8034 4145
rect 8000 4076 8002 4101
rect 8002 4076 8034 4101
rect 8000 4067 8034 4076
rect 8000 4007 8002 4028
rect 8002 4007 8034 4028
rect 8000 3994 8034 4007
rect 8000 3938 8002 3955
rect 8002 3938 8034 3955
rect 8000 3921 8034 3938
rect 8000 3869 8002 3882
rect 8002 3869 8034 3882
rect 8000 3848 8034 3869
rect 5878 3775 5912 3809
rect 6430 3775 6464 3809
rect 6509 3775 6543 3809
rect 6588 3775 6622 3809
rect 8000 3800 8002 3809
rect 8002 3800 8034 3809
rect 8000 3775 8034 3800
rect 3618 3735 3652 3769
rect 3618 3663 3652 3697
rect 3618 3591 3652 3625
rect 3618 3519 3652 3553
rect 3618 3447 3652 3481
rect 3618 3375 3652 3409
rect 3618 3303 3652 3337
rect 8000 3731 8002 3736
rect 8002 3731 8034 3736
rect 8000 3702 8034 3731
rect 8000 3662 8002 3663
rect 8002 3662 8034 3663
rect 8000 3629 8034 3662
rect 8000 3558 8034 3590
rect 8000 3556 8002 3558
rect 8002 3556 8034 3558
rect 8000 3489 8034 3517
rect 8000 3483 8002 3489
rect 8002 3483 8034 3489
rect 8000 3420 8034 3444
rect 8000 3410 8002 3420
rect 8002 3410 8034 3420
rect 8000 3351 8034 3371
rect 8000 3337 8002 3351
rect 8002 3337 8034 3351
rect 8000 3282 8034 3298
rect 8000 3264 8002 3282
rect 8002 3264 8034 3282
rect 8000 3213 8034 3225
rect 8000 3191 8002 3213
rect 8002 3191 8034 3213
rect 2684 3124 2718 3158
rect 2760 3124 2778 3158
rect 2778 3124 2794 3158
rect 2836 3124 2846 3158
rect 2846 3124 2870 3158
rect 2912 3124 2914 3158
rect 2914 3124 2946 3158
rect 2988 3124 3016 3158
rect 3016 3124 3022 3158
rect 3064 3124 3084 3158
rect 3084 3124 3098 3158
rect 3140 3124 3152 3158
rect 3152 3124 3174 3158
rect 3216 3124 3220 3158
rect 3220 3124 3250 3158
rect 3292 3124 3322 3158
rect 3322 3124 3326 3158
rect 3368 3124 3390 3158
rect 3390 3124 3402 3158
rect 3444 3124 3458 3158
rect 3458 3124 3478 3158
rect 3520 3124 3526 3158
rect 3526 3124 3554 3158
rect 3595 3124 3628 3158
rect 3628 3124 3629 3158
rect 3670 3124 3696 3158
rect 3696 3124 3704 3158
rect 3745 3124 3764 3158
rect 3764 3124 3779 3158
rect 3820 3124 3832 3158
rect 3832 3124 3854 3158
rect 8000 3144 8034 3152
rect 2487 2845 2488 2879
rect 2488 2845 2521 2879
rect 2559 2845 2590 2879
rect 2590 2845 2593 2879
rect 2487 2772 2488 2806
rect 2488 2772 2521 2806
rect 2559 2772 2590 2806
rect 2590 2772 2593 2806
rect 2487 2699 2488 2733
rect 2488 2699 2521 2733
rect 2559 2699 2590 2733
rect 2590 2699 2593 2733
rect 2487 2626 2488 2660
rect 2488 2626 2521 2660
rect 2559 2626 2590 2660
rect 2590 2626 2593 2660
rect 2487 2553 2488 2587
rect 2488 2553 2521 2587
rect 2559 2553 2590 2587
rect 2590 2553 2593 2587
rect 2487 2480 2488 2514
rect 2488 2480 2521 2514
rect 2559 2480 2590 2514
rect 2590 2480 2593 2514
rect 2487 2407 2488 2441
rect 2488 2407 2521 2441
rect 2559 2407 2590 2441
rect 2590 2407 2593 2441
rect 2487 2334 2488 2368
rect 2488 2334 2521 2368
rect 2559 2334 2590 2368
rect 2590 2334 2593 2368
rect 2487 2261 2488 2295
rect 2488 2261 2521 2295
rect 2559 2261 2590 2295
rect 2590 2261 2593 2295
rect 2487 2188 2488 2222
rect 2488 2188 2521 2222
rect 2559 2188 2590 2222
rect 2590 2188 2593 2222
rect 2487 2115 2488 2149
rect 2488 2115 2521 2149
rect 2559 2115 2590 2149
rect 2590 2115 2593 2149
rect 2487 2042 2488 2076
rect 2488 2042 2521 2076
rect 2559 2042 2590 2076
rect 2590 2042 2593 2076
rect 2487 1969 2488 2003
rect 2488 1969 2521 2003
rect 2559 1969 2590 2003
rect 2590 1969 2593 2003
rect 2487 1896 2488 1930
rect 2488 1896 2521 1930
rect 2559 1896 2590 1930
rect 2590 1896 2593 1930
rect 2487 1823 2488 1857
rect 2488 1823 2521 1857
rect 2559 1823 2590 1857
rect 2590 1823 2593 1857
rect 2487 1750 2488 1784
rect 2488 1750 2521 1784
rect 2559 1750 2590 1784
rect 2590 1750 2593 1784
rect 2487 1677 2488 1711
rect 2488 1677 2521 1711
rect 2559 1677 2590 1711
rect 2590 1677 2593 1711
rect 2487 1604 2488 1638
rect 2488 1604 2521 1638
rect 2559 1604 2590 1638
rect 2590 1604 2593 1638
rect 2487 1531 2488 1565
rect 2488 1531 2521 1565
rect 2559 1531 2590 1565
rect 2590 1531 2593 1565
rect 2487 1458 2488 1492
rect 2488 1458 2521 1492
rect 2559 1458 2590 1492
rect 2590 1458 2593 1492
rect 2487 1385 2488 1419
rect 2488 1385 2521 1419
rect 2559 1385 2590 1419
rect 2590 1385 2593 1419
rect 2487 1312 2488 1346
rect 2488 1312 2521 1346
rect 2559 1312 2590 1346
rect 2590 1312 2593 1346
rect 2487 1239 2488 1273
rect 2488 1239 2521 1273
rect 2559 1239 2590 1273
rect 2590 1239 2593 1273
rect 2487 1166 2488 1200
rect 2488 1166 2521 1200
rect 2559 1166 2590 1200
rect 2590 1166 2593 1200
rect 2487 1093 2488 1127
rect 2488 1093 2521 1127
rect 2559 1093 2590 1127
rect 2590 1093 2593 1127
rect 2487 1020 2488 1054
rect 2488 1020 2521 1054
rect 2559 1020 2590 1054
rect 2590 1020 2593 1054
rect 2487 947 2488 981
rect 2488 947 2521 981
rect 2559 947 2590 981
rect 2590 947 2593 981
rect 2487 874 2488 908
rect 2488 874 2521 908
rect 2559 874 2590 908
rect 2590 874 2593 908
rect 2487 801 2488 835
rect 2488 801 2521 835
rect 2559 801 2590 835
rect 2590 801 2593 835
rect 2487 728 2488 762
rect 2488 728 2521 762
rect 2559 728 2590 762
rect 2590 728 2593 762
rect 2487 655 2488 689
rect 2488 655 2521 689
rect 2559 655 2590 689
rect 2590 655 2593 689
rect 2487 582 2488 616
rect 2488 582 2521 616
rect 2559 582 2590 616
rect 2590 582 2593 616
rect 2487 509 2488 543
rect 2488 509 2521 543
rect 2559 509 2590 543
rect 2590 509 2593 543
rect 2487 436 2488 470
rect 2488 436 2521 470
rect 2559 436 2590 470
rect 2590 436 2593 470
rect 8000 3118 8002 3144
rect 8002 3118 8034 3144
rect 8000 3075 8034 3079
rect 8000 3045 8002 3075
rect 8002 3045 8034 3075
rect 8000 2972 8002 3006
rect 8002 2972 8034 3006
rect 8000 2903 8002 2933
rect 8002 2903 8034 2933
rect 8000 2899 8034 2903
rect 8000 2834 8002 2860
rect 8002 2834 8034 2860
rect 8000 2826 8034 2834
rect 8000 2765 8002 2787
rect 8002 2765 8034 2787
rect 8000 2753 8034 2765
rect 8000 2696 8002 2714
rect 8002 2696 8034 2714
rect 8000 2680 8034 2696
rect 8000 2627 8002 2641
rect 8002 2627 8034 2641
rect 8000 2607 8034 2627
rect 8000 2558 8002 2568
rect 8002 2558 8034 2568
rect 8000 2534 8034 2558
rect 8000 2489 8002 2495
rect 8002 2489 8034 2495
rect 8000 2461 8034 2489
rect 8000 2420 8002 2422
rect 8002 2420 8034 2422
rect 8000 2388 8034 2420
rect 8000 2316 8034 2349
rect 8000 2315 8002 2316
rect 8002 2315 8034 2316
rect 8000 2247 8034 2276
rect 8000 2242 8002 2247
rect 8002 2242 8034 2247
rect 8000 2178 8034 2203
rect 8000 2169 8002 2178
rect 8002 2169 8034 2178
rect 8000 2109 8034 2130
rect 8000 2096 8002 2109
rect 8002 2096 8034 2109
rect 8000 2040 8034 2057
rect 8000 2023 8002 2040
rect 8002 2023 8034 2040
rect 8000 1971 8034 1984
rect 8000 1950 8002 1971
rect 8002 1950 8034 1971
rect 8000 1902 8034 1911
rect 8000 1877 8002 1902
rect 8002 1877 8034 1902
rect 8000 1833 8034 1838
rect 8000 1804 8002 1833
rect 8002 1804 8034 1833
rect 8000 1764 8034 1765
rect 8000 1731 8002 1764
rect 8002 1731 8034 1764
rect 8000 1661 8002 1692
rect 8002 1661 8034 1692
rect 8000 1658 8034 1661
rect 8000 1592 8002 1619
rect 8002 1592 8034 1619
rect 8000 1585 8034 1592
rect 8000 1523 8002 1546
rect 8002 1523 8034 1546
rect 8000 1512 8034 1523
rect 8000 1454 8002 1473
rect 8002 1454 8034 1473
rect 8000 1439 8034 1454
rect 8000 1385 8002 1400
rect 8002 1385 8034 1400
rect 8000 1366 8034 1385
rect 8000 1316 8002 1327
rect 8002 1316 8034 1327
rect 8000 1293 8034 1316
rect 8000 1247 8002 1254
rect 8002 1247 8034 1254
rect 8000 1220 8034 1247
rect 8000 1178 8002 1181
rect 8002 1178 8034 1181
rect 8000 1147 8034 1178
rect 8000 1074 8034 1108
rect 8000 1005 8034 1035
rect 8000 1001 8002 1005
rect 8002 1001 8034 1005
rect 8000 936 8034 962
rect 8000 928 8002 936
rect 8002 928 8034 936
rect 8000 867 8034 889
rect 8000 855 8002 867
rect 8002 855 8034 867
rect 8000 798 8034 816
rect 8000 782 8002 798
rect 8002 782 8034 798
rect 8000 729 8034 743
rect 8000 709 8002 729
rect 8002 709 8034 729
rect 8000 660 8034 670
rect 8000 636 8002 660
rect 8002 636 8034 660
rect 8000 591 8034 597
rect 8000 563 8002 591
rect 8002 563 8034 591
rect 8000 522 8034 524
rect 8000 490 8002 522
rect 8002 490 8034 522
rect 8000 419 8002 451
rect 8002 419 8034 451
rect 8000 417 8034 419
rect 9752 39512 9786 39529
rect 9752 39495 9786 39512
rect 10559 39679 10593 39713
rect 10631 39679 10665 39713
rect 10559 39606 10593 39640
rect 10631 39606 10665 39640
rect 10559 39533 10593 39567
rect 10631 39533 10665 39567
rect 9752 39444 9786 39457
rect 9752 39423 9786 39444
rect 9752 39376 9786 39385
rect 9752 39351 9786 39376
rect 9752 39308 9786 39313
rect 9752 39279 9786 39308
rect 9752 39240 9786 39241
rect 9752 39207 9786 39240
rect 9752 39138 9786 39169
rect 9752 39135 9786 39138
rect 9752 39070 9786 39097
rect 9752 39063 9786 39070
rect 9752 39002 9786 39025
rect 9752 38991 9786 39002
rect 9752 38934 9786 38953
rect 9752 38919 9786 38934
rect 9752 38866 9786 38881
rect 9752 38847 9786 38866
rect 9752 38798 9786 38809
rect 9752 38775 9786 38798
rect 9752 38730 9786 38737
rect 9752 38703 9786 38730
rect 9752 38662 9786 38665
rect 9752 38631 9786 38662
rect 9752 38560 9786 38593
rect 9752 38559 9786 38560
rect 9752 38492 9786 38521
rect 9752 38487 9786 38492
rect 9752 38424 9786 38449
rect 9752 38415 9786 38424
rect 9752 38356 9786 38377
rect 9752 38343 9786 38356
rect 9752 38288 9786 38305
rect 9752 38271 9786 38288
rect 9752 38220 9786 38233
rect 9752 38199 9786 38220
rect 9752 38152 9786 38161
rect 9752 38127 9786 38152
rect 9752 38084 9786 38089
rect 9752 38055 9786 38084
rect 9752 38016 9786 38017
rect 9752 37983 9786 38016
rect 9752 37914 9786 37945
rect 9752 37911 9786 37914
rect 9752 37846 9786 37873
rect 9752 37839 9786 37846
rect 9752 37778 9786 37801
rect 9752 37767 9786 37778
rect 9752 37710 9786 37729
rect 9752 37695 9786 37710
rect 9752 37642 9786 37657
rect 9752 37623 9786 37642
rect 9752 37574 9786 37585
rect 9752 37551 9786 37574
rect 9752 37506 9786 37513
rect 9752 37479 9786 37506
rect 9752 37438 9786 37441
rect 9752 37407 9786 37438
rect 9752 37336 9786 37369
rect 9752 37335 9786 37336
rect 9752 37268 9786 37297
rect 9752 37263 9786 37268
rect 9752 37200 9786 37225
rect 9752 37191 9786 37200
rect 9752 37132 9786 37153
rect 9752 37119 9786 37132
rect 9752 37064 9786 37081
rect 9752 37047 9786 37064
rect 9752 36996 9786 37009
rect 9752 36975 9786 36996
rect 9752 36928 9786 36937
rect 9752 36903 9786 36928
rect 9752 36860 9786 36865
rect 9752 36831 9786 36860
rect 9752 36792 9786 36793
rect 9752 36759 9786 36792
rect 9752 36690 9786 36721
rect 9752 36687 9786 36690
rect 9752 36622 9786 36649
rect 9752 36615 9786 36622
rect 9752 36554 9786 36577
rect 9752 36543 9786 36554
rect 9752 36486 9786 36505
rect 9752 36471 9786 36486
rect 9752 36418 9786 36433
rect 9752 36399 9786 36418
rect 9752 36350 9786 36361
rect 9752 36327 9786 36350
rect 9752 36282 9786 36289
rect 9752 36255 9786 36282
rect 9752 36214 9786 36217
rect 9752 36183 9786 36214
rect 9752 36112 9786 36145
rect 9752 36111 9786 36112
rect 9752 36044 9786 36073
rect 9752 36039 9786 36044
rect 9752 35976 9786 36001
rect 9752 35967 9786 35976
rect 9752 35908 9786 35929
rect 9752 35895 9786 35908
rect 9752 35840 9786 35857
rect 9752 35823 9786 35840
rect 9752 35772 9786 35785
rect 9752 35751 9786 35772
rect 9752 35704 9786 35713
rect 9752 35679 9786 35704
rect 9752 35636 9786 35641
rect 9752 35607 9786 35636
rect 9752 35568 9786 35569
rect 9752 35535 9786 35568
rect 9752 35466 9786 35497
rect 9752 35463 9786 35466
rect 9752 35398 9786 35425
rect 9752 35391 9786 35398
rect 9752 35330 9786 35353
rect 9752 35319 9786 35330
rect 9752 35262 9786 35281
rect 9752 35247 9786 35262
rect 9752 35194 9786 35209
rect 9752 35175 9786 35194
rect 9752 35126 9786 35137
rect 9752 35103 9786 35126
rect 9752 35058 9786 35065
rect 9752 35031 9786 35058
rect 9752 34990 9786 34993
rect 9752 34959 9786 34990
rect 9752 34888 9786 34921
rect 9752 34887 9786 34888
rect 9752 34820 9786 34849
rect 9752 34815 9786 34820
rect 9752 34752 9786 34777
rect 9752 34743 9786 34752
rect 9752 34684 9786 34705
rect 9752 34671 9786 34684
rect 9752 34616 9786 34633
rect 9752 34599 9786 34616
rect 9752 34548 9786 34561
rect 9752 34527 9786 34548
rect 9752 34480 9786 34489
rect 9752 34455 9786 34480
rect 9752 34412 9786 34417
rect 9752 34383 9786 34412
rect 9752 34344 9786 34345
rect 9752 34311 9786 34344
rect 9752 34242 9786 34273
rect 9752 34239 9786 34242
rect 9752 34174 9786 34201
rect 9752 34167 9786 34174
rect 9752 34106 9786 34129
rect 9752 34095 9786 34106
rect 9752 34038 9786 34057
rect 9752 34023 9786 34038
rect 9752 33970 9786 33985
rect 9752 33951 9786 33970
rect 9752 33902 9786 33913
rect 9752 33879 9786 33902
rect 9752 33834 9786 33841
rect 9752 33807 9786 33834
rect 9752 33766 9786 33769
rect 9752 33735 9786 33766
rect 9752 33664 9786 33697
rect 9752 33663 9786 33664
rect 9752 33596 9786 33625
rect 9752 33591 9786 33596
rect 9752 33528 9786 33553
rect 9752 33519 9786 33528
rect 9752 33460 9786 33481
rect 9752 33447 9786 33460
rect 9752 33392 9786 33409
rect 9752 33375 9786 33392
rect 9752 33324 9786 33337
rect 9752 33303 9786 33324
rect 9752 33256 9786 33265
rect 9752 33231 9786 33256
rect 9752 33188 9786 33193
rect 9752 33159 9786 33188
rect 9752 33120 9786 33121
rect 9752 33087 9786 33120
rect 9752 33018 9786 33049
rect 9752 33015 9786 33018
rect 9752 32950 9786 32977
rect 9752 32943 9786 32950
rect 9752 32882 9786 32905
rect 9752 32871 9786 32882
rect 9752 32814 9786 32833
rect 9752 32799 9786 32814
rect 9752 32746 9786 32761
rect 9752 32727 9786 32746
rect 9752 32678 9786 32689
rect 9752 32655 9786 32678
rect 9752 32610 9786 32617
rect 9752 32583 9786 32610
rect 9752 32542 9786 32545
rect 9752 32511 9786 32542
rect 9752 32440 9786 32473
rect 9752 32439 9786 32440
rect 9752 32372 9786 32401
rect 9752 32367 9786 32372
rect 9752 32304 9786 32329
rect 9752 32295 9786 32304
rect 9752 32236 9786 32257
rect 9752 32223 9786 32236
rect 9752 32168 9786 32185
rect 9752 32151 9786 32168
rect 9752 32100 9786 32113
rect 9752 32079 9786 32100
rect 9752 32032 9786 32041
rect 9752 32007 9786 32032
rect 9752 31964 9786 31969
rect 9752 31935 9786 31964
rect 9752 31896 9786 31897
rect 9752 31863 9786 31896
rect 9752 31794 9786 31825
rect 9752 31791 9786 31794
rect 9752 31726 9786 31753
rect 9752 31719 9786 31726
rect 9752 31658 9786 31681
rect 9752 31647 9786 31658
rect 9752 31590 9786 31609
rect 9752 31575 9786 31590
rect 9752 31522 9786 31537
rect 9752 31503 9786 31522
rect 9752 31454 9786 31465
rect 9752 31431 9786 31454
rect 9752 31386 9786 31393
rect 9752 31359 9786 31386
rect 9752 31318 9786 31321
rect 9752 31287 9786 31318
rect 9752 31216 9786 31249
rect 9752 31215 9786 31216
rect 9752 31148 9786 31177
rect 9752 31143 9786 31148
rect 9752 31080 9786 31105
rect 9752 31071 9786 31080
rect 9752 31012 9786 31033
rect 9752 30999 9786 31012
rect 9752 30944 9786 30961
rect 9752 30927 9786 30944
rect 9752 30876 9786 30889
rect 9752 30855 9786 30876
rect 9752 30808 9786 30817
rect 9752 30783 9786 30808
rect 9752 30740 9786 30745
rect 9752 30711 9786 30740
rect 9752 30672 9786 30673
rect 9752 30639 9786 30672
rect 9752 30570 9786 30601
rect 9752 30567 9786 30570
rect 9752 30502 9786 30529
rect 9752 30495 9786 30502
rect 9752 30434 9786 30457
rect 9752 30423 9786 30434
rect 9752 30366 9786 30385
rect 9752 30351 9786 30366
rect 9752 30298 9786 30313
rect 9752 30279 9786 30298
rect 9752 30230 9786 30241
rect 9752 30207 9786 30230
rect 9752 30162 9786 30169
rect 9752 30135 9786 30162
rect 9752 30094 9786 30097
rect 9752 30063 9786 30094
rect 9752 29992 9786 30025
rect 9752 29991 9786 29992
rect 9752 29924 9786 29953
rect 9752 29919 9786 29924
rect 9752 29856 9786 29881
rect 9752 29847 9786 29856
rect 9752 29788 9786 29809
rect 9752 29775 9786 29788
rect 9752 29720 9786 29737
rect 9752 29703 9786 29720
rect 9752 29652 9786 29665
rect 9752 29631 9786 29652
rect 9752 29584 9786 29593
rect 9752 29559 9786 29584
rect 9752 29516 9786 29521
rect 9752 29487 9786 29516
rect 9752 29448 9786 29449
rect 9752 29415 9786 29448
rect 9752 29346 9786 29377
rect 9752 29343 9786 29346
rect 9752 29278 9786 29305
rect 9752 29271 9786 29278
rect 9752 29210 9786 29233
rect 9752 29199 9786 29210
rect 9752 29142 9786 29161
rect 9752 29127 9786 29142
rect 9752 29074 9786 29089
rect 9752 29055 9786 29074
rect 9752 29006 9786 29017
rect 9752 28983 9786 29006
rect 9752 28938 9786 28945
rect 9752 28911 9786 28938
rect 9752 28870 9786 28873
rect 9752 28839 9786 28870
rect 9752 28768 9786 28801
rect 9752 28767 9786 28768
rect 9752 28700 9786 28729
rect 9752 28695 9786 28700
rect 9752 28632 9786 28657
rect 9752 28623 9786 28632
rect 9752 28564 9786 28585
rect 9752 28551 9786 28564
rect 9752 28496 9786 28513
rect 9752 28479 9786 28496
rect 9752 28428 9786 28441
rect 9752 28407 9786 28428
rect 9752 28360 9786 28369
rect 9752 28335 9786 28360
rect 9752 28292 9786 28297
rect 9752 28263 9786 28292
rect 9752 28224 9786 28225
rect 9752 28191 9786 28224
rect 9752 28122 9786 28153
rect 9752 28119 9786 28122
rect 9752 28054 9786 28081
rect 9752 28047 9786 28054
rect 9752 27986 9786 28009
rect 9752 27975 9786 27986
rect 9752 27918 9786 27937
rect 9752 27903 9786 27918
rect 9752 27850 9786 27865
rect 9752 27831 9786 27850
rect 9752 27782 9786 27793
rect 9752 27759 9786 27782
rect 9752 27714 9786 27721
rect 9752 27687 9786 27714
rect 9752 27646 9786 27649
rect 9752 27615 9786 27646
rect 9752 27544 9786 27577
rect 9752 27543 9786 27544
rect 9752 27476 9786 27505
rect 9752 27471 9786 27476
rect 9752 27408 9786 27433
rect 9752 27399 9786 27408
rect 9752 27340 9786 27361
rect 9752 27327 9786 27340
rect 9752 27272 9786 27289
rect 9752 27255 9786 27272
rect 9752 27204 9786 27217
rect 9752 27183 9786 27204
rect 9752 27136 9786 27145
rect 9752 27111 9786 27136
rect 9752 27068 9786 27073
rect 9752 27039 9786 27068
rect 9752 27000 9786 27001
rect 9752 26967 9786 27000
rect 9752 26898 9786 26929
rect 9752 26895 9786 26898
rect 9752 26830 9786 26857
rect 9752 26823 9786 26830
rect 9752 26762 9786 26785
rect 9752 26751 9786 26762
rect 9752 26694 9786 26713
rect 9752 26679 9786 26694
rect 9752 26626 9786 26641
rect 9752 26607 9786 26626
rect 9752 26558 9786 26569
rect 9752 26535 9786 26558
rect 9752 26490 9786 26497
rect 9752 26463 9786 26490
rect 9752 26422 9786 26425
rect 9752 26391 9786 26422
rect 9752 26320 9786 26353
rect 9752 26319 9786 26320
rect 9752 26252 9786 26281
rect 9752 26247 9786 26252
rect 9752 26184 9786 26209
rect 9752 26175 9786 26184
rect 9752 26116 9786 26137
rect 9752 26103 9786 26116
rect 9752 26048 9786 26065
rect 9752 26031 9786 26048
rect 9752 25980 9786 25993
rect 9752 25959 9786 25980
rect 9752 25912 9786 25921
rect 9752 25887 9786 25912
rect 9752 25844 9786 25849
rect 9752 25815 9786 25844
rect 9752 25776 9786 25777
rect 9752 25743 9786 25776
rect 9752 25674 9786 25705
rect 9752 25671 9786 25674
rect 9752 25606 9786 25633
rect 9752 25599 9786 25606
rect 9752 25538 9786 25561
rect 9752 25527 9786 25538
rect 9752 25470 9786 25489
rect 9752 25455 9786 25470
rect 9752 25402 9786 25417
rect 9752 25383 9786 25402
rect 9752 25334 9786 25345
rect 9752 25311 9786 25334
rect 9752 25266 9786 25273
rect 9752 25239 9786 25266
rect 9752 25198 9786 25201
rect 9752 25167 9786 25198
rect 9752 25096 9786 25129
rect 9752 25095 9786 25096
rect 9752 25028 9786 25057
rect 9752 25023 9786 25028
rect 9752 24960 9786 24985
rect 9752 24951 9786 24960
rect 9752 24892 9786 24913
rect 9752 24879 9786 24892
rect 9752 24824 9786 24841
rect 9752 24807 9786 24824
rect 9752 24756 9786 24769
rect 9752 24735 9786 24756
rect 9752 24688 9786 24697
rect 9752 24663 9786 24688
rect 9752 24620 9786 24625
rect 9752 24591 9786 24620
rect 9752 24552 9786 24553
rect 9752 24519 9786 24552
rect 9752 24450 9786 24481
rect 9752 24447 9786 24450
rect 9752 24382 9786 24409
rect 9752 24375 9786 24382
rect 9752 24314 9786 24337
rect 9752 24303 9786 24314
rect 9752 24246 9786 24265
rect 9752 24231 9786 24246
rect 9752 24178 9786 24193
rect 9752 24159 9786 24178
rect 9752 24110 9786 24121
rect 9752 24087 9786 24110
rect 9752 24042 9786 24049
rect 9752 24015 9786 24042
rect 9752 23974 9786 23977
rect 9752 23943 9786 23974
rect 9752 23872 9786 23905
rect 9752 23871 9786 23872
rect 9752 23804 9786 23833
rect 9752 23799 9786 23804
rect 9752 23736 9786 23761
rect 9752 23727 9786 23736
rect 9752 23668 9786 23689
rect 9752 23655 9786 23668
rect 9752 23600 9786 23617
rect 9752 23583 9786 23600
rect 9752 23532 9786 23545
rect 9752 23511 9786 23532
rect 9752 23464 9786 23473
rect 9752 23439 9786 23464
rect 9752 23396 9786 23401
rect 9752 23367 9786 23396
rect 9752 23328 9786 23329
rect 9752 23295 9786 23328
rect 9752 23226 9786 23257
rect 9752 23223 9786 23226
rect 9752 23158 9786 23185
rect 9752 23151 9786 23158
rect 9752 23090 9786 23113
rect 9752 23079 9786 23090
rect 9752 23022 9786 23041
rect 9752 23007 9786 23022
rect 9752 22954 9786 22969
rect 9752 22935 9786 22954
rect 9752 22886 9786 22897
rect 9752 22863 9786 22886
rect 9752 22818 9786 22825
rect 9752 22791 9786 22818
rect 9752 22750 9786 22753
rect 9752 22719 9786 22750
rect 9752 22648 9786 22681
rect 9752 22647 9786 22648
rect 9752 22580 9786 22609
rect 9752 22575 9786 22580
rect 9752 22512 9786 22537
rect 9752 22503 9786 22512
rect 9752 22444 9786 22465
rect 9752 22431 9786 22444
rect 9752 22376 9786 22393
rect 9752 22359 9786 22376
rect 9752 22308 9786 22321
rect 9752 22287 9786 22308
rect 9752 22240 9786 22249
rect 9752 22215 9786 22240
rect 9752 22172 9786 22177
rect 9752 22143 9786 22172
rect 9752 22104 9786 22105
rect 9752 22071 9786 22104
rect 9752 22002 9786 22033
rect 9752 21999 9786 22002
rect 9752 21934 9786 21961
rect 9752 21927 9786 21934
rect 9752 21866 9786 21889
rect 9752 21855 9786 21866
rect 9752 21798 9786 21817
rect 9752 21783 9786 21798
rect 9752 21730 9786 21745
rect 9752 21711 9786 21730
rect 9752 21662 9786 21673
rect 9752 21639 9786 21662
rect 9752 21594 9786 21601
rect 9752 21567 9786 21594
rect 9752 21526 9786 21529
rect 9752 21495 9786 21526
rect 9752 21424 9786 21457
rect 9752 21423 9786 21424
rect 9752 21356 9786 21385
rect 9752 21351 9786 21356
rect 9752 21288 9786 21313
rect 9752 21279 9786 21288
rect 9752 21220 9786 21241
rect 9752 21207 9786 21220
rect 9752 21152 9786 21169
rect 9752 21135 9786 21152
rect 9752 21084 9786 21097
rect 9752 21063 9786 21084
rect 9752 21016 9786 21025
rect 9752 20991 9786 21016
rect 9752 20948 9786 20953
rect 9752 20919 9786 20948
rect 9752 20880 9786 20881
rect 9752 20847 9786 20880
rect 9752 20778 9786 20809
rect 9752 20775 9786 20778
rect 9752 20710 9786 20737
rect 9752 20703 9786 20710
rect 9752 20642 9786 20665
rect 9752 20631 9786 20642
rect 9752 20574 9786 20593
rect 9752 20559 9786 20574
rect 9752 20506 9786 20521
rect 9752 20487 9786 20506
rect 9752 20438 9786 20449
rect 9752 20415 9786 20438
rect 9752 20370 9786 20377
rect 9752 20343 9786 20370
rect 9752 20302 9786 20305
rect 9752 20271 9786 20302
rect 9752 20200 9786 20233
rect 9752 20199 9786 20200
rect 9752 20132 9786 20161
rect 9752 20127 9786 20132
rect 9752 20064 9786 20089
rect 9752 20055 9786 20064
rect 9752 19996 9786 20017
rect 9752 19983 9786 19996
rect 9752 19928 9786 19945
rect 9752 19911 9786 19928
rect 9752 19860 9786 19873
rect 9752 19839 9786 19860
rect 9752 19792 9786 19801
rect 9752 19767 9786 19792
rect 9752 19724 9786 19729
rect 9752 19695 9786 19724
rect 9752 19656 9786 19657
rect 9752 19623 9786 19656
rect 9752 19554 9786 19585
rect 9752 19551 9786 19554
rect 9752 19486 9786 19513
rect 9752 19479 9786 19486
rect 9752 19418 9786 19441
rect 9752 19407 9786 19418
rect 9752 19350 9786 19369
rect 9752 19335 9786 19350
rect 9752 19282 9786 19297
rect 9752 19263 9786 19282
rect 9752 19214 9786 19225
rect 9752 19191 9786 19214
rect 9752 19146 9786 19153
rect 9752 19119 9786 19146
rect 9752 19078 9786 19081
rect 9752 19047 9786 19078
rect 9752 18976 9786 19009
rect 9752 18975 9786 18976
rect 9752 18908 9786 18937
rect 9752 18903 9786 18908
rect 9752 18840 9786 18865
rect 9752 18831 9786 18840
rect 9752 18772 9786 18793
rect 9752 18759 9786 18772
rect 9752 18704 9786 18721
rect 9752 18687 9786 18704
rect 9752 18636 9786 18649
rect 9752 18615 9786 18636
rect 9752 18568 9786 18577
rect 9752 18543 9786 18568
rect 9752 18500 9786 18505
rect 9752 18471 9786 18500
rect 9752 18432 9786 18433
rect 9752 18399 9786 18432
rect 9752 18330 9786 18361
rect 9752 18327 9786 18330
rect 9752 18262 9786 18289
rect 9752 18255 9786 18262
rect 9752 18194 9786 18217
rect 9752 18183 9786 18194
rect 9752 18126 9786 18145
rect 9752 18111 9786 18126
rect 9752 18058 9786 18073
rect 9752 18039 9786 18058
rect 9752 17990 9786 18001
rect 9752 17967 9786 17990
rect 9752 17922 9786 17929
rect 9752 17895 9786 17922
rect 9752 17854 9786 17857
rect 9752 17823 9786 17854
rect 9752 17752 9786 17785
rect 9752 17751 9786 17752
rect 9752 17684 9786 17713
rect 9752 17679 9786 17684
rect 9752 17616 9786 17641
rect 9752 17607 9786 17616
rect 9752 17548 9786 17569
rect 9752 17535 9786 17548
rect 9752 17480 9786 17497
rect 9752 17463 9786 17480
rect 9752 17412 9786 17425
rect 9752 17391 9786 17412
rect 9752 17344 9786 17353
rect 9752 17319 9786 17344
rect 9752 17276 9786 17281
rect 9752 17247 9786 17276
rect 9752 17208 9786 17209
rect 9752 17175 9786 17208
rect 9752 17106 9786 17137
rect 9752 17103 9786 17106
rect 9752 17038 9786 17065
rect 9752 17031 9786 17038
rect 9752 16970 9786 16993
rect 9752 16959 9786 16970
rect 9752 16902 9786 16921
rect 9752 16887 9786 16902
rect 9752 16834 9786 16849
rect 9752 16815 9786 16834
rect 9752 16766 9786 16777
rect 9752 16743 9786 16766
rect 9752 16698 9786 16705
rect 9752 16671 9786 16698
rect 9752 16630 9786 16633
rect 9752 16599 9786 16630
rect 9752 16528 9786 16561
rect 9752 16527 9786 16528
rect 9752 16460 9786 16489
rect 9752 16455 9786 16460
rect 9752 16392 9786 16417
rect 9752 16383 9786 16392
rect 9752 16324 9786 16345
rect 9752 16311 9786 16324
rect 9752 16256 9786 16273
rect 9752 16239 9786 16256
rect 9752 16188 9786 16201
rect 9752 16167 9786 16188
rect 9752 16120 9786 16129
rect 9752 16095 9786 16120
rect 9752 16052 9786 16057
rect 9752 16023 9786 16052
rect 9752 15984 9786 15985
rect 9752 15951 9786 15984
rect 9752 15882 9786 15913
rect 9752 15879 9786 15882
rect 9752 15814 9786 15841
rect 9752 15807 9786 15814
rect 9752 15746 9786 15769
rect 9752 15735 9786 15746
rect 9752 15678 9786 15697
rect 9752 15663 9786 15678
rect 9752 15610 9786 15625
rect 9752 15591 9786 15610
rect 9752 15542 9786 15553
rect 9752 15519 9786 15542
rect 9752 15474 9786 15481
rect 9752 15447 9786 15474
rect 9752 15406 9786 15409
rect 9752 15375 9786 15406
rect 9752 15304 9786 15337
rect 9752 15303 9786 15304
rect 9752 15236 9786 15265
rect 9752 15231 9786 15236
rect 9752 15168 9786 15193
rect 9752 15159 9786 15168
rect 9752 15100 9786 15121
rect 9752 15087 9786 15100
rect 9752 15032 9786 15049
rect 9752 15015 9786 15032
rect 9752 14964 9786 14977
rect 9752 14943 9786 14964
rect 9752 14896 9786 14905
rect 9752 14871 9786 14896
rect 9752 14828 9786 14833
rect 9752 14799 9786 14828
rect 9752 14760 9786 14761
rect 9752 14727 9786 14760
rect 9752 14658 9786 14689
rect 9752 14655 9786 14658
rect 9752 14590 9786 14617
rect 9752 14583 9786 14590
rect 9752 14522 9786 14545
rect 9752 14511 9786 14522
rect 9752 14454 9786 14473
rect 9752 14439 9786 14454
rect 9752 14386 9786 14401
rect 9752 14367 9786 14386
rect 9752 14318 9786 14329
rect 9752 14295 9786 14318
rect 9752 14250 9786 14257
rect 9752 14223 9786 14250
rect 9752 14182 9786 14185
rect 9752 14151 9786 14182
rect 9752 14080 9786 14113
rect 9752 14079 9786 14080
rect 9752 14012 9786 14041
rect 9752 14007 9786 14012
rect 9752 13944 9786 13969
rect 9752 13935 9786 13944
rect 9752 13876 9786 13897
rect 9752 13863 9786 13876
rect 9752 13808 9786 13825
rect 9752 13791 9786 13808
rect 9752 13740 9786 13753
rect 9752 13719 9786 13740
rect 9752 13672 9786 13681
rect 9752 13647 9786 13672
rect 9752 13604 9786 13609
rect 9752 13575 9786 13604
rect 9752 13536 9786 13537
rect 9752 13503 9786 13536
rect 9752 13434 9786 13465
rect 9752 13431 9786 13434
rect 9752 13366 9786 13393
rect 9752 13359 9786 13366
rect 9752 13298 9786 13321
rect 9752 13287 9786 13298
rect 9752 13230 9786 13249
rect 9752 13215 9786 13230
rect 9752 13162 9786 13177
rect 9752 13143 9786 13162
rect 9752 13094 9786 13105
rect 9752 13071 9786 13094
rect 9752 13026 9786 13033
rect 9752 12999 9786 13026
rect 9752 12958 9786 12961
rect 9752 12927 9786 12958
rect 9752 12856 9786 12889
rect 9752 12855 9786 12856
rect 9752 12788 9786 12817
rect 9752 12783 9786 12788
rect 9752 12720 9786 12745
rect 9752 12711 9786 12720
rect 9752 12652 9786 12673
rect 9752 12639 9786 12652
rect 9752 12584 9786 12601
rect 9752 12567 9786 12584
rect 9752 12516 9786 12529
rect 9752 12495 9786 12516
rect 9752 12448 9786 12457
rect 9752 12423 9786 12448
rect 9752 12380 9786 12385
rect 9752 12351 9786 12380
rect 9752 12312 9786 12313
rect 9752 12279 9786 12312
rect 9752 12210 9786 12241
rect 9752 12207 9786 12210
rect 9752 12142 9786 12169
rect 9752 12135 9786 12142
rect 9752 12074 9786 12097
rect 9752 12063 9786 12074
rect 9752 12006 9786 12025
rect 9752 11991 9786 12006
rect 9752 11938 9786 11953
rect 9752 11919 9786 11938
rect 9752 11870 9786 11881
rect 9752 11847 9786 11870
rect 9752 11802 9786 11809
rect 9752 11775 9786 11802
rect 9752 11734 9786 11737
rect 9752 11703 9786 11734
rect 9752 11632 9786 11665
rect 9752 11631 9786 11632
rect 9752 11564 9786 11593
rect 9752 11559 9786 11564
rect 9752 11496 9786 11521
rect 9752 11487 9786 11496
rect 9752 11428 9786 11449
rect 9752 11415 9786 11428
rect 9752 11360 9786 11377
rect 9752 11343 9786 11360
rect 9752 11292 9786 11305
rect 9752 11271 9786 11292
rect 9752 11224 9786 11233
rect 9752 11199 9786 11224
rect 9752 11156 9786 11161
rect 9752 11127 9786 11156
rect 9752 11088 9786 11089
rect 9752 11055 9786 11088
rect 9752 10986 9786 11017
rect 9752 10983 9786 10986
rect 9752 10918 9786 10945
rect 9752 10911 9786 10918
rect 9752 10850 9786 10873
rect 9752 10839 9786 10850
rect 9752 10782 9786 10801
rect 9752 10767 9786 10782
rect 9752 10714 9786 10729
rect 9752 10695 9786 10714
rect 9752 10646 9786 10657
rect 9752 10623 9786 10646
rect 9752 10578 9786 10585
rect 9752 10551 9786 10578
rect 9752 10510 9786 10513
rect 9752 10479 9786 10510
rect 9752 10408 9786 10441
rect 9752 10407 9786 10408
rect 9752 10340 9786 10369
rect 9752 10335 9786 10340
rect 9752 10272 9786 10297
rect 9752 10263 9786 10272
rect 9752 10204 9786 10225
rect 9752 10191 9786 10204
rect 9752 10136 9786 10153
rect 9752 10119 9786 10136
rect 9752 10068 9786 10081
rect 9752 10047 9786 10068
rect 9752 10000 9786 10009
rect 9752 9975 9786 10000
rect 9752 9932 9786 9937
rect 9752 9903 9786 9932
rect 9752 9864 9786 9865
rect 9752 9831 9786 9864
rect 9752 9762 9786 9793
rect 9752 9759 9786 9762
rect 9752 9694 9786 9721
rect 9752 9687 9786 9694
rect 9752 9626 9786 9649
rect 9752 9615 9786 9626
rect 9752 9558 9786 9577
rect 9752 9543 9786 9558
rect 9752 9490 9786 9505
rect 9752 9471 9786 9490
rect 9752 9422 9786 9433
rect 9752 9399 9786 9422
rect 9752 9354 9786 9361
rect 9752 9327 9786 9354
rect 9752 9286 9786 9289
rect 9752 9255 9786 9286
rect 9752 9184 9786 9217
rect 9752 9183 9786 9184
rect 9752 9116 9786 9145
rect 9752 9111 9786 9116
rect 9752 9048 9786 9073
rect 9752 9039 9786 9048
rect 9752 8980 9786 9001
rect 9752 8967 9786 8980
rect 9752 8912 9786 8929
rect 9752 8895 9786 8912
rect 9752 8844 9786 8857
rect 9752 8823 9786 8844
rect 9752 8776 9786 8785
rect 9752 8751 9786 8776
rect 9752 8708 9786 8713
rect 9752 8679 9786 8708
rect 9752 8640 9786 8641
rect 9752 8607 9786 8640
rect 9752 8538 9786 8569
rect 9752 8535 9786 8538
rect 9752 8470 9786 8497
rect 9752 8463 9786 8470
rect 9752 8402 9786 8425
rect 9752 8391 9786 8402
rect 9752 8334 9786 8353
rect 9752 8319 9786 8334
rect 9752 8266 9786 8281
rect 9752 8247 9786 8266
rect 9752 8198 9786 8209
rect 9752 8175 9786 8198
rect 9752 8130 9786 8137
rect 9752 8103 9786 8130
rect 9752 8062 9786 8065
rect 9752 8031 9786 8062
rect 9752 7960 9786 7993
rect 9752 7959 9786 7960
rect 9752 7892 9786 7921
rect 9752 7887 9786 7892
rect 9752 7824 9786 7849
rect 9752 7815 9786 7824
rect 9752 7756 9786 7777
rect 9752 7743 9786 7756
rect 9752 7688 9786 7705
rect 9752 7671 9786 7688
rect 9752 7620 9786 7633
rect 9752 7599 9786 7620
rect 9752 7552 9786 7561
rect 9752 7527 9786 7552
rect 9752 7484 9786 7489
rect 9752 7455 9786 7484
rect 9752 7416 9786 7417
rect 9752 7383 9786 7416
rect 9752 7314 9786 7345
rect 9752 7311 9786 7314
rect 9752 7246 9786 7273
rect 9752 7239 9786 7246
rect 9752 7178 9786 7201
rect 9752 7167 9786 7178
rect 9752 7110 9786 7129
rect 9752 7095 9786 7110
rect 9752 7042 9786 7057
rect 9752 7023 9786 7042
rect 9752 6974 9786 6985
rect 9752 6951 9786 6974
rect 9752 6906 9786 6913
rect 9752 6879 9786 6906
rect 9752 6838 9786 6841
rect 9752 6807 9786 6838
rect 9752 6736 9786 6769
rect 9752 6735 9786 6736
rect 9752 6668 9786 6697
rect 9752 6663 9786 6668
rect 9752 6600 9786 6625
rect 9752 6591 9786 6600
rect 9752 6532 9786 6553
rect 9752 6519 9786 6532
rect 9752 6464 9786 6481
rect 9752 6447 9786 6464
rect 9752 6396 9786 6409
rect 9752 6375 9786 6396
rect 9752 6328 9786 6337
rect 9752 6303 9786 6328
rect 9752 6260 9786 6265
rect 9752 6231 9786 6260
rect 9752 6192 9786 6193
rect 9752 6159 9786 6192
rect 9752 6090 9786 6121
rect 9752 6087 9786 6090
rect 9752 6022 9786 6049
rect 9752 6015 9786 6022
rect 9752 5954 9786 5977
rect 9752 5943 9786 5954
rect 9752 5886 9786 5905
rect 9752 5871 9786 5886
rect 9752 5818 9786 5833
rect 9752 5799 9786 5818
rect 9752 5750 9786 5761
rect 9752 5727 9786 5750
rect 9752 5682 9786 5689
rect 9752 5655 9786 5682
rect 9752 5614 9786 5617
rect 9752 5583 9786 5614
rect 9752 5512 9786 5545
rect 9752 5511 9786 5512
rect 9752 5444 9786 5473
rect 9752 5439 9786 5444
rect 9752 5376 9786 5401
rect 9752 5367 9786 5376
rect 9752 5308 9786 5329
rect 9752 5295 9786 5308
rect 9752 5240 9786 5257
rect 9752 5223 9786 5240
rect 9752 5172 9786 5185
rect 9752 5151 9786 5172
rect 9752 5104 9786 5113
rect 9752 5079 9786 5104
rect 9752 5036 9786 5041
rect 9752 5007 9786 5036
rect 9752 4968 9786 4969
rect 9752 4935 9786 4968
rect 9752 4866 9786 4897
rect 9752 4863 9786 4866
rect 9752 4798 9786 4825
rect 9752 4791 9786 4798
rect 9752 4730 9786 4753
rect 9752 4719 9786 4730
rect 9752 4662 9786 4681
rect 9752 4647 9786 4662
rect 9752 4594 9786 4609
rect 9752 4575 9786 4594
rect 9752 4526 9786 4537
rect 9752 4503 9786 4526
rect 9752 4458 9786 4465
rect 9752 4431 9786 4458
rect 9752 4390 9786 4393
rect 9752 4359 9786 4390
rect 9752 4288 9786 4321
rect 9752 4287 9786 4288
rect 9752 4220 9786 4249
rect 9752 4215 9786 4220
rect 9752 4152 9786 4177
rect 9752 4143 9786 4152
rect 9752 4084 9786 4105
rect 9752 4071 9786 4084
rect 9752 4016 9786 4033
rect 9752 3999 9786 4016
rect 9752 3948 9786 3961
rect 9752 3927 9786 3948
rect 9752 3880 9786 3889
rect 9752 3855 9786 3880
rect 9752 3812 9786 3817
rect 9752 3783 9786 3812
rect 9752 3744 9786 3745
rect 9752 3711 9786 3744
rect 9752 3642 9786 3673
rect 9752 3639 9786 3642
rect 9752 3574 9786 3601
rect 9752 3567 9786 3574
rect 9752 3506 9786 3529
rect 9752 3495 9786 3506
rect 9752 3438 9786 3457
rect 9752 3423 9786 3438
rect 9752 3370 9786 3385
rect 9752 3351 9786 3370
rect 9752 3302 9786 3313
rect 9752 3279 9786 3302
rect 9752 3234 9786 3241
rect 9752 3207 9786 3234
rect 9752 3166 9786 3168
rect 9752 3134 9786 3166
rect 9752 3064 9786 3095
rect 9752 3061 9786 3064
rect 9752 2996 9786 3022
rect 9752 2988 9786 2996
rect 9752 2928 9786 2949
rect 9752 2915 9786 2928
rect 9752 2860 9786 2876
rect 9752 2842 9786 2860
rect 9752 2792 9786 2803
rect 9752 2769 9786 2792
rect 9752 2724 9786 2730
rect 9752 2696 9786 2724
rect 9752 2656 9786 2657
rect 9752 2623 9786 2656
rect 9752 2554 9786 2584
rect 9752 2550 9786 2554
rect 9752 2486 9786 2511
rect 9752 2477 9786 2486
rect 9752 2418 9786 2438
rect 9752 2404 9786 2418
rect 9752 2349 9786 2365
rect 9752 2331 9786 2349
rect 9752 2280 9786 2292
rect 9752 2258 9786 2280
rect 9752 2211 9786 2219
rect 9752 2185 9786 2211
rect 9752 2142 9786 2146
rect 9752 2112 9786 2142
rect 9752 2039 9786 2073
rect 9752 1970 9786 2000
rect 9752 1966 9786 1970
rect 9752 1901 9786 1927
rect 9752 1893 9786 1901
rect 9752 1832 9786 1854
rect 9752 1820 9786 1832
rect 9752 1763 9786 1781
rect 9752 1747 9786 1763
rect 9752 1694 9786 1708
rect 9752 1674 9786 1694
rect 9752 1625 9786 1635
rect 9752 1601 9786 1625
rect 9752 1556 9786 1562
rect 9752 1528 9786 1556
rect 9752 1487 9786 1489
rect 9752 1455 9786 1487
rect 9752 1383 9786 1416
rect 9752 1382 9786 1383
rect 10716 39752 10786 39784
rect 10786 39752 10820 39786
rect 10820 39752 10822 39786
rect 10716 39718 10822 39752
rect 10716 2487 10718 39718
rect 10718 2487 10820 39718
rect 10820 2487 10822 39718
rect 10716 2414 10718 2448
rect 10718 2414 10750 2448
rect 10788 2414 10820 2448
rect 10820 2414 10822 2448
rect 10716 2341 10718 2375
rect 10718 2341 10750 2375
rect 10788 2341 10820 2375
rect 10820 2341 10822 2375
rect 10716 2268 10718 2302
rect 10718 2268 10750 2302
rect 10788 2268 10820 2302
rect 10820 2268 10822 2302
rect 10716 2195 10718 2229
rect 10718 2195 10750 2229
rect 10788 2195 10820 2229
rect 10820 2195 10822 2229
rect 10716 2122 10718 2156
rect 10718 2122 10750 2156
rect 10788 2122 10820 2156
rect 10820 2122 10822 2156
rect 10716 2049 10718 2083
rect 10718 2049 10750 2083
rect 10788 2049 10820 2083
rect 10820 2049 10822 2083
rect 10716 1976 10718 2010
rect 10718 1976 10750 2010
rect 10788 1976 10820 2010
rect 10820 1976 10822 2010
rect 10716 1903 10718 1937
rect 10718 1903 10750 1937
rect 10788 1903 10820 1937
rect 10820 1903 10822 1937
rect 10716 1830 10718 1864
rect 10718 1830 10750 1864
rect 10788 1830 10820 1864
rect 10820 1830 10822 1864
rect 10716 1757 10718 1791
rect 10718 1757 10750 1791
rect 10788 1757 10820 1791
rect 10820 1757 10822 1791
rect 10716 1684 10718 1718
rect 10718 1684 10750 1718
rect 10788 1684 10820 1718
rect 10820 1684 10822 1718
rect 10716 1611 10718 1645
rect 10718 1611 10750 1645
rect 10788 1611 10820 1645
rect 10820 1611 10822 1645
rect 10716 1538 10718 1572
rect 10718 1538 10750 1572
rect 10788 1538 10820 1572
rect 10820 1538 10822 1572
rect 10716 1465 10718 1499
rect 10718 1465 10750 1499
rect 10788 1465 10820 1499
rect 10820 1465 10822 1499
rect 9752 1314 9786 1343
rect 9752 1309 9786 1314
rect 10137 1293 10243 1399
rect 10716 1392 10718 1426
rect 10718 1392 10750 1426
rect 10788 1392 10820 1426
rect 10820 1392 10822 1426
rect 10716 1319 10718 1353
rect 10718 1319 10750 1353
rect 10788 1319 10820 1353
rect 10820 1319 10822 1353
rect 9752 1245 9786 1270
rect 9752 1236 9786 1245
rect 9752 1176 9786 1197
rect 9752 1163 9786 1176
rect 9752 1107 9786 1124
rect 9752 1090 9786 1107
rect 9752 1038 9786 1051
rect 9752 1017 9786 1038
rect 9752 969 9786 978
rect 9752 944 9786 969
rect 9752 900 9786 905
rect 9752 871 9786 900
rect 9752 831 9786 832
rect 9752 798 9786 831
rect 9752 728 9786 759
rect 9752 725 9786 728
rect 9752 659 9786 686
rect 9752 652 9786 659
rect 9752 590 9786 613
rect 9752 579 9786 590
rect 9752 521 9786 540
rect 9752 506 9786 521
rect 9752 452 9786 467
rect 9752 433 9786 452
rect 8000 350 8002 378
rect 8002 350 8034 378
rect 8000 344 8034 350
rect 8000 281 8002 305
rect 8002 281 8034 305
rect 8000 271 8034 281
rect 8000 212 8002 232
rect 8002 212 8034 232
rect 8000 198 8034 212
rect 8000 143 8002 159
rect 8002 143 8034 159
rect 8000 125 8034 143
rect 10716 1246 10718 1280
rect 10718 1246 10750 1280
rect 10788 1246 10820 1280
rect 10820 1246 10822 1280
rect 10716 1173 10718 1207
rect 10718 1173 10750 1207
rect 10788 1173 10820 1207
rect 10820 1173 10822 1207
rect 10716 1100 10718 1134
rect 10718 1100 10750 1134
rect 10788 1100 10820 1134
rect 10820 1100 10822 1134
rect 10716 1027 10718 1061
rect 10718 1027 10750 1061
rect 10788 1027 10820 1061
rect 10820 1027 10822 1061
rect 10716 954 10718 988
rect 10718 954 10750 988
rect 10788 954 10820 988
rect 10820 954 10822 988
rect 10716 881 10718 915
rect 10718 881 10750 915
rect 10788 881 10820 915
rect 10820 881 10822 915
rect 10716 808 10718 842
rect 10718 808 10750 842
rect 10788 808 10820 842
rect 10820 808 10822 842
rect 10716 735 10718 769
rect 10718 735 10750 769
rect 10788 735 10820 769
rect 10820 735 10822 769
rect 10716 662 10718 696
rect 10718 662 10750 696
rect 10788 662 10820 696
rect 10820 662 10822 696
rect 10716 589 10718 623
rect 10718 589 10750 623
rect 10788 589 10820 623
rect 10820 589 10822 623
rect 10716 516 10718 550
rect 10718 516 10750 550
rect 10788 516 10820 550
rect 10820 516 10822 550
rect 10716 443 10718 477
rect 10718 443 10750 477
rect 10788 443 10820 477
rect 10820 443 10822 477
rect 10716 370 10718 404
rect 10718 370 10750 404
rect 10788 370 10820 404
rect 10820 370 10822 404
rect 10716 297 10718 331
rect 10718 297 10750 331
rect 10788 297 10820 331
rect 10820 297 10822 331
rect 10716 224 10718 258
rect 10718 224 10750 258
rect 10788 224 10820 258
rect 10820 224 10822 258
rect 10716 151 10718 185
rect 10718 151 10750 185
rect 10788 151 10820 185
rect 10820 151 10822 185
rect 8000 74 8002 86
rect 8002 74 8034 86
rect 8000 52 8034 74
rect 10716 108 10718 112
rect 10718 108 10750 112
rect 10788 108 10820 112
rect 10820 108 10822 112
rect 10716 78 10750 108
rect 10788 78 10822 108
<< metal1 >>
rect 366 39888 2599 39894
rect 366 39854 445 39888
rect 479 39854 518 39888
rect 552 39854 591 39888
rect 625 39854 664 39888
rect 698 39854 737 39888
rect 771 39854 810 39888
rect 844 39854 884 39888
rect 918 39854 958 39888
rect 992 39854 1032 39888
rect 1066 39854 1106 39888
rect 1140 39854 1216 39888
rect 1250 39854 1290 39888
rect 1324 39854 1364 39888
rect 1398 39854 1438 39888
rect 1472 39854 1512 39888
rect 1546 39854 1587 39888
rect 1621 39854 1662 39888
rect 1696 39854 1737 39888
rect 1771 39854 1812 39888
rect 1846 39854 1887 39888
rect 1921 39854 1962 39888
rect 1996 39854 2037 39888
rect 2071 39854 2112 39888
rect 2146 39854 2187 39888
rect 2221 39854 2262 39888
rect 2296 39854 2337 39888
rect 2371 39854 2412 39888
rect 2446 39854 2487 39888
rect 2521 39854 2599 39888
rect 366 39816 2599 39854
rect 366 39782 372 39816
rect 406 39782 444 39816
rect 478 39782 518 39816
rect 552 39782 591 39816
rect 625 39782 664 39816
rect 698 39782 737 39816
rect 771 39782 810 39816
rect 844 39782 884 39816
rect 918 39782 958 39816
rect 992 39782 1032 39816
rect 1066 39782 1106 39816
rect 1140 39782 1216 39816
rect 1250 39782 1290 39816
rect 1324 39782 1364 39816
rect 1398 39782 1438 39816
rect 1472 39782 1512 39816
rect 1546 39782 1587 39816
rect 1621 39782 1662 39816
rect 1696 39782 1737 39816
rect 1771 39782 1812 39816
rect 1846 39782 1887 39816
rect 1921 39782 1962 39816
rect 1996 39782 2037 39816
rect 2071 39782 2112 39816
rect 2146 39782 2187 39816
rect 2221 39782 2262 39816
rect 2296 39782 2337 39816
rect 2371 39782 2412 39816
rect 2446 39782 2487 39816
rect 366 39776 2487 39782
rect 366 39743 484 39776
rect 366 39709 372 39743
rect 406 39709 444 39743
rect 478 39709 484 39743
tri 484 39742 518 39776 nw
tri 2447 39742 2481 39776 ne
rect 2304 39719 2422 39725
rect 366 39670 484 39709
rect 366 39636 372 39670
rect 406 39636 444 39670
rect 478 39636 484 39670
rect 366 39597 484 39636
rect 366 39563 372 39597
rect 406 39563 444 39597
rect 478 39563 484 39597
rect 366 39524 484 39563
rect 366 39490 372 39524
rect 406 39490 444 39524
rect 478 39490 484 39524
rect 366 39451 484 39490
rect 366 39417 372 39451
rect 406 39417 444 39451
rect 478 39417 484 39451
rect 366 39378 484 39417
rect 366 39344 372 39378
rect 406 39344 444 39378
rect 478 39344 484 39378
rect 366 39305 484 39344
rect 366 39271 372 39305
rect 406 39271 444 39305
rect 478 39271 484 39305
rect 366 39232 484 39271
rect 366 39198 372 39232
rect 406 39198 444 39232
rect 478 39198 484 39232
rect 366 39159 484 39198
rect 366 39125 372 39159
rect 406 39125 444 39159
rect 478 39125 484 39159
rect 366 39086 484 39125
rect 366 39052 372 39086
rect 406 39052 444 39086
rect 478 39052 484 39086
rect 366 39013 484 39052
rect 366 38979 372 39013
rect 406 38979 444 39013
rect 478 38979 484 39013
rect 366 38940 484 38979
rect 366 38906 372 38940
rect 406 38906 444 38940
rect 478 38906 484 38940
rect 366 38867 484 38906
rect 366 38833 372 38867
rect 406 38833 444 38867
rect 478 38833 484 38867
rect 366 38794 484 38833
rect 366 38760 372 38794
rect 406 38760 444 38794
rect 478 38760 484 38794
rect 366 38721 484 38760
rect 366 38687 372 38721
rect 406 38687 444 38721
rect 478 38687 484 38721
rect 366 38648 484 38687
rect 366 38614 372 38648
rect 406 38614 444 38648
rect 478 38614 484 38648
rect 366 38575 484 38614
rect 366 38541 372 38575
rect 406 38541 444 38575
rect 478 38541 484 38575
rect 366 38502 484 38541
rect 366 38468 372 38502
rect 406 38468 444 38502
rect 478 38468 484 38502
rect 366 38429 484 38468
rect 366 38395 372 38429
rect 406 38395 444 38429
rect 478 38395 484 38429
rect 366 38356 484 38395
rect 366 38322 372 38356
rect 406 38322 444 38356
rect 478 38322 484 38356
rect 366 38283 484 38322
rect 366 38249 372 38283
rect 406 38249 444 38283
rect 478 38249 484 38283
rect 366 38210 484 38249
rect 366 38176 372 38210
rect 406 38176 444 38210
rect 478 38176 484 38210
rect 366 38137 484 38176
rect 366 38103 372 38137
rect 406 38103 444 38137
rect 478 38103 484 38137
rect 366 38064 484 38103
rect 366 38030 372 38064
rect 406 38030 444 38064
rect 478 38030 484 38064
rect 366 37991 484 38030
rect 366 37957 372 37991
rect 406 37957 444 37991
rect 478 37957 484 37991
rect 366 37918 484 37957
rect 366 37884 372 37918
rect 406 37884 444 37918
rect 478 37884 484 37918
rect 366 37845 484 37884
rect 366 37811 372 37845
rect 406 37811 444 37845
rect 478 37811 484 37845
rect 366 37772 484 37811
rect 366 37738 372 37772
rect 406 37738 444 37772
rect 478 37738 484 37772
rect 366 37699 484 37738
rect 366 37665 372 37699
rect 406 37665 444 37699
rect 478 37665 484 37699
rect 366 37626 484 37665
rect 366 37592 372 37626
rect 406 37592 444 37626
rect 478 37592 484 37626
rect 366 37553 484 37592
rect 366 37519 372 37553
rect 406 37519 444 37553
rect 478 37519 484 37553
rect 366 37480 484 37519
rect 366 37446 372 37480
rect 406 37446 444 37480
rect 478 37446 484 37480
rect 366 37407 484 37446
rect 366 37373 372 37407
rect 406 37373 444 37407
rect 478 37373 484 37407
rect 366 37334 484 37373
rect 366 436 372 37334
rect 478 436 484 37334
rect 512 39701 678 39713
rect 512 39667 566 39701
rect 600 39667 638 39701
rect 672 39667 678 39701
rect 512 39628 678 39667
rect 512 39594 566 39628
rect 600 39594 638 39628
rect 672 39594 678 39628
rect 512 39555 678 39594
rect 512 39521 566 39555
rect 600 39521 638 39555
rect 672 39521 678 39555
rect 2304 39667 2305 39719
rect 2357 39667 2369 39719
rect 2421 39667 2422 39719
rect 2304 39649 2422 39667
rect 2304 39597 2305 39649
rect 2357 39597 2369 39649
rect 2421 39597 2422 39649
rect 2304 39579 2422 39597
rect 2304 39527 2305 39579
rect 2357 39527 2369 39579
rect 2421 39527 2422 39579
rect 2304 39521 2422 39527
rect 512 39509 678 39521
rect 512 4455 628 39509
tri 628 39475 662 39509 nw
rect 656 26358 708 26364
rect 656 26294 708 26306
rect 656 6523 708 26242
rect 656 6459 708 6471
rect 656 4852 708 6407
rect 656 4788 708 4800
rect 656 4730 708 4736
rect 512 4333 628 4339
rect 366 398 484 436
rect 2481 2918 2487 39776
rect 2593 2918 2599 39816
rect 7994 39889 10828 39895
rect 7994 39855 8040 39889
rect 8074 39855 8116 39889
rect 8150 39855 8192 39889
rect 8226 39855 8268 39889
rect 8302 39855 8345 39889
rect 8379 39855 8422 39889
rect 8456 39855 8499 39889
rect 8533 39855 8576 39889
rect 8610 39855 8653 39889
rect 8687 39855 8730 39889
rect 8764 39855 8840 39889
rect 7994 39817 8840 39855
rect 7994 39783 8040 39817
rect 8074 39783 8116 39817
rect 8150 39783 8192 39817
rect 8226 39783 8268 39817
rect 8302 39783 8345 39817
rect 8379 39783 8422 39817
rect 8456 39783 8499 39817
rect 8533 39783 8576 39817
rect 8610 39783 8653 39817
rect 8687 39783 8730 39817
rect 8764 39783 8840 39817
rect 10458 39855 10497 39889
rect 10531 39855 10570 39889
rect 10604 39855 10643 39889
rect 10677 39855 10716 39889
rect 10750 39855 10828 39889
rect 10458 39817 10828 39855
rect 10458 39783 10497 39817
rect 10531 39783 10570 39817
rect 10604 39783 10643 39817
rect 10677 39783 10716 39817
rect 7994 39777 10716 39783
rect 7994 39745 8042 39777
tri 8042 39745 8074 39777 nw
rect 9746 39745 9792 39777
rect 7994 39742 8040 39745
tri 8040 39743 8042 39745 nw
rect 7994 39708 8000 39742
rect 8034 39708 8040 39742
rect 7994 39670 8040 39708
rect 7994 39636 8000 39670
rect 8034 39636 8040 39670
rect 5370 39614 7536 39620
rect 5370 39580 5402 39614
rect 5436 39580 5476 39614
rect 5510 39580 5550 39614
rect 5584 39580 5624 39614
rect 5658 39580 5698 39614
rect 5732 39580 5772 39614
rect 5806 39580 5846 39614
rect 5880 39580 5920 39614
rect 5954 39580 5994 39614
rect 6028 39580 6068 39614
rect 6102 39580 6142 39614
rect 6176 39580 6216 39614
rect 6250 39580 6290 39614
rect 6324 39580 6364 39614
rect 6398 39580 6438 39614
rect 6472 39580 6512 39614
rect 6546 39580 6586 39614
rect 6620 39580 6660 39614
rect 6694 39580 6734 39614
rect 6768 39580 6808 39614
rect 6842 39580 6882 39614
rect 6916 39580 6956 39614
rect 6990 39580 7030 39614
rect 7064 39580 7104 39614
rect 7138 39580 7178 39614
rect 7212 39580 7251 39614
rect 7285 39580 7324 39614
rect 7358 39580 7397 39614
rect 7431 39580 7470 39614
rect 7504 39580 7536 39614
rect 5370 39574 7536 39580
rect 5447 39564 7526 39574
tri 7526 39564 7536 39574 nw
rect 7994 39598 8040 39636
rect 7994 39564 8000 39598
rect 8034 39564 8040 39598
rect 5447 39533 7495 39564
tri 7495 39533 7526 39564 nw
rect 5447 39529 7491 39533
tri 7491 39529 7495 39533 nw
rect 5447 39526 7488 39529
tri 7488 39526 7491 39529 nw
rect 7994 39526 8040 39564
rect 5447 39521 7483 39526
tri 7483 39521 7488 39526 nw
rect 5447 39483 7470 39521
tri 7470 39508 7483 39521 nw
rect 7994 39492 8000 39526
rect 8034 39492 8040 39526
rect 8106 39719 8224 39725
rect 8106 39667 8107 39719
rect 8159 39667 8171 39719
rect 8223 39667 8224 39719
rect 8106 39649 8224 39667
rect 8106 39597 8107 39649
rect 8159 39597 8171 39649
rect 8223 39597 8224 39649
rect 8106 39579 8224 39597
rect 8106 39527 8107 39579
rect 8159 39527 8171 39579
rect 8223 39527 8224 39579
rect 8106 39521 8224 39527
rect 9558 39719 9676 39725
rect 9558 39667 9559 39719
rect 9611 39667 9623 39719
rect 9675 39667 9676 39719
rect 9558 39649 9676 39667
rect 9558 39597 9559 39649
rect 9611 39597 9623 39649
rect 9675 39597 9676 39649
rect 9558 39579 9676 39597
rect 9558 39527 9559 39579
rect 9611 39527 9623 39579
rect 9675 39527 9676 39579
rect 9558 39521 9676 39527
rect 9746 39711 9752 39745
rect 9786 39711 9792 39745
tri 10676 39743 10710 39777 ne
rect 9746 39673 9792 39711
rect 9746 39639 9752 39673
rect 9786 39639 9792 39673
rect 9746 39601 9792 39639
rect 9746 39567 9752 39601
rect 9786 39567 9792 39601
rect 9746 39529 9792 39567
rect 5447 39452 6207 39483
rect 7994 39454 8040 39492
rect 5447 39420 6209 39452
tri 6209 39420 6241 39452 nw
rect 7994 39420 8000 39454
rect 8034 39420 8040 39454
rect 5447 39270 6207 39420
tri 6207 39418 6209 39420 nw
rect 7994 39382 8040 39420
rect 5447 39218 5604 39270
rect 5656 39218 6207 39270
rect 5447 39206 6207 39218
rect 5447 39154 5604 39206
rect 5656 39154 6207 39206
rect 5447 39142 6207 39154
rect 5447 39090 5604 39142
rect 5656 39090 6207 39142
rect 5447 39078 6207 39090
rect 5447 39026 5604 39078
rect 5656 39068 6207 39078
rect 7526 39356 7572 39368
rect 7526 39322 7532 39356
rect 7566 39322 7572 39356
rect 7526 39284 7572 39322
rect 7526 39250 7532 39284
rect 7566 39250 7572 39284
rect 7526 39212 7572 39250
rect 7526 39178 7532 39212
rect 7566 39178 7572 39212
rect 7526 39140 7572 39178
rect 7526 39106 7532 39140
rect 7566 39106 7572 39140
tri 6207 39068 6215 39076 sw
rect 7526 39068 7572 39106
rect 5656 39042 6215 39068
tri 6215 39042 6241 39068 sw
rect 5656 39026 6207 39042
rect 5447 39014 6207 39026
rect 5447 38962 5604 39014
rect 5656 38962 6207 39014
rect 7526 39034 7532 39068
rect 7566 39034 7572 39068
rect 7526 38996 7572 39034
tri 6207 38962 6241 38996 nw
rect 7526 38962 7532 38996
rect 7566 38962 7572 38996
rect 5447 38950 6207 38962
rect 5447 38898 5604 38950
rect 5656 38898 6207 38950
rect 5447 38886 6207 38898
rect 5447 38834 5604 38886
rect 5656 38834 6207 38886
rect 5447 38822 6207 38834
rect 5447 38770 5604 38822
rect 5656 38770 6207 38822
rect 5447 38758 6207 38770
rect 5447 38706 5604 38758
rect 5656 38706 6207 38758
rect 5447 38694 6207 38706
rect 5447 38642 5604 38694
rect 5656 38642 6207 38694
rect 5447 38630 6207 38642
rect 5447 38578 5604 38630
rect 5656 38602 6207 38630
rect 7526 38924 7572 38962
rect 7526 38890 7532 38924
rect 7566 38890 7572 38924
rect 7526 38852 7572 38890
rect 7526 38818 7532 38852
rect 7566 38818 7572 38852
rect 7526 38780 7572 38818
rect 7526 38746 7532 38780
rect 7566 38746 7572 38780
rect 7526 38708 7572 38746
rect 7526 38674 7532 38708
rect 7566 38674 7572 38708
rect 7526 38636 7572 38674
tri 6207 38602 6225 38620 sw
rect 7526 38602 7532 38636
rect 7566 38602 7572 38636
rect 5656 38593 6225 38602
tri 6225 38593 6234 38602 sw
rect 5656 38590 6234 38593
tri 6234 38590 6237 38593 sw
rect 5656 38586 6237 38590
tri 6237 38586 6241 38590 sw
rect 5656 38578 6207 38586
rect 5447 38566 6207 38578
rect 5447 38514 5604 38566
rect 5656 38540 6207 38566
rect 7526 38564 7572 38602
rect 5656 38530 6231 38540
tri 6231 38530 6241 38540 nw
rect 7526 38530 7532 38564
rect 7566 38530 7572 38564
rect 5656 38521 6222 38530
tri 6222 38521 6231 38530 nw
rect 5656 38518 6219 38521
tri 6219 38518 6222 38521 nw
rect 5656 38514 6207 38518
rect 5447 38502 6207 38514
tri 6207 38506 6219 38518 nw
rect 5447 38450 5604 38502
rect 5656 38450 6207 38502
rect 5447 38438 6207 38450
rect 5447 38386 5604 38438
rect 5656 38386 6207 38438
rect 5447 38374 6207 38386
rect 5447 38322 5604 38374
rect 5656 38322 6207 38374
rect 5447 38310 6207 38322
rect 5447 38258 5604 38310
rect 5656 38258 6207 38310
rect 5447 38246 6207 38258
rect 5447 38194 5604 38246
rect 5656 38194 6207 38246
rect 5447 38182 6207 38194
rect 5447 38130 5604 38182
rect 5656 38161 6207 38182
rect 7526 38492 7572 38530
rect 7526 38458 7532 38492
rect 7566 38458 7572 38492
rect 7526 38420 7572 38458
rect 7526 38386 7532 38420
rect 7566 38386 7572 38420
rect 7526 38348 7572 38386
rect 7526 38314 7532 38348
rect 7566 38314 7572 38348
rect 7526 38276 7572 38314
rect 7526 38242 7532 38276
rect 7566 38242 7572 38276
rect 7526 38204 7572 38242
rect 7526 38170 7532 38204
rect 7566 38170 7572 38204
tri 6207 38161 6210 38164 sw
rect 5656 38158 6210 38161
tri 6210 38158 6213 38161 sw
rect 5656 38132 6213 38158
tri 6213 38132 6239 38158 sw
rect 7526 38132 7572 38170
rect 5656 38130 6239 38132
tri 6239 38130 6241 38132 sw
rect 5447 38118 6207 38130
rect 5447 38066 5604 38118
rect 5656 38084 6207 38118
rect 7526 38098 7532 38132
rect 7566 38098 7572 38132
rect 5656 38066 6217 38084
rect 5447 38060 6217 38066
tri 6217 38060 6241 38084 nw
rect 7526 38060 7572 38098
rect 5447 38054 6207 38060
rect 5447 38002 5604 38054
rect 5656 38002 6207 38054
tri 6207 38050 6217 38060 nw
rect 5447 37990 6207 38002
rect 5447 37938 5604 37990
rect 5656 37938 6207 37990
rect 5447 37926 6207 37938
rect 5447 37874 5604 37926
rect 5656 37874 6207 37926
rect 5447 37862 6207 37874
rect 5447 37810 5604 37862
rect 5656 37810 6207 37862
rect 5447 37798 6207 37810
rect 5447 37746 5604 37798
rect 5656 37746 6207 37798
rect 5447 37734 6207 37746
rect 5447 37682 5604 37734
rect 5656 37700 6207 37734
rect 7526 38026 7532 38060
rect 7566 38026 7572 38060
rect 7526 37988 7572 38026
rect 7526 37954 7532 37988
rect 7566 37954 7572 37988
rect 7526 37916 7572 37954
rect 7526 37882 7532 37916
rect 7566 37882 7572 37916
rect 7526 37844 7572 37882
rect 7526 37810 7532 37844
rect 7566 37810 7572 37844
rect 7526 37772 7572 37810
rect 7526 37738 7532 37772
rect 7566 37738 7572 37772
tri 6207 37700 6215 37708 sw
rect 7526 37700 7572 37738
rect 5656 37682 6215 37700
rect 5447 37674 6215 37682
tri 6215 37674 6241 37700 sw
rect 5447 37670 6207 37674
rect 5447 37618 5604 37670
rect 5656 37618 6207 37670
rect 7526 37666 7532 37700
rect 7566 37666 7572 37700
rect 7526 37628 7572 37666
rect 5447 37606 6207 37618
rect 5447 37554 5604 37606
rect 5656 37554 6207 37606
tri 6207 37594 6241 37628 nw
rect 7526 37594 7532 37628
rect 7566 37594 7572 37628
rect 5447 37542 6207 37554
rect 5447 37490 5604 37542
rect 5656 37490 6207 37542
rect 5447 37478 6207 37490
rect 5447 37426 5604 37478
rect 5656 37426 6207 37478
rect 5447 37414 6207 37426
rect 5447 37362 5604 37414
rect 5656 37362 6207 37414
rect 5447 37350 6207 37362
rect 5447 37298 5604 37350
rect 5656 37298 6207 37350
rect 5447 37286 6207 37298
rect 5447 37234 5604 37286
rect 5656 37234 6207 37286
rect 7526 37556 7572 37594
rect 7526 37522 7532 37556
rect 7566 37522 7572 37556
rect 7526 37484 7572 37522
rect 7526 37450 7532 37484
rect 7566 37450 7572 37484
rect 7526 37412 7572 37450
rect 7526 37378 7532 37412
rect 7566 37378 7572 37412
rect 7526 37340 7572 37378
rect 7526 37306 7532 37340
rect 7566 37306 7572 37340
rect 7526 37267 7572 37306
rect 5447 37233 6207 37234
tri 6207 37233 6226 37252 sw
rect 7526 37233 7532 37267
rect 7566 37233 7572 37267
rect 5447 37225 6226 37233
tri 6226 37225 6234 37233 sw
rect 5447 37222 6234 37225
tri 6234 37222 6237 37225 sw
rect 5447 37170 5604 37222
rect 5656 37218 6237 37222
tri 6237 37218 6241 37222 sw
rect 5656 37172 6207 37218
rect 7526 37194 7572 37233
rect 5656 37170 6229 37172
rect 5447 37160 6229 37170
tri 6229 37160 6241 37172 nw
rect 7526 37160 7532 37194
rect 7566 37160 7572 37194
rect 5447 37158 6222 37160
rect 5447 37106 5604 37158
rect 5656 37153 6222 37158
tri 6222 37153 6229 37160 nw
rect 5656 37150 6219 37153
tri 6219 37150 6222 37153 nw
rect 5656 37106 6207 37150
tri 6207 37138 6219 37150 nw
rect 5447 37094 6207 37106
rect 5447 37042 5604 37094
rect 5656 37042 6207 37094
rect 5447 37030 6207 37042
rect 5447 36978 5604 37030
rect 5656 36978 6207 37030
rect 5447 36966 6207 36978
rect 5447 36914 5604 36966
rect 5656 36914 6207 36966
rect 5447 36902 6207 36914
rect 5447 36850 5604 36902
rect 5656 36850 6207 36902
rect 5447 36838 6207 36850
rect 5447 36786 5604 36838
rect 5656 36795 6207 36838
rect 7526 37121 7572 37160
rect 7526 37087 7532 37121
rect 7566 37087 7572 37121
rect 7526 37048 7572 37087
rect 7526 37014 7532 37048
rect 7566 37014 7572 37048
rect 7526 36975 7572 37014
rect 7526 36941 7532 36975
rect 7566 36941 7572 36975
rect 7526 36902 7572 36941
rect 7526 36868 7532 36902
rect 7566 36868 7572 36902
rect 7526 36829 7572 36868
tri 6207 36795 6208 36796 sw
rect 7526 36795 7532 36829
rect 7566 36795 7572 36829
rect 5656 36793 6208 36795
tri 6208 36793 6210 36795 sw
rect 5656 36790 6210 36793
tri 6210 36790 6213 36793 sw
rect 5656 36786 6213 36790
rect 5447 36774 6213 36786
rect 5447 36722 5604 36774
rect 5656 36762 6213 36774
tri 6213 36762 6241 36790 sw
rect 5656 36722 6207 36762
rect 5447 36716 6207 36722
rect 7526 36756 7572 36795
rect 7526 36722 7532 36756
rect 7566 36722 7572 36756
rect 5447 36710 6209 36716
rect 5447 36658 5604 36710
rect 5656 36684 6209 36710
tri 6209 36684 6241 36716 nw
rect 5656 36683 6208 36684
tri 6208 36683 6209 36684 nw
rect 7526 36683 7572 36722
rect 5656 36658 6207 36683
tri 6207 36682 6208 36683 nw
rect 5447 36646 6207 36658
rect 5447 36594 5604 36646
rect 5656 36594 6207 36646
rect 5447 36582 6207 36594
rect 5447 36530 5604 36582
rect 5656 36530 6207 36582
rect 5447 36518 6207 36530
rect 5447 36466 5604 36518
rect 5656 36466 6207 36518
rect 5447 36454 6207 36466
rect 5447 36402 5604 36454
rect 5656 36402 6207 36454
rect 5447 36390 6207 36402
rect 5447 36338 5604 36390
rect 5656 36338 6207 36390
rect 7526 36649 7532 36683
rect 7566 36649 7572 36683
rect 7526 36610 7572 36649
rect 7526 36576 7532 36610
rect 7566 36576 7572 36610
rect 7526 36537 7572 36576
rect 7526 36503 7532 36537
rect 7566 36503 7572 36537
rect 7526 36464 7572 36503
rect 7526 36430 7532 36464
rect 7566 36430 7572 36464
rect 7526 36391 7572 36430
rect 7526 36357 7532 36391
rect 7566 36357 7572 36391
rect 5447 36326 6207 36338
rect 5447 36274 5604 36326
rect 5656 36324 6207 36326
tri 6207 36324 6223 36340 sw
rect 5656 36318 6223 36324
tri 6223 36318 6229 36324 sw
rect 7526 36318 7572 36357
rect 5656 36306 6229 36318
tri 6229 36306 6241 36318 sw
rect 5656 36274 6207 36306
rect 5447 36262 6207 36274
rect 5447 36210 5604 36262
rect 5656 36260 6207 36262
rect 7526 36284 7532 36318
rect 7566 36284 7572 36318
rect 5656 36252 6233 36260
tri 6233 36252 6241 36260 nw
rect 5656 36245 6226 36252
tri 6226 36245 6233 36252 nw
rect 7526 36245 7572 36284
rect 5656 36210 6207 36245
tri 6207 36226 6226 36245 nw
rect 5447 36198 6207 36210
rect 5447 36146 5604 36198
rect 5656 36146 6207 36198
rect 5447 36134 6207 36146
rect 5447 36082 5604 36134
rect 5656 36082 6207 36134
rect 5447 36070 6207 36082
rect 5447 36018 5604 36070
rect 5656 36018 6207 36070
rect 5447 36006 6207 36018
rect 5447 35954 5604 36006
rect 5656 35954 6207 36006
rect 5447 35942 6207 35954
rect 5447 35890 5604 35942
rect 5656 35890 6207 35942
rect 5447 35880 6207 35890
rect 7526 36211 7532 36245
rect 7566 36211 7572 36245
rect 7526 36172 7572 36211
rect 7526 36138 7532 36172
rect 7566 36138 7572 36172
rect 7526 36099 7572 36138
rect 7526 36065 7532 36099
rect 7566 36065 7572 36099
rect 7526 36026 7572 36065
rect 7526 35992 7532 36026
rect 7566 35992 7572 36026
rect 7526 35953 7572 35992
rect 7526 35919 7532 35953
rect 7566 35919 7572 35953
tri 6207 35880 6211 35884 sw
rect 7526 35880 7572 35919
rect 5447 35878 6211 35880
rect 5447 35826 5604 35878
rect 5656 35850 6211 35878
tri 6211 35850 6241 35880 sw
rect 5656 35826 6207 35850
rect 5447 35814 6207 35826
rect 5447 35762 5604 35814
rect 5656 35804 6207 35814
rect 7526 35846 7532 35880
rect 7566 35846 7572 35880
rect 7526 35807 7572 35846
rect 5656 35773 6210 35804
tri 6210 35773 6241 35804 nw
rect 7526 35773 7532 35807
rect 7566 35773 7572 35807
rect 5656 35762 6207 35773
tri 6207 35770 6210 35773 nw
rect 5447 35750 6207 35762
rect 5447 35698 5604 35750
rect 5656 35698 6207 35750
rect 5447 35686 6207 35698
rect 5447 35634 5604 35686
rect 5656 35634 6207 35686
rect 5447 35622 6207 35634
rect 5447 35570 5604 35622
rect 5656 35570 6207 35622
rect 5447 35558 6207 35570
rect 5447 35506 5604 35558
rect 5656 35506 6207 35558
rect 5447 35494 6207 35506
rect 5447 35442 5604 35494
rect 5656 35442 6207 35494
rect 5447 35430 6207 35442
rect 5447 35378 5604 35430
rect 5656 35408 6207 35430
rect 7526 35734 7572 35773
rect 7526 35700 7532 35734
rect 7566 35700 7572 35734
rect 7526 35661 7572 35700
rect 7526 35627 7532 35661
rect 7566 35627 7572 35661
rect 7526 35588 7572 35627
rect 7526 35554 7532 35588
rect 7566 35554 7572 35588
rect 7526 35515 7572 35554
rect 7526 35481 7532 35515
rect 7566 35481 7572 35515
rect 7526 35442 7572 35481
tri 6207 35408 6227 35428 sw
rect 7526 35408 7532 35442
rect 7566 35408 7572 35442
rect 5656 35394 6227 35408
tri 6227 35394 6241 35408 sw
rect 5656 35378 6207 35394
rect 5447 35366 6207 35378
rect 5447 35314 5604 35366
rect 5656 35348 6207 35366
rect 7526 35369 7572 35408
rect 5656 35335 6228 35348
tri 6228 35335 6241 35348 nw
rect 7526 35335 7532 35369
rect 7566 35335 7572 35369
rect 5656 35316 6209 35335
tri 6209 35316 6228 35335 nw
rect 5656 35314 6207 35316
tri 6207 35314 6209 35316 nw
rect 5447 35302 6207 35314
rect 5447 35250 5604 35302
rect 5656 35250 6207 35302
rect 5447 35238 6207 35250
rect 5447 35186 5604 35238
rect 5656 35186 6207 35238
rect 5447 35174 6207 35186
rect 5447 35122 5604 35174
rect 5656 35122 6207 35174
rect 5447 35110 6207 35122
rect 5447 35058 5604 35110
rect 5656 35058 6207 35110
rect 5447 35046 6207 35058
rect 5447 34994 5604 35046
rect 5656 34994 6207 35046
rect 5447 34982 6207 34994
rect 5447 34930 5604 34982
rect 5656 34970 6207 34982
rect 7526 35296 7572 35335
rect 7526 35262 7532 35296
rect 7566 35262 7572 35296
rect 7526 35223 7572 35262
rect 7526 35189 7532 35223
rect 7566 35189 7572 35223
rect 7526 35150 7572 35189
rect 7526 35116 7532 35150
rect 7566 35116 7572 35150
rect 7526 35077 7572 35116
rect 7526 35043 7532 35077
rect 7566 35043 7572 35077
rect 7526 35007 7572 35043
rect 7994 39348 8000 39382
rect 8034 39348 8040 39382
rect 7994 39310 8040 39348
rect 7994 39276 8000 39310
rect 8034 39276 8040 39310
rect 7994 39238 8040 39276
rect 7994 39204 8000 39238
rect 8034 39204 8040 39238
rect 7994 39166 8040 39204
rect 7994 39132 8000 39166
rect 8034 39132 8040 39166
rect 7994 39094 8040 39132
rect 7994 39060 8000 39094
rect 8034 39060 8040 39094
rect 7994 39022 8040 39060
rect 7994 38988 8000 39022
rect 8034 38988 8040 39022
rect 7994 38950 8040 38988
rect 7994 38916 8000 38950
rect 8034 38916 8040 38950
rect 7994 38878 8040 38916
rect 7994 38844 8000 38878
rect 8034 38844 8040 38878
rect 7994 38806 8040 38844
rect 7994 38772 8000 38806
rect 8034 38772 8040 38806
rect 7994 38734 8040 38772
rect 7994 38700 8000 38734
rect 8034 38700 8040 38734
rect 7994 38662 8040 38700
rect 7994 38628 8000 38662
rect 8034 38628 8040 38662
rect 7994 38590 8040 38628
rect 7994 38556 8000 38590
rect 8034 38556 8040 38590
rect 7994 38518 8040 38556
rect 7994 38484 8000 38518
rect 8034 38484 8040 38518
rect 7994 38446 8040 38484
rect 7994 38412 8000 38446
rect 8034 38412 8040 38446
rect 7994 38374 8040 38412
rect 7994 38340 8000 38374
rect 8034 38340 8040 38374
rect 7994 38302 8040 38340
rect 7994 38268 8000 38302
rect 8034 38268 8040 38302
rect 7994 38230 8040 38268
rect 7994 38196 8000 38230
rect 8034 38196 8040 38230
rect 7994 38158 8040 38196
rect 7994 38124 8000 38158
rect 8034 38124 8040 38158
rect 7994 38086 8040 38124
rect 7994 38052 8000 38086
rect 8034 38052 8040 38086
rect 7994 38014 8040 38052
rect 7994 37980 8000 38014
rect 8034 37980 8040 38014
rect 7994 37942 8040 37980
rect 7994 37908 8000 37942
rect 8034 37908 8040 37942
rect 7994 37870 8040 37908
rect 7994 37836 8000 37870
rect 8034 37836 8040 37870
rect 7994 37798 8040 37836
rect 7994 37764 8000 37798
rect 8034 37764 8040 37798
rect 7994 37726 8040 37764
rect 7994 37692 8000 37726
rect 8034 37692 8040 37726
rect 7994 37654 8040 37692
rect 7994 37620 8000 37654
rect 8034 37620 8040 37654
rect 7994 37582 8040 37620
rect 7994 37548 8000 37582
rect 8034 37548 8040 37582
rect 7994 37510 8040 37548
rect 7994 37476 8000 37510
rect 8034 37476 8040 37510
rect 7994 37438 8040 37476
rect 7994 37404 8000 37438
rect 8034 37404 8040 37438
rect 7994 37366 8040 37404
rect 7994 37332 8000 37366
rect 8034 37332 8040 37366
rect 7994 37294 8040 37332
rect 7994 37260 8000 37294
rect 8034 37260 8040 37294
rect 7994 37222 8040 37260
rect 7994 37188 8000 37222
rect 8034 37188 8040 37222
rect 7994 37150 8040 37188
rect 7994 37116 8000 37150
rect 8034 37116 8040 37150
rect 7994 37078 8040 37116
rect 7994 37044 8000 37078
rect 8034 37044 8040 37078
rect 7994 37006 8040 37044
rect 7994 36972 8000 37006
rect 8034 36972 8040 37006
rect 7994 36934 8040 36972
rect 7994 36900 8000 36934
rect 8034 36900 8040 36934
rect 7994 36862 8040 36900
rect 7994 36828 8000 36862
rect 8034 36828 8040 36862
rect 7994 36790 8040 36828
rect 7994 36756 8000 36790
rect 8034 36756 8040 36790
rect 7994 36718 8040 36756
rect 7994 36684 8000 36718
rect 8034 36684 8040 36718
rect 7994 36646 8040 36684
rect 7994 36612 8000 36646
rect 8034 36612 8040 36646
rect 7994 36574 8040 36612
rect 7994 36540 8000 36574
rect 8034 36540 8040 36574
rect 7994 36502 8040 36540
rect 7994 36468 8000 36502
rect 8034 36468 8040 36502
rect 7994 36430 8040 36468
rect 7994 36396 8000 36430
rect 8034 36396 8040 36430
rect 7994 36358 8040 36396
rect 7994 36324 8000 36358
rect 8034 36324 8040 36358
rect 7994 36286 8040 36324
rect 7994 36252 8000 36286
rect 8034 36252 8040 36286
rect 7994 36214 8040 36252
rect 7994 36180 8000 36214
rect 8034 36180 8040 36214
rect 7994 36142 8040 36180
rect 7994 36108 8000 36142
rect 8034 36108 8040 36142
rect 7994 36070 8040 36108
rect 7994 36036 8000 36070
rect 8034 36036 8040 36070
rect 7994 35998 8040 36036
rect 7994 35964 8000 35998
rect 8034 35964 8040 35998
rect 7994 35926 8040 35964
rect 7994 35892 8000 35926
rect 8034 35892 8040 35926
rect 7994 35854 8040 35892
rect 7994 35820 8000 35854
rect 8034 35820 8040 35854
rect 7994 35782 8040 35820
rect 7994 35748 8000 35782
rect 8034 35748 8040 35782
rect 7994 35710 8040 35748
rect 7994 35676 8000 35710
rect 8034 35676 8040 35710
rect 7994 35638 8040 35676
rect 7994 35604 8000 35638
rect 8034 35604 8040 35638
rect 7994 35566 8040 35604
rect 7994 35532 8000 35566
rect 8034 35532 8040 35566
rect 7994 35494 8040 35532
rect 7994 35460 8000 35494
rect 8034 35460 8040 35494
rect 7994 35422 8040 35460
rect 7994 35388 8000 35422
rect 8034 35388 8040 35422
rect 7994 35350 8040 35388
rect 7994 35316 8000 35350
rect 8034 35316 8040 35350
rect 7994 35278 8040 35316
rect 7994 35244 8000 35278
rect 8034 35244 8040 35278
rect 7994 35206 8040 35244
rect 7994 35172 8000 35206
rect 8034 35172 8040 35206
rect 7994 35134 8040 35172
rect 7994 35100 8000 35134
rect 8034 35100 8040 35134
rect 7994 35062 8040 35100
rect 7994 35028 8000 35062
rect 8034 35028 8040 35062
tri 7572 35007 7578 35013 sw
rect 7526 35004 7578 35007
rect 7526 35001 7532 35004
rect 7566 35001 7578 35004
tri 6207 34970 6209 34972 sw
rect 5656 34956 6209 34970
tri 6209 34956 6223 34970 sw
rect 5656 34938 6223 34956
tri 6223 34938 6241 34956 sw
rect 5656 34930 6207 34938
rect 5447 34918 6207 34930
rect 5447 34866 5604 34918
rect 5656 34892 6207 34918
rect 7526 34937 7578 34949
rect 5656 34884 6233 34892
tri 6233 34884 6241 34892 nw
rect 5656 34866 6207 34884
rect 5447 34854 6207 34866
tri 6207 34858 6233 34884 nw
rect 7526 34879 7578 34885
rect 7526 34858 7572 34879
tri 7572 34873 7578 34879 nw
rect 7994 34990 8040 35028
rect 9746 39495 9752 39529
rect 9786 39495 9792 39529
rect 10553 39719 10671 39725
rect 10553 39667 10554 39719
rect 10606 39667 10618 39719
rect 10670 39667 10671 39719
rect 10553 39649 10671 39667
rect 10553 39597 10554 39649
rect 10606 39597 10618 39649
rect 10670 39597 10671 39649
rect 10553 39579 10671 39597
rect 10553 39527 10554 39579
rect 10606 39527 10618 39579
rect 10670 39527 10671 39579
rect 10553 39521 10671 39527
rect 9746 39457 9792 39495
rect 9746 39423 9752 39457
rect 9786 39423 9792 39457
rect 9746 39385 9792 39423
rect 9746 39351 9752 39385
rect 9786 39351 9792 39385
rect 9746 39313 9792 39351
rect 9746 39279 9752 39313
rect 9786 39279 9792 39313
rect 9746 39241 9792 39279
rect 9746 39207 9752 39241
rect 9786 39207 9792 39241
rect 9746 39169 9792 39207
rect 9746 39135 9752 39169
rect 9786 39135 9792 39169
rect 9746 39097 9792 39135
rect 9746 39063 9752 39097
rect 9786 39063 9792 39097
rect 9746 39025 9792 39063
rect 9746 38991 9752 39025
rect 9786 38991 9792 39025
rect 9746 38953 9792 38991
rect 9746 38919 9752 38953
rect 9786 38919 9792 38953
rect 9746 38881 9792 38919
rect 9746 38847 9752 38881
rect 9786 38847 9792 38881
rect 9746 38809 9792 38847
rect 9746 38775 9752 38809
rect 9786 38775 9792 38809
rect 9746 38737 9792 38775
rect 9746 38703 9752 38737
rect 9786 38703 9792 38737
rect 9746 38665 9792 38703
rect 9746 38631 9752 38665
rect 9786 38631 9792 38665
rect 9746 38593 9792 38631
rect 9746 38559 9752 38593
rect 9786 38559 9792 38593
rect 9746 38521 9792 38559
rect 9746 38487 9752 38521
rect 9786 38487 9792 38521
rect 9746 38449 9792 38487
rect 9746 38415 9752 38449
rect 9786 38415 9792 38449
rect 9746 38377 9792 38415
rect 9746 38343 9752 38377
rect 9786 38343 9792 38377
rect 9746 38305 9792 38343
rect 9746 38271 9752 38305
rect 9786 38271 9792 38305
rect 9746 38233 9792 38271
rect 9746 38199 9752 38233
rect 9786 38199 9792 38233
rect 9746 38161 9792 38199
rect 9746 38127 9752 38161
rect 9786 38127 9792 38161
rect 9746 38089 9792 38127
rect 9746 38055 9752 38089
rect 9786 38055 9792 38089
rect 9746 38017 9792 38055
rect 9746 37983 9752 38017
rect 9786 37983 9792 38017
rect 9746 37945 9792 37983
rect 9746 37911 9752 37945
rect 9786 37911 9792 37945
rect 9746 37873 9792 37911
rect 9746 37839 9752 37873
rect 9786 37839 9792 37873
rect 9746 37801 9792 37839
rect 9746 37767 9752 37801
rect 9786 37767 9792 37801
rect 9746 37729 9792 37767
rect 9746 37695 9752 37729
rect 9786 37695 9792 37729
rect 9746 37657 9792 37695
rect 9746 37623 9752 37657
rect 9786 37623 9792 37657
rect 9746 37585 9792 37623
rect 9746 37551 9752 37585
rect 9786 37551 9792 37585
rect 9746 37513 9792 37551
rect 9746 37479 9752 37513
rect 9786 37479 9792 37513
rect 9746 37441 9792 37479
rect 9746 37407 9752 37441
rect 9786 37407 9792 37441
rect 9746 37369 9792 37407
rect 9746 37335 9752 37369
rect 9786 37335 9792 37369
rect 9746 37297 9792 37335
rect 9746 37263 9752 37297
rect 9786 37263 9792 37297
rect 9746 37225 9792 37263
rect 9746 37191 9752 37225
rect 9786 37191 9792 37225
rect 9746 37153 9792 37191
rect 9746 37119 9752 37153
rect 9786 37119 9792 37153
rect 9746 37081 9792 37119
rect 9746 37047 9752 37081
rect 9786 37047 9792 37081
rect 9746 37009 9792 37047
rect 9746 36975 9752 37009
rect 9786 36975 9792 37009
rect 9746 36937 9792 36975
rect 9746 36903 9752 36937
rect 9786 36903 9792 36937
rect 9746 36865 9792 36903
rect 9746 36831 9752 36865
rect 9786 36831 9792 36865
rect 9746 36793 9792 36831
rect 9746 36759 9752 36793
rect 9786 36759 9792 36793
rect 9746 36721 9792 36759
rect 9746 36687 9752 36721
rect 9786 36687 9792 36721
rect 9746 36649 9792 36687
rect 9746 36615 9752 36649
rect 9786 36615 9792 36649
rect 9746 36577 9792 36615
rect 9746 36543 9752 36577
rect 9786 36543 9792 36577
rect 9746 36505 9792 36543
rect 9746 36471 9752 36505
rect 9786 36471 9792 36505
rect 9746 36433 9792 36471
rect 9746 36399 9752 36433
rect 9786 36399 9792 36433
rect 9746 36361 9792 36399
rect 9746 36327 9752 36361
rect 9786 36327 9792 36361
rect 9746 36289 9792 36327
rect 9746 36255 9752 36289
rect 9786 36255 9792 36289
rect 9746 36217 9792 36255
rect 9746 36183 9752 36217
rect 9786 36183 9792 36217
rect 9746 36145 9792 36183
rect 9746 36111 9752 36145
rect 9786 36111 9792 36145
rect 9746 36073 9792 36111
rect 9746 36039 9752 36073
rect 9786 36039 9792 36073
rect 9746 36001 9792 36039
rect 9746 35967 9752 36001
rect 9786 35967 9792 36001
rect 9746 35929 9792 35967
rect 9746 35895 9752 35929
rect 9786 35895 9792 35929
rect 9746 35857 9792 35895
rect 9746 35823 9752 35857
rect 9786 35823 9792 35857
rect 9746 35785 9792 35823
rect 9746 35751 9752 35785
rect 9786 35751 9792 35785
rect 9746 35713 9792 35751
rect 9746 35679 9752 35713
rect 9786 35679 9792 35713
rect 9746 35641 9792 35679
rect 9746 35607 9752 35641
rect 9786 35607 9792 35641
rect 9746 35569 9792 35607
rect 9746 35535 9752 35569
rect 9786 35535 9792 35569
rect 9746 35497 9792 35535
rect 9746 35463 9752 35497
rect 9786 35463 9792 35497
rect 9746 35425 9792 35463
rect 9746 35391 9752 35425
rect 9786 35391 9792 35425
rect 9746 35353 9792 35391
rect 9746 35319 9752 35353
rect 9786 35319 9792 35353
rect 9746 35281 9792 35319
rect 9746 35247 9752 35281
rect 9786 35247 9792 35281
rect 9746 35209 9792 35247
rect 9746 35175 9752 35209
rect 9786 35175 9792 35209
rect 9746 35137 9792 35175
rect 9746 35103 9752 35137
rect 9786 35103 9792 35137
rect 9746 35065 9792 35103
rect 9746 35031 9752 35065
rect 9786 35031 9792 35065
rect 7994 34956 8000 34990
rect 8034 34956 8040 34990
rect 7994 34918 8040 34956
rect 7994 34884 8000 34918
rect 8034 34884 8040 34918
rect 5447 34802 5604 34854
rect 5656 34802 6207 34854
rect 5447 34790 6207 34802
rect 5447 34738 5604 34790
rect 5656 34738 6207 34790
rect 5447 34726 6207 34738
rect 5447 34674 5604 34726
rect 5656 34674 6207 34726
rect 5447 34662 6207 34674
rect 5447 34610 5604 34662
rect 5656 34610 6207 34662
rect 5447 34598 6207 34610
rect 5447 34546 5604 34598
rect 5656 34546 6207 34598
rect 5447 34534 6207 34546
rect 5447 34482 5604 34534
rect 5656 34493 6207 34534
rect 7526 34824 7532 34858
rect 7566 34824 7572 34858
rect 7526 34785 7572 34824
rect 7526 34751 7532 34785
rect 7566 34751 7572 34785
rect 7526 34712 7572 34751
rect 7526 34678 7532 34712
rect 7566 34678 7572 34712
rect 7526 34639 7572 34678
rect 7526 34605 7532 34639
rect 7566 34605 7572 34639
rect 7526 34566 7572 34605
rect 7526 34532 7532 34566
rect 7566 34532 7572 34566
tri 6207 34493 6230 34516 sw
rect 7526 34493 7572 34532
rect 5656 34482 6230 34493
tri 6230 34482 6241 34493 sw
rect 5447 34470 6207 34482
rect 5447 34418 5604 34470
rect 5656 34436 6207 34470
rect 7526 34459 7532 34493
rect 7566 34459 7572 34493
rect 5656 34420 6225 34436
tri 6225 34420 6241 34436 nw
rect 7526 34420 7572 34459
rect 5656 34418 6207 34420
rect 5447 34406 6207 34418
rect 5447 34354 5604 34406
rect 5656 34354 6207 34406
tri 6207 34402 6225 34420 nw
rect 5447 34342 6207 34354
rect 5447 34290 5604 34342
rect 5656 34290 6207 34342
rect 5447 34278 6207 34290
rect 5447 34226 5604 34278
rect 5656 34226 6207 34278
rect 5447 34214 6207 34226
rect 5447 34162 5604 34214
rect 5656 34162 6207 34214
rect 5447 34150 6207 34162
rect 5447 34098 5604 34150
rect 5656 34098 6207 34150
rect 5447 34086 6207 34098
rect 5447 34034 5604 34086
rect 5656 34057 6207 34086
rect 7526 34386 7532 34420
rect 7566 34386 7572 34420
rect 7526 34347 7572 34386
rect 7526 34313 7532 34347
rect 7566 34313 7572 34347
rect 7526 34274 7572 34313
rect 7526 34240 7532 34274
rect 7566 34240 7572 34274
rect 7526 34201 7572 34240
rect 7526 34167 7532 34201
rect 7566 34167 7572 34201
rect 7526 34128 7572 34167
rect 7526 34094 7532 34128
rect 7566 34094 7572 34128
tri 6207 34057 6210 34060 sw
rect 5656 34055 6210 34057
tri 6210 34055 6212 34057 sw
rect 7526 34055 7572 34094
rect 5656 34034 6212 34055
rect 5447 34026 6212 34034
tri 6212 34026 6241 34055 sw
rect 5447 34022 6207 34026
rect 5447 33970 5604 34022
rect 5656 33980 6207 34022
rect 7526 34021 7532 34055
rect 7566 34021 7572 34055
rect 7526 33982 7572 34021
rect 5656 33970 6209 33980
rect 5447 33958 6209 33970
rect 5447 33906 5604 33958
rect 5656 33948 6209 33958
tri 6209 33948 6241 33980 nw
rect 7526 33948 7532 33982
rect 7566 33948 7572 33982
rect 5656 33906 6207 33948
tri 6207 33946 6209 33948 nw
rect 5447 33894 6207 33906
rect 5447 33842 5604 33894
rect 5656 33842 6207 33894
rect 5447 33830 6207 33842
rect 5447 33778 5604 33830
rect 5656 33778 6207 33830
rect 5447 33766 6207 33778
rect 5447 33714 5604 33766
rect 5656 33714 6207 33766
rect 5447 33702 6207 33714
rect 5447 33650 5604 33702
rect 5656 33650 6207 33702
rect 5447 33638 6207 33650
rect 5447 33586 5604 33638
rect 5656 33586 6207 33638
rect 7526 33909 7572 33948
rect 7526 33875 7532 33909
rect 7566 33875 7572 33909
rect 7526 33836 7572 33875
rect 7526 33802 7532 33836
rect 7566 33802 7572 33836
rect 7526 33763 7572 33802
rect 7526 33729 7532 33763
rect 7566 33729 7572 33763
rect 7526 33690 7572 33729
rect 7526 33656 7532 33690
rect 7566 33656 7572 33690
rect 7526 33617 7572 33656
rect 5447 33583 6207 33586
tri 6207 33583 6228 33604 sw
rect 7526 33583 7532 33617
rect 7566 33583 7572 33617
rect 5447 33574 6228 33583
rect 5447 33522 5604 33574
rect 5656 33570 6228 33574
tri 6228 33570 6241 33583 sw
rect 5656 33524 6207 33570
rect 7526 33544 7572 33583
rect 5656 33522 6227 33524
rect 5447 33510 6227 33522
tri 6227 33510 6241 33524 nw
rect 7526 33510 7532 33544
rect 7566 33510 7572 33544
rect 5447 33458 5604 33510
rect 5656 33458 6207 33510
tri 6207 33490 6227 33510 nw
rect 5447 33446 6207 33458
rect 5447 33394 5604 33446
rect 5656 33394 6207 33446
rect 5447 33382 6207 33394
rect 5447 33330 5604 33382
rect 5656 33330 6207 33382
rect 5447 33318 6207 33330
rect 5447 33266 5604 33318
rect 5656 33266 6207 33318
rect 5447 33254 6207 33266
rect 5447 33202 5604 33254
rect 5656 33202 6207 33254
rect 5447 33190 6207 33202
rect 5447 33138 5604 33190
rect 5656 33145 6207 33190
rect 7526 33471 7572 33510
rect 7526 33437 7532 33471
rect 7566 33437 7572 33471
rect 7526 33398 7572 33437
rect 7526 33364 7532 33398
rect 7566 33364 7572 33398
rect 7526 33325 7572 33364
rect 7526 33291 7532 33325
rect 7566 33291 7572 33325
rect 7526 33252 7572 33291
rect 7526 33218 7532 33252
rect 7566 33218 7572 33252
rect 7526 33179 7572 33218
tri 6207 33145 6210 33148 sw
rect 7526 33145 7532 33179
rect 7566 33145 7572 33179
rect 5656 33138 6210 33145
rect 5447 33126 6210 33138
rect 5447 33074 5604 33126
rect 5656 33121 6210 33126
tri 6210 33121 6234 33145 sw
rect 5656 33118 6234 33121
tri 6234 33118 6237 33121 sw
rect 5656 33114 6237 33118
tri 6237 33114 6241 33118 sw
rect 5656 33074 6207 33114
rect 5447 33068 6207 33074
rect 7526 33106 7572 33145
rect 7526 33072 7532 33106
rect 7566 33072 7572 33106
rect 5447 33062 6222 33068
rect 5447 33010 5604 33062
rect 5656 33049 6222 33062
tri 6222 33049 6241 33068 nw
rect 5656 33046 6219 33049
tri 6219 33046 6222 33049 nw
rect 5656 33010 6207 33046
tri 6207 33034 6219 33046 nw
rect 5447 32998 6207 33010
rect 5447 32946 5604 32998
rect 5656 32946 6207 32998
rect 5447 32934 6207 32946
rect 5447 32882 5604 32934
rect 5656 32882 6207 32934
rect 5447 32870 6207 32882
rect 5447 32818 5604 32870
rect 5656 32818 6207 32870
rect 5447 32806 6207 32818
rect 5447 32754 5604 32806
rect 5656 32754 6207 32806
rect 5447 32742 6207 32754
rect 5447 32690 5604 32742
rect 5656 32690 6207 32742
rect 7526 33033 7572 33072
rect 7526 32999 7532 33033
rect 7566 32999 7572 33033
rect 7526 32960 7572 32999
rect 7526 32926 7532 32960
rect 7566 32926 7572 32960
rect 7526 32887 7572 32926
rect 7526 32853 7532 32887
rect 7566 32853 7572 32887
rect 7526 32814 7572 32853
rect 7526 32780 7532 32814
rect 7566 32780 7572 32814
rect 7526 32741 7572 32780
rect 7526 32707 7532 32741
rect 7566 32707 7572 32741
rect 7526 32695 7572 32707
rect 7994 34846 8040 34884
rect 7994 34812 8000 34846
rect 8034 34812 8040 34846
rect 7994 34774 8040 34812
rect 7994 34740 8000 34774
rect 8034 34740 8040 34774
rect 7994 34702 8040 34740
rect 7994 34668 8000 34702
rect 8034 34668 8040 34702
rect 7994 34630 8040 34668
rect 7994 34596 8000 34630
rect 8034 34596 8040 34630
rect 7994 34558 8040 34596
rect 7994 34524 8000 34558
rect 8034 34524 8040 34558
rect 7994 34486 8040 34524
rect 7994 34452 8000 34486
rect 8034 34452 8040 34486
rect 7994 34414 8040 34452
rect 7994 34380 8000 34414
rect 8034 34380 8040 34414
rect 7994 34342 8040 34380
rect 7994 34308 8000 34342
rect 8034 34308 8040 34342
rect 7994 34270 8040 34308
rect 7994 34236 8000 34270
rect 8034 34236 8040 34270
rect 7994 34198 8040 34236
rect 7994 34164 8000 34198
rect 8034 34164 8040 34198
rect 7994 34126 8040 34164
rect 7994 34092 8000 34126
rect 8034 34092 8040 34126
rect 7994 34054 8040 34092
rect 7994 34020 8000 34054
rect 8034 34020 8040 34054
rect 7994 33982 8040 34020
rect 7994 33948 8000 33982
rect 8034 33948 8040 33982
rect 7994 33910 8040 33948
rect 7994 33876 8000 33910
rect 8034 33876 8040 33910
rect 7994 33838 8040 33876
rect 7994 33804 8000 33838
rect 8034 33804 8040 33838
rect 7994 33766 8040 33804
rect 7994 33732 8000 33766
rect 8034 33732 8040 33766
rect 7994 33694 8040 33732
rect 7994 33660 8000 33694
rect 8034 33660 8040 33694
rect 7994 33622 8040 33660
rect 7994 33588 8000 33622
rect 8034 33588 8040 33622
rect 7994 33550 8040 33588
rect 7994 33516 8000 33550
rect 8034 33516 8040 33550
rect 7994 33478 8040 33516
rect 7994 33444 8000 33478
rect 8034 33444 8040 33478
rect 7994 33406 8040 33444
rect 7994 33372 8000 33406
rect 8034 33372 8040 33406
rect 7994 33334 8040 33372
rect 7994 33300 8000 33334
rect 8034 33300 8040 33334
rect 7994 33262 8040 33300
rect 7994 33228 8000 33262
rect 8034 33228 8040 33262
rect 7994 33190 8040 33228
rect 7994 33156 8000 33190
rect 8034 33156 8040 33190
rect 7994 33118 8040 33156
rect 7994 33084 8000 33118
rect 8034 33084 8040 33118
rect 7994 33046 8040 33084
rect 7994 33012 8000 33046
rect 8034 33012 8040 33046
rect 7994 32974 8040 33012
rect 7994 32940 8000 32974
rect 8034 32940 8040 32974
rect 7994 32902 8040 32940
rect 7994 32868 8000 32902
rect 8034 32868 8040 32902
rect 7994 32830 8040 32868
rect 7994 32796 8000 32830
rect 8034 32796 8040 32830
rect 7994 32758 8040 32796
rect 7994 32724 8000 32758
rect 8034 32724 8040 32758
rect 5447 32689 6207 32690
tri 6207 32689 6210 32692 sw
rect 5447 32686 6210 32689
tri 6210 32686 6213 32689 sw
rect 7994 32686 8040 32724
rect 5447 32677 6213 32686
rect 5447 32625 5604 32677
rect 5656 32658 6213 32677
tri 6213 32658 6241 32686 sw
rect 5656 32625 6207 32658
rect 5447 32612 6207 32625
rect 7994 32652 8000 32686
rect 8034 32652 8040 32686
rect 7994 32614 8040 32652
rect 5447 32560 5604 32612
rect 5656 32580 6209 32612
tri 6209 32580 6241 32612 nw
rect 7994 32580 8000 32614
rect 8034 32580 8040 32614
rect 5656 32560 6207 32580
tri 6207 32578 6209 32580 nw
rect 5447 32547 6207 32560
rect 5447 32495 5604 32547
rect 5656 32495 6207 32547
rect 5447 32482 6207 32495
rect 5447 32430 5604 32482
rect 5656 32430 6207 32482
rect 5447 32417 6207 32430
rect 5447 32365 5604 32417
rect 5656 32365 6207 32417
rect 5447 32352 6207 32365
rect 5447 32300 5604 32352
rect 5656 32300 6207 32352
rect 5447 32287 6207 32300
rect 5447 32235 5604 32287
rect 5656 32235 6207 32287
rect 7526 32539 7572 32551
rect 7526 32505 7532 32539
rect 7566 32505 7572 32539
rect 7526 32467 7572 32505
rect 7526 32433 7532 32467
rect 7566 32433 7572 32467
rect 7526 32395 7572 32433
rect 7526 32361 7532 32395
rect 7566 32361 7572 32395
rect 7526 32323 7572 32361
rect 7526 32289 7532 32323
rect 7566 32289 7572 32323
rect 7526 32251 7572 32289
rect 5447 32222 6207 32235
rect 5447 32170 5604 32222
rect 5656 32217 6207 32222
tri 6207 32217 6226 32236 sw
rect 7526 32217 7532 32251
rect 7566 32217 7572 32251
rect 5656 32202 6226 32217
tri 6226 32202 6241 32217 sw
rect 5656 32170 6207 32202
rect 5447 32157 6207 32170
rect 5447 32105 5604 32157
rect 5656 32156 6207 32157
rect 7526 32179 7572 32217
rect 5656 32145 6230 32156
tri 6230 32145 6241 32156 nw
rect 7526 32145 7532 32179
rect 7566 32145 7572 32179
rect 5656 32105 6207 32145
tri 6207 32122 6230 32145 nw
rect 5447 32092 6207 32105
rect 5447 32040 5604 32092
rect 5656 32040 6207 32092
rect 5447 32027 6207 32040
rect 5447 31975 5604 32027
rect 5656 31975 6207 32027
rect 5447 31962 6207 31975
rect 5447 31910 5604 31962
rect 5656 31910 6207 31962
rect 5447 31897 6207 31910
rect 5447 31845 5604 31897
rect 5656 31845 6207 31897
rect 5447 31832 6207 31845
rect 5447 31780 5604 31832
rect 5656 31780 6207 31832
rect 7526 32107 7572 32145
rect 7526 32073 7532 32107
rect 7566 32073 7572 32107
rect 7526 32035 7572 32073
rect 7526 32001 7532 32035
rect 7566 32001 7572 32035
rect 7526 31963 7572 32001
rect 7526 31929 7532 31963
rect 7566 31929 7572 31963
rect 7526 31891 7572 31929
rect 7526 31857 7532 31891
rect 7566 31857 7572 31891
rect 7526 31819 7572 31857
rect 7526 31785 7532 31819
rect 7566 31785 7572 31819
rect 5447 31767 6207 31780
rect 5447 31715 5604 31767
rect 5656 31753 6207 31767
tri 6207 31753 6234 31780 sw
rect 7526 31759 7572 31785
rect 7994 32542 8040 32580
rect 7994 32508 8000 32542
rect 8034 32508 8040 32542
rect 7994 32470 8040 32508
rect 7994 32436 8000 32470
rect 8034 32436 8040 32470
rect 7994 32398 8040 32436
rect 7994 32364 8000 32398
rect 8034 32364 8040 32398
rect 7994 32326 8040 32364
rect 7994 32292 8000 32326
rect 8034 32292 8040 32326
rect 7994 32254 8040 32292
rect 7994 32220 8000 32254
rect 8034 32220 8040 32254
rect 7994 32182 8040 32220
rect 7994 32148 8000 32182
rect 8034 32148 8040 32182
rect 7994 32110 8040 32148
rect 7994 32076 8000 32110
rect 8034 32076 8040 32110
rect 7994 32038 8040 32076
rect 7994 32004 8000 32038
rect 8034 32004 8040 32038
rect 7994 31966 8040 32004
rect 7994 31932 8000 31966
rect 8034 31932 8040 31966
rect 7994 31894 8040 31932
rect 7994 31860 8000 31894
rect 8034 31860 8040 31894
rect 7994 31822 8040 31860
rect 7994 31788 8000 31822
rect 8034 31788 8040 31822
tri 7572 31759 7578 31765 sw
rect 7526 31753 7578 31759
rect 5656 31750 6234 31753
tri 6234 31750 6237 31753 sw
rect 5656 31747 6237 31750
tri 6237 31747 6240 31750 sw
rect 5656 31746 6240 31747
tri 6240 31746 6241 31747 sw
rect 5656 31715 6207 31746
rect 5447 31702 6207 31715
rect 5447 31650 5604 31702
rect 5656 31700 6207 31702
rect 5656 31681 6222 31700
tri 6222 31681 6241 31700 nw
rect 7526 31689 7578 31701
rect 5656 31678 6219 31681
tri 6219 31678 6222 31681 nw
rect 5656 31675 6216 31678
tri 6216 31675 6219 31678 nw
rect 5656 31650 6207 31675
tri 6207 31666 6216 31675 nw
rect 5447 31637 6207 31650
rect 5447 31585 5604 31637
rect 5656 31585 6207 31637
rect 5447 31572 6207 31585
rect 5447 31520 5604 31572
rect 5656 31520 6207 31572
rect 5447 31507 6207 31520
rect 5447 31455 5604 31507
rect 5656 31455 6207 31507
rect 5447 31442 6207 31455
rect 5447 31390 5604 31442
rect 5656 31390 6207 31442
rect 5447 31377 6207 31390
rect 5447 31325 5604 31377
rect 5656 31325 6207 31377
rect 5447 31321 6207 31325
rect 7526 31631 7578 31637
rect 7526 31603 7572 31631
tri 7572 31625 7578 31631 nw
rect 7994 31750 8040 31788
rect 8760 35001 8860 35007
rect 8760 34949 8784 35001
rect 8836 34949 8860 35001
rect 8760 34937 8860 34949
rect 8760 34885 8784 34937
rect 8836 34885 8860 34937
rect 7994 31716 8000 31750
rect 8034 31716 8040 31750
rect 7994 31678 8040 31716
rect 7994 31644 8000 31678
rect 8034 31644 8040 31678
rect 7526 31569 7532 31603
rect 7566 31569 7572 31603
rect 7526 31531 7572 31569
rect 7526 31497 7532 31531
rect 7566 31497 7572 31531
rect 7526 31459 7572 31497
rect 7526 31425 7532 31459
rect 7566 31425 7572 31459
rect 7526 31387 7572 31425
rect 7526 31353 7532 31387
rect 7566 31353 7572 31387
tri 6207 31321 6210 31324 sw
rect 5447 31318 6210 31321
tri 6210 31318 6213 31321 sw
rect 5447 31315 6213 31318
tri 6213 31315 6216 31318 sw
rect 7526 31315 7572 31353
rect 5447 31312 6216 31315
rect 5447 31260 5604 31312
rect 5656 31290 6216 31312
tri 6216 31290 6241 31315 sw
rect 5656 31260 6207 31290
rect 5447 31247 6207 31260
rect 5447 31195 5604 31247
rect 5656 31244 6207 31247
rect 7526 31281 7532 31315
rect 7566 31281 7572 31315
rect 5656 31243 6240 31244
tri 6240 31243 6241 31244 nw
rect 7526 31243 7572 31281
rect 5656 31195 6207 31243
tri 6207 31210 6240 31243 nw
rect 5447 31182 6207 31195
rect 5447 31130 5604 31182
rect 5656 31130 6207 31182
rect 5447 31117 6207 31130
rect 5447 31065 5604 31117
rect 5656 31065 6207 31117
rect 5447 31052 6207 31065
rect 5447 31000 5604 31052
rect 5656 31000 6207 31052
rect 5447 30987 6207 31000
rect 5447 30935 5604 30987
rect 5656 30935 6207 30987
rect 5447 30922 6207 30935
rect 5447 30870 5604 30922
rect 5656 30870 6207 30922
rect 5447 30857 6207 30870
rect 7526 31209 7532 31243
rect 7566 31209 7572 31243
rect 7526 31171 7572 31209
rect 7526 31137 7532 31171
rect 7566 31137 7572 31171
rect 7526 31099 7572 31137
rect 7526 31065 7532 31099
rect 7566 31065 7572 31099
rect 7526 31026 7572 31065
rect 7526 30992 7532 31026
rect 7566 30992 7572 31026
rect 7526 30953 7572 30992
rect 7526 30919 7532 30953
rect 7566 30919 7572 30953
rect 7526 30880 7572 30919
rect 5447 30805 5604 30857
rect 5656 30846 6207 30857
tri 6207 30846 6229 30868 sw
rect 7526 30846 7532 30880
rect 7566 30846 7572 30880
rect 5656 30834 6229 30846
tri 6229 30834 6241 30846 sw
rect 5656 30805 6207 30834
rect 5447 30792 6207 30805
rect 5447 30740 5604 30792
rect 5656 30788 6207 30792
rect 7526 30807 7572 30846
rect 5656 30773 6226 30788
tri 6226 30773 6241 30788 nw
rect 7526 30773 7532 30807
rect 7566 30773 7572 30807
rect 5656 30740 6207 30773
tri 6207 30754 6226 30773 nw
rect 5447 30727 6207 30740
rect 5447 30675 5604 30727
rect 5656 30675 6207 30727
rect 5447 30662 6207 30675
rect 5447 30610 5604 30662
rect 5656 30610 6207 30662
rect 5447 30597 6207 30610
rect 5447 30545 5604 30597
rect 5656 30545 6207 30597
rect 5447 30532 6207 30545
rect 5447 30480 5604 30532
rect 5656 30480 6207 30532
rect 5447 30467 6207 30480
rect 5447 30415 5604 30467
rect 5656 30415 6207 30467
rect 5447 30408 6207 30415
rect 7526 30734 7572 30773
rect 7526 30700 7532 30734
rect 7566 30700 7572 30734
rect 7526 30661 7572 30700
rect 7526 30627 7532 30661
rect 7566 30627 7572 30661
rect 7526 30588 7572 30627
rect 7526 30554 7532 30588
rect 7566 30554 7572 30588
rect 7526 30515 7572 30554
rect 7526 30481 7532 30515
rect 7566 30481 7572 30515
rect 7526 30442 7572 30481
tri 6207 30408 6211 30412 sw
rect 7526 30408 7532 30442
rect 7566 30408 7572 30442
rect 5447 30402 6211 30408
rect 5447 30350 5604 30402
rect 5656 30396 6211 30402
tri 6211 30396 6223 30408 sw
rect 7526 30396 7572 30408
rect 7994 31606 8040 31644
rect 7994 31572 8000 31606
rect 8034 31572 8040 31606
rect 7994 31534 8040 31572
rect 7994 31500 8000 31534
rect 8034 31500 8040 31534
rect 7994 31462 8040 31500
rect 7994 31428 8000 31462
rect 8034 31428 8040 31462
rect 7994 31390 8040 31428
rect 7994 31356 8000 31390
rect 8034 31356 8040 31390
rect 7994 31318 8040 31356
rect 7994 31284 8000 31318
rect 8034 31284 8040 31318
rect 7994 31246 8040 31284
rect 7994 31212 8000 31246
rect 8034 31212 8040 31246
rect 7994 31174 8040 31212
rect 7994 31140 8000 31174
rect 8034 31140 8040 31174
rect 7994 31102 8040 31140
rect 7994 31068 8000 31102
rect 8034 31068 8040 31102
rect 7994 31030 8040 31068
rect 7994 30996 8000 31030
rect 8034 30996 8040 31030
rect 7994 30958 8040 30996
rect 7994 30924 8000 30958
rect 8034 30924 8040 30958
rect 7994 30886 8040 30924
rect 7994 30852 8000 30886
rect 8034 30852 8040 30886
rect 7994 30814 8040 30852
rect 7994 30780 8000 30814
rect 8034 30780 8040 30814
rect 7994 30742 8040 30780
rect 7994 30708 8000 30742
rect 8034 30708 8040 30742
rect 7994 30670 8040 30708
rect 7994 30636 8000 30670
rect 8034 30636 8040 30670
rect 7994 30598 8040 30636
rect 7994 30564 8000 30598
rect 8034 30564 8040 30598
rect 7994 30526 8040 30564
rect 7994 30492 8000 30526
rect 8034 30492 8040 30526
rect 7994 30454 8040 30492
rect 7994 30420 8000 30454
rect 8034 30420 8040 30454
rect 5656 30385 6223 30396
tri 6223 30385 6234 30396 sw
rect 5656 30382 6234 30385
tri 6234 30382 6237 30385 sw
rect 7994 30382 8040 30420
rect 5656 30378 6237 30382
tri 6237 30378 6241 30382 sw
rect 5656 30350 6207 30378
rect 5447 30332 6207 30350
rect 7994 30348 8000 30382
rect 8034 30348 8040 30382
rect 7994 30310 8040 30348
rect 7994 30276 8000 30310
rect 8034 30276 8040 30310
rect 7994 30238 8040 30276
rect 7994 30204 8000 30238
rect 8034 30204 8040 30238
rect 7994 30166 8040 30204
rect 7994 30132 8000 30166
rect 8034 30132 8040 30166
rect 7994 30094 8040 30132
rect 6800 30034 7605 30062
tri 7527 30025 7536 30034 ne
rect 7536 30025 7605 30034
tri 7536 30022 7539 30025 ne
rect 7539 30022 7605 30025
tri 7539 30006 7555 30022 ne
rect 7555 30006 7605 30022
rect 6945 29988 7472 30006
tri 7472 29988 7490 30006 sw
tri 7555 29988 7573 30006 ne
rect 7573 29988 7605 30006
rect 6945 29978 7490 29988
tri 7444 29953 7469 29978 ne
rect 7469 29953 7490 29978
tri 7490 29953 7525 29988 sw
tri 7573 29984 7577 29988 ne
tri 7469 29950 7472 29953 ne
rect 7472 29950 7525 29953
rect 7017 29936 7368 29950
tri 7368 29936 7382 29950 sw
tri 7472 29936 7486 29950 ne
rect 7486 29936 7525 29950
rect 7017 29922 7382 29936
tri 7334 29916 7340 29922 ne
rect 7340 29916 7382 29922
tri 7382 29916 7402 29936 sw
tri 7486 29928 7494 29936 ne
rect 7494 29928 7525 29936
tri 7494 29925 7497 29928 ne
tri 7340 29911 7345 29916 ne
rect 7345 29911 7402 29916
tri 7402 29911 7407 29916 sw
rect 5708 29859 5714 29911
rect 5766 29859 5801 29911
rect 5853 29859 5859 29911
tri 7345 29894 7362 29911 ne
rect 7362 29894 7407 29911
rect 5708 29835 5859 29859
rect 5708 29783 5714 29835
rect 5766 29783 5801 29835
rect 5853 29783 5859 29835
rect 6769 29888 7131 29894
rect 6769 29854 6781 29888
rect 6815 29854 6853 29888
rect 6887 29854 7013 29888
rect 7047 29854 7085 29888
rect 7119 29854 7131 29888
tri 7362 29881 7375 29894 ne
rect 7375 29881 7407 29894
tri 7407 29881 7437 29911 sw
tri 7375 29878 7378 29881 ne
rect 7378 29878 7437 29881
tri 7437 29878 7440 29881 sw
tri 7378 29874 7382 29878 ne
rect 7382 29874 7440 29878
tri 7440 29874 7444 29878 sw
rect 6769 29848 7131 29854
rect 6769 29844 6847 29848
tri 6847 29844 6851 29848 nw
tri 6893 29844 6897 29848 ne
rect 6897 29844 7003 29848
tri 7003 29844 7007 29848 nw
tri 7049 29844 7053 29848 ne
rect 7053 29844 7131 29848
tri 7382 29844 7412 29874 ne
rect 7412 29844 7444 29874
rect 5708 29772 5859 29783
tri 5859 29772 5877 29790 sw
rect 5708 29756 5877 29772
tri 5877 29756 5893 29772 sw
rect 5708 29737 5993 29756
tri 5993 29737 6012 29756 sw
rect 5708 29734 6012 29737
tri 6012 29734 6015 29737 sw
rect 5708 29729 6015 29734
tri 6015 29729 6020 29734 sw
rect 5708 29704 6020 29729
tri 6020 29704 6045 29729 sw
rect 5708 29700 5889 29704
tri 5889 29700 5893 29704 nw
tri 5971 29700 5975 29704 ne
rect 5975 29700 6045 29704
tri 6045 29700 6049 29704 sw
rect 5708 29692 5881 29700
tri 5881 29692 5889 29700 nw
tri 5975 29692 5983 29700 ne
rect 5983 29692 6049 29700
tri 6049 29692 6057 29700 sw
rect 5708 29689 5878 29692
tri 5878 29689 5881 29692 nw
tri 5983 29689 5986 29692 ne
rect 5986 29689 6057 29692
tri 6057 29689 6060 29692 sw
rect 5708 29603 5859 29689
tri 5859 29670 5878 29689 nw
tri 5986 29670 6005 29689 ne
rect 6005 29670 6060 29689
tri 6060 29670 6079 29689 sw
tri 6183 29670 6202 29689 se
rect 6202 29670 6250 29694
tri 6005 29665 6010 29670 ne
rect 6010 29665 6079 29670
tri 6079 29665 6084 29670 sw
tri 6178 29665 6183 29670 se
rect 6183 29665 6250 29670
tri 6250 29665 6274 29689 sw
tri 6336 29665 6360 29689 se
rect 6360 29665 6406 29694
tri 6406 29665 6430 29689 sw
tri 6492 29665 6516 29689 se
rect 6516 29665 6564 29694
tri 6564 29665 6588 29689 sw
tri 6745 29665 6769 29689 se
rect 6769 29665 6817 29844
tri 6817 29814 6847 29844 nw
tri 6897 29814 6927 29844 ne
rect 6927 29746 6973 29844
tri 6973 29814 7003 29844 nw
tri 7053 29814 7083 29844 ne
tri 6817 29665 6841 29689 sw
tri 6903 29665 6927 29689 se
rect 6927 29665 6973 29694
tri 6973 29665 6997 29689 sw
tri 7059 29665 7083 29689 se
rect 7083 29665 7131 29844
tri 7412 29840 7416 29844 ne
tri 7383 29700 7416 29733 se
rect 7416 29700 7444 29844
rect 7497 29844 7525 29928
rect 7577 29916 7605 29988
rect 7994 30060 8000 30094
rect 8034 30060 8040 30094
rect 7994 30022 8040 30060
rect 7994 29988 8000 30022
rect 8034 29988 8040 30022
rect 7994 29950 8040 29988
tri 7605 29916 7617 29928 sw
rect 7994 29916 8000 29950
rect 8034 29916 8040 29950
rect 7577 29911 7617 29916
tri 7617 29911 7622 29916 sw
rect 7577 29894 7622 29911
tri 7622 29894 7639 29911 sw
tri 7525 29844 7529 29848 sw
rect 7497 29814 7529 29844
tri 7529 29814 7559 29844 sw
rect 7577 29842 7583 29894
rect 7635 29842 7647 29894
rect 7699 29842 7705 29894
rect 7994 29878 8040 29916
rect 7994 29844 8000 29878
rect 8034 29844 8040 29878
rect 7497 29762 7503 29814
rect 7555 29762 7567 29814
rect 7619 29762 7625 29814
rect 7994 29806 8040 29844
rect 7994 29772 8000 29806
rect 8034 29772 8040 29806
tri 7382 29699 7383 29700 se
rect 7383 29699 7444 29700
tri 6010 29662 6013 29665 ne
rect 6013 29662 6084 29665
tri 6084 29662 6087 29665 sw
tri 6175 29662 6178 29665 se
rect 6178 29662 6274 29665
tri 6274 29662 6277 29665 sw
tri 6333 29662 6336 29665 se
rect 6336 29662 6430 29665
tri 6430 29662 6433 29665 sw
tri 6489 29662 6492 29665 se
rect 6492 29662 6588 29665
tri 6588 29662 6591 29665 sw
tri 6742 29662 6745 29665 se
rect 6745 29662 6841 29665
tri 6841 29662 6844 29665 sw
tri 6900 29662 6903 29665 se
rect 6903 29662 6997 29665
tri 6997 29662 7000 29665 sw
tri 7056 29662 7059 29665 se
rect 7059 29662 7131 29665
tri 6013 29655 6020 29662 ne
rect 6020 29655 6087 29662
tri 6087 29655 6094 29662 sw
tri 6168 29655 6175 29662 se
rect 6175 29655 6277 29662
tri 6277 29655 6284 29662 sw
tri 6326 29655 6333 29662 se
rect 6333 29655 6433 29662
tri 6433 29655 6440 29662 sw
tri 6482 29655 6489 29662 se
rect 6489 29655 6591 29662
tri 6591 29655 6598 29662 sw
tri 6735 29655 6742 29662 se
rect 6742 29655 6844 29662
tri 6844 29655 6851 29662 sw
tri 6893 29655 6900 29662 se
rect 6900 29655 7000 29662
tri 7000 29655 7007 29662 sw
tri 7049 29655 7056 29662 se
rect 7056 29655 7131 29662
tri 6020 29647 6028 29655 ne
rect 6028 29647 7131 29655
rect 7316 29647 7322 29699
rect 7374 29647 7386 29699
rect 7438 29647 7444 29699
rect 7994 29734 8040 29772
rect 7994 29700 8000 29734
rect 8034 29700 8040 29734
rect 7994 29662 8040 29700
tri 6028 29628 6047 29647 ne
rect 6047 29628 7131 29647
tri 6047 29605 6070 29628 ne
rect 6070 29605 7131 29628
tri 5859 29603 5861 29605 sw
tri 6070 29603 6072 29605 ne
rect 6072 29603 7131 29605
rect 7994 29628 8000 29662
rect 8034 29628 8040 29662
rect 5708 29593 5861 29603
tri 5861 29593 5871 29603 sw
rect 5708 29590 5871 29593
tri 5871 29590 5874 29593 sw
rect 7994 29590 8040 29628
rect 5708 29571 5874 29590
tri 5874 29571 5893 29590 sw
rect 5708 29565 7489 29571
rect 5708 29531 5850 29565
rect 5884 29531 5923 29565
rect 5957 29531 5996 29565
rect 6030 29531 6069 29565
rect 6103 29531 6142 29565
rect 6176 29531 6215 29565
rect 6249 29531 6288 29565
rect 6322 29531 6361 29565
rect 6395 29531 6434 29565
rect 6468 29531 6507 29565
rect 6541 29531 6579 29565
rect 6613 29531 6651 29565
rect 6685 29531 6723 29565
rect 6757 29531 6795 29565
rect 6829 29531 6867 29565
rect 6901 29531 6939 29565
rect 6973 29531 7011 29565
rect 7045 29531 7083 29565
rect 7117 29531 7155 29565
rect 7189 29531 7227 29565
rect 7261 29531 7299 29565
rect 7333 29531 7371 29565
rect 7405 29531 7443 29565
rect 7477 29531 7489 29565
rect 5708 29525 7489 29531
rect 5708 29521 5889 29525
tri 5889 29521 5893 29525 nw
tri 7409 29521 7413 29525 ne
rect 7413 29521 7489 29525
rect 5708 29518 5886 29521
tri 5886 29518 5889 29521 nw
tri 7413 29518 7416 29521 ne
rect 7416 29518 7489 29521
rect 5708 29233 5859 29518
tri 5859 29491 5886 29518 nw
tri 7416 29491 7443 29518 ne
rect 7443 29425 7489 29518
rect 7994 29556 8000 29590
rect 8034 29556 8040 29590
rect 7994 29518 8040 29556
rect 7994 29484 8000 29518
rect 8034 29484 8040 29518
rect 7994 29446 8040 29484
rect 7994 29412 8000 29446
rect 8034 29412 8040 29446
rect 7994 29374 8040 29412
rect 7994 29340 8000 29374
rect 8034 29340 8040 29374
rect 7994 29302 8040 29340
rect 7994 29268 8000 29302
rect 8034 29268 8040 29302
tri 5859 29233 5860 29234 sw
rect 5708 29230 5860 29233
tri 5860 29230 5863 29233 sw
rect 7994 29230 8040 29268
rect 5708 29200 5863 29230
tri 5863 29200 5893 29230 sw
rect 5708 29194 6715 29200
rect 5708 29160 5939 29194
rect 5973 29160 6020 29194
rect 6054 29160 6101 29194
rect 6135 29160 6182 29194
rect 6216 29160 6263 29194
rect 6297 29160 6344 29194
rect 6378 29160 6425 29194
rect 6459 29160 6505 29194
rect 6539 29160 6585 29194
rect 6619 29160 6715 29194
rect 5708 29154 6715 29160
rect 5708 29124 5863 29154
tri 5863 29124 5893 29154 nw
tri 6635 29124 6665 29154 ne
rect 6665 29124 6715 29154
rect 5708 28836 5859 29124
tri 5859 29120 5863 29124 nw
tri 6665 29120 6669 29124 ne
rect 6669 29012 6715 29124
rect 6883 29194 7085 29200
rect 6883 29160 6946 29194
rect 6980 29160 7018 29194
rect 7052 29160 7085 29194
rect 6883 29154 7085 29160
rect 6883 29124 6933 29154
tri 6933 29124 6963 29154 nw
tri 7005 29124 7035 29154 ne
rect 7035 29124 7085 29154
rect 6883 29073 6929 29124
tri 6929 29120 6933 29124 nw
tri 7035 29120 7039 29124 ne
rect 7039 29078 7085 29124
rect 7249 29194 7451 29200
rect 7249 29160 7314 29194
rect 7348 29160 7386 29194
rect 7420 29160 7451 29194
rect 7249 29154 7451 29160
rect 7249 29124 7299 29154
tri 7299 29124 7329 29154 nw
tri 7371 29124 7401 29154 ne
rect 7401 29124 7451 29154
rect 7249 29040 7295 29124
tri 7295 29120 7299 29124 nw
tri 7401 29120 7405 29124 ne
rect 7405 29025 7451 29124
rect 7994 29196 8000 29230
rect 8034 29196 8040 29230
rect 7994 29158 8040 29196
rect 7994 29124 8000 29158
rect 8034 29124 8040 29158
rect 7994 29086 8040 29124
rect 7994 29052 8000 29086
rect 8034 29052 8040 29086
rect 7994 29014 8040 29052
rect 7994 28980 8000 29014
rect 8034 28980 8040 29014
rect 7994 28942 8040 28980
rect 7994 28908 8000 28942
rect 8034 28908 8040 28942
rect 6883 28870 6929 28896
tri 6929 28870 6930 28871 sw
tri 7038 28870 7039 28871 se
rect 7039 28870 7085 28896
tri 5859 28836 5885 28862 sw
rect 6883 28837 6930 28870
tri 6930 28837 6963 28870 sw
tri 7005 28837 7038 28870 se
rect 7038 28837 7085 28870
rect 5708 28828 5885 28836
tri 5885 28828 5893 28836 sw
rect 5708 28822 6715 28828
rect 5708 28788 5939 28822
rect 5973 28788 6020 28822
rect 6054 28788 6101 28822
rect 6135 28788 6182 28822
rect 6216 28788 6263 28822
rect 6297 28788 6344 28822
rect 6378 28788 6425 28822
rect 6459 28788 6505 28822
rect 6539 28788 6585 28822
rect 6619 28788 6715 28822
rect 5708 28782 6715 28788
rect 5708 28764 5875 28782
tri 5875 28764 5893 28782 nw
tri 6635 28764 6653 28782 ne
rect 6653 28764 6715 28782
rect 5708 28441 5859 28764
tri 5859 28748 5875 28764 nw
tri 6653 28748 6669 28764 ne
rect 6669 28640 6715 28764
rect 6883 28822 7085 28837
rect 6883 28788 6946 28822
rect 6980 28788 7018 28822
rect 7052 28788 7085 28822
rect 6883 28782 7085 28788
rect 6883 28764 6945 28782
tri 6945 28764 6963 28782 nw
tri 7005 28764 7023 28782 ne
rect 7023 28764 7085 28782
rect 6883 28710 6929 28764
tri 6929 28748 6945 28764 nw
tri 7023 28748 7039 28764 ne
rect 7039 28715 7085 28764
rect 7994 28870 8040 28908
rect 7994 28836 8000 28870
rect 8034 28836 8040 28870
rect 7994 28798 8040 28836
rect 7994 28764 8000 28798
rect 8034 28764 8040 28798
rect 7994 28726 8040 28764
rect 7994 28692 8000 28726
rect 8034 28692 8040 28726
rect 7994 28654 8040 28692
rect 7994 28620 8000 28654
rect 8034 28620 8040 28654
rect 7994 28582 8040 28620
rect 7994 28548 8000 28582
rect 8034 28548 8040 28582
tri 5859 28441 5882 28464 sw
tri 6860 28441 6883 28464 se
rect 6883 28441 6929 28533
rect 7994 28510 8040 28548
tri 6929 28441 6952 28464 sw
tri 7226 28441 7249 28464 se
rect 7249 28441 7295 28496
tri 7295 28441 7318 28464 sw
tri 7382 28441 7405 28464 se
rect 7405 28441 7451 28496
rect 5708 28438 5882 28441
tri 5882 28438 5885 28441 sw
tri 6857 28438 6860 28441 se
rect 6860 28438 6952 28441
tri 6952 28438 6955 28441 sw
tri 7223 28438 7226 28441 se
rect 7226 28438 7318 28441
tri 7318 28438 7321 28441 sw
tri 7379 28438 7382 28441 se
rect 7382 28438 7451 28441
rect 5708 28430 5885 28438
tri 5885 28430 5893 28438 sw
tri 6849 28430 6857 28438 se
rect 6857 28430 6955 28438
tri 6955 28430 6963 28438 sw
tri 7215 28430 7223 28438 se
rect 7223 28430 7321 28438
tri 7321 28430 7329 28438 sw
tri 7371 28430 7379 28438 se
rect 7379 28430 7451 28438
rect 5708 28424 7451 28430
rect 5708 28390 5867 28424
rect 5901 28390 5943 28424
rect 5977 28390 6019 28424
rect 6053 28390 6095 28424
rect 6129 28390 6171 28424
rect 6205 28390 6246 28424
rect 6280 28390 6321 28424
rect 6355 28390 6396 28424
rect 6430 28390 6471 28424
rect 6505 28390 6546 28424
rect 6580 28390 6621 28424
rect 6655 28390 6696 28424
rect 6730 28390 6771 28424
rect 6805 28390 6846 28424
rect 6880 28390 6921 28424
rect 6955 28390 6996 28424
rect 7030 28390 7071 28424
rect 7105 28390 7146 28424
rect 7180 28390 7221 28424
rect 7255 28390 7296 28424
rect 7330 28390 7371 28424
rect 7405 28390 7451 28424
rect 5708 28301 7451 28390
rect 7994 28476 8000 28510
rect 8034 28476 8040 28510
rect 7994 28438 8040 28476
rect 7994 28404 8000 28438
rect 8034 28404 8040 28438
rect 7994 28366 8040 28404
rect 7994 28332 8000 28366
rect 8034 28332 8040 28366
rect 7994 28294 8040 28332
rect 7994 28260 8000 28294
rect 8034 28260 8040 28294
rect 7994 28222 8040 28260
rect 7994 28188 8000 28222
rect 8034 28188 8040 28222
rect 7994 28150 8040 28188
rect 7994 28116 8000 28150
rect 8034 28116 8040 28150
rect 7994 28078 8040 28116
rect 7994 28044 8000 28078
rect 8034 28044 8040 28078
rect 7994 28006 8040 28044
rect 7994 27972 8000 28006
rect 8034 27972 8040 28006
rect 7994 27934 8040 27972
rect 7994 27900 8000 27934
rect 8034 27900 8040 27934
rect 7994 27862 8040 27900
rect 7994 27828 8000 27862
rect 8034 27828 8040 27862
rect 7994 27790 8040 27828
rect 7994 27756 8000 27790
rect 8034 27756 8040 27790
rect 7994 27718 8040 27756
rect 7994 27684 8000 27718
rect 8034 27684 8040 27718
rect 7994 27646 8040 27684
rect 7994 27612 8000 27646
rect 8034 27612 8040 27646
rect 7994 27574 8040 27612
rect 7994 27540 8000 27574
rect 8034 27540 8040 27574
rect 7994 27502 8040 27540
rect 7994 27468 8000 27502
rect 8034 27468 8040 27502
rect 7994 27430 8040 27468
rect 7994 27396 8000 27430
rect 8034 27396 8040 27430
rect 7994 27358 8040 27396
rect 7994 27324 8000 27358
rect 8034 27324 8040 27358
rect 6733 27280 7800 27310
rect 6733 27228 6739 27280
rect 6791 27228 6806 27280
rect 6858 27228 6873 27280
rect 6925 27228 6940 27280
rect 6992 27228 7007 27280
rect 7059 27228 7074 27280
rect 7126 27228 7141 27280
rect 7193 27228 7208 27280
rect 7260 27228 7275 27280
rect 7327 27228 7342 27280
rect 7394 27228 7409 27280
rect 7461 27228 7476 27280
rect 7528 27228 7543 27280
rect 7595 27228 7610 27280
rect 7662 27228 7676 27280
rect 7728 27228 7742 27280
rect 7794 27228 7800 27280
rect 6733 27197 7800 27228
rect 2819 27126 4669 27138
rect 2819 27092 2825 27126
rect 2859 27092 4669 27126
rect 2819 27086 4669 27092
rect 4721 27086 4736 27138
rect 4788 27086 4803 27138
rect 4855 27086 4870 27138
rect 4922 27086 4937 27138
rect 4989 27086 5004 27138
rect 5056 27086 5071 27138
rect 5123 27086 5138 27138
rect 5190 27086 5205 27138
rect 5257 27086 5272 27138
rect 5324 27086 5339 27138
rect 5391 27086 5406 27138
rect 5458 27086 5473 27138
rect 5525 27086 5539 27138
rect 5591 27086 5605 27138
rect 5657 27088 6117 27138
rect 5657 27086 5929 27088
rect 2819 27060 5929 27086
rect 2819 27054 4669 27060
rect 2819 27020 2825 27054
rect 2859 27020 4669 27054
rect 2819 27008 4669 27020
rect 4721 27008 4736 27060
rect 4788 27008 4803 27060
rect 4855 27008 4870 27060
rect 4922 27008 4937 27060
rect 4989 27008 5004 27060
rect 5056 27008 5071 27060
rect 5123 27008 5138 27060
rect 5190 27008 5205 27060
rect 5257 27008 5272 27060
rect 5324 27008 5339 27060
rect 5391 27008 5406 27060
rect 5458 27008 5473 27060
rect 5525 27008 5539 27060
rect 5591 27008 5605 27060
rect 5657 27054 5929 27060
rect 5963 27054 6071 27088
rect 6105 27054 6117 27088
rect 5657 27008 6117 27054
rect 6473 27008 6479 27124
rect 6595 27008 6603 27124
rect 6473 27006 6603 27008
rect 6831 27091 6961 27097
rect 6831 26985 6843 27091
rect 6949 26985 6961 27091
rect 6831 26853 6961 26985
rect 7305 27080 7436 27197
rect 7305 26974 7318 27080
rect 7424 26974 7436 27080
rect 7305 26968 7436 26974
rect 7669 27080 7800 27197
rect 7669 26974 7682 27080
rect 7788 26974 7800 27080
rect 7669 26968 7800 26974
rect 7994 27286 8040 27324
rect 7994 27252 8000 27286
rect 8034 27252 8040 27286
rect 7994 27214 8040 27252
rect 7994 27180 8000 27214
rect 8034 27180 8040 27214
rect 7994 27142 8040 27180
rect 7994 27108 8000 27142
rect 8034 27108 8040 27142
rect 7994 27070 8040 27108
rect 7994 27036 8000 27070
rect 8034 27036 8040 27070
rect 7994 26998 8040 27036
rect 3452 26520 3489 26781
rect 5710 26451 6961 26853
rect 7994 26964 8000 26998
rect 8034 26964 8040 26998
rect 7994 26926 8040 26964
rect 7994 26892 8000 26926
rect 8034 26892 8040 26926
rect 7994 26854 8040 26892
rect 7994 26820 8000 26854
rect 8034 26820 8040 26854
rect 7994 26782 8040 26820
rect 7994 26748 8000 26782
rect 8034 26748 8040 26782
rect 7994 26710 8040 26748
rect 7994 26676 8000 26710
rect 8034 26676 8040 26710
rect 7994 26638 8040 26676
rect 7994 26604 8000 26638
rect 8034 26604 8040 26638
rect 7994 26566 8040 26604
rect 7994 26532 8000 26566
rect 8034 26532 8040 26566
rect 7994 26494 8040 26532
rect 7994 26460 8000 26494
rect 8034 26460 8040 26494
rect 7994 26422 8040 26460
rect 7994 26388 8000 26422
rect 8034 26388 8040 26422
rect 7994 26350 8040 26388
rect 7994 26316 8000 26350
rect 8034 26316 8040 26350
rect 7994 26278 8040 26316
rect 7994 26244 8000 26278
rect 8034 26244 8040 26278
rect 7994 26206 8040 26244
rect 7994 26172 8000 26206
rect 8034 26172 8040 26206
rect 7994 26134 8040 26172
rect 7994 26100 8000 26134
rect 8034 26100 8040 26134
rect 7994 26062 8040 26100
rect 7994 26028 8000 26062
rect 8034 26028 8040 26062
rect 7994 25990 8040 26028
rect 7994 25956 8000 25990
rect 8034 25956 8040 25990
rect 7994 25918 8040 25956
rect 7994 25884 8000 25918
rect 8034 25884 8040 25918
rect 7994 25846 8040 25884
rect 7994 25812 8000 25846
rect 8034 25812 8040 25846
rect 7994 25774 8040 25812
rect 7994 25740 8000 25774
rect 8034 25740 8040 25774
rect 7994 25702 8040 25740
rect 7994 25668 8000 25702
rect 8034 25668 8040 25702
rect 7994 25630 8040 25668
rect 7994 25596 8000 25630
rect 8034 25596 8040 25630
rect 7994 25558 8040 25596
rect 7994 25524 8000 25558
rect 8034 25524 8040 25558
rect 7994 25486 8040 25524
rect 7994 25452 8000 25486
rect 8034 25452 8040 25486
rect 7994 25414 8040 25452
rect 7994 25380 8000 25414
rect 8034 25380 8040 25414
rect 7994 25342 8040 25380
rect 7994 25308 8000 25342
rect 8034 25308 8040 25342
rect 7994 25270 8040 25308
rect 7994 25236 8000 25270
rect 8034 25236 8040 25270
rect 7994 25198 8040 25236
rect 7994 25164 8000 25198
rect 8034 25164 8040 25198
rect 7994 25126 8040 25164
rect 7994 25092 8000 25126
rect 8034 25092 8040 25126
rect 7994 25054 8040 25092
rect 7994 25020 8000 25054
rect 8034 25020 8040 25054
rect 7994 24982 8040 25020
rect 7994 24948 8000 24982
rect 8034 24948 8040 24982
rect 7994 24910 8040 24948
rect 7994 24876 8000 24910
rect 8034 24876 8040 24910
rect 7994 24838 8040 24876
rect 7994 24804 8000 24838
rect 8034 24804 8040 24838
rect 7994 24766 8040 24804
rect 7994 24732 8000 24766
rect 8034 24732 8040 24766
rect 7994 24694 8040 24732
rect 7994 24660 8000 24694
rect 8034 24660 8040 24694
rect 7994 24622 8040 24660
rect 7994 24588 8000 24622
rect 8034 24588 8040 24622
rect 7994 24550 8040 24588
tri 7988 24523 7994 24529 se
rect 7994 24516 8000 24550
rect 8034 24516 8040 24550
rect 7994 24478 8040 24516
rect 7994 24444 8000 24478
rect 8034 24444 8040 24478
rect 7994 24406 8040 24444
rect 7994 24372 8000 24406
rect 8034 24372 8040 24406
rect 7994 24341 8040 24372
tri 7988 24337 7992 24341 ne
rect 7992 24337 8040 24341
tri 7992 24335 7994 24337 ne
rect 7994 24334 8040 24337
rect 7994 24300 8000 24334
rect 8034 24300 8040 24334
rect 7994 24262 8040 24300
rect 7994 24228 8000 24262
rect 8034 24228 8040 24262
rect 7994 24190 8040 24228
rect 7994 24156 8000 24190
rect 8034 24156 8040 24190
rect 7994 24118 8040 24156
rect 7994 24084 8000 24118
rect 8034 24084 8040 24118
rect 7994 24046 8040 24084
rect 7994 24012 8000 24046
rect 8034 24012 8040 24046
rect 7994 23974 8040 24012
rect 7994 23940 8000 23974
rect 8034 23940 8040 23974
rect 7994 23902 8040 23940
rect 7994 23868 8000 23902
rect 8034 23868 8040 23902
rect 7994 23830 8040 23868
rect 7994 23796 8000 23830
rect 8034 23796 8040 23830
rect 7994 23758 8040 23796
rect 7994 23724 8000 23758
rect 8034 23724 8040 23758
rect 7994 23686 8040 23724
rect 7994 23652 8000 23686
rect 8034 23652 8040 23686
rect 7994 23614 8040 23652
rect 7994 23580 8000 23614
rect 8034 23580 8040 23614
rect 7994 23542 8040 23580
rect 7994 23508 8000 23542
rect 8034 23508 8040 23542
rect 7994 23470 8040 23508
rect 7994 23436 8000 23470
rect 8034 23436 8040 23470
rect 7994 23398 8040 23436
rect 7994 23364 8000 23398
rect 8034 23364 8040 23398
rect 7994 23326 8040 23364
tri 7064 23292 7074 23302 se
tri 7040 23268 7064 23292 se
rect 7064 23268 7074 23292
tri 7192 23292 7202 23302 sw
rect 7994 23292 8000 23326
rect 8034 23292 8040 23326
rect 7192 23268 7202 23292
tri 7202 23268 7226 23292 sw
rect 7994 23254 8040 23292
rect 7994 23220 8000 23254
rect 8034 23220 8040 23254
rect 7994 23182 8040 23220
rect 7994 23148 8000 23182
rect 8034 23148 8040 23182
rect 7994 23110 8040 23148
rect 7994 23076 8000 23110
rect 8034 23076 8040 23110
rect 7994 23038 8040 23076
rect 7994 23004 8000 23038
rect 8034 23004 8040 23038
rect 7994 22966 8040 23004
rect 7994 22932 8000 22966
rect 8034 22932 8040 22966
rect 7994 22894 8040 22932
rect 7994 22860 8000 22894
rect 8034 22860 8040 22894
rect 7994 22822 8040 22860
rect 7994 22788 8000 22822
rect 8034 22788 8040 22822
rect 7994 22750 8040 22788
rect 7994 22716 8000 22750
rect 8034 22716 8040 22750
rect 7994 22678 8040 22716
rect 7994 22644 8000 22678
rect 8034 22644 8040 22678
rect 7994 22606 8040 22644
rect 7994 22572 8000 22606
rect 8034 22572 8040 22606
rect 7994 22534 8040 22572
rect 7994 22500 8000 22534
rect 8034 22500 8040 22534
rect 7994 22462 8040 22500
rect 7994 22428 8000 22462
rect 8034 22428 8040 22462
rect 7994 22390 8040 22428
rect 7994 22356 8000 22390
rect 8034 22356 8040 22390
rect 7994 22318 8040 22356
rect 7994 22284 8000 22318
rect 8034 22284 8040 22318
rect 7994 22246 8040 22284
rect 7994 22212 8000 22246
rect 8034 22212 8040 22246
rect 7994 22174 8040 22212
rect 7994 22140 8000 22174
rect 8034 22140 8040 22174
rect 6077 22079 6083 22131
rect 6135 22079 6147 22131
rect 6199 22119 6790 22131
rect 6199 22085 6442 22119
rect 6476 22085 6517 22119
rect 6551 22085 6592 22119
rect 6626 22085 6667 22119
rect 6701 22085 6742 22119
rect 6776 22085 6790 22119
rect 6199 22079 6790 22085
tri 6396 22068 6407 22079 ne
rect 6407 22068 6499 22079
tri 6499 22068 6510 22079 nw
tri 6552 22068 6563 22079 ne
rect 6563 22068 6655 22079
tri 6655 22068 6666 22079 nw
tri 6708 22068 6719 22079 ne
rect 6719 22068 6790 22079
tri 6407 22045 6430 22068 ne
rect 6430 21960 6476 22068
tri 6476 22045 6499 22068 nw
tri 6563 22045 6586 22068 ne
rect 6586 21960 6632 22068
tri 6632 22045 6655 22068 nw
tri 6719 22045 6742 22068 ne
rect 6430 21636 6476 21718
tri 6476 21636 6484 21644 sw
tri 6578 21636 6586 21644 se
rect 6586 21636 6632 21718
tri 6632 21636 6640 21644 sw
tri 6734 21636 6742 21644 se
rect 6742 21636 6790 22068
rect 6430 21610 6484 21636
tri 6484 21610 6510 21636 sw
tri 6552 21610 6578 21636 se
rect 6578 21610 6640 21636
tri 6640 21610 6666 21636 sw
tri 6708 21610 6734 21636 se
rect 6734 21610 6790 21636
rect 6430 21604 6790 21610
rect 6430 21570 6442 21604
rect 6476 21570 6514 21604
rect 6548 21570 6672 21604
rect 6706 21570 6744 21604
rect 6778 21570 6790 21604
rect 6430 21564 6790 21570
rect 7994 22102 8040 22140
rect 7994 22068 8000 22102
rect 8034 22068 8040 22102
rect 7994 22030 8040 22068
rect 7994 21996 8000 22030
rect 8034 21996 8040 22030
rect 7994 21958 8040 21996
rect 7994 21924 8000 21958
rect 8034 21924 8040 21958
rect 7994 21886 8040 21924
rect 7994 21852 8000 21886
rect 8034 21852 8040 21886
rect 7994 21814 8040 21852
rect 7994 21780 8000 21814
rect 8034 21780 8040 21814
rect 7994 21742 8040 21780
rect 7994 21708 8000 21742
rect 8034 21708 8040 21742
rect 7994 21670 8040 21708
rect 7994 21636 8000 21670
rect 8034 21636 8040 21670
rect 7994 21598 8040 21636
rect 7994 21564 8000 21598
rect 8034 21564 8040 21598
rect 7994 21526 8040 21564
rect 7994 21492 8000 21526
rect 8034 21492 8040 21526
rect 7994 21454 8040 21492
rect 6669 21374 6675 21426
rect 6727 21374 6739 21426
rect 6791 21374 6797 21426
rect 7994 21420 8000 21454
rect 8034 21420 8040 21454
rect 7994 21382 8040 21420
rect 7994 21348 8000 21382
rect 8034 21348 8040 21382
rect 6586 21294 6592 21346
rect 6644 21294 6656 21346
rect 6708 21294 6714 21346
rect 7994 21310 8040 21348
rect 7994 21276 8000 21310
rect 8034 21276 8040 21310
rect 6417 21214 6423 21266
rect 6475 21214 6487 21266
rect 6539 21214 6545 21266
rect 7994 21238 8040 21276
rect 7994 21204 8000 21238
rect 8034 21204 8040 21238
rect 7994 21166 8040 21204
rect 7994 21132 8000 21166
rect 8034 21132 8040 21166
rect 7994 21094 8040 21132
rect 7994 21060 8000 21094
rect 8034 21060 8040 21094
rect 7994 21022 8040 21060
rect 7994 20988 8000 21022
rect 8034 20988 8040 21022
rect 7994 20950 8040 20988
rect 7994 20916 8000 20950
rect 8034 20916 8040 20950
rect 7994 20878 8040 20916
rect 7994 20844 8000 20878
rect 8034 20844 8040 20878
rect 7994 20806 8040 20844
rect 7994 20772 8000 20806
rect 8034 20772 8040 20806
rect 7994 20734 8040 20772
rect 7994 20700 8000 20734
rect 8034 20700 8040 20734
rect 7994 20662 8040 20700
rect 7994 20628 8000 20662
rect 8034 20628 8040 20662
rect 7994 20590 8040 20628
rect 7994 20556 8000 20590
rect 8034 20556 8040 20590
rect 7994 20518 8040 20556
rect 7994 20484 8000 20518
rect 8034 20484 8040 20518
rect 7994 20446 8040 20484
rect 7994 20412 8000 20446
rect 8034 20412 8040 20446
rect 7994 20374 8040 20412
rect 7994 20340 8000 20374
rect 8034 20340 8040 20374
rect 7994 20302 8040 20340
rect 7994 20268 8000 20302
rect 8034 20268 8040 20302
rect 7994 20230 8040 20268
rect 7994 20196 8000 20230
rect 8034 20196 8040 20230
rect 7994 20158 8040 20196
rect 7994 20124 8000 20158
rect 8034 20124 8040 20158
rect 7994 20086 8040 20124
rect 7994 20052 8000 20086
rect 8034 20052 8040 20086
rect 7994 20014 8040 20052
rect 7994 19980 8000 20014
rect 8034 19980 8040 20014
rect 7994 19942 8040 19980
rect 7994 19908 8000 19942
rect 8034 19908 8040 19942
rect 7994 19870 8040 19908
rect 7994 19836 8000 19870
rect 8034 19836 8040 19870
rect 7994 19798 8040 19836
rect 7994 19764 8000 19798
rect 8034 19764 8040 19798
rect 7994 19726 8040 19764
rect 7994 19692 8000 19726
rect 8034 19692 8040 19726
rect 7994 19654 8040 19692
rect 7994 19620 8000 19654
rect 8034 19620 8040 19654
rect 7994 19582 8040 19620
rect 7994 19548 8000 19582
rect 8034 19548 8040 19582
rect 7994 19510 8040 19548
rect 7994 19476 8000 19510
rect 8034 19476 8040 19510
rect 7994 19438 8040 19476
rect 7994 19404 8000 19438
rect 8034 19404 8040 19438
rect 7994 19366 8040 19404
rect 7994 19332 8000 19366
rect 8034 19332 8040 19366
rect 7994 19294 8040 19332
rect 7994 19260 8000 19294
rect 8034 19260 8040 19294
rect 7994 19222 8040 19260
rect 7994 19188 8000 19222
rect 8034 19188 8040 19222
rect 7994 19150 8040 19188
rect 7994 19116 8000 19150
rect 8034 19116 8040 19150
rect 7994 19078 8040 19116
rect 7994 19044 8000 19078
rect 8034 19044 8040 19078
rect 7994 19006 8040 19044
rect 7994 18972 8000 19006
rect 8034 18972 8040 19006
rect 7994 18934 8040 18972
rect 7994 18900 8000 18934
rect 8034 18900 8040 18934
rect 7994 18862 8040 18900
rect 7994 18828 8000 18862
rect 8034 18828 8040 18862
rect 7994 18790 8040 18828
rect 7994 18756 8000 18790
rect 8034 18756 8040 18790
rect 7994 18718 8040 18756
rect 7994 18684 8000 18718
rect 8034 18684 8040 18718
rect 7994 18646 8040 18684
rect 7994 18612 8000 18646
rect 8034 18612 8040 18646
rect 7994 18574 8040 18612
rect 7994 18540 8000 18574
rect 8034 18540 8040 18574
rect 7994 18502 8040 18540
rect 7994 18468 8000 18502
rect 8034 18468 8040 18502
rect 7994 18430 8040 18468
rect 7994 18396 8000 18430
rect 8034 18396 8040 18430
rect 7994 18358 8040 18396
rect 7994 18324 8000 18358
rect 8034 18324 8040 18358
rect 7994 18286 8040 18324
rect 7994 18252 8000 18286
rect 8034 18252 8040 18286
rect 7994 18214 8040 18252
rect 7994 18180 8000 18214
rect 8034 18180 8040 18214
rect 7994 18142 8040 18180
rect 7994 18108 8000 18142
rect 8034 18108 8040 18142
rect 7994 18070 8040 18108
rect 7994 18036 8000 18070
rect 8034 18036 8040 18070
rect 7994 17998 8040 18036
rect 7994 17964 8000 17998
rect 8034 17964 8040 17998
rect 7994 17926 8040 17964
rect 7994 17892 8000 17926
rect 8034 17892 8040 17926
rect 7994 17854 8040 17892
rect 7994 17820 8000 17854
rect 8034 17820 8040 17854
rect 7994 17782 8040 17820
rect 7994 17748 8000 17782
rect 8034 17748 8040 17782
rect 7994 17710 8040 17748
rect 7994 17676 8000 17710
rect 8034 17676 8040 17710
rect 7994 17638 8040 17676
rect 7994 17604 8000 17638
rect 8034 17604 8040 17638
rect 7994 17566 8040 17604
rect 7994 17532 8000 17566
rect 8034 17532 8040 17566
rect 7994 17494 8040 17532
rect 7994 17460 8000 17494
rect 8034 17460 8040 17494
rect 7994 17422 8040 17460
rect 7994 17388 8000 17422
rect 8034 17388 8040 17422
rect 7994 17350 8040 17388
rect 7994 17316 8000 17350
rect 8034 17316 8040 17350
rect 7994 17278 8040 17316
rect 7994 17244 8000 17278
rect 8034 17244 8040 17278
rect 7994 17206 8040 17244
rect 7994 17172 8000 17206
rect 8034 17172 8040 17206
rect 7994 17134 8040 17172
rect 7994 17100 8000 17134
rect 8034 17100 8040 17134
rect 7994 17062 8040 17100
rect 7994 17028 8000 17062
rect 8034 17028 8040 17062
rect 7994 16990 8040 17028
rect 7994 16956 8000 16990
rect 8034 16956 8040 16990
rect 7994 16918 8040 16956
rect 7994 16884 8000 16918
rect 8034 16884 8040 16918
rect 7994 16846 8040 16884
rect 7994 16812 8000 16846
rect 8034 16812 8040 16846
rect 7994 16774 8040 16812
rect 7994 16740 8000 16774
rect 8034 16740 8040 16774
rect 7994 16702 8040 16740
rect 7994 16668 8000 16702
rect 8034 16668 8040 16702
rect 7994 16630 8040 16668
rect 7994 16596 8000 16630
rect 8034 16596 8040 16630
rect 7994 16558 8040 16596
rect 7994 16524 8000 16558
rect 8034 16524 8040 16558
rect 7994 16486 8040 16524
rect 7994 16452 8000 16486
rect 8034 16452 8040 16486
rect 7994 16414 8040 16452
rect 7994 16380 8000 16414
rect 8034 16380 8040 16414
rect 7994 16342 8040 16380
rect 7994 16308 8000 16342
rect 8034 16308 8040 16342
rect 7994 16270 8040 16308
rect 7994 16236 8000 16270
rect 8034 16236 8040 16270
rect 7994 16198 8040 16236
rect 7994 16164 8000 16198
rect 8034 16164 8040 16198
rect 7994 16126 8040 16164
rect 7994 16092 8000 16126
rect 8034 16092 8040 16126
rect 7994 16054 8040 16092
rect 7994 16020 8000 16054
rect 8034 16020 8040 16054
rect 7994 15982 8040 16020
rect 7994 15948 8000 15982
rect 8034 15948 8040 15982
rect 7994 15910 8040 15948
rect 7994 15876 8000 15910
rect 8034 15876 8040 15910
rect 7994 15838 8040 15876
rect 7994 15804 8000 15838
rect 8034 15804 8040 15838
rect 7994 15766 8040 15804
rect 7994 15732 8000 15766
rect 8034 15732 8040 15766
rect 7994 15694 8040 15732
rect 7994 15660 8000 15694
rect 8034 15660 8040 15694
rect 7994 15622 8040 15660
rect 7994 15588 8000 15622
rect 8034 15588 8040 15622
rect 7994 15550 8040 15588
rect 7994 15516 8000 15550
rect 8034 15516 8040 15550
rect 7994 15478 8040 15516
rect 7994 15444 8000 15478
rect 8034 15444 8040 15478
rect 7994 15406 8040 15444
rect 7994 15372 8000 15406
rect 8034 15372 8040 15406
rect 7994 15334 8040 15372
rect 7994 15300 8000 15334
rect 8034 15300 8040 15334
rect 7994 15262 8040 15300
rect 7994 15228 8000 15262
rect 8034 15228 8040 15262
rect 7994 15190 8040 15228
rect 7994 15156 8000 15190
rect 8034 15156 8040 15190
rect 7994 15118 8040 15156
rect 7994 15084 8000 15118
rect 8034 15084 8040 15118
rect 7994 15046 8040 15084
rect 7994 15012 8000 15046
rect 8034 15012 8040 15046
rect 7994 14974 8040 15012
rect 7994 14940 8000 14974
rect 8034 14940 8040 14974
rect 7994 14902 8040 14940
rect 7994 14868 8000 14902
rect 8034 14868 8040 14902
rect 7994 14830 8040 14868
rect 7994 14796 8000 14830
rect 8034 14796 8040 14830
rect 7994 14758 8040 14796
rect 7994 14724 8000 14758
rect 8034 14724 8040 14758
rect 7994 14686 8040 14724
rect 7994 14652 8000 14686
rect 8034 14652 8040 14686
rect 7994 14614 8040 14652
rect 7994 14580 8000 14614
rect 8034 14580 8040 14614
rect 7994 14542 8040 14580
rect 7994 14508 8000 14542
rect 8034 14508 8040 14542
rect 7994 14470 8040 14508
rect 7994 14436 8000 14470
rect 8034 14436 8040 14470
rect 7994 14398 8040 14436
rect 7994 14364 8000 14398
rect 8034 14364 8040 14398
rect 7994 14326 8040 14364
rect 7994 14292 8000 14326
rect 8034 14292 8040 14326
rect 7994 14254 8040 14292
rect 7994 14220 8000 14254
rect 8034 14220 8040 14254
rect 7994 14182 8040 14220
rect 7994 14148 8000 14182
rect 8034 14148 8040 14182
rect 7994 14110 8040 14148
rect 7994 14076 8000 14110
rect 8034 14076 8040 14110
rect 7994 14038 8040 14076
rect 7994 14004 8000 14038
rect 8034 14004 8040 14038
rect 7994 13966 8040 14004
rect 7994 13932 8000 13966
rect 8034 13932 8040 13966
rect 7994 13894 8040 13932
rect 7994 13860 8000 13894
rect 8034 13860 8040 13894
rect 7994 13822 8040 13860
rect 7994 13788 8000 13822
rect 8034 13788 8040 13822
rect 7994 13750 8040 13788
rect 7994 13716 8000 13750
rect 8034 13716 8040 13750
rect 7994 13678 8040 13716
rect 7994 13644 8000 13678
rect 8034 13644 8040 13678
rect 7994 13606 8040 13644
rect 7994 13572 8000 13606
rect 8034 13572 8040 13606
rect 7994 13534 8040 13572
rect 7994 13500 8000 13534
rect 8034 13500 8040 13534
rect 7994 13462 8040 13500
rect 7994 13428 8000 13462
rect 8034 13428 8040 13462
rect 7994 13390 8040 13428
rect 7994 13356 8000 13390
rect 8034 13356 8040 13390
rect 7994 13318 8040 13356
rect 7994 13284 8000 13318
rect 8034 13284 8040 13318
rect 7994 13246 8040 13284
rect 7994 13212 8000 13246
rect 8034 13212 8040 13246
rect 7994 13174 8040 13212
rect 7994 13140 8000 13174
rect 8034 13140 8040 13174
rect 7994 13102 8040 13140
rect 7994 13068 8000 13102
rect 8034 13068 8040 13102
rect 7994 13030 8040 13068
rect 7994 12996 8000 13030
rect 8034 12996 8040 13030
rect 7994 12958 8040 12996
rect 7994 12924 8000 12958
rect 8034 12924 8040 12958
rect 7994 12886 8040 12924
rect 7994 12852 8000 12886
rect 8034 12852 8040 12886
rect 7994 12814 8040 12852
rect 7994 12780 8000 12814
rect 8034 12780 8040 12814
rect 7994 12742 8040 12780
rect 7994 12708 8000 12742
rect 8034 12708 8040 12742
rect 7994 12670 8040 12708
rect 7994 12636 8000 12670
rect 8034 12636 8040 12670
rect 7994 12598 8040 12636
rect 7994 12564 8000 12598
rect 8034 12564 8040 12598
rect 7994 12526 8040 12564
rect 7994 12492 8000 12526
rect 8034 12492 8040 12526
rect 7994 12454 8040 12492
rect 7994 12420 8000 12454
rect 8034 12420 8040 12454
rect 7994 12382 8040 12420
rect 7994 12348 8000 12382
rect 8034 12348 8040 12382
rect 7994 12310 8040 12348
rect 7994 12276 8000 12310
rect 8034 12276 8040 12310
rect 7994 12238 8040 12276
rect 7994 12204 8000 12238
rect 8034 12204 8040 12238
rect 7994 12166 8040 12204
rect 7994 12132 8000 12166
rect 8034 12132 8040 12166
rect 7994 12094 8040 12132
rect 7994 12060 8000 12094
rect 8034 12060 8040 12094
rect 7994 12022 8040 12060
rect 7994 11988 8000 12022
rect 8034 11988 8040 12022
rect 7994 11950 8040 11988
rect 7994 11916 8000 11950
rect 8034 11916 8040 11950
rect 7994 11878 8040 11916
rect 7994 11844 8000 11878
rect 8034 11844 8040 11878
rect 7994 11806 8040 11844
rect 7994 11772 8000 11806
rect 8034 11772 8040 11806
rect 7994 11734 8040 11772
rect 7994 11700 8000 11734
rect 8034 11700 8040 11734
rect 7994 11662 8040 11700
rect 7994 11628 8000 11662
rect 8034 11628 8040 11662
rect 7994 11590 8040 11628
rect 7994 11556 8000 11590
rect 8034 11556 8040 11590
rect 7994 11518 8040 11556
rect 8068 31753 8120 31759
rect 8068 31689 8120 31701
rect 8068 11537 8120 31637
rect 8760 27130 8860 34885
rect 9746 34993 9792 35031
rect 9746 34959 9752 34993
rect 9786 34959 9792 34993
rect 9746 34921 9792 34959
rect 9746 34887 9752 34921
rect 9786 34887 9792 34921
rect 9746 34849 9792 34887
rect 9746 34815 9752 34849
rect 9786 34815 9792 34849
rect 9746 34777 9792 34815
rect 9746 34743 9752 34777
rect 9786 34743 9792 34777
rect 9746 34705 9792 34743
rect 9746 34671 9752 34705
rect 9786 34671 9792 34705
rect 9746 34633 9792 34671
rect 9746 34599 9752 34633
rect 9786 34599 9792 34633
rect 9746 34561 9792 34599
rect 9746 34527 9752 34561
rect 9786 34527 9792 34561
rect 9746 34489 9792 34527
rect 9746 34455 9752 34489
rect 9786 34455 9792 34489
rect 9746 34417 9792 34455
rect 9746 34383 9752 34417
rect 9786 34383 9792 34417
rect 9746 34345 9792 34383
rect 9746 34311 9752 34345
rect 9786 34311 9792 34345
rect 9746 34273 9792 34311
rect 9746 34239 9752 34273
rect 9786 34239 9792 34273
rect 9746 34201 9792 34239
rect 9746 34167 9752 34201
rect 9786 34167 9792 34201
rect 9746 34129 9792 34167
rect 9746 34095 9752 34129
rect 9786 34095 9792 34129
rect 9746 34057 9792 34095
rect 9746 34023 9752 34057
rect 9786 34023 9792 34057
rect 9746 33985 9792 34023
rect 9746 33951 9752 33985
rect 9786 33951 9792 33985
rect 9746 33913 9792 33951
rect 9746 33879 9752 33913
rect 9786 33879 9792 33913
rect 9746 33841 9792 33879
rect 9746 33807 9752 33841
rect 9786 33807 9792 33841
rect 9746 33769 9792 33807
rect 9746 33735 9752 33769
rect 9786 33735 9792 33769
rect 9746 33697 9792 33735
rect 9746 33663 9752 33697
rect 9786 33663 9792 33697
rect 9746 33625 9792 33663
rect 9746 33591 9752 33625
rect 9786 33591 9792 33625
rect 9746 33553 9792 33591
rect 9746 33519 9752 33553
rect 9786 33519 9792 33553
rect 9746 33481 9792 33519
rect 9746 33447 9752 33481
rect 9786 33447 9792 33481
rect 9746 33409 9792 33447
rect 9746 33375 9752 33409
rect 9786 33375 9792 33409
rect 9746 33337 9792 33375
rect 9746 33303 9752 33337
rect 9786 33303 9792 33337
rect 9746 33265 9792 33303
rect 9746 33231 9752 33265
rect 9786 33231 9792 33265
rect 9746 33193 9792 33231
rect 9746 33159 9752 33193
rect 9786 33159 9792 33193
rect 9746 33121 9792 33159
rect 9746 33087 9752 33121
rect 9786 33087 9792 33121
rect 9746 33049 9792 33087
rect 9746 33015 9752 33049
rect 9786 33015 9792 33049
rect 9746 32977 9792 33015
rect 9746 32943 9752 32977
rect 9786 32943 9792 32977
rect 9746 32905 9792 32943
rect 9746 32871 9752 32905
rect 9786 32871 9792 32905
rect 9746 32833 9792 32871
rect 9746 32799 9752 32833
rect 9786 32799 9792 32833
rect 9746 32761 9792 32799
rect 9746 32727 9752 32761
rect 9786 32727 9792 32761
rect 9746 32689 9792 32727
rect 9746 32655 9752 32689
rect 9786 32655 9792 32689
rect 9746 32617 9792 32655
rect 9746 32583 9752 32617
rect 9786 32583 9792 32617
rect 9746 32545 9792 32583
rect 9746 32511 9752 32545
rect 9786 32511 9792 32545
rect 9746 32473 9792 32511
rect 9746 32439 9752 32473
rect 9786 32439 9792 32473
rect 9746 32401 9792 32439
rect 9746 32367 9752 32401
rect 9786 32367 9792 32401
rect 9746 32329 9792 32367
rect 9746 32295 9752 32329
rect 9786 32295 9792 32329
rect 9746 32257 9792 32295
rect 9746 32223 9752 32257
rect 9786 32223 9792 32257
rect 9746 32185 9792 32223
rect 9746 32151 9752 32185
rect 9786 32151 9792 32185
rect 9746 32113 9792 32151
rect 9746 32079 9752 32113
rect 9786 32079 9792 32113
rect 9746 32041 9792 32079
rect 9746 32007 9752 32041
rect 9786 32007 9792 32041
rect 9746 31969 9792 32007
rect 9746 31935 9752 31969
rect 9786 31935 9792 31969
rect 9746 31897 9792 31935
rect 9746 31863 9752 31897
rect 9786 31863 9792 31897
rect 9746 31825 9792 31863
rect 9746 31791 9752 31825
rect 9786 31791 9792 31825
rect 9746 31753 9792 31791
rect 9746 31719 9752 31753
rect 9786 31719 9792 31753
rect 9746 31681 9792 31719
rect 9746 31647 9752 31681
rect 9786 31647 9792 31681
rect 9746 31609 9792 31647
rect 9746 31575 9752 31609
rect 9786 31575 9792 31609
rect 9746 31537 9792 31575
rect 9746 31503 9752 31537
rect 9786 31503 9792 31537
rect 9746 31465 9792 31503
rect 9746 31431 9752 31465
rect 9786 31431 9792 31465
rect 9746 31393 9792 31431
rect 9746 31359 9752 31393
rect 9786 31359 9792 31393
rect 9746 31321 9792 31359
rect 9746 31287 9752 31321
rect 9786 31287 9792 31321
rect 9746 31249 9792 31287
rect 9746 31215 9752 31249
rect 9786 31215 9792 31249
rect 9746 31177 9792 31215
rect 9746 31143 9752 31177
rect 9786 31143 9792 31177
rect 9746 31105 9792 31143
rect 9746 31071 9752 31105
rect 9786 31071 9792 31105
rect 9746 31033 9792 31071
rect 9746 30999 9752 31033
rect 9786 30999 9792 31033
rect 9746 30961 9792 30999
rect 9746 30927 9752 30961
rect 9786 30927 9792 30961
rect 9746 30889 9792 30927
rect 9746 30855 9752 30889
rect 9786 30855 9792 30889
rect 9746 30817 9792 30855
rect 9746 30783 9752 30817
rect 9786 30783 9792 30817
rect 9746 30745 9792 30783
rect 9746 30711 9752 30745
rect 9786 30711 9792 30745
rect 9746 30673 9792 30711
rect 9746 30639 9752 30673
rect 9786 30639 9792 30673
rect 9746 30601 9792 30639
rect 9746 30567 9752 30601
rect 9786 30567 9792 30601
rect 9746 30529 9792 30567
rect 9746 30495 9752 30529
rect 9786 30495 9792 30529
rect 9746 30457 9792 30495
rect 9746 30423 9752 30457
rect 9786 30423 9792 30457
rect 9746 30385 9792 30423
rect 9746 30351 9752 30385
rect 9786 30351 9792 30385
rect 9746 30313 9792 30351
rect 9746 30279 9752 30313
rect 9786 30279 9792 30313
rect 9746 30241 9792 30279
rect 9746 30207 9752 30241
rect 9786 30207 9792 30241
rect 9746 30169 9792 30207
rect 9746 30135 9752 30169
rect 9786 30135 9792 30169
rect 9746 30097 9792 30135
rect 9746 30063 9752 30097
rect 9786 30063 9792 30097
rect 9746 30025 9792 30063
rect 9746 29991 9752 30025
rect 9786 29991 9792 30025
rect 9746 29953 9792 29991
rect 9746 29919 9752 29953
rect 9786 29919 9792 29953
rect 9088 29842 9094 29894
rect 9146 29842 9158 29894
rect 9210 29842 9216 29894
rect 9746 29881 9792 29919
rect 9746 29847 9752 29881
rect 9786 29847 9792 29881
rect 9008 29808 9060 29814
rect 9008 29744 9060 29756
rect 8760 27078 8784 27130
rect 8836 27078 8860 27130
rect 8760 27066 8860 27078
rect 8760 27014 8784 27066
rect 8836 27014 8860 27066
rect 8760 26358 8860 27014
rect 8760 26306 8784 26358
rect 8836 26306 8860 26358
rect 8760 26294 8860 26306
rect 8760 26242 8784 26294
rect 8836 26242 8860 26294
rect 8760 26236 8860 26242
rect 8928 29693 8980 29699
rect 8928 29629 8980 29641
tri 8925 21457 8928 21460 se
rect 8928 21457 8980 29577
tri 8894 21426 8925 21457 se
rect 8803 21374 8809 21426
rect 8861 21374 8873 21426
rect 8925 21374 8980 21457
rect 9008 21416 9060 29692
rect 9008 21352 9060 21364
rect 9008 21294 9060 21300
rect 9088 29809 9141 29842
tri 9141 29809 9174 29842 nw
rect 9746 29809 9792 29847
rect 9088 21279 9140 29809
tri 9140 29808 9141 29809 nw
rect 9746 29775 9752 29809
rect 9786 29775 9792 29809
rect 9746 29737 9792 29775
rect 9746 29703 9752 29737
rect 9786 29703 9792 29737
rect 9746 29665 9792 29703
rect 9746 29631 9752 29665
rect 9786 29631 9792 29665
rect 9746 29593 9792 29631
rect 9746 29559 9752 29593
rect 9786 29559 9792 29593
rect 9746 29521 9792 29559
rect 9746 29487 9752 29521
rect 9786 29487 9792 29521
rect 9746 29449 9792 29487
rect 9746 29415 9752 29449
rect 9786 29415 9792 29449
rect 9746 29377 9792 29415
rect 9746 29343 9752 29377
rect 9786 29343 9792 29377
rect 9746 29305 9792 29343
rect 9746 29271 9752 29305
rect 9786 29271 9792 29305
rect 9746 29233 9792 29271
rect 9746 29199 9752 29233
rect 9786 29199 9792 29233
rect 9746 29161 9792 29199
rect 9746 29127 9752 29161
rect 9786 29127 9792 29161
rect 9746 29089 9792 29127
rect 9746 29055 9752 29089
rect 9786 29055 9792 29089
rect 9746 29017 9792 29055
rect 9746 28983 9752 29017
rect 9786 28983 9792 29017
rect 9746 28945 9792 28983
rect 9746 28911 9752 28945
rect 9786 28911 9792 28945
rect 9746 28873 9792 28911
rect 9746 28839 9752 28873
rect 9786 28839 9792 28873
rect 9746 28801 9792 28839
rect 9746 28767 9752 28801
rect 9786 28767 9792 28801
rect 9746 28729 9792 28767
rect 9746 28695 9752 28729
rect 9786 28695 9792 28729
rect 9746 28657 9792 28695
rect 9746 28623 9752 28657
rect 9786 28623 9792 28657
rect 9746 28585 9792 28623
rect 9746 28551 9752 28585
rect 9786 28551 9792 28585
rect 9746 28513 9792 28551
rect 9746 28479 9752 28513
rect 9786 28479 9792 28513
rect 9746 28441 9792 28479
rect 9746 28407 9752 28441
rect 9786 28407 9792 28441
rect 9746 28369 9792 28407
rect 9746 28335 9752 28369
rect 9786 28335 9792 28369
rect 9746 28297 9792 28335
rect 9746 28263 9752 28297
rect 9786 28263 9792 28297
rect 9746 28225 9792 28263
rect 9746 28191 9752 28225
rect 9786 28191 9792 28225
rect 9746 28153 9792 28191
rect 9746 28119 9752 28153
rect 9786 28119 9792 28153
rect 9746 28081 9792 28119
rect 9746 28047 9752 28081
rect 9786 28047 9792 28081
rect 9746 28009 9792 28047
rect 9746 27975 9752 28009
rect 9786 27975 9792 28009
rect 9746 27937 9792 27975
rect 9746 27903 9752 27937
rect 9786 27903 9792 27937
rect 9746 27865 9792 27903
rect 9746 27831 9752 27865
rect 9786 27831 9792 27865
rect 9746 27793 9792 27831
rect 9746 27759 9752 27793
rect 9786 27759 9792 27793
rect 9746 27721 9792 27759
rect 9746 27687 9752 27721
rect 9786 27687 9792 27721
rect 9746 27649 9792 27687
rect 9746 27615 9752 27649
rect 9786 27615 9792 27649
rect 9746 27577 9792 27615
rect 9746 27543 9752 27577
rect 9786 27543 9792 27577
rect 9746 27505 9792 27543
rect 9746 27471 9752 27505
rect 9786 27471 9792 27505
rect 9746 27433 9792 27471
rect 9746 27399 9752 27433
rect 9786 27399 9792 27433
rect 9746 27361 9792 27399
rect 9746 27327 9752 27361
rect 9786 27327 9792 27361
rect 9746 27289 9792 27327
rect 9746 27255 9752 27289
rect 9786 27255 9792 27289
rect 9746 27217 9792 27255
rect 9746 27183 9752 27217
rect 9786 27183 9792 27217
rect 9746 27145 9792 27183
rect 9746 27111 9752 27145
rect 9786 27111 9792 27145
rect 9746 27073 9792 27111
rect 9746 27039 9752 27073
rect 9786 27039 9792 27073
rect 9746 27001 9792 27039
rect 9746 26967 9752 27001
rect 9786 26967 9792 27001
rect 9746 26929 9792 26967
rect 9746 26895 9752 26929
rect 9786 26895 9792 26929
rect 9746 26857 9792 26895
rect 9746 26823 9752 26857
rect 9786 26823 9792 26857
rect 9746 26785 9792 26823
rect 9746 26751 9752 26785
rect 9786 26751 9792 26785
rect 9746 26713 9792 26751
rect 9746 26679 9752 26713
rect 9786 26679 9792 26713
rect 9746 26641 9792 26679
rect 9746 26607 9752 26641
rect 9786 26607 9792 26641
rect 9746 26569 9792 26607
rect 9746 26535 9752 26569
rect 9786 26535 9792 26569
rect 9746 26497 9792 26535
rect 9746 26463 9752 26497
rect 9786 26463 9792 26497
rect 9746 26425 9792 26463
rect 9746 26391 9752 26425
rect 9786 26391 9792 26425
rect 9746 26353 9792 26391
rect 9746 26319 9752 26353
rect 9786 26319 9792 26353
rect 9746 26281 9792 26319
rect 9746 26247 9752 26281
rect 9786 26247 9792 26281
rect 9746 26209 9792 26247
rect 9746 26175 9752 26209
rect 9786 26175 9792 26209
rect 9746 26137 9792 26175
rect 9746 26103 9752 26137
rect 9786 26103 9792 26137
rect 9746 26065 9792 26103
rect 9746 26031 9752 26065
rect 9786 26031 9792 26065
rect 9746 25993 9792 26031
rect 9746 25959 9752 25993
rect 9786 25959 9792 25993
rect 9746 25921 9792 25959
rect 9746 25887 9752 25921
rect 9786 25887 9792 25921
rect 9746 25849 9792 25887
rect 9746 25815 9752 25849
rect 9786 25815 9792 25849
rect 9746 25777 9792 25815
rect 9746 25743 9752 25777
rect 9786 25743 9792 25777
rect 9746 25705 9792 25743
rect 9746 25671 9752 25705
rect 9786 25671 9792 25705
rect 9746 25633 9792 25671
rect 9746 25599 9752 25633
rect 9786 25599 9792 25633
rect 9746 25561 9792 25599
rect 9746 25527 9752 25561
rect 9786 25527 9792 25561
rect 9746 25489 9792 25527
rect 9746 25455 9752 25489
rect 9786 25455 9792 25489
rect 9746 25417 9792 25455
rect 9746 25383 9752 25417
rect 9786 25383 9792 25417
rect 9746 25345 9792 25383
rect 9746 25311 9752 25345
rect 9786 25311 9792 25345
rect 9746 25273 9792 25311
rect 9746 25239 9752 25273
rect 9786 25239 9792 25273
rect 9746 25201 9792 25239
rect 9746 25167 9752 25201
rect 9786 25167 9792 25201
rect 9746 25129 9792 25167
rect 9746 25095 9752 25129
rect 9786 25095 9792 25129
rect 9746 25057 9792 25095
rect 9746 25023 9752 25057
rect 9786 25023 9792 25057
rect 9746 24985 9792 25023
rect 9746 24951 9752 24985
rect 9786 24951 9792 24985
rect 9746 24913 9792 24951
rect 9746 24879 9752 24913
rect 9786 24879 9792 24913
rect 9746 24841 9792 24879
rect 9746 24807 9752 24841
rect 9786 24807 9792 24841
rect 9746 24769 9792 24807
rect 9746 24735 9752 24769
rect 9786 24735 9792 24769
rect 9746 24697 9792 24735
rect 9746 24663 9752 24697
rect 9786 24663 9792 24697
rect 9746 24625 9792 24663
rect 9746 24591 9752 24625
rect 9786 24591 9792 24625
rect 9746 24553 9792 24591
rect 9746 24519 9752 24553
rect 9786 24519 9792 24553
rect 9746 24481 9792 24519
rect 9746 24447 9752 24481
rect 9786 24447 9792 24481
rect 9746 24409 9792 24447
rect 9746 24375 9752 24409
rect 9786 24375 9792 24409
rect 9746 24337 9792 24375
rect 9746 24303 9752 24337
rect 9786 24303 9792 24337
rect 9746 24265 9792 24303
rect 9746 24231 9752 24265
rect 9786 24231 9792 24265
rect 9746 24193 9792 24231
rect 9746 24159 9752 24193
rect 9786 24159 9792 24193
rect 9746 24121 9792 24159
rect 9746 24087 9752 24121
rect 9786 24087 9792 24121
rect 9746 24049 9792 24087
rect 9746 24015 9752 24049
rect 9786 24015 9792 24049
rect 9746 23977 9792 24015
rect 9746 23943 9752 23977
rect 9786 23943 9792 23977
rect 9746 23905 9792 23943
rect 9746 23871 9752 23905
rect 9786 23871 9792 23905
rect 9746 23833 9792 23871
rect 9746 23799 9752 23833
rect 9786 23799 9792 23833
rect 9746 23761 9792 23799
rect 9746 23727 9752 23761
rect 9786 23727 9792 23761
rect 9746 23689 9792 23727
rect 9746 23655 9752 23689
rect 9786 23655 9792 23689
rect 9746 23617 9792 23655
rect 9746 23583 9752 23617
rect 9786 23583 9792 23617
rect 9746 23545 9792 23583
rect 9746 23511 9752 23545
rect 9786 23511 9792 23545
rect 9746 23473 9792 23511
rect 9746 23439 9752 23473
rect 9786 23439 9792 23473
rect 9746 23401 9792 23439
rect 9746 23367 9752 23401
rect 9786 23367 9792 23401
rect 9746 23329 9792 23367
rect 9746 23295 9752 23329
rect 9786 23295 9792 23329
rect 9746 23257 9792 23295
rect 9746 23223 9752 23257
rect 9786 23223 9792 23257
rect 9746 23185 9792 23223
rect 9746 23151 9752 23185
rect 9786 23151 9792 23185
rect 9746 23113 9792 23151
rect 9746 23079 9752 23113
rect 9786 23079 9792 23113
rect 9746 23041 9792 23079
rect 9746 23007 9752 23041
rect 9786 23007 9792 23041
rect 9746 22969 9792 23007
rect 9746 22935 9752 22969
rect 9786 22935 9792 22969
rect 9746 22897 9792 22935
rect 9746 22863 9752 22897
rect 9786 22863 9792 22897
rect 9746 22825 9792 22863
rect 9746 22791 9752 22825
rect 9786 22791 9792 22825
rect 9746 22753 9792 22791
rect 9746 22719 9752 22753
rect 9786 22719 9792 22753
rect 9746 22681 9792 22719
rect 9746 22647 9752 22681
rect 9786 22647 9792 22681
rect 9746 22609 9792 22647
rect 9746 22575 9752 22609
rect 9786 22575 9792 22609
rect 9746 22537 9792 22575
rect 9746 22503 9752 22537
rect 9786 22503 9792 22537
rect 9746 22465 9792 22503
rect 9746 22431 9752 22465
rect 9786 22431 9792 22465
rect 9746 22393 9792 22431
rect 9746 22359 9752 22393
rect 9786 22359 9792 22393
rect 9746 22321 9792 22359
rect 9746 22287 9752 22321
rect 9786 22287 9792 22321
rect 9746 22249 9792 22287
rect 9746 22215 9752 22249
rect 9786 22215 9792 22249
rect 9746 22177 9792 22215
rect 9746 22143 9752 22177
rect 9786 22143 9792 22177
rect 9746 22105 9792 22143
rect 9746 22071 9752 22105
rect 9786 22071 9792 22105
rect 9746 22033 9792 22071
rect 9746 21999 9752 22033
rect 9786 21999 9792 22033
rect 9746 21961 9792 21999
rect 9746 21927 9752 21961
rect 9786 21927 9792 21961
rect 9746 21889 9792 21927
rect 9746 21855 9752 21889
rect 9786 21855 9792 21889
rect 9746 21817 9792 21855
rect 9746 21783 9752 21817
rect 9786 21783 9792 21817
rect 9746 21745 9792 21783
rect 9746 21711 9752 21745
rect 9786 21711 9792 21745
rect 9746 21673 9792 21711
rect 9746 21639 9752 21673
rect 9786 21639 9792 21673
rect 9746 21601 9792 21639
rect 9746 21567 9752 21601
rect 9786 21567 9792 21601
rect 9746 21529 9792 21567
rect 9746 21495 9752 21529
rect 9786 21495 9792 21529
rect 9746 21457 9792 21495
rect 9746 21423 9752 21457
rect 9786 21423 9792 21457
rect 9746 21385 9792 21423
rect 9746 21351 9752 21385
rect 9786 21351 9792 21385
rect 9746 21313 9792 21351
tri 9140 21279 9161 21300 sw
rect 9746 21279 9752 21313
rect 9786 21279 9792 21313
rect 9088 21266 9161 21279
tri 9161 21266 9174 21279 sw
rect 9088 21214 9094 21266
rect 9146 21214 9158 21266
rect 9210 21214 9216 21266
rect 9746 21241 9792 21279
rect 9746 21207 9752 21241
rect 9786 21207 9792 21241
rect 9746 21169 9792 21207
rect 9746 21135 9752 21169
rect 9786 21135 9792 21169
rect 9746 21097 9792 21135
rect 9746 21063 9752 21097
rect 9786 21063 9792 21097
rect 9746 21025 9792 21063
rect 9746 20991 9752 21025
rect 9786 20991 9792 21025
rect 9746 20953 9792 20991
rect 9746 20919 9752 20953
rect 9786 20919 9792 20953
rect 9746 20881 9792 20919
rect 9746 20847 9752 20881
rect 9786 20847 9792 20881
rect 9746 20809 9792 20847
rect 9746 20775 9752 20809
rect 9786 20775 9792 20809
rect 9746 20737 9792 20775
rect 9746 20703 9752 20737
rect 9786 20703 9792 20737
rect 9746 20665 9792 20703
rect 9746 20631 9752 20665
rect 9786 20631 9792 20665
rect 9746 20593 9792 20631
rect 9746 20559 9752 20593
rect 9786 20559 9792 20593
rect 9746 20521 9792 20559
rect 9746 20487 9752 20521
rect 9786 20487 9792 20521
rect 9746 20449 9792 20487
rect 9746 20415 9752 20449
rect 9786 20415 9792 20449
rect 9746 20377 9792 20415
rect 9746 20343 9752 20377
rect 9786 20343 9792 20377
rect 9746 20305 9792 20343
rect 9746 20271 9752 20305
rect 9786 20271 9792 20305
rect 9746 20233 9792 20271
rect 9746 20199 9752 20233
rect 9786 20199 9792 20233
rect 9746 20161 9792 20199
rect 9746 20127 9752 20161
rect 9786 20127 9792 20161
rect 9746 20089 9792 20127
rect 9746 20055 9752 20089
rect 9786 20055 9792 20089
rect 9746 20017 9792 20055
rect 9746 19983 9752 20017
rect 9786 19983 9792 20017
rect 9746 19945 9792 19983
rect 9746 19911 9752 19945
rect 9786 19911 9792 19945
rect 9746 19873 9792 19911
rect 9746 19839 9752 19873
rect 9786 19839 9792 19873
rect 9746 19801 9792 19839
rect 9746 19767 9752 19801
rect 9786 19767 9792 19801
rect 9746 19729 9792 19767
rect 9746 19695 9752 19729
rect 9786 19695 9792 19729
rect 9746 19657 9792 19695
rect 9746 19623 9752 19657
rect 9786 19623 9792 19657
rect 9746 19585 9792 19623
rect 9746 19551 9752 19585
rect 9786 19551 9792 19585
rect 9746 19513 9792 19551
rect 9746 19479 9752 19513
rect 9786 19479 9792 19513
rect 9746 19441 9792 19479
rect 9746 19407 9752 19441
rect 9786 19407 9792 19441
rect 9746 19369 9792 19407
rect 9746 19335 9752 19369
rect 9786 19335 9792 19369
rect 9746 19297 9792 19335
rect 9746 19263 9752 19297
rect 9786 19263 9792 19297
rect 9746 19225 9792 19263
rect 9746 19191 9752 19225
rect 9786 19191 9792 19225
rect 9746 19153 9792 19191
rect 9746 19119 9752 19153
rect 9786 19119 9792 19153
rect 9746 19081 9792 19119
rect 9746 19047 9752 19081
rect 9786 19047 9792 19081
rect 9746 19009 9792 19047
rect 9746 18975 9752 19009
rect 9786 18975 9792 19009
rect 9746 18937 9792 18975
rect 9746 18903 9752 18937
rect 9786 18903 9792 18937
rect 9746 18865 9792 18903
rect 9746 18831 9752 18865
rect 9786 18831 9792 18865
rect 9746 18793 9792 18831
rect 9746 18759 9752 18793
rect 9786 18759 9792 18793
rect 9746 18721 9792 18759
rect 9746 18687 9752 18721
rect 9786 18687 9792 18721
rect 9746 18649 9792 18687
rect 9746 18615 9752 18649
rect 9786 18615 9792 18649
rect 9746 18577 9792 18615
rect 9746 18543 9752 18577
rect 9786 18543 9792 18577
rect 9746 18505 9792 18543
rect 9746 18471 9752 18505
rect 9786 18471 9792 18505
rect 9746 18433 9792 18471
rect 9746 18399 9752 18433
rect 9786 18399 9792 18433
rect 9746 18361 9792 18399
rect 9746 18327 9752 18361
rect 9786 18327 9792 18361
rect 9746 18289 9792 18327
rect 9746 18255 9752 18289
rect 9786 18255 9792 18289
rect 9746 18217 9792 18255
rect 9746 18183 9752 18217
rect 9786 18183 9792 18217
rect 9746 18145 9792 18183
rect 9746 18111 9752 18145
rect 9786 18111 9792 18145
rect 9746 18073 9792 18111
rect 9746 18039 9752 18073
rect 9786 18039 9792 18073
rect 9746 18001 9792 18039
rect 9746 17967 9752 18001
rect 9786 17967 9792 18001
rect 9746 17929 9792 17967
rect 9746 17895 9752 17929
rect 9786 17895 9792 17929
rect 9746 17857 9792 17895
rect 9746 17823 9752 17857
rect 9786 17823 9792 17857
rect 9746 17785 9792 17823
rect 9746 17751 9752 17785
rect 9786 17751 9792 17785
rect 9746 17713 9792 17751
rect 9746 17679 9752 17713
rect 9786 17679 9792 17713
rect 9746 17641 9792 17679
rect 9746 17607 9752 17641
rect 9786 17607 9792 17641
rect 9746 17569 9792 17607
rect 9746 17535 9752 17569
rect 9786 17535 9792 17569
rect 9746 17497 9792 17535
rect 9746 17463 9752 17497
rect 9786 17463 9792 17497
rect 9746 17425 9792 17463
rect 9746 17391 9752 17425
rect 9786 17391 9792 17425
rect 9746 17353 9792 17391
rect 9746 17319 9752 17353
rect 9786 17319 9792 17353
rect 9746 17281 9792 17319
rect 9746 17247 9752 17281
rect 9786 17247 9792 17281
rect 9746 17209 9792 17247
rect 9746 17175 9752 17209
rect 9786 17175 9792 17209
rect 9746 17137 9792 17175
rect 9746 17103 9752 17137
rect 9786 17103 9792 17137
rect 9746 17065 9792 17103
rect 9746 17031 9752 17065
rect 9786 17031 9792 17065
rect 9746 16993 9792 17031
rect 9746 16959 9752 16993
rect 9786 16959 9792 16993
rect 9746 16921 9792 16959
rect 9746 16887 9752 16921
rect 9786 16887 9792 16921
rect 9746 16849 9792 16887
rect 9746 16815 9752 16849
rect 9786 16815 9792 16849
rect 9746 16777 9792 16815
rect 9746 16743 9752 16777
rect 9786 16743 9792 16777
rect 9746 16705 9792 16743
rect 9746 16671 9752 16705
rect 9786 16671 9792 16705
rect 9746 16633 9792 16671
rect 9746 16599 9752 16633
rect 9786 16599 9792 16633
rect 9746 16561 9792 16599
rect 9746 16527 9752 16561
rect 9786 16527 9792 16561
rect 9746 16489 9792 16527
rect 9746 16455 9752 16489
rect 9786 16455 9792 16489
rect 9746 16417 9792 16455
rect 9746 16383 9752 16417
rect 9786 16383 9792 16417
rect 9746 16345 9792 16383
rect 9746 16311 9752 16345
rect 9786 16311 9792 16345
rect 9746 16273 9792 16311
rect 9746 16239 9752 16273
rect 9786 16239 9792 16273
rect 9746 16201 9792 16239
rect 9746 16167 9752 16201
rect 9786 16167 9792 16201
rect 9746 16129 9792 16167
rect 9746 16095 9752 16129
rect 9786 16095 9792 16129
rect 9746 16057 9792 16095
rect 9746 16023 9752 16057
rect 9786 16023 9792 16057
rect 9746 15985 9792 16023
rect 9746 15951 9752 15985
rect 9786 15951 9792 15985
rect 9746 15913 9792 15951
rect 9746 15879 9752 15913
rect 9786 15879 9792 15913
rect 9746 15841 9792 15879
rect 9746 15807 9752 15841
rect 9786 15807 9792 15841
rect 9746 15769 9792 15807
rect 9746 15735 9752 15769
rect 9786 15735 9792 15769
rect 9746 15697 9792 15735
rect 9746 15663 9752 15697
rect 9786 15663 9792 15697
rect 9746 15625 9792 15663
rect 9746 15591 9752 15625
rect 9786 15591 9792 15625
rect 9746 15553 9792 15591
rect 9746 15519 9752 15553
rect 9786 15519 9792 15553
rect 9746 15481 9792 15519
rect 9746 15447 9752 15481
rect 9786 15447 9792 15481
rect 9746 15409 9792 15447
rect 9746 15375 9752 15409
rect 9786 15375 9792 15409
rect 9746 15337 9792 15375
rect 9746 15303 9752 15337
rect 9786 15303 9792 15337
rect 9746 15265 9792 15303
rect 9746 15231 9752 15265
rect 9786 15231 9792 15265
rect 9746 15193 9792 15231
rect 9746 15159 9752 15193
rect 9786 15159 9792 15193
rect 9746 15121 9792 15159
rect 9746 15087 9752 15121
rect 9786 15087 9792 15121
rect 9746 15049 9792 15087
rect 9746 15015 9752 15049
rect 9786 15015 9792 15049
rect 9746 14977 9792 15015
rect 9746 14943 9752 14977
rect 9786 14943 9792 14977
rect 9746 14905 9792 14943
rect 9746 14871 9752 14905
rect 9786 14871 9792 14905
rect 9746 14833 9792 14871
rect 9746 14799 9752 14833
rect 9786 14799 9792 14833
rect 9746 14761 9792 14799
rect 9746 14727 9752 14761
rect 9786 14727 9792 14761
rect 9746 14689 9792 14727
rect 9746 14655 9752 14689
rect 9786 14655 9792 14689
rect 9746 14617 9792 14655
rect 9746 14583 9752 14617
rect 9786 14583 9792 14617
rect 9746 14545 9792 14583
rect 9746 14511 9752 14545
rect 9786 14511 9792 14545
rect 9746 14473 9792 14511
rect 9746 14439 9752 14473
rect 9786 14439 9792 14473
rect 9746 14401 9792 14439
rect 9746 14367 9752 14401
rect 9786 14367 9792 14401
rect 9746 14329 9792 14367
rect 9746 14295 9752 14329
rect 9786 14295 9792 14329
rect 9746 14257 9792 14295
rect 9746 14223 9752 14257
rect 9786 14223 9792 14257
rect 9746 14185 9792 14223
rect 9746 14151 9752 14185
rect 9786 14151 9792 14185
rect 9746 14113 9792 14151
rect 9746 14079 9752 14113
rect 9786 14079 9792 14113
rect 9746 14041 9792 14079
rect 9746 14007 9752 14041
rect 9786 14007 9792 14041
rect 9746 13969 9792 14007
rect 9746 13935 9752 13969
rect 9786 13935 9792 13969
rect 9746 13897 9792 13935
rect 9746 13863 9752 13897
rect 9786 13863 9792 13897
rect 9746 13825 9792 13863
rect 9746 13791 9752 13825
rect 9786 13791 9792 13825
rect 9746 13753 9792 13791
rect 9746 13719 9752 13753
rect 9786 13719 9792 13753
rect 9746 13681 9792 13719
rect 9746 13647 9752 13681
rect 9786 13647 9792 13681
rect 9746 13609 9792 13647
rect 9746 13575 9752 13609
rect 9786 13575 9792 13609
rect 9746 13537 9792 13575
rect 9746 13503 9752 13537
rect 9786 13503 9792 13537
rect 9746 13465 9792 13503
rect 9746 13431 9752 13465
rect 9786 13431 9792 13465
rect 9746 13393 9792 13431
rect 9746 13359 9752 13393
rect 9786 13359 9792 13393
rect 9746 13321 9792 13359
rect 9746 13287 9752 13321
rect 9786 13287 9792 13321
rect 9746 13249 9792 13287
rect 9746 13215 9752 13249
rect 9786 13215 9792 13249
rect 9746 13177 9792 13215
rect 9746 13143 9752 13177
rect 9786 13143 9792 13177
rect 9746 13105 9792 13143
rect 9746 13071 9752 13105
rect 9786 13071 9792 13105
rect 9746 13033 9792 13071
rect 9746 12999 9752 13033
rect 9786 12999 9792 13033
rect 9746 12961 9792 12999
rect 9746 12927 9752 12961
rect 9786 12927 9792 12961
rect 9746 12889 9792 12927
rect 9746 12855 9752 12889
rect 9786 12855 9792 12889
rect 9746 12817 9792 12855
rect 9746 12783 9752 12817
rect 9786 12783 9792 12817
rect 9746 12745 9792 12783
rect 9746 12711 9752 12745
rect 9786 12711 9792 12745
rect 9746 12673 9792 12711
rect 9746 12639 9752 12673
rect 9786 12639 9792 12673
rect 9746 12601 9792 12639
rect 9746 12567 9752 12601
rect 9786 12567 9792 12601
rect 9746 12529 9792 12567
rect 9746 12495 9752 12529
rect 9786 12495 9792 12529
rect 9746 12457 9792 12495
rect 9746 12423 9752 12457
rect 9786 12423 9792 12457
rect 9746 12385 9792 12423
rect 9746 12351 9752 12385
rect 9786 12351 9792 12385
rect 9746 12313 9792 12351
rect 9746 12279 9752 12313
rect 9786 12279 9792 12313
rect 9746 12241 9792 12279
rect 9746 12207 9752 12241
rect 9786 12207 9792 12241
rect 9746 12169 9792 12207
rect 9746 12135 9752 12169
rect 9786 12135 9792 12169
rect 9746 12097 9792 12135
rect 9746 12063 9752 12097
rect 9786 12063 9792 12097
rect 9746 12025 9792 12063
rect 9746 11991 9752 12025
rect 9786 11991 9792 12025
rect 9746 11953 9792 11991
rect 9746 11919 9752 11953
rect 9786 11919 9792 11953
rect 9746 11881 9792 11919
rect 9746 11847 9752 11881
rect 9786 11847 9792 11881
rect 9746 11809 9792 11847
rect 9746 11775 9752 11809
rect 9786 11775 9792 11809
rect 9746 11737 9792 11775
rect 9746 11703 9752 11737
rect 9786 11703 9792 11737
rect 9746 11665 9792 11703
rect 9746 11631 9752 11665
rect 9786 11631 9792 11665
rect 9746 11593 9792 11631
rect 9746 11559 9752 11593
rect 9786 11559 9792 11593
tri 8068 11521 8084 11537 ne
rect 8084 11521 8120 11537
tri 8120 11521 8158 11559 sw
rect 9746 11521 9792 11559
rect 7994 11484 8000 11518
rect 8034 11484 8040 11518
tri 8084 11499 8106 11521 ne
rect 8106 11499 8158 11521
tri 8158 11499 8180 11521 sw
tri 8106 11487 8118 11499 ne
rect 8118 11487 8180 11499
tri 8118 11485 8120 11487 ne
rect 8120 11485 8180 11487
rect 7994 11446 8040 11484
tri 8120 11477 8128 11485 ne
rect 7994 11412 8000 11446
rect 8034 11412 8040 11446
rect 2796 11399 7477 11405
rect 2796 11365 2879 11399
rect 2913 11365 2956 11399
rect 2990 11365 3033 11399
rect 3067 11365 3110 11399
rect 3144 11365 3188 11399
rect 3222 11365 3266 11399
rect 3300 11365 3344 11399
rect 3378 11365 3422 11399
rect 3456 11365 3500 11399
rect 3534 11365 3578 11399
rect 3612 11365 3656 11399
rect 3690 11365 3766 11399
rect 3800 11365 3839 11399
rect 3873 11365 3912 11399
rect 3946 11365 3985 11399
rect 4019 11365 4058 11399
rect 4092 11365 4131 11399
rect 4165 11365 4204 11399
rect 4238 11365 4277 11399
rect 4311 11365 4350 11399
rect 4384 11365 4423 11399
rect 4457 11365 4496 11399
rect 4530 11365 4569 11399
rect 4603 11365 4642 11399
rect 4676 11365 4715 11399
rect 4749 11365 4788 11399
rect 4822 11365 4861 11399
rect 4895 11365 4934 11399
rect 4968 11365 5007 11399
rect 5041 11365 5080 11399
rect 5114 11365 5153 11399
rect 5187 11365 5226 11399
rect 5260 11365 5299 11399
rect 5333 11365 5372 11399
rect 5406 11365 5445 11399
rect 5479 11365 5518 11399
rect 5552 11365 5591 11399
rect 5625 11365 5664 11399
rect 5698 11365 5737 11399
rect 5771 11365 5811 11399
rect 5845 11365 5885 11399
rect 5919 11365 5959 11399
rect 5993 11365 6033 11399
rect 6067 11365 6107 11399
rect 6141 11365 6181 11399
rect 6215 11365 6255 11399
rect 6289 11365 6329 11399
rect 6363 11365 6403 11399
rect 6437 11365 6477 11399
rect 6511 11365 6551 11399
rect 6585 11365 6625 11399
rect 6659 11365 6699 11399
rect 6733 11365 6773 11399
rect 6807 11365 6847 11399
rect 6881 11365 6921 11399
rect 6955 11365 6995 11399
rect 7029 11365 7069 11399
rect 7103 11365 7143 11399
rect 7177 11365 7217 11399
rect 7251 11365 7291 11399
rect 7325 11365 7365 11399
rect 7399 11365 7477 11399
rect 2796 11359 7477 11365
rect 2796 11340 2857 11359
tri 2857 11340 2876 11359 nw
tri 7397 11340 7416 11359 ne
rect 7416 11340 7477 11359
rect 2796 11327 2842 11340
rect 2796 11293 2802 11327
rect 2836 11293 2842 11327
tri 2842 11325 2857 11340 nw
tri 7416 11325 7431 11340 ne
rect 7431 11325 7477 11340
rect 2796 11254 2842 11293
rect 2796 11220 2802 11254
rect 2836 11220 2842 11254
rect 2796 11181 2842 11220
rect 2796 11147 2802 11181
rect 2836 11147 2842 11181
rect 2796 11108 2842 11147
rect 2796 11074 2802 11108
rect 2836 11074 2842 11108
rect 2796 11035 2842 11074
rect 2796 11001 2802 11035
rect 2836 11001 2842 11035
rect 2796 10962 2842 11001
rect 2796 10928 2802 10962
rect 2836 10928 2842 10962
rect 2796 10889 2842 10928
rect 2796 10855 2802 10889
rect 2836 10855 2842 10889
rect 2796 10816 2842 10855
rect 2796 10782 2802 10816
rect 2836 10782 2842 10816
rect 2796 10743 2842 10782
rect 2796 10709 2802 10743
rect 2836 10709 2842 10743
rect 2796 10670 2842 10709
rect 2796 10636 2802 10670
rect 2836 10636 2842 10670
rect 2796 10597 2842 10636
rect 2796 10563 2802 10597
rect 2836 10563 2842 10597
rect 2796 10524 2842 10563
rect 2796 10490 2802 10524
rect 2836 10490 2842 10524
rect 2796 10451 2842 10490
rect 2796 10417 2802 10451
rect 2836 10417 2842 10451
rect 2796 10378 2842 10417
rect 2796 10344 2802 10378
rect 2836 10344 2842 10378
rect 2796 10305 2842 10344
rect 2796 10271 2802 10305
rect 2836 10271 2842 10305
rect 2796 10232 2842 10271
rect 2796 10198 2802 10232
rect 2836 10198 2842 10232
rect 2796 10159 2842 10198
rect 2796 10125 2802 10159
rect 2836 10125 2842 10159
rect 2796 10086 2842 10125
rect 2796 10052 2802 10086
rect 2836 10052 2842 10086
rect 2796 10013 2842 10052
rect 2796 9979 2802 10013
rect 2836 9979 2842 10013
rect 2796 9940 2842 9979
rect 2796 9906 2802 9940
rect 2836 9906 2842 9940
rect 2796 9867 2842 9906
rect 2796 9833 2802 9867
rect 2836 9833 2842 9867
rect 2796 9794 2842 9833
rect 2796 9760 2802 9794
rect 2836 9760 2842 9794
rect 2796 9721 2842 9760
rect 2796 9687 2802 9721
rect 2836 9687 2842 9721
rect 2796 9648 2842 9687
rect 2796 9614 2802 9648
rect 2836 9614 2842 9648
rect 2796 9575 2842 9614
rect 2796 9541 2802 9575
rect 2836 9541 2842 9575
rect 2796 9502 2842 9541
rect 2796 9468 2802 9502
rect 2836 9468 2842 9502
rect 2796 9429 2842 9468
rect 2796 9395 2802 9429
rect 2836 9395 2842 9429
rect 2796 9356 2842 9395
rect 2796 9322 2802 9356
rect 2836 9322 2842 9356
rect 2796 9283 2842 9322
rect 2796 9249 2802 9283
rect 2836 9249 2842 9283
rect 2796 9210 2842 9249
rect 2796 9176 2802 9210
rect 2836 9176 2842 9210
rect 2796 9137 2842 9176
rect 2796 9103 2802 9137
rect 2836 9103 2842 9137
rect 2796 9064 2842 9103
rect 2796 9030 2802 9064
rect 2836 9030 2842 9064
rect 2796 8991 2842 9030
rect 2796 8957 2802 8991
rect 2836 8957 2842 8991
rect 2796 8918 2842 8957
rect 2796 8884 2802 8918
rect 2836 8884 2842 8918
rect 2796 8845 2842 8884
rect 2796 8811 2802 8845
rect 2836 8811 2842 8845
rect 2796 8772 2842 8811
rect 2796 8738 2802 8772
rect 2836 8738 2842 8772
rect 2796 8699 2842 8738
rect 2796 8665 2802 8699
rect 2836 8665 2842 8699
rect 2796 8626 2842 8665
rect 2796 8592 2802 8626
rect 2836 8592 2842 8626
rect 2796 8553 2842 8592
rect 2796 8519 2802 8553
rect 2836 8519 2842 8553
rect 2796 8480 2842 8519
rect 2796 8446 2802 8480
rect 2836 8446 2842 8480
rect 2796 8407 2842 8446
rect 2796 8373 2802 8407
rect 2836 8373 2842 8407
rect 2796 8334 2842 8373
rect 2796 8300 2802 8334
rect 2836 8300 2842 8334
rect 2796 8261 2842 8300
rect 2796 8227 2802 8261
rect 2836 8227 2842 8261
rect 2796 8188 2842 8227
rect 2796 8154 2802 8188
rect 2836 8154 2842 8188
rect 2796 8115 2842 8154
rect 7431 11291 7437 11325
rect 7471 11291 7477 11325
rect 7431 11251 7477 11291
rect 7431 11217 7437 11251
rect 7471 11217 7477 11251
rect 7431 11177 7477 11217
rect 7431 11143 7437 11177
rect 7471 11143 7477 11177
rect 7431 11103 7477 11143
rect 7431 11069 7437 11103
rect 7471 11069 7477 11103
rect 7431 11029 7477 11069
rect 7431 10995 7437 11029
rect 7471 10995 7477 11029
rect 7431 10955 7477 10995
rect 7431 10921 7437 10955
rect 7471 10921 7477 10955
rect 7431 10880 7477 10921
rect 7431 10846 7437 10880
rect 7471 10846 7477 10880
rect 7431 10805 7477 10846
rect 7431 10771 7437 10805
rect 7471 10771 7477 10805
rect 7431 10730 7477 10771
rect 7431 10696 7437 10730
rect 7471 10696 7477 10730
rect 7431 10655 7477 10696
rect 7431 10621 7437 10655
rect 7471 10621 7477 10655
rect 7431 10580 7477 10621
rect 7431 10546 7437 10580
rect 7471 10546 7477 10580
rect 7431 10505 7477 10546
rect 7431 10471 7437 10505
rect 7471 10471 7477 10505
rect 7431 10401 7477 10471
rect 7431 10367 7437 10401
rect 7471 10367 7477 10401
rect 7431 10328 7477 10367
rect 7431 10294 7437 10328
rect 7471 10294 7477 10328
rect 7431 10255 7477 10294
rect 7431 10221 7437 10255
rect 7471 10221 7477 10255
rect 7431 10182 7477 10221
rect 7431 10148 7437 10182
rect 7471 10148 7477 10182
rect 7431 10108 7477 10148
rect 7431 10074 7437 10108
rect 7471 10074 7477 10108
rect 7431 10034 7477 10074
rect 7431 10000 7437 10034
rect 7471 10000 7477 10034
rect 7431 9960 7477 10000
rect 7431 9926 7437 9960
rect 7471 9926 7477 9960
rect 7431 9886 7477 9926
rect 7431 9852 7437 9886
rect 7471 9852 7477 9886
rect 7431 9812 7477 9852
rect 7431 9778 7437 9812
rect 7471 9778 7477 9812
rect 7431 9738 7477 9778
rect 7431 9704 7437 9738
rect 7471 9704 7477 9738
rect 7431 9664 7477 9704
rect 7431 9630 7437 9664
rect 7471 9630 7477 9664
rect 7431 9590 7477 9630
rect 7431 9556 7437 9590
rect 7471 9556 7477 9590
rect 7431 9516 7477 9556
rect 7431 9482 7437 9516
rect 7471 9482 7477 9516
rect 7431 9442 7477 9482
rect 7431 9408 7437 9442
rect 7471 9408 7477 9442
rect 7431 9368 7477 9408
rect 7431 9334 7437 9368
rect 7471 9334 7477 9368
rect 7431 9294 7477 9334
rect 7431 9260 7437 9294
rect 7471 9260 7477 9294
rect 7431 9220 7477 9260
rect 7431 9186 7437 9220
rect 7471 9186 7477 9220
rect 7431 9146 7477 9186
rect 7431 9112 7437 9146
rect 7471 9112 7477 9146
rect 7431 9072 7477 9112
rect 7431 9038 7437 9072
rect 7471 9038 7477 9072
rect 7431 8998 7477 9038
rect 7431 8964 7437 8998
rect 7471 8964 7477 8998
rect 7431 8924 7477 8964
rect 7431 8890 7437 8924
rect 7471 8890 7477 8924
rect 7431 8850 7477 8890
rect 7431 8816 7437 8850
rect 7471 8816 7477 8850
rect 7431 8776 7477 8816
rect 7431 8742 7437 8776
rect 7471 8742 7477 8776
rect 7431 8702 7477 8742
rect 7431 8668 7437 8702
rect 7471 8668 7477 8702
rect 7431 8628 7477 8668
rect 7431 8594 7437 8628
rect 7471 8594 7477 8628
rect 7431 8554 7477 8594
rect 7431 8520 7437 8554
rect 7471 8520 7477 8554
rect 7431 8480 7477 8520
rect 7431 8446 7437 8480
rect 7471 8446 7477 8480
rect 7431 8406 7477 8446
rect 7431 8372 7437 8406
rect 7471 8372 7477 8406
rect 7431 8332 7477 8372
rect 7431 8298 7437 8332
rect 7471 8298 7477 8332
rect 7431 8258 7477 8298
rect 7431 8224 7437 8258
rect 7471 8224 7477 8258
rect 7431 8184 7477 8224
rect 7431 8150 7437 8184
rect 7471 8150 7477 8184
rect 2796 8081 2802 8115
rect 2836 8081 2842 8115
rect 2796 8042 2842 8081
rect 2796 8008 2802 8042
rect 2836 8008 2842 8042
rect 2796 7969 2842 8008
rect 2796 7935 2802 7969
rect 2836 7935 2842 7969
rect 2796 7896 2842 7935
rect 2796 7862 2802 7896
rect 2836 7862 2842 7896
rect 2796 7823 2842 7862
rect 2796 7789 2802 7823
rect 2836 7789 2842 7823
rect 2796 7750 2842 7789
rect 2796 7716 2802 7750
rect 2836 7716 2842 7750
rect 6744 8094 6790 8126
rect 7431 8118 7477 8150
rect 6744 8060 6750 8094
rect 6784 8060 6790 8094
rect 7016 8112 7477 8118
rect 7016 8078 7048 8112
rect 7082 8078 7126 8112
rect 7160 8078 7204 8112
rect 7238 8078 7282 8112
rect 7316 8078 7360 8112
rect 7394 8078 7477 8112
rect 7016 8072 7477 8078
rect 7994 11374 8040 11412
rect 7994 11340 8000 11374
rect 8034 11340 8040 11374
rect 7994 11302 8040 11340
rect 7994 11268 8000 11302
rect 8034 11268 8040 11302
rect 7994 11230 8040 11268
rect 7994 11196 8000 11230
rect 8034 11196 8040 11230
rect 7994 11158 8040 11196
rect 7994 11124 8000 11158
rect 8034 11124 8040 11158
rect 7994 11086 8040 11124
rect 7994 11052 8000 11086
rect 8034 11052 8040 11086
rect 7994 11014 8040 11052
rect 7994 10980 8000 11014
rect 8034 10980 8040 11014
rect 7994 10942 8040 10980
rect 7994 10908 8000 10942
rect 8034 10908 8040 10942
rect 7994 10870 8040 10908
rect 7994 10836 8000 10870
rect 8034 10836 8040 10870
rect 7994 10798 8040 10836
rect 7994 10764 8000 10798
rect 8034 10764 8040 10798
rect 7994 10726 8040 10764
rect 7994 10692 8000 10726
rect 8034 10692 8040 10726
rect 7994 10654 8040 10692
rect 7994 10620 8000 10654
rect 8034 10620 8040 10654
rect 7994 10582 8040 10620
rect 7994 10548 8000 10582
rect 8034 10548 8040 10582
rect 7994 10510 8040 10548
rect 7994 10476 8000 10510
rect 8034 10476 8040 10510
rect 7994 10438 8040 10476
rect 7994 10404 8000 10438
rect 8034 10404 8040 10438
rect 7994 10366 8040 10404
rect 7994 10332 8000 10366
rect 8034 10332 8040 10366
rect 7994 10294 8040 10332
rect 7994 10260 8000 10294
rect 8034 10260 8040 10294
rect 7994 10222 8040 10260
rect 7994 10188 8000 10222
rect 8034 10188 8040 10222
rect 7994 10150 8040 10188
rect 7994 10116 8000 10150
rect 8034 10116 8040 10150
rect 7994 10078 8040 10116
rect 7994 10044 8000 10078
rect 8034 10044 8040 10078
rect 7994 10006 8040 10044
rect 7994 9972 8000 10006
rect 8034 9972 8040 10006
rect 7994 9934 8040 9972
rect 7994 9900 8000 9934
rect 8034 9900 8040 9934
rect 7994 9862 8040 9900
rect 7994 9828 8000 9862
rect 8034 9828 8040 9862
rect 7994 9790 8040 9828
rect 7994 9756 8000 9790
rect 8034 9756 8040 9790
rect 7994 9718 8040 9756
rect 7994 9684 8000 9718
rect 8034 9684 8040 9718
rect 7994 9646 8040 9684
rect 7994 9612 8000 9646
rect 8034 9612 8040 9646
rect 7994 9574 8040 9612
rect 7994 9540 8000 9574
rect 8034 9540 8040 9574
rect 7994 9502 8040 9540
rect 7994 9468 8000 9502
rect 8034 9468 8040 9502
rect 7994 9430 8040 9468
rect 7994 9396 8000 9430
rect 8034 9396 8040 9430
rect 7994 9358 8040 9396
rect 7994 9324 8000 9358
rect 8034 9324 8040 9358
rect 7994 9286 8040 9324
rect 7994 9252 8000 9286
rect 8034 9252 8040 9286
rect 7994 9214 8040 9252
rect 7994 9180 8000 9214
rect 8034 9180 8040 9214
rect 7994 9142 8040 9180
rect 7994 9108 8000 9142
rect 8034 9108 8040 9142
rect 7994 9070 8040 9108
rect 7994 9036 8000 9070
rect 8034 9036 8040 9070
rect 7994 8998 8040 9036
rect 7994 8964 8000 8998
rect 8034 8964 8040 8998
rect 7994 8926 8040 8964
rect 7994 8892 8000 8926
rect 8034 8892 8040 8926
rect 7994 8854 8040 8892
rect 7994 8820 8000 8854
rect 8034 8820 8040 8854
rect 7994 8782 8040 8820
rect 7994 8748 8000 8782
rect 8034 8748 8040 8782
rect 7994 8710 8040 8748
rect 7994 8676 8000 8710
rect 8034 8676 8040 8710
rect 7994 8638 8040 8676
rect 7994 8604 8000 8638
rect 8034 8604 8040 8638
rect 7994 8566 8040 8604
rect 7994 8532 8000 8566
rect 8034 8532 8040 8566
rect 7994 8494 8040 8532
rect 7994 8460 8000 8494
rect 8034 8460 8040 8494
rect 7994 8422 8040 8460
rect 7994 8388 8000 8422
rect 8034 8388 8040 8422
rect 7994 8350 8040 8388
rect 7994 8316 8000 8350
rect 8034 8316 8040 8350
rect 7994 8278 8040 8316
rect 7994 8244 8000 8278
rect 8034 8244 8040 8278
rect 7994 8206 8040 8244
rect 7994 8172 8000 8206
rect 8034 8172 8040 8206
rect 7994 8134 8040 8172
rect 7994 8100 8000 8134
rect 8034 8100 8040 8134
rect 6744 7992 6790 8060
rect 6744 7958 6750 7992
rect 6784 7958 6790 7992
rect 6744 7888 6790 7958
rect 6744 7854 6750 7888
rect 6784 7854 6790 7888
rect 6744 7815 6790 7854
rect 6744 7781 6750 7815
rect 6784 7781 6790 7815
rect 6744 7742 6790 7781
rect 2796 7677 2842 7716
rect 2796 7643 2802 7677
rect 2836 7643 2842 7677
rect 2796 7604 2842 7643
rect 2796 7570 2802 7604
rect 2836 7570 2842 7604
rect 2796 7531 2842 7570
rect 2796 7497 2802 7531
rect 2836 7497 2842 7531
rect 2796 7458 2842 7497
rect 2796 7424 2802 7458
rect 2836 7424 2842 7458
rect 2796 7385 2842 7424
rect 2796 7351 2802 7385
rect 2836 7351 2842 7385
rect 2796 7312 2842 7351
rect 2796 7278 2802 7312
rect 2836 7278 2842 7312
rect 2796 7239 2842 7278
rect 2796 7205 2802 7239
rect 2836 7205 2842 7239
rect 2796 7166 2842 7205
rect 2796 7132 2802 7166
rect 2836 7132 2842 7166
rect 2796 7093 2842 7132
rect 2796 7059 2802 7093
rect 2836 7059 2842 7093
rect 2796 7020 2842 7059
rect 2796 6986 2802 7020
rect 2836 6986 2842 7020
rect 2796 6947 2842 6986
rect 2796 6913 2802 6947
rect 2836 6913 2842 6947
rect 2796 6874 2842 6913
rect 2796 6840 2802 6874
rect 2836 6840 2842 6874
rect 2796 6801 2842 6840
rect 2796 6767 2802 6801
rect 2836 6767 2842 6801
rect 2796 6729 2842 6767
rect 2796 6695 2802 6729
rect 2836 6695 2842 6729
rect 2796 6657 2842 6695
rect 2796 6623 2802 6657
rect 2836 6623 2842 6657
rect 2796 6585 2842 6623
rect 2796 6551 2802 6585
rect 2836 6551 2842 6585
rect 2796 6513 2842 6551
rect 2796 6479 2802 6513
rect 2836 6479 2842 6513
rect 2796 6441 2842 6479
rect 2796 6407 2802 6441
rect 2836 6407 2842 6441
rect 2796 6369 2842 6407
rect 2796 6335 2802 6369
rect 2836 6335 2842 6369
rect 2796 6297 2842 6335
rect 2796 6263 2802 6297
rect 2836 6263 2842 6297
rect 2796 6225 2842 6263
rect 2796 6191 2802 6225
rect 2836 6191 2842 6225
rect 2796 6153 2842 6191
rect 2796 6119 2802 6153
rect 2836 6119 2842 6153
rect 2796 6081 2842 6119
rect 2796 6047 2802 6081
rect 2836 6047 2842 6081
rect 2796 6009 2842 6047
rect 2796 5975 2802 6009
rect 2836 5975 2842 6009
rect 2796 5937 2842 5975
rect 2796 5903 2802 5937
rect 2836 5903 2842 5937
rect 2796 5865 2842 5903
rect 2796 5831 2802 5865
rect 2836 5831 2842 5865
rect 2796 5793 2842 5831
rect 2796 5759 2802 5793
rect 2836 5759 2842 5793
rect 2796 5721 2842 5759
rect 2796 5687 2802 5721
rect 2836 5687 2842 5721
rect 2796 5649 2842 5687
rect 2796 5615 2802 5649
rect 2836 5615 2842 5649
rect 2796 5577 2842 5615
rect 2796 5543 2802 5577
rect 2836 5543 2842 5577
rect 2796 5505 2842 5543
rect 2796 5471 2802 5505
rect 2836 5471 2842 5505
rect 2796 5433 2842 5471
rect 2796 5399 2802 5433
rect 2836 5399 2842 5433
rect 2796 5361 2842 5399
rect 2796 5327 2802 5361
rect 2836 5327 2842 5361
rect 2796 5289 2842 5327
rect 2796 5255 2802 5289
rect 2836 5255 2842 5289
rect 3076 7723 6533 7729
rect 3076 7689 3164 7723
rect 3198 7689 3246 7723
rect 3280 7689 3328 7723
rect 3362 7689 3411 7723
rect 3445 7689 3494 7723
rect 3528 7689 3604 7723
rect 3638 7689 3676 7723
rect 3710 7689 3748 7723
rect 3782 7689 3820 7723
rect 3854 7689 3892 7723
rect 3926 7689 3964 7723
rect 3998 7689 4036 7723
rect 4070 7689 4108 7723
rect 4142 7689 4180 7723
rect 4214 7689 4252 7723
rect 4286 7689 4324 7723
rect 4358 7689 4396 7723
rect 4430 7689 4468 7723
rect 4502 7689 4540 7723
rect 4574 7689 4612 7723
rect 4646 7689 4684 7723
rect 4718 7710 4756 7723
rect 4790 7710 4828 7723
rect 4862 7710 4900 7723
rect 4934 7710 4972 7723
rect 5006 7710 5044 7723
rect 5078 7710 5116 7723
rect 5150 7710 5188 7723
rect 5222 7710 5260 7723
rect 4718 7689 4728 7710
rect 4790 7689 4800 7710
rect 4862 7689 4871 7710
rect 4934 7689 4942 7710
rect 5006 7689 5013 7710
rect 5078 7689 5084 7710
rect 5150 7689 5155 7710
rect 5222 7689 5226 7710
rect 5294 7689 5332 7723
rect 5366 7689 5404 7723
rect 5438 7689 5476 7723
rect 5510 7689 5548 7723
rect 5582 7689 5620 7723
rect 5654 7719 5692 7723
rect 5726 7719 5764 7723
rect 5798 7719 5836 7723
rect 5870 7689 5908 7723
rect 5942 7689 5980 7723
rect 6014 7689 6053 7723
rect 6087 7689 6126 7723
rect 6160 7700 6199 7723
rect 6233 7700 6272 7723
rect 6306 7700 6345 7723
rect 6379 7700 6418 7723
rect 6160 7689 6197 7700
rect 3076 7683 4728 7689
rect 3076 7669 3142 7683
tri 3142 7669 3156 7683 nw
tri 4688 7669 4702 7683 ne
rect 4702 7669 4728 7683
rect 3076 7651 3124 7669
tri 3124 7651 3142 7669 nw
tri 4702 7651 4720 7669 ne
rect 4720 7658 4728 7669
rect 4780 7658 4800 7689
rect 4852 7658 4871 7689
rect 4923 7658 4942 7689
rect 4994 7658 5013 7689
rect 5065 7658 5084 7689
rect 5136 7658 5155 7689
rect 5207 7658 5226 7689
rect 5278 7683 5649 7689
rect 5278 7669 5410 7683
tri 5410 7669 5424 7683 nw
tri 5614 7669 5628 7683 ne
rect 5628 7669 5649 7683
rect 5278 7658 5391 7669
rect 4720 7651 5391 7658
rect 3076 7617 3082 7651
rect 3116 7617 3122 7651
tri 3122 7649 3124 7651 nw
tri 4720 7649 4722 7651 ne
rect 3076 7577 3122 7617
rect 3076 7543 3082 7577
rect 3116 7543 3122 7577
rect 3076 7503 3122 7543
rect 3076 7469 3082 7503
rect 3116 7469 3122 7503
rect 3076 7429 3122 7469
rect 4722 7636 5350 7651
rect 4722 7584 4728 7636
rect 4780 7584 4800 7636
rect 4852 7584 4871 7636
rect 4923 7584 4942 7636
rect 4994 7584 5013 7636
rect 5065 7584 5084 7636
rect 5136 7584 5155 7636
rect 5207 7584 5226 7636
rect 5278 7617 5350 7636
rect 5384 7650 5391 7651
tri 5391 7650 5410 7669 nw
tri 5628 7650 5647 7669 ne
rect 5647 7667 5649 7669
rect 5701 7667 5723 7689
rect 5775 7667 5797 7689
rect 5849 7683 6197 7689
rect 5849 7669 5870 7683
tri 5870 7669 5884 7683 nw
tri 6162 7669 6176 7683 ne
rect 6176 7669 6197 7683
rect 5849 7667 5851 7669
rect 5647 7650 5851 7667
tri 5851 7650 5870 7669 nw
tri 6176 7650 6195 7669 ne
rect 6195 7650 6197 7669
rect 5384 7617 5390 7650
tri 5390 7649 5391 7650 nw
tri 5647 7649 5648 7650 ne
rect 5278 7584 5390 7617
rect 4722 7578 5390 7584
rect 4722 7562 5350 7578
rect 4722 7510 4728 7562
rect 4780 7510 4800 7562
rect 4852 7510 4871 7562
rect 4923 7510 4942 7562
rect 4994 7510 5013 7562
rect 5065 7510 5084 7562
rect 5136 7510 5155 7562
rect 5207 7510 5226 7562
rect 5278 7544 5350 7562
rect 5384 7544 5390 7578
rect 5278 7510 5390 7544
rect 4722 7505 5390 7510
rect 4722 7488 5350 7505
rect 3076 7395 3082 7429
rect 3116 7395 3122 7429
rect 3076 7355 3122 7395
rect 3076 7321 3082 7355
rect 3116 7321 3122 7355
rect 3076 7281 3122 7321
rect 3262 7286 4554 7457
rect 4722 7436 4728 7488
rect 4780 7436 4800 7488
rect 4852 7436 4871 7488
rect 4923 7436 4942 7488
rect 4994 7436 5013 7488
rect 5065 7436 5084 7488
rect 5136 7436 5155 7488
rect 5207 7436 5226 7488
rect 5278 7471 5350 7488
rect 5384 7471 5390 7505
rect 5278 7436 5390 7471
rect 4722 7432 5390 7436
rect 4722 7414 5350 7432
rect 4722 7362 4728 7414
rect 4780 7362 4800 7414
rect 4852 7362 4871 7414
rect 4923 7362 4942 7414
rect 4994 7362 5013 7414
rect 5065 7362 5084 7414
rect 5136 7362 5155 7414
rect 5207 7362 5226 7414
rect 5278 7398 5350 7414
rect 5384 7398 5390 7432
rect 5278 7362 5390 7398
rect 4722 7359 5390 7362
rect 4722 7340 5350 7359
rect 4722 7288 4728 7340
rect 4780 7288 4800 7340
rect 4852 7288 4871 7340
rect 4923 7288 4942 7340
rect 4994 7288 5013 7340
rect 5065 7288 5084 7340
rect 5136 7288 5155 7340
rect 5207 7288 5226 7340
rect 5278 7325 5350 7340
rect 5384 7325 5390 7359
rect 5278 7288 5390 7325
rect 4722 7286 5390 7288
rect 5648 7644 5850 7650
tri 5850 7649 5851 7650 nw
tri 6195 7649 6196 7650 ne
rect 5648 7592 5649 7644
rect 5701 7592 5723 7644
rect 5775 7592 5797 7644
rect 5849 7592 5850 7644
rect 5648 7569 5850 7592
rect 5648 7517 5649 7569
rect 5701 7517 5723 7569
rect 5775 7517 5797 7569
rect 5849 7517 5850 7569
rect 5648 7494 5850 7517
rect 5648 7442 5649 7494
rect 5701 7442 5723 7494
rect 5775 7442 5797 7494
rect 5849 7442 5850 7494
rect 5648 7419 5850 7442
rect 5648 7367 5649 7419
rect 5701 7367 5723 7419
rect 5775 7367 5797 7419
rect 5849 7367 5850 7419
rect 5648 7344 5850 7367
rect 5648 7292 5649 7344
rect 5701 7292 5723 7344
rect 5775 7292 5797 7344
rect 5849 7292 5850 7344
rect 5648 7286 5850 7292
rect 6196 7648 6197 7650
rect 6249 7648 6271 7700
rect 6323 7648 6345 7700
rect 6397 7689 6418 7700
rect 6452 7689 6481 7723
rect 6397 7671 6481 7689
rect 6397 7650 6533 7671
rect 6397 7648 6490 7650
rect 6524 7648 6533 7650
rect 6196 7629 6481 7648
rect 6196 7577 6197 7629
rect 6249 7577 6271 7629
rect 6323 7577 6345 7629
rect 6397 7596 6481 7629
rect 6397 7577 6533 7596
rect 6196 7573 6490 7577
rect 6524 7573 6533 7577
rect 6196 7558 6481 7573
rect 6196 7506 6197 7558
rect 6249 7506 6271 7558
rect 6323 7506 6345 7558
rect 6397 7521 6481 7558
rect 6397 7506 6533 7521
rect 6196 7504 6533 7506
rect 6196 7497 6490 7504
rect 6524 7497 6533 7504
rect 6196 7487 6481 7497
rect 6196 7435 6197 7487
rect 6249 7435 6271 7487
rect 6323 7435 6345 7487
rect 6397 7445 6481 7487
rect 6397 7435 6533 7445
rect 6196 7431 6533 7435
rect 6196 7421 6490 7431
rect 6524 7421 6533 7431
rect 6196 7416 6481 7421
rect 6196 7364 6197 7416
rect 6249 7364 6271 7416
rect 6323 7364 6345 7416
rect 6397 7369 6481 7416
rect 6397 7364 6533 7369
rect 6196 7358 6533 7364
rect 6196 7345 6490 7358
rect 6524 7345 6533 7358
rect 6196 7293 6197 7345
rect 6249 7293 6271 7345
rect 6323 7293 6345 7345
rect 6397 7293 6481 7345
rect 3076 7247 3082 7281
rect 3116 7247 3122 7281
tri 5310 7252 5344 7286 ne
rect 5344 7252 5350 7286
rect 5384 7252 5390 7286
rect 3076 7207 3122 7247
rect 3076 7173 3082 7207
rect 3116 7173 3122 7207
rect 3076 7133 3122 7173
rect 3076 7099 3082 7133
rect 3116 7099 3122 7133
rect 3076 7059 3122 7099
rect 3076 7025 3082 7059
rect 3116 7025 3122 7059
rect 3076 6985 3122 7025
rect 3076 6951 3082 6985
rect 3116 6951 3122 6985
rect 3076 6911 3122 6951
rect 3076 6877 3082 6911
rect 3116 6877 3122 6911
rect 3076 6837 3122 6877
rect 3076 6803 3082 6837
rect 3116 6803 3122 6837
rect 3076 6763 3122 6803
rect 3076 6729 3082 6763
rect 3116 6729 3122 6763
rect 3076 6689 3122 6729
rect 3076 6655 3082 6689
rect 3116 6655 3122 6689
rect 3076 6615 3122 6655
rect 3076 6581 3082 6615
rect 3116 6581 3122 6615
rect 3076 6542 3122 6581
rect 3076 6508 3082 6542
rect 3116 6508 3122 6542
rect 3076 6469 3122 6508
rect 3076 6435 3082 6469
rect 3116 6435 3122 6469
rect 3076 6396 3122 6435
rect 3076 6362 3082 6396
rect 3116 6362 3122 6396
rect 3076 6323 3122 6362
rect 3076 6289 3082 6323
rect 3116 6289 3122 6323
rect 3076 6250 3122 6289
rect 3076 6216 3082 6250
rect 3116 6216 3122 6250
rect 3076 6177 3122 6216
rect 3076 6143 3082 6177
rect 3116 6143 3122 6177
rect 3076 6104 3122 6143
rect 3076 6070 3082 6104
rect 3116 6070 3122 6104
rect 3076 6031 3122 6070
rect 3076 5997 3082 6031
rect 3116 5997 3122 6031
rect 3076 5958 3122 5997
rect 3076 5924 3082 5958
rect 3116 5924 3122 5958
rect 3076 5885 3122 5924
rect 3076 5851 3082 5885
rect 3116 5851 3122 5885
rect 3076 5812 3122 5851
rect 3076 5778 3082 5812
rect 3116 5778 3122 5812
rect 3076 5739 3122 5778
rect 3076 5705 3082 5739
rect 3116 5705 3122 5739
rect 3847 7193 3899 7249
rect 3847 7159 3856 7193
rect 3890 7159 3899 7193
rect 3847 7119 3899 7159
rect 3847 7085 3856 7119
rect 3890 7085 3899 7119
rect 3847 7045 3899 7085
rect 3847 7011 3856 7045
rect 3890 7011 3899 7045
rect 3847 6971 3899 7011
rect 3847 6937 3856 6971
rect 3890 6937 3899 6971
rect 3847 6897 3899 6937
rect 3847 6863 3856 6897
rect 3890 6863 3899 6897
rect 3847 6823 3899 6863
rect 3847 6789 3856 6823
rect 3890 6789 3899 6823
rect 3847 6749 3899 6789
rect 3847 6715 3856 6749
rect 3890 6715 3899 6749
rect 3847 6675 3899 6715
rect 3847 6641 3856 6675
rect 3890 6641 3899 6675
rect 3847 6601 3899 6641
rect 3847 6567 3856 6601
rect 3890 6567 3899 6601
rect 3847 6527 3899 6567
rect 3847 6523 3856 6527
rect 3890 6523 3899 6527
rect 3847 6459 3899 6471
rect 3847 6377 3899 6407
rect 3847 6343 3856 6377
rect 3890 6343 3899 6377
rect 3847 6302 3899 6343
rect 3847 6268 3856 6302
rect 3890 6268 3899 6302
rect 3847 6227 3899 6268
rect 3847 6193 3856 6227
rect 3890 6193 3899 6227
rect 3847 6152 3899 6193
rect 3847 6118 3856 6152
rect 3890 6118 3899 6152
rect 3847 6077 3899 6118
rect 3847 6043 3856 6077
rect 3890 6043 3899 6077
rect 3847 6002 3899 6043
rect 3847 5968 3856 6002
rect 3890 5968 3899 6002
rect 3847 5927 3899 5968
rect 3847 5893 3856 5927
rect 3890 5893 3899 5927
rect 3847 5852 3899 5893
rect 3847 5818 3856 5852
rect 3890 5818 3899 5852
rect 3847 5777 3899 5818
rect 3847 5743 3856 5777
rect 3890 5743 3899 5777
rect 3847 5731 3899 5743
rect 4577 7193 4629 7249
rect 4577 7159 4586 7193
rect 4620 7159 4629 7193
rect 4577 7119 4629 7159
rect 4577 7085 4586 7119
rect 4620 7085 4629 7119
rect 4577 7045 4629 7085
rect 4577 7011 4586 7045
rect 4620 7011 4629 7045
rect 4577 6971 4629 7011
rect 4577 6937 4586 6971
rect 4620 6937 4629 6971
rect 4577 6897 4629 6937
rect 4577 6863 4586 6897
rect 4620 6863 4629 6897
rect 4577 6823 4629 6863
rect 4577 6789 4586 6823
rect 4620 6789 4629 6823
rect 4577 6749 4629 6789
rect 4577 6715 4586 6749
rect 4620 6715 4629 6749
rect 4577 6675 4629 6715
rect 4577 6641 4586 6675
rect 4620 6641 4629 6675
rect 4577 6601 4629 6641
rect 4577 6567 4586 6601
rect 4620 6567 4629 6601
rect 4577 6527 4629 6567
rect 4577 6523 4586 6527
rect 4620 6523 4629 6527
rect 4577 6459 4629 6471
rect 4577 6377 4629 6407
rect 4577 6343 4586 6377
rect 4620 6343 4629 6377
rect 4577 6302 4629 6343
rect 4577 6268 4586 6302
rect 4620 6268 4629 6302
rect 4577 6227 4629 6268
rect 4577 6193 4586 6227
rect 4620 6193 4629 6227
rect 4577 6152 4629 6193
rect 4577 6118 4586 6152
rect 4620 6118 4629 6152
rect 4577 6077 4629 6118
rect 4577 6043 4586 6077
rect 4620 6043 4629 6077
rect 4577 6002 4629 6043
rect 4577 5968 4586 6002
rect 4620 5968 4629 6002
rect 4577 5927 4629 5968
rect 4577 5893 4586 5927
rect 4620 5893 4629 5927
rect 4577 5852 4629 5893
rect 4577 5818 4586 5852
rect 4620 5818 4629 5852
rect 4577 5777 4629 5818
rect 4577 5743 4586 5777
rect 4620 5743 4629 5777
rect 4577 5731 4629 5743
rect 5344 7213 5390 7252
rect 5344 7179 5350 7213
rect 5384 7179 5390 7213
rect 5653 7181 5699 7286
rect 6196 7285 6533 7293
rect 6196 7251 6490 7285
rect 6524 7251 6533 7285
rect 6196 7212 6533 7251
rect 5344 7140 5390 7179
rect 5344 7106 5350 7140
rect 5384 7106 5390 7140
rect 6196 7178 6490 7212
rect 6524 7178 6533 7212
rect 6196 7139 6533 7178
rect 6196 7137 6490 7139
rect 6391 7129 6490 7137
rect 5344 7067 5390 7106
tri 6447 7105 6471 7129 ne
rect 6471 7105 6490 7129
rect 6524 7105 6533 7139
tri 6471 7095 6481 7105 ne
rect 5344 7033 5350 7067
rect 5384 7033 5390 7067
rect 6481 7066 6533 7105
rect 5344 6994 5390 7033
rect 5344 6960 5350 6994
rect 5384 6960 5390 6994
rect 5344 6921 5390 6960
rect 5344 6887 5350 6921
rect 5384 6887 5390 6921
rect 5344 6848 5390 6887
rect 5344 6814 5350 6848
rect 5384 6814 5390 6848
rect 5344 6775 5390 6814
rect 5344 6741 5350 6775
rect 5384 6741 5390 6775
rect 5344 6702 5390 6741
rect 5344 6668 5350 6702
rect 5384 6668 5390 6702
rect 5344 6629 5390 6668
rect 5344 6595 5350 6629
rect 5384 6595 5390 6629
rect 6094 7046 6146 7058
rect 6094 7012 6100 7046
rect 6134 7012 6146 7046
rect 6094 6954 6146 7012
rect 6094 6920 6100 6954
rect 6134 6920 6146 6954
rect 6094 6862 6146 6920
rect 6094 6828 6100 6862
rect 6134 6828 6146 6862
rect 6094 6770 6146 6828
rect 6094 6736 6100 6770
rect 6134 6736 6146 6770
rect 6094 6628 6146 6736
rect 6481 7032 6490 7066
rect 6524 7032 6533 7066
rect 6481 6993 6533 7032
rect 6481 6959 6490 6993
rect 6524 6959 6533 6993
rect 6481 6920 6533 6959
rect 6481 6886 6490 6920
rect 6524 6886 6533 6920
rect 6481 6847 6533 6886
rect 6481 6813 6490 6847
rect 6524 6813 6533 6847
rect 6481 6774 6533 6813
rect 6481 6740 6490 6774
rect 6524 6740 6533 6774
rect 6196 6671 6269 6723
rect 6321 6671 6369 6723
rect 6421 6671 6427 6723
rect 6481 6701 6533 6740
rect 6481 6667 6490 6701
rect 6524 6667 6533 6701
tri 6146 6628 6161 6643 sw
rect 6481 6628 6533 6667
rect 6094 6609 6161 6628
tri 6161 6609 6180 6628 sw
rect 5344 6556 5390 6595
rect 5344 6522 5350 6556
rect 5384 6522 5390 6556
rect 5344 6483 5390 6522
rect 5344 6449 5350 6483
rect 5384 6449 5390 6483
rect 5809 6589 5861 6595
rect 6094 6557 6401 6609
tri 6293 6555 6295 6557 ne
rect 6295 6555 6399 6557
tri 6399 6555 6401 6557 nw
rect 6481 6594 6490 6628
rect 6524 6594 6533 6628
rect 6481 6555 6533 6594
rect 5809 6525 5861 6537
tri 6295 6523 6327 6555 ne
rect 5809 6467 5861 6473
rect 6091 6506 6156 6518
rect 6091 6472 6100 6506
rect 6134 6472 6156 6506
rect 5344 6409 5390 6449
rect 5344 6375 5350 6409
rect 5384 6375 5390 6409
rect 5344 6335 5390 6375
rect 5344 6301 5350 6335
rect 5384 6301 5390 6335
rect 5344 6261 5390 6301
rect 5344 6227 5350 6261
rect 5384 6227 5390 6261
rect 5344 6187 5390 6227
rect 5344 6153 5350 6187
rect 5384 6153 5390 6187
rect 5344 6113 5390 6153
rect 5344 6079 5350 6113
rect 5384 6079 5390 6113
rect 5344 6039 5390 6079
rect 6091 6430 6156 6472
rect 6091 6396 6100 6430
rect 6134 6396 6156 6430
rect 6091 6354 6156 6396
rect 6091 6320 6100 6354
rect 6134 6320 6156 6354
rect 6091 6278 6156 6320
rect 6091 6272 6100 6278
rect 6134 6272 6156 6278
rect 6143 6220 6156 6272
rect 6091 6202 6156 6220
rect 6091 6199 6100 6202
rect 6134 6199 6156 6202
rect 6143 6147 6156 6199
rect 6091 6126 6156 6147
rect 6143 6074 6156 6126
rect 6327 6228 6379 6555
tri 6379 6535 6399 6555 nw
rect 6327 6164 6379 6176
rect 6327 6106 6379 6112
rect 6481 6521 6490 6555
rect 6524 6521 6533 6555
rect 6481 6482 6533 6521
rect 6481 6448 6490 6482
rect 6524 6448 6533 6482
rect 6481 6409 6533 6448
rect 6481 6375 6490 6409
rect 6524 6375 6533 6409
rect 6481 6335 6533 6375
rect 6481 6301 6490 6335
rect 6524 6301 6533 6335
rect 6481 6261 6533 6301
rect 6481 6227 6490 6261
rect 6524 6227 6533 6261
rect 6481 6187 6533 6227
rect 6481 6153 6490 6187
rect 6524 6153 6533 6187
rect 6481 6113 6533 6153
rect 6091 6053 6156 6074
rect 5344 6005 5350 6039
rect 5384 6005 5390 6039
rect 5344 5965 5390 6005
rect 5344 5931 5350 5965
rect 5384 5931 5390 5965
rect 5344 5891 5390 5931
rect 5344 5857 5350 5891
rect 5384 5857 5390 5891
rect 5344 5817 5390 5857
rect 5344 5783 5350 5817
rect 5384 5783 5390 5817
rect 5344 5743 5390 5783
rect 3076 5666 3122 5705
rect 5344 5709 5350 5743
rect 5384 5709 5390 5743
rect 3076 5632 3082 5666
rect 3116 5632 3122 5666
rect 3076 5593 3122 5632
rect 3262 5625 3488 5677
rect 3540 5625 3552 5677
rect 3604 5625 3824 5677
tri 3688 5595 3718 5625 ne
rect 3718 5595 3824 5625
rect 3076 5559 3082 5593
rect 3116 5559 3122 5593
tri 3718 5592 3721 5595 ne
rect 3076 5520 3122 5559
rect 3076 5486 3082 5520
rect 3116 5486 3122 5520
rect 3076 5447 3122 5486
rect 3076 5413 3082 5447
rect 3116 5413 3122 5447
rect 3076 5374 3122 5413
rect 3076 5340 3082 5374
rect 3116 5340 3122 5374
rect 3076 5339 3122 5340
tri 3122 5339 3127 5344 sw
rect 3076 5333 3127 5339
tri 3127 5333 3133 5339 sw
rect 3076 5310 3133 5333
tri 3133 5310 3156 5333 sw
rect 3076 5301 3533 5310
rect 3585 5301 3597 5310
rect 3076 5267 3154 5301
rect 3188 5267 3240 5301
rect 3274 5267 3326 5301
rect 3360 5267 3412 5301
rect 3446 5267 3498 5301
rect 3532 5267 3533 5301
rect 3076 5258 3533 5267
rect 3585 5258 3597 5267
rect 3649 5258 3655 5310
rect 2796 5217 2842 5255
rect 2796 5183 2802 5217
rect 2836 5183 2842 5217
rect 2796 5145 2842 5183
rect 2796 5111 2802 5145
rect 2836 5111 2842 5145
rect 2796 5079 2842 5111
tri 2842 5079 2847 5084 sw
rect 2796 5076 2847 5079
tri 2847 5076 2850 5079 sw
rect 2796 5073 2850 5076
rect 2796 5039 2802 5073
rect 2836 5050 2850 5073
tri 2850 5050 2876 5076 sw
rect 2836 5041 3533 5050
rect 2836 5039 2899 5041
rect 2796 5007 2899 5039
rect 2933 5007 2977 5041
rect 3011 5007 3056 5041
rect 3090 5007 3135 5041
rect 3169 5007 3214 5041
rect 3248 5007 3293 5041
rect 3327 5007 3372 5041
rect 3406 5007 3451 5041
rect 3485 5007 3530 5041
rect 2796 4998 3533 5007
rect 3585 4998 3597 5050
rect 3649 4998 3655 5050
rect 2791 4894 3533 4903
rect 2791 4860 2803 4894
rect 2837 4860 2876 4894
rect 2910 4860 2949 4894
rect 2983 4860 3022 4894
rect 3056 4860 3095 4894
rect 3129 4860 3168 4894
rect 3202 4860 3241 4894
rect 3275 4860 3314 4894
rect 3348 4860 3387 4894
rect 3421 4860 3461 4894
rect 3495 4860 3533 4894
rect 2791 4851 3533 4860
rect 3585 4851 3597 4903
rect 3649 4851 3655 4903
rect 3120 4730 3126 4782
rect 3178 4773 3220 4782
rect 3272 4773 3314 4782
rect 3366 4773 3591 4782
rect 3178 4739 3215 4773
rect 3272 4739 3298 4773
rect 3366 4739 3381 4773
rect 3415 4739 3463 4773
rect 3497 4739 3545 4773
rect 3579 4739 3591 4773
rect 3178 4730 3220 4739
rect 3272 4730 3314 4739
rect 3366 4730 3591 4739
rect 2985 4633 3037 4645
rect 2985 4599 2994 4633
rect 3028 4599 3037 4633
rect 2985 4561 3037 4599
rect 2985 4527 2994 4561
rect 3028 4527 3037 4561
rect 2985 4489 3037 4527
rect 2985 4455 2994 4489
rect 3028 4455 3037 4489
rect 2985 4391 2994 4403
rect 3028 4391 3037 4403
rect 2985 4311 2994 4339
rect 3028 4311 3037 4339
rect 2985 4273 3037 4311
rect 2985 4239 2994 4273
rect 3028 4239 3037 4273
rect 2985 4201 3037 4239
rect 2985 4167 2994 4201
rect 3028 4167 3037 4201
rect 2985 4129 3037 4167
rect 2985 4095 2994 4129
rect 3028 4095 3037 4129
rect 2985 4057 3037 4095
rect 2985 4023 2994 4057
rect 3028 4023 3037 4057
rect 2985 3985 3037 4023
rect 2985 3951 2994 3985
rect 3028 3951 3037 3985
rect 2985 3913 3037 3951
rect 2985 3879 2994 3913
rect 3028 3879 3037 3913
rect 2985 3841 3037 3879
rect 2985 3807 2994 3841
rect 3028 3807 3037 3841
rect 2985 3769 3037 3807
rect 2985 3735 2994 3769
rect 3028 3735 3037 3769
rect 2985 3697 3037 3735
rect 2985 3663 2994 3697
rect 3028 3663 3037 3697
rect 2985 3625 3037 3663
rect 2985 3591 2994 3625
rect 3028 3591 3037 3625
rect 2985 3553 3037 3591
rect 2985 3519 2994 3553
rect 3028 3519 3037 3553
rect 2985 3481 3037 3519
rect 2985 3447 2994 3481
rect 3028 3447 3037 3481
rect 2985 3409 3037 3447
rect 2985 3375 2994 3409
rect 3028 3375 3037 3409
rect 2985 3337 3037 3375
rect 2985 3303 2994 3337
rect 3028 3303 3037 3337
rect 2985 3291 3037 3303
rect 3141 4633 3193 4645
rect 3141 4599 3150 4633
rect 3184 4599 3193 4633
rect 3141 4561 3193 4599
rect 3141 4527 3150 4561
rect 3184 4527 3193 4561
rect 3141 4489 3193 4527
rect 3141 4455 3150 4489
rect 3184 4455 3193 4489
rect 3141 4417 3193 4455
rect 3141 4383 3150 4417
rect 3184 4383 3193 4417
rect 3141 4345 3193 4383
rect 3141 4311 3150 4345
rect 3184 4311 3193 4345
rect 3141 4273 3193 4311
rect 3141 4241 3150 4273
rect 3184 4241 3193 4273
rect 3141 4177 3150 4189
rect 3184 4177 3193 4189
rect 3141 4095 3150 4125
rect 3184 4095 3193 4125
rect 3141 4057 3193 4095
rect 3141 4023 3150 4057
rect 3184 4023 3193 4057
rect 3141 3985 3193 4023
rect 3141 3951 3150 3985
rect 3184 3951 3193 3985
rect 3141 3913 3193 3951
rect 3141 3879 3150 3913
rect 3184 3879 3193 3913
rect 3141 3841 3193 3879
rect 3141 3807 3150 3841
rect 3184 3807 3193 3841
rect 3141 3769 3193 3807
rect 3141 3735 3150 3769
rect 3184 3735 3193 3769
rect 3141 3697 3193 3735
rect 3141 3663 3150 3697
rect 3184 3663 3193 3697
rect 3141 3625 3193 3663
rect 3141 3591 3150 3625
rect 3184 3591 3193 3625
rect 3141 3553 3193 3591
rect 3141 3519 3150 3553
rect 3184 3519 3193 3553
rect 3141 3481 3193 3519
rect 3141 3447 3150 3481
rect 3184 3447 3193 3481
rect 3141 3409 3193 3447
rect 3141 3375 3150 3409
rect 3184 3375 3193 3409
rect 3141 3337 3193 3375
rect 3141 3303 3150 3337
rect 3184 3303 3193 3337
rect 3141 3291 3193 3303
rect 3297 4633 3349 4645
rect 3297 4599 3306 4633
rect 3340 4599 3349 4633
rect 3297 4561 3349 4599
rect 3297 4527 3306 4561
rect 3340 4527 3349 4561
rect 3297 4489 3349 4527
rect 3297 4455 3306 4489
rect 3340 4455 3349 4489
rect 3297 4391 3306 4403
rect 3340 4391 3349 4403
rect 3297 4311 3306 4339
rect 3340 4311 3349 4339
rect 3297 4273 3349 4311
rect 3297 4239 3306 4273
rect 3340 4239 3349 4273
rect 3297 4201 3349 4239
rect 3297 4167 3306 4201
rect 3340 4167 3349 4201
rect 3297 4129 3349 4167
rect 3297 4095 3306 4129
rect 3340 4095 3349 4129
rect 3297 4057 3349 4095
rect 3297 4023 3306 4057
rect 3340 4023 3349 4057
rect 3297 3985 3349 4023
rect 3297 3951 3306 3985
rect 3340 3951 3349 3985
rect 3297 3913 3349 3951
rect 3297 3879 3306 3913
rect 3340 3879 3349 3913
rect 3297 3841 3349 3879
rect 3297 3807 3306 3841
rect 3340 3807 3349 3841
rect 3297 3769 3349 3807
rect 3297 3735 3306 3769
rect 3340 3735 3349 3769
rect 3297 3697 3349 3735
rect 3297 3663 3306 3697
rect 3340 3663 3349 3697
rect 3297 3625 3349 3663
rect 3297 3591 3306 3625
rect 3340 3591 3349 3625
rect 3297 3553 3349 3591
rect 3297 3519 3306 3553
rect 3340 3519 3349 3553
rect 3297 3481 3349 3519
rect 3297 3447 3306 3481
rect 3340 3447 3349 3481
rect 3297 3409 3349 3447
rect 3297 3375 3306 3409
rect 3340 3375 3349 3409
rect 3297 3337 3349 3375
rect 3297 3303 3306 3337
rect 3340 3303 3349 3337
rect 3297 3291 3349 3303
rect 3453 4633 3505 4645
rect 3453 4599 3462 4633
rect 3496 4599 3505 4633
rect 3453 4561 3505 4599
rect 3453 4527 3462 4561
rect 3496 4527 3505 4561
rect 3453 4489 3505 4527
rect 3453 4455 3462 4489
rect 3496 4455 3505 4489
rect 3453 4417 3505 4455
rect 3453 4383 3462 4417
rect 3496 4383 3505 4417
rect 3453 4345 3505 4383
rect 3453 4311 3462 4345
rect 3496 4311 3505 4345
rect 3453 4273 3505 4311
rect 3453 4241 3462 4273
rect 3496 4241 3505 4273
rect 3453 4177 3462 4189
rect 3496 4177 3505 4189
rect 3453 4095 3462 4125
rect 3496 4095 3505 4125
rect 3453 4057 3505 4095
rect 3453 4023 3462 4057
rect 3496 4023 3505 4057
rect 3453 3985 3505 4023
rect 3453 3951 3462 3985
rect 3496 3951 3505 3985
rect 3453 3913 3505 3951
rect 3453 3879 3462 3913
rect 3496 3879 3505 3913
rect 3453 3841 3505 3879
rect 3453 3807 3462 3841
rect 3496 3807 3505 3841
rect 3453 3769 3505 3807
rect 3453 3735 3462 3769
rect 3496 3735 3505 3769
rect 3453 3697 3505 3735
rect 3453 3663 3462 3697
rect 3496 3663 3505 3697
rect 3453 3625 3505 3663
rect 3453 3591 3462 3625
rect 3496 3591 3505 3625
rect 3453 3553 3505 3591
rect 3453 3519 3462 3553
rect 3496 3519 3505 3553
rect 3453 3481 3505 3519
rect 3453 3447 3462 3481
rect 3496 3447 3505 3481
rect 3453 3409 3505 3447
rect 3453 3375 3462 3409
rect 3496 3375 3505 3409
rect 3453 3337 3505 3375
rect 3453 3303 3462 3337
rect 3496 3303 3505 3337
rect 3453 3291 3505 3303
rect 3609 4633 3661 4645
rect 3609 4599 3618 4633
rect 3652 4599 3661 4633
rect 3609 4561 3661 4599
rect 3609 4527 3618 4561
rect 3652 4527 3661 4561
rect 3609 4489 3661 4527
rect 3609 4455 3618 4489
rect 3652 4455 3661 4489
rect 3609 4391 3618 4403
rect 3652 4391 3661 4403
rect 3609 4311 3618 4339
rect 3652 4311 3661 4339
rect 3609 4273 3661 4311
rect 3609 4239 3618 4273
rect 3652 4239 3661 4273
rect 3609 4201 3661 4239
rect 3609 4167 3618 4201
rect 3652 4167 3661 4201
rect 3609 4129 3661 4167
rect 3609 4095 3618 4129
rect 3652 4095 3661 4129
rect 3721 4241 3824 5595
rect 3991 5476 5284 5676
rect 5344 5669 5390 5709
rect 5543 6033 5595 6039
rect 5543 5969 5595 5981
rect 5543 5748 5595 5917
rect 6143 6001 6156 6053
rect 6091 5979 6156 6001
rect 6143 5927 6156 5979
rect 6091 5905 6156 5927
rect 6143 5853 6156 5905
rect 6091 5831 6156 5853
rect 5543 5742 5775 5748
rect 5543 5708 5657 5742
rect 5691 5708 5729 5742
rect 5763 5708 5775 5742
rect 5543 5702 5775 5708
rect 5344 5635 5350 5669
rect 5384 5635 5390 5669
rect 5344 5595 5390 5635
rect 5344 5561 5350 5595
rect 5384 5561 5390 5595
rect 5344 5521 5390 5561
rect 5344 5487 5350 5521
rect 5384 5487 5390 5521
rect 5344 5447 5390 5487
rect 5809 5459 5855 5787
rect 6143 5779 6156 5831
rect 6481 6079 6490 6113
rect 6524 6079 6533 6113
rect 6481 6039 6533 6079
rect 6481 6005 6490 6039
rect 6524 6005 6533 6039
rect 6481 5965 6533 6005
rect 6481 5931 6490 5965
rect 6524 5931 6533 5965
rect 6481 5891 6533 5931
rect 6481 5857 6490 5891
rect 6524 5857 6533 5891
rect 6481 5817 6533 5857
rect 6481 5783 6490 5817
rect 6524 5783 6533 5817
tri 6085 5487 6091 5493 se
rect 6091 5487 6156 5779
tri 6471 5771 6481 5781 se
rect 6481 5771 6533 5783
tri 6447 5747 6471 5771 se
rect 6471 5747 6533 5771
rect 6396 5743 6533 5747
rect 6396 5709 6490 5743
rect 6524 5709 6533 5743
rect 6396 5701 6533 5709
tri 6447 5698 6450 5701 ne
rect 6450 5698 6533 5701
tri 6450 5669 6479 5698 ne
rect 6479 5669 6533 5698
tri 6479 5667 6481 5669 ne
tri 6077 5479 6085 5487 se
rect 6085 5479 6156 5487
tri 6057 5459 6077 5479 se
rect 6077 5459 6156 5479
rect 5344 5413 5350 5447
rect 5384 5413 5390 5447
rect 5344 5373 5390 5413
tri 5339 5339 5344 5344 se
rect 5344 5339 5350 5373
rect 5384 5339 5390 5373
rect 5647 5427 6156 5459
rect 5647 5375 5653 5427
rect 5705 5375 5717 5427
rect 5769 5375 6034 5427
rect 6086 5375 6098 5427
rect 6150 5375 6156 5427
rect 5647 5366 6156 5375
rect 6481 5635 6490 5669
rect 6524 5635 6533 5669
rect 6481 5595 6533 5635
rect 6481 5561 6490 5595
rect 6524 5561 6533 5595
rect 6481 5521 6533 5561
rect 6481 5487 6490 5521
rect 6524 5487 6533 5521
rect 6481 5447 6533 5487
rect 6481 5413 6490 5447
rect 6524 5413 6533 5447
rect 6481 5373 6533 5413
tri 5390 5339 5395 5344 sw
tri 6476 5339 6481 5344 se
rect 6481 5339 6490 5373
rect 6524 5339 6533 5373
tri 5333 5333 5339 5339 se
rect 5339 5333 5395 5339
tri 5395 5333 5401 5339 sw
tri 6470 5333 6476 5339 se
rect 6476 5333 6533 5339
tri 5310 5310 5333 5333 se
rect 5333 5310 5401 5333
tri 5401 5310 5424 5333 sw
tri 6447 5310 6470 5333 se
rect 6470 5310 6533 5333
rect 3880 5258 3886 5310
rect 3938 5301 3950 5310
rect 4002 5301 6533 5310
rect 4026 5267 4066 5301
rect 4100 5267 4140 5301
rect 4174 5267 4214 5301
rect 4248 5267 4288 5301
rect 4322 5267 4362 5301
rect 4396 5267 4436 5301
rect 4470 5267 4510 5301
rect 4544 5267 4584 5301
rect 4618 5267 4658 5301
rect 4692 5267 4732 5301
rect 4766 5267 4806 5301
rect 4840 5267 4880 5301
rect 4914 5267 4954 5301
rect 4988 5267 5028 5301
rect 5062 5267 5102 5301
rect 5136 5267 5176 5301
rect 5210 5267 5249 5301
rect 5283 5267 5322 5301
rect 5356 5267 5395 5301
rect 5429 5267 5468 5301
rect 5502 5267 5541 5301
rect 5575 5267 5614 5301
rect 5648 5267 5687 5301
rect 5721 5267 5760 5301
rect 5794 5267 5833 5301
rect 5867 5267 5906 5301
rect 5940 5267 5979 5301
rect 6013 5267 6052 5301
rect 6086 5267 6125 5301
rect 6159 5267 6198 5301
rect 6232 5267 6271 5301
rect 6305 5267 6344 5301
rect 6378 5267 6417 5301
rect 6451 5267 6533 5301
rect 3938 5258 3950 5267
rect 4002 5258 6533 5267
rect 6744 7708 6750 7742
rect 6784 7708 6790 7742
rect 6744 7669 6790 7708
rect 6744 7635 6750 7669
rect 6784 7635 6790 7669
rect 6744 7596 6790 7635
rect 6744 7562 6750 7596
rect 6784 7562 6790 7596
rect 6744 7523 6790 7562
rect 6744 7489 6750 7523
rect 6784 7489 6790 7523
rect 6744 7450 6790 7489
rect 6744 7416 6750 7450
rect 6784 7416 6790 7450
rect 6744 7377 6790 7416
rect 6744 7343 6750 7377
rect 6784 7343 6790 7377
rect 6744 7304 6790 7343
rect 6744 7270 6750 7304
rect 6784 7270 6790 7304
rect 6744 7231 6790 7270
rect 6744 7197 6750 7231
rect 6784 7197 6790 7231
rect 6744 7158 6790 7197
rect 6744 7124 6750 7158
rect 6784 7124 6790 7158
rect 6744 7085 6790 7124
rect 6744 7051 6750 7085
rect 6784 7051 6790 7085
rect 6744 7012 6790 7051
rect 6744 6978 6750 7012
rect 6784 6978 6790 7012
rect 6744 6939 6790 6978
rect 6744 6905 6750 6939
rect 6784 6905 6790 6939
rect 6744 6866 6790 6905
rect 6744 6832 6750 6866
rect 6784 6832 6790 6866
rect 6744 6793 6790 6832
rect 7994 8062 8040 8100
rect 7994 8028 8000 8062
rect 8034 8028 8040 8062
rect 7994 7990 8040 8028
rect 7994 7956 8000 7990
rect 8034 7956 8040 7990
rect 7994 7918 8040 7956
rect 7994 7884 8000 7918
rect 8034 7884 8040 7918
rect 7994 7846 8040 7884
rect 7994 7812 8000 7846
rect 8034 7812 8040 7846
rect 7994 7774 8040 7812
rect 7994 7740 8000 7774
rect 8034 7740 8040 7774
rect 7994 7702 8040 7740
rect 7994 7668 8000 7702
rect 8034 7668 8040 7702
rect 7994 7630 8040 7668
rect 7994 7596 8000 7630
rect 8034 7596 8040 7630
rect 7994 7558 8040 7596
rect 7994 7524 8000 7558
rect 8034 7524 8040 7558
rect 7994 7486 8040 7524
rect 7994 7452 8000 7486
rect 8034 7452 8040 7486
rect 7994 7414 8040 7452
rect 7994 7380 8000 7414
rect 8034 7380 8040 7414
rect 7994 7342 8040 7380
rect 7994 7308 8000 7342
rect 8034 7308 8040 7342
rect 7994 7270 8040 7308
rect 7994 7236 8000 7270
rect 8034 7236 8040 7270
rect 7994 7198 8040 7236
rect 7994 7164 8000 7198
rect 8034 7164 8040 7198
rect 7994 7126 8040 7164
rect 7994 7092 8000 7126
rect 8034 7092 8040 7126
rect 7994 7054 8040 7092
rect 7994 7020 8000 7054
rect 8034 7020 8040 7054
rect 7994 6982 8040 7020
rect 7994 6948 8000 6982
rect 8034 6948 8040 6982
rect 7994 6910 8040 6948
rect 7994 6876 8000 6910
rect 8034 6876 8040 6910
rect 7994 6838 8040 6876
rect 7994 6804 8000 6838
rect 8034 6804 8040 6838
rect 6744 6759 6750 6793
rect 6784 6759 6790 6793
rect 6744 6720 6790 6759
rect 6744 6686 6750 6720
rect 6784 6686 6790 6720
rect 6744 6647 6790 6686
rect 6744 6613 6750 6647
rect 6784 6613 6790 6647
rect 6744 6574 6790 6613
rect 6744 6540 6750 6574
rect 6784 6540 6790 6574
rect 6744 6501 6790 6540
rect 6744 6467 6750 6501
rect 6784 6467 6790 6501
rect 6744 6428 6790 6467
rect 6744 6394 6750 6428
rect 6784 6394 6790 6428
rect 6744 6355 6790 6394
rect 6744 6321 6750 6355
rect 6784 6321 6790 6355
rect 6744 6282 6790 6321
rect 6744 6248 6750 6282
rect 6784 6248 6790 6282
rect 6744 6209 6790 6248
rect 6744 6175 6750 6209
rect 6784 6175 6790 6209
rect 6744 6136 6790 6175
rect 6744 6102 6750 6136
rect 6784 6102 6790 6136
rect 6744 6063 6790 6102
rect 6744 6029 6750 6063
rect 6784 6029 6790 6063
rect 6744 5990 6790 6029
rect 6744 5956 6750 5990
rect 6784 5956 6790 5990
rect 6744 5917 6790 5956
rect 6744 5883 6750 5917
rect 6784 5883 6790 5917
rect 6744 5844 6790 5883
rect 6744 5810 6750 5844
rect 6784 5810 6790 5844
rect 6744 5771 6790 5810
rect 6744 5737 6750 5771
rect 6784 5737 6790 5771
rect 6744 5698 6790 5737
rect 6744 5664 6750 5698
rect 6784 5664 6790 5698
rect 6744 5625 6790 5664
rect 6744 5591 6750 5625
rect 6784 5591 6790 5625
rect 6744 5552 6790 5591
rect 6744 5518 6750 5552
rect 6784 5518 6790 5552
rect 6744 5479 6790 5518
rect 6744 5445 6750 5479
rect 6784 5445 6790 5479
rect 6744 5406 6790 5445
rect 6744 5372 6750 5406
rect 6784 5372 6790 5406
rect 6744 5333 6790 5372
rect 6744 5299 6750 5333
rect 6784 5299 6790 5333
rect 6744 5260 6790 5299
rect 6744 5226 6750 5260
rect 6784 5226 6790 5260
rect 6744 5187 6790 5226
rect 6744 5153 6750 5187
rect 6784 5153 6790 5187
rect 6744 5113 6790 5153
tri 6742 5079 6744 5081 se
rect 6744 5079 6750 5113
rect 6784 5079 6790 5113
tri 6739 5076 6742 5079 se
rect 6742 5076 6790 5079
tri 6713 5050 6739 5076 se
rect 6739 5050 6790 5076
rect 3721 4189 3746 4241
rect 3798 4189 3824 4241
rect 3721 4177 3824 4189
rect 3721 4125 3746 4177
rect 3798 4125 3824 4177
rect 3721 4119 3824 4125
rect 3856 4998 3886 5050
rect 3938 5041 3950 5050
rect 4002 5047 4056 5050
tri 4056 5047 4059 5050 sw
tri 6710 5047 6713 5050 se
rect 6713 5047 6790 5050
rect 4002 5041 6790 5047
rect 4025 5007 4064 5041
rect 4098 5007 4137 5041
rect 4171 5007 4210 5041
rect 4244 5007 4283 5041
rect 4317 5007 4356 5041
rect 4390 5007 4429 5041
rect 4463 5007 4502 5041
rect 4536 5007 4575 5041
rect 4609 5007 4648 5041
rect 4682 5007 4721 5041
rect 4755 5007 4794 5041
rect 4828 5007 4867 5041
rect 4901 5007 4940 5041
rect 4974 5007 5013 5041
rect 5047 5007 5086 5041
rect 5120 5007 5159 5041
rect 5193 5007 5232 5041
rect 5266 5007 5305 5041
rect 5339 5007 5378 5041
rect 5412 5007 5451 5041
rect 5485 5007 5524 5041
rect 5558 5007 5597 5041
rect 5631 5007 5670 5041
rect 5704 5007 5742 5041
rect 5776 5007 5814 5041
rect 5848 5007 5874 5041
rect 3938 4998 3950 5007
rect 4002 5001 5874 5007
rect 4002 4998 4058 5001
rect 3856 4969 4058 4998
tri 4058 4969 4090 5001 nw
tri 5839 4969 5871 5001 ne
rect 5871 4989 5874 5001
rect 5926 4989 5942 5041
rect 5994 4989 6010 5041
rect 6064 5007 6078 5041
rect 6136 5007 6146 5041
rect 6208 5007 6214 5041
rect 6280 5007 6318 5041
rect 6352 5007 6390 5041
rect 6424 5007 6462 5041
rect 6496 5007 6534 5041
rect 6568 5007 6606 5041
rect 6640 5007 6678 5041
rect 6712 5007 6790 5041
rect 6062 4989 6078 5007
rect 6130 4989 6146 5007
rect 6198 4989 6214 5007
rect 6266 5001 6790 5007
rect 7784 6793 7875 6799
rect 7784 6741 7792 6793
rect 7844 6741 7875 6793
rect 7784 6729 7875 6741
rect 7784 6677 7792 6729
rect 7844 6677 7875 6729
rect 6266 4989 6269 5001
rect 5871 4971 6269 4989
rect 5871 4969 5874 4971
rect 3856 4932 4056 4969
tri 4056 4967 4058 4969 nw
tri 5871 4967 5873 4969 ne
tri 4056 4932 4058 4934 sw
tri 5871 4932 5873 4934 se
rect 5873 4932 5874 4969
rect 3856 4903 4058 4932
rect 3856 4851 3886 4903
rect 3938 4851 3950 4903
rect 4002 4900 4058 4903
tri 4058 4900 4090 4932 sw
tri 5839 4900 5871 4932 se
rect 5871 4919 5874 4932
rect 5926 4919 5942 4971
rect 5994 4919 6010 4971
rect 6062 4919 6078 4971
rect 6130 4919 6146 4971
rect 6198 4919 6214 4971
rect 6266 4969 6269 4971
tri 6269 4969 6301 5001 nw
rect 6266 4932 6267 4969
tri 6267 4967 6269 4969 nw
tri 6267 4932 6269 4934 sw
rect 6266 4919 6269 4932
rect 5871 4901 6269 4919
rect 5871 4900 5874 4901
rect 4002 4894 5874 4900
rect 5926 4894 5942 4901
rect 5994 4894 6010 4901
rect 6062 4894 6078 4901
rect 6130 4894 6146 4901
rect 6198 4894 6214 4901
rect 6266 4900 6269 4901
tri 6269 4900 6301 4932 sw
rect 6266 4894 6763 4900
rect 4002 4860 4038 4894
rect 4072 4860 4111 4894
rect 4145 4860 4184 4894
rect 4218 4860 4257 4894
rect 4291 4860 4330 4894
rect 4364 4860 4403 4894
rect 4437 4860 4476 4894
rect 4510 4860 4549 4894
rect 4583 4860 4622 4894
rect 4656 4860 4695 4894
rect 4729 4860 4768 4894
rect 4802 4860 4841 4894
rect 4875 4860 4914 4894
rect 4948 4860 4987 4894
rect 5021 4860 5060 4894
rect 5094 4860 5133 4894
rect 5167 4860 5205 4894
rect 5239 4860 5277 4894
rect 5311 4860 5349 4894
rect 5383 4860 5421 4894
rect 5455 4860 5493 4894
rect 5527 4860 5565 4894
rect 5599 4860 5637 4894
rect 5671 4860 5709 4894
rect 5743 4860 5781 4894
rect 5815 4860 5853 4894
rect 5994 4860 5997 4894
rect 6062 4860 6069 4894
rect 6130 4860 6141 4894
rect 6198 4860 6213 4894
rect 6266 4860 6285 4894
rect 6319 4860 6357 4894
rect 6391 4860 6429 4894
rect 6463 4860 6501 4894
rect 6535 4860 6573 4894
rect 6607 4860 6645 4894
rect 6679 4860 6717 4894
rect 6751 4860 6763 4894
rect 4002 4854 5874 4860
rect 4002 4851 4061 4854
rect 3856 4825 4061 4851
tri 4061 4825 4090 4854 nw
tri 5838 4825 5867 4854 ne
rect 5867 4849 5874 4854
rect 5926 4849 5942 4860
rect 5994 4849 6010 4860
rect 6062 4849 6078 4860
rect 6130 4849 6146 4860
rect 6198 4849 6214 4860
rect 6266 4854 6763 4860
rect 6266 4849 6640 4854
rect 5867 4831 6640 4849
rect 5867 4825 5874 4831
rect 3856 4822 4058 4825
tri 4058 4822 4061 4825 nw
tri 5867 4822 5870 4825 ne
rect 5870 4822 5874 4825
rect 3609 4057 3661 4095
rect 3609 4023 3618 4057
rect 3652 4023 3661 4057
rect 3609 3985 3661 4023
rect 3609 3951 3618 3985
rect 3652 3951 3661 3985
rect 3609 3913 3661 3951
rect 3609 3879 3618 3913
rect 3652 3879 3661 3913
rect 3609 3841 3661 3879
rect 3609 3807 3618 3841
rect 3652 3807 3661 3841
rect 3609 3769 3661 3807
rect 3609 3735 3618 3769
rect 3652 3735 3661 3769
rect 3609 3697 3661 3735
rect 3609 3663 3618 3697
rect 3652 3663 3661 3697
rect 3609 3625 3661 3663
rect 3609 3591 3618 3625
rect 3652 3591 3661 3625
rect 3609 3553 3661 3591
rect 3609 3519 3618 3553
rect 3652 3519 3661 3553
rect 3609 3481 3661 3519
rect 3609 3447 3618 3481
rect 3652 3447 3661 3481
rect 3609 3409 3661 3447
rect 3609 3375 3618 3409
rect 3652 3375 3661 3409
rect 3609 3337 3661 3375
rect 3609 3303 3618 3337
rect 3652 3303 3661 3337
rect 3609 3291 3661 3303
rect 3856 3915 4056 4822
tri 4056 4820 4058 4822 nw
tri 5870 4820 5872 4822 ne
rect 5872 4779 5874 4822
rect 5926 4779 5942 4831
rect 5994 4779 6010 4831
rect 6062 4779 6078 4831
rect 6130 4779 6146 4831
rect 6198 4779 6214 4831
rect 6266 4825 6640 4831
tri 6640 4825 6669 4854 nw
rect 6266 4822 6637 4825
tri 6637 4822 6640 4825 nw
rect 6266 4779 6635 4822
tri 6635 4820 6637 4822 nw
rect 5872 4761 6635 4779
rect 5872 4709 5874 4761
rect 5926 4709 5942 4761
rect 5994 4709 6010 4761
rect 6062 4709 6078 4761
rect 6130 4709 6146 4761
rect 6198 4709 6214 4761
rect 6266 4721 6635 4761
rect 6266 4709 6430 4721
rect 5872 4691 6430 4709
rect 4216 4679 4265 4691
rect 4216 4645 4222 4679
rect 4256 4645 4265 4679
rect 4216 4537 4265 4645
rect 4216 4503 4222 4537
rect 4256 4503 4265 4537
rect 4216 4347 4265 4503
rect 5872 4639 5874 4691
rect 5926 4639 5942 4691
rect 5994 4639 6010 4691
rect 6062 4639 6078 4691
rect 6130 4639 6146 4691
rect 6198 4639 6214 4691
rect 6266 4687 6430 4691
rect 6464 4687 6509 4721
rect 6543 4687 6588 4721
rect 6622 4687 6635 4721
rect 6266 4681 6635 4687
rect 6266 4678 6454 4681
tri 6454 4678 6457 4681 nw
rect 6266 4644 6420 4678
tri 6420 4644 6454 4678 nw
rect 6266 4639 6385 4644
rect 5872 4620 6385 4639
rect 5872 4568 5874 4620
rect 5926 4568 5942 4620
rect 5994 4568 6010 4620
rect 6062 4568 6078 4620
rect 6130 4568 6146 4620
rect 6198 4568 6214 4620
rect 6266 4609 6385 4620
tri 6385 4609 6420 4644 nw
rect 6266 4606 6382 4609
tri 6382 4606 6385 4609 nw
rect 6266 4572 6348 4606
tri 6348 4572 6382 4606 nw
rect 6266 4568 6313 4572
rect 5872 4549 6313 4568
rect 5872 4497 5874 4549
rect 5926 4497 5942 4549
rect 5994 4497 6010 4549
rect 6062 4497 6078 4549
rect 6130 4497 6146 4549
rect 6198 4497 6214 4549
rect 6266 4537 6313 4549
tri 6313 4537 6348 4572 nw
rect 6266 4534 6310 4537
tri 6310 4534 6313 4537 nw
rect 6266 4500 6276 4534
tri 6276 4500 6310 4534 nw
rect 6266 4497 6267 4500
rect 5872 4491 6267 4497
tri 6267 4491 6276 4500 nw
rect 6327 4458 6379 4464
rect 4322 4443 4650 4453
rect 4702 4443 4714 4453
rect 4766 4443 5684 4453
rect 4322 4409 4334 4443
rect 4368 4409 4407 4443
rect 4441 4409 4480 4443
rect 4514 4409 4553 4443
rect 4587 4409 4626 4443
rect 4766 4409 4772 4443
rect 4806 4409 4845 4443
rect 4879 4409 4918 4443
rect 4952 4409 4990 4443
rect 5024 4409 5062 4443
rect 5096 4409 5134 4443
rect 5168 4409 5206 4443
rect 5240 4409 5278 4443
rect 5312 4409 5350 4443
rect 5384 4409 5422 4443
rect 5456 4409 5494 4443
rect 5528 4409 5566 4443
rect 5600 4409 5638 4443
rect 5672 4409 5684 4443
rect 4322 4401 4650 4409
rect 4702 4401 4714 4409
rect 4766 4401 5684 4409
rect 6327 4388 6379 4406
rect 4216 4313 4222 4347
rect 4256 4313 4265 4347
rect 4216 4205 4265 4313
rect 4216 4171 4222 4205
rect 4256 4171 4265 4205
rect 4216 4159 4265 4171
rect 5802 4347 5918 4366
rect 5802 4313 5878 4347
rect 5912 4313 5918 4347
rect 5802 4205 5918 4313
rect 5802 4171 5878 4205
rect 5912 4171 5918 4205
rect 5802 4159 5918 4171
rect 6327 4318 6379 4336
rect 7784 4303 7875 6677
rect 6327 4249 6379 4266
rect 6418 4265 6483 4271
rect 6535 4265 6547 4271
rect 6599 4265 6634 4271
rect 6418 4231 6430 4265
rect 6464 4231 6483 4265
rect 6543 4231 6547 4265
rect 6622 4231 6634 4265
rect 6418 4225 6483 4231
rect 6477 4219 6483 4225
rect 6535 4219 6547 4231
rect 6599 4225 6634 4231
rect 7784 4251 7823 4303
rect 7784 4239 7875 4251
rect 6599 4219 6605 4225
rect 6327 4193 6336 4197
rect 6370 4193 6379 4197
rect 6327 4180 6379 4193
tri 5791 4075 5802 4086 se
rect 5802 4075 5905 4159
tri 5771 4055 5791 4075 se
rect 5791 4055 5905 4075
rect 4223 4049 5653 4055
rect 5705 4049 5717 4055
rect 5769 4049 5905 4055
rect 4223 4015 4293 4049
rect 4327 4015 4367 4049
rect 4401 4015 4441 4049
rect 4475 4015 4515 4049
rect 4549 4015 4588 4049
rect 4622 4015 4661 4049
rect 4695 4015 4734 4049
rect 4768 4015 4807 4049
rect 4841 4015 4880 4049
rect 4914 4015 4953 4049
rect 4987 4015 5026 4049
rect 5060 4015 5099 4049
rect 5133 4015 5172 4049
rect 5206 4015 5245 4049
rect 5279 4015 5318 4049
rect 5352 4015 5391 4049
rect 5425 4015 5464 4049
rect 5498 4015 5537 4049
rect 5571 4015 5610 4049
rect 5644 4015 5653 4049
rect 5790 4015 5905 4049
rect 4223 4009 5653 4015
rect 5647 4003 5653 4009
rect 5705 4003 5717 4015
rect 5769 4009 5905 4015
rect 6327 4117 6336 4128
rect 6370 4117 6379 4128
rect 6327 4111 6379 4117
rect 6327 4042 6336 4059
rect 6370 4042 6379 4059
rect 5769 4003 5775 4009
rect 7784 4187 7823 4239
rect 7784 4039 7875 4187
rect 7994 6766 8040 6804
rect 7994 6732 8000 6766
rect 8034 6732 8040 6766
rect 7994 6694 8040 6732
rect 7994 6660 8000 6694
rect 8034 6660 8040 6694
rect 7994 6622 8040 6660
rect 7994 6588 8000 6622
rect 8034 6588 8040 6622
rect 7994 6550 8040 6588
rect 7994 6516 8000 6550
rect 8034 6516 8040 6550
rect 7994 6478 8040 6516
rect 7994 6444 8000 6478
rect 8034 6444 8040 6478
rect 8128 6589 8180 11485
rect 8128 6525 8180 6537
rect 8128 6467 8180 6473
rect 9746 11487 9752 11521
rect 9786 11487 9792 11521
rect 9746 11449 9792 11487
rect 9746 11415 9752 11449
rect 9786 11415 9792 11449
rect 9746 11377 9792 11415
rect 9746 11343 9752 11377
rect 9786 11343 9792 11377
rect 9746 11305 9792 11343
rect 9746 11271 9752 11305
rect 9786 11271 9792 11305
rect 9746 11233 9792 11271
rect 9746 11199 9752 11233
rect 9786 11199 9792 11233
rect 9746 11161 9792 11199
rect 9746 11127 9752 11161
rect 9786 11127 9792 11161
rect 9746 11089 9792 11127
rect 9746 11055 9752 11089
rect 9786 11055 9792 11089
rect 9746 11017 9792 11055
rect 9746 10983 9752 11017
rect 9786 10983 9792 11017
rect 9746 10945 9792 10983
rect 9746 10911 9752 10945
rect 9786 10911 9792 10945
rect 9746 10873 9792 10911
rect 9746 10839 9752 10873
rect 9786 10839 9792 10873
rect 9746 10801 9792 10839
rect 9746 10767 9752 10801
rect 9786 10767 9792 10801
rect 9746 10729 9792 10767
rect 9746 10695 9752 10729
rect 9786 10695 9792 10729
rect 9746 10657 9792 10695
rect 9746 10623 9752 10657
rect 9786 10623 9792 10657
rect 9746 10585 9792 10623
rect 9746 10551 9752 10585
rect 9786 10551 9792 10585
rect 9746 10513 9792 10551
rect 9746 10479 9752 10513
rect 9786 10479 9792 10513
rect 9746 10441 9792 10479
rect 9746 10407 9752 10441
rect 9786 10407 9792 10441
rect 9746 10369 9792 10407
rect 9746 10335 9752 10369
rect 9786 10335 9792 10369
rect 9746 10297 9792 10335
rect 9746 10263 9752 10297
rect 9786 10263 9792 10297
rect 9746 10225 9792 10263
rect 9746 10191 9752 10225
rect 9786 10191 9792 10225
rect 9746 10153 9792 10191
rect 9746 10119 9752 10153
rect 9786 10119 9792 10153
rect 9746 10081 9792 10119
rect 9746 10047 9752 10081
rect 9786 10047 9792 10081
rect 9746 10009 9792 10047
rect 9746 9975 9752 10009
rect 9786 9975 9792 10009
rect 9746 9937 9792 9975
rect 9746 9903 9752 9937
rect 9786 9903 9792 9937
rect 9746 9865 9792 9903
rect 9746 9831 9752 9865
rect 9786 9831 9792 9865
rect 9746 9793 9792 9831
rect 9746 9759 9752 9793
rect 9786 9759 9792 9793
rect 9746 9721 9792 9759
rect 9746 9687 9752 9721
rect 9786 9687 9792 9721
rect 9746 9649 9792 9687
rect 9746 9615 9752 9649
rect 9786 9615 9792 9649
rect 9746 9577 9792 9615
rect 9746 9543 9752 9577
rect 9786 9543 9792 9577
rect 9746 9505 9792 9543
rect 9746 9471 9752 9505
rect 9786 9471 9792 9505
rect 9746 9433 9792 9471
rect 9746 9399 9752 9433
rect 9786 9399 9792 9433
rect 9746 9361 9792 9399
rect 9746 9327 9752 9361
rect 9786 9327 9792 9361
rect 9746 9289 9792 9327
rect 9746 9255 9752 9289
rect 9786 9255 9792 9289
rect 9746 9217 9792 9255
rect 9746 9183 9752 9217
rect 9786 9183 9792 9217
rect 9746 9145 9792 9183
rect 9746 9111 9752 9145
rect 9786 9111 9792 9145
rect 9746 9073 9792 9111
rect 9746 9039 9752 9073
rect 9786 9039 9792 9073
rect 9746 9001 9792 9039
rect 9746 8967 9752 9001
rect 9786 8967 9792 9001
rect 9746 8929 9792 8967
rect 9746 8895 9752 8929
rect 9786 8895 9792 8929
rect 9746 8857 9792 8895
rect 9746 8823 9752 8857
rect 9786 8823 9792 8857
rect 9746 8785 9792 8823
rect 9746 8751 9752 8785
rect 9786 8751 9792 8785
rect 9746 8713 9792 8751
rect 9746 8679 9752 8713
rect 9786 8679 9792 8713
rect 9746 8641 9792 8679
rect 9746 8607 9752 8641
rect 9786 8607 9792 8641
rect 9746 8569 9792 8607
rect 9746 8535 9752 8569
rect 9786 8535 9792 8569
rect 9746 8497 9792 8535
rect 9746 8463 9752 8497
rect 9786 8463 9792 8497
rect 9746 8425 9792 8463
rect 9746 8391 9752 8425
rect 9786 8391 9792 8425
rect 9746 8353 9792 8391
rect 9746 8319 9752 8353
rect 9786 8319 9792 8353
rect 9746 8281 9792 8319
rect 9746 8247 9752 8281
rect 9786 8247 9792 8281
rect 9746 8209 9792 8247
rect 9746 8175 9752 8209
rect 9786 8175 9792 8209
rect 9746 8137 9792 8175
rect 9746 8103 9752 8137
rect 9786 8103 9792 8137
rect 9746 8065 9792 8103
rect 9746 8031 9752 8065
rect 9786 8031 9792 8065
rect 9746 7993 9792 8031
rect 9746 7959 9752 7993
rect 9786 7959 9792 7993
rect 9746 7921 9792 7959
rect 9746 7887 9752 7921
rect 9786 7887 9792 7921
rect 9746 7849 9792 7887
rect 9746 7815 9752 7849
rect 9786 7815 9792 7849
rect 9746 7777 9792 7815
rect 9746 7743 9752 7777
rect 9786 7743 9792 7777
rect 9746 7705 9792 7743
rect 9746 7671 9752 7705
rect 9786 7671 9792 7705
rect 9746 7633 9792 7671
rect 9746 7599 9752 7633
rect 9786 7599 9792 7633
rect 9746 7561 9792 7599
rect 9746 7527 9752 7561
rect 9786 7527 9792 7561
rect 9746 7489 9792 7527
rect 9746 7455 9752 7489
rect 9786 7455 9792 7489
rect 9746 7417 9792 7455
rect 9746 7383 9752 7417
rect 9786 7383 9792 7417
rect 9746 7345 9792 7383
rect 9746 7311 9752 7345
rect 9786 7311 9792 7345
rect 9746 7273 9792 7311
rect 9746 7239 9752 7273
rect 9786 7239 9792 7273
rect 9746 7201 9792 7239
rect 9746 7167 9752 7201
rect 9786 7167 9792 7201
rect 9746 7129 9792 7167
rect 9746 7095 9752 7129
rect 9786 7095 9792 7129
rect 9746 7057 9792 7095
rect 9746 7023 9752 7057
rect 9786 7023 9792 7057
rect 9746 6985 9792 7023
rect 9746 6951 9752 6985
rect 9786 6951 9792 6985
rect 9746 6913 9792 6951
rect 9746 6879 9752 6913
rect 9786 6879 9792 6913
rect 9746 6841 9792 6879
rect 9746 6807 9752 6841
rect 9786 6807 9792 6841
rect 9746 6769 9792 6807
rect 9746 6735 9752 6769
rect 9786 6735 9792 6769
rect 9746 6697 9792 6735
rect 9746 6663 9752 6697
rect 9786 6663 9792 6697
rect 9746 6625 9792 6663
rect 9746 6591 9752 6625
rect 9786 6591 9792 6625
rect 9746 6553 9792 6591
rect 9746 6519 9752 6553
rect 9786 6519 9792 6553
rect 9746 6481 9792 6519
rect 7994 6406 8040 6444
rect 7994 6372 8000 6406
rect 8034 6372 8040 6406
rect 7994 6334 8040 6372
rect 7994 6300 8000 6334
rect 8034 6300 8040 6334
rect 7994 6262 8040 6300
rect 7994 6228 8000 6262
rect 8034 6228 8040 6262
rect 7994 6190 8040 6228
rect 7994 6156 8000 6190
rect 8034 6156 8040 6190
rect 7994 6118 8040 6156
rect 7994 6084 8000 6118
rect 8034 6084 8040 6118
rect 7994 6046 8040 6084
rect 7994 6012 8000 6046
rect 8034 6012 8040 6046
rect 7994 5974 8040 6012
rect 7994 5940 8000 5974
rect 8034 5940 8040 5974
rect 7994 5902 8040 5940
rect 7994 5868 8000 5902
rect 8034 5868 8040 5902
rect 7994 5830 8040 5868
rect 7994 5796 8000 5830
rect 8034 5796 8040 5830
rect 7994 5758 8040 5796
rect 7994 5724 8000 5758
rect 8034 5724 8040 5758
rect 7994 5686 8040 5724
rect 7994 5652 8000 5686
rect 8034 5652 8040 5686
rect 7994 5614 8040 5652
rect 7994 5580 8000 5614
rect 8034 5580 8040 5614
rect 7994 5542 8040 5580
rect 7994 5508 8000 5542
rect 8034 5508 8040 5542
rect 7994 5470 8040 5508
rect 7994 5436 8000 5470
rect 8034 5436 8040 5470
rect 7994 5398 8040 5436
rect 7994 5364 8000 5398
rect 8034 5364 8040 5398
rect 7994 5326 8040 5364
rect 7994 5292 8000 5326
rect 8034 5292 8040 5326
rect 7994 5254 8040 5292
rect 7994 5220 8000 5254
rect 8034 5220 8040 5254
rect 7994 5182 8040 5220
rect 7994 5148 8000 5182
rect 8034 5148 8040 5182
rect 7994 5110 8040 5148
rect 7994 5076 8000 5110
rect 8034 5076 8040 5110
rect 7994 5038 8040 5076
rect 7994 5004 8000 5038
rect 8034 5004 8040 5038
rect 7994 4966 8040 5004
rect 7994 4932 8000 4966
rect 8034 4932 8040 4966
rect 7994 4894 8040 4932
rect 7994 4860 8000 4894
rect 8034 4860 8040 4894
rect 7994 4822 8040 4860
rect 7994 4788 8000 4822
rect 8034 4788 8040 4822
rect 7994 4750 8040 4788
rect 7994 4716 8000 4750
rect 8034 4716 8040 4750
rect 7994 4678 8040 4716
rect 7994 4644 8000 4678
rect 8034 4644 8040 4678
rect 7994 4606 8040 4644
rect 7994 4572 8000 4606
rect 8034 4572 8040 4606
rect 7994 4534 8040 4572
rect 7994 4500 8000 4534
rect 8034 4500 8040 4534
rect 7994 4462 8040 4500
rect 7994 4428 8000 4462
rect 8034 4428 8040 4462
rect 7994 4390 8040 4428
rect 7994 4356 8000 4390
rect 8034 4356 8040 4390
rect 7994 4318 8040 4356
rect 7994 4284 8000 4318
rect 8034 4284 8040 4318
rect 7994 4246 8040 4284
rect 7994 4212 8000 4246
rect 8034 4212 8040 4246
rect 7994 4174 8040 4212
rect 7994 4140 8000 4174
rect 8034 4140 8040 4174
rect 7994 4101 8040 4140
rect 7994 4067 8000 4101
rect 8034 4067 8040 4101
rect 6327 3973 6336 3990
rect 6370 3973 6379 3990
rect 4160 3949 4206 3961
tri 4056 3915 4068 3927 sw
tri 4148 3915 4160 3927 se
rect 4160 3915 4166 3949
rect 4200 3915 4206 3949
rect 3856 3893 4068 3915
tri 4068 3893 4090 3915 sw
tri 4126 3893 4148 3915 se
rect 4148 3893 4206 3915
rect 3856 3809 4206 3893
rect 3856 3775 4166 3809
rect 4200 3775 4206 3809
rect 3856 3763 4206 3775
rect 3856 3745 4188 3763
tri 4188 3745 4206 3763 nw
rect 4973 3955 5101 3967
rect 4973 3921 5022 3955
rect 5056 3921 5101 3955
rect 4973 3880 5101 3921
rect 4973 3846 5022 3880
rect 5056 3846 5101 3880
rect 4973 3805 5101 3846
rect 4973 3771 5022 3805
rect 5056 3771 5101 3805
rect 3856 3736 4179 3745
tri 4179 3736 4188 3745 nw
rect 3856 3702 4145 3736
tri 4145 3702 4179 3736 nw
rect 4973 3703 5101 3771
rect 5872 3955 5879 3967
rect 5872 3921 5878 3955
rect 5872 3915 5879 3921
rect 5931 3915 5962 3967
rect 6014 3915 6045 3967
rect 6097 3915 6127 3967
rect 6179 3915 6209 3967
rect 6261 3915 6268 3967
rect 5872 3891 6268 3915
rect 5872 3882 5879 3891
rect 5872 3848 5878 3882
rect 5872 3839 5879 3848
rect 5931 3839 5962 3891
rect 6014 3839 6045 3891
rect 6097 3839 6127 3891
rect 6179 3839 6209 3891
rect 6261 3839 6268 3891
rect 6327 3889 6336 3921
rect 6370 3889 6379 3921
rect 6327 3877 6379 3889
rect 7994 4028 8040 4067
rect 7994 3994 8000 4028
rect 8034 3994 8040 4028
rect 7994 3955 8040 3994
rect 7994 3921 8000 3955
rect 8034 3921 8040 3955
rect 7994 3882 8040 3921
rect 7994 3848 8000 3882
rect 8034 3848 8040 3882
rect 5872 3817 6268 3839
tri 6268 3817 6299 3848 sw
rect 5872 3815 6299 3817
tri 6299 3815 6301 3817 sw
rect 5872 3809 5879 3815
rect 5872 3775 5878 3809
rect 5872 3763 5879 3775
rect 5931 3763 5962 3815
rect 6014 3763 6045 3815
rect 6097 3763 6127 3815
rect 6179 3763 6209 3815
rect 6261 3809 6673 3815
rect 6261 3775 6430 3809
rect 6464 3775 6509 3809
rect 6543 3775 6588 3809
rect 6622 3775 6673 3809
rect 6261 3763 6673 3775
rect 5872 3749 6673 3763
rect 7994 3809 8040 3848
rect 7994 3775 8000 3809
rect 8034 3775 8040 3809
rect 3856 3673 4116 3702
tri 4116 3673 4145 3702 nw
rect 3856 3663 4106 3673
tri 4106 3663 4116 3673 nw
rect 3856 3651 4094 3663
tri 4094 3651 4106 3663 nw
rect 4973 3651 4979 3703
rect 5031 3651 5043 3703
rect 5095 3651 5101 3703
rect 7994 3736 8040 3775
rect 7994 3702 8000 3736
rect 8034 3702 8040 3736
rect 7994 3663 8040 3702
rect 3856 3629 4072 3651
tri 4072 3629 4094 3651 nw
rect 7994 3629 8000 3663
rect 8034 3629 8040 3663
tri 3849 3191 3856 3198 se
rect 3856 3191 4056 3629
tri 4056 3613 4072 3629 nw
tri 3826 3168 3849 3191 se
rect 3849 3168 4056 3191
tri 3822 3164 3826 3168 se
rect 3826 3164 4056 3168
rect 2672 3158 4056 3164
rect 2672 3124 2684 3158
rect 2718 3124 2760 3158
rect 2794 3124 2836 3158
rect 2870 3124 2912 3158
rect 2946 3124 2988 3158
rect 3022 3124 3064 3158
rect 3098 3124 3140 3158
rect 3174 3124 3216 3158
rect 3250 3124 3292 3158
rect 3326 3124 3368 3158
rect 3402 3124 3444 3158
rect 3478 3124 3520 3158
rect 3554 3124 3595 3158
rect 3629 3124 3670 3158
rect 3704 3124 3745 3158
rect 3779 3124 3820 3158
rect 3854 3124 4056 3158
rect 2672 3118 4056 3124
rect 7994 3590 8040 3629
rect 7994 3556 8000 3590
rect 8034 3556 8040 3590
rect 7994 3517 8040 3556
rect 7994 3483 8000 3517
rect 8034 3483 8040 3517
rect 7994 3444 8040 3483
rect 7994 3410 8000 3444
rect 8034 3410 8040 3444
rect 7994 3371 8040 3410
rect 7994 3337 8000 3371
rect 8034 3337 8040 3371
rect 7994 3298 8040 3337
rect 7994 3264 8000 3298
rect 8034 3264 8040 3298
rect 7994 3225 8040 3264
rect 7994 3191 8000 3225
rect 8034 3191 8040 3225
rect 7994 3152 8040 3191
rect 7994 3118 8000 3152
rect 8034 3118 8040 3152
rect 2481 2879 2599 2918
rect 2481 2845 2487 2879
rect 2521 2845 2559 2879
rect 2593 2845 2599 2879
rect 2481 2806 2599 2845
rect 2481 2772 2487 2806
rect 2521 2772 2559 2806
rect 2593 2772 2599 2806
rect 2481 2733 2599 2772
rect 2481 2699 2487 2733
rect 2521 2699 2559 2733
rect 2593 2699 2599 2733
rect 2481 2660 2599 2699
rect 2481 2626 2487 2660
rect 2521 2626 2559 2660
rect 2593 2626 2599 2660
rect 2481 2587 2599 2626
rect 2481 2553 2487 2587
rect 2521 2553 2559 2587
rect 2593 2553 2599 2587
rect 2481 2514 2599 2553
rect 2481 2480 2487 2514
rect 2521 2480 2559 2514
rect 2593 2480 2599 2514
rect 2481 2441 2599 2480
rect 2481 2407 2487 2441
rect 2521 2407 2559 2441
rect 2593 2407 2599 2441
rect 2481 2368 2599 2407
rect 2481 2334 2487 2368
rect 2521 2334 2559 2368
rect 2593 2334 2599 2368
rect 2481 2295 2599 2334
rect 2481 2261 2487 2295
rect 2521 2261 2559 2295
rect 2593 2261 2599 2295
rect 2481 2222 2599 2261
rect 2481 2188 2487 2222
rect 2521 2188 2559 2222
rect 2593 2188 2599 2222
rect 2481 2149 2599 2188
rect 2481 2115 2487 2149
rect 2521 2115 2559 2149
rect 2593 2115 2599 2149
rect 2481 2076 2599 2115
rect 2481 2042 2487 2076
rect 2521 2042 2559 2076
rect 2593 2042 2599 2076
rect 2481 2003 2599 2042
rect 2481 1969 2487 2003
rect 2521 1969 2559 2003
rect 2593 1969 2599 2003
rect 2481 1930 2599 1969
rect 2481 1896 2487 1930
rect 2521 1896 2559 1930
rect 2593 1896 2599 1930
rect 2481 1857 2599 1896
rect 2481 1823 2487 1857
rect 2521 1823 2559 1857
rect 2593 1823 2599 1857
rect 2481 1784 2599 1823
rect 2481 1750 2487 1784
rect 2521 1750 2559 1784
rect 2593 1750 2599 1784
rect 2481 1711 2599 1750
rect 2481 1677 2487 1711
rect 2521 1677 2559 1711
rect 2593 1677 2599 1711
rect 2481 1638 2599 1677
rect 2481 1604 2487 1638
rect 2521 1604 2559 1638
rect 2593 1604 2599 1638
rect 2481 1565 2599 1604
rect 2481 1531 2487 1565
rect 2521 1531 2559 1565
rect 2593 1531 2599 1565
rect 2481 1492 2599 1531
rect 2481 1458 2487 1492
rect 2521 1458 2559 1492
rect 2593 1458 2599 1492
rect 2481 1419 2599 1458
rect 2481 1385 2487 1419
rect 2521 1385 2559 1419
rect 2593 1385 2599 1419
rect 2481 1346 2599 1385
rect 2481 1312 2487 1346
rect 2521 1312 2559 1346
rect 2593 1312 2599 1346
rect 2481 1273 2599 1312
rect 2481 1239 2487 1273
rect 2521 1239 2559 1273
rect 2593 1239 2599 1273
rect 2481 1200 2599 1239
rect 2481 1166 2487 1200
rect 2521 1166 2559 1200
rect 2593 1166 2599 1200
rect 2481 1127 2599 1166
rect 2481 1093 2487 1127
rect 2521 1093 2559 1127
rect 2593 1093 2599 1127
rect 2481 1054 2599 1093
rect 2481 1020 2487 1054
rect 2521 1020 2559 1054
rect 2593 1020 2599 1054
rect 2481 981 2599 1020
rect 2481 947 2487 981
rect 2521 947 2559 981
rect 2593 947 2599 981
rect 2481 908 2599 947
rect 2481 874 2487 908
rect 2521 874 2559 908
rect 2593 874 2599 908
rect 2481 835 2599 874
rect 2481 801 2487 835
rect 2521 801 2559 835
rect 2593 801 2599 835
rect 2481 762 2599 801
rect 2481 728 2487 762
rect 2521 728 2559 762
rect 2593 728 2599 762
rect 2481 689 2599 728
rect 2481 655 2487 689
rect 2521 655 2559 689
rect 2593 655 2599 689
rect 2481 616 2599 655
rect 2481 582 2487 616
rect 2521 582 2559 616
rect 2593 582 2599 616
rect 2481 543 2599 582
rect 2481 509 2487 543
rect 2521 509 2559 543
rect 2593 509 2599 543
rect 2481 470 2599 509
rect 2481 436 2487 470
rect 2521 436 2559 470
rect 2593 436 2599 470
rect 2481 398 2599 436
rect 7994 3079 8040 3118
rect 7994 3045 8000 3079
rect 8034 3045 8040 3079
rect 7994 3006 8040 3045
rect 7994 2972 8000 3006
rect 8034 2972 8040 3006
rect 7994 2933 8040 2972
rect 7994 2899 8000 2933
rect 8034 2899 8040 2933
rect 7994 2860 8040 2899
rect 7994 2826 8000 2860
rect 8034 2826 8040 2860
rect 7994 2787 8040 2826
rect 7994 2753 8000 2787
rect 8034 2753 8040 2787
rect 7994 2714 8040 2753
rect 7994 2680 8000 2714
rect 8034 2680 8040 2714
rect 7994 2641 8040 2680
rect 7994 2607 8000 2641
rect 8034 2607 8040 2641
rect 7994 2568 8040 2607
rect 7994 2534 8000 2568
rect 8034 2534 8040 2568
rect 7994 2495 8040 2534
rect 7994 2461 8000 2495
rect 8034 2461 8040 2495
rect 7994 2422 8040 2461
rect 7994 2388 8000 2422
rect 8034 2388 8040 2422
rect 7994 2349 8040 2388
rect 7994 2315 8000 2349
rect 8034 2315 8040 2349
rect 7994 2276 8040 2315
rect 7994 2242 8000 2276
rect 8034 2242 8040 2276
rect 7994 2203 8040 2242
rect 7994 2169 8000 2203
rect 8034 2169 8040 2203
rect 7994 2130 8040 2169
rect 7994 2096 8000 2130
rect 8034 2096 8040 2130
rect 7994 2057 8040 2096
rect 7994 2023 8000 2057
rect 8034 2023 8040 2057
rect 7994 1984 8040 2023
rect 7994 1950 8000 1984
rect 8034 1950 8040 1984
rect 7994 1911 8040 1950
rect 7994 1877 8000 1911
rect 8034 1877 8040 1911
rect 7994 1838 8040 1877
rect 7994 1804 8000 1838
rect 8034 1804 8040 1838
rect 7994 1765 8040 1804
rect 7994 1731 8000 1765
rect 8034 1731 8040 1765
rect 7994 1692 8040 1731
rect 7994 1658 8000 1692
rect 8034 1658 8040 1692
rect 7994 1619 8040 1658
rect 7994 1585 8000 1619
rect 8034 1585 8040 1619
rect 7994 1546 8040 1585
rect 7994 1512 8000 1546
rect 8034 1512 8040 1546
rect 7994 1473 8040 1512
rect 7994 1439 8000 1473
rect 8034 1439 8040 1473
rect 7994 1400 8040 1439
rect 7994 1366 8000 1400
rect 8034 1366 8040 1400
rect 7994 1327 8040 1366
rect 7994 1293 8000 1327
rect 8034 1293 8040 1327
rect 7994 1254 8040 1293
rect 7994 1220 8000 1254
rect 8034 1220 8040 1254
rect 7994 1181 8040 1220
rect 7994 1147 8000 1181
rect 8034 1147 8040 1181
rect 7994 1108 8040 1147
rect 7994 1074 8000 1108
rect 8034 1074 8040 1108
rect 7994 1035 8040 1074
rect 7994 1001 8000 1035
rect 8034 1001 8040 1035
rect 7994 962 8040 1001
rect 7994 928 8000 962
rect 8034 928 8040 962
rect 7994 889 8040 928
rect 7994 855 8000 889
rect 8034 855 8040 889
rect 7994 816 8040 855
rect 7994 782 8000 816
rect 8034 782 8040 816
rect 7994 743 8040 782
rect 7994 709 8000 743
rect 8034 709 8040 743
rect 7994 670 8040 709
rect 7994 636 8000 670
rect 8034 636 8040 670
rect 7994 597 8040 636
rect 7994 563 8000 597
rect 8034 563 8040 597
rect 7994 524 8040 563
rect 7994 490 8000 524
rect 8034 490 8040 524
rect 7994 451 8040 490
rect 7994 417 8000 451
rect 8034 417 8040 451
rect 7994 378 8040 417
rect 9746 6447 9752 6481
rect 9786 6447 9792 6481
rect 9746 6409 9792 6447
rect 9746 6375 9752 6409
rect 9786 6375 9792 6409
rect 9746 6337 9792 6375
rect 9746 6303 9752 6337
rect 9786 6303 9792 6337
rect 9746 6265 9792 6303
rect 9746 6231 9752 6265
rect 9786 6231 9792 6265
rect 9746 6193 9792 6231
rect 9746 6159 9752 6193
rect 9786 6159 9792 6193
rect 9746 6121 9792 6159
rect 9746 6087 9752 6121
rect 9786 6087 9792 6121
rect 9746 6049 9792 6087
rect 9746 6015 9752 6049
rect 9786 6015 9792 6049
rect 9746 5977 9792 6015
rect 9746 5943 9752 5977
rect 9786 5943 9792 5977
rect 9746 5905 9792 5943
rect 9746 5871 9752 5905
rect 9786 5871 9792 5905
rect 9746 5833 9792 5871
rect 9746 5799 9752 5833
rect 9786 5799 9792 5833
rect 9746 5761 9792 5799
rect 9746 5727 9752 5761
rect 9786 5727 9792 5761
rect 9746 5689 9792 5727
rect 9746 5655 9752 5689
rect 9786 5655 9792 5689
rect 9746 5617 9792 5655
rect 9746 5583 9752 5617
rect 9786 5583 9792 5617
rect 9746 5545 9792 5583
rect 9746 5511 9752 5545
rect 9786 5511 9792 5545
rect 9746 5473 9792 5511
rect 9746 5439 9752 5473
rect 9786 5439 9792 5473
rect 9746 5401 9792 5439
rect 9746 5367 9752 5401
rect 9786 5367 9792 5401
rect 9746 5329 9792 5367
rect 9746 5295 9752 5329
rect 9786 5295 9792 5329
rect 9746 5257 9792 5295
rect 9746 5223 9752 5257
rect 9786 5223 9792 5257
rect 9746 5185 9792 5223
rect 9746 5151 9752 5185
rect 9786 5151 9792 5185
rect 9746 5113 9792 5151
rect 9746 5079 9752 5113
rect 9786 5079 9792 5113
rect 9746 5041 9792 5079
rect 9746 5007 9752 5041
rect 9786 5007 9792 5041
rect 9746 4969 9792 5007
rect 9746 4935 9752 4969
rect 9786 4935 9792 4969
rect 9746 4897 9792 4935
rect 9746 4863 9752 4897
rect 9786 4863 9792 4897
rect 9746 4825 9792 4863
rect 9746 4791 9752 4825
rect 9786 4791 9792 4825
rect 9746 4753 9792 4791
rect 9746 4719 9752 4753
rect 9786 4719 9792 4753
rect 9746 4681 9792 4719
rect 9746 4647 9752 4681
rect 9786 4647 9792 4681
rect 9746 4609 9792 4647
rect 9746 4575 9752 4609
rect 9786 4575 9792 4609
rect 9746 4537 9792 4575
rect 9746 4503 9752 4537
rect 9786 4503 9792 4537
rect 9746 4465 9792 4503
rect 9746 4431 9752 4465
rect 9786 4431 9792 4465
rect 9746 4393 9792 4431
rect 9746 4359 9752 4393
rect 9786 4359 9792 4393
rect 9746 4321 9792 4359
rect 9746 4287 9752 4321
rect 9786 4287 9792 4321
rect 9746 4249 9792 4287
rect 9746 4215 9752 4249
rect 9786 4215 9792 4249
rect 9746 4177 9792 4215
rect 9746 4143 9752 4177
rect 9786 4143 9792 4177
rect 9746 4105 9792 4143
rect 9746 4071 9752 4105
rect 9786 4071 9792 4105
rect 9746 4033 9792 4071
rect 9746 3999 9752 4033
rect 9786 3999 9792 4033
rect 9746 3961 9792 3999
rect 9746 3927 9752 3961
rect 9786 3927 9792 3961
rect 9746 3889 9792 3927
rect 9746 3855 9752 3889
rect 9786 3855 9792 3889
rect 9746 3817 9792 3855
rect 9746 3783 9752 3817
rect 9786 3783 9792 3817
rect 9746 3745 9792 3783
rect 9746 3711 9752 3745
rect 9786 3711 9792 3745
rect 9746 3673 9792 3711
rect 9746 3639 9752 3673
rect 9786 3639 9792 3673
rect 9746 3601 9792 3639
rect 9746 3567 9752 3601
rect 9786 3567 9792 3601
rect 9746 3529 9792 3567
rect 9746 3495 9752 3529
rect 9786 3495 9792 3529
rect 9746 3457 9792 3495
rect 9746 3423 9752 3457
rect 9786 3423 9792 3457
rect 9746 3385 9792 3423
rect 9746 3351 9752 3385
rect 9786 3351 9792 3385
rect 9746 3313 9792 3351
rect 9746 3279 9752 3313
rect 9786 3279 9792 3313
rect 9746 3241 9792 3279
rect 9746 3207 9752 3241
rect 9786 3207 9792 3241
rect 9746 3168 9792 3207
rect 9746 3134 9752 3168
rect 9786 3134 9792 3168
rect 9746 3095 9792 3134
rect 9746 3061 9752 3095
rect 9786 3061 9792 3095
rect 9746 3022 9792 3061
rect 9746 2988 9752 3022
rect 9786 2988 9792 3022
rect 9746 2949 9792 2988
rect 9746 2915 9752 2949
rect 9786 2915 9792 2949
rect 9746 2876 9792 2915
rect 9746 2842 9752 2876
rect 9786 2842 9792 2876
rect 9746 2803 9792 2842
rect 9746 2769 9752 2803
rect 9786 2769 9792 2803
rect 9746 2730 9792 2769
rect 9746 2696 9752 2730
rect 9786 2696 9792 2730
rect 9746 2657 9792 2696
rect 9746 2623 9752 2657
rect 9786 2623 9792 2657
rect 9746 2584 9792 2623
rect 9746 2550 9752 2584
rect 9786 2550 9792 2584
rect 9746 2511 9792 2550
rect 9746 2477 9752 2511
rect 9786 2477 9792 2511
rect 9746 2438 9792 2477
rect 9746 2404 9752 2438
rect 9786 2404 9792 2438
rect 9746 2365 9792 2404
rect 9746 2331 9752 2365
rect 9786 2331 9792 2365
rect 9746 2292 9792 2331
rect 9746 2258 9752 2292
rect 9786 2258 9792 2292
rect 9746 2219 9792 2258
rect 9746 2185 9752 2219
rect 9786 2185 9792 2219
rect 9746 2146 9792 2185
rect 9746 2112 9752 2146
rect 9786 2112 9792 2146
rect 9746 2073 9792 2112
rect 9746 2039 9752 2073
rect 9786 2039 9792 2073
rect 9746 2000 9792 2039
rect 9746 1966 9752 2000
rect 9786 1966 9792 2000
rect 9746 1927 9792 1966
rect 9746 1893 9752 1927
rect 9786 1893 9792 1927
rect 9746 1854 9792 1893
rect 9746 1820 9752 1854
rect 9786 1820 9792 1854
rect 9746 1781 9792 1820
rect 9746 1747 9752 1781
rect 9786 1747 9792 1781
rect 9746 1708 9792 1747
rect 9746 1674 9752 1708
rect 9786 1674 9792 1708
rect 9746 1635 9792 1674
rect 9746 1601 9752 1635
rect 9786 1601 9792 1635
rect 9746 1562 9792 1601
rect 9746 1528 9752 1562
rect 9786 1528 9792 1562
rect 9746 1489 9792 1528
rect 9746 1455 9752 1489
rect 9786 1455 9792 1489
rect 9746 1416 9792 1455
rect 9746 1382 9752 1416
rect 9786 1382 9792 1416
rect 9746 1343 9792 1382
rect 9746 1309 9752 1343
rect 9786 1309 9792 1343
rect 9746 1270 9792 1309
rect 9746 1236 9752 1270
rect 9786 1236 9792 1270
rect 10131 3514 10249 3520
rect 10183 3462 10197 3514
rect 10131 3450 10249 3462
rect 10183 3398 10197 3450
rect 10131 1399 10249 3398
rect 10131 1293 10137 1399
rect 10243 1293 10249 1399
rect 10131 1260 10249 1293
rect 10710 2487 10716 39777
rect 10822 2487 10828 39817
rect 10710 2448 10828 2487
rect 10710 2414 10716 2448
rect 10750 2414 10788 2448
rect 10822 2414 10828 2448
rect 10710 2375 10828 2414
rect 10710 2341 10716 2375
rect 10750 2341 10788 2375
rect 10822 2341 10828 2375
rect 10710 2302 10828 2341
rect 10710 2268 10716 2302
rect 10750 2268 10788 2302
rect 10822 2268 10828 2302
rect 10710 2229 10828 2268
rect 10710 2195 10716 2229
rect 10750 2195 10788 2229
rect 10822 2195 10828 2229
rect 10710 2156 10828 2195
rect 10710 2122 10716 2156
rect 10750 2122 10788 2156
rect 10822 2122 10828 2156
rect 10710 2083 10828 2122
rect 10710 2049 10716 2083
rect 10750 2049 10788 2083
rect 10822 2049 10828 2083
rect 10710 2010 10828 2049
rect 10710 1976 10716 2010
rect 10750 1976 10788 2010
rect 10822 1976 10828 2010
rect 10710 1937 10828 1976
rect 10710 1903 10716 1937
rect 10750 1903 10788 1937
rect 10822 1903 10828 1937
rect 10710 1864 10828 1903
rect 10710 1830 10716 1864
rect 10750 1830 10788 1864
rect 10822 1830 10828 1864
rect 10710 1791 10828 1830
rect 10710 1757 10716 1791
rect 10750 1757 10788 1791
rect 10822 1757 10828 1791
rect 10710 1718 10828 1757
rect 10710 1684 10716 1718
rect 10750 1684 10788 1718
rect 10822 1684 10828 1718
rect 10710 1645 10828 1684
rect 10710 1611 10716 1645
rect 10750 1611 10788 1645
rect 10822 1611 10828 1645
rect 10710 1572 10828 1611
rect 10710 1538 10716 1572
rect 10750 1538 10788 1572
rect 10822 1538 10828 1572
rect 10710 1499 10828 1538
rect 10710 1465 10716 1499
rect 10750 1465 10788 1499
rect 10822 1465 10828 1499
rect 10710 1426 10828 1465
rect 10710 1392 10716 1426
rect 10750 1392 10788 1426
rect 10822 1392 10828 1426
rect 10710 1353 10828 1392
rect 10710 1319 10716 1353
rect 10750 1319 10788 1353
rect 10822 1319 10828 1353
rect 10710 1280 10828 1319
rect 9746 1197 9792 1236
rect 9746 1163 9752 1197
rect 9786 1163 9792 1197
rect 9746 1124 9792 1163
rect 9746 1090 9752 1124
rect 9786 1090 9792 1124
rect 9746 1051 9792 1090
rect 9746 1017 9752 1051
rect 9786 1017 9792 1051
rect 9746 978 9792 1017
rect 9746 944 9752 978
rect 9786 944 9792 978
rect 9746 905 9792 944
rect 9746 871 9752 905
rect 9786 871 9792 905
rect 9746 832 9792 871
rect 9746 798 9752 832
rect 9786 798 9792 832
rect 9746 759 9792 798
rect 9746 725 9752 759
rect 9786 725 9792 759
rect 9746 686 9792 725
rect 9746 652 9752 686
rect 9786 652 9792 686
rect 9746 613 9792 652
rect 9746 579 9752 613
rect 9786 579 9792 613
rect 9746 540 9792 579
rect 9746 506 9752 540
rect 9786 506 9792 540
rect 9746 467 9792 506
rect 9746 433 9752 467
rect 9786 433 9792 467
rect 9746 401 9792 433
rect 10710 1246 10716 1280
rect 10750 1246 10788 1280
rect 10822 1246 10828 1280
rect 10710 1207 10828 1246
rect 10710 1173 10716 1207
rect 10750 1173 10788 1207
rect 10822 1173 10828 1207
rect 10710 1134 10828 1173
rect 10710 1100 10716 1134
rect 10750 1100 10788 1134
rect 10822 1100 10828 1134
rect 10710 1061 10828 1100
rect 10710 1027 10716 1061
rect 10750 1027 10788 1061
rect 10822 1027 10828 1061
rect 10710 988 10828 1027
rect 10710 954 10716 988
rect 10750 954 10788 988
rect 10822 954 10828 988
rect 10710 915 10828 954
rect 10710 881 10716 915
rect 10750 881 10788 915
rect 10822 881 10828 915
rect 10710 842 10828 881
rect 10710 808 10716 842
rect 10750 808 10788 842
rect 10822 808 10828 842
rect 10710 769 10828 808
rect 10710 735 10716 769
rect 10750 735 10788 769
rect 10822 735 10828 769
rect 10710 696 10828 735
rect 10710 662 10716 696
rect 10750 662 10788 696
rect 10822 662 10828 696
rect 10710 623 10828 662
rect 10710 589 10716 623
rect 10750 589 10788 623
rect 10822 589 10828 623
rect 10710 550 10828 589
rect 10710 516 10716 550
rect 10750 516 10788 550
rect 10822 516 10828 550
rect 10710 477 10828 516
rect 10710 443 10716 477
rect 10750 443 10788 477
rect 10822 443 10828 477
rect 10710 404 10828 443
rect 7994 344 8000 378
rect 8034 344 8040 378
rect 7994 305 8040 344
rect 7994 271 8000 305
rect 8034 271 8040 305
rect 7994 232 8040 271
rect 7994 198 8000 232
rect 8034 198 8040 232
rect 7994 159 8040 198
rect 7994 125 8000 159
rect 8034 125 8040 159
rect 7994 86 8040 125
rect 7994 52 8000 86
rect 8034 52 8040 86
rect 7994 40 8040 52
rect 10710 370 10716 404
rect 10750 370 10788 404
rect 10822 370 10828 404
rect 10710 331 10828 370
rect 10710 297 10716 331
rect 10750 297 10788 331
rect 10822 297 10828 331
rect 10710 258 10828 297
rect 10710 224 10716 258
rect 10750 224 10788 258
rect 10822 224 10828 258
rect 10710 185 10828 224
rect 10710 151 10716 185
rect 10750 151 10788 185
rect 10822 151 10828 185
rect 10710 112 10828 151
rect 10710 78 10716 112
rect 10750 78 10788 112
rect 10822 78 10828 112
rect 10710 40 10828 78
<< via1 >>
rect 2305 39713 2357 39719
rect 2305 39679 2310 39713
rect 2310 39679 2344 39713
rect 2344 39679 2357 39713
rect 2305 39667 2357 39679
rect 2369 39713 2421 39719
rect 2369 39679 2382 39713
rect 2382 39679 2416 39713
rect 2416 39679 2421 39713
rect 2369 39667 2421 39679
rect 2305 39640 2357 39649
rect 2305 39606 2310 39640
rect 2310 39606 2344 39640
rect 2344 39606 2357 39640
rect 2305 39597 2357 39606
rect 2369 39640 2421 39649
rect 2369 39606 2382 39640
rect 2382 39606 2416 39640
rect 2416 39606 2421 39640
rect 2369 39597 2421 39606
rect 2305 39567 2357 39579
rect 2305 39533 2310 39567
rect 2310 39533 2344 39567
rect 2344 39533 2357 39567
rect 2305 39527 2357 39533
rect 2369 39567 2421 39579
rect 2369 39533 2382 39567
rect 2382 39533 2416 39567
rect 2416 39533 2421 39567
rect 2369 39527 2421 39533
rect 656 26306 708 26358
rect 656 26242 708 26294
rect 656 6471 708 6523
rect 656 6407 708 6459
rect 656 4800 708 4852
rect 656 4736 708 4788
rect 512 4339 628 4455
rect 8107 39713 8159 39719
rect 8107 39679 8112 39713
rect 8112 39679 8146 39713
rect 8146 39679 8159 39713
rect 8107 39667 8159 39679
rect 8171 39713 8223 39719
rect 8171 39679 8184 39713
rect 8184 39679 8218 39713
rect 8218 39679 8223 39713
rect 8171 39667 8223 39679
rect 8107 39640 8159 39649
rect 8107 39606 8112 39640
rect 8112 39606 8146 39640
rect 8146 39606 8159 39640
rect 8107 39597 8159 39606
rect 8171 39640 8223 39649
rect 8171 39606 8184 39640
rect 8184 39606 8218 39640
rect 8218 39606 8223 39640
rect 8171 39597 8223 39606
rect 8107 39567 8159 39579
rect 8107 39533 8112 39567
rect 8112 39533 8146 39567
rect 8146 39533 8159 39567
rect 8107 39527 8159 39533
rect 8171 39567 8223 39579
rect 8171 39533 8184 39567
rect 8184 39533 8218 39567
rect 8218 39533 8223 39567
rect 8171 39527 8223 39533
rect 9559 39713 9611 39719
rect 9559 39679 9564 39713
rect 9564 39679 9598 39713
rect 9598 39679 9611 39713
rect 9559 39667 9611 39679
rect 9623 39713 9675 39719
rect 9623 39679 9636 39713
rect 9636 39679 9670 39713
rect 9670 39679 9675 39713
rect 9623 39667 9675 39679
rect 9559 39640 9611 39649
rect 9559 39606 9564 39640
rect 9564 39606 9598 39640
rect 9598 39606 9611 39640
rect 9559 39597 9611 39606
rect 9623 39640 9675 39649
rect 9623 39606 9636 39640
rect 9636 39606 9670 39640
rect 9670 39606 9675 39640
rect 9623 39597 9675 39606
rect 9559 39567 9611 39579
rect 9559 39533 9564 39567
rect 9564 39533 9598 39567
rect 9598 39533 9611 39567
rect 9559 39527 9611 39533
rect 9623 39567 9675 39579
rect 9623 39533 9636 39567
rect 9636 39533 9670 39567
rect 9670 39533 9675 39567
rect 9623 39527 9675 39533
rect 5604 39218 5656 39270
rect 5604 39154 5656 39206
rect 5604 39090 5656 39142
rect 5604 39026 5656 39078
rect 5604 38962 5656 39014
rect 5604 38898 5656 38950
rect 5604 38834 5656 38886
rect 5604 38770 5656 38822
rect 5604 38706 5656 38758
rect 5604 38642 5656 38694
rect 5604 38578 5656 38630
rect 5604 38514 5656 38566
rect 5604 38450 5656 38502
rect 5604 38386 5656 38438
rect 5604 38322 5656 38374
rect 5604 38258 5656 38310
rect 5604 38194 5656 38246
rect 5604 38130 5656 38182
rect 5604 38066 5656 38118
rect 5604 38002 5656 38054
rect 5604 37938 5656 37990
rect 5604 37874 5656 37926
rect 5604 37810 5656 37862
rect 5604 37746 5656 37798
rect 5604 37682 5656 37734
rect 5604 37618 5656 37670
rect 5604 37554 5656 37606
rect 5604 37490 5656 37542
rect 5604 37426 5656 37478
rect 5604 37362 5656 37414
rect 5604 37298 5656 37350
rect 5604 37234 5656 37286
rect 5604 37170 5656 37222
rect 5604 37106 5656 37158
rect 5604 37042 5656 37094
rect 5604 36978 5656 37030
rect 5604 36914 5656 36966
rect 5604 36850 5656 36902
rect 5604 36786 5656 36838
rect 5604 36722 5656 36774
rect 5604 36658 5656 36710
rect 5604 36594 5656 36646
rect 5604 36530 5656 36582
rect 5604 36466 5656 36518
rect 5604 36402 5656 36454
rect 5604 36338 5656 36390
rect 5604 36274 5656 36326
rect 5604 36210 5656 36262
rect 5604 36146 5656 36198
rect 5604 36082 5656 36134
rect 5604 36018 5656 36070
rect 5604 35954 5656 36006
rect 5604 35890 5656 35942
rect 5604 35826 5656 35878
rect 5604 35762 5656 35814
rect 5604 35698 5656 35750
rect 5604 35634 5656 35686
rect 5604 35570 5656 35622
rect 5604 35506 5656 35558
rect 5604 35442 5656 35494
rect 5604 35378 5656 35430
rect 5604 35314 5656 35366
rect 5604 35250 5656 35302
rect 5604 35186 5656 35238
rect 5604 35122 5656 35174
rect 5604 35058 5656 35110
rect 5604 34994 5656 35046
rect 5604 34930 5656 34982
rect 7526 34970 7532 35001
rect 7532 34970 7566 35001
rect 7566 34970 7578 35001
rect 7526 34949 7578 34970
rect 5604 34866 5656 34918
rect 7526 34931 7578 34937
rect 7526 34897 7532 34931
rect 7532 34897 7566 34931
rect 7566 34897 7578 34931
rect 7526 34885 7578 34897
rect 10554 39713 10606 39719
rect 10554 39679 10559 39713
rect 10559 39679 10593 39713
rect 10593 39679 10606 39713
rect 10554 39667 10606 39679
rect 10618 39713 10670 39719
rect 10618 39679 10631 39713
rect 10631 39679 10665 39713
rect 10665 39679 10670 39713
rect 10618 39667 10670 39679
rect 10554 39640 10606 39649
rect 10554 39606 10559 39640
rect 10559 39606 10593 39640
rect 10593 39606 10606 39640
rect 10554 39597 10606 39606
rect 10618 39640 10670 39649
rect 10618 39606 10631 39640
rect 10631 39606 10665 39640
rect 10665 39606 10670 39640
rect 10618 39597 10670 39606
rect 10554 39567 10606 39579
rect 10554 39533 10559 39567
rect 10559 39533 10593 39567
rect 10593 39533 10606 39567
rect 10554 39527 10606 39533
rect 10618 39567 10670 39579
rect 10618 39533 10631 39567
rect 10631 39533 10665 39567
rect 10665 39533 10670 39567
rect 10618 39527 10670 39533
rect 5604 34802 5656 34854
rect 5604 34738 5656 34790
rect 5604 34674 5656 34726
rect 5604 34610 5656 34662
rect 5604 34546 5656 34598
rect 5604 34482 5656 34534
rect 5604 34418 5656 34470
rect 5604 34354 5656 34406
rect 5604 34290 5656 34342
rect 5604 34226 5656 34278
rect 5604 34162 5656 34214
rect 5604 34098 5656 34150
rect 5604 34034 5656 34086
rect 5604 33970 5656 34022
rect 5604 33906 5656 33958
rect 5604 33842 5656 33894
rect 5604 33778 5656 33830
rect 5604 33714 5656 33766
rect 5604 33650 5656 33702
rect 5604 33586 5656 33638
rect 5604 33522 5656 33574
rect 5604 33458 5656 33510
rect 5604 33394 5656 33446
rect 5604 33330 5656 33382
rect 5604 33266 5656 33318
rect 5604 33202 5656 33254
rect 5604 33138 5656 33190
rect 5604 33074 5656 33126
rect 5604 33010 5656 33062
rect 5604 32946 5656 32998
rect 5604 32882 5656 32934
rect 5604 32818 5656 32870
rect 5604 32754 5656 32806
rect 5604 32690 5656 32742
rect 5604 32625 5656 32677
rect 5604 32560 5656 32612
rect 5604 32495 5656 32547
rect 5604 32430 5656 32482
rect 5604 32365 5656 32417
rect 5604 32300 5656 32352
rect 5604 32235 5656 32287
rect 5604 32170 5656 32222
rect 5604 32105 5656 32157
rect 5604 32040 5656 32092
rect 5604 31975 5656 32027
rect 5604 31910 5656 31962
rect 5604 31845 5656 31897
rect 5604 31780 5656 31832
rect 5604 31715 5656 31767
rect 7526 31747 7578 31753
rect 5604 31650 5656 31702
rect 7526 31713 7532 31747
rect 7532 31713 7566 31747
rect 7566 31713 7578 31747
rect 7526 31701 7578 31713
rect 7526 31675 7578 31689
rect 5604 31585 5656 31637
rect 5604 31520 5656 31572
rect 5604 31455 5656 31507
rect 5604 31390 5656 31442
rect 5604 31325 5656 31377
rect 7526 31641 7532 31675
rect 7532 31641 7566 31675
rect 7566 31641 7578 31675
rect 7526 31637 7578 31641
rect 8784 34949 8836 35001
rect 8784 34885 8836 34937
rect 5604 31260 5656 31312
rect 5604 31195 5656 31247
rect 5604 31130 5656 31182
rect 5604 31065 5656 31117
rect 5604 31000 5656 31052
rect 5604 30935 5656 30987
rect 5604 30870 5656 30922
rect 5604 30805 5656 30857
rect 5604 30740 5656 30792
rect 5604 30675 5656 30727
rect 5604 30610 5656 30662
rect 5604 30545 5656 30597
rect 5604 30480 5656 30532
rect 5604 30415 5656 30467
rect 5604 30350 5656 30402
rect 5714 29859 5766 29911
rect 5801 29859 5853 29911
rect 5714 29783 5766 29835
rect 5801 29783 5853 29835
rect 7583 29842 7635 29894
rect 7647 29842 7699 29894
rect 7503 29762 7555 29814
rect 7567 29762 7619 29814
rect 7322 29647 7374 29699
rect 7386 29647 7438 29699
rect 6739 27228 6791 27280
rect 6806 27228 6858 27280
rect 6873 27228 6925 27280
rect 6940 27228 6992 27280
rect 7007 27228 7059 27280
rect 7074 27228 7126 27280
rect 7141 27228 7193 27280
rect 7208 27228 7260 27280
rect 7275 27228 7327 27280
rect 7342 27228 7394 27280
rect 7409 27228 7461 27280
rect 7476 27228 7528 27280
rect 7543 27228 7595 27280
rect 7610 27228 7662 27280
rect 7676 27228 7728 27280
rect 7742 27228 7794 27280
rect 4669 27086 4721 27138
rect 4736 27086 4788 27138
rect 4803 27086 4855 27138
rect 4870 27086 4922 27138
rect 4937 27086 4989 27138
rect 5004 27086 5056 27138
rect 5071 27086 5123 27138
rect 5138 27086 5190 27138
rect 5205 27086 5257 27138
rect 5272 27086 5324 27138
rect 5339 27086 5391 27138
rect 5406 27086 5458 27138
rect 5473 27086 5525 27138
rect 5539 27086 5591 27138
rect 5605 27086 5657 27138
rect 4669 27008 4721 27060
rect 4736 27008 4788 27060
rect 4803 27008 4855 27060
rect 4870 27008 4922 27060
rect 4937 27008 4989 27060
rect 5004 27008 5056 27060
rect 5071 27008 5123 27060
rect 5138 27008 5190 27060
rect 5205 27008 5257 27060
rect 5272 27008 5324 27060
rect 5339 27008 5391 27060
rect 5406 27008 5458 27060
rect 5473 27008 5525 27060
rect 5539 27008 5591 27060
rect 5605 27008 5657 27060
rect 6479 27118 6595 27124
rect 6479 27012 6485 27118
rect 6485 27012 6591 27118
rect 6591 27012 6595 27118
rect 6479 27008 6595 27012
rect 6083 22079 6135 22131
rect 6147 22079 6199 22131
rect 6675 21374 6727 21426
rect 6739 21374 6791 21426
rect 6592 21294 6644 21346
rect 6656 21294 6708 21346
rect 6423 21214 6475 21266
rect 6487 21214 6539 21266
rect 8068 31701 8120 31753
rect 8068 31637 8120 31689
rect 9094 29842 9146 29894
rect 9158 29842 9210 29894
rect 9008 29756 9060 29808
rect 8784 27078 8836 27130
rect 8784 27014 8836 27066
rect 8784 26306 8836 26358
rect 8784 26242 8836 26294
rect 8928 29641 8980 29693
rect 8928 29577 8980 29629
rect 8809 21374 8861 21426
rect 8873 21374 8925 21426
rect 9008 29692 9060 29744
rect 9008 21364 9060 21416
rect 9008 21300 9060 21352
rect 9094 21214 9146 21266
rect 9158 21214 9210 21266
rect 4728 7689 4756 7710
rect 4756 7689 4780 7710
rect 4800 7689 4828 7710
rect 4828 7689 4852 7710
rect 4871 7689 4900 7710
rect 4900 7689 4923 7710
rect 4942 7689 4972 7710
rect 4972 7689 4994 7710
rect 5013 7689 5044 7710
rect 5044 7689 5065 7710
rect 5084 7689 5116 7710
rect 5116 7689 5136 7710
rect 5155 7689 5188 7710
rect 5188 7689 5207 7710
rect 5226 7689 5260 7710
rect 5260 7689 5278 7710
rect 5649 7689 5654 7719
rect 5654 7689 5692 7719
rect 5692 7689 5701 7719
rect 5723 7689 5726 7719
rect 5726 7689 5764 7719
rect 5764 7689 5775 7719
rect 5797 7689 5798 7719
rect 5798 7689 5836 7719
rect 5836 7689 5849 7719
rect 6197 7689 6199 7700
rect 6199 7689 6233 7700
rect 6233 7689 6249 7700
rect 4728 7658 4780 7689
rect 4800 7658 4852 7689
rect 4871 7658 4923 7689
rect 4942 7658 4994 7689
rect 5013 7658 5065 7689
rect 5084 7658 5136 7689
rect 5155 7658 5207 7689
rect 5226 7658 5278 7689
rect 4728 7584 4780 7636
rect 4800 7584 4852 7636
rect 4871 7584 4923 7636
rect 4942 7584 4994 7636
rect 5013 7584 5065 7636
rect 5084 7584 5136 7636
rect 5155 7584 5207 7636
rect 5226 7584 5278 7636
rect 5649 7667 5701 7689
rect 5723 7667 5775 7689
rect 5797 7667 5849 7689
rect 4728 7510 4780 7562
rect 4800 7510 4852 7562
rect 4871 7510 4923 7562
rect 4942 7510 4994 7562
rect 5013 7510 5065 7562
rect 5084 7510 5136 7562
rect 5155 7510 5207 7562
rect 5226 7510 5278 7562
rect 4728 7436 4780 7488
rect 4800 7436 4852 7488
rect 4871 7436 4923 7488
rect 4942 7436 4994 7488
rect 5013 7436 5065 7488
rect 5084 7436 5136 7488
rect 5155 7436 5207 7488
rect 5226 7436 5278 7488
rect 4728 7362 4780 7414
rect 4800 7362 4852 7414
rect 4871 7362 4923 7414
rect 4942 7362 4994 7414
rect 5013 7362 5065 7414
rect 5084 7362 5136 7414
rect 5155 7362 5207 7414
rect 5226 7362 5278 7414
rect 4728 7288 4780 7340
rect 4800 7288 4852 7340
rect 4871 7288 4923 7340
rect 4942 7288 4994 7340
rect 5013 7288 5065 7340
rect 5084 7288 5136 7340
rect 5155 7288 5207 7340
rect 5226 7288 5278 7340
rect 5649 7592 5701 7644
rect 5723 7592 5775 7644
rect 5797 7592 5849 7644
rect 5649 7517 5701 7569
rect 5723 7517 5775 7569
rect 5797 7517 5849 7569
rect 5649 7442 5701 7494
rect 5723 7442 5775 7494
rect 5797 7442 5849 7494
rect 5649 7367 5701 7419
rect 5723 7367 5775 7419
rect 5797 7367 5849 7419
rect 5649 7292 5701 7344
rect 5723 7292 5775 7344
rect 5797 7292 5849 7344
rect 6197 7648 6249 7689
rect 6271 7689 6272 7700
rect 6272 7689 6306 7700
rect 6306 7689 6323 7700
rect 6271 7648 6323 7689
rect 6345 7689 6379 7700
rect 6379 7689 6397 7700
rect 6345 7648 6397 7689
rect 6481 7671 6533 7723
rect 6197 7577 6249 7629
rect 6271 7577 6323 7629
rect 6345 7577 6397 7629
rect 6481 7616 6490 7648
rect 6490 7616 6524 7648
rect 6524 7616 6533 7648
rect 6481 7596 6533 7616
rect 6197 7506 6249 7558
rect 6271 7506 6323 7558
rect 6345 7506 6397 7558
rect 6481 7543 6490 7573
rect 6490 7543 6524 7573
rect 6524 7543 6533 7573
rect 6481 7521 6533 7543
rect 6197 7435 6249 7487
rect 6271 7435 6323 7487
rect 6345 7435 6397 7487
rect 6481 7470 6490 7497
rect 6490 7470 6524 7497
rect 6524 7470 6533 7497
rect 6481 7445 6533 7470
rect 6197 7364 6249 7416
rect 6271 7364 6323 7416
rect 6345 7364 6397 7416
rect 6481 7397 6490 7421
rect 6490 7397 6524 7421
rect 6524 7397 6533 7421
rect 6481 7369 6533 7397
rect 6197 7293 6249 7345
rect 6271 7293 6323 7345
rect 6345 7293 6397 7345
rect 6481 7324 6490 7345
rect 6490 7324 6524 7345
rect 6524 7324 6533 7345
rect 6481 7293 6533 7324
rect 3847 6493 3856 6523
rect 3856 6493 3890 6523
rect 3890 6493 3899 6523
rect 3847 6471 3899 6493
rect 3847 6452 3899 6459
rect 3847 6418 3856 6452
rect 3856 6418 3890 6452
rect 3890 6418 3899 6452
rect 3847 6407 3899 6418
rect 4577 6493 4586 6523
rect 4586 6493 4620 6523
rect 4620 6493 4629 6523
rect 4577 6471 4629 6493
rect 4577 6452 4629 6459
rect 4577 6418 4586 6452
rect 4586 6418 4620 6452
rect 4620 6418 4629 6452
rect 4577 6407 4629 6418
rect 6269 6671 6321 6723
rect 6369 6671 6421 6723
rect 5809 6537 5861 6589
rect 5809 6473 5861 6525
rect 6091 6244 6100 6272
rect 6100 6244 6134 6272
rect 6134 6244 6143 6272
rect 6091 6220 6143 6244
rect 6091 6168 6100 6199
rect 6100 6168 6134 6199
rect 6134 6168 6143 6199
rect 6091 6147 6143 6168
rect 6091 6092 6100 6126
rect 6100 6092 6134 6126
rect 6134 6092 6143 6126
rect 6091 6074 6143 6092
rect 6327 6176 6379 6228
rect 6327 6112 6379 6164
rect 6091 6050 6143 6053
rect 3488 5625 3540 5677
rect 3552 5625 3604 5677
rect 3533 5301 3585 5310
rect 3597 5301 3649 5310
rect 3533 5267 3583 5301
rect 3583 5267 3585 5301
rect 3597 5267 3617 5301
rect 3617 5267 3649 5301
rect 3533 5258 3585 5267
rect 3597 5258 3649 5267
rect 3533 5041 3585 5050
rect 3533 5007 3564 5041
rect 3564 5007 3585 5041
rect 3533 4998 3585 5007
rect 3597 5041 3649 5050
rect 3597 5007 3609 5041
rect 3609 5007 3643 5041
rect 3643 5007 3649 5041
rect 3597 4998 3649 5007
rect 3533 4894 3585 4903
rect 3533 4860 3535 4894
rect 3535 4860 3569 4894
rect 3569 4860 3585 4894
rect 3533 4851 3585 4860
rect 3597 4894 3649 4903
rect 3597 4860 3609 4894
rect 3609 4860 3643 4894
rect 3643 4860 3649 4894
rect 3597 4851 3649 4860
rect 3126 4773 3178 4782
rect 3220 4773 3272 4782
rect 3314 4773 3366 4782
rect 3126 4739 3132 4773
rect 3132 4739 3166 4773
rect 3166 4739 3178 4773
rect 3220 4739 3249 4773
rect 3249 4739 3272 4773
rect 3314 4739 3332 4773
rect 3332 4739 3366 4773
rect 3126 4730 3178 4739
rect 3220 4730 3272 4739
rect 3314 4730 3366 4739
rect 2985 4417 3037 4455
rect 2985 4403 2994 4417
rect 2994 4403 3028 4417
rect 3028 4403 3037 4417
rect 2985 4383 2994 4391
rect 2994 4383 3028 4391
rect 3028 4383 3037 4391
rect 2985 4345 3037 4383
rect 2985 4339 2994 4345
rect 2994 4339 3028 4345
rect 3028 4339 3037 4345
rect 3141 4239 3150 4241
rect 3150 4239 3184 4241
rect 3184 4239 3193 4241
rect 3141 4201 3193 4239
rect 3141 4189 3150 4201
rect 3150 4189 3184 4201
rect 3184 4189 3193 4201
rect 3141 4167 3150 4177
rect 3150 4167 3184 4177
rect 3184 4167 3193 4177
rect 3141 4129 3193 4167
rect 3141 4125 3150 4129
rect 3150 4125 3184 4129
rect 3184 4125 3193 4129
rect 3297 4417 3349 4455
rect 3297 4403 3306 4417
rect 3306 4403 3340 4417
rect 3340 4403 3349 4417
rect 3297 4383 3306 4391
rect 3306 4383 3340 4391
rect 3340 4383 3349 4391
rect 3297 4345 3349 4383
rect 3297 4339 3306 4345
rect 3306 4339 3340 4345
rect 3340 4339 3349 4345
rect 3453 4239 3462 4241
rect 3462 4239 3496 4241
rect 3496 4239 3505 4241
rect 3453 4201 3505 4239
rect 3453 4189 3462 4201
rect 3462 4189 3496 4201
rect 3496 4189 3505 4201
rect 3453 4167 3462 4177
rect 3462 4167 3496 4177
rect 3496 4167 3505 4177
rect 3453 4129 3505 4167
rect 3453 4125 3462 4129
rect 3462 4125 3496 4129
rect 3496 4125 3505 4129
rect 3609 4417 3661 4455
rect 3609 4403 3618 4417
rect 3618 4403 3652 4417
rect 3652 4403 3661 4417
rect 3609 4383 3618 4391
rect 3618 4383 3652 4391
rect 3652 4383 3661 4391
rect 3609 4345 3661 4383
rect 3609 4339 3618 4345
rect 3618 4339 3652 4345
rect 3652 4339 3661 4345
rect 5543 5981 5595 6033
rect 5543 5917 5595 5969
rect 6091 6016 6100 6050
rect 6100 6016 6134 6050
rect 6134 6016 6143 6050
rect 6091 6001 6143 6016
rect 6091 5973 6143 5979
rect 6091 5939 6100 5973
rect 6100 5939 6134 5973
rect 6134 5939 6143 5973
rect 6091 5927 6143 5939
rect 6091 5896 6143 5905
rect 6091 5862 6100 5896
rect 6100 5862 6134 5896
rect 6134 5862 6143 5896
rect 6091 5853 6143 5862
rect 6091 5819 6143 5831
rect 6091 5785 6100 5819
rect 6100 5785 6134 5819
rect 6134 5785 6143 5819
rect 6091 5779 6143 5785
rect 5653 5375 5705 5427
rect 5717 5375 5769 5427
rect 6034 5375 6086 5427
rect 6098 5375 6150 5427
rect 3886 5301 3938 5310
rect 3950 5301 4002 5310
rect 3886 5267 3918 5301
rect 3918 5267 3938 5301
rect 3950 5267 3952 5301
rect 3952 5267 3992 5301
rect 3992 5267 4002 5301
rect 3886 5258 3938 5267
rect 3950 5258 4002 5267
rect 3746 4189 3798 4241
rect 3746 4125 3798 4177
rect 3886 5041 3938 5050
rect 3950 5041 4002 5050
rect 3886 5007 3918 5041
rect 3918 5007 3938 5041
rect 3950 5007 3952 5041
rect 3952 5007 3991 5041
rect 3991 5007 4002 5041
rect 5874 5007 5886 5041
rect 5886 5007 5920 5041
rect 5920 5007 5926 5041
rect 3886 4998 3938 5007
rect 3950 4998 4002 5007
rect 5874 4989 5926 5007
rect 5942 5007 5958 5041
rect 5958 5007 5992 5041
rect 5992 5007 5994 5041
rect 5942 4989 5994 5007
rect 6010 5007 6030 5041
rect 6030 5007 6062 5041
rect 6078 5007 6102 5041
rect 6102 5007 6130 5041
rect 6146 5007 6174 5041
rect 6174 5007 6198 5041
rect 6214 5007 6246 5041
rect 6246 5007 6266 5041
rect 6010 4989 6062 5007
rect 6078 4989 6130 5007
rect 6146 4989 6198 5007
rect 6214 4989 6266 5007
rect 7792 6741 7844 6793
rect 7792 6677 7844 6729
rect 3886 4894 3938 4903
rect 3886 4860 3892 4894
rect 3892 4860 3926 4894
rect 3926 4860 3938 4894
rect 3886 4851 3938 4860
rect 3950 4894 4002 4903
rect 5874 4919 5926 4971
rect 5942 4919 5994 4971
rect 6010 4919 6062 4971
rect 6078 4919 6130 4971
rect 6146 4919 6198 4971
rect 6214 4919 6266 4971
rect 5874 4894 5926 4901
rect 5942 4894 5994 4901
rect 6010 4894 6062 4901
rect 6078 4894 6130 4901
rect 6146 4894 6198 4901
rect 6214 4894 6266 4901
rect 3950 4860 3965 4894
rect 3965 4860 3999 4894
rect 3999 4860 4002 4894
rect 5874 4860 5887 4894
rect 5887 4860 5925 4894
rect 5925 4860 5926 4894
rect 5942 4860 5959 4894
rect 5959 4860 5994 4894
rect 6010 4860 6031 4894
rect 6031 4860 6062 4894
rect 6078 4860 6103 4894
rect 6103 4860 6130 4894
rect 6146 4860 6175 4894
rect 6175 4860 6198 4894
rect 6214 4860 6247 4894
rect 6247 4860 6266 4894
rect 3950 4851 4002 4860
rect 5874 4849 5926 4860
rect 5942 4849 5994 4860
rect 6010 4849 6062 4860
rect 6078 4849 6130 4860
rect 6146 4849 6198 4860
rect 6214 4849 6266 4860
rect 5874 4779 5926 4831
rect 5942 4779 5994 4831
rect 6010 4779 6062 4831
rect 6078 4779 6130 4831
rect 6146 4779 6198 4831
rect 6214 4779 6266 4831
rect 5874 4709 5926 4761
rect 5942 4709 5994 4761
rect 6010 4709 6062 4761
rect 6078 4709 6130 4761
rect 6146 4709 6198 4761
rect 6214 4709 6266 4761
rect 5874 4679 5926 4691
rect 5874 4645 5878 4679
rect 5878 4645 5912 4679
rect 5912 4645 5926 4679
rect 5874 4639 5926 4645
rect 5942 4639 5994 4691
rect 6010 4639 6062 4691
rect 6078 4639 6130 4691
rect 6146 4639 6198 4691
rect 6214 4639 6266 4691
rect 5874 4568 5926 4620
rect 5942 4568 5994 4620
rect 6010 4568 6062 4620
rect 6078 4568 6130 4620
rect 6146 4568 6198 4620
rect 6214 4568 6266 4620
rect 5874 4537 5926 4549
rect 5874 4503 5878 4537
rect 5878 4503 5912 4537
rect 5912 4503 5926 4537
rect 5874 4497 5926 4503
rect 5942 4497 5994 4549
rect 6010 4497 6062 4549
rect 6078 4497 6130 4549
rect 6146 4497 6198 4549
rect 6214 4497 6266 4549
rect 4650 4443 4702 4453
rect 4714 4443 4766 4453
rect 4650 4409 4660 4443
rect 4660 4409 4699 4443
rect 4699 4409 4702 4443
rect 4714 4409 4733 4443
rect 4733 4409 4766 4443
rect 4650 4401 4702 4409
rect 4714 4401 4766 4409
rect 6327 4452 6379 4458
rect 6327 4418 6336 4452
rect 6336 4418 6370 4452
rect 6370 4418 6379 4452
rect 6327 4406 6379 4418
rect 6327 4377 6379 4388
rect 6327 4343 6336 4377
rect 6336 4343 6370 4377
rect 6370 4343 6379 4377
rect 6327 4336 6379 4343
rect 6327 4302 6379 4318
rect 6327 4268 6336 4302
rect 6336 4268 6370 4302
rect 6370 4268 6379 4302
rect 6327 4266 6379 4268
rect 6327 4227 6379 4249
rect 6327 4197 6336 4227
rect 6336 4197 6370 4227
rect 6370 4197 6379 4227
rect 6483 4265 6535 4271
rect 6547 4265 6599 4271
rect 6483 4231 6509 4265
rect 6509 4231 6535 4265
rect 6547 4231 6588 4265
rect 6588 4231 6599 4265
rect 6483 4219 6535 4231
rect 6547 4219 6599 4231
rect 7823 4251 7875 4303
rect 5653 4049 5705 4055
rect 5717 4049 5769 4055
rect 5653 4015 5683 4049
rect 5683 4015 5705 4049
rect 5717 4015 5756 4049
rect 5756 4015 5769 4049
rect 5653 4003 5705 4015
rect 5717 4003 5769 4015
rect 6327 4151 6379 4180
rect 6327 4128 6336 4151
rect 6336 4128 6370 4151
rect 6370 4128 6379 4151
rect 6327 4075 6379 4111
rect 6327 4059 6336 4075
rect 6336 4059 6370 4075
rect 6370 4059 6379 4075
rect 6327 4041 6336 4042
rect 6336 4041 6370 4042
rect 6370 4041 6379 4042
rect 6327 3999 6379 4041
rect 7823 4187 7875 4239
rect 8128 6537 8180 6589
rect 8128 6473 8180 6525
rect 6327 3990 6336 3999
rect 6336 3990 6370 3999
rect 6370 3990 6379 3999
rect 5879 3955 5931 3967
rect 5879 3921 5912 3955
rect 5912 3921 5931 3955
rect 5879 3915 5931 3921
rect 5962 3915 6014 3967
rect 6045 3915 6097 3967
rect 6127 3915 6179 3967
rect 6209 3915 6261 3967
rect 5879 3882 5931 3891
rect 5879 3848 5912 3882
rect 5912 3848 5931 3882
rect 5879 3839 5931 3848
rect 5962 3839 6014 3891
rect 6045 3839 6097 3891
rect 6127 3839 6179 3891
rect 6209 3839 6261 3891
rect 6327 3965 6336 3973
rect 6336 3965 6370 3973
rect 6370 3965 6379 3973
rect 6327 3923 6379 3965
rect 6327 3921 6336 3923
rect 6336 3921 6370 3923
rect 6370 3921 6379 3923
rect 5879 3809 5931 3815
rect 5879 3775 5912 3809
rect 5912 3775 5931 3809
rect 5879 3763 5931 3775
rect 5962 3763 6014 3815
rect 6045 3763 6097 3815
rect 6127 3763 6179 3815
rect 6209 3763 6261 3815
rect 4979 3651 5031 3703
rect 5043 3651 5095 3703
rect 10131 3462 10183 3514
rect 10197 3462 10249 3514
rect 10131 3398 10183 3450
rect 10197 3398 10249 3450
<< metal2 >>
rect 2303 39719 8224 39725
rect 2303 39667 2305 39719
rect 2357 39667 2369 39719
rect 2421 39667 8107 39719
rect 8159 39667 8171 39719
rect 8223 39667 8224 39719
rect 2303 39649 8224 39667
rect 2303 39597 2305 39649
rect 2357 39597 2369 39649
rect 2421 39597 8107 39649
rect 8159 39597 8171 39649
rect 8223 39597 8224 39649
rect 2303 39579 8224 39597
rect 2303 39527 2305 39579
rect 2357 39527 2369 39579
rect 2421 39527 8107 39579
rect 8159 39527 8171 39579
rect 8223 39527 8224 39579
rect 2303 39521 8224 39527
rect 9559 39719 10670 39725
rect 9611 39667 9623 39719
rect 9675 39667 10554 39719
rect 10606 39667 10618 39719
rect 9559 39649 10670 39667
rect 9611 39597 9623 39649
rect 9675 39597 10554 39649
rect 10606 39597 10618 39649
rect 9559 39579 10670 39597
rect 9611 39527 9623 39579
rect 9675 39527 10554 39579
rect 10606 39527 10618 39579
rect 9559 39521 10670 39527
rect 5595 39270 5663 39276
rect 5595 39267 5604 39270
rect 5656 39267 5663 39270
rect 5595 39211 5602 39267
rect 5658 39211 5663 39267
rect 5595 39206 5663 39211
rect 5595 39187 5604 39206
rect 5656 39187 5663 39206
rect 5595 39131 5602 39187
rect 5658 39131 5663 39187
rect 5595 39107 5604 39131
rect 5656 39107 5663 39131
rect 5595 39051 5602 39107
rect 5658 39051 5663 39107
rect 5595 39027 5604 39051
rect 5656 39027 5663 39051
rect 5595 38971 5602 39027
rect 5658 38971 5663 39027
rect 5595 38962 5604 38971
rect 5656 38962 5663 38971
rect 5595 38950 5663 38962
rect 5595 38947 5604 38950
rect 5656 38947 5663 38950
rect 5595 38891 5602 38947
rect 5658 38891 5663 38947
rect 5595 38886 5663 38891
rect 5595 38867 5604 38886
rect 5656 38867 5663 38886
rect 5595 38811 5602 38867
rect 5658 38811 5663 38867
rect 5595 38787 5604 38811
rect 5656 38787 5663 38811
rect 5595 38731 5602 38787
rect 5658 38731 5663 38787
rect 5595 38707 5604 38731
rect 5656 38707 5663 38731
rect 5595 38651 5602 38707
rect 5658 38651 5663 38707
rect 5595 38642 5604 38651
rect 5656 38642 5663 38651
rect 5595 38630 5663 38642
rect 5595 38627 5604 38630
rect 5656 38627 5663 38630
rect 5595 38571 5602 38627
rect 5658 38571 5663 38627
rect 5595 38566 5663 38571
rect 5595 38547 5604 38566
rect 5656 38547 5663 38566
rect 5595 38491 5602 38547
rect 5658 38491 5663 38547
rect 5595 38467 5604 38491
rect 5656 38467 5663 38491
rect 5595 38411 5602 38467
rect 5658 38411 5663 38467
rect 5595 38387 5604 38411
rect 5656 38387 5663 38411
rect 5595 38331 5602 38387
rect 5658 38331 5663 38387
rect 5595 38322 5604 38331
rect 5656 38322 5663 38331
rect 5595 38310 5663 38322
rect 5595 38307 5604 38310
rect 5656 38307 5663 38310
rect 5595 38251 5602 38307
rect 5658 38251 5663 38307
rect 5595 38246 5663 38251
rect 5595 38227 5604 38246
rect 5656 38227 5663 38246
rect 5595 38171 5602 38227
rect 5658 38171 5663 38227
rect 5595 38147 5604 38171
rect 5656 38147 5663 38171
rect 5595 38091 5602 38147
rect 5658 38091 5663 38147
rect 5595 38067 5604 38091
rect 5656 38067 5663 38091
rect 5595 38011 5602 38067
rect 5658 38011 5663 38067
rect 5595 38002 5604 38011
rect 5656 38002 5663 38011
rect 5595 37990 5663 38002
rect 5595 37987 5604 37990
rect 5656 37987 5663 37990
rect 5595 37931 5602 37987
rect 5658 37931 5663 37987
rect 5595 37926 5663 37931
rect 5595 37907 5604 37926
rect 5656 37907 5663 37926
rect 5595 37851 5602 37907
rect 5658 37851 5663 37907
rect 5595 37827 5604 37851
rect 5656 37827 5663 37851
rect 5595 37771 5602 37827
rect 5658 37771 5663 37827
rect 5595 37747 5604 37771
rect 5656 37747 5663 37771
rect 5595 37691 5602 37747
rect 5658 37691 5663 37747
rect 5595 37682 5604 37691
rect 5656 37682 5663 37691
rect 5595 37670 5663 37682
rect 5595 37667 5604 37670
rect 5656 37667 5663 37670
rect 5595 37611 5602 37667
rect 5658 37611 5663 37667
rect 5595 37606 5663 37611
rect 5595 37587 5604 37606
rect 5656 37587 5663 37606
rect 5595 37531 5602 37587
rect 5658 37531 5663 37587
rect 5595 37507 5604 37531
rect 5656 37507 5663 37531
rect 5595 37451 5602 37507
rect 5658 37451 5663 37507
rect 5595 37427 5604 37451
rect 5656 37427 5663 37451
rect 5595 37371 5602 37427
rect 5658 37371 5663 37427
rect 5595 37362 5604 37371
rect 5656 37362 5663 37371
rect 5595 37350 5663 37362
rect 5595 37347 5604 37350
rect 5656 37347 5663 37350
rect 5595 37291 5602 37347
rect 5658 37291 5663 37347
rect 5595 37286 5663 37291
rect 5595 37267 5604 37286
rect 5656 37267 5663 37286
rect 5595 37211 5602 37267
rect 5658 37211 5663 37267
rect 5595 37187 5604 37211
rect 5656 37187 5663 37211
rect 5595 37131 5602 37187
rect 5658 37131 5663 37187
rect 5595 37107 5604 37131
rect 5656 37107 5663 37131
rect 5595 37051 5602 37107
rect 5658 37051 5663 37107
rect 5595 37042 5604 37051
rect 5656 37042 5663 37051
rect 5595 37030 5663 37042
rect 5595 37027 5604 37030
rect 5656 37027 5663 37030
rect 5595 36971 5602 37027
rect 5658 36971 5663 37027
rect 5595 36966 5663 36971
rect 5595 36947 5604 36966
rect 5656 36947 5663 36966
rect 5595 36891 5602 36947
rect 5658 36891 5663 36947
rect 5595 36867 5604 36891
rect 5656 36867 5663 36891
rect 5595 36811 5602 36867
rect 5658 36811 5663 36867
rect 5595 36787 5604 36811
rect 5656 36787 5663 36811
rect 5595 36731 5602 36787
rect 5658 36731 5663 36787
rect 5595 36722 5604 36731
rect 5656 36722 5663 36731
rect 5595 36710 5663 36722
rect 5595 36707 5604 36710
rect 5656 36707 5663 36710
rect 5595 36651 5602 36707
rect 5658 36651 5663 36707
rect 5595 36646 5663 36651
rect 5595 36627 5604 36646
rect 5656 36627 5663 36646
rect 5595 36571 5602 36627
rect 5658 36571 5663 36627
rect 5595 36547 5604 36571
rect 5656 36547 5663 36571
rect 5595 36491 5602 36547
rect 5658 36491 5663 36547
rect 5595 36467 5604 36491
rect 5656 36467 5663 36491
rect 5595 36411 5602 36467
rect 5658 36411 5663 36467
rect 5595 36402 5604 36411
rect 5656 36402 5663 36411
rect 5595 36390 5663 36402
rect 5595 36387 5604 36390
rect 5656 36387 5663 36390
rect 5595 36331 5602 36387
rect 5658 36331 5663 36387
rect 5595 36326 5663 36331
rect 5595 36307 5604 36326
rect 5656 36307 5663 36326
rect 5595 36251 5602 36307
rect 5658 36251 5663 36307
rect 5595 36227 5604 36251
rect 5656 36227 5663 36251
rect 5595 36171 5602 36227
rect 5658 36171 5663 36227
rect 5595 36147 5604 36171
rect 5656 36147 5663 36171
rect 5595 36091 5602 36147
rect 5658 36091 5663 36147
rect 5595 36082 5604 36091
rect 5656 36082 5663 36091
rect 5595 36070 5663 36082
rect 5595 36067 5604 36070
rect 5656 36067 5663 36070
rect 5595 36011 5602 36067
rect 5658 36011 5663 36067
rect 5595 36006 5663 36011
rect 5595 35986 5604 36006
rect 5656 35986 5663 36006
rect 5595 35930 5602 35986
rect 5658 35930 5663 35986
rect 5595 35905 5604 35930
rect 5656 35905 5663 35930
rect 5595 35849 5602 35905
rect 5658 35849 5663 35905
rect 5595 35826 5604 35849
rect 5656 35826 5663 35849
rect 5595 35824 5663 35826
rect 5595 35768 5602 35824
rect 5658 35768 5663 35824
rect 5595 35762 5604 35768
rect 5656 35762 5663 35768
rect 5595 35750 5663 35762
rect 5595 35743 5604 35750
rect 5656 35743 5663 35750
rect 5595 35687 5602 35743
rect 5658 35687 5663 35743
rect 5595 35686 5663 35687
rect 5595 35662 5604 35686
rect 5656 35662 5663 35686
rect 5595 35606 5602 35662
rect 5658 35606 5663 35662
rect 5595 35581 5604 35606
rect 5656 35581 5663 35606
rect 5595 35525 5602 35581
rect 5658 35525 5663 35581
rect 5595 35506 5604 35525
rect 5656 35506 5663 35525
rect 5595 35500 5663 35506
rect 5595 35444 5602 35500
rect 5658 35444 5663 35500
rect 5595 35442 5604 35444
rect 5656 35442 5663 35444
rect 5595 35430 5663 35442
rect 5595 35419 5604 35430
rect 5656 35419 5663 35430
rect 5595 35363 5602 35419
rect 5658 35363 5663 35419
rect 5595 35338 5604 35363
rect 5656 35338 5663 35363
rect 5595 35282 5602 35338
rect 5658 35282 5663 35338
rect 5595 35257 5604 35282
rect 5656 35257 5663 35282
rect 5595 35201 5602 35257
rect 5658 35201 5663 35257
rect 5595 35186 5604 35201
rect 5656 35186 5663 35201
rect 5595 35176 5663 35186
rect 5595 35120 5602 35176
rect 5658 35120 5663 35176
rect 5595 35110 5663 35120
rect 5595 35095 5604 35110
rect 5656 35095 5663 35110
rect 5595 35039 5602 35095
rect 5658 35039 5663 35095
rect 5595 35014 5604 35039
rect 5656 35014 5663 35039
rect 5595 34958 5602 35014
rect 5658 34958 5663 35014
rect 5595 34933 5604 34958
rect 5656 34933 5663 34958
rect 5595 34877 5602 34933
rect 5658 34877 5663 34933
rect 7526 35001 8860 35007
rect 7578 34949 8784 35001
rect 8836 34949 8860 35001
rect 7526 34937 8860 34949
rect 7578 34885 8784 34937
rect 8836 34885 8860 34937
rect 7526 34879 8860 34885
rect 5595 34866 5604 34877
rect 5656 34866 5663 34877
rect 5595 34854 5663 34866
rect 5595 34852 5604 34854
rect 5656 34852 5663 34854
rect 5595 34796 5602 34852
rect 5658 34796 5663 34852
rect 5595 34790 5663 34796
rect 5595 34771 5604 34790
rect 5656 34771 5663 34790
rect 5595 34715 5602 34771
rect 5658 34715 5663 34771
rect 5595 34690 5604 34715
rect 5656 34690 5663 34715
rect 5595 34634 5602 34690
rect 5658 34634 5663 34690
rect 5595 34610 5604 34634
rect 5656 34610 5663 34634
rect 5595 34609 5663 34610
rect 5595 34553 5602 34609
rect 5658 34553 5663 34609
rect 5595 34546 5604 34553
rect 5656 34546 5663 34553
rect 5595 34534 5663 34546
rect 5595 34528 5604 34534
rect 5656 34528 5663 34534
rect 5595 34472 5602 34528
rect 5658 34472 5663 34528
rect 5595 34470 5663 34472
rect 5595 34447 5604 34470
rect 5656 34447 5663 34470
rect 5595 34391 5602 34447
rect 5658 34391 5663 34447
rect 5595 34366 5604 34391
rect 5656 34366 5663 34391
rect 5595 34310 5602 34366
rect 5658 34310 5663 34366
rect 5595 34290 5604 34310
rect 5656 34290 5663 34310
rect 5595 34285 5663 34290
rect 5595 34229 5602 34285
rect 5658 34229 5663 34285
rect 5595 34226 5604 34229
rect 5656 34226 5663 34229
rect 5595 34214 5663 34226
rect 5595 34204 5604 34214
rect 5656 34204 5663 34214
rect 5595 34148 5602 34204
rect 5658 34148 5663 34204
rect 5595 34123 5604 34148
rect 5656 34123 5663 34148
rect 5595 34067 5602 34123
rect 5658 34067 5663 34123
rect 5595 34042 5604 34067
rect 5656 34042 5663 34067
rect 5595 33986 5602 34042
rect 5658 33986 5663 34042
rect 5595 33970 5604 33986
rect 5656 33970 5663 33986
rect 5595 33961 5663 33970
rect 5595 33905 5602 33961
rect 5658 33905 5663 33961
rect 5595 33894 5663 33905
rect 5595 33880 5604 33894
rect 5656 33880 5663 33894
rect 5595 33824 5602 33880
rect 5658 33824 5663 33880
rect 5595 33799 5604 33824
rect 5656 33799 5663 33824
rect 5595 33743 5602 33799
rect 5658 33743 5663 33799
rect 5595 33718 5604 33743
rect 5656 33718 5663 33743
rect 5595 33662 5602 33718
rect 5658 33662 5663 33718
rect 5595 33650 5604 33662
rect 5656 33650 5663 33662
rect 5595 33638 5663 33650
rect 5595 33637 5604 33638
rect 5656 33637 5663 33638
rect 5595 33581 5602 33637
rect 5658 33581 5663 33637
rect 5595 33574 5663 33581
rect 5595 33556 5604 33574
rect 5656 33556 5663 33574
rect 5595 33500 5602 33556
rect 5658 33500 5663 33556
rect 5595 33475 5604 33500
rect 5656 33475 5663 33500
rect 5595 33419 5602 33475
rect 5658 33419 5663 33475
rect 5595 33394 5604 33419
rect 5656 33394 5663 33419
rect 5595 33338 5602 33394
rect 5658 33338 5663 33394
rect 5595 33330 5604 33338
rect 5656 33330 5663 33338
rect 5595 33318 5663 33330
rect 5595 33313 5604 33318
rect 5656 33313 5663 33318
rect 5595 33257 5602 33313
rect 5658 33257 5663 33313
rect 5595 33254 5663 33257
rect 5595 33232 5604 33254
rect 5656 33232 5663 33254
rect 5595 33176 5602 33232
rect 5658 33176 5663 33232
rect 5595 33151 5604 33176
rect 5656 33151 5663 33176
rect 5595 33095 5602 33151
rect 5658 33095 5663 33151
rect 5595 33074 5604 33095
rect 5656 33074 5663 33095
rect 5595 33070 5663 33074
rect 5595 33014 5602 33070
rect 5658 33014 5663 33070
rect 5595 33010 5604 33014
rect 5656 33010 5663 33014
rect 5595 32998 5663 33010
rect 5595 32989 5604 32998
rect 5656 32989 5663 32998
rect 5595 32933 5602 32989
rect 5658 32933 5663 32989
rect 5595 32908 5604 32933
rect 5656 32908 5663 32933
rect 5595 32852 5602 32908
rect 5658 32852 5663 32908
rect 5595 32827 5604 32852
rect 5656 32827 5663 32852
rect 5595 32771 5602 32827
rect 5658 32771 5663 32827
rect 5595 32754 5604 32771
rect 5656 32754 5663 32771
rect 5595 32746 5663 32754
rect 5595 32690 5602 32746
rect 5658 32690 5663 32746
rect 5595 32677 5663 32690
rect 5595 32665 5604 32677
rect 5656 32665 5663 32677
rect 5595 32609 5602 32665
rect 5658 32609 5663 32665
rect 5595 32584 5604 32609
rect 5656 32584 5663 32609
rect 5595 32528 5602 32584
rect 5658 32528 5663 32584
rect 5595 32503 5604 32528
rect 5656 32503 5663 32528
rect 5595 32447 5602 32503
rect 5658 32447 5663 32503
rect 5595 32430 5604 32447
rect 5656 32430 5663 32447
rect 5595 32422 5663 32430
rect 5595 32366 5602 32422
rect 5658 32366 5663 32422
rect 5595 32365 5604 32366
rect 5656 32365 5663 32366
rect 5595 32352 5663 32365
rect 5595 32341 5604 32352
rect 5656 32341 5663 32352
rect 5595 32285 5602 32341
rect 5658 32285 5663 32341
rect 5595 32260 5604 32285
rect 5656 32260 5663 32285
rect 5595 32204 5602 32260
rect 5658 32204 5663 32260
rect 5595 32179 5604 32204
rect 5656 32179 5663 32204
rect 5595 32123 5602 32179
rect 5658 32123 5663 32179
rect 5595 32105 5604 32123
rect 5656 32105 5663 32123
rect 5595 32098 5663 32105
rect 5595 32042 5602 32098
rect 5658 32042 5663 32098
rect 5595 32040 5604 32042
rect 5656 32040 5663 32042
rect 5595 32027 5663 32040
rect 5595 32017 5604 32027
rect 5656 32017 5663 32027
rect 5595 31961 5602 32017
rect 5658 31961 5663 32017
rect 5595 31936 5604 31961
rect 5656 31936 5663 31961
rect 5595 31880 5602 31936
rect 5658 31880 5663 31936
rect 5595 31855 5604 31880
rect 5656 31855 5663 31880
rect 5595 31799 5602 31855
rect 5658 31799 5663 31855
rect 5595 31780 5604 31799
rect 5656 31780 5663 31799
rect 5595 31774 5663 31780
rect 5595 31718 5602 31774
rect 5658 31718 5663 31774
rect 5595 31715 5604 31718
rect 5656 31715 5663 31718
rect 5595 31702 5663 31715
rect 5595 31693 5604 31702
rect 5656 31693 5663 31702
rect 5595 31637 5602 31693
rect 5658 31637 5663 31693
rect 5595 31612 5604 31637
rect 5656 31612 5663 31637
rect 7526 31753 8120 31759
rect 7578 31701 8068 31753
rect 7526 31689 8120 31701
rect 7578 31637 8068 31689
rect 7526 31631 8120 31637
rect 5595 31556 5602 31612
rect 5658 31556 5663 31612
rect 5595 31531 5604 31556
rect 5656 31531 5663 31556
rect 5595 31475 5602 31531
rect 5658 31475 5663 31531
rect 5595 31455 5604 31475
rect 5656 31455 5663 31475
rect 5595 31450 5663 31455
rect 5595 31394 5602 31450
rect 5658 31394 5663 31450
rect 5595 31390 5604 31394
rect 5656 31390 5663 31394
rect 5595 31377 5663 31390
rect 5595 31369 5604 31377
rect 5656 31369 5663 31377
rect 5595 31313 5602 31369
rect 5658 31313 5663 31369
rect 5595 31312 5663 31313
rect 5595 31288 5604 31312
rect 5656 31288 5663 31312
rect 5595 31232 5602 31288
rect 5658 31232 5663 31288
rect 5595 31207 5604 31232
rect 5656 31207 5663 31232
rect 5595 31151 5602 31207
rect 5658 31151 5663 31207
rect 5595 31130 5604 31151
rect 5656 31130 5663 31151
rect 5595 31126 5663 31130
rect 5595 31070 5602 31126
rect 5658 31070 5663 31126
rect 5595 31065 5604 31070
rect 5656 31065 5663 31070
rect 5595 31052 5663 31065
rect 5595 31045 5604 31052
rect 5656 31045 5663 31052
rect 5595 30989 5602 31045
rect 5658 30989 5663 31045
rect 5595 30987 5663 30989
rect 5595 30964 5604 30987
rect 5656 30964 5663 30987
rect 5595 30908 5602 30964
rect 5658 30908 5663 30964
rect 5595 30883 5604 30908
rect 5656 30883 5663 30908
rect 5595 30827 5602 30883
rect 5658 30827 5663 30883
rect 5595 30805 5604 30827
rect 5656 30805 5663 30827
rect 5595 30802 5663 30805
rect 5595 30746 5602 30802
rect 5658 30746 5663 30802
rect 5595 30740 5604 30746
rect 5656 30740 5663 30746
rect 5595 30727 5663 30740
rect 5595 30721 5604 30727
rect 5656 30721 5663 30727
rect 5595 30665 5602 30721
rect 5658 30665 5663 30721
rect 5595 30662 5663 30665
rect 5595 30640 5604 30662
rect 5656 30640 5663 30662
rect 5595 30584 5602 30640
rect 5658 30584 5663 30640
rect 5595 30559 5604 30584
rect 5656 30559 5663 30584
rect 5595 30503 5602 30559
rect 5658 30503 5663 30559
rect 5595 30480 5604 30503
rect 5656 30480 5663 30503
rect 5595 30478 5663 30480
rect 5595 30422 5602 30478
rect 5658 30422 5663 30478
rect 5595 30415 5604 30422
rect 5656 30415 5663 30422
rect 5595 30402 5663 30415
rect 5595 30397 5604 30402
rect 5656 30397 5663 30402
rect 5595 30341 5602 30397
rect 5658 30341 5663 30397
rect 5595 30332 5663 30341
rect 5610 29859 5714 29911
rect 5766 29859 5801 29911
rect 5853 29859 5859 29911
rect 5610 29835 5859 29859
rect 7577 29842 7583 29894
rect 7635 29842 7647 29894
rect 7699 29842 9094 29894
rect 9146 29842 9158 29894
rect 9210 29842 9216 29894
rect 5610 29783 5714 29835
rect 5766 29783 5801 29835
rect 5853 29783 5859 29835
rect 7497 29762 7503 29814
rect 7555 29762 7567 29814
rect 7619 29808 9060 29814
rect 7619 29762 9008 29808
tri 8974 29756 8980 29762 ne
rect 8980 29756 9008 29762
tri 8980 29744 8992 29756 ne
rect 8992 29744 9060 29756
tri 8992 29728 9008 29744 ne
rect 7316 29647 7322 29699
rect 7374 29647 7386 29699
rect 7438 29693 8980 29699
rect 7438 29647 8928 29693
rect 9008 29686 9060 29692
rect 8928 29629 8980 29641
rect 8928 29571 8980 29577
rect 6733 27282 7800 27310
rect 6733 27280 6742 27282
rect 6798 27280 6825 27282
rect 6881 27280 6908 27282
rect 6964 27280 6991 27282
rect 7047 27280 7074 27282
rect 7130 27280 7157 27282
rect 7213 27280 7240 27282
rect 7296 27280 7323 27282
rect 7379 27280 7406 27282
rect 7462 27280 7489 27282
rect 7545 27280 7571 27282
rect 7627 27280 7653 27282
rect 7709 27280 7735 27282
rect 7791 27280 7800 27282
rect 6733 27228 6739 27280
rect 6798 27228 6806 27280
rect 7059 27228 7074 27280
rect 7130 27228 7141 27280
rect 7394 27228 7406 27280
rect 7462 27228 7476 27280
rect 7728 27228 7735 27280
rect 7794 27228 7800 27280
rect 6733 27226 6742 27228
rect 6798 27226 6825 27228
rect 6881 27226 6908 27228
rect 6964 27226 6991 27228
rect 7047 27226 7074 27228
rect 7130 27226 7157 27228
rect 7213 27226 7240 27228
rect 7296 27226 7323 27228
rect 7379 27226 7406 27228
rect 7462 27226 7489 27228
rect 7545 27226 7571 27228
rect 7627 27226 7653 27228
rect 7709 27226 7735 27228
rect 7791 27226 7800 27228
rect 6733 27197 7800 27226
rect 4663 27086 4669 27138
rect 4721 27101 4736 27138
rect 4788 27101 4803 27138
rect 4855 27101 4870 27138
rect 4922 27101 4937 27138
rect 4728 27086 4736 27101
rect 4922 27086 4926 27101
rect 4989 27086 5004 27138
rect 5056 27101 5071 27138
rect 5123 27101 5138 27138
rect 5190 27101 5205 27138
rect 5257 27101 5272 27138
rect 5066 27086 5071 27101
rect 5257 27086 5262 27101
rect 5324 27086 5339 27138
rect 5391 27101 5406 27138
rect 5458 27101 5473 27138
rect 5525 27101 5539 27138
rect 5591 27101 5605 27138
rect 5402 27086 5406 27101
rect 5591 27086 5598 27101
rect 5657 27086 5663 27138
rect 4663 27060 4672 27086
rect 4728 27060 4757 27086
rect 4813 27060 4842 27086
rect 4898 27060 4926 27086
rect 4982 27060 5010 27086
rect 5066 27060 5094 27086
rect 5150 27060 5178 27086
rect 5234 27060 5262 27086
rect 5318 27060 5346 27086
rect 5402 27060 5430 27086
rect 5486 27060 5514 27086
rect 5570 27060 5598 27086
rect 5654 27060 5663 27086
rect 4663 27008 4669 27060
rect 4728 27045 4736 27060
rect 4922 27045 4926 27060
rect 4721 27008 4736 27045
rect 4788 27008 4803 27045
rect 4855 27008 4870 27045
rect 4922 27008 4937 27045
rect 4989 27008 5004 27060
rect 5066 27045 5071 27060
rect 5257 27045 5262 27060
rect 5056 27008 5071 27045
rect 5123 27008 5138 27045
rect 5190 27008 5205 27045
rect 5257 27008 5272 27045
rect 5324 27008 5339 27060
rect 5402 27045 5406 27060
rect 5591 27045 5598 27060
rect 5391 27008 5406 27045
rect 5458 27008 5473 27045
rect 5525 27008 5539 27045
rect 5591 27008 5605 27045
rect 5657 27008 5663 27060
rect 6473 27130 8860 27136
rect 6473 27124 8784 27130
rect 6473 27008 6479 27124
rect 6595 27078 8784 27124
rect 8836 27078 8860 27130
rect 6595 27066 8860 27078
rect 6595 27014 8784 27066
rect 8836 27014 8860 27066
rect 6595 27008 8860 27014
rect 656 26358 8860 26364
rect 708 26306 8784 26358
rect 8836 26306 8860 26358
rect 656 26294 8860 26306
rect 708 26242 8784 26294
rect 8836 26242 8860 26294
rect 656 26236 8860 26242
rect 6077 22131 6086 22133
rect 6142 22131 6166 22133
rect 6077 22079 6083 22131
rect 6142 22079 6147 22131
rect 6077 22077 6086 22079
rect 6142 22077 6166 22079
rect 6222 22077 6231 22133
rect 6610 21374 6675 21426
rect 6727 21374 6739 21426
rect 6791 21374 8809 21426
rect 8861 21374 8873 21426
rect 8925 21374 8931 21426
rect 9008 21416 9060 21422
tri 9002 21374 9008 21380 se
tri 8992 21364 9002 21374 se
rect 9002 21364 9008 21374
tri 8980 21352 8992 21364 se
rect 8992 21352 9060 21364
tri 8974 21346 8980 21352 se
rect 8980 21346 9008 21352
rect 6457 21294 6592 21346
rect 6644 21294 6656 21346
rect 6708 21300 9008 21346
rect 6708 21294 9060 21300
rect 6417 21214 6423 21266
rect 6475 21214 6487 21266
rect 6539 21214 9094 21266
rect 9146 21214 9158 21266
rect 9210 21214 9216 21266
rect 4722 7727 6533 7729
rect 4722 7710 5110 7727
rect 5166 7710 5192 7727
rect 5248 7710 5274 7727
rect 4722 7658 4728 7710
rect 4780 7658 4800 7710
rect 4852 7658 4871 7710
rect 4923 7658 4942 7710
rect 4994 7658 5013 7710
rect 5065 7658 5084 7710
rect 5330 7671 5355 7727
rect 5411 7671 5436 7727
rect 5492 7671 5517 7727
rect 5573 7671 5598 7727
rect 5654 7723 6533 7727
rect 5654 7719 6481 7723
rect 5136 7658 5155 7671
rect 5207 7658 5226 7671
rect 5278 7667 5649 7671
rect 5701 7667 5723 7719
rect 5775 7667 5797 7719
rect 5849 7700 6481 7719
rect 5849 7667 6197 7700
rect 5278 7658 6197 7667
rect 4722 7648 6197 7658
rect 6249 7648 6271 7700
rect 6323 7648 6345 7700
rect 6397 7671 6481 7700
rect 6397 7648 6533 7671
rect 4722 7644 6481 7648
rect 4722 7636 5649 7644
rect 4722 7584 4728 7636
rect 4780 7584 4800 7636
rect 4852 7584 4871 7636
rect 4923 7584 4942 7636
rect 4994 7584 5013 7636
rect 5065 7584 5084 7636
rect 5136 7631 5155 7636
rect 5207 7631 5226 7636
rect 5278 7631 5649 7636
rect 4722 7575 5110 7584
rect 5166 7575 5192 7584
rect 5248 7575 5274 7584
rect 5330 7575 5355 7631
rect 5411 7575 5436 7631
rect 5492 7575 5517 7631
rect 5573 7575 5598 7631
rect 5701 7592 5723 7644
rect 5775 7592 5797 7644
rect 5849 7629 6481 7644
rect 5849 7592 6197 7629
rect 5654 7577 6197 7592
rect 6249 7577 6271 7629
rect 6323 7577 6345 7629
rect 6397 7596 6481 7629
rect 6397 7577 6533 7596
rect 5654 7575 6533 7577
rect 4722 7573 6533 7575
rect 4722 7569 6481 7573
rect 4722 7562 5649 7569
rect 4722 7510 4728 7562
rect 4780 7510 4800 7562
rect 4852 7510 4871 7562
rect 4923 7510 4942 7562
rect 4994 7510 5013 7562
rect 5065 7510 5084 7562
rect 5136 7535 5155 7562
rect 5207 7535 5226 7562
rect 5278 7535 5649 7562
rect 4722 7488 5110 7510
rect 5166 7488 5192 7510
rect 5248 7488 5274 7510
rect 4722 7436 4728 7488
rect 4780 7436 4800 7488
rect 4852 7436 4871 7488
rect 4923 7436 4942 7488
rect 4994 7436 5013 7488
rect 5065 7436 5084 7488
rect 5330 7479 5355 7535
rect 5411 7479 5436 7535
rect 5492 7479 5517 7535
rect 5573 7479 5598 7535
rect 5701 7517 5723 7569
rect 5775 7517 5797 7569
rect 5849 7558 6481 7569
rect 5849 7517 6197 7558
rect 5654 7506 6197 7517
rect 6249 7506 6271 7558
rect 6323 7506 6345 7558
rect 6397 7521 6481 7558
rect 6397 7506 6533 7521
rect 5654 7497 6533 7506
rect 5654 7494 6481 7497
rect 5136 7439 5155 7479
rect 5207 7439 5226 7479
rect 5278 7442 5649 7479
rect 5701 7442 5723 7494
rect 5775 7442 5797 7494
rect 5849 7487 6481 7494
rect 5849 7442 6197 7487
rect 5278 7439 6197 7442
rect 4722 7414 5110 7436
rect 5166 7414 5192 7436
rect 5248 7414 5274 7436
rect 4722 7362 4728 7414
rect 4780 7362 4800 7414
rect 4852 7362 4871 7414
rect 4923 7362 4942 7414
rect 4994 7362 5013 7414
rect 5065 7362 5084 7414
rect 5330 7383 5355 7439
rect 5411 7383 5436 7439
rect 5492 7383 5517 7439
rect 5573 7383 5598 7439
rect 5654 7435 6197 7439
rect 6249 7435 6271 7487
rect 6323 7435 6345 7487
rect 6397 7445 6481 7487
rect 6397 7435 6533 7445
rect 5654 7421 6533 7435
rect 5654 7419 6481 7421
rect 5136 7362 5155 7383
rect 5207 7362 5226 7383
rect 5278 7367 5649 7383
rect 5701 7367 5723 7419
rect 5775 7367 5797 7419
rect 5849 7416 6481 7419
rect 5849 7367 6197 7416
rect 5278 7364 6197 7367
rect 6249 7364 6271 7416
rect 6323 7364 6345 7416
rect 6397 7369 6481 7416
rect 6397 7364 6533 7369
rect 5278 7362 6533 7364
rect 4722 7345 6533 7362
rect 4722 7344 6197 7345
rect 4722 7343 5649 7344
rect 4722 7340 5110 7343
rect 5166 7340 5192 7343
rect 5248 7340 5274 7343
rect 4722 7288 4728 7340
rect 4780 7288 4800 7340
rect 4852 7288 4871 7340
rect 4923 7288 4942 7340
rect 4994 7288 5013 7340
rect 5065 7288 5084 7340
rect 4722 7287 5110 7288
rect 5166 7287 5192 7288
rect 5248 7287 5274 7288
rect 5330 7287 5355 7343
rect 5411 7287 5436 7343
rect 5492 7287 5517 7343
rect 5573 7287 5598 7343
rect 5701 7292 5723 7344
rect 5775 7292 5797 7344
rect 5849 7293 6197 7344
rect 6249 7293 6271 7345
rect 6323 7293 6345 7345
rect 6397 7293 6481 7345
rect 5849 7292 6533 7293
rect 5654 7287 6533 7292
rect 4722 7286 6533 7287
rect 7792 6793 7844 6799
tri 7776 6741 7792 6757 se
tri 7764 6729 7776 6741 se
rect 7776 6729 7844 6741
tri 7758 6723 7764 6729 se
rect 7764 6723 7792 6729
rect 6263 6671 6269 6723
rect 6321 6671 6369 6723
rect 6421 6677 7792 6723
rect 6421 6671 7844 6677
rect 5809 6589 5861 6595
rect 656 6523 4637 6529
rect 708 6471 3847 6523
rect 3899 6471 4577 6523
rect 4629 6471 4637 6523
rect 656 6459 4637 6471
rect 5809 6525 5861 6537
rect 8128 6589 8180 6595
rect 8128 6525 8180 6537
rect 5861 6473 8128 6519
rect 5809 6467 8180 6473
rect 708 6407 3847 6459
rect 3899 6407 4577 6459
rect 4629 6407 4637 6459
rect 656 6401 4637 6407
rect 6028 6272 6156 6278
rect 6028 6220 6091 6272
rect 6143 6220 6156 6272
rect 6028 6199 6156 6220
rect 6028 6147 6091 6199
rect 6143 6147 6156 6199
rect 6028 6126 6156 6147
rect 6028 6074 6091 6126
rect 6143 6074 6156 6126
rect 6028 6053 6156 6074
tri 3689 6033 3695 6039 se
rect 3695 6033 5595 6039
tri 3637 5981 3689 6033 se
rect 3689 5981 5543 6033
tri 3635 5979 3637 5981 se
rect 3637 5979 5595 5981
tri 3625 5969 3635 5979 se
rect 3635 5969 5595 5979
tri 3573 5917 3625 5969 se
rect 3625 5917 5543 5969
tri 3567 5911 3573 5917 se
rect 3573 5911 5595 5917
rect 6028 6001 6091 6053
rect 6143 6001 6156 6053
rect 6028 5979 6156 6001
rect 6028 5927 6091 5979
rect 6143 5927 6156 5979
tri 3561 5905 3567 5911 se
rect 3567 5905 3743 5911
tri 3743 5905 3749 5911 nw
rect 6028 5905 6156 5927
tri 3513 5857 3561 5905 se
rect 3561 5857 3695 5905
tri 3695 5857 3743 5905 nw
tri 3509 5853 3513 5857 se
rect 3513 5853 3691 5857
tri 3691 5853 3695 5857 nw
rect 6028 5853 6091 5905
rect 6143 5853 6156 5905
tri 3487 5831 3509 5853 se
rect 3509 5831 3669 5853
tri 3669 5831 3691 5853 nw
rect 6028 5831 6156 5853
tri 3482 5826 3487 5831 se
rect 3487 5826 3664 5831
tri 3664 5826 3669 5831 nw
rect 3482 5779 3617 5826
tri 3617 5779 3664 5826 nw
rect 6028 5779 6091 5831
rect 6143 5779 6156 5831
rect 3482 5677 3610 5779
tri 3610 5772 3617 5779 nw
rect 3482 5625 3488 5677
rect 3540 5625 3552 5677
rect 3604 5625 3610 5677
rect 6028 5427 6156 5779
rect 5647 5375 5653 5427
rect 5705 5375 5717 5427
rect 5769 5375 5775 5427
rect 6028 5375 6034 5427
rect 6086 5375 6098 5427
rect 6150 5375 6156 5427
rect 6327 6228 6379 6234
rect 6327 6164 6379 6176
rect 3527 5258 3533 5310
rect 3585 5258 3597 5310
rect 3649 5258 3886 5310
rect 3938 5258 3950 5310
rect 4002 5258 4008 5310
rect 3527 4998 3533 5050
rect 3585 4998 3597 5050
rect 3649 4998 3886 5050
rect 3938 4998 3950 5050
rect 4002 4998 4008 5050
rect 656 4852 708 4858
rect 3527 4851 3533 4903
rect 3585 4851 3597 4903
rect 3649 4851 3886 4903
rect 3938 4851 3950 4903
rect 4002 4851 4008 4903
rect 656 4788 708 4800
tri 708 4782 742 4816 sw
rect 708 4736 3126 4782
rect 656 4730 3126 4736
rect 3178 4730 3220 4782
rect 3272 4730 3314 4782
rect 3366 4730 3372 4782
rect 512 4455 3828 4461
rect 628 4403 2985 4455
rect 3037 4403 3297 4455
rect 3349 4403 3609 4455
rect 3661 4403 3828 4455
rect 628 4391 3828 4403
rect 628 4339 2985 4391
rect 3037 4339 3297 4391
rect 3349 4339 3609 4391
rect 3661 4339 3828 4391
rect 512 4333 3828 4339
rect 4644 4401 4650 4453
rect 4702 4401 4714 4453
rect 4766 4401 4772 4453
tri 4593 4266 4644 4317 se
rect 4644 4266 4772 4401
tri 4576 4249 4593 4266 se
rect 4593 4249 4772 4266
tri 4574 4247 4576 4249 se
rect 4576 4247 4772 4249
rect 3141 4241 4772 4247
rect 3193 4189 3453 4241
rect 3505 4189 3746 4241
rect 3798 4189 4772 4241
rect 3141 4177 4772 4189
rect 3193 4125 3453 4177
rect 3505 4125 3746 4177
rect 3798 4125 4772 4177
rect 3141 4119 4772 4125
rect 5647 4055 5775 5375
rect 5647 4003 5653 4055
rect 5705 4003 5717 4055
rect 5769 4003 5775 4055
rect 5647 4002 5775 4003
rect 5873 5041 6267 5047
rect 5873 4982 5874 5041
rect 5926 5038 5942 5041
rect 5994 5038 6010 5041
rect 6062 5038 6078 5041
rect 6130 5038 6146 5041
rect 6198 5038 6214 5041
rect 5930 4989 5942 5038
rect 6198 4989 6210 5038
rect 5930 4982 5958 4989
rect 6014 4982 6042 4989
rect 6098 4982 6126 4989
rect 6182 4982 6210 4989
rect 6266 4982 6267 5041
rect 5873 4971 6267 4982
rect 5873 4902 5874 4971
rect 5926 4958 5942 4971
rect 5994 4958 6010 4971
rect 6062 4958 6078 4971
rect 6130 4958 6146 4971
rect 6198 4958 6214 4971
rect 5930 4919 5942 4958
rect 6198 4919 6210 4958
rect 5930 4902 5958 4919
rect 6014 4902 6042 4919
rect 6098 4902 6126 4919
rect 6182 4902 6210 4919
rect 6266 4902 6267 4971
rect 5873 4901 6267 4902
rect 5873 4639 5874 4901
rect 5926 4878 5942 4901
rect 5994 4878 6010 4901
rect 6062 4878 6078 4901
rect 6130 4878 6146 4901
rect 6198 4878 6214 4901
rect 5930 4849 5942 4878
rect 6198 4849 6210 4878
rect 5930 4831 5958 4849
rect 6014 4831 6042 4849
rect 6098 4831 6126 4849
rect 6182 4831 6210 4849
rect 5930 4822 5942 4831
rect 6198 4822 6210 4831
rect 5926 4798 5942 4822
rect 5994 4798 6010 4822
rect 6062 4798 6078 4822
rect 6130 4798 6146 4822
rect 6198 4798 6214 4822
rect 5930 4779 5942 4798
rect 6198 4779 6210 4798
rect 5930 4761 5958 4779
rect 6014 4761 6042 4779
rect 6098 4761 6126 4779
rect 6182 4761 6210 4779
rect 5930 4742 5942 4761
rect 6198 4742 6210 4761
rect 5926 4718 5942 4742
rect 5994 4718 6010 4742
rect 6062 4718 6078 4742
rect 6130 4718 6146 4742
rect 6198 4718 6214 4742
rect 5930 4709 5942 4718
rect 6198 4709 6210 4718
rect 5930 4691 5958 4709
rect 6014 4691 6042 4709
rect 6098 4691 6126 4709
rect 6182 4691 6210 4709
rect 5930 4662 5942 4691
rect 6198 4662 6210 4691
rect 5926 4639 5942 4662
rect 5994 4639 6010 4662
rect 6062 4639 6078 4662
rect 6130 4639 6146 4662
rect 6198 4639 6214 4662
rect 6266 4639 6267 4901
rect 5873 4638 6267 4639
rect 5873 4568 5874 4638
rect 5930 4620 5958 4638
rect 6014 4620 6042 4638
rect 6098 4620 6126 4638
rect 6182 4620 6210 4638
rect 5930 4582 5942 4620
rect 6198 4582 6210 4620
rect 5926 4568 5942 4582
rect 5994 4568 6010 4582
rect 6062 4568 6078 4582
rect 6130 4568 6146 4582
rect 6198 4568 6214 4582
rect 6266 4568 6267 4638
rect 5873 4557 6267 4568
rect 5873 4497 5874 4557
rect 5930 4549 5958 4557
rect 6014 4549 6042 4557
rect 6098 4549 6126 4557
rect 6182 4549 6210 4557
rect 5930 4501 5942 4549
rect 6198 4501 6210 4549
rect 5926 4497 5942 4501
rect 5994 4497 6010 4501
rect 6062 4497 6078 4501
rect 6130 4497 6146 4501
rect 6198 4497 6214 4501
rect 6266 4497 6267 4557
rect 5873 4476 6267 4497
rect 5873 4420 5874 4476
rect 5930 4420 5958 4476
rect 6014 4420 6042 4476
rect 6098 4420 6126 4476
rect 6182 4420 6210 4476
rect 6266 4420 6267 4476
rect 5873 4395 6267 4420
rect 5873 4339 5874 4395
rect 5930 4339 5958 4395
rect 6014 4339 6042 4395
rect 6098 4339 6126 4395
rect 6182 4339 6210 4395
rect 6266 4339 6267 4395
rect 5873 4314 6267 4339
rect 5873 4258 5874 4314
rect 5930 4258 5958 4314
rect 6014 4258 6042 4314
rect 6098 4258 6126 4314
rect 6182 4258 6210 4314
rect 6266 4258 6267 4314
rect 5873 4233 6267 4258
rect 5873 4177 5874 4233
rect 5930 4177 5958 4233
rect 6014 4177 6042 4233
rect 6098 4177 6126 4233
rect 6182 4177 6210 4233
rect 6266 4177 6267 4233
rect 5873 4152 6267 4177
rect 5873 4096 5874 4152
rect 5930 4096 5958 4152
rect 6014 4096 6042 4152
rect 6098 4096 6126 4152
rect 6182 4096 6210 4152
rect 6266 4096 6267 4152
rect 5873 4071 6267 4096
rect 5873 4015 5874 4071
rect 5930 4015 5958 4071
rect 6014 4015 6042 4071
rect 6098 4015 6126 4071
rect 6182 4015 6210 4071
rect 6266 4015 6267 4071
rect 5873 3990 6267 4015
rect 5873 3934 5874 3990
rect 5930 3967 5958 3990
rect 5931 3934 5958 3967
rect 6014 3934 6042 3990
rect 6098 3934 6126 3990
rect 6182 3967 6210 3990
rect 6182 3934 6209 3967
rect 6266 3934 6267 3990
rect 5873 3915 5879 3934
rect 5931 3915 5962 3934
rect 6014 3915 6045 3934
rect 6097 3915 6127 3934
rect 6179 3915 6209 3934
rect 6261 3915 6267 3934
rect 5873 3909 6267 3915
rect 5873 3853 5874 3909
rect 5930 3891 5958 3909
rect 5931 3853 5958 3891
rect 6014 3853 6042 3909
rect 6098 3853 6126 3909
rect 6182 3891 6210 3909
rect 6182 3853 6209 3891
rect 6266 3853 6267 3909
rect 5873 3839 5879 3853
rect 5931 3839 5962 3853
rect 6014 3839 6045 3853
rect 6097 3839 6127 3853
rect 6179 3839 6209 3853
rect 6261 3839 6267 3853
rect 5873 3828 6267 3839
rect 5873 3772 5874 3828
rect 5930 3815 5958 3828
rect 5931 3772 5958 3815
rect 6014 3772 6042 3828
rect 6098 3772 6126 3828
rect 6182 3815 6210 3828
rect 6182 3772 6209 3815
rect 6266 3772 6267 3828
rect 5873 3763 5879 3772
rect 5931 3763 5962 3772
rect 6014 3763 6045 3772
rect 6097 3763 6127 3772
rect 6179 3763 6209 3772
rect 6261 3763 6267 3772
rect 6327 4458 6379 6112
rect 6327 4388 6379 4406
rect 6327 4318 6379 4336
tri 7821 4303 7823 4305 se
rect 7823 4303 7875 4309
tri 7789 4271 7821 4303 se
rect 7821 4271 7823 4303
rect 6327 4249 6379 4266
rect 6418 4225 6483 4271
rect 6477 4219 6483 4225
rect 6535 4219 6547 4271
rect 6599 4251 7823 4271
rect 6599 4239 7875 4251
rect 6599 4225 7823 4239
rect 6599 4219 6605 4225
tri 7789 4219 7795 4225 ne
rect 7795 4219 7823 4225
rect 6327 4180 6379 4197
tri 7795 4191 7823 4219 ne
rect 7823 4181 7875 4187
rect 6327 4111 6379 4128
rect 6327 4042 6379 4059
rect 6327 3973 6379 3990
tri 6293 3703 6327 3737 se
rect 6327 3703 6379 3921
rect 4973 3651 4979 3703
rect 5031 3651 5043 3703
rect 5095 3651 6379 3703
rect 5823 3514 10249 3520
rect 5823 3484 10131 3514
rect 5823 3428 5832 3484
rect 5888 3428 5953 3484
rect 6009 3428 6074 3484
rect 6130 3428 6195 3484
rect 6251 3428 6316 3484
rect 6372 3428 6437 3484
rect 6493 3428 6558 3484
rect 6614 3462 10131 3484
rect 10183 3462 10197 3514
rect 6614 3450 10249 3462
rect 6614 3428 10131 3450
rect 5823 3398 10131 3428
rect 10183 3398 10197 3450
rect 5823 3392 10249 3398
<< via2 >>
rect 5602 39218 5604 39267
rect 5604 39218 5656 39267
rect 5656 39218 5658 39267
rect 5602 39211 5658 39218
rect 5602 39154 5604 39187
rect 5604 39154 5656 39187
rect 5656 39154 5658 39187
rect 5602 39142 5658 39154
rect 5602 39131 5604 39142
rect 5604 39131 5656 39142
rect 5656 39131 5658 39142
rect 5602 39090 5604 39107
rect 5604 39090 5656 39107
rect 5656 39090 5658 39107
rect 5602 39078 5658 39090
rect 5602 39051 5604 39078
rect 5604 39051 5656 39078
rect 5656 39051 5658 39078
rect 5602 39026 5604 39027
rect 5604 39026 5656 39027
rect 5656 39026 5658 39027
rect 5602 39014 5658 39026
rect 5602 38971 5604 39014
rect 5604 38971 5656 39014
rect 5656 38971 5658 39014
rect 5602 38898 5604 38947
rect 5604 38898 5656 38947
rect 5656 38898 5658 38947
rect 5602 38891 5658 38898
rect 5602 38834 5604 38867
rect 5604 38834 5656 38867
rect 5656 38834 5658 38867
rect 5602 38822 5658 38834
rect 5602 38811 5604 38822
rect 5604 38811 5656 38822
rect 5656 38811 5658 38822
rect 5602 38770 5604 38787
rect 5604 38770 5656 38787
rect 5656 38770 5658 38787
rect 5602 38758 5658 38770
rect 5602 38731 5604 38758
rect 5604 38731 5656 38758
rect 5656 38731 5658 38758
rect 5602 38706 5604 38707
rect 5604 38706 5656 38707
rect 5656 38706 5658 38707
rect 5602 38694 5658 38706
rect 5602 38651 5604 38694
rect 5604 38651 5656 38694
rect 5656 38651 5658 38694
rect 5602 38578 5604 38627
rect 5604 38578 5656 38627
rect 5656 38578 5658 38627
rect 5602 38571 5658 38578
rect 5602 38514 5604 38547
rect 5604 38514 5656 38547
rect 5656 38514 5658 38547
rect 5602 38502 5658 38514
rect 5602 38491 5604 38502
rect 5604 38491 5656 38502
rect 5656 38491 5658 38502
rect 5602 38450 5604 38467
rect 5604 38450 5656 38467
rect 5656 38450 5658 38467
rect 5602 38438 5658 38450
rect 5602 38411 5604 38438
rect 5604 38411 5656 38438
rect 5656 38411 5658 38438
rect 5602 38386 5604 38387
rect 5604 38386 5656 38387
rect 5656 38386 5658 38387
rect 5602 38374 5658 38386
rect 5602 38331 5604 38374
rect 5604 38331 5656 38374
rect 5656 38331 5658 38374
rect 5602 38258 5604 38307
rect 5604 38258 5656 38307
rect 5656 38258 5658 38307
rect 5602 38251 5658 38258
rect 5602 38194 5604 38227
rect 5604 38194 5656 38227
rect 5656 38194 5658 38227
rect 5602 38182 5658 38194
rect 5602 38171 5604 38182
rect 5604 38171 5656 38182
rect 5656 38171 5658 38182
rect 5602 38130 5604 38147
rect 5604 38130 5656 38147
rect 5656 38130 5658 38147
rect 5602 38118 5658 38130
rect 5602 38091 5604 38118
rect 5604 38091 5656 38118
rect 5656 38091 5658 38118
rect 5602 38066 5604 38067
rect 5604 38066 5656 38067
rect 5656 38066 5658 38067
rect 5602 38054 5658 38066
rect 5602 38011 5604 38054
rect 5604 38011 5656 38054
rect 5656 38011 5658 38054
rect 5602 37938 5604 37987
rect 5604 37938 5656 37987
rect 5656 37938 5658 37987
rect 5602 37931 5658 37938
rect 5602 37874 5604 37907
rect 5604 37874 5656 37907
rect 5656 37874 5658 37907
rect 5602 37862 5658 37874
rect 5602 37851 5604 37862
rect 5604 37851 5656 37862
rect 5656 37851 5658 37862
rect 5602 37810 5604 37827
rect 5604 37810 5656 37827
rect 5656 37810 5658 37827
rect 5602 37798 5658 37810
rect 5602 37771 5604 37798
rect 5604 37771 5656 37798
rect 5656 37771 5658 37798
rect 5602 37746 5604 37747
rect 5604 37746 5656 37747
rect 5656 37746 5658 37747
rect 5602 37734 5658 37746
rect 5602 37691 5604 37734
rect 5604 37691 5656 37734
rect 5656 37691 5658 37734
rect 5602 37618 5604 37667
rect 5604 37618 5656 37667
rect 5656 37618 5658 37667
rect 5602 37611 5658 37618
rect 5602 37554 5604 37587
rect 5604 37554 5656 37587
rect 5656 37554 5658 37587
rect 5602 37542 5658 37554
rect 5602 37531 5604 37542
rect 5604 37531 5656 37542
rect 5656 37531 5658 37542
rect 5602 37490 5604 37507
rect 5604 37490 5656 37507
rect 5656 37490 5658 37507
rect 5602 37478 5658 37490
rect 5602 37451 5604 37478
rect 5604 37451 5656 37478
rect 5656 37451 5658 37478
rect 5602 37426 5604 37427
rect 5604 37426 5656 37427
rect 5656 37426 5658 37427
rect 5602 37414 5658 37426
rect 5602 37371 5604 37414
rect 5604 37371 5656 37414
rect 5656 37371 5658 37414
rect 5602 37298 5604 37347
rect 5604 37298 5656 37347
rect 5656 37298 5658 37347
rect 5602 37291 5658 37298
rect 5602 37234 5604 37267
rect 5604 37234 5656 37267
rect 5656 37234 5658 37267
rect 5602 37222 5658 37234
rect 5602 37211 5604 37222
rect 5604 37211 5656 37222
rect 5656 37211 5658 37222
rect 5602 37170 5604 37187
rect 5604 37170 5656 37187
rect 5656 37170 5658 37187
rect 5602 37158 5658 37170
rect 5602 37131 5604 37158
rect 5604 37131 5656 37158
rect 5656 37131 5658 37158
rect 5602 37106 5604 37107
rect 5604 37106 5656 37107
rect 5656 37106 5658 37107
rect 5602 37094 5658 37106
rect 5602 37051 5604 37094
rect 5604 37051 5656 37094
rect 5656 37051 5658 37094
rect 5602 36978 5604 37027
rect 5604 36978 5656 37027
rect 5656 36978 5658 37027
rect 5602 36971 5658 36978
rect 5602 36914 5604 36947
rect 5604 36914 5656 36947
rect 5656 36914 5658 36947
rect 5602 36902 5658 36914
rect 5602 36891 5604 36902
rect 5604 36891 5656 36902
rect 5656 36891 5658 36902
rect 5602 36850 5604 36867
rect 5604 36850 5656 36867
rect 5656 36850 5658 36867
rect 5602 36838 5658 36850
rect 5602 36811 5604 36838
rect 5604 36811 5656 36838
rect 5656 36811 5658 36838
rect 5602 36786 5604 36787
rect 5604 36786 5656 36787
rect 5656 36786 5658 36787
rect 5602 36774 5658 36786
rect 5602 36731 5604 36774
rect 5604 36731 5656 36774
rect 5656 36731 5658 36774
rect 5602 36658 5604 36707
rect 5604 36658 5656 36707
rect 5656 36658 5658 36707
rect 5602 36651 5658 36658
rect 5602 36594 5604 36627
rect 5604 36594 5656 36627
rect 5656 36594 5658 36627
rect 5602 36582 5658 36594
rect 5602 36571 5604 36582
rect 5604 36571 5656 36582
rect 5656 36571 5658 36582
rect 5602 36530 5604 36547
rect 5604 36530 5656 36547
rect 5656 36530 5658 36547
rect 5602 36518 5658 36530
rect 5602 36491 5604 36518
rect 5604 36491 5656 36518
rect 5656 36491 5658 36518
rect 5602 36466 5604 36467
rect 5604 36466 5656 36467
rect 5656 36466 5658 36467
rect 5602 36454 5658 36466
rect 5602 36411 5604 36454
rect 5604 36411 5656 36454
rect 5656 36411 5658 36454
rect 5602 36338 5604 36387
rect 5604 36338 5656 36387
rect 5656 36338 5658 36387
rect 5602 36331 5658 36338
rect 5602 36274 5604 36307
rect 5604 36274 5656 36307
rect 5656 36274 5658 36307
rect 5602 36262 5658 36274
rect 5602 36251 5604 36262
rect 5604 36251 5656 36262
rect 5656 36251 5658 36262
rect 5602 36210 5604 36227
rect 5604 36210 5656 36227
rect 5656 36210 5658 36227
rect 5602 36198 5658 36210
rect 5602 36171 5604 36198
rect 5604 36171 5656 36198
rect 5656 36171 5658 36198
rect 5602 36146 5604 36147
rect 5604 36146 5656 36147
rect 5656 36146 5658 36147
rect 5602 36134 5658 36146
rect 5602 36091 5604 36134
rect 5604 36091 5656 36134
rect 5656 36091 5658 36134
rect 5602 36018 5604 36067
rect 5604 36018 5656 36067
rect 5656 36018 5658 36067
rect 5602 36011 5658 36018
rect 5602 35954 5604 35986
rect 5604 35954 5656 35986
rect 5656 35954 5658 35986
rect 5602 35942 5658 35954
rect 5602 35930 5604 35942
rect 5604 35930 5656 35942
rect 5656 35930 5658 35942
rect 5602 35890 5604 35905
rect 5604 35890 5656 35905
rect 5656 35890 5658 35905
rect 5602 35878 5658 35890
rect 5602 35849 5604 35878
rect 5604 35849 5656 35878
rect 5656 35849 5658 35878
rect 5602 35814 5658 35824
rect 5602 35768 5604 35814
rect 5604 35768 5656 35814
rect 5656 35768 5658 35814
rect 5602 35698 5604 35743
rect 5604 35698 5656 35743
rect 5656 35698 5658 35743
rect 5602 35687 5658 35698
rect 5602 35634 5604 35662
rect 5604 35634 5656 35662
rect 5656 35634 5658 35662
rect 5602 35622 5658 35634
rect 5602 35606 5604 35622
rect 5604 35606 5656 35622
rect 5656 35606 5658 35622
rect 5602 35570 5604 35581
rect 5604 35570 5656 35581
rect 5656 35570 5658 35581
rect 5602 35558 5658 35570
rect 5602 35525 5604 35558
rect 5604 35525 5656 35558
rect 5656 35525 5658 35558
rect 5602 35494 5658 35500
rect 5602 35444 5604 35494
rect 5604 35444 5656 35494
rect 5656 35444 5658 35494
rect 5602 35378 5604 35419
rect 5604 35378 5656 35419
rect 5656 35378 5658 35419
rect 5602 35366 5658 35378
rect 5602 35363 5604 35366
rect 5604 35363 5656 35366
rect 5656 35363 5658 35366
rect 5602 35314 5604 35338
rect 5604 35314 5656 35338
rect 5656 35314 5658 35338
rect 5602 35302 5658 35314
rect 5602 35282 5604 35302
rect 5604 35282 5656 35302
rect 5656 35282 5658 35302
rect 5602 35250 5604 35257
rect 5604 35250 5656 35257
rect 5656 35250 5658 35257
rect 5602 35238 5658 35250
rect 5602 35201 5604 35238
rect 5604 35201 5656 35238
rect 5656 35201 5658 35238
rect 5602 35174 5658 35176
rect 5602 35122 5604 35174
rect 5604 35122 5656 35174
rect 5656 35122 5658 35174
rect 5602 35120 5658 35122
rect 5602 35058 5604 35095
rect 5604 35058 5656 35095
rect 5656 35058 5658 35095
rect 5602 35046 5658 35058
rect 5602 35039 5604 35046
rect 5604 35039 5656 35046
rect 5656 35039 5658 35046
rect 5602 34994 5604 35014
rect 5604 34994 5656 35014
rect 5656 34994 5658 35014
rect 5602 34982 5658 34994
rect 5602 34958 5604 34982
rect 5604 34958 5656 34982
rect 5656 34958 5658 34982
rect 5602 34930 5604 34933
rect 5604 34930 5656 34933
rect 5656 34930 5658 34933
rect 5602 34918 5658 34930
rect 5602 34877 5604 34918
rect 5604 34877 5656 34918
rect 5656 34877 5658 34918
rect 5602 34802 5604 34852
rect 5604 34802 5656 34852
rect 5656 34802 5658 34852
rect 5602 34796 5658 34802
rect 5602 34738 5604 34771
rect 5604 34738 5656 34771
rect 5656 34738 5658 34771
rect 5602 34726 5658 34738
rect 5602 34715 5604 34726
rect 5604 34715 5656 34726
rect 5656 34715 5658 34726
rect 5602 34674 5604 34690
rect 5604 34674 5656 34690
rect 5656 34674 5658 34690
rect 5602 34662 5658 34674
rect 5602 34634 5604 34662
rect 5604 34634 5656 34662
rect 5656 34634 5658 34662
rect 5602 34598 5658 34609
rect 5602 34553 5604 34598
rect 5604 34553 5656 34598
rect 5656 34553 5658 34598
rect 5602 34482 5604 34528
rect 5604 34482 5656 34528
rect 5656 34482 5658 34528
rect 5602 34472 5658 34482
rect 5602 34418 5604 34447
rect 5604 34418 5656 34447
rect 5656 34418 5658 34447
rect 5602 34406 5658 34418
rect 5602 34391 5604 34406
rect 5604 34391 5656 34406
rect 5656 34391 5658 34406
rect 5602 34354 5604 34366
rect 5604 34354 5656 34366
rect 5656 34354 5658 34366
rect 5602 34342 5658 34354
rect 5602 34310 5604 34342
rect 5604 34310 5656 34342
rect 5656 34310 5658 34342
rect 5602 34278 5658 34285
rect 5602 34229 5604 34278
rect 5604 34229 5656 34278
rect 5656 34229 5658 34278
rect 5602 34162 5604 34204
rect 5604 34162 5656 34204
rect 5656 34162 5658 34204
rect 5602 34150 5658 34162
rect 5602 34148 5604 34150
rect 5604 34148 5656 34150
rect 5656 34148 5658 34150
rect 5602 34098 5604 34123
rect 5604 34098 5656 34123
rect 5656 34098 5658 34123
rect 5602 34086 5658 34098
rect 5602 34067 5604 34086
rect 5604 34067 5656 34086
rect 5656 34067 5658 34086
rect 5602 34034 5604 34042
rect 5604 34034 5656 34042
rect 5656 34034 5658 34042
rect 5602 34022 5658 34034
rect 5602 33986 5604 34022
rect 5604 33986 5656 34022
rect 5656 33986 5658 34022
rect 5602 33958 5658 33961
rect 5602 33906 5604 33958
rect 5604 33906 5656 33958
rect 5656 33906 5658 33958
rect 5602 33905 5658 33906
rect 5602 33842 5604 33880
rect 5604 33842 5656 33880
rect 5656 33842 5658 33880
rect 5602 33830 5658 33842
rect 5602 33824 5604 33830
rect 5604 33824 5656 33830
rect 5656 33824 5658 33830
rect 5602 33778 5604 33799
rect 5604 33778 5656 33799
rect 5656 33778 5658 33799
rect 5602 33766 5658 33778
rect 5602 33743 5604 33766
rect 5604 33743 5656 33766
rect 5656 33743 5658 33766
rect 5602 33714 5604 33718
rect 5604 33714 5656 33718
rect 5656 33714 5658 33718
rect 5602 33702 5658 33714
rect 5602 33662 5604 33702
rect 5604 33662 5656 33702
rect 5656 33662 5658 33702
rect 5602 33586 5604 33637
rect 5604 33586 5656 33637
rect 5656 33586 5658 33637
rect 5602 33581 5658 33586
rect 5602 33522 5604 33556
rect 5604 33522 5656 33556
rect 5656 33522 5658 33556
rect 5602 33510 5658 33522
rect 5602 33500 5604 33510
rect 5604 33500 5656 33510
rect 5656 33500 5658 33510
rect 5602 33458 5604 33475
rect 5604 33458 5656 33475
rect 5656 33458 5658 33475
rect 5602 33446 5658 33458
rect 5602 33419 5604 33446
rect 5604 33419 5656 33446
rect 5656 33419 5658 33446
rect 5602 33382 5658 33394
rect 5602 33338 5604 33382
rect 5604 33338 5656 33382
rect 5656 33338 5658 33382
rect 5602 33266 5604 33313
rect 5604 33266 5656 33313
rect 5656 33266 5658 33313
rect 5602 33257 5658 33266
rect 5602 33202 5604 33232
rect 5604 33202 5656 33232
rect 5656 33202 5658 33232
rect 5602 33190 5658 33202
rect 5602 33176 5604 33190
rect 5604 33176 5656 33190
rect 5656 33176 5658 33190
rect 5602 33138 5604 33151
rect 5604 33138 5656 33151
rect 5656 33138 5658 33151
rect 5602 33126 5658 33138
rect 5602 33095 5604 33126
rect 5604 33095 5656 33126
rect 5656 33095 5658 33126
rect 5602 33062 5658 33070
rect 5602 33014 5604 33062
rect 5604 33014 5656 33062
rect 5656 33014 5658 33062
rect 5602 32946 5604 32989
rect 5604 32946 5656 32989
rect 5656 32946 5658 32989
rect 5602 32934 5658 32946
rect 5602 32933 5604 32934
rect 5604 32933 5656 32934
rect 5656 32933 5658 32934
rect 5602 32882 5604 32908
rect 5604 32882 5656 32908
rect 5656 32882 5658 32908
rect 5602 32870 5658 32882
rect 5602 32852 5604 32870
rect 5604 32852 5656 32870
rect 5656 32852 5658 32870
rect 5602 32818 5604 32827
rect 5604 32818 5656 32827
rect 5656 32818 5658 32827
rect 5602 32806 5658 32818
rect 5602 32771 5604 32806
rect 5604 32771 5656 32806
rect 5656 32771 5658 32806
rect 5602 32742 5658 32746
rect 5602 32690 5604 32742
rect 5604 32690 5656 32742
rect 5656 32690 5658 32742
rect 5602 32625 5604 32665
rect 5604 32625 5656 32665
rect 5656 32625 5658 32665
rect 5602 32612 5658 32625
rect 5602 32609 5604 32612
rect 5604 32609 5656 32612
rect 5656 32609 5658 32612
rect 5602 32560 5604 32584
rect 5604 32560 5656 32584
rect 5656 32560 5658 32584
rect 5602 32547 5658 32560
rect 5602 32528 5604 32547
rect 5604 32528 5656 32547
rect 5656 32528 5658 32547
rect 5602 32495 5604 32503
rect 5604 32495 5656 32503
rect 5656 32495 5658 32503
rect 5602 32482 5658 32495
rect 5602 32447 5604 32482
rect 5604 32447 5656 32482
rect 5656 32447 5658 32482
rect 5602 32417 5658 32422
rect 5602 32366 5604 32417
rect 5604 32366 5656 32417
rect 5656 32366 5658 32417
rect 5602 32300 5604 32341
rect 5604 32300 5656 32341
rect 5656 32300 5658 32341
rect 5602 32287 5658 32300
rect 5602 32285 5604 32287
rect 5604 32285 5656 32287
rect 5656 32285 5658 32287
rect 5602 32235 5604 32260
rect 5604 32235 5656 32260
rect 5656 32235 5658 32260
rect 5602 32222 5658 32235
rect 5602 32204 5604 32222
rect 5604 32204 5656 32222
rect 5656 32204 5658 32222
rect 5602 32170 5604 32179
rect 5604 32170 5656 32179
rect 5656 32170 5658 32179
rect 5602 32157 5658 32170
rect 5602 32123 5604 32157
rect 5604 32123 5656 32157
rect 5656 32123 5658 32157
rect 5602 32092 5658 32098
rect 5602 32042 5604 32092
rect 5604 32042 5656 32092
rect 5656 32042 5658 32092
rect 5602 31975 5604 32017
rect 5604 31975 5656 32017
rect 5656 31975 5658 32017
rect 5602 31962 5658 31975
rect 5602 31961 5604 31962
rect 5604 31961 5656 31962
rect 5656 31961 5658 31962
rect 5602 31910 5604 31936
rect 5604 31910 5656 31936
rect 5656 31910 5658 31936
rect 5602 31897 5658 31910
rect 5602 31880 5604 31897
rect 5604 31880 5656 31897
rect 5656 31880 5658 31897
rect 5602 31845 5604 31855
rect 5604 31845 5656 31855
rect 5656 31845 5658 31855
rect 5602 31832 5658 31845
rect 5602 31799 5604 31832
rect 5604 31799 5656 31832
rect 5656 31799 5658 31832
rect 5602 31767 5658 31774
rect 5602 31718 5604 31767
rect 5604 31718 5656 31767
rect 5656 31718 5658 31767
rect 5602 31650 5604 31693
rect 5604 31650 5656 31693
rect 5656 31650 5658 31693
rect 5602 31637 5658 31650
rect 5602 31585 5604 31612
rect 5604 31585 5656 31612
rect 5656 31585 5658 31612
rect 5602 31572 5658 31585
rect 5602 31556 5604 31572
rect 5604 31556 5656 31572
rect 5656 31556 5658 31572
rect 5602 31520 5604 31531
rect 5604 31520 5656 31531
rect 5656 31520 5658 31531
rect 5602 31507 5658 31520
rect 5602 31475 5604 31507
rect 5604 31475 5656 31507
rect 5656 31475 5658 31507
rect 5602 31442 5658 31450
rect 5602 31394 5604 31442
rect 5604 31394 5656 31442
rect 5656 31394 5658 31442
rect 5602 31325 5604 31369
rect 5604 31325 5656 31369
rect 5656 31325 5658 31369
rect 5602 31313 5658 31325
rect 5602 31260 5604 31288
rect 5604 31260 5656 31288
rect 5656 31260 5658 31288
rect 5602 31247 5658 31260
rect 5602 31232 5604 31247
rect 5604 31232 5656 31247
rect 5656 31232 5658 31247
rect 5602 31195 5604 31207
rect 5604 31195 5656 31207
rect 5656 31195 5658 31207
rect 5602 31182 5658 31195
rect 5602 31151 5604 31182
rect 5604 31151 5656 31182
rect 5656 31151 5658 31182
rect 5602 31117 5658 31126
rect 5602 31070 5604 31117
rect 5604 31070 5656 31117
rect 5656 31070 5658 31117
rect 5602 31000 5604 31045
rect 5604 31000 5656 31045
rect 5656 31000 5658 31045
rect 5602 30989 5658 31000
rect 5602 30935 5604 30964
rect 5604 30935 5656 30964
rect 5656 30935 5658 30964
rect 5602 30922 5658 30935
rect 5602 30908 5604 30922
rect 5604 30908 5656 30922
rect 5656 30908 5658 30922
rect 5602 30870 5604 30883
rect 5604 30870 5656 30883
rect 5656 30870 5658 30883
rect 5602 30857 5658 30870
rect 5602 30827 5604 30857
rect 5604 30827 5656 30857
rect 5656 30827 5658 30857
rect 5602 30792 5658 30802
rect 5602 30746 5604 30792
rect 5604 30746 5656 30792
rect 5656 30746 5658 30792
rect 5602 30675 5604 30721
rect 5604 30675 5656 30721
rect 5656 30675 5658 30721
rect 5602 30665 5658 30675
rect 5602 30610 5604 30640
rect 5604 30610 5656 30640
rect 5656 30610 5658 30640
rect 5602 30597 5658 30610
rect 5602 30584 5604 30597
rect 5604 30584 5656 30597
rect 5656 30584 5658 30597
rect 5602 30545 5604 30559
rect 5604 30545 5656 30559
rect 5656 30545 5658 30559
rect 5602 30532 5658 30545
rect 5602 30503 5604 30532
rect 5604 30503 5656 30532
rect 5656 30503 5658 30532
rect 5602 30467 5658 30478
rect 5602 30422 5604 30467
rect 5604 30422 5656 30467
rect 5656 30422 5658 30467
rect 5602 30350 5604 30397
rect 5604 30350 5656 30397
rect 5656 30350 5658 30397
rect 5602 30341 5658 30350
rect 6742 27280 6798 27282
rect 6825 27280 6881 27282
rect 6908 27280 6964 27282
rect 6991 27280 7047 27282
rect 7074 27280 7130 27282
rect 7157 27280 7213 27282
rect 7240 27280 7296 27282
rect 7323 27280 7379 27282
rect 7406 27280 7462 27282
rect 7489 27280 7545 27282
rect 7571 27280 7627 27282
rect 7653 27280 7709 27282
rect 7735 27280 7791 27282
rect 6742 27228 6791 27280
rect 6791 27228 6798 27280
rect 6825 27228 6858 27280
rect 6858 27228 6873 27280
rect 6873 27228 6881 27280
rect 6908 27228 6925 27280
rect 6925 27228 6940 27280
rect 6940 27228 6964 27280
rect 6991 27228 6992 27280
rect 6992 27228 7007 27280
rect 7007 27228 7047 27280
rect 7074 27228 7126 27280
rect 7126 27228 7130 27280
rect 7157 27228 7193 27280
rect 7193 27228 7208 27280
rect 7208 27228 7213 27280
rect 7240 27228 7260 27280
rect 7260 27228 7275 27280
rect 7275 27228 7296 27280
rect 7323 27228 7327 27280
rect 7327 27228 7342 27280
rect 7342 27228 7379 27280
rect 7406 27228 7409 27280
rect 7409 27228 7461 27280
rect 7461 27228 7462 27280
rect 7489 27228 7528 27280
rect 7528 27228 7543 27280
rect 7543 27228 7545 27280
rect 7571 27228 7595 27280
rect 7595 27228 7610 27280
rect 7610 27228 7627 27280
rect 7653 27228 7662 27280
rect 7662 27228 7676 27280
rect 7676 27228 7709 27280
rect 7735 27228 7742 27280
rect 7742 27228 7791 27280
rect 6742 27226 6798 27228
rect 6825 27226 6881 27228
rect 6908 27226 6964 27228
rect 6991 27226 7047 27228
rect 7074 27226 7130 27228
rect 7157 27226 7213 27228
rect 7240 27226 7296 27228
rect 7323 27226 7379 27228
rect 7406 27226 7462 27228
rect 7489 27226 7545 27228
rect 7571 27226 7627 27228
rect 7653 27226 7709 27228
rect 7735 27226 7791 27228
rect 4672 27086 4721 27101
rect 4721 27086 4728 27101
rect 4757 27086 4788 27101
rect 4788 27086 4803 27101
rect 4803 27086 4813 27101
rect 4842 27086 4855 27101
rect 4855 27086 4870 27101
rect 4870 27086 4898 27101
rect 4926 27086 4937 27101
rect 4937 27086 4982 27101
rect 5010 27086 5056 27101
rect 5056 27086 5066 27101
rect 5094 27086 5123 27101
rect 5123 27086 5138 27101
rect 5138 27086 5150 27101
rect 5178 27086 5190 27101
rect 5190 27086 5205 27101
rect 5205 27086 5234 27101
rect 5262 27086 5272 27101
rect 5272 27086 5318 27101
rect 5346 27086 5391 27101
rect 5391 27086 5402 27101
rect 5430 27086 5458 27101
rect 5458 27086 5473 27101
rect 5473 27086 5486 27101
rect 5514 27086 5525 27101
rect 5525 27086 5539 27101
rect 5539 27086 5570 27101
rect 5598 27086 5605 27101
rect 5605 27086 5654 27101
rect 4672 27060 4728 27086
rect 4757 27060 4813 27086
rect 4842 27060 4898 27086
rect 4926 27060 4982 27086
rect 5010 27060 5066 27086
rect 5094 27060 5150 27086
rect 5178 27060 5234 27086
rect 5262 27060 5318 27086
rect 5346 27060 5402 27086
rect 5430 27060 5486 27086
rect 5514 27060 5570 27086
rect 5598 27060 5654 27086
rect 4672 27045 4721 27060
rect 4721 27045 4728 27060
rect 4757 27045 4788 27060
rect 4788 27045 4803 27060
rect 4803 27045 4813 27060
rect 4842 27045 4855 27060
rect 4855 27045 4870 27060
rect 4870 27045 4898 27060
rect 4926 27045 4937 27060
rect 4937 27045 4982 27060
rect 5010 27045 5056 27060
rect 5056 27045 5066 27060
rect 5094 27045 5123 27060
rect 5123 27045 5138 27060
rect 5138 27045 5150 27060
rect 5178 27045 5190 27060
rect 5190 27045 5205 27060
rect 5205 27045 5234 27060
rect 5262 27045 5272 27060
rect 5272 27045 5318 27060
rect 5346 27045 5391 27060
rect 5391 27045 5402 27060
rect 5430 27045 5458 27060
rect 5458 27045 5473 27060
rect 5473 27045 5486 27060
rect 5514 27045 5525 27060
rect 5525 27045 5539 27060
rect 5539 27045 5570 27060
rect 5598 27045 5605 27060
rect 5605 27045 5654 27060
rect 6086 22131 6142 22133
rect 6166 22131 6222 22133
rect 6086 22079 6135 22131
rect 6135 22079 6142 22131
rect 6166 22079 6199 22131
rect 6199 22079 6222 22131
rect 6086 22077 6142 22079
rect 6166 22077 6222 22079
rect 5110 7710 5166 7727
rect 5192 7710 5248 7727
rect 5274 7710 5330 7727
rect 5110 7671 5136 7710
rect 5136 7671 5155 7710
rect 5155 7671 5166 7710
rect 5192 7671 5207 7710
rect 5207 7671 5226 7710
rect 5226 7671 5248 7710
rect 5274 7671 5278 7710
rect 5278 7671 5330 7710
rect 5355 7671 5411 7727
rect 5436 7671 5492 7727
rect 5517 7671 5573 7727
rect 5598 7719 5654 7727
rect 5598 7671 5649 7719
rect 5649 7671 5654 7719
rect 5110 7584 5136 7631
rect 5136 7584 5155 7631
rect 5155 7584 5166 7631
rect 5192 7584 5207 7631
rect 5207 7584 5226 7631
rect 5226 7584 5248 7631
rect 5274 7584 5278 7631
rect 5278 7584 5330 7631
rect 5110 7575 5166 7584
rect 5192 7575 5248 7584
rect 5274 7575 5330 7584
rect 5355 7575 5411 7631
rect 5436 7575 5492 7631
rect 5517 7575 5573 7631
rect 5598 7592 5649 7631
rect 5649 7592 5654 7631
rect 5598 7575 5654 7592
rect 5110 7510 5136 7535
rect 5136 7510 5155 7535
rect 5155 7510 5166 7535
rect 5192 7510 5207 7535
rect 5207 7510 5226 7535
rect 5226 7510 5248 7535
rect 5274 7510 5278 7535
rect 5278 7510 5330 7535
rect 5110 7488 5166 7510
rect 5192 7488 5248 7510
rect 5274 7488 5330 7510
rect 5110 7479 5136 7488
rect 5136 7479 5155 7488
rect 5155 7479 5166 7488
rect 5192 7479 5207 7488
rect 5207 7479 5226 7488
rect 5226 7479 5248 7488
rect 5274 7479 5278 7488
rect 5278 7479 5330 7488
rect 5355 7479 5411 7535
rect 5436 7479 5492 7535
rect 5517 7479 5573 7535
rect 5598 7517 5649 7535
rect 5649 7517 5654 7535
rect 5598 7494 5654 7517
rect 5598 7479 5649 7494
rect 5649 7479 5654 7494
rect 5110 7436 5136 7439
rect 5136 7436 5155 7439
rect 5155 7436 5166 7439
rect 5192 7436 5207 7439
rect 5207 7436 5226 7439
rect 5226 7436 5248 7439
rect 5274 7436 5278 7439
rect 5278 7436 5330 7439
rect 5110 7414 5166 7436
rect 5192 7414 5248 7436
rect 5274 7414 5330 7436
rect 5110 7383 5136 7414
rect 5136 7383 5155 7414
rect 5155 7383 5166 7414
rect 5192 7383 5207 7414
rect 5207 7383 5226 7414
rect 5226 7383 5248 7414
rect 5274 7383 5278 7414
rect 5278 7383 5330 7414
rect 5355 7383 5411 7439
rect 5436 7383 5492 7439
rect 5517 7383 5573 7439
rect 5598 7419 5654 7439
rect 5598 7383 5649 7419
rect 5649 7383 5654 7419
rect 5110 7340 5166 7343
rect 5192 7340 5248 7343
rect 5274 7340 5330 7343
rect 5110 7288 5136 7340
rect 5136 7288 5155 7340
rect 5155 7288 5166 7340
rect 5192 7288 5207 7340
rect 5207 7288 5226 7340
rect 5226 7288 5248 7340
rect 5274 7288 5278 7340
rect 5278 7288 5330 7340
rect 5110 7287 5166 7288
rect 5192 7287 5248 7288
rect 5274 7287 5330 7288
rect 5355 7287 5411 7343
rect 5436 7287 5492 7343
rect 5517 7287 5573 7343
rect 5598 7292 5649 7343
rect 5649 7292 5654 7343
rect 5598 7287 5654 7292
rect 5874 4989 5926 5038
rect 5926 4989 5930 5038
rect 5958 4989 5994 5038
rect 5994 4989 6010 5038
rect 6010 4989 6014 5038
rect 6042 4989 6062 5038
rect 6062 4989 6078 5038
rect 6078 4989 6098 5038
rect 6126 4989 6130 5038
rect 6130 4989 6146 5038
rect 6146 4989 6182 5038
rect 6210 4989 6214 5038
rect 6214 4989 6266 5038
rect 5874 4982 5930 4989
rect 5958 4982 6014 4989
rect 6042 4982 6098 4989
rect 6126 4982 6182 4989
rect 6210 4982 6266 4989
rect 5874 4919 5926 4958
rect 5926 4919 5930 4958
rect 5958 4919 5994 4958
rect 5994 4919 6010 4958
rect 6010 4919 6014 4958
rect 6042 4919 6062 4958
rect 6062 4919 6078 4958
rect 6078 4919 6098 4958
rect 6126 4919 6130 4958
rect 6130 4919 6146 4958
rect 6146 4919 6182 4958
rect 6210 4919 6214 4958
rect 6214 4919 6266 4958
rect 5874 4902 5930 4919
rect 5958 4902 6014 4919
rect 6042 4902 6098 4919
rect 6126 4902 6182 4919
rect 6210 4902 6266 4919
rect 5874 4849 5926 4878
rect 5926 4849 5930 4878
rect 5958 4849 5994 4878
rect 5994 4849 6010 4878
rect 6010 4849 6014 4878
rect 6042 4849 6062 4878
rect 6062 4849 6078 4878
rect 6078 4849 6098 4878
rect 6126 4849 6130 4878
rect 6130 4849 6146 4878
rect 6146 4849 6182 4878
rect 6210 4849 6214 4878
rect 6214 4849 6266 4878
rect 5874 4831 5930 4849
rect 5958 4831 6014 4849
rect 6042 4831 6098 4849
rect 6126 4831 6182 4849
rect 6210 4831 6266 4849
rect 5874 4822 5926 4831
rect 5926 4822 5930 4831
rect 5958 4822 5994 4831
rect 5994 4822 6010 4831
rect 6010 4822 6014 4831
rect 6042 4822 6062 4831
rect 6062 4822 6078 4831
rect 6078 4822 6098 4831
rect 6126 4822 6130 4831
rect 6130 4822 6146 4831
rect 6146 4822 6182 4831
rect 6210 4822 6214 4831
rect 6214 4822 6266 4831
rect 5874 4779 5926 4798
rect 5926 4779 5930 4798
rect 5958 4779 5994 4798
rect 5994 4779 6010 4798
rect 6010 4779 6014 4798
rect 6042 4779 6062 4798
rect 6062 4779 6078 4798
rect 6078 4779 6098 4798
rect 6126 4779 6130 4798
rect 6130 4779 6146 4798
rect 6146 4779 6182 4798
rect 6210 4779 6214 4798
rect 6214 4779 6266 4798
rect 5874 4761 5930 4779
rect 5958 4761 6014 4779
rect 6042 4761 6098 4779
rect 6126 4761 6182 4779
rect 6210 4761 6266 4779
rect 5874 4742 5926 4761
rect 5926 4742 5930 4761
rect 5958 4742 5994 4761
rect 5994 4742 6010 4761
rect 6010 4742 6014 4761
rect 6042 4742 6062 4761
rect 6062 4742 6078 4761
rect 6078 4742 6098 4761
rect 6126 4742 6130 4761
rect 6130 4742 6146 4761
rect 6146 4742 6182 4761
rect 6210 4742 6214 4761
rect 6214 4742 6266 4761
rect 5874 4709 5926 4718
rect 5926 4709 5930 4718
rect 5958 4709 5994 4718
rect 5994 4709 6010 4718
rect 6010 4709 6014 4718
rect 6042 4709 6062 4718
rect 6062 4709 6078 4718
rect 6078 4709 6098 4718
rect 6126 4709 6130 4718
rect 6130 4709 6146 4718
rect 6146 4709 6182 4718
rect 6210 4709 6214 4718
rect 6214 4709 6266 4718
rect 5874 4691 5930 4709
rect 5958 4691 6014 4709
rect 6042 4691 6098 4709
rect 6126 4691 6182 4709
rect 6210 4691 6266 4709
rect 5874 4662 5926 4691
rect 5926 4662 5930 4691
rect 5958 4662 5994 4691
rect 5994 4662 6010 4691
rect 6010 4662 6014 4691
rect 6042 4662 6062 4691
rect 6062 4662 6078 4691
rect 6078 4662 6098 4691
rect 6126 4662 6130 4691
rect 6130 4662 6146 4691
rect 6146 4662 6182 4691
rect 6210 4662 6214 4691
rect 6214 4662 6266 4691
rect 5874 4620 5930 4638
rect 5958 4620 6014 4638
rect 6042 4620 6098 4638
rect 6126 4620 6182 4638
rect 6210 4620 6266 4638
rect 5874 4582 5926 4620
rect 5926 4582 5930 4620
rect 5958 4582 5994 4620
rect 5994 4582 6010 4620
rect 6010 4582 6014 4620
rect 6042 4582 6062 4620
rect 6062 4582 6078 4620
rect 6078 4582 6098 4620
rect 6126 4582 6130 4620
rect 6130 4582 6146 4620
rect 6146 4582 6182 4620
rect 6210 4582 6214 4620
rect 6214 4582 6266 4620
rect 5874 4549 5930 4557
rect 5958 4549 6014 4557
rect 6042 4549 6098 4557
rect 6126 4549 6182 4557
rect 6210 4549 6266 4557
rect 5874 4501 5926 4549
rect 5926 4501 5930 4549
rect 5958 4501 5994 4549
rect 5994 4501 6010 4549
rect 6010 4501 6014 4549
rect 6042 4501 6062 4549
rect 6062 4501 6078 4549
rect 6078 4501 6098 4549
rect 6126 4501 6130 4549
rect 6130 4501 6146 4549
rect 6146 4501 6182 4549
rect 6210 4501 6214 4549
rect 6214 4501 6266 4549
rect 5874 4420 5930 4476
rect 5958 4420 6014 4476
rect 6042 4420 6098 4476
rect 6126 4420 6182 4476
rect 6210 4420 6266 4476
rect 5874 4339 5930 4395
rect 5958 4339 6014 4395
rect 6042 4339 6098 4395
rect 6126 4339 6182 4395
rect 6210 4339 6266 4395
rect 5874 4258 5930 4314
rect 5958 4258 6014 4314
rect 6042 4258 6098 4314
rect 6126 4258 6182 4314
rect 6210 4258 6266 4314
rect 5874 4177 5930 4233
rect 5958 4177 6014 4233
rect 6042 4177 6098 4233
rect 6126 4177 6182 4233
rect 6210 4177 6266 4233
rect 5874 4096 5930 4152
rect 5958 4096 6014 4152
rect 6042 4096 6098 4152
rect 6126 4096 6182 4152
rect 6210 4096 6266 4152
rect 5874 4015 5930 4071
rect 5958 4015 6014 4071
rect 6042 4015 6098 4071
rect 6126 4015 6182 4071
rect 6210 4015 6266 4071
rect 5874 3967 5930 3990
rect 5958 3967 6014 3990
rect 5874 3934 5879 3967
rect 5879 3934 5930 3967
rect 5958 3934 5962 3967
rect 5962 3934 6014 3967
rect 6042 3967 6098 3990
rect 6042 3934 6045 3967
rect 6045 3934 6097 3967
rect 6097 3934 6098 3967
rect 6126 3967 6182 3990
rect 6210 3967 6266 3990
rect 6126 3934 6127 3967
rect 6127 3934 6179 3967
rect 6179 3934 6182 3967
rect 6210 3934 6261 3967
rect 6261 3934 6266 3967
rect 5874 3891 5930 3909
rect 5958 3891 6014 3909
rect 5874 3853 5879 3891
rect 5879 3853 5930 3891
rect 5958 3853 5962 3891
rect 5962 3853 6014 3891
rect 6042 3891 6098 3909
rect 6042 3853 6045 3891
rect 6045 3853 6097 3891
rect 6097 3853 6098 3891
rect 6126 3891 6182 3909
rect 6210 3891 6266 3909
rect 6126 3853 6127 3891
rect 6127 3853 6179 3891
rect 6179 3853 6182 3891
rect 6210 3853 6261 3891
rect 6261 3853 6266 3891
rect 5874 3815 5930 3828
rect 5958 3815 6014 3828
rect 5874 3772 5879 3815
rect 5879 3772 5930 3815
rect 5958 3772 5962 3815
rect 5962 3772 6014 3815
rect 6042 3815 6098 3828
rect 6042 3772 6045 3815
rect 6045 3772 6097 3815
rect 6097 3772 6098 3815
rect 6126 3815 6182 3828
rect 6210 3815 6266 3828
rect 6126 3772 6127 3815
rect 6127 3772 6179 3815
rect 6179 3772 6182 3815
rect 6210 3772 6261 3815
rect 6261 3772 6266 3815
rect 5832 3428 5888 3484
rect 5953 3428 6009 3484
rect 6074 3428 6130 3484
rect 6195 3428 6251 3484
rect 6316 3428 6372 3484
rect 6437 3428 6493 3484
rect 6558 3428 6614 3484
<< metal3 >>
rect 4663 39267 5663 40000
rect 4663 39211 5602 39267
rect 5658 39211 5663 39267
rect 4663 39187 5663 39211
rect 4663 39131 5602 39187
rect 5658 39131 5663 39187
rect 4663 39107 5663 39131
rect 4663 39051 5602 39107
rect 5658 39051 5663 39107
rect 4663 39027 5663 39051
rect 4663 38971 5602 39027
rect 5658 38971 5663 39027
rect 4663 38947 5663 38971
rect 4663 38891 5602 38947
rect 5658 38891 5663 38947
rect 4663 38867 5663 38891
rect 4663 38811 5602 38867
rect 5658 38811 5663 38867
rect 4663 38787 5663 38811
rect 4663 38731 5602 38787
rect 5658 38731 5663 38787
rect 4663 38707 5663 38731
rect 4663 38651 5602 38707
rect 5658 38651 5663 38707
rect 4663 38627 5663 38651
rect 4663 38571 5602 38627
rect 5658 38571 5663 38627
rect 4663 38547 5663 38571
rect 4663 38491 5602 38547
rect 5658 38491 5663 38547
rect 4663 38467 5663 38491
rect 4663 38411 5602 38467
rect 5658 38411 5663 38467
rect 4663 38387 5663 38411
rect 4663 38331 5602 38387
rect 5658 38331 5663 38387
rect 4663 38307 5663 38331
rect 4663 38251 5602 38307
rect 5658 38251 5663 38307
rect 4663 38227 5663 38251
rect 4663 38171 5602 38227
rect 5658 38171 5663 38227
rect 4663 38147 5663 38171
rect 4663 38091 5602 38147
rect 5658 38091 5663 38147
rect 4663 38067 5663 38091
rect 4663 38011 5602 38067
rect 5658 38011 5663 38067
rect 4663 37987 5663 38011
rect 4663 37931 5602 37987
rect 5658 37931 5663 37987
rect 4663 37907 5663 37931
rect 4663 37851 5602 37907
rect 5658 37851 5663 37907
rect 4663 37827 5663 37851
rect 4663 37771 5602 37827
rect 5658 37771 5663 37827
rect 4663 37747 5663 37771
rect 4663 37691 5602 37747
rect 5658 37691 5663 37747
rect 4663 37667 5663 37691
rect 4663 37611 5602 37667
rect 5658 37611 5663 37667
rect 4663 37587 5663 37611
rect 4663 37531 5602 37587
rect 5658 37531 5663 37587
rect 4663 37507 5663 37531
rect 4663 37451 5602 37507
rect 5658 37451 5663 37507
rect 4663 37427 5663 37451
rect 4663 37371 5602 37427
rect 5658 37371 5663 37427
rect 4663 37347 5663 37371
rect 4663 37291 5602 37347
rect 5658 37291 5663 37347
rect 4663 37267 5663 37291
rect 4663 37211 5602 37267
rect 5658 37211 5663 37267
rect 4663 37187 5663 37211
rect 4663 37131 5602 37187
rect 5658 37131 5663 37187
rect 4663 37107 5663 37131
rect 4663 37051 5602 37107
rect 5658 37051 5663 37107
rect 4663 37027 5663 37051
rect 4663 36971 5602 37027
rect 5658 36971 5663 37027
rect 4663 36947 5663 36971
rect 4663 36891 5602 36947
rect 5658 36891 5663 36947
rect 4663 36867 5663 36891
rect 4663 36811 5602 36867
rect 5658 36811 5663 36867
rect 4663 36787 5663 36811
rect 4663 36731 5602 36787
rect 5658 36731 5663 36787
rect 4663 36707 5663 36731
rect 4663 36651 5602 36707
rect 5658 36651 5663 36707
rect 4663 36627 5663 36651
rect 4663 36571 5602 36627
rect 5658 36571 5663 36627
rect 4663 36547 5663 36571
rect 4663 36491 5602 36547
rect 5658 36491 5663 36547
rect 4663 36467 5663 36491
rect 4663 36411 5602 36467
rect 5658 36411 5663 36467
rect 4663 36387 5663 36411
rect 4663 36331 5602 36387
rect 5658 36331 5663 36387
rect 4663 36307 5663 36331
rect 4663 36251 5602 36307
rect 5658 36251 5663 36307
rect 4663 36227 5663 36251
rect 4663 36171 5602 36227
rect 5658 36171 5663 36227
rect 4663 36147 5663 36171
rect 4663 36091 5602 36147
rect 5658 36091 5663 36147
rect 4663 36067 5663 36091
rect 4663 36011 5602 36067
rect 5658 36011 5663 36067
rect 4663 35986 5663 36011
rect 4663 35930 5602 35986
rect 5658 35930 5663 35986
rect 4663 35905 5663 35930
rect 4663 35849 5602 35905
rect 5658 35849 5663 35905
rect 4663 35824 5663 35849
rect 4663 35768 5602 35824
rect 5658 35768 5663 35824
rect 4663 35743 5663 35768
rect 4663 35687 5602 35743
rect 5658 35687 5663 35743
rect 4663 35662 5663 35687
rect 4663 35606 5602 35662
rect 5658 35606 5663 35662
rect 4663 35581 5663 35606
rect 4663 35525 5602 35581
rect 5658 35525 5663 35581
rect 4663 35500 5663 35525
rect 4663 35444 5602 35500
rect 5658 35444 5663 35500
rect 4663 35419 5663 35444
rect 4663 35363 5602 35419
rect 5658 35363 5663 35419
rect 4663 35338 5663 35363
rect 4663 35282 5602 35338
rect 5658 35282 5663 35338
rect 4663 35257 5663 35282
rect 4663 35201 5602 35257
rect 5658 35201 5663 35257
rect 4663 35176 5663 35201
rect 4663 35120 5602 35176
rect 5658 35120 5663 35176
rect 4663 35095 5663 35120
rect 4663 35039 5602 35095
rect 5658 35039 5663 35095
rect 4663 35014 5663 35039
rect 4663 34958 5602 35014
rect 5658 34958 5663 35014
rect 4663 34933 5663 34958
rect 4663 34877 5602 34933
rect 5658 34877 5663 34933
rect 4663 34852 5663 34877
rect 4663 34796 5602 34852
rect 5658 34796 5663 34852
rect 4663 34771 5663 34796
rect 4663 34715 5602 34771
rect 5658 34715 5663 34771
rect 4663 34690 5663 34715
rect 4663 34634 5602 34690
rect 5658 34634 5663 34690
rect 4663 34609 5663 34634
rect 4663 34553 5602 34609
rect 5658 34553 5663 34609
rect 4663 34528 5663 34553
rect 4663 34472 5602 34528
rect 5658 34472 5663 34528
rect 4663 34447 5663 34472
rect 4663 34391 5602 34447
rect 5658 34391 5663 34447
rect 4663 34366 5663 34391
rect 4663 34310 5602 34366
rect 5658 34310 5663 34366
rect 4663 34285 5663 34310
rect 4663 34229 5602 34285
rect 5658 34229 5663 34285
rect 4663 34204 5663 34229
rect 4663 34148 5602 34204
rect 5658 34148 5663 34204
rect 4663 34123 5663 34148
rect 4663 34067 5602 34123
rect 5658 34067 5663 34123
rect 4663 34042 5663 34067
rect 4663 33986 5602 34042
rect 5658 33986 5663 34042
rect 4663 33961 5663 33986
rect 4663 33905 5602 33961
rect 5658 33905 5663 33961
rect 4663 33880 5663 33905
rect 4663 33824 5602 33880
rect 5658 33824 5663 33880
rect 4663 33799 5663 33824
rect 4663 33743 5602 33799
rect 5658 33743 5663 33799
rect 4663 33718 5663 33743
rect 4663 33662 5602 33718
rect 5658 33662 5663 33718
rect 4663 33637 5663 33662
rect 4663 33581 5602 33637
rect 5658 33581 5663 33637
rect 4663 33556 5663 33581
rect 4663 33500 5602 33556
rect 5658 33500 5663 33556
rect 4663 33475 5663 33500
rect 4663 33419 5602 33475
rect 5658 33419 5663 33475
rect 4663 33394 5663 33419
rect 4663 33338 5602 33394
rect 5658 33338 5663 33394
rect 4663 33313 5663 33338
rect 4663 33257 5602 33313
rect 5658 33257 5663 33313
rect 4663 33232 5663 33257
rect 4663 33176 5602 33232
rect 5658 33176 5663 33232
rect 4663 33151 5663 33176
rect 4663 33095 5602 33151
rect 5658 33095 5663 33151
rect 4663 33070 5663 33095
rect 4663 33014 5602 33070
rect 5658 33014 5663 33070
rect 4663 32989 5663 33014
rect 4663 32933 5602 32989
rect 5658 32933 5663 32989
rect 4663 32908 5663 32933
rect 4663 32852 5602 32908
rect 5658 32852 5663 32908
rect 4663 32827 5663 32852
rect 4663 32771 5602 32827
rect 5658 32771 5663 32827
rect 4663 32746 5663 32771
rect 4663 32690 5602 32746
rect 5658 32690 5663 32746
rect 4663 32665 5663 32690
rect 4663 32609 5602 32665
rect 5658 32609 5663 32665
rect 4663 32584 5663 32609
rect 4663 32528 5602 32584
rect 5658 32528 5663 32584
rect 4663 32503 5663 32528
rect 4663 32447 5602 32503
rect 5658 32447 5663 32503
rect 4663 32422 5663 32447
rect 4663 32366 5602 32422
rect 5658 32366 5663 32422
rect 4663 32341 5663 32366
rect 4663 32285 5602 32341
rect 5658 32285 5663 32341
rect 4663 32260 5663 32285
rect 4663 32204 5602 32260
rect 5658 32204 5663 32260
rect 4663 32179 5663 32204
rect 4663 32123 5602 32179
rect 5658 32123 5663 32179
rect 4663 32098 5663 32123
rect 4663 32042 5602 32098
rect 5658 32042 5663 32098
rect 4663 32017 5663 32042
rect 4663 31961 5602 32017
rect 5658 31961 5663 32017
rect 4663 31936 5663 31961
rect 4663 31880 5602 31936
rect 5658 31880 5663 31936
rect 4663 31855 5663 31880
rect 4663 31799 5602 31855
rect 5658 31799 5663 31855
rect 4663 31774 5663 31799
rect 4663 31718 5602 31774
rect 5658 31718 5663 31774
rect 4663 31693 5663 31718
rect 4663 31637 5602 31693
rect 5658 31637 5663 31693
rect 4663 31612 5663 31637
rect 4663 31556 5602 31612
rect 5658 31556 5663 31612
rect 4663 31531 5663 31556
rect 4663 31475 5602 31531
rect 5658 31475 5663 31531
rect 4663 31450 5663 31475
rect 4663 31394 5602 31450
rect 5658 31394 5663 31450
rect 4663 31369 5663 31394
rect 4663 31313 5602 31369
rect 5658 31313 5663 31369
rect 4663 31288 5663 31313
rect 4663 31232 5602 31288
rect 5658 31232 5663 31288
rect 4663 31207 5663 31232
rect 4663 31151 5602 31207
rect 5658 31151 5663 31207
rect 4663 31126 5663 31151
rect 4663 31070 5602 31126
rect 5658 31070 5663 31126
rect 4663 31045 5663 31070
rect 4663 30989 5602 31045
rect 5658 30989 5663 31045
rect 4663 30964 5663 30989
rect 4663 30908 5602 30964
rect 5658 30908 5663 30964
rect 4663 30883 5663 30908
rect 4663 30827 5602 30883
rect 5658 30827 5663 30883
rect 4663 30802 5663 30827
rect 4663 30746 5602 30802
rect 5658 30746 5663 30802
rect 4663 30721 5663 30746
rect 4663 30665 5602 30721
rect 5658 30665 5663 30721
rect 4663 30640 5663 30665
rect 4663 30584 5602 30640
rect 5658 30584 5663 30640
rect 4663 30559 5663 30584
rect 4663 30503 5602 30559
rect 5658 30503 5663 30559
rect 4663 30478 5663 30503
rect 4663 30422 5602 30478
rect 5658 30422 5663 30478
rect 4663 30397 5663 30422
rect 4663 30341 5602 30397
rect 5658 30341 5663 30397
rect 4663 27101 5663 30341
rect 4663 27045 4672 27101
rect 4728 27045 4757 27101
rect 4813 27045 4842 27101
rect 4898 27045 4926 27101
rect 4982 27045 5010 27101
rect 5066 27045 5094 27101
rect 5150 27045 5178 27101
rect 5234 27045 5262 27101
rect 5318 27045 5346 27101
rect 5402 27045 5430 27101
rect 5486 27045 5514 27101
rect 5570 27045 5598 27101
rect 5654 27045 5663 27101
rect 4663 7727 5663 27045
rect 4663 7671 5110 7727
rect 5166 7671 5192 7727
rect 5248 7671 5274 7727
rect 5330 7671 5355 7727
rect 5411 7671 5436 7727
rect 5492 7671 5517 7727
rect 5573 7671 5598 7727
rect 5654 7671 5663 7727
rect 4663 7631 5663 7671
rect 4663 7575 5110 7631
rect 5166 7575 5192 7631
rect 5248 7575 5274 7631
rect 5330 7575 5355 7631
rect 5411 7575 5436 7631
rect 5492 7575 5517 7631
rect 5573 7575 5598 7631
rect 5654 7575 5663 7631
rect 4663 7535 5663 7575
rect 4663 7479 5110 7535
rect 5166 7479 5192 7535
rect 5248 7479 5274 7535
rect 5330 7479 5355 7535
rect 5411 7479 5436 7535
rect 5492 7479 5517 7535
rect 5573 7479 5598 7535
rect 5654 7479 5663 7535
rect 4663 7439 5663 7479
rect 4663 7383 5110 7439
rect 5166 7383 5192 7439
rect 5248 7383 5274 7439
rect 5330 7383 5355 7439
rect 5411 7383 5436 7439
rect 5492 7383 5517 7439
rect 5573 7383 5598 7439
rect 5654 7383 5663 7439
rect 4663 7343 5663 7383
rect 4663 7287 5110 7343
rect 5166 7287 5192 7343
rect 5248 7287 5274 7343
rect 5330 7287 5355 7343
rect 5411 7287 5436 7343
rect 5492 7287 5517 7343
rect 5573 7287 5598 7343
rect 5654 7287 5663 7343
rect 4663 14 5663 7287
rect 5823 22133 6623 40000
rect 6737 27282 7796 27287
rect 6737 27226 6742 27282
rect 6798 27226 6825 27282
rect 6881 27226 6908 27282
rect 6964 27226 6991 27282
rect 7047 27226 7074 27282
rect 7130 27226 7157 27282
rect 7213 27226 7240 27282
rect 7296 27226 7323 27282
rect 7379 27226 7406 27282
rect 7462 27226 7489 27282
rect 7545 27226 7571 27282
rect 7627 27226 7653 27282
rect 7709 27226 7735 27282
rect 7791 27226 7796 27282
rect 6737 27221 7796 27226
rect 5823 22077 6086 22133
rect 6142 22077 6166 22133
rect 6222 22077 6623 22133
rect 5823 5038 6623 22077
rect 5823 4982 5874 5038
rect 5930 4982 5958 5038
rect 6014 4982 6042 5038
rect 6098 4982 6126 5038
rect 6182 4982 6210 5038
rect 6266 4982 6623 5038
rect 5823 4958 6623 4982
rect 5823 4902 5874 4958
rect 5930 4902 5958 4958
rect 6014 4902 6042 4958
rect 6098 4902 6126 4958
rect 6182 4902 6210 4958
rect 6266 4902 6623 4958
rect 5823 4878 6623 4902
rect 5823 4822 5874 4878
rect 5930 4822 5958 4878
rect 6014 4822 6042 4878
rect 6098 4822 6126 4878
rect 6182 4822 6210 4878
rect 6266 4822 6623 4878
rect 5823 4798 6623 4822
rect 5823 4742 5874 4798
rect 5930 4742 5958 4798
rect 6014 4742 6042 4798
rect 6098 4742 6126 4798
rect 6182 4742 6210 4798
rect 6266 4742 6623 4798
rect 5823 4718 6623 4742
rect 5823 4662 5874 4718
rect 5930 4662 5958 4718
rect 6014 4662 6042 4718
rect 6098 4662 6126 4718
rect 6182 4662 6210 4718
rect 6266 4662 6623 4718
rect 5823 4638 6623 4662
rect 5823 4582 5874 4638
rect 5930 4582 5958 4638
rect 6014 4582 6042 4638
rect 6098 4582 6126 4638
rect 6182 4582 6210 4638
rect 6266 4582 6623 4638
rect 5823 4557 6623 4582
rect 5823 4501 5874 4557
rect 5930 4501 5958 4557
rect 6014 4501 6042 4557
rect 6098 4501 6126 4557
rect 6182 4501 6210 4557
rect 6266 4501 6623 4557
rect 5823 4476 6623 4501
rect 5823 4420 5874 4476
rect 5930 4420 5958 4476
rect 6014 4420 6042 4476
rect 6098 4420 6126 4476
rect 6182 4420 6210 4476
rect 6266 4420 6623 4476
rect 5823 4395 6623 4420
rect 5823 4339 5874 4395
rect 5930 4339 5958 4395
rect 6014 4339 6042 4395
rect 6098 4339 6126 4395
rect 6182 4339 6210 4395
rect 6266 4339 6623 4395
rect 5823 4314 6623 4339
rect 5823 4258 5874 4314
rect 5930 4258 5958 4314
rect 6014 4258 6042 4314
rect 6098 4258 6126 4314
rect 6182 4258 6210 4314
rect 6266 4258 6623 4314
rect 5823 4233 6623 4258
rect 5823 4177 5874 4233
rect 5930 4177 5958 4233
rect 6014 4177 6042 4233
rect 6098 4177 6126 4233
rect 6182 4177 6210 4233
rect 6266 4177 6623 4233
rect 5823 4152 6623 4177
rect 5823 4096 5874 4152
rect 5930 4096 5958 4152
rect 6014 4096 6042 4152
rect 6098 4096 6126 4152
rect 6182 4096 6210 4152
rect 6266 4096 6623 4152
rect 5823 4071 6623 4096
rect 5823 4015 5874 4071
rect 5930 4015 5958 4071
rect 6014 4015 6042 4071
rect 6098 4015 6126 4071
rect 6182 4015 6210 4071
rect 6266 4015 6623 4071
rect 5823 3990 6623 4015
rect 5823 3934 5874 3990
rect 5930 3934 5958 3990
rect 6014 3934 6042 3990
rect 6098 3934 6126 3990
rect 6182 3934 6210 3990
rect 6266 3934 6623 3990
rect 5823 3909 6623 3934
rect 5823 3853 5874 3909
rect 5930 3853 5958 3909
rect 6014 3853 6042 3909
rect 6098 3853 6126 3909
rect 6182 3853 6210 3909
rect 6266 3853 6623 3909
rect 5823 3828 6623 3853
rect 5823 3772 5874 3828
rect 5930 3772 5958 3828
rect 6014 3772 6042 3828
rect 6098 3772 6126 3828
rect 6182 3772 6210 3828
rect 6266 3772 6623 3828
rect 5823 3484 6623 3772
rect 5823 3428 5832 3484
rect 5888 3428 5953 3484
rect 6009 3428 6074 3484
rect 6130 3428 6195 3484
rect 6251 3428 6316 3484
rect 6372 3428 6437 3484
rect 6493 3428 6558 3484
rect 6614 3428 6623 3484
rect 5823 14 6623 3428
use nfet_CDNS_52468879185886  nfet_CDNS_52468879185886_0
timestamp 1707688321
transform 1 0 6822 0 -1 29806
box -82 -32 338 182
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_0
timestamp 1707688321
transform 0 -1 4538 1 0 5681
box -82 -32 1682 632
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_1
timestamp 1707688321
transform 0 -1 5268 1 0 5681
box -82 -32 1682 632
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_2
timestamp 1707688321
transform 0 -1 3808 1 0 5681
box -82 -32 1682 632
use nfet_CDNS_52468879185889  nfet_CDNS_52468879185889_0
timestamp 1707688321
transform 1 0 5838 0 1 29284
box -82 -32 1682 232
use nfet_CDNS_52468879185893  nfet_CDNS_52468879185893_0
timestamp 1707688321
transform 0 1 5484 1 0 30383
box -82 -32 9146 2032
use nfet_CDNS_52468879185906  nfet_CDNS_52468879185906_0
timestamp 1707688321
transform 1 0 7300 0 1 28512
box -82 -32 182 632
use nfet_CDNS_52468879185907  nfet_CDNS_52468879185907_0
timestamp 1707688321
transform 1 0 6934 0 1 28912
box -82 -32 182 232
use nfet_CDNS_52468879185907  nfet_CDNS_52468879185907_1
timestamp 1707688321
transform 1 0 6934 0 1 28540
box -82 -32 182 232
use nfet_CDNS_52468879185908  nfet_CDNS_52468879185908_0
timestamp 1707688321
transform -1 0 5804 0 -1 7190
box -82 -32 182 1432
use nfet_CDNS_52468879185909  nfet_CDNS_52468879185909_0
timestamp 1707688321
transform 0 -1 6382 1 0 5752
box -82 -32 882 232
use nfet_CDNS_52468879185909  nfet_CDNS_52468879185909_1
timestamp 1707688321
transform 1 0 5864 0 1 28912
box -82 -32 882 232
use nfet_CDNS_52468879185909  nfet_CDNS_52468879185909_2
timestamp 1707688321
transform 1 0 5864 0 1 28540
box -82 -32 882 232
use nfet_CDNS_52468879185910  nfet_CDNS_52468879185910_0
timestamp 1707688321
transform 0 -1 6382 1 0 6724
box -82 -32 482 232
use pfet_CDNS_52468879185895  pfet_CDNS_52468879185895_0
timestamp 1707688321
transform 1 0 6481 0 -1 21952
box -122 -66 378 366
use pfet_CDNS_52468879185902  pfet_CDNS_52468879185902_0
timestamp 1707688321
transform 1 0 3039 0 1 3291
box -119 -66 687 1466
use pfet_CDNS_52468879185903  pfet_CDNS_52468879185903_0
timestamp 1707688321
transform 0 -1 6618 1 0 3820
box -119 -66 975 266
use pfet_CDNS_52468879185904  pfet_CDNS_52468879185904_0
timestamp 1707688321
transform 1 0 4267 0 1 4491
box -119 -66 1719 266
use pfet_CDNS_52468879185904  pfet_CDNS_52468879185904_1
timestamp 1707688321
transform 1 0 4267 0 1 4161
box -119 -66 1719 266
use pfet_CDNS_52468879185905  pfet_CDNS_52468879185905_0
timestamp 1707688321
transform 1 0 4211 0 1 3767
box -119 -66 1775 266
use PYbentRes_CDNS_52468879185900  PYbentRes_CDNS_52468879185900_0
timestamp 1707688321
transform 0 -1 8198 -1 0 39549
box -50 -1458 38933 66
use PYres_CDNS_52468879185901  PYres_CDNS_52468879185901_0
timestamp 1707688321
transform 1 0 2875 0 1 27044
box -50 0 3177 66
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1707688321
transform 1 0 3440 0 -1 26854
box 0 0 2270 404
use sky130_fd_io__top_pwrdetv2_res1  sky130_fd_io__top_pwrdetv2_res1_0
timestamp 1707688321
transform 1 0 526 0 1 192
box 0 0 1912 39433
use sky130_fd_io__top_pwrdetv2_res6  sky130_fd_io__top_pwrdetv2_res6_0
timestamp 1707688321
transform 1 0 9836 0 1 1275
box 0 0 832 38350
use sky130_fd_io__top_pwrdetv2_res7  sky130_fd_io__top_pwrdetv2_res7_0
timestamp 1707688321
transform 1 0 7315 0 1 23547
box 0 0 472 3549
use sky130_fd_io__top_pwrdetv2_res7  sky130_fd_io__top_pwrdetv2_res7_1
timestamp 1707688321
transform 1 0 6489 0 1 23547
box 0 0 472 3549
<< labels >>
flabel comment s 6619 7255 6619 7255 0 FreeSans 600 90 0 0 condiode
flabel metal1 s 7795 4328 7870 4461 3 FreeSans 520 0 0 0 out
port 1 nsew
flabel metal1 s 3452 26520 3489 26781 3 FreeSans 520 0 0 0 vddd
port 2 nsew
flabel metal3 s 4663 39534 5663 39838 3 FreeSans 520 0 0 0 vssa
port 4 nsew
flabel metal3 s 5823 39464 6623 39822 3 FreeSans 520 0 0 0 vddio_q
port 5 nsew
<< properties >>
string GDS_END 7534530
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6699176
string path 186.350 238.750 186.350 284.550 161.550 284.550 
<< end >>
