magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 80 80 1870 1870
<< nwell >>
rect 70 1880 286 1950
rect 1664 1880 1880 1950
rect 0 1664 1950 1880
rect 70 286 286 1664
rect 1664 286 1880 1664
rect 0 70 1950 286
rect 70 0 286 70
rect 1664 0 1880 70
<< pbase >>
rect 286 286 1664 1664
<< mvnmos >>
tri 862 1125 888 1151 se
rect 888 1125 1063 1151
tri 1063 1125 1089 1151 sw
tri 850 1113 862 1125 se
rect 862 1113 888 1125
tri 888 1113 900 1125 nw
tri 1051 1113 1063 1125 ne
rect 1063 1113 1089 1125
tri 1089 1113 1101 1125 sw
tri 831 1094 850 1113 se
rect 850 1094 869 1113
tri 869 1094 888 1113 nw
tri 1063 1094 1082 1113 ne
rect 1082 1094 1101 1113
tri 1101 1094 1120 1113 sw
tri 799 1062 831 1094 se
rect 831 1062 837 1094
tri 837 1062 869 1094 nw
tri 1082 1063 1113 1094 ne
rect 1113 1063 1120 1094
tri 1120 1063 1151 1094 sw
rect 799 899 825 1062
tri 825 1050 837 1062 nw
tri 825 899 826 900 sw
rect 799 888 826 899
tri 826 888 837 899 sw
tri 1113 1051 1125 1063 ne
tri 799 856 831 888 ne
rect 831 856 837 888
tri 837 856 869 888 sw
tri 1113 887 1125 899 se
rect 1125 887 1151 1063
tri 1082 856 1113 887 se
rect 1113 856 1120 887
tri 1120 856 1151 887 nw
tri 831 837 850 856 ne
rect 850 837 869 856
tri 869 837 888 856 sw
tri 1063 837 1082 856 se
rect 1082 837 1101 856
tri 1101 837 1120 856 nw
tri 850 825 862 837 ne
rect 862 825 888 837
tri 888 825 900 837 sw
tri 1051 825 1063 837 se
rect 1063 825 1089 837
tri 1089 825 1101 837 nw
tri 862 799 888 825 ne
rect 888 799 1063 825
tri 1063 799 1089 825 nw
<< mvpmos >>
rect 512 1151 1438 1437
rect 512 1125 862 1151
tri 862 1125 888 1151 nw
tri 1063 1125 1089 1151 ne
rect 1089 1125 1438 1151
rect 512 1113 850 1125
tri 850 1113 862 1125 nw
tri 1089 1113 1101 1125 ne
rect 1101 1113 1438 1125
rect 512 1094 831 1113
tri 831 1094 850 1113 nw
tri 1101 1094 1120 1113 ne
rect 1120 1094 1438 1113
rect 512 856 799 1094
tri 799 1062 831 1094 nw
tri 1120 1063 1151 1094 ne
tri 799 856 831 888 sw
tri 1120 856 1151 887 se
rect 1151 856 1438 1094
rect 512 837 831 856
tri 831 837 850 856 sw
tri 1101 837 1120 856 se
rect 1120 837 1438 856
rect 512 825 850 837
tri 850 825 862 837 sw
tri 1089 825 1101 837 se
rect 1101 825 1438 837
rect 512 799 862 825
tri 862 799 888 825 sw
tri 1063 799 1089 825 se
rect 1089 799 1438 825
rect 512 512 1438 799
<< mvndiff >>
tri 888 1113 900 1125 se
rect 900 1113 1051 1125
tri 1051 1113 1063 1125 sw
tri 869 1094 888 1113 se
rect 888 1094 1063 1113
tri 1063 1094 1082 1113 sw
tri 837 1062 869 1094 se
rect 869 1063 1082 1094
tri 1082 1063 1113 1094 sw
rect 869 1062 1113 1063
tri 825 1050 837 1062 se
rect 837 1060 1113 1062
rect 837 1050 890 1060
rect 825 900 890 1050
tri 825 899 826 900 ne
rect 826 899 890 900
tri 826 888 837 899 ne
rect 837 890 890 899
rect 1060 1051 1113 1060
tri 1113 1051 1125 1063 sw
rect 1060 899 1125 1051
rect 1060 890 1113 899
rect 837 888 1113 890
tri 837 856 869 888 ne
rect 869 887 1113 888
tri 1113 887 1125 899 nw
rect 869 856 1082 887
tri 1082 856 1113 887 nw
tri 869 837 888 856 ne
rect 888 837 1063 856
tri 1063 837 1082 856 nw
tri 888 825 900 837 ne
rect 900 825 1051 837
tri 1051 825 1063 837 nw
<< mvndiffc >>
rect 890 890 1060 1060
<< mvpsubdiff >>
rect 372 1570 1578 1577
rect 372 1536 448 1570
rect 482 1536 516 1570
rect 550 1536 584 1570
rect 618 1536 652 1570
rect 686 1536 720 1570
rect 754 1536 788 1570
rect 822 1536 856 1570
rect 890 1536 924 1570
rect 958 1536 992 1570
rect 1026 1536 1060 1570
rect 1094 1536 1128 1570
rect 1162 1536 1196 1570
rect 1230 1536 1264 1570
rect 1298 1536 1332 1570
rect 1366 1536 1400 1570
rect 1434 1536 1468 1570
rect 1502 1536 1578 1570
rect 372 1502 1578 1536
rect 372 1468 380 1502
rect 414 1468 1536 1502
rect 1570 1468 1578 1502
rect 372 1437 1578 1468
rect 372 1434 512 1437
rect 372 1400 380 1434
rect 414 1400 512 1434
rect 372 1366 512 1400
rect 372 1332 380 1366
rect 414 1332 512 1366
rect 372 1298 512 1332
rect 372 1264 380 1298
rect 414 1264 512 1298
rect 372 1230 512 1264
rect 372 1196 380 1230
rect 414 1196 512 1230
rect 372 779 512 1196
rect 1438 1434 1578 1437
rect 1438 1400 1536 1434
rect 1570 1400 1578 1434
rect 1438 1366 1578 1400
rect 1438 1332 1536 1366
rect 1570 1332 1578 1366
rect 1438 1298 1578 1332
rect 1438 1264 1536 1298
rect 1570 1264 1578 1298
rect 1438 1230 1578 1264
rect 1438 1196 1536 1230
rect 1570 1196 1578 1230
rect 1438 1162 1578 1196
rect 1438 1128 1536 1162
rect 1570 1128 1578 1162
rect 1438 1094 1578 1128
rect 1438 1060 1536 1094
rect 1570 1060 1578 1094
rect 1438 1026 1578 1060
rect 1438 992 1536 1026
rect 1570 992 1578 1026
rect 1438 958 1578 992
rect 1438 924 1536 958
rect 1570 924 1578 958
rect 1438 890 1578 924
rect 1438 856 1536 890
rect 1570 856 1578 890
rect 1438 822 1578 856
rect 372 745 380 779
rect 414 745 512 779
rect 372 711 512 745
rect 372 677 380 711
rect 414 677 512 711
rect 372 643 512 677
rect 372 609 380 643
rect 414 609 512 643
rect 372 575 512 609
rect 372 541 380 575
rect 414 541 512 575
rect 372 512 512 541
rect 1438 788 1536 822
rect 1570 788 1578 822
rect 1438 754 1578 788
rect 1438 720 1536 754
rect 1570 720 1578 754
rect 1438 686 1578 720
rect 1438 652 1536 686
rect 1570 652 1578 686
rect 1438 618 1578 652
rect 1438 584 1536 618
rect 1570 584 1578 618
rect 1438 550 1578 584
rect 1438 516 1536 550
rect 1570 516 1578 550
rect 1438 512 1578 516
rect 372 507 1578 512
rect 372 473 380 507
rect 414 482 1578 507
rect 414 473 1536 482
rect 372 448 1536 473
rect 1570 448 1578 482
rect 372 414 1578 448
rect 372 380 448 414
rect 482 380 516 414
rect 550 380 584 414
rect 618 380 652 414
rect 686 380 720 414
rect 754 380 788 414
rect 822 380 856 414
rect 890 380 924 414
rect 958 380 992 414
rect 1026 380 1060 414
rect 1094 380 1128 414
rect 1162 380 1196 414
rect 1230 380 1264 414
rect 1298 380 1332 414
rect 1366 380 1400 414
rect 1434 380 1468 414
rect 1502 380 1578 414
rect 372 372 1578 380
<< mvnsubdiff >>
rect 137 1789 1813 1813
rect 137 1755 243 1789
rect 277 1755 311 1789
rect 345 1755 379 1789
rect 413 1755 447 1789
rect 481 1755 515 1789
rect 549 1755 583 1789
rect 617 1755 651 1789
rect 685 1755 719 1789
rect 753 1755 787 1789
rect 821 1755 855 1789
rect 889 1755 923 1789
rect 957 1755 991 1789
rect 1025 1755 1059 1789
rect 1093 1755 1127 1789
rect 1161 1755 1195 1789
rect 1229 1755 1263 1789
rect 1297 1755 1331 1789
rect 1365 1755 1399 1789
rect 1433 1755 1467 1789
rect 1501 1755 1535 1789
rect 1569 1755 1604 1789
rect 1638 1755 1673 1789
rect 1707 1755 1813 1789
rect 137 1731 1813 1755
rect 137 1707 219 1731
rect 137 1673 161 1707
rect 195 1673 219 1707
rect 137 1638 219 1673
rect 137 1604 161 1638
rect 195 1604 219 1638
rect 137 1569 219 1604
rect 1731 1707 1813 1731
rect 1731 1673 1755 1707
rect 1789 1673 1813 1707
rect 1731 1638 1813 1673
rect 1731 1604 1755 1638
rect 1789 1604 1813 1638
rect 137 1535 161 1569
rect 195 1535 219 1569
rect 137 1501 219 1535
rect 137 1467 161 1501
rect 195 1467 219 1501
rect 137 1433 219 1467
rect 137 1399 161 1433
rect 195 1399 219 1433
rect 137 1365 219 1399
rect 137 1331 161 1365
rect 195 1331 219 1365
rect 137 1297 219 1331
rect 137 1263 161 1297
rect 195 1263 219 1297
rect 137 1229 219 1263
rect 137 1195 161 1229
rect 195 1195 219 1229
rect 137 1161 219 1195
rect 137 1127 161 1161
rect 195 1127 219 1161
rect 137 1093 219 1127
rect 137 1059 161 1093
rect 195 1059 219 1093
rect 137 1025 219 1059
rect 137 991 161 1025
rect 195 991 219 1025
rect 137 957 219 991
rect 137 923 161 957
rect 195 923 219 957
rect 137 889 219 923
rect 137 855 161 889
rect 195 855 219 889
rect 137 821 219 855
rect 137 787 161 821
rect 195 787 219 821
rect 137 753 219 787
rect 137 719 161 753
rect 195 719 219 753
rect 137 685 219 719
rect 137 651 161 685
rect 195 651 219 685
rect 137 617 219 651
rect 137 583 161 617
rect 195 583 219 617
rect 137 549 219 583
rect 137 515 161 549
rect 195 515 219 549
rect 137 481 219 515
rect 137 447 161 481
rect 195 447 219 481
rect 137 413 219 447
rect 137 379 161 413
rect 195 379 219 413
rect 137 345 219 379
rect 1731 1569 1813 1604
rect 1731 1535 1755 1569
rect 1789 1535 1813 1569
rect 1731 1501 1813 1535
rect 1731 1467 1755 1501
rect 1789 1467 1813 1501
rect 1731 1433 1813 1467
rect 1731 1399 1755 1433
rect 1789 1399 1813 1433
rect 1731 1365 1813 1399
rect 1731 1331 1755 1365
rect 1789 1331 1813 1365
rect 1731 1297 1813 1331
rect 1731 1263 1755 1297
rect 1789 1263 1813 1297
rect 1731 1229 1813 1263
rect 1731 1195 1755 1229
rect 1789 1195 1813 1229
rect 1731 1161 1813 1195
rect 1731 1127 1755 1161
rect 1789 1127 1813 1161
rect 1731 1093 1813 1127
rect 1731 1059 1755 1093
rect 1789 1059 1813 1093
rect 1731 1025 1813 1059
rect 1731 991 1755 1025
rect 1789 991 1813 1025
rect 1731 957 1813 991
rect 1731 923 1755 957
rect 1789 923 1813 957
rect 1731 889 1813 923
rect 1731 855 1755 889
rect 1789 855 1813 889
rect 1731 821 1813 855
rect 1731 787 1755 821
rect 1789 787 1813 821
rect 1731 753 1813 787
rect 1731 719 1755 753
rect 1789 719 1813 753
rect 1731 685 1813 719
rect 1731 651 1755 685
rect 1789 651 1813 685
rect 1731 617 1813 651
rect 1731 583 1755 617
rect 1789 583 1813 617
rect 1731 549 1813 583
rect 1731 515 1755 549
rect 1789 515 1813 549
rect 1731 481 1813 515
rect 1731 447 1755 481
rect 1789 447 1813 481
rect 1731 413 1813 447
rect 1731 379 1755 413
rect 1789 379 1813 413
rect 137 311 161 345
rect 195 311 219 345
rect 137 277 219 311
rect 137 243 161 277
rect 195 243 219 277
rect 137 219 219 243
rect 1731 345 1813 379
rect 1731 311 1755 345
rect 1789 311 1813 345
rect 1731 277 1813 311
rect 1731 243 1755 277
rect 1789 243 1813 277
rect 1731 219 1813 243
rect 137 195 1813 219
rect 137 161 243 195
rect 277 161 311 195
rect 345 161 379 195
rect 413 161 447 195
rect 481 161 515 195
rect 549 161 583 195
rect 617 161 651 195
rect 685 161 719 195
rect 753 161 787 195
rect 821 161 855 195
rect 889 161 923 195
rect 957 161 991 195
rect 1025 161 1059 195
rect 1093 161 1127 195
rect 1161 161 1195 195
rect 1229 161 1263 195
rect 1297 161 1331 195
rect 1365 161 1399 195
rect 1433 161 1467 195
rect 1501 161 1535 195
rect 1569 161 1604 195
rect 1638 161 1673 195
rect 1707 161 1813 195
rect 137 137 1813 161
<< mvpsubdiffcont >>
rect 448 1536 482 1570
rect 516 1536 550 1570
rect 584 1536 618 1570
rect 652 1536 686 1570
rect 720 1536 754 1570
rect 788 1536 822 1570
rect 856 1536 890 1570
rect 924 1536 958 1570
rect 992 1536 1026 1570
rect 1060 1536 1094 1570
rect 1128 1536 1162 1570
rect 1196 1536 1230 1570
rect 1264 1536 1298 1570
rect 1332 1536 1366 1570
rect 1400 1536 1434 1570
rect 1468 1536 1502 1570
rect 380 1468 414 1502
rect 1536 1468 1570 1502
rect 380 1400 414 1434
rect 380 1332 414 1366
rect 380 1264 414 1298
rect 380 1196 414 1230
rect 1536 1400 1570 1434
rect 1536 1332 1570 1366
rect 1536 1264 1570 1298
rect 1536 1196 1570 1230
rect 1536 1128 1570 1162
rect 1536 1060 1570 1094
rect 1536 992 1570 1026
rect 1536 924 1570 958
rect 1536 856 1570 890
rect 380 745 414 779
rect 380 677 414 711
rect 380 609 414 643
rect 380 541 414 575
rect 1536 788 1570 822
rect 1536 720 1570 754
rect 1536 652 1570 686
rect 1536 584 1570 618
rect 1536 516 1570 550
rect 380 473 414 507
rect 1536 448 1570 482
rect 448 380 482 414
rect 516 380 550 414
rect 584 380 618 414
rect 652 380 686 414
rect 720 380 754 414
rect 788 380 822 414
rect 856 380 890 414
rect 924 380 958 414
rect 992 380 1026 414
rect 1060 380 1094 414
rect 1128 380 1162 414
rect 1196 380 1230 414
rect 1264 380 1298 414
rect 1332 380 1366 414
rect 1400 380 1434 414
rect 1468 380 1502 414
<< mvnsubdiffcont >>
rect 243 1755 277 1789
rect 311 1755 345 1789
rect 379 1755 413 1789
rect 447 1755 481 1789
rect 515 1755 549 1789
rect 583 1755 617 1789
rect 651 1755 685 1789
rect 719 1755 753 1789
rect 787 1755 821 1789
rect 855 1755 889 1789
rect 923 1755 957 1789
rect 991 1755 1025 1789
rect 1059 1755 1093 1789
rect 1127 1755 1161 1789
rect 1195 1755 1229 1789
rect 1263 1755 1297 1789
rect 1331 1755 1365 1789
rect 1399 1755 1433 1789
rect 1467 1755 1501 1789
rect 1535 1755 1569 1789
rect 1604 1755 1638 1789
rect 1673 1755 1707 1789
rect 161 1673 195 1707
rect 161 1604 195 1638
rect 1755 1673 1789 1707
rect 1755 1604 1789 1638
rect 161 1535 195 1569
rect 161 1467 195 1501
rect 161 1399 195 1433
rect 161 1331 195 1365
rect 161 1263 195 1297
rect 161 1195 195 1229
rect 161 1127 195 1161
rect 161 1059 195 1093
rect 161 991 195 1025
rect 161 923 195 957
rect 161 855 195 889
rect 161 787 195 821
rect 161 719 195 753
rect 161 651 195 685
rect 161 583 195 617
rect 161 515 195 549
rect 161 447 195 481
rect 161 379 195 413
rect 1755 1535 1789 1569
rect 1755 1467 1789 1501
rect 1755 1399 1789 1433
rect 1755 1331 1789 1365
rect 1755 1263 1789 1297
rect 1755 1195 1789 1229
rect 1755 1127 1789 1161
rect 1755 1059 1789 1093
rect 1755 991 1789 1025
rect 1755 923 1789 957
rect 1755 855 1789 889
rect 1755 787 1789 821
rect 1755 719 1789 753
rect 1755 651 1789 685
rect 1755 583 1789 617
rect 1755 515 1789 549
rect 1755 447 1789 481
rect 1755 379 1789 413
rect 161 311 195 345
rect 161 243 195 277
rect 1755 311 1789 345
rect 1755 243 1789 277
rect 243 161 277 195
rect 311 161 345 195
rect 379 161 413 195
rect 447 161 481 195
rect 515 161 549 195
rect 583 161 617 195
rect 651 161 685 195
rect 719 161 753 195
rect 787 161 821 195
rect 855 161 889 195
rect 923 161 957 195
rect 991 161 1025 195
rect 1059 161 1093 195
rect 1127 161 1161 195
rect 1195 161 1229 195
rect 1263 161 1297 195
rect 1331 161 1365 195
rect 1399 161 1433 195
rect 1467 161 1501 195
rect 1535 161 1569 195
rect 1604 161 1638 195
rect 1673 161 1707 195
<< poly >>
rect 261 1025 372 1041
rect 261 991 277 1025
rect 311 991 372 1025
rect 261 957 372 991
rect 261 923 277 957
rect 311 923 372 957
rect 261 907 372 923
<< polycont >>
rect 277 991 311 1025
rect 277 923 311 957
<< locali >>
rect 137 1789 1813 1813
rect 137 1755 243 1789
rect 293 1755 311 1789
rect 366 1755 379 1789
rect 439 1755 447 1789
rect 512 1755 515 1789
rect 549 1755 551 1789
rect 617 1755 625 1789
rect 685 1755 699 1789
rect 753 1755 773 1789
rect 821 1755 847 1789
rect 889 1755 921 1789
rect 957 1755 991 1789
rect 1029 1755 1059 1789
rect 1103 1755 1127 1789
rect 1177 1755 1195 1789
rect 1251 1755 1263 1789
rect 1325 1755 1331 1789
rect 1433 1755 1439 1789
rect 1501 1755 1513 1789
rect 1569 1755 1587 1789
rect 1638 1755 1661 1789
rect 1707 1755 1813 1789
rect 137 1731 1813 1755
rect 137 1707 219 1731
rect 137 1662 161 1707
rect 195 1662 219 1707
rect 137 1638 219 1662
rect 137 1588 161 1638
rect 195 1588 219 1638
rect 1731 1707 1813 1731
rect 1731 1662 1755 1707
rect 1789 1662 1813 1707
rect 1731 1638 1813 1662
rect 137 1569 219 1588
rect 137 1514 161 1569
rect 195 1514 219 1569
rect 137 1501 219 1514
rect 137 1440 161 1501
rect 195 1440 219 1501
rect 137 1433 219 1440
rect 137 1366 161 1433
rect 195 1366 219 1433
rect 137 1365 219 1366
rect 137 1331 161 1365
rect 195 1331 219 1365
rect 137 1326 219 1331
rect 137 1263 161 1326
rect 195 1263 219 1326
rect 137 1252 219 1263
rect 137 1195 161 1252
rect 195 1195 219 1252
rect 137 1178 219 1195
rect 137 1127 161 1178
rect 195 1127 219 1178
rect 332 1593 1616 1616
rect 332 1559 414 1593
rect 448 1570 487 1593
rect 521 1570 560 1593
rect 594 1570 633 1593
rect 667 1570 706 1593
rect 740 1570 779 1593
rect 813 1570 852 1593
rect 886 1570 924 1593
rect 958 1570 996 1593
rect 1030 1570 1068 1593
rect 1102 1570 1140 1593
rect 1174 1570 1212 1593
rect 1246 1570 1284 1593
rect 1318 1570 1356 1593
rect 1390 1570 1428 1593
rect 1462 1570 1616 1593
rect 332 1536 448 1559
rect 482 1559 487 1570
rect 550 1559 560 1570
rect 618 1559 633 1570
rect 686 1559 706 1570
rect 754 1559 779 1570
rect 822 1559 852 1570
rect 482 1536 516 1559
rect 550 1536 584 1559
rect 618 1536 652 1559
rect 686 1536 720 1559
rect 754 1536 788 1559
rect 822 1536 856 1559
rect 890 1536 924 1570
rect 958 1536 992 1570
rect 1030 1559 1060 1570
rect 1102 1559 1128 1570
rect 1174 1559 1196 1570
rect 1246 1559 1264 1570
rect 1318 1559 1332 1570
rect 1390 1559 1400 1570
rect 1462 1559 1468 1570
rect 1026 1536 1060 1559
rect 1094 1536 1128 1559
rect 1162 1536 1196 1559
rect 1230 1536 1264 1559
rect 1298 1536 1332 1559
rect 1366 1536 1400 1559
rect 1434 1536 1468 1559
rect 1502 1536 1616 1570
rect 332 1522 414 1536
rect 332 1488 355 1522
rect 389 1502 414 1522
rect 332 1468 380 1488
rect 332 1437 414 1468
rect 332 1403 355 1437
rect 389 1434 414 1437
rect 332 1400 380 1403
rect 332 1366 414 1400
rect 332 1352 380 1366
rect 332 1318 355 1352
rect 389 1318 414 1332
rect 332 1298 414 1318
rect 332 1267 380 1298
rect 332 1233 355 1267
rect 389 1233 414 1264
rect 332 1230 414 1233
rect 332 1196 380 1230
rect 332 1182 414 1196
rect 332 1148 355 1182
rect 389 1148 414 1182
rect 332 1136 414 1148
rect 1536 1534 1616 1536
rect 1536 1502 1559 1534
rect 1593 1500 1616 1534
rect 1570 1468 1616 1500
rect 1536 1461 1616 1468
rect 1536 1434 1559 1461
rect 1593 1427 1616 1461
rect 1570 1400 1616 1427
rect 1536 1388 1616 1400
rect 1536 1366 1559 1388
rect 1593 1354 1616 1388
rect 1570 1332 1616 1354
rect 1536 1315 1616 1332
rect 1536 1298 1559 1315
rect 1593 1281 1616 1315
rect 1570 1264 1616 1281
rect 1536 1242 1616 1264
rect 1536 1230 1559 1242
rect 1593 1208 1616 1242
rect 1570 1196 1616 1208
rect 1536 1170 1616 1196
rect 1536 1162 1559 1170
rect 1593 1136 1616 1170
rect 137 1104 219 1127
rect 137 1059 161 1104
rect 195 1059 219 1104
rect 1570 1128 1616 1136
rect 1536 1098 1616 1128
rect 1536 1094 1559 1098
rect 137 1030 219 1059
rect 137 991 161 1030
rect 195 991 219 1030
rect 137 957 219 991
rect 137 922 161 957
rect 195 922 219 957
rect 137 889 219 922
rect 137 848 161 889
rect 195 848 219 889
rect 261 1042 295 1076
rect 329 1042 367 1076
rect 401 1042 439 1076
rect 473 1060 1076 1076
rect 473 1042 890 1060
rect 261 1025 890 1042
rect 261 991 277 1025
rect 311 992 890 1025
rect 261 958 295 991
rect 329 958 367 992
rect 401 958 439 992
rect 473 958 890 992
rect 261 957 890 958
rect 261 923 277 957
rect 311 923 890 957
rect 261 908 890 923
rect 261 874 295 908
rect 329 874 367 908
rect 401 874 439 908
rect 473 890 890 908
rect 1060 890 1076 1060
rect 473 874 1076 890
rect 1593 1064 1616 1098
rect 1570 1060 1616 1064
rect 1536 1026 1616 1060
rect 1593 992 1616 1026
rect 1536 958 1616 992
rect 1570 954 1616 958
rect 1536 920 1559 924
rect 1593 920 1616 954
rect 1536 890 1616 920
rect 1570 882 1616 890
rect 137 821 219 848
rect 137 774 161 821
rect 195 774 219 821
rect 1536 848 1559 856
rect 1593 848 1616 882
rect 1536 822 1616 848
rect 137 753 219 774
rect 137 700 161 753
rect 195 700 219 753
rect 137 685 219 700
rect 137 626 161 685
rect 195 626 219 685
rect 137 617 219 626
rect 137 552 161 617
rect 195 552 219 617
rect 137 549 219 552
rect 137 515 161 549
rect 195 515 219 549
rect 137 512 219 515
rect 137 447 161 512
rect 195 447 219 512
rect 137 439 219 447
rect 137 379 161 439
rect 195 379 219 439
rect 137 366 219 379
rect 137 311 161 366
rect 195 311 219 366
rect 332 801 414 813
rect 332 767 355 801
rect 389 779 414 801
rect 332 745 380 767
rect 332 714 414 745
rect 332 680 355 714
rect 389 711 414 714
rect 332 677 380 680
rect 332 643 414 677
rect 332 626 380 643
rect 332 592 355 626
rect 389 592 414 609
rect 332 575 414 592
rect 332 541 380 575
rect 332 538 414 541
rect 332 504 355 538
rect 389 507 414 538
rect 332 473 380 504
rect 332 450 414 473
rect 332 416 355 450
rect 389 416 414 450
rect 332 414 414 416
rect 1570 810 1616 822
rect 1536 776 1559 788
rect 1593 776 1616 810
rect 1536 754 1616 776
rect 1570 738 1616 754
rect 1536 704 1559 720
rect 1593 704 1616 738
rect 1536 686 1616 704
rect 1570 666 1616 686
rect 1536 632 1559 652
rect 1593 632 1616 666
rect 1536 618 1616 632
rect 1570 594 1616 618
rect 1536 560 1559 584
rect 1593 560 1616 594
rect 1536 550 1616 560
rect 1570 522 1616 550
rect 1536 488 1559 516
rect 1593 488 1616 522
rect 1536 482 1616 488
rect 1570 448 1616 482
rect 1536 414 1616 448
rect 332 380 448 414
rect 482 391 516 414
rect 550 391 584 414
rect 618 391 652 414
rect 686 391 720 414
rect 754 391 788 414
rect 822 391 856 414
rect 890 391 924 414
rect 958 391 992 414
rect 482 380 486 391
rect 550 380 558 391
rect 618 380 630 391
rect 686 380 702 391
rect 754 380 774 391
rect 822 380 846 391
rect 890 380 918 391
rect 958 380 990 391
rect 1026 380 1060 414
rect 1094 391 1128 414
rect 1162 391 1196 414
rect 1230 391 1264 414
rect 1298 391 1332 414
rect 1366 391 1400 414
rect 1434 391 1468 414
rect 1502 391 1616 414
rect 1096 380 1128 391
rect 1169 380 1196 391
rect 1242 380 1264 391
rect 1315 380 1332 391
rect 1388 380 1400 391
rect 1461 380 1468 391
rect 332 357 486 380
rect 520 357 558 380
rect 592 357 630 380
rect 664 357 702 380
rect 736 357 774 380
rect 808 357 846 380
rect 880 357 918 380
rect 952 357 990 380
rect 1024 357 1062 380
rect 1096 357 1135 380
rect 1169 357 1208 380
rect 1242 357 1281 380
rect 1315 357 1354 380
rect 1388 357 1427 380
rect 1461 357 1500 380
rect 1534 357 1616 391
rect 332 334 1616 357
rect 1731 1588 1755 1638
rect 1789 1588 1813 1638
rect 1731 1569 1813 1588
rect 1731 1514 1755 1569
rect 1789 1514 1813 1569
rect 1731 1501 1813 1514
rect 1731 1440 1755 1501
rect 1789 1440 1813 1501
rect 1731 1433 1813 1440
rect 1731 1366 1755 1433
rect 1789 1366 1813 1433
rect 1731 1365 1813 1366
rect 1731 1331 1755 1365
rect 1789 1331 1813 1365
rect 1731 1326 1813 1331
rect 1731 1263 1755 1326
rect 1789 1263 1813 1326
rect 1731 1252 1813 1263
rect 1731 1195 1755 1252
rect 1789 1195 1813 1252
rect 1731 1178 1813 1195
rect 1731 1127 1755 1178
rect 1789 1127 1813 1178
rect 1731 1104 1813 1127
rect 1731 1059 1755 1104
rect 1789 1059 1813 1104
rect 1731 1030 1813 1059
rect 1731 991 1755 1030
rect 1789 991 1813 1030
rect 1731 957 1813 991
rect 1731 922 1755 957
rect 1789 922 1813 957
rect 1731 889 1813 922
rect 1731 848 1755 889
rect 1789 848 1813 889
rect 1731 821 1813 848
rect 1731 774 1755 821
rect 1789 774 1813 821
rect 1731 753 1813 774
rect 1731 700 1755 753
rect 1789 700 1813 753
rect 1731 685 1813 700
rect 1731 626 1755 685
rect 1789 626 1813 685
rect 1731 617 1813 626
rect 1731 552 1755 617
rect 1789 552 1813 617
rect 1731 549 1813 552
rect 1731 515 1755 549
rect 1789 515 1813 549
rect 1731 512 1813 515
rect 1731 447 1755 512
rect 1789 447 1813 512
rect 1731 439 1813 447
rect 1731 379 1755 439
rect 1789 379 1813 439
rect 1731 366 1813 379
rect 137 293 219 311
rect 137 243 161 293
rect 195 243 219 293
rect 137 219 219 243
rect 1731 311 1755 366
rect 1789 311 1813 366
rect 1731 293 1813 311
rect 1731 243 1755 293
rect 1789 243 1813 293
rect 1731 219 1813 243
rect 137 195 1813 219
rect 137 161 243 195
rect 293 161 311 195
rect 366 161 379 195
rect 439 161 447 195
rect 512 161 515 195
rect 549 161 551 195
rect 617 161 625 195
rect 685 161 699 195
rect 753 161 773 195
rect 821 161 847 195
rect 889 161 921 195
rect 957 161 991 195
rect 1029 161 1059 195
rect 1103 161 1127 195
rect 1177 161 1195 195
rect 1251 161 1263 195
rect 1325 161 1331 195
rect 1433 161 1439 195
rect 1501 161 1513 195
rect 1569 161 1587 195
rect 1638 161 1661 195
rect 1707 161 1813 195
rect 137 137 1813 161
<< viali >>
rect 259 1755 277 1789
rect 277 1755 293 1789
rect 332 1755 345 1789
rect 345 1755 366 1789
rect 405 1755 413 1789
rect 413 1755 439 1789
rect 478 1755 481 1789
rect 481 1755 512 1789
rect 551 1755 583 1789
rect 583 1755 585 1789
rect 625 1755 651 1789
rect 651 1755 659 1789
rect 699 1755 719 1789
rect 719 1755 733 1789
rect 773 1755 787 1789
rect 787 1755 807 1789
rect 847 1755 855 1789
rect 855 1755 881 1789
rect 921 1755 923 1789
rect 923 1755 955 1789
rect 995 1755 1025 1789
rect 1025 1755 1029 1789
rect 1069 1755 1093 1789
rect 1093 1755 1103 1789
rect 1143 1755 1161 1789
rect 1161 1755 1177 1789
rect 1217 1755 1229 1789
rect 1229 1755 1251 1789
rect 1291 1755 1297 1789
rect 1297 1755 1325 1789
rect 1365 1755 1399 1789
rect 1439 1755 1467 1789
rect 1467 1755 1473 1789
rect 1513 1755 1535 1789
rect 1535 1755 1547 1789
rect 1587 1755 1604 1789
rect 1604 1755 1621 1789
rect 1661 1755 1673 1789
rect 1673 1755 1695 1789
rect 161 1673 195 1696
rect 161 1662 195 1673
rect 161 1604 195 1622
rect 161 1588 195 1604
rect 1755 1673 1789 1696
rect 1755 1662 1789 1673
rect 161 1535 195 1548
rect 161 1514 195 1535
rect 161 1467 195 1474
rect 161 1440 195 1467
rect 161 1399 195 1400
rect 161 1366 195 1399
rect 161 1297 195 1326
rect 161 1292 195 1297
rect 161 1229 195 1252
rect 161 1218 195 1229
rect 161 1161 195 1178
rect 161 1144 195 1161
rect 414 1559 448 1593
rect 487 1570 521 1593
rect 560 1570 594 1593
rect 633 1570 667 1593
rect 706 1570 740 1593
rect 779 1570 813 1593
rect 852 1570 886 1593
rect 924 1570 958 1593
rect 996 1570 1030 1593
rect 1068 1570 1102 1593
rect 1140 1570 1174 1593
rect 1212 1570 1246 1593
rect 1284 1570 1318 1593
rect 1356 1570 1390 1593
rect 1428 1570 1462 1593
rect 487 1559 516 1570
rect 516 1559 521 1570
rect 560 1559 584 1570
rect 584 1559 594 1570
rect 633 1559 652 1570
rect 652 1559 667 1570
rect 706 1559 720 1570
rect 720 1559 740 1570
rect 779 1559 788 1570
rect 788 1559 813 1570
rect 852 1559 856 1570
rect 856 1559 886 1570
rect 924 1559 958 1570
rect 996 1559 1026 1570
rect 1026 1559 1030 1570
rect 1068 1559 1094 1570
rect 1094 1559 1102 1570
rect 1140 1559 1162 1570
rect 1162 1559 1174 1570
rect 1212 1559 1230 1570
rect 1230 1559 1246 1570
rect 1284 1559 1298 1570
rect 1298 1559 1318 1570
rect 1356 1559 1366 1570
rect 1366 1559 1390 1570
rect 1428 1559 1434 1570
rect 1434 1559 1462 1570
rect 355 1502 389 1522
rect 355 1488 380 1502
rect 380 1488 389 1502
rect 355 1434 389 1437
rect 355 1403 380 1434
rect 380 1403 389 1434
rect 355 1332 380 1352
rect 380 1332 389 1352
rect 355 1318 389 1332
rect 355 1264 380 1267
rect 380 1264 389 1267
rect 355 1233 389 1264
rect 355 1148 389 1182
rect 1559 1502 1593 1534
rect 1559 1500 1570 1502
rect 1570 1500 1593 1502
rect 1559 1434 1593 1461
rect 1559 1427 1570 1434
rect 1570 1427 1593 1434
rect 1559 1366 1593 1388
rect 1559 1354 1570 1366
rect 1570 1354 1593 1366
rect 1559 1298 1593 1315
rect 1559 1281 1570 1298
rect 1570 1281 1593 1298
rect 1559 1230 1593 1242
rect 1559 1208 1570 1230
rect 1570 1208 1593 1230
rect 1559 1162 1593 1170
rect 1559 1136 1570 1162
rect 1570 1136 1593 1162
rect 161 1093 195 1104
rect 161 1070 195 1093
rect 1559 1094 1593 1098
rect 161 1025 195 1030
rect 161 996 195 1025
rect 161 923 195 956
rect 161 922 195 923
rect 161 855 195 882
rect 161 848 195 855
rect 295 1042 329 1076
rect 367 1042 401 1076
rect 439 1042 473 1076
rect 295 991 311 992
rect 311 991 329 992
rect 295 958 329 991
rect 367 958 401 992
rect 439 958 473 992
rect 295 874 329 908
rect 367 874 401 908
rect 439 874 473 908
rect 1559 1064 1570 1094
rect 1570 1064 1593 1094
rect 1559 992 1570 1026
rect 1570 992 1593 1026
rect 1559 924 1570 954
rect 1570 924 1593 954
rect 1559 920 1593 924
rect 161 787 195 808
rect 161 774 195 787
rect 1559 856 1570 882
rect 1570 856 1593 882
rect 1559 848 1593 856
rect 161 719 195 734
rect 161 700 195 719
rect 161 651 195 660
rect 161 626 195 651
rect 161 583 195 586
rect 161 552 195 583
rect 161 481 195 512
rect 161 478 195 481
rect 161 413 195 439
rect 161 405 195 413
rect 161 345 195 366
rect 161 332 195 345
rect 355 779 389 801
rect 355 767 380 779
rect 380 767 389 779
rect 355 711 389 714
rect 355 680 380 711
rect 380 680 389 711
rect 355 609 380 626
rect 380 609 389 626
rect 355 592 389 609
rect 355 507 389 538
rect 355 504 380 507
rect 380 504 389 507
rect 355 416 389 450
rect 1559 788 1570 810
rect 1570 788 1593 810
rect 1559 776 1593 788
rect 1559 720 1570 738
rect 1570 720 1593 738
rect 1559 704 1593 720
rect 1559 652 1570 666
rect 1570 652 1593 666
rect 1559 632 1593 652
rect 1559 584 1570 594
rect 1570 584 1593 594
rect 1559 560 1593 584
rect 1559 516 1570 522
rect 1570 516 1593 522
rect 1559 488 1593 516
rect 486 380 516 391
rect 516 380 520 391
rect 558 380 584 391
rect 584 380 592 391
rect 630 380 652 391
rect 652 380 664 391
rect 702 380 720 391
rect 720 380 736 391
rect 774 380 788 391
rect 788 380 808 391
rect 846 380 856 391
rect 856 380 880 391
rect 918 380 924 391
rect 924 380 952 391
rect 990 380 992 391
rect 992 380 1024 391
rect 1062 380 1094 391
rect 1094 380 1096 391
rect 1135 380 1162 391
rect 1162 380 1169 391
rect 1208 380 1230 391
rect 1230 380 1242 391
rect 1281 380 1298 391
rect 1298 380 1315 391
rect 1354 380 1366 391
rect 1366 380 1388 391
rect 1427 380 1434 391
rect 1434 380 1461 391
rect 1500 380 1502 391
rect 1502 380 1534 391
rect 486 357 520 380
rect 558 357 592 380
rect 630 357 664 380
rect 702 357 736 380
rect 774 357 808 380
rect 846 357 880 380
rect 918 357 952 380
rect 990 357 1024 380
rect 1062 357 1096 380
rect 1135 357 1169 380
rect 1208 357 1242 380
rect 1281 357 1315 380
rect 1354 357 1388 380
rect 1427 357 1461 380
rect 1500 357 1534 380
rect 1755 1604 1789 1622
rect 1755 1588 1789 1604
rect 1755 1535 1789 1548
rect 1755 1514 1789 1535
rect 1755 1467 1789 1474
rect 1755 1440 1789 1467
rect 1755 1399 1789 1400
rect 1755 1366 1789 1399
rect 1755 1297 1789 1326
rect 1755 1292 1789 1297
rect 1755 1229 1789 1252
rect 1755 1218 1789 1229
rect 1755 1161 1789 1178
rect 1755 1144 1789 1161
rect 1755 1093 1789 1104
rect 1755 1070 1789 1093
rect 1755 1025 1789 1030
rect 1755 996 1789 1025
rect 1755 923 1789 956
rect 1755 922 1789 923
rect 1755 855 1789 882
rect 1755 848 1789 855
rect 1755 787 1789 808
rect 1755 774 1789 787
rect 1755 719 1789 734
rect 1755 700 1789 719
rect 1755 651 1789 660
rect 1755 626 1789 651
rect 1755 583 1789 586
rect 1755 552 1789 583
rect 1755 481 1789 512
rect 1755 478 1789 481
rect 1755 413 1789 439
rect 1755 405 1789 413
rect 161 277 195 293
rect 161 259 195 277
rect 1755 345 1789 366
rect 1755 332 1789 345
rect 1755 277 1789 293
rect 1755 259 1789 277
rect 259 161 277 195
rect 277 161 293 195
rect 332 161 345 195
rect 345 161 366 195
rect 405 161 413 195
rect 413 161 439 195
rect 478 161 481 195
rect 481 161 512 195
rect 551 161 583 195
rect 583 161 585 195
rect 625 161 651 195
rect 651 161 659 195
rect 699 161 719 195
rect 719 161 733 195
rect 773 161 787 195
rect 787 161 807 195
rect 847 161 855 195
rect 855 161 881 195
rect 921 161 923 195
rect 923 161 955 195
rect 995 161 1025 195
rect 1025 161 1029 195
rect 1069 161 1093 195
rect 1093 161 1103 195
rect 1143 161 1161 195
rect 1161 161 1177 195
rect 1217 161 1229 195
rect 1229 161 1251 195
rect 1291 161 1297 195
rect 1297 161 1325 195
rect 1365 161 1399 195
rect 1439 161 1467 195
rect 1467 161 1473 195
rect 1513 161 1535 195
rect 1535 161 1547 195
rect 1587 161 1604 195
rect 1604 161 1621 195
rect 1661 161 1673 195
rect 1673 161 1695 195
<< metal1 >>
rect 142 1789 1808 1809
rect 142 1755 259 1789
rect 293 1755 332 1789
rect 366 1755 405 1789
rect 439 1755 478 1789
rect 512 1755 551 1789
rect 585 1755 625 1789
rect 659 1755 699 1789
rect 733 1755 773 1789
rect 807 1755 847 1789
rect 881 1755 921 1789
rect 955 1755 995 1789
rect 1029 1755 1069 1789
rect 1103 1755 1143 1789
rect 1177 1755 1217 1789
rect 1251 1755 1291 1789
rect 1325 1755 1365 1789
rect 1399 1755 1439 1789
rect 1473 1755 1513 1789
rect 1547 1755 1587 1789
rect 1621 1755 1661 1789
rect 1695 1755 1808 1789
rect 142 1737 1808 1755
rect 142 1696 214 1737
rect 142 1662 161 1696
rect 195 1662 214 1696
rect 142 1622 214 1662
rect 142 1588 161 1622
rect 195 1588 214 1622
rect 1736 1696 1808 1737
rect 1736 1662 1755 1696
rect 1789 1662 1808 1696
rect 1736 1622 1808 1662
rect 142 1548 214 1588
rect 142 1514 161 1548
rect 195 1514 214 1548
rect 142 1474 214 1514
rect 142 1440 161 1474
rect 195 1440 214 1474
rect 142 1400 214 1440
rect 142 1366 161 1400
rect 195 1366 214 1400
rect 142 1326 214 1366
rect 142 1292 161 1326
rect 195 1292 214 1326
rect 142 1252 214 1292
rect 142 1218 161 1252
rect 195 1218 214 1252
rect 142 1178 214 1218
rect 142 1144 161 1178
rect 195 1144 214 1178
rect 142 1104 214 1144
rect 336 1593 1612 1612
rect 336 1559 414 1593
rect 448 1559 487 1593
rect 521 1559 560 1593
rect 594 1559 633 1593
rect 667 1559 706 1593
rect 740 1559 779 1593
rect 813 1559 852 1593
rect 886 1559 924 1593
rect 958 1559 996 1593
rect 1030 1559 1068 1593
rect 1102 1559 1140 1593
rect 1174 1559 1212 1593
rect 1246 1559 1284 1593
rect 1318 1559 1356 1593
rect 1390 1559 1428 1593
rect 1462 1559 1612 1593
rect 336 1540 1612 1559
rect 336 1522 408 1540
rect 336 1488 355 1522
rect 389 1488 408 1522
rect 336 1437 408 1488
rect 336 1403 355 1437
rect 389 1403 408 1437
rect 336 1352 408 1403
rect 336 1318 355 1352
rect 389 1318 408 1352
rect 336 1267 408 1318
rect 336 1233 355 1267
rect 389 1233 408 1267
rect 336 1182 408 1233
rect 336 1148 355 1182
rect 389 1148 408 1182
rect 336 1136 408 1148
rect 1540 1534 1612 1540
rect 1540 1500 1559 1534
rect 1593 1500 1612 1534
rect 1540 1461 1612 1500
rect 1540 1427 1559 1461
rect 1593 1427 1612 1461
rect 1540 1388 1612 1427
rect 1540 1354 1559 1388
rect 1593 1354 1612 1388
rect 1540 1315 1612 1354
rect 1540 1281 1559 1315
rect 1593 1281 1612 1315
rect 1540 1242 1612 1281
rect 1540 1208 1559 1242
rect 1593 1208 1612 1242
rect 1540 1170 1612 1208
rect 1540 1136 1559 1170
rect 1593 1136 1612 1170
rect 142 1070 161 1104
rect 195 1070 214 1104
rect 1540 1098 1612 1136
rect 142 1030 214 1070
rect 142 996 161 1030
rect 195 996 214 1030
rect 142 956 214 996
rect 142 922 161 956
rect 195 922 214 956
rect 142 882 214 922
rect 142 848 161 882
rect 195 848 214 882
rect 289 1076 479 1088
rect 289 1042 295 1076
rect 329 1042 367 1076
rect 401 1042 439 1076
rect 473 1042 479 1076
rect 289 992 479 1042
rect 289 958 295 992
rect 329 958 367 992
rect 401 958 439 992
rect 473 958 479 992
rect 289 908 479 958
rect 289 874 295 908
rect 329 874 367 908
rect 401 874 439 908
rect 473 874 479 908
rect 289 862 479 874
rect 1540 1064 1559 1098
rect 1593 1064 1612 1098
rect 1540 1026 1612 1064
rect 1540 992 1559 1026
rect 1593 992 1612 1026
rect 1540 954 1612 992
rect 1540 920 1559 954
rect 1593 920 1612 954
rect 1540 882 1612 920
rect 142 808 214 848
rect 1540 848 1559 882
rect 1593 848 1612 882
rect 142 774 161 808
rect 195 774 214 808
rect 142 734 214 774
rect 142 700 161 734
rect 195 700 214 734
rect 142 660 214 700
rect 142 626 161 660
rect 195 626 214 660
rect 142 586 214 626
rect 142 552 161 586
rect 195 552 214 586
rect 142 512 214 552
rect 142 478 161 512
rect 195 478 214 512
rect 142 439 214 478
rect 142 405 161 439
rect 195 405 214 439
rect 142 366 214 405
rect 142 332 161 366
rect 195 332 214 366
rect 336 801 408 813
rect 336 767 355 801
rect 389 767 408 801
rect 336 714 408 767
rect 336 680 355 714
rect 389 680 408 714
rect 336 626 408 680
rect 336 592 355 626
rect 389 592 408 626
rect 336 538 408 592
rect 336 504 355 538
rect 389 504 408 538
rect 336 450 408 504
rect 336 416 355 450
rect 389 416 408 450
rect 336 410 408 416
rect 1540 810 1612 848
rect 1540 776 1559 810
rect 1593 776 1612 810
rect 1540 738 1612 776
rect 1540 704 1559 738
rect 1593 704 1612 738
rect 1540 666 1612 704
rect 1540 632 1559 666
rect 1593 632 1612 666
rect 1540 594 1612 632
rect 1540 560 1559 594
rect 1593 560 1612 594
rect 1540 522 1612 560
rect 1540 488 1559 522
rect 1593 488 1612 522
rect 1540 410 1612 488
rect 336 391 1612 410
rect 336 357 486 391
rect 520 357 558 391
rect 592 357 630 391
rect 664 357 702 391
rect 736 357 774 391
rect 808 357 846 391
rect 880 357 918 391
rect 952 357 990 391
rect 1024 357 1062 391
rect 1096 357 1135 391
rect 1169 357 1208 391
rect 1242 357 1281 391
rect 1315 357 1354 391
rect 1388 357 1427 391
rect 1461 357 1500 391
rect 1534 357 1612 391
rect 336 338 1612 357
rect 1736 1588 1755 1622
rect 1789 1588 1808 1622
rect 1736 1548 1808 1588
rect 1736 1514 1755 1548
rect 1789 1514 1808 1548
rect 1736 1474 1808 1514
rect 1736 1440 1755 1474
rect 1789 1440 1808 1474
rect 1736 1400 1808 1440
rect 1736 1366 1755 1400
rect 1789 1366 1808 1400
rect 1736 1326 1808 1366
rect 1736 1292 1755 1326
rect 1789 1292 1808 1326
rect 1736 1252 1808 1292
rect 1736 1218 1755 1252
rect 1789 1218 1808 1252
rect 1736 1178 1808 1218
rect 1736 1144 1755 1178
rect 1789 1144 1808 1178
rect 1736 1104 1808 1144
rect 1736 1070 1755 1104
rect 1789 1070 1808 1104
rect 1736 1030 1808 1070
rect 1736 996 1755 1030
rect 1789 996 1808 1030
rect 1736 956 1808 996
rect 1736 922 1755 956
rect 1789 922 1808 956
rect 1736 882 1808 922
rect 1736 848 1755 882
rect 1789 848 1808 882
rect 1736 808 1808 848
rect 1736 774 1755 808
rect 1789 774 1808 808
rect 1736 734 1808 774
rect 1736 700 1755 734
rect 1789 700 1808 734
rect 1736 660 1808 700
rect 1736 626 1755 660
rect 1789 626 1808 660
rect 1736 586 1808 626
rect 1736 552 1755 586
rect 1789 552 1808 586
rect 1736 512 1808 552
rect 1736 478 1755 512
rect 1789 478 1808 512
rect 1736 439 1808 478
rect 1736 405 1755 439
rect 1789 405 1808 439
rect 1736 366 1808 405
rect 142 293 214 332
rect 142 259 161 293
rect 195 259 214 293
rect 142 214 214 259
rect 1736 332 1755 366
rect 1789 332 1808 366
rect 1736 293 1808 332
rect 1736 259 1755 293
rect 1789 259 1808 293
rect 1736 214 1808 259
rect 142 195 1808 214
rect 142 161 259 195
rect 293 161 332 195
rect 366 161 405 195
rect 439 161 478 195
rect 512 161 551 195
rect 585 161 625 195
rect 659 161 699 195
rect 733 161 773 195
rect 807 161 847 195
rect 881 161 921 195
rect 955 161 995 195
rect 1029 161 1069 195
rect 1103 161 1143 195
rect 1177 161 1217 195
rect 1251 161 1291 195
rect 1325 161 1365 195
rect 1399 161 1439 195
rect 1473 161 1513 195
rect 1547 161 1587 195
rect 1621 161 1661 195
rect 1695 161 1808 195
rect 142 142 1808 161
<< labels >>
flabel metal1 s 289 862 479 1088 0 FreeSans 44 0 0 0 E
port 2 nsew
flabel metal1 s 354 1336 394 1421 0 FreeSans 44 0 0 0 B
port 3 nsew
flabel metal1 s 477 1758 1474 1786 0 FreeSans 44 0 0 0 C
port 4 nsew
<< properties >>
string GDS_END 9109982
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9086230
string gencell sky130_fd_pr__npn_11v0_W1p00L1p00
string library sky130
string parameter m=1
string path 4.450 44.925 4.450 3.825 
<< end >>
