##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 17:43:22 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RegFile
  CLASS BLOCK ;
  SIZE 240.1200 BY 219.6400 ;
  FOREIGN RegFile 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 309.824 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 472.416 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 219.3100 14.1150 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.104 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 175.136 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 270.384 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 219.3100 12.7350 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.9298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.304 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 85.696 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 132.384 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 219.3100 11.3550 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.0515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.3398 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.616 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 219.3100 10.4350 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.0405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.7552 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.576 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 219.3100 25.1550 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 219.3100 23.7750 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.8533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.0955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.759 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.208 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 166.288 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 253.272 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 219.3100 22.3950 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 219.3100 21.0150 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.388 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.8625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.142 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 219.3100 19.6350 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 21.9603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 109.631 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 51.9048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 277.296 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 219.3100 18.2550 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 257.92 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 390.72 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 219.3100 16.8750 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.757 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.504 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 86.464 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 133.536 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 219.3100 15.4950 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.5999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.7896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 219.3100 35.7350 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 26.5462 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 132.654 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.8216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.99 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 219.3100 34.3550 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.6596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 233.792 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 219.3100 33.4350 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 219.3100 32.0550 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 23.2912 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 116.379 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 219.3100 30.6750 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 176.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 269.328 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 219.3100 29.2950 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.38 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 219.3100 27.9150 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.6264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.014 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 219.3100 26.5350 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 219.3100 57.3550 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.5708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 219.3100 56.4350 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.6849 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.384 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 50.032 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 78.888 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 219.3100 55.0550 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.6392 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.832 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 126.544 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 193.656 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 219.3100 53.6750 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.934 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 219.3100 52.2950 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.63 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 219.3100 50.9150 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.686 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.56 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 219.3100 49.5350 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 219.3100 48.1550 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.388 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 219.3100 46.7750 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.866 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 219.3100 45.3950 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 24.7528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 123.687 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 219.3100 44.0150 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.6008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.216 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 75.424 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 116.976 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 219.3100 42.6350 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.9987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.8225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 219.3100 41.2550 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4184 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.502 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 219.3100 39.8750 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3772 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.414 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 219.3100 38.4950 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.842 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 219.3100 37.1150 219.6400 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.8728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.722 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 219.3100 79.4350 219.6400 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 214.528 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 325.632 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 219.3100 78.0550 219.6400 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.6084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 219.3100 76.6750 219.6400 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.7878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 197.88 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 37.888 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 60.672 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 219.3100 75.2950 219.6400 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 219.3100 73.9150 219.6400 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.558 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 219.3100 72.5350 219.6400 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 219.3100 71.1550 219.6400 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.092 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 85.3825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.6578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 219.3100 69.7750 219.6400 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.202 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 219.3100 68.3950 219.6400 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.148 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 219.3100 67.0150 219.6400 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.4898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.416 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 219.3100 65.6350 219.6400 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 219.3100 64.2550 219.6400 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.3288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.526 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 219.3100 62.8750 219.6400 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.9352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.558 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 219.3100 61.4950 219.6400 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.7438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.312 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 148.288 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 226.272 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 219.3100 60.1150 219.6400 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.0088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.392 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 65.64 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 219.3100 58.7350 219.6400 ;
    END
  END NN4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.7641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.189 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0991 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 0.0000 14.1150 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.4062 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 142.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.3516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.816 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 0.0000 12.7350 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.9238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 49.272 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.872 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 140.56 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 214.68 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 0.0000 11.3550 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.281 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7488 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.3905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.555 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.9298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.4836 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.3035 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7488 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.9266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.709 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 17.8044 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.5421 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 0.0000 25.1550 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.6199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.8776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 86.3143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 460.279 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 0.0000 23.7750 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.7488 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 298 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 450.84 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 443.362 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 824.778 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 0.0000 22.3950 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.2888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.552 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.5616 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 125.104 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 191.496 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 189.18 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 356.766 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 0.0000 21.0150 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.788 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.8625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.8018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.9398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.4521 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 123.319 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 0.0000 19.6350 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.1705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.739 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.567 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 351.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 0.0000 18.2550 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 22.7595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.508 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.5448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.9028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 13.4927 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 70.0256 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 0.0000 16.8750 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 17.2675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.1665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8227 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.1219 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 154.119 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.62605 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.913 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.296 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.1376 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 128.416 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 196.464 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 0.0000 35.7350 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.708 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4255 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.9195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 26.4232 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 141.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 0.0000 34.3550 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5273 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 0.0000 33.4350 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.0587 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 296.464 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 0.0000 32.0550 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.8648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.624 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.5048 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 209.68 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 318.36 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 0.0000 30.6750 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 12.4023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.7225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.0998 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6531 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.696 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.5048 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 34.576 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 55.704 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 0.0000 29.2950 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4565 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 0.0000 27.9150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.2016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.1889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.0855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.264 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 0.0000 26.5350 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.6338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 233.184 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 67.2198 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 356.221 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 0.0000 57.3550 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.0136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 75.2454 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 401.038 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 21.4996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 107.384 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.636 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.34094 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.0189 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.2308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4568 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 343.239 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0593 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.1108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 74.4028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.791 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.4375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.017 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 4.04296 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 19.6215 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.0092 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.472 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 107.44 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 165 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 176.513 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 384.392 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 0.0000 49.5350 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.974 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.7925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 20.043 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.4795 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 0.0000 48.1550 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.94 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.11758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.2842 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 0.0000 46.7750 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.8139 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.8985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.5658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.5738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.424 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 62.512 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 97.608 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 104.209 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 232.917 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 0.0000 45.3950 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9167 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 48.928 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 79.8672 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 168.836 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 0.0000 44.0150 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.9758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 65.8587 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 347.972 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 0.0000 42.6350 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.9606 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 0.0000 41.2550 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.7908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.688 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 0.0000 39.8750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.952 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.1304 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 114.064 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 174.936 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 0.0000 38.4950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8015 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.544 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 0.0000 37.1150 0.3300 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 29.3508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 146.636 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 40.4037 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 199.63 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 0.0000 79.4350 0.3300 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.8798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 476.382 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 0.0000 78.0550 0.3300 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.7465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 88.3422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 471.216 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 0.0000 76.6750 0.3300 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.7032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.632 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.9837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.297 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 0.0000 75.2950 0.3300 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.358 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 26.6403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 132.913 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.52512 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.8909 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 25.366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 35.0373 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 173.474 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.66 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 83.5127 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 441.993 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.956 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.2838 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.628 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 293.15 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2142 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.252 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.2192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 23.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.174 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 32.3033 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 160.054 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.5306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.312 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 30.16 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 49.08 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 107.988 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 417.389 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.2692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.834 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.18916 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.1919 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.5666 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.504 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 179.552 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 277.008 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 253.535 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 427.917 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.2854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.63 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.9275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.4674 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 81.403 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 0.0000 61.4950 0.3300 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 27.6104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 137.721 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0675 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 0.0000 60.1150 0.3300 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.31705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.373 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.7216 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.4935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.7587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.8408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.288 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 0.0000 58.7350 0.3300 ;
    END
  END NN4END[0]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.813 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.1068 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 84.7600 240.1200 84.9000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 83.4000 240.1200 83.5400 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7196 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.437 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.105 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.32 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 81.7000 240.1200 81.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3094 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.386 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.8898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.216 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 80.3400 240.1200 80.4800 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.4305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 96.6600 240.1200 96.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7211 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.3265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.7968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.72 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 94.9600 240.1200 95.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 93.6000 240.1200 93.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 92.2400 240.1200 92.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.1916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 90.5400 240.1200 90.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.942 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 89.1800 240.1200 89.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.59 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 87.8200 240.1200 87.9600 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.8685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 86.1200 240.1200 86.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5661 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.992 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 108.2200 240.1200 108.3600 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 106.8600 240.1200 107.0000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 105.5000 240.1200 105.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 103.8000 240.1200 103.9400 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 102.4400 240.1200 102.5800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.8572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.06 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 101.0800 240.1200 101.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.0668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.368 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 72.112 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 112.008 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 99.3800 240.1200 99.5200 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.8214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.144 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 98.0200 240.1200 98.1600 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 132.0200 240.1200 132.1600 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.2038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.224 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 130.3200 240.1200 130.4600 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.9758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.008 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 128.9600 240.1200 129.1000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.346 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 127.6000 240.1200 127.7400 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.5622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.467 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 125.9000 240.1200 126.0400 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 124.5400 240.1200 124.6800 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.736 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 149.968 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 228.792 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 123.1800 240.1200 123.3200 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 279.664 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 423.336 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 121.4800 240.1200 121.6200 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.0152 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.732 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 120.1200 240.1200 120.2600 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 118.7600 240.1200 118.9000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.7726 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.637 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 117.0600 240.1200 117.2000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 253.504 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 384.096 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 115.7000 240.1200 115.8400 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.9875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 257.584 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 390.216 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 114.3400 240.1200 114.4800 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.9546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.24 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 266.752 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 403.968 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 112.6400 240.1200 112.7800 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.668 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.061 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.3048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.304 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 257.92 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 390.72 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 111.2800 240.1200 111.4200 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 109.9200 240.1200 110.0600 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4879 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.0618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.8 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 149.7000 240.1200 149.8400 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 148.0000 240.1200 148.1400 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 146.6400 240.1200 146.7800 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.216 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 145.2800 240.1200 145.4200 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.868 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 143.5800 240.1200 143.7200 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 142.2200 240.1200 142.3600 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.128 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 87.568 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 135.192 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 140.8600 240.1200 141.0000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.0448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.998 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 139.1600 240.1200 139.3000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.806 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.103 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.9726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.48 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 137.8000 240.1200 137.9400 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3367 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.163 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.0068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.048 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 258.688 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 391.872 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 136.4400 240.1200 136.5800 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 134.7400 240.1200 134.8800 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.7505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.4085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 133.3800 240.1200 133.5200 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 35.9606 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.0844 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.4233 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 373.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.7600 0.4850 84.9000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.9067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.1167 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0844 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8481 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.4000 0.4850 83.5400 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.288 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.0614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.7000 0.4850 81.8400 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.475 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.3400 0.4850 80.4800 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.963 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.4716 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.707 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.6600 0.4850 96.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.936 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 19.0423 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.968 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.9600 0.4850 95.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4158 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.8178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 340.832 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 92.3756 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 488.769 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.6998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 85.8936 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 453.572 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.2400 0.4850 92.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.7138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.763 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8533 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.803 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.955 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.5688 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 175.472 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 270.888 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 243.92 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 399.234 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.1800 0.4850 89.3200 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.8958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 10.9279 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 55.1805 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.8200 0.4850 87.9600 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.6979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0925 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6799 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.4835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4974 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 66.4721 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 16.3685 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 82.4182 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.1200 0.4850 86.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.1412 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 250.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 380.28 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.4866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.813 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.5858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.5000 0.4850 105.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9504 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9504 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.5192 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.849 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.71 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.4400 0.4850 102.5800 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.455 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 109.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.264 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.7028 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 79.072 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 122.448 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.0800 0.4850 101.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.3800 0.4850 99.5200 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6076 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.877 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.0200 0.4850 98.1600 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.4488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 123.232 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 188.688 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 217.528 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 517.301 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 12.5345 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.6155 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.49212 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0296 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.9600 0.4850 129.1000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.078 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.48189 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8694 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.6000 0.4850 127.7400 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.352 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 117.724 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 623.83 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.9000 0.4850 126.0400 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.729 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.8474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.3422 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.156 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.5400 0.4850 124.6800 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1217 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.16539 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.2869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.1800 0.4850 123.3200 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.43785 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.7582 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.4800 0.4850 121.6200 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5489 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.2108 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.82175 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.9818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.34593 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 4.19596 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.0600 0.4850 117.2000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.56189 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.3785 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.7000 0.4850 115.8400 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.288 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.378 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 27.952 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 45.768 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.3400 0.4850 114.4800 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.1926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.176 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.378 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 195.76 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 297.48 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.6400 0.4850 112.7800 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.0846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.392 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.2800 0.4850 111.4200 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.1833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.6375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.5884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 211.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.5977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 62.7095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.208 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 74.32 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 115.32 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 107.717 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 188.995 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.7000 0.4850 149.8400 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 48.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 256.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 28.2514 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.269 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.0000 0.4850 148.1400 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.6077 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.409 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.6400 0.4850 146.7800 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.28 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.63596 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.6397 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.2800 0.4850 145.4200 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 21.3127 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 106.29 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.5800 0.4850 143.7200 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.22 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.528 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 112.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 173.28 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 182.798 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 390.341 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.471 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 21.1358 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.443 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.8600 0.4850 141.0000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.3322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.435 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.9174 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 62.0532 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.1600 0.4850 139.3000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.5646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.304 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.1755 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 355.545 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.8000 0.4850 137.9400 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1293 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.3922 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.1707 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 161.461 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.4400 0.4850 136.5800 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.4552 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.3818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.712 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.7400 0.4850 134.8800 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.8435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 2.4552 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.4194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.024 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 48.928 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 77.232 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.2944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.6238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.464 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.0345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.033 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.6824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 122.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.556 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 0.0000 106.1150 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 0.0000 104.7350 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.3235 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.488 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 0.0000 103.3550 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.7326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 0.0000 102.4350 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.4594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.528 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 0.0000 101.0550 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0412 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.088 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 0.0000 99.6750 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1374 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 0.0000 98.2950 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.248 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 0.0000 96.9150 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 0.0000 95.5350 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 0.0000 94.1550 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 0.0000 92.7750 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.488 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 0.0000 91.3950 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.9272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 84.5215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.71 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.432 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 0.0000 90.0150 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.448 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.1625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.1218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 225.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 0.0000 88.6350 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.9364 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 0.0000 87.2550 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.1732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.748 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.24 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 0.0000 127.7350 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.5836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 0.0000 126.3550 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.9226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.528 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 0.0000 125.4350 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.1516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 0.0000 124.0550 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.907 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.4575 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.986 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 0.0000 122.6750 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.1744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.358 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 0.0000 121.2950 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1984 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.6314 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 0.0000 119.9150 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 261.448 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 143.872 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 219.648 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 0.0000 118.5350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0492 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 210.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 0.0000 117.1550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.4696 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.2705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.202 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.892 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 0.0000 115.7750 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.2514 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 0.0000 114.3950 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.8332 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 0.0000 113.0150 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 91.8435 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 0.0000 111.6350 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7461 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 305.328 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 0.0000 110.2550 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.5772 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.8085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.77 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 0.0000 108.8750 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.0698 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.384 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 128.416 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 196.464 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 0.0000 107.4950 0.3300 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.528 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 0.0000 149.3550 0.3300 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.66385 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.781 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.0485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.3112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.438 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 0.0000 148.4350 0.3300 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.0524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.024 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 0.0000 147.0550 0.3300 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.989 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.5546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 0.0000 145.6750 0.3300 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0588 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.956 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 0.0000 144.2950 0.3300 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.0892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.3685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.006 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 0.0000 142.9150 0.3300 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.3128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.68 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 185.824 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 282.576 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 0.0000 141.5350 0.3300 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.6558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.176 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 89.008 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 137.352 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 0.0000 140.1550 0.3300 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.1749 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.6706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.184 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 0.0000 138.7750 0.3300 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.8604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 0.0000 137.3950 0.3300 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9336 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.484 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 0.0000 136.0150 0.3300 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.8494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.608 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 0.0000 134.6350 0.3300 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.6745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.3657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.6575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.332 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.5014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 0.0000 133.2550 0.3300 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.0212 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.0285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.248 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.122 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 0.0000 131.8750 0.3300 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.3814 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 0.0000 130.4950 0.3300 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2592 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.2185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2907 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.7396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 223.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 0.0000 129.1150 0.3300 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.4261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.8415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.134 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5415 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 219.3100 84.4950 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.4701 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 219.3100 83.1150 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9689 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 219.3100 81.7350 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.512 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 66.3165 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 356.976 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 219.3100 80.3550 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.0718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.5661 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 369.668 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 219.3100 106.1150 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.7919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.7465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.0898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 24.6789 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 130.234 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 219.3100 104.7350 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.0766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 190.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 59.6763 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.677 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 219.3100 103.3550 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0232 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.2546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 60.585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4653 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.1704 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 219.3100 102.4350 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.9228 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.6 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.7488 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 132.064 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 201.936 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 191.516 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 336.521 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 219.3100 101.0550 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 22.4397 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 121.588 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 219.3100 99.6750 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5115 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.13663 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.0781 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 4.58242 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 21.0842 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.76 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.5444 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 96.1818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 219.3100 98.2950 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1307 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.1306 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 336.917 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 219.3100 96.9150 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.1536 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.9717 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 219.3100 95.5350 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7849 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.4704 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 219.3100 94.1550 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5721 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.897 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.424 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 219.3100 92.7750 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1922 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.456 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 219.3100 91.3950 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.8462 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 92 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.5192 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 109.648 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 168.312 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 219.3100 90.0150 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5048 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 219.3100 88.6350 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.5858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.136 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.5012 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 41.2 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 65.64 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 219.3100 87.2550 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5084 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.7084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.856 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 219.3100 85.8750 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.6192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.456 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 131.728 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 201.432 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 215.27 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 466.54 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 219.3100 127.7350 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.8818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.0753 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 388.075 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 219.3100 126.3550 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5672 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.7585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.7 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.99293 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.5764 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 219.3100 125.4350 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.056 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4934 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.6559 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 219.3100 124.0550 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.8892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 64.3685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2656 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.21 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.15327 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.4626 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 219.3100 122.6750 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.0916 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.304 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 78.736 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 121.944 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 122.935 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 248.176 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 219.3100 121.2950 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.18405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.0856 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.3505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3276 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.52 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.26923 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.9515 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 219.3100 119.9150 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.6484 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.1645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.3432 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.598 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.0609 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.5138 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 219.3100 118.5350 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.1944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.8945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.928 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.13724 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.2916 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 219.3100 117.1550 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.4488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.63 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.3941 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.5758 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 219.3100 115.7750 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.196 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.7094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 219.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 57.76 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 90.48 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 97.8304 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 222.675 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 219.3100 114.3950 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.0644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.6051 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 164.134 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 219.3100 113.0150 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.5137 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.1615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9834 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 219.3100 111.6350 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.95285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.4138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.552 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.1376 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 57.76 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 90.48 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 219.3100 110.2550 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8289 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 219.3100 108.8750 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.7536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0586 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 219.3100 107.4950 219.6400 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.398 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.916 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 21.0343 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 103.941 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 219.3100 149.3550 219.6400 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.1825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.0608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.3941 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 309.811 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 219.3100 148.4350 219.6400 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.3595 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.969 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 219.3100 147.0550 219.6400 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.5432 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 82.6385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.68855 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6519 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 219.3100 145.6750 219.6400 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 11.8585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 60.6613 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 219.3100 144.2950 219.6400 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.318 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.668 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.04397 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.27 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 219.3100 142.9150 219.6400 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2473 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.41525 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.672 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 52.576 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 82.704 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 147.27 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 515.801 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 219.3100 141.5350 219.6400 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2734 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 24.8723 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 130.603 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 219.3100 140.1550 219.6400 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.1948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.99 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.714 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.43529 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.7138 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 219.3100 138.7750 219.6400 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.1634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 199.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 59.6114 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 315.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 219.3100 137.3950 219.6400 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0704 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.79232 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 7.567 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 219.3100 136.0150 219.6400 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.0028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.8995 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5272 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.13582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 219.3100 134.6350 219.6400 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.853 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 219.3100 133.2550 219.6400 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.1397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 219.3100 131.8750 219.6400 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.4242 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 71.9355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.8023 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.7225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.0124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 219.3100 130.4950 219.6400 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3744 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.2965 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.744 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.5616 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 68.8 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 107.04 LAYER met5  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 219.3100 129.1150 219.6400 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.3008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.616 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 222.256 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 337.224 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.631 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.84 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.6862 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.6800 0.4850 12.8200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.879 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.04 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.3200 0.4850 11.4600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.969 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.8584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 208.656 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.9600 0.4850 10.1000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.242 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 148.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.1306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.512 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 78.736 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 121.944 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.5800 0.4850 24.7200 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.364 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.8800 0.4850 23.0200 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.2848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.656 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.5200 0.4850 21.6600 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.23 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.7358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 340.96 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 515.28 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.718 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.878 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 239.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.0958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.856 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 85.36 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 131.88 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.1000 0.4850 17.2400 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.4638 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.944 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.22 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.8400 0.4850 37.9800 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.0108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 290.704 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 439.896 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.55 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.6578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.52 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 339.952 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 513.768 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.7800 0.4850 34.9200 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2954 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.316 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.1914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.4200 0.4850 33.5600 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 256.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.7200 0.4850 31.8600 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.7664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.04 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 36.784 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 59.016 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.3600 0.4850 30.5000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.0000 0.4850 29.1400 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.391 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 155.248 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 236.712 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.3000 0.4850 61.4400 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4229 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.4528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.0102 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.2400 0.4850 58.3800 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.439 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 49.0258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 262.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.712 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 26.848 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 44.112 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.8800 0.4850 57.0200 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.834 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.692 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.8200 0.4850 53.9600 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.3996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.772 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7388 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.468 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.1000 0.4850 51.2400 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.4000 0.4850 49.5400 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.0400 0.4850 48.1800 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.604 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.794 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.343 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.4197 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.408 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 19.12 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.9800 0.4850 45.1200 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3906 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.792 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 229.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 35.4216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.856 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.2600 0.4850 42.4000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.3486 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 47.521 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 253.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.144 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 36.784 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 59.016 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.2000 0.4850 39.3400 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 37.864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 202.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.9800 0.4850 79.1200 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.009 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 53.359 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 285.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.6200 0.4850 77.7600 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.976 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 272.608 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 412.752 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.9200 0.4850 76.0600 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.038 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.5600 0.4850 74.7000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.2000 0.4850 73.3400 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.45 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.368 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 289.6 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 438.24 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.5000 0.4850 71.6400 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.132 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.4616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.082 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.7800 0.4850 68.9200 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.7956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.634 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.7200 0.4850 65.8600 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 32.158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.9706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.992 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 56.656 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 88.824 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.3600 0.4850 64.5000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 231.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.6600 0.4850 62.8000 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1267 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.792 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3212 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5403 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.432 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.07 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 63.28 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 98.76 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 14.0400 240.1200 14.1800 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.07 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.6664 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 353.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 12.6800 240.1200 12.8200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 69.7248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 374.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 11.3200 240.1200 11.4600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.7486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0477 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.8076 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.184 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 9.9600 240.1200 10.1000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 30.9287 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 157.712 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.261145 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 25.9400 240.1200 26.0800 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.1521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.3735 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 15.5999 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.2424 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.416 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 28.3471 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 145.49 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 29.2465 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.92 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 24.5800 240.1200 24.7200 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.7538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.5838 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 154.509 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.183704 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 22.8800 240.1200 23.0200 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.427 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.3028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.96 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.5616 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 44.512 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 70.608 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 106.667 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 339.195 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 21.5200 240.1200 21.6600 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.2696 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.444 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.4454 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.7737 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 20.1600 240.1200 20.3000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.8007 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 431.913 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.284714 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 18.4600 240.1200 18.6000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1281 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.7518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.688 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.7632 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 55.552 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 87.168 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 132.157 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 407.483 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 17.1000 240.1200 17.2400 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0078 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.76 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.8122 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.88 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.2154 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.904 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 15.7400 240.1200 15.8800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.5306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 37.8400 240.1200 37.9800 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.168 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 36.1400 240.1200 36.2800 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.62 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.7104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 181.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 34.7800 240.1200 34.9200 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.219 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.4 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.5156 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 75.424 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 116.976 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 33.4200 240.1200 33.5600 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.7028 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.1295 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 54.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 31.7200 240.1200 31.8600 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3284 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.4248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 30.3600 240.1200 30.5000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.237 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1412 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 29.0000 240.1200 29.1400 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6027 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3104 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 27.3000 240.1200 27.4400 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.1672 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.44 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.3102 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.952 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 61.3000 240.1200 61.4400 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 20.1518 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 106.993 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 59.9400 240.1200 60.0800 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.457 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.721 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.9882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.424 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 75.424 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 116.976 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 149.589 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 405.096 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 58.2400 240.1200 58.3800 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.853 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.705 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 9.00485 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 49.4141 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 56.8800 240.1200 57.0200 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.4109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.6575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 104.128 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 160.032 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 168.8 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 360.808 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 55.5200 240.1200 55.6600 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.748 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.514 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.41576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.62963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 53.8200 240.1200 53.9600 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.83 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.409 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 97.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 52.4600 240.1200 52.6000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.68687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.9535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 51.1000 240.1200 51.2400 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.264 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.26195 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.7697 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 49.4000 240.1200 49.5400 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.85468 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8424 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 48.0400 240.1200 48.1800 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.38364 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.2458 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 46.6800 240.1200 46.8200 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.748 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.514 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 1.41576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 5.62963 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 44.9800 240.1200 45.1200 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.751 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.17 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 63.912 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.378 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 58.864 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 92.136 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 43.6200 240.1200 43.7600 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2537 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.957 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 0.378 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 59.968 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 93.792 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 42.2600 240.1200 42.4000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.5496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.872 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 40.5600 240.1200 40.7000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.11 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 39.2000 240.1200 39.3400 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.315 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.4307 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.6135 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 78.9800 240.1200 79.1200 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.23 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.2824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.5051 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 77.6200 240.1200 77.7600 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.843 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.633 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.2036 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.568 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 76.528 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 118.632 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 146.466 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 388.665 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 75.9200 240.1200 76.0600 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.81818 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 43.5596 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 74.5600 240.1200 74.7000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7185 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.07751 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.9448 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 73.2000 240.1200 73.3400 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.1534 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.6547 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.751 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 71.5000 240.1200 71.6400 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.82 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.6162 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 101.168 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.1749 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.865 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 70.1400 240.1200 70.2800 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 14.8187 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 76.536 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 68.7800 240.1200 68.9200 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.853 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.473 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 70.666 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 67.0800 240.1200 67.2200 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.086 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8694 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.6545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 65.7200 240.1200 65.8600 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0592 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.1694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 170 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 64.3600 240.1200 64.5000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.12 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.439 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.323 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8003 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.216 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.0592 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 88.672 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 136.848 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 62.6600 240.1200 62.8000 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.0424 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 140.096 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 201.28 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 305.76 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met5  ;
    ANTENNAMAXAREACAR 52.3 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 110.664 LAYER met5  ;
    PORT
      LAYER met4 ;
        RECT 89.5500 0.0000 89.8500 0.8000 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 217.476 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met2  ;
    ANTENNAMAXAREACAR 42.4854 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 207.238 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.5400 0.4850 209.6800 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 45.8767 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 229.835 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.562875 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.8400 0.4850 207.9800 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.276 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met2  ;
    ANTENNAMAXAREACAR 33.1721 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.506709 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 34.5317 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 167.595 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.548637 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.1567 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.968 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 38.5027 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.94 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.1400 0.4850 206.2800 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4939 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.2024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.032 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 44.512 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 70.608 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 100.745 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 471.847 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.4400 0.4850 204.5800 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 65.7882 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 355.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 57.6107 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 305.58 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.7400 0.4850 202.8800 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.141 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.8694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met4  ;
    ANTENNAMAXAREACAR 55.7653 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.437 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 1.53396 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 65.488 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 102.072 LAYER met5  ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 143.209 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 665.099 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 201.0400 0.4850 201.1800 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.5248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.144 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 47.824 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 75.576 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 64.7679 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 267.987 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 199.0000 0.4850 199.1400 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.605 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.9479 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 79.9206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.737 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.3000 0.4850 197.4400 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 39.3978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 67.7476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 355.333 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.09371 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.6000 0.4850 195.7400 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.17 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.175 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.8099 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 52.7934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.339 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.08323 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.9000 0.4850 194.0400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.427 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.096 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 56.656 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 88.824 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 70.0435 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 286.731 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.2000 0.4850 192.3400 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.233 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.0978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 77.304 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.186 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.1600 0.4850 190.3000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.913 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 51.136 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 80.544 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 74.5703 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 310.329 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.4600 0.4850 188.6000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.5558 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.976 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 161.888 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 250.512 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 93.425 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 265.902 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.7600 0.4850 186.9000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.282 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0605 LAYER met2  ;
    ANTENNAMAXAREACAR 26.4191 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.681725 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.928 LAYER met3  ;
    ANTENNAGATEAREA 1.0605 LAYER met3  ;
    ANTENNAMAXAREACAR 26.7784 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 129.716 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.757162 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.5576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 38.4648 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.695 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.757162 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 185.0600 0.4850 185.2000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1757 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.3833 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.296 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 26.0793 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 128.522 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.551831 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.0192 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.984 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0671 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.404 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.3600 0.4850 183.5000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.4432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.096 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 60.6445 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 306.513 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.03082 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.088 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 68.4672 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 348.9 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.03082 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.3200 0.4850 181.4600 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.382 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.1023 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 96.3026 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 502.684 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.6200 0.4850 179.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8453 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 36.9266 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 179.342 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 40.3763 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 198.474 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.732075 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.1962 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.8 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 75.2017 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 397.696 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.9200 0.4850 178.0600 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.9302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.33 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2904 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.941 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.648218 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.77 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.24 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 35.4832 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.459 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 28.5867 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.28 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 72.4857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 375.188 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.2200 0.4850 176.3600 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.917 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.2675 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 64.6751 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.89 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.5200 0.4850 174.6600 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.6396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.005 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met2  ;
    ANTENNAMAXAREACAR 32.9272 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 159.151 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.515094 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 33.9511 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 165.199 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.565409 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.9854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 108 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0646 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.64 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.4800 0.4850 172.6200 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.136 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.0198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.784 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 82.048 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 126.912 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 118.568 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 501.432 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.7800 0.4850 170.9200 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.0767 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 200.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 42.6504 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.773 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 169.0800 0.4850 169.2200 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5409 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4255 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.1782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 48.5357 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.243 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00764 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.3800 0.4850 167.5200 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.5075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6965 LAYER met2  ;
    ANTENNAMAXAREACAR 28.5243 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 137.932 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.488358 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.032 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.304 LAYER met3  ;
    ANTENNAGATEAREA 1.6965 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7221 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 144.595 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.511936 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 55.6242 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.693 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.807547 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.6800 0.4850 165.8200 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.4985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.728 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 98.1975 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 504.199 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.87673 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5861 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.608 LAYER met4  ;
    ANTENNAGATEAREA 0.954 LAYER met4  ;
    ANTENNAMAXAREACAR 110.342 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 565.633 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 1.54759 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 27.952 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 45.768 LAYER met5  ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 120.291 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 581.923 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.6400 0.4850 163.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2261 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.979 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0729 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 149.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 55.4746 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 287.523 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.9400 0.4850 162.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.6758 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 159.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 81.2562 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 423.419 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80 LAYER met4  ;
    ANTENNAGATEAREA 1.8555 LAYER met4  ;
    ANTENNAMAXAREACAR 89.615 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 466.534 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 1.17134 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 97.856 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 154.464 LAYER met5  ;
    ANTENNAGATEAREA 2.8095 LAYER met5  ;
    ANTENNAMAXAREACAR 124.445 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 521.514 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.2400 0.4850 160.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.257 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 79.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.8095 LAYER met4  ;
    ANTENNAMAXAREACAR 38.2027 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 189.789 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.5400 0.4850 158.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.018 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.747 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.9417 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met4  ;
    ANTENNAMAXAREACAR 68.025 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 353.581 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.8400 0.4850 156.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.451 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3924 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.776 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 73.216 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 113.664 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6505 LAYER met5  ;
    ANTENNAMAXAREACAR 72.0469 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 264.251 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.1400 0.4850 155.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.276 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 209.5400 240.1200 209.6800 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5358 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.9286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 207.8400 240.1200 207.9800 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.3691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.6195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 206.1400 240.1200 206.2800 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.043 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.976 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 204.4400 240.1200 204.5800 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.385 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 202.7400 240.1200 202.8800 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6869 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3265 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 201.0400 240.1200 201.1800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.261 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 199.0000 240.1200 199.1400 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.339 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 197.3000 240.1200 197.4400 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.459 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.4824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 293.192 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 80.944 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 125.256 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 195.6000 240.1200 195.7400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.0515 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.862 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.1406 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 183.024 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 193.9000 240.1200 194.0400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 15.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 192.2000 240.1200 192.3400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 190.1600 240.1200 190.3000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 188.4600 240.1200 188.6000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.704 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 186.7600 240.1200 186.9000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.944 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 185.0600 240.1200 185.2000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.767 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.373 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 183.3600 240.1200 183.5000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.701 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.872 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.4422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 181.3200 240.1200 181.4600 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.265 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 179.6200 240.1200 179.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 177.9200 240.1200 178.0600 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 176.2200 240.1200 176.3600 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 174.5200 240.1200 174.6600 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.322 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 172.4800 240.1200 172.6200 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.2308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 220.368 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 170.7800 240.1200 170.9200 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 169.0800 240.1200 169.2200 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.6628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 206.672 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 167.3800 240.1200 167.5200 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.45345 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 22.432 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 37.488 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 165.6800 240.1200 165.8200 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7126 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.337 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 163.6400 240.1200 163.7800 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.207 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 161.9400 240.1200 162.0800 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.6463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.9525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.7458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 160.2400 240.1200 160.3800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.503 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.0746 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.88 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 1.782 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 76.528 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 118.632 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 158.5400 240.1200 158.6800 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.8058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 156.8400 240.1200 156.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6486 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.017 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 155.1400 240.1200 155.2800 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.17104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.3152 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.9200 0.0000 210.0600 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.521 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.689 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.9526 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.0828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 405.368 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 206.7000 0.0000 206.8400 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.6628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 335.88 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 6.976 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 14.304 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 12.1223 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 27.9589 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 203.9400 0.0000 204.0800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5428 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.553 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.2024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.032 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 90.88 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 140.16 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met5  ;
    ANTENNAMAXAREACAR 184.488 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 511.045 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 201.1800 0.0000 201.3200 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.215 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.914 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.7676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.4831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 386.652 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 197.5000 0.0000 197.6400 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.9099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 124.324 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 34.423 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 170.575 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 195.2000 0.0000 195.3400 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.283 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.633 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.7318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.1439 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 402.725 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 192.4400 0.0000 192.5800 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.044 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.655 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 25.8414 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.9665 LAYER met4  ;
    ANTENNAMAXAREACAR 48.738 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 242.775 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 0.0000 189.8200 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.7958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.18 LAYER met3  ;
    ANTENNAMAXAREACAR 23.0772 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 109.34 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.684277 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.6998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.536 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.3727 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 132.339 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.684277 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 186.4600 0.0000 186.6000 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1826 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.752 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 105.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 28.9334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.646 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.693657 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 183.7000 0.0000 183.8400 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9638 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.292 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.6275 LAYER met2  ;
    ANTENNAMAXAREACAR 33.7275 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 157.102 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.671118 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAGATEAREA 1.6275 LAYER met3  ;
    ANTENNAMAXAREACAR 36.5595 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 172.492 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.695696 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.4443 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.776 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.9143 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.318 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.695696 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 180.9400 0.0000 181.0800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.0446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 30.2999 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.345 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.681884 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 178.1800 0.0000 178.3200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.3948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 38.7256 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 190.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.645305 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.9600 0.0000 175.1000 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 29.6216 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 147.152 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.870881 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.2000 0.0000 172.3400 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3286 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.482 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.9209 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 41.7065 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 169.4400 0.0000 169.5800 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.847 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9505 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.5181 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.709434 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.112 LAYER met3  ;
    ANTENNAGATEAREA 2.544 LAYER met3  ;
    ANTENNAMAXAREACAR 21.6771 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 105.101 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.725157 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.136 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 41.848 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 207.982 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.730948 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 166.2200 0.0000 166.3600 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.366 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.8146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.5408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.6485 LAYER met4  ;
    ANTENNAMAXAREACAR 45.2212 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.921 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 1.08988 LAYER via4  ;
    ANTENNAPARTIALMETALAREA 131.728 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 201.432 LAYER met5  ;
    ANTENNAGATEAREA 5.2845 LAYER met5  ;
    ANTENNAMAXAREACAR 70.1484 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 272.039 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 163.4600 0.0000 163.6000 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.327 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 37.1396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 179.294 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.232 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 39.4289 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.237 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.732075 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.0139 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 285.088 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 49.4609 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 246.185 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 160.7000 0.0000 160.8400 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.6877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.8485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1815 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 108.994 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.669182 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.7253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.12 LAYER met3  ;
    ANTENNAGATEAREA 1.908 LAYER met3  ;
    ANTENNAMAXAREACAR 31.9044 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 155.051 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.690147 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.6138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 247.968 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 46.1593 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.612 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.9400 0.0000 158.0800 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.044 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 24.3181 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.894 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.677803 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 0.0000 155.3200 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.665 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.046 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.0226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.9200 219.1550 210.0600 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0758 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.982 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.52 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 206.7000 219.1550 206.8400 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 203.9400 219.1550 204.0800 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5254 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.348 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.165 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 201.1800 219.1550 201.3200 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 197.9600 219.1550 198.1000 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.817 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.831 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.7822 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.72 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 195.2000 219.1550 195.3400 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.3075 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.4400 219.1550 192.5800 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.8894 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 123.488 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 219.1550 189.8200 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.2823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.4600 219.1550 186.6000 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.9955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 104.752 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 183.7000 219.1550 183.8400 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.8523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.0355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.9400 219.1550 181.0800 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 178.1800 219.1550 178.3200 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.9600 219.1550 175.1000 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.986 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.4798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.696 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 172.2000 219.1550 172.3400 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1845 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.9800 219.1550 169.1200 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.6800 219.1550 166.8200 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.0235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.4600 219.1550 163.6000 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7685 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 160.7000 219.1550 160.8400 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1515 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 157.4800 219.1550 157.6200 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.8223 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.8855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 219.1550 155.3200 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 234.5600 8.4300 ;
        RECT 5.5600 210.5300 234.5600 213.5300 ;
        RECT 5.5600 12.3400 8.5600 12.8200 ;
        RECT 5.5600 17.7800 8.5600 18.2600 ;
        RECT 55.1200 17.7800 56.1200 18.2600 ;
        RECT 55.1200 12.3400 56.1200 12.8200 ;
        RECT 5.5600 23.2200 8.5600 23.7000 ;
        RECT 5.5600 34.1000 8.5600 34.5800 ;
        RECT 5.5600 28.6600 8.5600 29.1400 ;
        RECT 5.5600 39.5400 8.5600 40.0200 ;
        RECT 5.5600 44.9800 8.5600 45.4600 ;
        RECT 55.1200 34.1000 56.1200 34.5800 ;
        RECT 55.1200 28.6600 56.1200 29.1400 ;
        RECT 55.1200 23.2200 56.1200 23.7000 ;
        RECT 55.1200 44.9800 56.1200 45.4600 ;
        RECT 55.1200 39.5400 56.1200 40.0200 ;
        RECT 100.1200 17.7800 101.1200 18.2600 ;
        RECT 100.1200 12.3400 101.1200 12.8200 ;
        RECT 100.1200 34.1000 101.1200 34.5800 ;
        RECT 100.1200 28.6600 101.1200 29.1400 ;
        RECT 100.1200 23.2200 101.1200 23.7000 ;
        RECT 100.1200 44.9800 101.1200 45.4600 ;
        RECT 100.1200 39.5400 101.1200 40.0200 ;
        RECT 5.5600 55.8600 8.5600 56.3400 ;
        RECT 5.5600 50.4200 8.5600 50.9000 ;
        RECT 5.5600 61.3000 8.5600 61.7800 ;
        RECT 5.5600 72.1800 8.5600 72.6600 ;
        RECT 5.5600 66.7400 8.5600 67.2200 ;
        RECT 5.5600 77.6200 8.5600 78.1000 ;
        RECT 55.1200 61.3000 56.1200 61.7800 ;
        RECT 55.1200 55.8600 56.1200 56.3400 ;
        RECT 55.1200 50.4200 56.1200 50.9000 ;
        RECT 55.1200 77.6200 56.1200 78.1000 ;
        RECT 55.1200 72.1800 56.1200 72.6600 ;
        RECT 55.1200 66.7400 56.1200 67.2200 ;
        RECT 5.5600 83.0600 8.5600 83.5400 ;
        RECT 5.5600 93.9400 8.5600 94.4200 ;
        RECT 5.5600 88.5000 8.5600 88.9800 ;
        RECT 5.5600 99.3800 8.5600 99.8600 ;
        RECT 5.5600 104.8200 8.5600 105.3000 ;
        RECT 55.1200 93.9400 56.1200 94.4200 ;
        RECT 55.1200 88.5000 56.1200 88.9800 ;
        RECT 55.1200 83.0600 56.1200 83.5400 ;
        RECT 55.1200 104.8200 56.1200 105.3000 ;
        RECT 55.1200 99.3800 56.1200 99.8600 ;
        RECT 100.1200 61.3000 101.1200 61.7800 ;
        RECT 100.1200 55.8600 101.1200 56.3400 ;
        RECT 100.1200 50.4200 101.1200 50.9000 ;
        RECT 100.1200 77.6200 101.1200 78.1000 ;
        RECT 100.1200 72.1800 101.1200 72.6600 ;
        RECT 100.1200 66.7400 101.1200 67.2200 ;
        RECT 100.1200 93.9400 101.1200 94.4200 ;
        RECT 100.1200 88.5000 101.1200 88.9800 ;
        RECT 100.1200 83.0600 101.1200 83.5400 ;
        RECT 100.1200 104.8200 101.1200 105.3000 ;
        RECT 100.1200 99.3800 101.1200 99.8600 ;
        RECT 145.1200 17.7800 146.1200 18.2600 ;
        RECT 145.1200 12.3400 146.1200 12.8200 ;
        RECT 145.1200 34.1000 146.1200 34.5800 ;
        RECT 145.1200 28.6600 146.1200 29.1400 ;
        RECT 145.1200 23.2200 146.1200 23.7000 ;
        RECT 145.1200 44.9800 146.1200 45.4600 ;
        RECT 145.1200 39.5400 146.1200 40.0200 ;
        RECT 190.1200 17.7800 191.1200 18.2600 ;
        RECT 190.1200 12.3400 191.1200 12.8200 ;
        RECT 231.5600 17.7800 234.5600 18.2600 ;
        RECT 231.5600 12.3400 234.5600 12.8200 ;
        RECT 190.1200 34.1000 191.1200 34.5800 ;
        RECT 190.1200 28.6600 191.1200 29.1400 ;
        RECT 190.1200 23.2200 191.1200 23.7000 ;
        RECT 190.1200 44.9800 191.1200 45.4600 ;
        RECT 190.1200 39.5400 191.1200 40.0200 ;
        RECT 231.5600 23.2200 234.5600 23.7000 ;
        RECT 231.5600 28.6600 234.5600 29.1400 ;
        RECT 231.5600 34.1000 234.5600 34.5800 ;
        RECT 231.5600 44.9800 234.5600 45.4600 ;
        RECT 231.5600 39.5400 234.5600 40.0200 ;
        RECT 145.1200 61.3000 146.1200 61.7800 ;
        RECT 145.1200 55.8600 146.1200 56.3400 ;
        RECT 145.1200 50.4200 146.1200 50.9000 ;
        RECT 145.1200 77.6200 146.1200 78.1000 ;
        RECT 145.1200 72.1800 146.1200 72.6600 ;
        RECT 145.1200 66.7400 146.1200 67.2200 ;
        RECT 145.1200 93.9400 146.1200 94.4200 ;
        RECT 145.1200 88.5000 146.1200 88.9800 ;
        RECT 145.1200 83.0600 146.1200 83.5400 ;
        RECT 145.1200 104.8200 146.1200 105.3000 ;
        RECT 145.1200 99.3800 146.1200 99.8600 ;
        RECT 190.1200 61.3000 191.1200 61.7800 ;
        RECT 190.1200 55.8600 191.1200 56.3400 ;
        RECT 190.1200 50.4200 191.1200 50.9000 ;
        RECT 190.1200 77.6200 191.1200 78.1000 ;
        RECT 190.1200 72.1800 191.1200 72.6600 ;
        RECT 190.1200 66.7400 191.1200 67.2200 ;
        RECT 231.5600 55.8600 234.5600 56.3400 ;
        RECT 231.5600 50.4200 234.5600 50.9000 ;
        RECT 231.5600 61.3000 234.5600 61.7800 ;
        RECT 231.5600 77.6200 234.5600 78.1000 ;
        RECT 231.5600 72.1800 234.5600 72.6600 ;
        RECT 231.5600 66.7400 234.5600 67.2200 ;
        RECT 190.1200 93.9400 191.1200 94.4200 ;
        RECT 190.1200 88.5000 191.1200 88.9800 ;
        RECT 190.1200 83.0600 191.1200 83.5400 ;
        RECT 190.1200 104.8200 191.1200 105.3000 ;
        RECT 190.1200 99.3800 191.1200 99.8600 ;
        RECT 231.5600 83.0600 234.5600 83.5400 ;
        RECT 231.5600 88.5000 234.5600 88.9800 ;
        RECT 231.5600 93.9400 234.5600 94.4200 ;
        RECT 231.5600 104.8200 234.5600 105.3000 ;
        RECT 231.5600 99.3800 234.5600 99.8600 ;
        RECT 5.5600 115.7000 8.5600 116.1800 ;
        RECT 5.5600 110.2600 8.5600 110.7400 ;
        RECT 5.5600 121.1400 8.5600 121.6200 ;
        RECT 5.5600 132.0200 8.5600 132.5000 ;
        RECT 5.5600 126.5800 8.5600 127.0600 ;
        RECT 5.5600 137.4600 8.5600 137.9400 ;
        RECT 55.1200 121.1400 56.1200 121.6200 ;
        RECT 55.1200 115.7000 56.1200 116.1800 ;
        RECT 55.1200 110.2600 56.1200 110.7400 ;
        RECT 55.1200 137.4600 56.1200 137.9400 ;
        RECT 55.1200 132.0200 56.1200 132.5000 ;
        RECT 55.1200 126.5800 56.1200 127.0600 ;
        RECT 5.5600 142.9000 8.5600 143.3800 ;
        RECT 5.5600 153.7800 8.5600 154.2600 ;
        RECT 5.5600 148.3400 8.5600 148.8200 ;
        RECT 5.5600 159.2200 8.5600 159.7000 ;
        RECT 5.5600 164.6600 8.5600 165.1400 ;
        RECT 55.1200 153.7800 56.1200 154.2600 ;
        RECT 55.1200 148.3400 56.1200 148.8200 ;
        RECT 55.1200 142.9000 56.1200 143.3800 ;
        RECT 55.1200 164.6600 56.1200 165.1400 ;
        RECT 55.1200 159.2200 56.1200 159.7000 ;
        RECT 100.1200 121.1400 101.1200 121.6200 ;
        RECT 100.1200 115.7000 101.1200 116.1800 ;
        RECT 100.1200 110.2600 101.1200 110.7400 ;
        RECT 100.1200 137.4600 101.1200 137.9400 ;
        RECT 100.1200 132.0200 101.1200 132.5000 ;
        RECT 100.1200 126.5800 101.1200 127.0600 ;
        RECT 100.1200 153.7800 101.1200 154.2600 ;
        RECT 100.1200 148.3400 101.1200 148.8200 ;
        RECT 100.1200 142.9000 101.1200 143.3800 ;
        RECT 100.1200 164.6600 101.1200 165.1400 ;
        RECT 100.1200 159.2200 101.1200 159.7000 ;
        RECT 5.5600 175.5400 8.5600 176.0200 ;
        RECT 5.5600 170.1000 8.5600 170.5800 ;
        RECT 5.5600 180.9800 8.5600 181.4600 ;
        RECT 5.5600 191.8600 8.5600 192.3400 ;
        RECT 5.5600 186.4200 8.5600 186.9000 ;
        RECT 5.5600 197.3000 8.5600 197.7800 ;
        RECT 55.1200 180.9800 56.1200 181.4600 ;
        RECT 55.1200 175.5400 56.1200 176.0200 ;
        RECT 55.1200 170.1000 56.1200 170.5800 ;
        RECT 55.1200 197.3000 56.1200 197.7800 ;
        RECT 55.1200 191.8600 56.1200 192.3400 ;
        RECT 55.1200 186.4200 56.1200 186.9000 ;
        RECT 5.5600 202.7400 8.5600 203.2200 ;
        RECT 5.5600 208.1800 8.5600 208.6600 ;
        RECT 55.1200 208.1800 56.1200 208.6600 ;
        RECT 55.1200 202.7400 56.1200 203.2200 ;
        RECT 100.1200 180.9800 101.1200 181.4600 ;
        RECT 100.1200 175.5400 101.1200 176.0200 ;
        RECT 100.1200 170.1000 101.1200 170.5800 ;
        RECT 100.1200 197.3000 101.1200 197.7800 ;
        RECT 100.1200 191.8600 101.1200 192.3400 ;
        RECT 100.1200 186.4200 101.1200 186.9000 ;
        RECT 100.1200 208.1800 101.1200 208.6600 ;
        RECT 100.1200 202.7400 101.1200 203.2200 ;
        RECT 145.1200 121.1400 146.1200 121.6200 ;
        RECT 145.1200 115.7000 146.1200 116.1800 ;
        RECT 145.1200 110.2600 146.1200 110.7400 ;
        RECT 145.1200 137.4600 146.1200 137.9400 ;
        RECT 145.1200 132.0200 146.1200 132.5000 ;
        RECT 145.1200 126.5800 146.1200 127.0600 ;
        RECT 145.1200 153.7800 146.1200 154.2600 ;
        RECT 145.1200 148.3400 146.1200 148.8200 ;
        RECT 145.1200 142.9000 146.1200 143.3800 ;
        RECT 145.1200 164.6600 146.1200 165.1400 ;
        RECT 145.1200 159.2200 146.1200 159.7000 ;
        RECT 190.1200 121.1400 191.1200 121.6200 ;
        RECT 190.1200 115.7000 191.1200 116.1800 ;
        RECT 190.1200 110.2600 191.1200 110.7400 ;
        RECT 190.1200 137.4600 191.1200 137.9400 ;
        RECT 190.1200 132.0200 191.1200 132.5000 ;
        RECT 190.1200 126.5800 191.1200 127.0600 ;
        RECT 231.5600 115.7000 234.5600 116.1800 ;
        RECT 231.5600 110.2600 234.5600 110.7400 ;
        RECT 231.5600 121.1400 234.5600 121.6200 ;
        RECT 231.5600 137.4600 234.5600 137.9400 ;
        RECT 231.5600 132.0200 234.5600 132.5000 ;
        RECT 231.5600 126.5800 234.5600 127.0600 ;
        RECT 190.1200 153.7800 191.1200 154.2600 ;
        RECT 190.1200 148.3400 191.1200 148.8200 ;
        RECT 190.1200 142.9000 191.1200 143.3800 ;
        RECT 190.1200 164.6600 191.1200 165.1400 ;
        RECT 190.1200 159.2200 191.1200 159.7000 ;
        RECT 231.5600 142.9000 234.5600 143.3800 ;
        RECT 231.5600 148.3400 234.5600 148.8200 ;
        RECT 231.5600 153.7800 234.5600 154.2600 ;
        RECT 231.5600 164.6600 234.5600 165.1400 ;
        RECT 231.5600 159.2200 234.5600 159.7000 ;
        RECT 145.1200 180.9800 146.1200 181.4600 ;
        RECT 145.1200 175.5400 146.1200 176.0200 ;
        RECT 145.1200 170.1000 146.1200 170.5800 ;
        RECT 145.1200 197.3000 146.1200 197.7800 ;
        RECT 145.1200 191.8600 146.1200 192.3400 ;
        RECT 145.1200 186.4200 146.1200 186.9000 ;
        RECT 145.1200 208.1800 146.1200 208.6600 ;
        RECT 145.1200 202.7400 146.1200 203.2200 ;
        RECT 190.1200 180.9800 191.1200 181.4600 ;
        RECT 190.1200 175.5400 191.1200 176.0200 ;
        RECT 190.1200 170.1000 191.1200 170.5800 ;
        RECT 190.1200 197.3000 191.1200 197.7800 ;
        RECT 190.1200 191.8600 191.1200 192.3400 ;
        RECT 190.1200 186.4200 191.1200 186.9000 ;
        RECT 231.5600 175.5400 234.5600 176.0200 ;
        RECT 231.5600 170.1000 234.5600 170.5800 ;
        RECT 231.5600 180.9800 234.5600 181.4600 ;
        RECT 231.5600 197.3000 234.5600 197.7800 ;
        RECT 231.5600 191.8600 234.5600 192.3400 ;
        RECT 231.5600 186.4200 234.5600 186.9000 ;
        RECT 190.1200 208.1800 191.1200 208.6600 ;
        RECT 190.1200 202.7400 191.1200 203.2200 ;
        RECT 231.5600 208.1800 234.5600 208.6600 ;
        RECT 231.5600 202.7400 234.5600 203.2200 ;
      LAYER met4 ;
        RECT 5.5600 5.4300 8.5600 213.5300 ;
        RECT 231.5600 5.4300 234.5600 213.5300 ;
        RECT 55.1200 5.4300 56.1200 213.5300 ;
        RECT 100.1200 5.4300 101.1200 213.5300 ;
        RECT 145.1200 5.4300 146.1200 213.5300 ;
        RECT 190.1200 5.4300 191.1200 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5600 1.4300 238.5600 4.4300 ;
        RECT 1.5600 214.5300 238.5600 217.5300 ;
        RECT 12.3200 9.6200 13.3200 10.1000 ;
        RECT 1.5600 9.6200 4.5600 10.1000 ;
        RECT 12.3200 15.0600 13.3200 15.5400 ;
        RECT 1.5600 15.0600 4.5600 15.5400 ;
        RECT 57.3200 15.0600 58.3200 15.5400 ;
        RECT 57.3200 9.6200 58.3200 10.1000 ;
        RECT 1.5600 20.5000 4.5600 20.9800 ;
        RECT 1.5600 25.9400 4.5600 26.4200 ;
        RECT 12.3200 20.5000 13.3200 20.9800 ;
        RECT 12.3200 25.9400 13.3200 26.4200 ;
        RECT 12.3200 31.3800 13.3200 31.8600 ;
        RECT 1.5600 31.3800 4.5600 31.8600 ;
        RECT 12.3200 42.2600 13.3200 42.7400 ;
        RECT 1.5600 42.2600 4.5600 42.7400 ;
        RECT 12.3200 36.8200 13.3200 37.3000 ;
        RECT 1.5600 36.8200 4.5600 37.3000 ;
        RECT 12.3200 47.7000 13.3200 48.1800 ;
        RECT 1.5600 47.7000 4.5600 48.1800 ;
        RECT 57.3200 31.3800 58.3200 31.8600 ;
        RECT 57.3200 25.9400 58.3200 26.4200 ;
        RECT 57.3200 20.5000 58.3200 20.9800 ;
        RECT 57.3200 47.7000 58.3200 48.1800 ;
        RECT 57.3200 42.2600 58.3200 42.7400 ;
        RECT 57.3200 36.8200 58.3200 37.3000 ;
        RECT 102.3200 15.0600 103.3200 15.5400 ;
        RECT 102.3200 9.6200 103.3200 10.1000 ;
        RECT 102.3200 31.3800 103.3200 31.8600 ;
        RECT 102.3200 25.9400 103.3200 26.4200 ;
        RECT 102.3200 20.5000 103.3200 20.9800 ;
        RECT 102.3200 47.7000 103.3200 48.1800 ;
        RECT 102.3200 42.2600 103.3200 42.7400 ;
        RECT 102.3200 36.8200 103.3200 37.3000 ;
        RECT 12.3200 53.1400 13.3200 53.6200 ;
        RECT 1.5600 53.1400 4.5600 53.6200 ;
        RECT 1.5600 58.5800 4.5600 59.0600 ;
        RECT 1.5600 64.0200 4.5600 64.5000 ;
        RECT 12.3200 58.5800 13.3200 59.0600 ;
        RECT 12.3200 64.0200 13.3200 64.5000 ;
        RECT 12.3200 69.4600 13.3200 69.9400 ;
        RECT 1.5600 69.4600 4.5600 69.9400 ;
        RECT 12.3200 74.9000 13.3200 75.3800 ;
        RECT 1.5600 74.9000 4.5600 75.3800 ;
        RECT 57.3200 64.0200 58.3200 64.5000 ;
        RECT 57.3200 58.5800 58.3200 59.0600 ;
        RECT 57.3200 53.1400 58.3200 53.6200 ;
        RECT 57.3200 74.9000 58.3200 75.3800 ;
        RECT 57.3200 69.4600 58.3200 69.9400 ;
        RECT 1.5600 80.3400 4.5600 80.8200 ;
        RECT 1.5600 85.7800 4.5600 86.2600 ;
        RECT 12.3200 80.3400 13.3200 80.8200 ;
        RECT 12.3200 85.7800 13.3200 86.2600 ;
        RECT 12.3200 91.2200 13.3200 91.7000 ;
        RECT 1.5600 91.2200 4.5600 91.7000 ;
        RECT 12.3200 102.1000 13.3200 102.5800 ;
        RECT 1.5600 102.1000 4.5600 102.5800 ;
        RECT 12.3200 96.6600 13.3200 97.1400 ;
        RECT 1.5600 96.6600 4.5600 97.1400 ;
        RECT 12.3200 107.5400 13.3200 108.0200 ;
        RECT 1.5600 107.5400 4.5600 108.0200 ;
        RECT 57.3200 91.2200 58.3200 91.7000 ;
        RECT 57.3200 85.7800 58.3200 86.2600 ;
        RECT 57.3200 80.3400 58.3200 80.8200 ;
        RECT 57.3200 107.5400 58.3200 108.0200 ;
        RECT 57.3200 102.1000 58.3200 102.5800 ;
        RECT 57.3200 96.6600 58.3200 97.1400 ;
        RECT 102.3200 64.0200 103.3200 64.5000 ;
        RECT 102.3200 58.5800 103.3200 59.0600 ;
        RECT 102.3200 53.1400 103.3200 53.6200 ;
        RECT 102.3200 74.9000 103.3200 75.3800 ;
        RECT 102.3200 69.4600 103.3200 69.9400 ;
        RECT 102.3200 91.2200 103.3200 91.7000 ;
        RECT 102.3200 85.7800 103.3200 86.2600 ;
        RECT 102.3200 80.3400 103.3200 80.8200 ;
        RECT 102.3200 107.5400 103.3200 108.0200 ;
        RECT 102.3200 102.1000 103.3200 102.5800 ;
        RECT 102.3200 96.6600 103.3200 97.1400 ;
        RECT 147.3200 15.0600 148.3200 15.5400 ;
        RECT 147.3200 9.6200 148.3200 10.1000 ;
        RECT 147.3200 31.3800 148.3200 31.8600 ;
        RECT 147.3200 25.9400 148.3200 26.4200 ;
        RECT 147.3200 20.5000 148.3200 20.9800 ;
        RECT 147.3200 47.7000 148.3200 48.1800 ;
        RECT 147.3200 42.2600 148.3200 42.7400 ;
        RECT 147.3200 36.8200 148.3200 37.3000 ;
        RECT 192.3200 15.0600 193.3200 15.5400 ;
        RECT 192.3200 9.6200 193.3200 10.1000 ;
        RECT 235.5600 15.0600 238.5600 15.5400 ;
        RECT 235.5600 9.6200 238.5600 10.1000 ;
        RECT 192.3200 31.3800 193.3200 31.8600 ;
        RECT 192.3200 25.9400 193.3200 26.4200 ;
        RECT 192.3200 20.5000 193.3200 20.9800 ;
        RECT 192.3200 47.7000 193.3200 48.1800 ;
        RECT 192.3200 42.2600 193.3200 42.7400 ;
        RECT 192.3200 36.8200 193.3200 37.3000 ;
        RECT 235.5600 25.9400 238.5600 26.4200 ;
        RECT 235.5600 20.5000 238.5600 20.9800 ;
        RECT 235.5600 31.3800 238.5600 31.8600 ;
        RECT 235.5600 47.7000 238.5600 48.1800 ;
        RECT 235.5600 42.2600 238.5600 42.7400 ;
        RECT 235.5600 36.8200 238.5600 37.3000 ;
        RECT 147.3200 64.0200 148.3200 64.5000 ;
        RECT 147.3200 58.5800 148.3200 59.0600 ;
        RECT 147.3200 53.1400 148.3200 53.6200 ;
        RECT 147.3200 74.9000 148.3200 75.3800 ;
        RECT 147.3200 69.4600 148.3200 69.9400 ;
        RECT 147.3200 91.2200 148.3200 91.7000 ;
        RECT 147.3200 85.7800 148.3200 86.2600 ;
        RECT 147.3200 80.3400 148.3200 80.8200 ;
        RECT 147.3200 107.5400 148.3200 108.0200 ;
        RECT 147.3200 102.1000 148.3200 102.5800 ;
        RECT 147.3200 96.6600 148.3200 97.1400 ;
        RECT 192.3200 64.0200 193.3200 64.5000 ;
        RECT 192.3200 58.5800 193.3200 59.0600 ;
        RECT 192.3200 53.1400 193.3200 53.6200 ;
        RECT 192.3200 74.9000 193.3200 75.3800 ;
        RECT 192.3200 69.4600 193.3200 69.9400 ;
        RECT 235.5600 53.1400 238.5600 53.6200 ;
        RECT 235.5600 64.0200 238.5600 64.5000 ;
        RECT 235.5600 58.5800 238.5600 59.0600 ;
        RECT 235.5600 74.9000 238.5600 75.3800 ;
        RECT 235.5600 69.4600 238.5600 69.9400 ;
        RECT 192.3200 91.2200 193.3200 91.7000 ;
        RECT 192.3200 85.7800 193.3200 86.2600 ;
        RECT 192.3200 80.3400 193.3200 80.8200 ;
        RECT 192.3200 107.5400 193.3200 108.0200 ;
        RECT 192.3200 102.1000 193.3200 102.5800 ;
        RECT 192.3200 96.6600 193.3200 97.1400 ;
        RECT 235.5600 85.7800 238.5600 86.2600 ;
        RECT 235.5600 80.3400 238.5600 80.8200 ;
        RECT 235.5600 91.2200 238.5600 91.7000 ;
        RECT 235.5600 107.5400 238.5600 108.0200 ;
        RECT 235.5600 102.1000 238.5600 102.5800 ;
        RECT 235.5600 96.6600 238.5600 97.1400 ;
        RECT 12.3200 112.9800 13.3200 113.4600 ;
        RECT 1.5600 112.9800 4.5600 113.4600 ;
        RECT 1.5600 118.4200 4.5600 118.9000 ;
        RECT 1.5600 123.8600 4.5600 124.3400 ;
        RECT 12.3200 118.4200 13.3200 118.9000 ;
        RECT 12.3200 123.8600 13.3200 124.3400 ;
        RECT 12.3200 129.3000 13.3200 129.7800 ;
        RECT 1.5600 129.3000 4.5600 129.7800 ;
        RECT 12.3200 134.7400 13.3200 135.2200 ;
        RECT 1.5600 134.7400 4.5600 135.2200 ;
        RECT 57.3200 123.8600 58.3200 124.3400 ;
        RECT 57.3200 118.4200 58.3200 118.9000 ;
        RECT 57.3200 112.9800 58.3200 113.4600 ;
        RECT 57.3200 134.7400 58.3200 135.2200 ;
        RECT 57.3200 129.3000 58.3200 129.7800 ;
        RECT 1.5600 140.1800 4.5600 140.6600 ;
        RECT 1.5600 145.6200 4.5600 146.1000 ;
        RECT 12.3200 140.1800 13.3200 140.6600 ;
        RECT 12.3200 145.6200 13.3200 146.1000 ;
        RECT 12.3200 151.0600 13.3200 151.5400 ;
        RECT 1.5600 151.0600 4.5600 151.5400 ;
        RECT 12.3200 161.9400 13.3200 162.4200 ;
        RECT 1.5600 161.9400 4.5600 162.4200 ;
        RECT 12.3200 156.5000 13.3200 156.9800 ;
        RECT 1.5600 156.5000 4.5600 156.9800 ;
        RECT 12.3200 167.3800 13.3200 167.8600 ;
        RECT 1.5600 167.3800 4.5600 167.8600 ;
        RECT 57.3200 151.0600 58.3200 151.5400 ;
        RECT 57.3200 145.6200 58.3200 146.1000 ;
        RECT 57.3200 140.1800 58.3200 140.6600 ;
        RECT 57.3200 167.3800 58.3200 167.8600 ;
        RECT 57.3200 161.9400 58.3200 162.4200 ;
        RECT 57.3200 156.5000 58.3200 156.9800 ;
        RECT 102.3200 123.8600 103.3200 124.3400 ;
        RECT 102.3200 118.4200 103.3200 118.9000 ;
        RECT 102.3200 112.9800 103.3200 113.4600 ;
        RECT 102.3200 134.7400 103.3200 135.2200 ;
        RECT 102.3200 129.3000 103.3200 129.7800 ;
        RECT 102.3200 151.0600 103.3200 151.5400 ;
        RECT 102.3200 145.6200 103.3200 146.1000 ;
        RECT 102.3200 140.1800 103.3200 140.6600 ;
        RECT 102.3200 167.3800 103.3200 167.8600 ;
        RECT 102.3200 161.9400 103.3200 162.4200 ;
        RECT 102.3200 156.5000 103.3200 156.9800 ;
        RECT 12.3200 172.8200 13.3200 173.3000 ;
        RECT 1.5600 172.8200 4.5600 173.3000 ;
        RECT 1.5600 178.2600 4.5600 178.7400 ;
        RECT 1.5600 183.7000 4.5600 184.1800 ;
        RECT 12.3200 178.2600 13.3200 178.7400 ;
        RECT 12.3200 183.7000 13.3200 184.1800 ;
        RECT 12.3200 189.1400 13.3200 189.6200 ;
        RECT 1.5600 189.1400 4.5600 189.6200 ;
        RECT 12.3200 194.5800 13.3200 195.0600 ;
        RECT 1.5600 194.5800 4.5600 195.0600 ;
        RECT 57.3200 183.7000 58.3200 184.1800 ;
        RECT 57.3200 178.2600 58.3200 178.7400 ;
        RECT 57.3200 172.8200 58.3200 173.3000 ;
        RECT 57.3200 194.5800 58.3200 195.0600 ;
        RECT 57.3200 189.1400 58.3200 189.6200 ;
        RECT 1.5600 200.0200 4.5600 200.5000 ;
        RECT 1.5600 205.4600 4.5600 205.9400 ;
        RECT 12.3200 200.0200 13.3200 200.5000 ;
        RECT 12.3200 205.4600 13.3200 205.9400 ;
        RECT 57.3200 205.4600 58.3200 205.9400 ;
        RECT 57.3200 200.0200 58.3200 200.5000 ;
        RECT 102.3200 183.7000 103.3200 184.1800 ;
        RECT 102.3200 178.2600 103.3200 178.7400 ;
        RECT 102.3200 172.8200 103.3200 173.3000 ;
        RECT 102.3200 194.5800 103.3200 195.0600 ;
        RECT 102.3200 189.1400 103.3200 189.6200 ;
        RECT 102.3200 205.4600 103.3200 205.9400 ;
        RECT 102.3200 200.0200 103.3200 200.5000 ;
        RECT 147.3200 123.8600 148.3200 124.3400 ;
        RECT 147.3200 118.4200 148.3200 118.9000 ;
        RECT 147.3200 112.9800 148.3200 113.4600 ;
        RECT 147.3200 134.7400 148.3200 135.2200 ;
        RECT 147.3200 129.3000 148.3200 129.7800 ;
        RECT 147.3200 151.0600 148.3200 151.5400 ;
        RECT 147.3200 145.6200 148.3200 146.1000 ;
        RECT 147.3200 140.1800 148.3200 140.6600 ;
        RECT 147.3200 167.3800 148.3200 167.8600 ;
        RECT 147.3200 161.9400 148.3200 162.4200 ;
        RECT 147.3200 156.5000 148.3200 156.9800 ;
        RECT 192.3200 123.8600 193.3200 124.3400 ;
        RECT 192.3200 118.4200 193.3200 118.9000 ;
        RECT 192.3200 112.9800 193.3200 113.4600 ;
        RECT 192.3200 134.7400 193.3200 135.2200 ;
        RECT 192.3200 129.3000 193.3200 129.7800 ;
        RECT 235.5600 112.9800 238.5600 113.4600 ;
        RECT 235.5600 123.8600 238.5600 124.3400 ;
        RECT 235.5600 118.4200 238.5600 118.9000 ;
        RECT 235.5600 134.7400 238.5600 135.2200 ;
        RECT 235.5600 129.3000 238.5600 129.7800 ;
        RECT 192.3200 151.0600 193.3200 151.5400 ;
        RECT 192.3200 145.6200 193.3200 146.1000 ;
        RECT 192.3200 140.1800 193.3200 140.6600 ;
        RECT 192.3200 167.3800 193.3200 167.8600 ;
        RECT 192.3200 161.9400 193.3200 162.4200 ;
        RECT 192.3200 156.5000 193.3200 156.9800 ;
        RECT 235.5600 145.6200 238.5600 146.1000 ;
        RECT 235.5600 140.1800 238.5600 140.6600 ;
        RECT 235.5600 151.0600 238.5600 151.5400 ;
        RECT 235.5600 167.3800 238.5600 167.8600 ;
        RECT 235.5600 161.9400 238.5600 162.4200 ;
        RECT 235.5600 156.5000 238.5600 156.9800 ;
        RECT 147.3200 183.7000 148.3200 184.1800 ;
        RECT 147.3200 178.2600 148.3200 178.7400 ;
        RECT 147.3200 172.8200 148.3200 173.3000 ;
        RECT 147.3200 194.5800 148.3200 195.0600 ;
        RECT 147.3200 189.1400 148.3200 189.6200 ;
        RECT 147.3200 205.4600 148.3200 205.9400 ;
        RECT 147.3200 200.0200 148.3200 200.5000 ;
        RECT 192.3200 183.7000 193.3200 184.1800 ;
        RECT 192.3200 178.2600 193.3200 178.7400 ;
        RECT 192.3200 172.8200 193.3200 173.3000 ;
        RECT 192.3200 194.5800 193.3200 195.0600 ;
        RECT 192.3200 189.1400 193.3200 189.6200 ;
        RECT 235.5600 172.8200 238.5600 173.3000 ;
        RECT 235.5600 183.7000 238.5600 184.1800 ;
        RECT 235.5600 178.2600 238.5600 178.7400 ;
        RECT 235.5600 194.5800 238.5600 195.0600 ;
        RECT 235.5600 189.1400 238.5600 189.6200 ;
        RECT 192.3200 205.4600 193.3200 205.9400 ;
        RECT 192.3200 200.0200 193.3200 200.5000 ;
        RECT 235.5600 205.4600 238.5600 205.9400 ;
        RECT 235.5600 200.0200 238.5600 200.5000 ;
      LAYER met4 ;
        RECT 1.5600 1.4300 4.5600 217.5300 ;
        RECT 235.5600 1.4300 238.5600 217.5300 ;
        RECT 12.3200 1.4300 13.3200 217.5300 ;
        RECT 57.3200 1.4300 58.3200 217.5300 ;
        RECT 102.3200 1.4300 103.3200 217.5300 ;
        RECT 147.3200 1.4300 148.3200 217.5300 ;
        RECT 192.3200 1.4300 193.3200 217.5300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.5250 219.1400 240.1200 219.6400 ;
      RECT 148.6050 219.1400 149.0150 219.6400 ;
      RECT 147.2250 219.1400 148.0950 219.6400 ;
      RECT 145.8450 219.1400 146.7150 219.6400 ;
      RECT 144.4650 219.1400 145.3350 219.6400 ;
      RECT 143.0850 219.1400 143.9550 219.6400 ;
      RECT 141.7050 219.1400 142.5750 219.6400 ;
      RECT 140.3250 219.1400 141.1950 219.6400 ;
      RECT 138.9450 219.1400 139.8150 219.6400 ;
      RECT 137.5650 219.1400 138.4350 219.6400 ;
      RECT 136.1850 219.1400 137.0550 219.6400 ;
      RECT 134.8050 219.1400 135.6750 219.6400 ;
      RECT 133.4250 219.1400 134.2950 219.6400 ;
      RECT 132.0450 219.1400 132.9150 219.6400 ;
      RECT 130.6650 219.1400 131.5350 219.6400 ;
      RECT 129.2850 219.1400 130.1550 219.6400 ;
      RECT 127.9050 219.1400 128.7750 219.6400 ;
      RECT 126.5250 219.1400 127.3950 219.6400 ;
      RECT 125.6050 219.1400 126.0150 219.6400 ;
      RECT 124.2250 219.1400 125.0950 219.6400 ;
      RECT 122.8450 219.1400 123.7150 219.6400 ;
      RECT 121.4650 219.1400 122.3350 219.6400 ;
      RECT 120.0850 219.1400 120.9550 219.6400 ;
      RECT 118.7050 219.1400 119.5750 219.6400 ;
      RECT 117.3250 219.1400 118.1950 219.6400 ;
      RECT 115.9450 219.1400 116.8150 219.6400 ;
      RECT 114.5650 219.1400 115.4350 219.6400 ;
      RECT 113.1850 219.1400 114.0550 219.6400 ;
      RECT 111.8050 219.1400 112.6750 219.6400 ;
      RECT 110.4250 219.1400 111.2950 219.6400 ;
      RECT 109.0450 219.1400 109.9150 219.6400 ;
      RECT 107.6650 219.1400 108.5350 219.6400 ;
      RECT 106.2850 219.1400 107.1550 219.6400 ;
      RECT 104.9050 219.1400 105.7750 219.6400 ;
      RECT 103.5250 219.1400 104.3950 219.6400 ;
      RECT 102.6050 219.1400 103.0150 219.6400 ;
      RECT 101.2250 219.1400 102.0950 219.6400 ;
      RECT 99.8450 219.1400 100.7150 219.6400 ;
      RECT 98.4650 219.1400 99.3350 219.6400 ;
      RECT 97.0850 219.1400 97.9550 219.6400 ;
      RECT 95.7050 219.1400 96.5750 219.6400 ;
      RECT 94.3250 219.1400 95.1950 219.6400 ;
      RECT 92.9450 219.1400 93.8150 219.6400 ;
      RECT 91.5650 219.1400 92.4350 219.6400 ;
      RECT 90.1850 219.1400 91.0550 219.6400 ;
      RECT 88.8050 219.1400 89.6750 219.6400 ;
      RECT 87.4250 219.1400 88.2950 219.6400 ;
      RECT 86.0450 219.1400 86.9150 219.6400 ;
      RECT 84.6650 219.1400 85.5350 219.6400 ;
      RECT 83.2850 219.1400 84.1550 219.6400 ;
      RECT 81.9050 219.1400 82.7750 219.6400 ;
      RECT 80.5250 219.1400 81.3950 219.6400 ;
      RECT 79.6050 219.1400 80.0150 219.6400 ;
      RECT 78.2250 219.1400 79.0950 219.6400 ;
      RECT 76.8450 219.1400 77.7150 219.6400 ;
      RECT 75.4650 219.1400 76.3350 219.6400 ;
      RECT 74.0850 219.1400 74.9550 219.6400 ;
      RECT 72.7050 219.1400 73.5750 219.6400 ;
      RECT 71.3250 219.1400 72.1950 219.6400 ;
      RECT 69.9450 219.1400 70.8150 219.6400 ;
      RECT 68.5650 219.1400 69.4350 219.6400 ;
      RECT 67.1850 219.1400 68.0550 219.6400 ;
      RECT 65.8050 219.1400 66.6750 219.6400 ;
      RECT 64.4250 219.1400 65.2950 219.6400 ;
      RECT 63.0450 219.1400 63.9150 219.6400 ;
      RECT 61.6650 219.1400 62.5350 219.6400 ;
      RECT 60.2850 219.1400 61.1550 219.6400 ;
      RECT 58.9050 219.1400 59.7750 219.6400 ;
      RECT 57.5250 219.1400 58.3950 219.6400 ;
      RECT 56.6050 219.1400 57.0150 219.6400 ;
      RECT 55.2250 219.1400 56.0950 219.6400 ;
      RECT 53.8450 219.1400 54.7150 219.6400 ;
      RECT 52.4650 219.1400 53.3350 219.6400 ;
      RECT 51.0850 219.1400 51.9550 219.6400 ;
      RECT 49.7050 219.1400 50.5750 219.6400 ;
      RECT 48.3250 219.1400 49.1950 219.6400 ;
      RECT 46.9450 219.1400 47.8150 219.6400 ;
      RECT 45.5650 219.1400 46.4350 219.6400 ;
      RECT 44.1850 219.1400 45.0550 219.6400 ;
      RECT 42.8050 219.1400 43.6750 219.6400 ;
      RECT 41.4250 219.1400 42.2950 219.6400 ;
      RECT 40.0450 219.1400 40.9150 219.6400 ;
      RECT 38.6650 219.1400 39.5350 219.6400 ;
      RECT 37.2850 219.1400 38.1550 219.6400 ;
      RECT 35.9050 219.1400 36.7750 219.6400 ;
      RECT 34.5250 219.1400 35.3950 219.6400 ;
      RECT 33.6050 219.1400 34.0150 219.6400 ;
      RECT 32.2250 219.1400 33.0950 219.6400 ;
      RECT 30.8450 219.1400 31.7150 219.6400 ;
      RECT 29.4650 219.1400 30.3350 219.6400 ;
      RECT 28.0850 219.1400 28.9550 219.6400 ;
      RECT 26.7050 219.1400 27.5750 219.6400 ;
      RECT 25.3250 219.1400 26.1950 219.6400 ;
      RECT 23.9450 219.1400 24.8150 219.6400 ;
      RECT 22.5650 219.1400 23.4350 219.6400 ;
      RECT 21.1850 219.1400 22.0550 219.6400 ;
      RECT 19.8050 219.1400 20.6750 219.6400 ;
      RECT 18.4250 219.1400 19.2950 219.6400 ;
      RECT 17.0450 219.1400 17.9150 219.6400 ;
      RECT 15.6650 219.1400 16.5350 219.6400 ;
      RECT 14.2850 219.1400 15.1550 219.6400 ;
      RECT 12.9050 219.1400 13.7750 219.6400 ;
      RECT 11.5250 219.1400 12.3950 219.6400 ;
      RECT 10.6050 219.1400 11.0150 219.6400 ;
      RECT 0.0000 219.1400 10.0950 219.6400 ;
      RECT 0.0000 0.5000 240.1200 219.1400 ;
      RECT 149.5250 0.0000 240.1200 0.5000 ;
      RECT 148.6050 0.0000 149.0150 0.5000 ;
      RECT 147.2250 0.0000 148.0950 0.5000 ;
      RECT 145.8450 0.0000 146.7150 0.5000 ;
      RECT 144.4650 0.0000 145.3350 0.5000 ;
      RECT 143.0850 0.0000 143.9550 0.5000 ;
      RECT 141.7050 0.0000 142.5750 0.5000 ;
      RECT 140.3250 0.0000 141.1950 0.5000 ;
      RECT 138.9450 0.0000 139.8150 0.5000 ;
      RECT 137.5650 0.0000 138.4350 0.5000 ;
      RECT 136.1850 0.0000 137.0550 0.5000 ;
      RECT 134.8050 0.0000 135.6750 0.5000 ;
      RECT 133.4250 0.0000 134.2950 0.5000 ;
      RECT 132.0450 0.0000 132.9150 0.5000 ;
      RECT 130.6650 0.0000 131.5350 0.5000 ;
      RECT 129.2850 0.0000 130.1550 0.5000 ;
      RECT 127.9050 0.0000 128.7750 0.5000 ;
      RECT 126.5250 0.0000 127.3950 0.5000 ;
      RECT 125.6050 0.0000 126.0150 0.5000 ;
      RECT 124.2250 0.0000 125.0950 0.5000 ;
      RECT 122.8450 0.0000 123.7150 0.5000 ;
      RECT 121.4650 0.0000 122.3350 0.5000 ;
      RECT 120.0850 0.0000 120.9550 0.5000 ;
      RECT 118.7050 0.0000 119.5750 0.5000 ;
      RECT 117.3250 0.0000 118.1950 0.5000 ;
      RECT 115.9450 0.0000 116.8150 0.5000 ;
      RECT 114.5650 0.0000 115.4350 0.5000 ;
      RECT 113.1850 0.0000 114.0550 0.5000 ;
      RECT 111.8050 0.0000 112.6750 0.5000 ;
      RECT 110.4250 0.0000 111.2950 0.5000 ;
      RECT 109.0450 0.0000 109.9150 0.5000 ;
      RECT 107.6650 0.0000 108.5350 0.5000 ;
      RECT 106.2850 0.0000 107.1550 0.5000 ;
      RECT 104.9050 0.0000 105.7750 0.5000 ;
      RECT 103.5250 0.0000 104.3950 0.5000 ;
      RECT 102.6050 0.0000 103.0150 0.5000 ;
      RECT 101.2250 0.0000 102.0950 0.5000 ;
      RECT 99.8450 0.0000 100.7150 0.5000 ;
      RECT 98.4650 0.0000 99.3350 0.5000 ;
      RECT 97.0850 0.0000 97.9550 0.5000 ;
      RECT 95.7050 0.0000 96.5750 0.5000 ;
      RECT 94.3250 0.0000 95.1950 0.5000 ;
      RECT 92.9450 0.0000 93.8150 0.5000 ;
      RECT 91.5650 0.0000 92.4350 0.5000 ;
      RECT 90.1850 0.0000 91.0550 0.5000 ;
      RECT 88.8050 0.0000 89.6750 0.5000 ;
      RECT 87.4250 0.0000 88.2950 0.5000 ;
      RECT 86.0450 0.0000 86.9150 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.6050 0.0000 80.0150 0.5000 ;
      RECT 78.2250 0.0000 79.0950 0.5000 ;
      RECT 76.8450 0.0000 77.7150 0.5000 ;
      RECT 75.4650 0.0000 76.3350 0.5000 ;
      RECT 74.0850 0.0000 74.9550 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 61.6650 0.0000 62.5350 0.5000 ;
      RECT 60.2850 0.0000 61.1550 0.5000 ;
      RECT 58.9050 0.0000 59.7750 0.5000 ;
      RECT 57.5250 0.0000 58.3950 0.5000 ;
      RECT 56.6050 0.0000 57.0150 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 49.7050 0.0000 50.5750 0.5000 ;
      RECT 48.3250 0.0000 49.1950 0.5000 ;
      RECT 46.9450 0.0000 47.8150 0.5000 ;
      RECT 45.5650 0.0000 46.4350 0.5000 ;
      RECT 44.1850 0.0000 45.0550 0.5000 ;
      RECT 42.8050 0.0000 43.6750 0.5000 ;
      RECT 41.4250 0.0000 42.2950 0.5000 ;
      RECT 40.0450 0.0000 40.9150 0.5000 ;
      RECT 38.6650 0.0000 39.5350 0.5000 ;
      RECT 37.2850 0.0000 38.1550 0.5000 ;
      RECT 35.9050 0.0000 36.7750 0.5000 ;
      RECT 34.5250 0.0000 35.3950 0.5000 ;
      RECT 33.6050 0.0000 34.0150 0.5000 ;
      RECT 32.2250 0.0000 33.0950 0.5000 ;
      RECT 30.8450 0.0000 31.7150 0.5000 ;
      RECT 29.4650 0.0000 30.3350 0.5000 ;
      RECT 28.0850 0.0000 28.9550 0.5000 ;
      RECT 26.7050 0.0000 27.5750 0.5000 ;
      RECT 25.3250 0.0000 26.1950 0.5000 ;
      RECT 23.9450 0.0000 24.8150 0.5000 ;
      RECT 22.5650 0.0000 23.4350 0.5000 ;
      RECT 21.1850 0.0000 22.0550 0.5000 ;
      RECT 19.8050 0.0000 20.6750 0.5000 ;
      RECT 18.4250 0.0000 19.2950 0.5000 ;
      RECT 17.0450 0.0000 17.9150 0.5000 ;
      RECT 15.6650 0.0000 16.5350 0.5000 ;
      RECT 14.2850 0.0000 15.1550 0.5000 ;
      RECT 12.9050 0.0000 13.7750 0.5000 ;
      RECT 11.5250 0.0000 12.3950 0.5000 ;
      RECT 10.6050 0.0000 11.0150 0.5000 ;
      RECT 0.0000 0.0000 10.0950 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 240.1200 219.6400 ;
    LAYER met2 ;
      RECT 210.2000 219.0150 240.1200 219.6400 ;
      RECT 206.9800 219.0150 209.7800 219.6400 ;
      RECT 204.2200 219.0150 206.5600 219.6400 ;
      RECT 201.4600 219.0150 203.8000 219.6400 ;
      RECT 198.2400 219.0150 201.0400 219.6400 ;
      RECT 195.4800 219.0150 197.8200 219.6400 ;
      RECT 192.7200 219.0150 195.0600 219.6400 ;
      RECT 189.9600 219.0150 192.3000 219.6400 ;
      RECT 186.7400 219.0150 189.5400 219.6400 ;
      RECT 183.9800 219.0150 186.3200 219.6400 ;
      RECT 181.2200 219.0150 183.5600 219.6400 ;
      RECT 178.4600 219.0150 180.8000 219.6400 ;
      RECT 175.2400 219.0150 178.0400 219.6400 ;
      RECT 172.4800 219.0150 174.8200 219.6400 ;
      RECT 169.2600 219.0150 172.0600 219.6400 ;
      RECT 166.9600 219.0150 168.8400 219.6400 ;
      RECT 163.7400 219.0150 166.5400 219.6400 ;
      RECT 160.9800 219.0150 163.3200 219.6400 ;
      RECT 157.7600 219.0150 160.5600 219.6400 ;
      RECT 155.4600 219.0150 157.3400 219.6400 ;
      RECT 0.0000 219.0150 155.0400 219.6400 ;
      RECT 0.0000 209.8200 240.1200 219.0150 ;
      RECT 0.6250 209.4000 239.4950 209.8200 ;
      RECT 0.0000 208.1200 240.1200 209.4000 ;
      RECT 0.6250 207.7000 239.4950 208.1200 ;
      RECT 0.0000 206.4200 240.1200 207.7000 ;
      RECT 0.6250 206.0000 239.4950 206.4200 ;
      RECT 0.0000 204.7200 240.1200 206.0000 ;
      RECT 0.6250 204.3000 239.4950 204.7200 ;
      RECT 0.0000 203.0200 240.1200 204.3000 ;
      RECT 0.6250 202.6000 239.4950 203.0200 ;
      RECT 0.0000 201.3200 240.1200 202.6000 ;
      RECT 0.6250 200.9000 239.4950 201.3200 ;
      RECT 0.0000 199.2800 240.1200 200.9000 ;
      RECT 0.6250 198.8600 239.4950 199.2800 ;
      RECT 0.0000 197.5800 240.1200 198.8600 ;
      RECT 0.6250 197.1600 239.4950 197.5800 ;
      RECT 0.0000 195.8800 240.1200 197.1600 ;
      RECT 0.6250 195.4600 239.4950 195.8800 ;
      RECT 0.0000 194.1800 240.1200 195.4600 ;
      RECT 0.6250 193.7600 239.4950 194.1800 ;
      RECT 0.0000 192.4800 240.1200 193.7600 ;
      RECT 0.6250 192.0600 239.4950 192.4800 ;
      RECT 0.0000 190.4400 240.1200 192.0600 ;
      RECT 0.6250 190.0200 239.4950 190.4400 ;
      RECT 0.0000 188.7400 240.1200 190.0200 ;
      RECT 0.6250 188.3200 239.4950 188.7400 ;
      RECT 0.0000 187.0400 240.1200 188.3200 ;
      RECT 0.6250 186.6200 239.4950 187.0400 ;
      RECT 0.0000 185.3400 240.1200 186.6200 ;
      RECT 0.6250 184.9200 239.4950 185.3400 ;
      RECT 0.0000 183.6400 240.1200 184.9200 ;
      RECT 0.6250 183.2200 239.4950 183.6400 ;
      RECT 0.0000 181.6000 240.1200 183.2200 ;
      RECT 0.6250 181.1800 239.4950 181.6000 ;
      RECT 0.0000 179.9000 240.1200 181.1800 ;
      RECT 0.6250 179.4800 239.4950 179.9000 ;
      RECT 0.0000 178.2000 240.1200 179.4800 ;
      RECT 0.6250 177.7800 239.4950 178.2000 ;
      RECT 0.0000 176.5000 240.1200 177.7800 ;
      RECT 0.6250 176.0800 239.4950 176.5000 ;
      RECT 0.0000 174.8000 240.1200 176.0800 ;
      RECT 0.6250 174.3800 239.4950 174.8000 ;
      RECT 0.0000 172.7600 240.1200 174.3800 ;
      RECT 0.6250 172.3400 239.4950 172.7600 ;
      RECT 0.0000 171.0600 240.1200 172.3400 ;
      RECT 0.6250 170.6400 239.4950 171.0600 ;
      RECT 0.0000 169.3600 240.1200 170.6400 ;
      RECT 0.6250 168.9400 239.4950 169.3600 ;
      RECT 0.0000 167.6600 240.1200 168.9400 ;
      RECT 0.6250 167.2400 239.4950 167.6600 ;
      RECT 0.0000 165.9600 240.1200 167.2400 ;
      RECT 0.6250 165.5400 239.4950 165.9600 ;
      RECT 0.0000 163.9200 240.1200 165.5400 ;
      RECT 0.6250 163.5000 239.4950 163.9200 ;
      RECT 0.0000 162.2200 240.1200 163.5000 ;
      RECT 0.6250 161.8000 239.4950 162.2200 ;
      RECT 0.0000 160.5200 240.1200 161.8000 ;
      RECT 0.6250 160.1000 239.4950 160.5200 ;
      RECT 0.0000 158.8200 240.1200 160.1000 ;
      RECT 0.6250 158.4000 239.4950 158.8200 ;
      RECT 0.0000 157.1200 240.1200 158.4000 ;
      RECT 0.6250 156.7000 239.4950 157.1200 ;
      RECT 0.0000 155.4200 240.1200 156.7000 ;
      RECT 0.6250 155.0000 239.4950 155.4200 ;
      RECT 0.0000 149.9800 240.1200 155.0000 ;
      RECT 0.6250 149.5600 239.4950 149.9800 ;
      RECT 0.0000 148.2800 240.1200 149.5600 ;
      RECT 0.6250 147.8600 239.4950 148.2800 ;
      RECT 0.0000 146.9200 240.1200 147.8600 ;
      RECT 0.6250 146.5000 239.4950 146.9200 ;
      RECT 0.0000 145.5600 240.1200 146.5000 ;
      RECT 0.6250 145.1400 239.4950 145.5600 ;
      RECT 0.0000 143.8600 240.1200 145.1400 ;
      RECT 0.6250 143.4400 239.4950 143.8600 ;
      RECT 0.0000 142.5000 240.1200 143.4400 ;
      RECT 0.6250 142.0800 239.4950 142.5000 ;
      RECT 0.0000 141.1400 240.1200 142.0800 ;
      RECT 0.6250 140.7200 239.4950 141.1400 ;
      RECT 0.0000 139.4400 240.1200 140.7200 ;
      RECT 0.6250 139.0200 239.4950 139.4400 ;
      RECT 0.0000 138.0800 240.1200 139.0200 ;
      RECT 0.6250 137.6600 239.4950 138.0800 ;
      RECT 0.0000 136.7200 240.1200 137.6600 ;
      RECT 0.6250 136.3000 239.4950 136.7200 ;
      RECT 0.0000 135.0200 240.1200 136.3000 ;
      RECT 0.6250 134.6000 239.4950 135.0200 ;
      RECT 0.0000 133.6600 240.1200 134.6000 ;
      RECT 0.6250 133.2400 239.4950 133.6600 ;
      RECT 0.0000 132.3000 240.1200 133.2400 ;
      RECT 0.6250 131.8800 239.4950 132.3000 ;
      RECT 0.0000 130.6000 240.1200 131.8800 ;
      RECT 0.6250 130.1800 239.4950 130.6000 ;
      RECT 0.0000 129.2400 240.1200 130.1800 ;
      RECT 0.6250 128.8200 239.4950 129.2400 ;
      RECT 0.0000 127.8800 240.1200 128.8200 ;
      RECT 0.6250 127.4600 239.4950 127.8800 ;
      RECT 0.0000 126.1800 240.1200 127.4600 ;
      RECT 0.6250 125.7600 239.4950 126.1800 ;
      RECT 0.0000 124.8200 240.1200 125.7600 ;
      RECT 0.6250 124.4000 239.4950 124.8200 ;
      RECT 0.0000 123.4600 240.1200 124.4000 ;
      RECT 0.6250 123.0400 239.4950 123.4600 ;
      RECT 0.0000 121.7600 240.1200 123.0400 ;
      RECT 0.6250 121.3400 239.4950 121.7600 ;
      RECT 0.0000 120.4000 240.1200 121.3400 ;
      RECT 0.6250 119.9800 239.4950 120.4000 ;
      RECT 0.0000 119.0400 240.1200 119.9800 ;
      RECT 0.6250 118.6200 239.4950 119.0400 ;
      RECT 0.0000 117.3400 240.1200 118.6200 ;
      RECT 0.6250 116.9200 239.4950 117.3400 ;
      RECT 0.0000 115.9800 240.1200 116.9200 ;
      RECT 0.6250 115.5600 239.4950 115.9800 ;
      RECT 0.0000 114.6200 240.1200 115.5600 ;
      RECT 0.6250 114.2000 239.4950 114.6200 ;
      RECT 0.0000 112.9200 240.1200 114.2000 ;
      RECT 0.6250 112.5000 239.4950 112.9200 ;
      RECT 0.0000 111.5600 240.1200 112.5000 ;
      RECT 0.6250 111.1400 239.4950 111.5600 ;
      RECT 0.0000 110.2000 240.1200 111.1400 ;
      RECT 0.6250 109.7800 239.4950 110.2000 ;
      RECT 0.0000 108.5000 240.1200 109.7800 ;
      RECT 0.6250 108.0800 239.4950 108.5000 ;
      RECT 0.0000 107.1400 240.1200 108.0800 ;
      RECT 0.6250 106.7200 239.4950 107.1400 ;
      RECT 0.0000 105.7800 240.1200 106.7200 ;
      RECT 0.6250 105.3600 239.4950 105.7800 ;
      RECT 0.0000 104.0800 240.1200 105.3600 ;
      RECT 0.6250 103.6600 239.4950 104.0800 ;
      RECT 0.0000 102.7200 240.1200 103.6600 ;
      RECT 0.6250 102.3000 239.4950 102.7200 ;
      RECT 0.0000 101.3600 240.1200 102.3000 ;
      RECT 0.6250 100.9400 239.4950 101.3600 ;
      RECT 0.0000 99.6600 240.1200 100.9400 ;
      RECT 0.6250 99.2400 239.4950 99.6600 ;
      RECT 0.0000 98.3000 240.1200 99.2400 ;
      RECT 0.6250 97.8800 239.4950 98.3000 ;
      RECT 0.0000 96.9400 240.1200 97.8800 ;
      RECT 0.6250 96.5200 239.4950 96.9400 ;
      RECT 0.0000 95.2400 240.1200 96.5200 ;
      RECT 0.6250 94.8200 239.4950 95.2400 ;
      RECT 0.0000 93.8800 240.1200 94.8200 ;
      RECT 0.6250 93.4600 239.4950 93.8800 ;
      RECT 0.0000 92.5200 240.1200 93.4600 ;
      RECT 0.6250 92.1000 239.4950 92.5200 ;
      RECT 0.0000 90.8200 240.1200 92.1000 ;
      RECT 0.6250 90.4000 239.4950 90.8200 ;
      RECT 0.0000 89.4600 240.1200 90.4000 ;
      RECT 0.6250 89.0400 239.4950 89.4600 ;
      RECT 0.0000 88.1000 240.1200 89.0400 ;
      RECT 0.6250 87.6800 239.4950 88.1000 ;
      RECT 0.0000 86.4000 240.1200 87.6800 ;
      RECT 0.6250 85.9800 239.4950 86.4000 ;
      RECT 0.0000 85.0400 240.1200 85.9800 ;
      RECT 0.6250 84.6200 239.4950 85.0400 ;
      RECT 0.0000 83.6800 240.1200 84.6200 ;
      RECT 0.6250 83.2600 239.4950 83.6800 ;
      RECT 0.0000 81.9800 240.1200 83.2600 ;
      RECT 0.6250 81.5600 239.4950 81.9800 ;
      RECT 0.0000 80.6200 240.1200 81.5600 ;
      RECT 0.6250 80.2000 239.4950 80.6200 ;
      RECT 0.0000 79.2600 240.1200 80.2000 ;
      RECT 0.6250 78.8400 239.4950 79.2600 ;
      RECT 0.0000 77.9000 240.1200 78.8400 ;
      RECT 0.6250 77.4800 239.4950 77.9000 ;
      RECT 0.0000 76.2000 240.1200 77.4800 ;
      RECT 0.6250 75.7800 239.4950 76.2000 ;
      RECT 0.0000 74.8400 240.1200 75.7800 ;
      RECT 0.6250 74.4200 239.4950 74.8400 ;
      RECT 0.0000 73.4800 240.1200 74.4200 ;
      RECT 0.6250 73.0600 239.4950 73.4800 ;
      RECT 0.0000 71.7800 240.1200 73.0600 ;
      RECT 0.6250 71.3600 239.4950 71.7800 ;
      RECT 0.0000 70.4200 240.1200 71.3600 ;
      RECT 0.6250 70.0000 239.4950 70.4200 ;
      RECT 0.0000 69.0600 240.1200 70.0000 ;
      RECT 0.6250 68.6400 239.4950 69.0600 ;
      RECT 0.0000 67.3600 240.1200 68.6400 ;
      RECT 0.6250 66.9400 239.4950 67.3600 ;
      RECT 0.0000 66.0000 240.1200 66.9400 ;
      RECT 0.6250 65.5800 239.4950 66.0000 ;
      RECT 0.0000 64.6400 240.1200 65.5800 ;
      RECT 0.6250 64.2200 239.4950 64.6400 ;
      RECT 0.0000 62.9400 240.1200 64.2200 ;
      RECT 0.6250 62.5200 239.4950 62.9400 ;
      RECT 0.0000 61.5800 240.1200 62.5200 ;
      RECT 0.6250 61.1600 239.4950 61.5800 ;
      RECT 0.0000 60.2200 240.1200 61.1600 ;
      RECT 0.6250 59.8000 239.4950 60.2200 ;
      RECT 0.0000 58.5200 240.1200 59.8000 ;
      RECT 0.6250 58.1000 239.4950 58.5200 ;
      RECT 0.0000 57.1600 240.1200 58.1000 ;
      RECT 0.6250 56.7400 239.4950 57.1600 ;
      RECT 0.0000 55.8000 240.1200 56.7400 ;
      RECT 0.6250 55.3800 239.4950 55.8000 ;
      RECT 0.0000 54.1000 240.1200 55.3800 ;
      RECT 0.6250 53.6800 239.4950 54.1000 ;
      RECT 0.0000 52.7400 240.1200 53.6800 ;
      RECT 0.6250 52.3200 239.4950 52.7400 ;
      RECT 0.0000 51.3800 240.1200 52.3200 ;
      RECT 0.6250 50.9600 239.4950 51.3800 ;
      RECT 0.0000 49.6800 240.1200 50.9600 ;
      RECT 0.6250 49.2600 239.4950 49.6800 ;
      RECT 0.0000 48.3200 240.1200 49.2600 ;
      RECT 0.6250 47.9000 239.4950 48.3200 ;
      RECT 0.0000 46.9600 240.1200 47.9000 ;
      RECT 0.6250 46.5400 239.4950 46.9600 ;
      RECT 0.0000 45.2600 240.1200 46.5400 ;
      RECT 0.6250 44.8400 239.4950 45.2600 ;
      RECT 0.0000 43.9000 240.1200 44.8400 ;
      RECT 0.6250 43.4800 239.4950 43.9000 ;
      RECT 0.0000 42.5400 240.1200 43.4800 ;
      RECT 0.6250 42.1200 239.4950 42.5400 ;
      RECT 0.0000 40.8400 240.1200 42.1200 ;
      RECT 0.6250 40.4200 239.4950 40.8400 ;
      RECT 0.0000 39.4800 240.1200 40.4200 ;
      RECT 0.6250 39.0600 239.4950 39.4800 ;
      RECT 0.0000 38.1200 240.1200 39.0600 ;
      RECT 0.6250 37.7000 239.4950 38.1200 ;
      RECT 0.0000 36.4200 240.1200 37.7000 ;
      RECT 0.6250 36.0000 239.4950 36.4200 ;
      RECT 0.0000 35.0600 240.1200 36.0000 ;
      RECT 0.6250 34.6400 239.4950 35.0600 ;
      RECT 0.0000 33.7000 240.1200 34.6400 ;
      RECT 0.6250 33.2800 239.4950 33.7000 ;
      RECT 0.0000 32.0000 240.1200 33.2800 ;
      RECT 0.6250 31.5800 239.4950 32.0000 ;
      RECT 0.0000 30.6400 240.1200 31.5800 ;
      RECT 0.6250 30.2200 239.4950 30.6400 ;
      RECT 0.0000 29.2800 240.1200 30.2200 ;
      RECT 0.6250 28.8600 239.4950 29.2800 ;
      RECT 0.0000 27.5800 240.1200 28.8600 ;
      RECT 0.6250 27.1600 239.4950 27.5800 ;
      RECT 0.0000 26.2200 240.1200 27.1600 ;
      RECT 0.6250 25.8000 239.4950 26.2200 ;
      RECT 0.0000 24.8600 240.1200 25.8000 ;
      RECT 0.6250 24.4400 239.4950 24.8600 ;
      RECT 0.0000 23.1600 240.1200 24.4400 ;
      RECT 0.6250 22.7400 239.4950 23.1600 ;
      RECT 0.0000 21.8000 240.1200 22.7400 ;
      RECT 0.6250 21.3800 239.4950 21.8000 ;
      RECT 0.0000 20.4400 240.1200 21.3800 ;
      RECT 0.6250 20.0200 239.4950 20.4400 ;
      RECT 0.0000 18.7400 240.1200 20.0200 ;
      RECT 0.6250 18.3200 239.4950 18.7400 ;
      RECT 0.0000 17.3800 240.1200 18.3200 ;
      RECT 0.6250 16.9600 239.4950 17.3800 ;
      RECT 0.0000 16.0200 240.1200 16.9600 ;
      RECT 0.6250 15.6000 239.4950 16.0200 ;
      RECT 0.0000 14.3200 240.1200 15.6000 ;
      RECT 0.6250 13.9000 239.4950 14.3200 ;
      RECT 0.0000 12.9600 240.1200 13.9000 ;
      RECT 0.6250 12.5400 239.4950 12.9600 ;
      RECT 0.0000 11.6000 240.1200 12.5400 ;
      RECT 0.6250 11.1800 239.4950 11.6000 ;
      RECT 0.0000 10.2400 240.1200 11.1800 ;
      RECT 0.6250 9.8200 239.4950 10.2400 ;
      RECT 0.0000 0.6250 240.1200 9.8200 ;
      RECT 210.2000 0.0000 240.1200 0.6250 ;
      RECT 206.9800 0.0000 209.7800 0.6250 ;
      RECT 204.2200 0.0000 206.5600 0.6250 ;
      RECT 201.4600 0.0000 203.8000 0.6250 ;
      RECT 197.7800 0.0000 201.0400 0.6250 ;
      RECT 195.4800 0.0000 197.3600 0.6250 ;
      RECT 192.7200 0.0000 195.0600 0.6250 ;
      RECT 189.9600 0.0000 192.3000 0.6250 ;
      RECT 186.7400 0.0000 189.5400 0.6250 ;
      RECT 183.9800 0.0000 186.3200 0.6250 ;
      RECT 181.2200 0.0000 183.5600 0.6250 ;
      RECT 178.4600 0.0000 180.8000 0.6250 ;
      RECT 175.2400 0.0000 178.0400 0.6250 ;
      RECT 172.4800 0.0000 174.8200 0.6250 ;
      RECT 169.7200 0.0000 172.0600 0.6250 ;
      RECT 166.5000 0.0000 169.3000 0.6250 ;
      RECT 163.7400 0.0000 166.0800 0.6250 ;
      RECT 160.9800 0.0000 163.3200 0.6250 ;
      RECT 158.2200 0.0000 160.5600 0.6250 ;
      RECT 155.4600 0.0000 157.8000 0.6250 ;
      RECT 0.0000 0.0000 155.0400 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 217.8300 240.1200 219.6400 ;
      RECT 238.8600 214.2300 240.1200 217.8300 ;
      RECT 0.0000 214.2300 1.2600 217.8300 ;
      RECT 0.0000 213.8300 240.1200 214.2300 ;
      RECT 234.8600 210.2300 240.1200 213.8300 ;
      RECT 0.0000 210.2300 5.2600 213.8300 ;
      RECT 0.0000 208.9600 240.1200 210.2300 ;
      RECT 234.8600 207.8800 240.1200 208.9600 ;
      RECT 191.4200 207.8800 231.2600 208.9600 ;
      RECT 146.4200 207.8800 189.8200 208.9600 ;
      RECT 101.4200 207.8800 144.8200 208.9600 ;
      RECT 56.4200 207.8800 99.8200 208.9600 ;
      RECT 8.8600 207.8800 54.8200 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 240.1200 207.8800 ;
      RECT 238.8600 205.1600 240.1200 206.2400 ;
      RECT 193.6200 205.1600 235.2600 206.2400 ;
      RECT 148.6200 205.1600 192.0200 206.2400 ;
      RECT 103.6200 205.1600 147.0200 206.2400 ;
      RECT 58.6200 205.1600 102.0200 206.2400 ;
      RECT 13.6200 205.1600 57.0200 206.2400 ;
      RECT 4.8600 205.1600 12.0200 206.2400 ;
      RECT 0.0000 205.1600 1.2600 206.2400 ;
      RECT 0.0000 203.5200 240.1200 205.1600 ;
      RECT 234.8600 202.4400 240.1200 203.5200 ;
      RECT 191.4200 202.4400 231.2600 203.5200 ;
      RECT 146.4200 202.4400 189.8200 203.5200 ;
      RECT 101.4200 202.4400 144.8200 203.5200 ;
      RECT 56.4200 202.4400 99.8200 203.5200 ;
      RECT 8.8600 202.4400 54.8200 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 240.1200 202.4400 ;
      RECT 238.8600 199.7200 240.1200 200.8000 ;
      RECT 193.6200 199.7200 235.2600 200.8000 ;
      RECT 148.6200 199.7200 192.0200 200.8000 ;
      RECT 103.6200 199.7200 147.0200 200.8000 ;
      RECT 58.6200 199.7200 102.0200 200.8000 ;
      RECT 13.6200 199.7200 57.0200 200.8000 ;
      RECT 4.8600 199.7200 12.0200 200.8000 ;
      RECT 0.0000 199.7200 1.2600 200.8000 ;
      RECT 0.0000 198.0800 240.1200 199.7200 ;
      RECT 234.8600 197.0000 240.1200 198.0800 ;
      RECT 191.4200 197.0000 231.2600 198.0800 ;
      RECT 146.4200 197.0000 189.8200 198.0800 ;
      RECT 101.4200 197.0000 144.8200 198.0800 ;
      RECT 56.4200 197.0000 99.8200 198.0800 ;
      RECT 8.8600 197.0000 54.8200 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 240.1200 197.0000 ;
      RECT 238.8600 194.2800 240.1200 195.3600 ;
      RECT 193.6200 194.2800 235.2600 195.3600 ;
      RECT 148.6200 194.2800 192.0200 195.3600 ;
      RECT 103.6200 194.2800 147.0200 195.3600 ;
      RECT 58.6200 194.2800 102.0200 195.3600 ;
      RECT 13.6200 194.2800 57.0200 195.3600 ;
      RECT 4.8600 194.2800 12.0200 195.3600 ;
      RECT 0.0000 194.2800 1.2600 195.3600 ;
      RECT 0.0000 192.6400 240.1200 194.2800 ;
      RECT 234.8600 191.5600 240.1200 192.6400 ;
      RECT 191.4200 191.5600 231.2600 192.6400 ;
      RECT 146.4200 191.5600 189.8200 192.6400 ;
      RECT 101.4200 191.5600 144.8200 192.6400 ;
      RECT 56.4200 191.5600 99.8200 192.6400 ;
      RECT 8.8600 191.5600 54.8200 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 240.1200 191.5600 ;
      RECT 238.8600 188.8400 240.1200 189.9200 ;
      RECT 193.6200 188.8400 235.2600 189.9200 ;
      RECT 148.6200 188.8400 192.0200 189.9200 ;
      RECT 103.6200 188.8400 147.0200 189.9200 ;
      RECT 58.6200 188.8400 102.0200 189.9200 ;
      RECT 13.6200 188.8400 57.0200 189.9200 ;
      RECT 4.8600 188.8400 12.0200 189.9200 ;
      RECT 0.0000 188.8400 1.2600 189.9200 ;
      RECT 0.0000 187.2000 240.1200 188.8400 ;
      RECT 234.8600 186.1200 240.1200 187.2000 ;
      RECT 191.4200 186.1200 231.2600 187.2000 ;
      RECT 146.4200 186.1200 189.8200 187.2000 ;
      RECT 101.4200 186.1200 144.8200 187.2000 ;
      RECT 56.4200 186.1200 99.8200 187.2000 ;
      RECT 8.8600 186.1200 54.8200 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 240.1200 186.1200 ;
      RECT 238.8600 183.4000 240.1200 184.4800 ;
      RECT 193.6200 183.4000 235.2600 184.4800 ;
      RECT 148.6200 183.4000 192.0200 184.4800 ;
      RECT 103.6200 183.4000 147.0200 184.4800 ;
      RECT 58.6200 183.4000 102.0200 184.4800 ;
      RECT 13.6200 183.4000 57.0200 184.4800 ;
      RECT 4.8600 183.4000 12.0200 184.4800 ;
      RECT 0.0000 183.4000 1.2600 184.4800 ;
      RECT 0.0000 181.7600 240.1200 183.4000 ;
      RECT 234.8600 180.6800 240.1200 181.7600 ;
      RECT 191.4200 180.6800 231.2600 181.7600 ;
      RECT 146.4200 180.6800 189.8200 181.7600 ;
      RECT 101.4200 180.6800 144.8200 181.7600 ;
      RECT 56.4200 180.6800 99.8200 181.7600 ;
      RECT 8.8600 180.6800 54.8200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 240.1200 180.6800 ;
      RECT 238.8600 177.9600 240.1200 179.0400 ;
      RECT 193.6200 177.9600 235.2600 179.0400 ;
      RECT 148.6200 177.9600 192.0200 179.0400 ;
      RECT 103.6200 177.9600 147.0200 179.0400 ;
      RECT 58.6200 177.9600 102.0200 179.0400 ;
      RECT 13.6200 177.9600 57.0200 179.0400 ;
      RECT 4.8600 177.9600 12.0200 179.0400 ;
      RECT 0.0000 177.9600 1.2600 179.0400 ;
      RECT 0.0000 176.3200 240.1200 177.9600 ;
      RECT 234.8600 175.2400 240.1200 176.3200 ;
      RECT 191.4200 175.2400 231.2600 176.3200 ;
      RECT 146.4200 175.2400 189.8200 176.3200 ;
      RECT 101.4200 175.2400 144.8200 176.3200 ;
      RECT 56.4200 175.2400 99.8200 176.3200 ;
      RECT 8.8600 175.2400 54.8200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 240.1200 175.2400 ;
      RECT 238.8600 172.5200 240.1200 173.6000 ;
      RECT 193.6200 172.5200 235.2600 173.6000 ;
      RECT 148.6200 172.5200 192.0200 173.6000 ;
      RECT 103.6200 172.5200 147.0200 173.6000 ;
      RECT 58.6200 172.5200 102.0200 173.6000 ;
      RECT 13.6200 172.5200 57.0200 173.6000 ;
      RECT 4.8600 172.5200 12.0200 173.6000 ;
      RECT 0.0000 172.5200 1.2600 173.6000 ;
      RECT 0.0000 170.8800 240.1200 172.5200 ;
      RECT 234.8600 169.8000 240.1200 170.8800 ;
      RECT 191.4200 169.8000 231.2600 170.8800 ;
      RECT 146.4200 169.8000 189.8200 170.8800 ;
      RECT 101.4200 169.8000 144.8200 170.8800 ;
      RECT 56.4200 169.8000 99.8200 170.8800 ;
      RECT 8.8600 169.8000 54.8200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 240.1200 169.8000 ;
      RECT 238.8600 167.0800 240.1200 168.1600 ;
      RECT 193.6200 167.0800 235.2600 168.1600 ;
      RECT 148.6200 167.0800 192.0200 168.1600 ;
      RECT 103.6200 167.0800 147.0200 168.1600 ;
      RECT 58.6200 167.0800 102.0200 168.1600 ;
      RECT 13.6200 167.0800 57.0200 168.1600 ;
      RECT 4.8600 167.0800 12.0200 168.1600 ;
      RECT 0.0000 167.0800 1.2600 168.1600 ;
      RECT 0.0000 165.4400 240.1200 167.0800 ;
      RECT 234.8600 164.3600 240.1200 165.4400 ;
      RECT 191.4200 164.3600 231.2600 165.4400 ;
      RECT 146.4200 164.3600 189.8200 165.4400 ;
      RECT 101.4200 164.3600 144.8200 165.4400 ;
      RECT 56.4200 164.3600 99.8200 165.4400 ;
      RECT 8.8600 164.3600 54.8200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 240.1200 164.3600 ;
      RECT 238.8600 161.6400 240.1200 162.7200 ;
      RECT 193.6200 161.6400 235.2600 162.7200 ;
      RECT 148.6200 161.6400 192.0200 162.7200 ;
      RECT 103.6200 161.6400 147.0200 162.7200 ;
      RECT 58.6200 161.6400 102.0200 162.7200 ;
      RECT 13.6200 161.6400 57.0200 162.7200 ;
      RECT 4.8600 161.6400 12.0200 162.7200 ;
      RECT 0.0000 161.6400 1.2600 162.7200 ;
      RECT 0.0000 160.0000 240.1200 161.6400 ;
      RECT 234.8600 158.9200 240.1200 160.0000 ;
      RECT 191.4200 158.9200 231.2600 160.0000 ;
      RECT 146.4200 158.9200 189.8200 160.0000 ;
      RECT 101.4200 158.9200 144.8200 160.0000 ;
      RECT 56.4200 158.9200 99.8200 160.0000 ;
      RECT 8.8600 158.9200 54.8200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 240.1200 158.9200 ;
      RECT 238.8600 156.2000 240.1200 157.2800 ;
      RECT 193.6200 156.2000 235.2600 157.2800 ;
      RECT 148.6200 156.2000 192.0200 157.2800 ;
      RECT 103.6200 156.2000 147.0200 157.2800 ;
      RECT 58.6200 156.2000 102.0200 157.2800 ;
      RECT 13.6200 156.2000 57.0200 157.2800 ;
      RECT 4.8600 156.2000 12.0200 157.2800 ;
      RECT 0.0000 156.2000 1.2600 157.2800 ;
      RECT 0.0000 154.5600 240.1200 156.2000 ;
      RECT 234.8600 153.4800 240.1200 154.5600 ;
      RECT 191.4200 153.4800 231.2600 154.5600 ;
      RECT 146.4200 153.4800 189.8200 154.5600 ;
      RECT 101.4200 153.4800 144.8200 154.5600 ;
      RECT 56.4200 153.4800 99.8200 154.5600 ;
      RECT 8.8600 153.4800 54.8200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 240.1200 153.4800 ;
      RECT 238.8600 150.7600 240.1200 151.8400 ;
      RECT 193.6200 150.7600 235.2600 151.8400 ;
      RECT 148.6200 150.7600 192.0200 151.8400 ;
      RECT 103.6200 150.7600 147.0200 151.8400 ;
      RECT 58.6200 150.7600 102.0200 151.8400 ;
      RECT 13.6200 150.7600 57.0200 151.8400 ;
      RECT 4.8600 150.7600 12.0200 151.8400 ;
      RECT 0.0000 150.7600 1.2600 151.8400 ;
      RECT 0.0000 149.1200 240.1200 150.7600 ;
      RECT 234.8600 148.0400 240.1200 149.1200 ;
      RECT 191.4200 148.0400 231.2600 149.1200 ;
      RECT 146.4200 148.0400 189.8200 149.1200 ;
      RECT 101.4200 148.0400 144.8200 149.1200 ;
      RECT 56.4200 148.0400 99.8200 149.1200 ;
      RECT 8.8600 148.0400 54.8200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 240.1200 148.0400 ;
      RECT 238.8600 145.3200 240.1200 146.4000 ;
      RECT 193.6200 145.3200 235.2600 146.4000 ;
      RECT 148.6200 145.3200 192.0200 146.4000 ;
      RECT 103.6200 145.3200 147.0200 146.4000 ;
      RECT 58.6200 145.3200 102.0200 146.4000 ;
      RECT 13.6200 145.3200 57.0200 146.4000 ;
      RECT 4.8600 145.3200 12.0200 146.4000 ;
      RECT 0.0000 145.3200 1.2600 146.4000 ;
      RECT 0.0000 143.6800 240.1200 145.3200 ;
      RECT 234.8600 142.6000 240.1200 143.6800 ;
      RECT 191.4200 142.6000 231.2600 143.6800 ;
      RECT 146.4200 142.6000 189.8200 143.6800 ;
      RECT 101.4200 142.6000 144.8200 143.6800 ;
      RECT 56.4200 142.6000 99.8200 143.6800 ;
      RECT 8.8600 142.6000 54.8200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 240.1200 142.6000 ;
      RECT 238.8600 139.8800 240.1200 140.9600 ;
      RECT 193.6200 139.8800 235.2600 140.9600 ;
      RECT 148.6200 139.8800 192.0200 140.9600 ;
      RECT 103.6200 139.8800 147.0200 140.9600 ;
      RECT 58.6200 139.8800 102.0200 140.9600 ;
      RECT 13.6200 139.8800 57.0200 140.9600 ;
      RECT 4.8600 139.8800 12.0200 140.9600 ;
      RECT 0.0000 139.8800 1.2600 140.9600 ;
      RECT 0.0000 138.2400 240.1200 139.8800 ;
      RECT 234.8600 137.1600 240.1200 138.2400 ;
      RECT 191.4200 137.1600 231.2600 138.2400 ;
      RECT 146.4200 137.1600 189.8200 138.2400 ;
      RECT 101.4200 137.1600 144.8200 138.2400 ;
      RECT 56.4200 137.1600 99.8200 138.2400 ;
      RECT 8.8600 137.1600 54.8200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 240.1200 137.1600 ;
      RECT 238.8600 134.4400 240.1200 135.5200 ;
      RECT 193.6200 134.4400 235.2600 135.5200 ;
      RECT 148.6200 134.4400 192.0200 135.5200 ;
      RECT 103.6200 134.4400 147.0200 135.5200 ;
      RECT 58.6200 134.4400 102.0200 135.5200 ;
      RECT 13.6200 134.4400 57.0200 135.5200 ;
      RECT 4.8600 134.4400 12.0200 135.5200 ;
      RECT 0.0000 134.4400 1.2600 135.5200 ;
      RECT 0.0000 132.8000 240.1200 134.4400 ;
      RECT 234.8600 131.7200 240.1200 132.8000 ;
      RECT 191.4200 131.7200 231.2600 132.8000 ;
      RECT 146.4200 131.7200 189.8200 132.8000 ;
      RECT 101.4200 131.7200 144.8200 132.8000 ;
      RECT 56.4200 131.7200 99.8200 132.8000 ;
      RECT 8.8600 131.7200 54.8200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 240.1200 131.7200 ;
      RECT 238.8600 129.0000 240.1200 130.0800 ;
      RECT 193.6200 129.0000 235.2600 130.0800 ;
      RECT 148.6200 129.0000 192.0200 130.0800 ;
      RECT 103.6200 129.0000 147.0200 130.0800 ;
      RECT 58.6200 129.0000 102.0200 130.0800 ;
      RECT 13.6200 129.0000 57.0200 130.0800 ;
      RECT 4.8600 129.0000 12.0200 130.0800 ;
      RECT 0.0000 129.0000 1.2600 130.0800 ;
      RECT 0.0000 127.3600 240.1200 129.0000 ;
      RECT 234.8600 126.2800 240.1200 127.3600 ;
      RECT 191.4200 126.2800 231.2600 127.3600 ;
      RECT 146.4200 126.2800 189.8200 127.3600 ;
      RECT 101.4200 126.2800 144.8200 127.3600 ;
      RECT 56.4200 126.2800 99.8200 127.3600 ;
      RECT 8.8600 126.2800 54.8200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 240.1200 126.2800 ;
      RECT 238.8600 123.5600 240.1200 124.6400 ;
      RECT 193.6200 123.5600 235.2600 124.6400 ;
      RECT 148.6200 123.5600 192.0200 124.6400 ;
      RECT 103.6200 123.5600 147.0200 124.6400 ;
      RECT 58.6200 123.5600 102.0200 124.6400 ;
      RECT 13.6200 123.5600 57.0200 124.6400 ;
      RECT 4.8600 123.5600 12.0200 124.6400 ;
      RECT 0.0000 123.5600 1.2600 124.6400 ;
      RECT 0.0000 121.9200 240.1200 123.5600 ;
      RECT 234.8600 120.8400 240.1200 121.9200 ;
      RECT 191.4200 120.8400 231.2600 121.9200 ;
      RECT 146.4200 120.8400 189.8200 121.9200 ;
      RECT 101.4200 120.8400 144.8200 121.9200 ;
      RECT 56.4200 120.8400 99.8200 121.9200 ;
      RECT 8.8600 120.8400 54.8200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 240.1200 120.8400 ;
      RECT 238.8600 118.1200 240.1200 119.2000 ;
      RECT 193.6200 118.1200 235.2600 119.2000 ;
      RECT 148.6200 118.1200 192.0200 119.2000 ;
      RECT 103.6200 118.1200 147.0200 119.2000 ;
      RECT 58.6200 118.1200 102.0200 119.2000 ;
      RECT 13.6200 118.1200 57.0200 119.2000 ;
      RECT 4.8600 118.1200 12.0200 119.2000 ;
      RECT 0.0000 118.1200 1.2600 119.2000 ;
      RECT 0.0000 116.4800 240.1200 118.1200 ;
      RECT 234.8600 115.4000 240.1200 116.4800 ;
      RECT 191.4200 115.4000 231.2600 116.4800 ;
      RECT 146.4200 115.4000 189.8200 116.4800 ;
      RECT 101.4200 115.4000 144.8200 116.4800 ;
      RECT 56.4200 115.4000 99.8200 116.4800 ;
      RECT 8.8600 115.4000 54.8200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 240.1200 115.4000 ;
      RECT 238.8600 112.6800 240.1200 113.7600 ;
      RECT 193.6200 112.6800 235.2600 113.7600 ;
      RECT 148.6200 112.6800 192.0200 113.7600 ;
      RECT 103.6200 112.6800 147.0200 113.7600 ;
      RECT 58.6200 112.6800 102.0200 113.7600 ;
      RECT 13.6200 112.6800 57.0200 113.7600 ;
      RECT 4.8600 112.6800 12.0200 113.7600 ;
      RECT 0.0000 112.6800 1.2600 113.7600 ;
      RECT 0.0000 111.0400 240.1200 112.6800 ;
      RECT 234.8600 109.9600 240.1200 111.0400 ;
      RECT 191.4200 109.9600 231.2600 111.0400 ;
      RECT 146.4200 109.9600 189.8200 111.0400 ;
      RECT 101.4200 109.9600 144.8200 111.0400 ;
      RECT 56.4200 109.9600 99.8200 111.0400 ;
      RECT 8.8600 109.9600 54.8200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 240.1200 109.9600 ;
      RECT 238.8600 107.2400 240.1200 108.3200 ;
      RECT 193.6200 107.2400 235.2600 108.3200 ;
      RECT 148.6200 107.2400 192.0200 108.3200 ;
      RECT 103.6200 107.2400 147.0200 108.3200 ;
      RECT 58.6200 107.2400 102.0200 108.3200 ;
      RECT 13.6200 107.2400 57.0200 108.3200 ;
      RECT 4.8600 107.2400 12.0200 108.3200 ;
      RECT 0.0000 107.2400 1.2600 108.3200 ;
      RECT 0.0000 105.6000 240.1200 107.2400 ;
      RECT 234.8600 104.5200 240.1200 105.6000 ;
      RECT 191.4200 104.5200 231.2600 105.6000 ;
      RECT 146.4200 104.5200 189.8200 105.6000 ;
      RECT 101.4200 104.5200 144.8200 105.6000 ;
      RECT 56.4200 104.5200 99.8200 105.6000 ;
      RECT 8.8600 104.5200 54.8200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 240.1200 104.5200 ;
      RECT 238.8600 101.8000 240.1200 102.8800 ;
      RECT 193.6200 101.8000 235.2600 102.8800 ;
      RECT 148.6200 101.8000 192.0200 102.8800 ;
      RECT 103.6200 101.8000 147.0200 102.8800 ;
      RECT 58.6200 101.8000 102.0200 102.8800 ;
      RECT 13.6200 101.8000 57.0200 102.8800 ;
      RECT 4.8600 101.8000 12.0200 102.8800 ;
      RECT 0.0000 101.8000 1.2600 102.8800 ;
      RECT 0.0000 100.1600 240.1200 101.8000 ;
      RECT 234.8600 99.0800 240.1200 100.1600 ;
      RECT 191.4200 99.0800 231.2600 100.1600 ;
      RECT 146.4200 99.0800 189.8200 100.1600 ;
      RECT 101.4200 99.0800 144.8200 100.1600 ;
      RECT 56.4200 99.0800 99.8200 100.1600 ;
      RECT 8.8600 99.0800 54.8200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 240.1200 99.0800 ;
      RECT 238.8600 96.3600 240.1200 97.4400 ;
      RECT 193.6200 96.3600 235.2600 97.4400 ;
      RECT 148.6200 96.3600 192.0200 97.4400 ;
      RECT 103.6200 96.3600 147.0200 97.4400 ;
      RECT 58.6200 96.3600 102.0200 97.4400 ;
      RECT 13.6200 96.3600 57.0200 97.4400 ;
      RECT 4.8600 96.3600 12.0200 97.4400 ;
      RECT 0.0000 96.3600 1.2600 97.4400 ;
      RECT 0.0000 94.7200 240.1200 96.3600 ;
      RECT 234.8600 93.6400 240.1200 94.7200 ;
      RECT 191.4200 93.6400 231.2600 94.7200 ;
      RECT 146.4200 93.6400 189.8200 94.7200 ;
      RECT 101.4200 93.6400 144.8200 94.7200 ;
      RECT 56.4200 93.6400 99.8200 94.7200 ;
      RECT 8.8600 93.6400 54.8200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 240.1200 93.6400 ;
      RECT 238.8600 90.9200 240.1200 92.0000 ;
      RECT 193.6200 90.9200 235.2600 92.0000 ;
      RECT 148.6200 90.9200 192.0200 92.0000 ;
      RECT 103.6200 90.9200 147.0200 92.0000 ;
      RECT 58.6200 90.9200 102.0200 92.0000 ;
      RECT 13.6200 90.9200 57.0200 92.0000 ;
      RECT 4.8600 90.9200 12.0200 92.0000 ;
      RECT 0.0000 90.9200 1.2600 92.0000 ;
      RECT 0.0000 89.2800 240.1200 90.9200 ;
      RECT 234.8600 88.2000 240.1200 89.2800 ;
      RECT 191.4200 88.2000 231.2600 89.2800 ;
      RECT 146.4200 88.2000 189.8200 89.2800 ;
      RECT 101.4200 88.2000 144.8200 89.2800 ;
      RECT 56.4200 88.2000 99.8200 89.2800 ;
      RECT 8.8600 88.2000 54.8200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 240.1200 88.2000 ;
      RECT 238.8600 85.4800 240.1200 86.5600 ;
      RECT 193.6200 85.4800 235.2600 86.5600 ;
      RECT 148.6200 85.4800 192.0200 86.5600 ;
      RECT 103.6200 85.4800 147.0200 86.5600 ;
      RECT 58.6200 85.4800 102.0200 86.5600 ;
      RECT 13.6200 85.4800 57.0200 86.5600 ;
      RECT 4.8600 85.4800 12.0200 86.5600 ;
      RECT 0.0000 85.4800 1.2600 86.5600 ;
      RECT 0.0000 83.8400 240.1200 85.4800 ;
      RECT 234.8600 82.7600 240.1200 83.8400 ;
      RECT 191.4200 82.7600 231.2600 83.8400 ;
      RECT 146.4200 82.7600 189.8200 83.8400 ;
      RECT 101.4200 82.7600 144.8200 83.8400 ;
      RECT 56.4200 82.7600 99.8200 83.8400 ;
      RECT 8.8600 82.7600 54.8200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 240.1200 82.7600 ;
      RECT 238.8600 80.0400 240.1200 81.1200 ;
      RECT 193.6200 80.0400 235.2600 81.1200 ;
      RECT 148.6200 80.0400 192.0200 81.1200 ;
      RECT 103.6200 80.0400 147.0200 81.1200 ;
      RECT 58.6200 80.0400 102.0200 81.1200 ;
      RECT 13.6200 80.0400 57.0200 81.1200 ;
      RECT 4.8600 80.0400 12.0200 81.1200 ;
      RECT 0.0000 80.0400 1.2600 81.1200 ;
      RECT 0.0000 78.4000 240.1200 80.0400 ;
      RECT 234.8600 77.3200 240.1200 78.4000 ;
      RECT 191.4200 77.3200 231.2600 78.4000 ;
      RECT 146.4200 77.3200 189.8200 78.4000 ;
      RECT 101.4200 77.3200 144.8200 78.4000 ;
      RECT 56.4200 77.3200 99.8200 78.4000 ;
      RECT 8.8600 77.3200 54.8200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 240.1200 77.3200 ;
      RECT 238.8600 74.6000 240.1200 75.6800 ;
      RECT 193.6200 74.6000 235.2600 75.6800 ;
      RECT 148.6200 74.6000 192.0200 75.6800 ;
      RECT 103.6200 74.6000 147.0200 75.6800 ;
      RECT 58.6200 74.6000 102.0200 75.6800 ;
      RECT 13.6200 74.6000 57.0200 75.6800 ;
      RECT 4.8600 74.6000 12.0200 75.6800 ;
      RECT 0.0000 74.6000 1.2600 75.6800 ;
      RECT 0.0000 72.9600 240.1200 74.6000 ;
      RECT 234.8600 71.8800 240.1200 72.9600 ;
      RECT 191.4200 71.8800 231.2600 72.9600 ;
      RECT 146.4200 71.8800 189.8200 72.9600 ;
      RECT 101.4200 71.8800 144.8200 72.9600 ;
      RECT 56.4200 71.8800 99.8200 72.9600 ;
      RECT 8.8600 71.8800 54.8200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 240.1200 71.8800 ;
      RECT 238.8600 69.1600 240.1200 70.2400 ;
      RECT 193.6200 69.1600 235.2600 70.2400 ;
      RECT 148.6200 69.1600 192.0200 70.2400 ;
      RECT 103.6200 69.1600 147.0200 70.2400 ;
      RECT 58.6200 69.1600 102.0200 70.2400 ;
      RECT 13.6200 69.1600 57.0200 70.2400 ;
      RECT 4.8600 69.1600 12.0200 70.2400 ;
      RECT 0.0000 69.1600 1.2600 70.2400 ;
      RECT 0.0000 67.5200 240.1200 69.1600 ;
      RECT 234.8600 66.4400 240.1200 67.5200 ;
      RECT 191.4200 66.4400 231.2600 67.5200 ;
      RECT 146.4200 66.4400 189.8200 67.5200 ;
      RECT 101.4200 66.4400 144.8200 67.5200 ;
      RECT 56.4200 66.4400 99.8200 67.5200 ;
      RECT 8.8600 66.4400 54.8200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 240.1200 66.4400 ;
      RECT 238.8600 63.7200 240.1200 64.8000 ;
      RECT 193.6200 63.7200 235.2600 64.8000 ;
      RECT 148.6200 63.7200 192.0200 64.8000 ;
      RECT 103.6200 63.7200 147.0200 64.8000 ;
      RECT 58.6200 63.7200 102.0200 64.8000 ;
      RECT 13.6200 63.7200 57.0200 64.8000 ;
      RECT 4.8600 63.7200 12.0200 64.8000 ;
      RECT 0.0000 63.7200 1.2600 64.8000 ;
      RECT 0.0000 62.0800 240.1200 63.7200 ;
      RECT 234.8600 61.0000 240.1200 62.0800 ;
      RECT 191.4200 61.0000 231.2600 62.0800 ;
      RECT 146.4200 61.0000 189.8200 62.0800 ;
      RECT 101.4200 61.0000 144.8200 62.0800 ;
      RECT 56.4200 61.0000 99.8200 62.0800 ;
      RECT 8.8600 61.0000 54.8200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 240.1200 61.0000 ;
      RECT 238.8600 58.2800 240.1200 59.3600 ;
      RECT 193.6200 58.2800 235.2600 59.3600 ;
      RECT 148.6200 58.2800 192.0200 59.3600 ;
      RECT 103.6200 58.2800 147.0200 59.3600 ;
      RECT 58.6200 58.2800 102.0200 59.3600 ;
      RECT 13.6200 58.2800 57.0200 59.3600 ;
      RECT 4.8600 58.2800 12.0200 59.3600 ;
      RECT 0.0000 58.2800 1.2600 59.3600 ;
      RECT 0.0000 56.6400 240.1200 58.2800 ;
      RECT 234.8600 55.5600 240.1200 56.6400 ;
      RECT 191.4200 55.5600 231.2600 56.6400 ;
      RECT 146.4200 55.5600 189.8200 56.6400 ;
      RECT 101.4200 55.5600 144.8200 56.6400 ;
      RECT 56.4200 55.5600 99.8200 56.6400 ;
      RECT 8.8600 55.5600 54.8200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 240.1200 55.5600 ;
      RECT 238.8600 52.8400 240.1200 53.9200 ;
      RECT 193.6200 52.8400 235.2600 53.9200 ;
      RECT 148.6200 52.8400 192.0200 53.9200 ;
      RECT 103.6200 52.8400 147.0200 53.9200 ;
      RECT 58.6200 52.8400 102.0200 53.9200 ;
      RECT 13.6200 52.8400 57.0200 53.9200 ;
      RECT 4.8600 52.8400 12.0200 53.9200 ;
      RECT 0.0000 52.8400 1.2600 53.9200 ;
      RECT 0.0000 51.2000 240.1200 52.8400 ;
      RECT 234.8600 50.1200 240.1200 51.2000 ;
      RECT 191.4200 50.1200 231.2600 51.2000 ;
      RECT 146.4200 50.1200 189.8200 51.2000 ;
      RECT 101.4200 50.1200 144.8200 51.2000 ;
      RECT 56.4200 50.1200 99.8200 51.2000 ;
      RECT 8.8600 50.1200 54.8200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 240.1200 50.1200 ;
      RECT 238.8600 47.4000 240.1200 48.4800 ;
      RECT 193.6200 47.4000 235.2600 48.4800 ;
      RECT 148.6200 47.4000 192.0200 48.4800 ;
      RECT 103.6200 47.4000 147.0200 48.4800 ;
      RECT 58.6200 47.4000 102.0200 48.4800 ;
      RECT 13.6200 47.4000 57.0200 48.4800 ;
      RECT 4.8600 47.4000 12.0200 48.4800 ;
      RECT 0.0000 47.4000 1.2600 48.4800 ;
      RECT 0.0000 45.7600 240.1200 47.4000 ;
      RECT 234.8600 44.6800 240.1200 45.7600 ;
      RECT 191.4200 44.6800 231.2600 45.7600 ;
      RECT 146.4200 44.6800 189.8200 45.7600 ;
      RECT 101.4200 44.6800 144.8200 45.7600 ;
      RECT 56.4200 44.6800 99.8200 45.7600 ;
      RECT 8.8600 44.6800 54.8200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 240.1200 44.6800 ;
      RECT 238.8600 41.9600 240.1200 43.0400 ;
      RECT 193.6200 41.9600 235.2600 43.0400 ;
      RECT 148.6200 41.9600 192.0200 43.0400 ;
      RECT 103.6200 41.9600 147.0200 43.0400 ;
      RECT 58.6200 41.9600 102.0200 43.0400 ;
      RECT 13.6200 41.9600 57.0200 43.0400 ;
      RECT 4.8600 41.9600 12.0200 43.0400 ;
      RECT 0.0000 41.9600 1.2600 43.0400 ;
      RECT 0.0000 40.3200 240.1200 41.9600 ;
      RECT 234.8600 39.2400 240.1200 40.3200 ;
      RECT 191.4200 39.2400 231.2600 40.3200 ;
      RECT 146.4200 39.2400 189.8200 40.3200 ;
      RECT 101.4200 39.2400 144.8200 40.3200 ;
      RECT 56.4200 39.2400 99.8200 40.3200 ;
      RECT 8.8600 39.2400 54.8200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 240.1200 39.2400 ;
      RECT 238.8600 36.5200 240.1200 37.6000 ;
      RECT 193.6200 36.5200 235.2600 37.6000 ;
      RECT 148.6200 36.5200 192.0200 37.6000 ;
      RECT 103.6200 36.5200 147.0200 37.6000 ;
      RECT 58.6200 36.5200 102.0200 37.6000 ;
      RECT 13.6200 36.5200 57.0200 37.6000 ;
      RECT 4.8600 36.5200 12.0200 37.6000 ;
      RECT 0.0000 36.5200 1.2600 37.6000 ;
      RECT 0.0000 34.8800 240.1200 36.5200 ;
      RECT 234.8600 33.8000 240.1200 34.8800 ;
      RECT 191.4200 33.8000 231.2600 34.8800 ;
      RECT 146.4200 33.8000 189.8200 34.8800 ;
      RECT 101.4200 33.8000 144.8200 34.8800 ;
      RECT 56.4200 33.8000 99.8200 34.8800 ;
      RECT 8.8600 33.8000 54.8200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 240.1200 33.8000 ;
      RECT 238.8600 31.0800 240.1200 32.1600 ;
      RECT 193.6200 31.0800 235.2600 32.1600 ;
      RECT 148.6200 31.0800 192.0200 32.1600 ;
      RECT 103.6200 31.0800 147.0200 32.1600 ;
      RECT 58.6200 31.0800 102.0200 32.1600 ;
      RECT 13.6200 31.0800 57.0200 32.1600 ;
      RECT 4.8600 31.0800 12.0200 32.1600 ;
      RECT 0.0000 31.0800 1.2600 32.1600 ;
      RECT 0.0000 29.4400 240.1200 31.0800 ;
      RECT 234.8600 28.3600 240.1200 29.4400 ;
      RECT 191.4200 28.3600 231.2600 29.4400 ;
      RECT 146.4200 28.3600 189.8200 29.4400 ;
      RECT 101.4200 28.3600 144.8200 29.4400 ;
      RECT 56.4200 28.3600 99.8200 29.4400 ;
      RECT 8.8600 28.3600 54.8200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 240.1200 28.3600 ;
      RECT 238.8600 25.6400 240.1200 26.7200 ;
      RECT 193.6200 25.6400 235.2600 26.7200 ;
      RECT 148.6200 25.6400 192.0200 26.7200 ;
      RECT 103.6200 25.6400 147.0200 26.7200 ;
      RECT 58.6200 25.6400 102.0200 26.7200 ;
      RECT 13.6200 25.6400 57.0200 26.7200 ;
      RECT 4.8600 25.6400 12.0200 26.7200 ;
      RECT 0.0000 25.6400 1.2600 26.7200 ;
      RECT 0.0000 24.0000 240.1200 25.6400 ;
      RECT 234.8600 22.9200 240.1200 24.0000 ;
      RECT 191.4200 22.9200 231.2600 24.0000 ;
      RECT 146.4200 22.9200 189.8200 24.0000 ;
      RECT 101.4200 22.9200 144.8200 24.0000 ;
      RECT 56.4200 22.9200 99.8200 24.0000 ;
      RECT 8.8600 22.9200 54.8200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 240.1200 22.9200 ;
      RECT 238.8600 20.2000 240.1200 21.2800 ;
      RECT 193.6200 20.2000 235.2600 21.2800 ;
      RECT 148.6200 20.2000 192.0200 21.2800 ;
      RECT 103.6200 20.2000 147.0200 21.2800 ;
      RECT 58.6200 20.2000 102.0200 21.2800 ;
      RECT 13.6200 20.2000 57.0200 21.2800 ;
      RECT 4.8600 20.2000 12.0200 21.2800 ;
      RECT 0.0000 20.2000 1.2600 21.2800 ;
      RECT 0.0000 18.5600 240.1200 20.2000 ;
      RECT 234.8600 17.4800 240.1200 18.5600 ;
      RECT 191.4200 17.4800 231.2600 18.5600 ;
      RECT 146.4200 17.4800 189.8200 18.5600 ;
      RECT 101.4200 17.4800 144.8200 18.5600 ;
      RECT 56.4200 17.4800 99.8200 18.5600 ;
      RECT 8.8600 17.4800 54.8200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 240.1200 17.4800 ;
      RECT 238.8600 14.7600 240.1200 15.8400 ;
      RECT 193.6200 14.7600 235.2600 15.8400 ;
      RECT 148.6200 14.7600 192.0200 15.8400 ;
      RECT 103.6200 14.7600 147.0200 15.8400 ;
      RECT 58.6200 14.7600 102.0200 15.8400 ;
      RECT 13.6200 14.7600 57.0200 15.8400 ;
      RECT 4.8600 14.7600 12.0200 15.8400 ;
      RECT 0.0000 14.7600 1.2600 15.8400 ;
      RECT 0.0000 13.1200 240.1200 14.7600 ;
      RECT 234.8600 12.0400 240.1200 13.1200 ;
      RECT 191.4200 12.0400 231.2600 13.1200 ;
      RECT 146.4200 12.0400 189.8200 13.1200 ;
      RECT 101.4200 12.0400 144.8200 13.1200 ;
      RECT 56.4200 12.0400 99.8200 13.1200 ;
      RECT 8.8600 12.0400 54.8200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 240.1200 12.0400 ;
      RECT 238.8600 9.3200 240.1200 10.4000 ;
      RECT 193.6200 9.3200 235.2600 10.4000 ;
      RECT 148.6200 9.3200 192.0200 10.4000 ;
      RECT 103.6200 9.3200 147.0200 10.4000 ;
      RECT 58.6200 9.3200 102.0200 10.4000 ;
      RECT 13.6200 9.3200 57.0200 10.4000 ;
      RECT 4.8600 9.3200 12.0200 10.4000 ;
      RECT 0.0000 9.3200 1.2600 10.4000 ;
      RECT 0.0000 8.7300 240.1200 9.3200 ;
      RECT 234.8600 5.1300 240.1200 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 240.1200 5.1300 ;
      RECT 238.8600 1.1300 240.1200 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 240.1200 1.1300 ;
    LAYER met4 ;
      RECT 0.0000 217.8300 240.1200 219.6400 ;
      RECT 193.6200 213.8300 235.2600 217.8300 ;
      RECT 148.6200 213.8300 192.0200 217.8300 ;
      RECT 103.6200 213.8300 147.0200 217.8300 ;
      RECT 58.6200 213.8300 102.0200 217.8300 ;
      RECT 13.6200 213.8300 57.0200 217.8300 ;
      RECT 4.8600 213.8300 12.0200 217.8300 ;
      RECT 234.8600 5.1300 235.2600 213.8300 ;
      RECT 193.6200 5.1300 231.2600 213.8300 ;
      RECT 191.4200 5.1300 192.0200 213.8300 ;
      RECT 148.6200 5.1300 189.8200 213.8300 ;
      RECT 146.4200 5.1300 147.0200 213.8300 ;
      RECT 103.6200 5.1300 144.8200 213.8300 ;
      RECT 101.4200 5.1300 102.0200 213.8300 ;
      RECT 58.6200 5.1300 99.8200 213.8300 ;
      RECT 56.4200 5.1300 57.0200 213.8300 ;
      RECT 13.6200 5.1300 54.8200 213.8300 ;
      RECT 8.8600 5.1300 12.0200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 238.8600 1.1300 240.1200 217.8300 ;
      RECT 193.6200 1.1300 235.2600 5.1300 ;
      RECT 148.6200 1.1300 192.0200 5.1300 ;
      RECT 103.6200 1.1300 147.0200 5.1300 ;
      RECT 58.6200 1.1300 102.0200 5.1300 ;
      RECT 13.6200 1.1300 57.0200 5.1300 ;
      RECT 4.8600 1.1300 12.0200 5.1300 ;
      RECT 0.0000 1.1300 1.2600 217.8300 ;
      RECT 0.0000 1.1000 240.1200 1.1300 ;
      RECT 90.1500 0.0000 240.1200 1.1000 ;
      RECT 0.0000 0.0000 89.2500 1.1000 ;
    LAYER met5 ;
      RECT 0.0000 0.0000 240.1200 219.6400 ;
  END
END RegFile

END LIBRARY
