magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 366 157 827 203
rect 1 21 827 157
rect 30 -17 64 21
<< locali >>
rect 659 353 725 425
rect 98 153 156 335
rect 381 325 725 353
rect 381 289 811 325
rect 190 153 256 255
rect 765 171 811 289
rect 659 127 811 171
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 369 69 493
rect 103 369 190 527
rect 17 123 64 369
rect 224 353 282 493
rect 320 421 362 493
rect 396 455 462 527
rect 496 459 811 493
rect 496 421 625 459
rect 320 387 625 421
rect 759 359 811 459
rect 224 289 347 353
rect 290 255 347 289
rect 290 205 593 255
rect 649 205 731 255
rect 17 56 69 123
rect 290 119 346 205
rect 103 17 170 119
rect 204 51 346 119
rect 380 131 625 171
rect 380 51 434 131
rect 468 17 534 97
rect 568 93 625 131
rect 568 55 810 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< obsm1 >>
rect 17 252 76 261
rect 664 252 722 261
rect 17 224 722 252
rect 17 215 76 224
rect 664 215 722 224
<< labels >>
rlabel locali s 98 153 156 335 6 A
port 1 nsew signal input
rlabel locali s 190 153 256 255 6 TE_B
port 2 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 827 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 366 157 827 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 659 127 811 171 6 Z
port 7 nsew signal output
rlabel locali s 765 171 811 289 6 Z
port 7 nsew signal output
rlabel locali s 381 289 811 325 6 Z
port 7 nsew signal output
rlabel locali s 381 325 725 353 6 Z
port 7 nsew signal output
rlabel locali s 659 353 725 425 6 Z
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2931524
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2924328
<< end >>
