magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -82 -26 282 226
<< mvnmos >>
rect 0 0 200 200
<< mvndiff >>
rect -56 182 0 200
rect -56 148 -45 182
rect -11 148 0 182
rect -56 114 0 148
rect -56 80 -45 114
rect -11 80 0 114
rect -56 46 0 80
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 200 182 256 200
rect 200 148 211 182
rect 245 148 256 182
rect 200 114 256 148
rect 200 80 211 114
rect 245 80 256 114
rect 200 46 256 80
rect 200 12 211 46
rect 245 12 256 46
rect 200 0 256 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 211 148 245 182
rect 211 80 245 114
rect 211 12 245 46
<< poly >>
rect 0 200 200 232
rect 0 -32 200 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 211 182 245 198
rect 211 114 245 148
rect 211 46 245 80
rect 211 -4 245 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_1
timestamp 1707688321
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 228 97 228 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85636082
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85635188
<< end >>
