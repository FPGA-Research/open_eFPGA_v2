magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -79 -26 207 226
<< nmos >>
rect 0 0 36 200
rect 92 0 128 200
<< ndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 36 182 92 200
rect 36 148 47 182
rect 81 148 92 182
rect 36 114 92 148
rect 36 80 47 114
rect 81 80 92 114
rect 36 46 92 80
rect 36 12 47 46
rect 81 12 92 46
rect 36 0 92 12
rect 128 182 181 200
rect 128 148 139 182
rect 173 148 181 182
rect 128 114 181 148
rect 128 80 139 114
rect 173 80 181 114
rect 128 46 181 80
rect 128 12 139 46
rect 173 12 181 46
rect 128 0 181 12
<< ndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 47 148 81 182
rect 47 80 81 114
rect 47 12 81 46
rect 139 148 173 182
rect 139 80 173 114
rect 139 12 173 46
<< poly >>
rect 0 200 36 226
rect 92 200 128 226
rect 0 -26 36 0
rect 92 -26 128 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 47 182 81 198
rect 47 114 81 148
rect 47 46 81 80
rect 47 -4 81 12
rect 139 182 173 198
rect 139 114 173 148
rect 139 46 173 80
rect 139 -4 173 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1707688321
transform 1 0 36 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_1
timestamp 1707688321
transform 1 0 128 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 64 97 64 97 0 FreeSans 300 0 0 0 D
flabel comment s 156 97 156 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 79588968
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79587642
<< end >>
