magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 2727 1126 2895
rect 0 168 168 2727
rect 958 168 1126 2727
rect 0 0 1126 168
<< pwell >>
rect 228 2581 898 2667
rect 228 314 314 2581
rect 812 314 898 2581
rect 228 228 898 314
<< mvpsubdiff >>
rect 254 2607 278 2641
rect 312 2607 351 2641
rect 385 2607 423 2641
rect 457 2607 495 2641
rect 529 2607 567 2641
rect 601 2607 701 2641
rect 735 2617 872 2641
rect 735 2607 838 2617
rect 254 2547 288 2607
rect 254 2478 288 2513
rect 254 2409 288 2444
rect 254 2340 288 2375
rect 254 2271 288 2306
rect 254 2202 288 2237
rect 254 2132 288 2168
rect 254 2062 288 2098
rect 254 1992 288 2028
rect 254 1922 288 1958
rect 254 1852 288 1888
rect 254 1782 288 1818
rect 254 1712 288 1748
rect 254 1642 288 1678
rect 254 1572 288 1608
rect 254 1502 288 1538
rect 838 2547 872 2583
rect 838 2477 872 2513
rect 838 2407 872 2443
rect 838 2337 872 2373
rect 838 2267 872 2303
rect 838 2197 872 2233
rect 838 2127 872 2163
rect 838 2057 872 2093
rect 838 1987 872 2023
rect 838 1917 872 1953
rect 838 1847 872 1883
rect 838 1777 872 1813
rect 838 1707 872 1743
rect 838 1637 872 1673
rect 838 1567 872 1603
rect 254 1432 288 1468
rect 838 1497 872 1533
rect 254 1362 288 1398
rect 254 1292 288 1328
rect 254 1222 288 1258
rect 254 1152 288 1188
rect 254 1082 288 1118
rect 254 1012 288 1048
rect 254 942 288 978
rect 254 872 288 908
rect 254 802 288 838
rect 254 732 288 768
rect 254 662 288 698
rect 254 592 288 628
rect 254 522 288 558
rect 254 452 288 488
rect 254 382 288 418
rect 838 1427 872 1463
rect 838 1357 872 1393
rect 838 1287 872 1323
rect 838 1217 872 1253
rect 838 1147 872 1183
rect 838 1077 872 1113
rect 838 1007 872 1043
rect 838 937 872 973
rect 838 867 872 903
rect 838 797 872 833
rect 838 727 872 763
rect 838 658 872 693
rect 838 589 872 624
rect 838 520 872 555
rect 838 451 872 486
rect 254 312 288 348
rect 838 382 872 417
rect 838 288 872 348
rect 288 278 360 288
rect 254 254 360 278
rect 394 254 435 288
rect 469 254 510 288
rect 544 254 586 288
rect 620 254 662 288
rect 696 254 738 288
rect 772 254 814 288
rect 848 254 872 288
<< mvnsubdiff >>
rect 68 2794 1058 2828
rect 68 2678 102 2794
rect 68 2609 102 2644
rect 68 2540 102 2575
rect 68 2471 102 2506
rect 68 2401 102 2437
rect 68 2331 102 2367
rect 68 2261 102 2297
rect 68 2191 102 2227
rect 68 2121 102 2157
rect 68 2051 102 2087
rect 68 1981 102 2017
rect 68 1911 102 1947
rect 68 1841 102 1877
rect 68 1771 102 1807
rect 68 1701 102 1737
rect 68 1631 102 1667
rect 68 1561 102 1597
rect 68 1491 102 1527
rect 68 1421 102 1457
rect 68 1351 102 1387
rect 68 1281 102 1317
rect 68 1211 102 1247
rect 68 1141 102 1177
rect 68 1071 102 1107
rect 68 1001 102 1037
rect 68 931 102 967
rect 68 861 102 897
rect 68 791 102 827
rect 68 721 102 757
rect 68 651 102 687
rect 68 581 102 617
rect 68 511 102 547
rect 68 441 102 477
rect 68 371 102 407
rect 68 301 102 337
rect 68 231 102 267
rect 68 101 102 197
rect 1024 101 1058 2794
rect 68 67 203 101
rect 237 67 277 101
rect 311 67 351 101
rect 385 67 425 101
rect 459 67 499 101
rect 533 67 573 101
rect 607 67 647 101
rect 681 67 721 101
rect 755 67 796 101
rect 830 67 871 101
rect 905 67 946 101
rect 980 67 1058 101
<< mvpsubdiffcont >>
rect 278 2607 312 2641
rect 351 2607 385 2641
rect 423 2607 457 2641
rect 495 2607 529 2641
rect 567 2607 601 2641
rect 701 2607 735 2641
rect 254 2513 288 2547
rect 254 2444 288 2478
rect 254 2375 288 2409
rect 254 2306 288 2340
rect 254 2237 288 2271
rect 254 2168 288 2202
rect 254 2098 288 2132
rect 254 2028 288 2062
rect 254 1958 288 1992
rect 254 1888 288 1922
rect 254 1818 288 1852
rect 254 1748 288 1782
rect 254 1678 288 1712
rect 254 1608 288 1642
rect 254 1538 288 1572
rect 838 2583 872 2617
rect 838 2513 872 2547
rect 838 2443 872 2477
rect 838 2373 872 2407
rect 838 2303 872 2337
rect 838 2233 872 2267
rect 838 2163 872 2197
rect 838 2093 872 2127
rect 838 2023 872 2057
rect 838 1953 872 1987
rect 838 1883 872 1917
rect 838 1813 872 1847
rect 838 1743 872 1777
rect 838 1673 872 1707
rect 838 1603 872 1637
rect 838 1533 872 1567
rect 254 1468 288 1502
rect 838 1463 872 1497
rect 254 1398 288 1432
rect 254 1328 288 1362
rect 254 1258 288 1292
rect 254 1188 288 1222
rect 254 1118 288 1152
rect 254 1048 288 1082
rect 254 978 288 1012
rect 254 908 288 942
rect 254 838 288 872
rect 254 768 288 802
rect 254 698 288 732
rect 254 628 288 662
rect 254 558 288 592
rect 254 488 288 522
rect 254 418 288 452
rect 838 1393 872 1427
rect 838 1323 872 1357
rect 838 1253 872 1287
rect 838 1183 872 1217
rect 838 1113 872 1147
rect 838 1043 872 1077
rect 838 973 872 1007
rect 838 903 872 937
rect 838 833 872 867
rect 838 763 872 797
rect 838 693 872 727
rect 838 624 872 658
rect 838 555 872 589
rect 838 486 872 520
rect 838 417 872 451
rect 254 348 288 382
rect 838 348 872 382
rect 254 278 288 312
rect 360 254 394 288
rect 435 254 469 288
rect 510 254 544 288
rect 586 254 620 288
rect 662 254 696 288
rect 738 254 772 288
rect 814 254 848 288
<< mvnsubdiffcont >>
rect 68 2644 102 2678
rect 68 2575 102 2609
rect 68 2506 102 2540
rect 68 2437 102 2471
rect 68 2367 102 2401
rect 68 2297 102 2331
rect 68 2227 102 2261
rect 68 2157 102 2191
rect 68 2087 102 2121
rect 68 2017 102 2051
rect 68 1947 102 1981
rect 68 1877 102 1911
rect 68 1807 102 1841
rect 68 1737 102 1771
rect 68 1667 102 1701
rect 68 1597 102 1631
rect 68 1527 102 1561
rect 68 1457 102 1491
rect 68 1387 102 1421
rect 68 1317 102 1351
rect 68 1247 102 1281
rect 68 1177 102 1211
rect 68 1107 102 1141
rect 68 1037 102 1071
rect 68 967 102 1001
rect 68 897 102 931
rect 68 827 102 861
rect 68 757 102 791
rect 68 687 102 721
rect 68 617 102 651
rect 68 547 102 581
rect 68 477 102 511
rect 68 407 102 441
rect 68 337 102 371
rect 68 267 102 301
rect 68 197 102 231
rect 203 67 237 101
rect 277 67 311 101
rect 351 67 385 101
rect 425 67 459 101
rect 499 67 533 101
rect 573 67 607 101
rect 647 67 681 101
rect 721 67 755 101
rect 796 67 830 101
rect 871 67 905 101
rect 946 67 980 101
<< poly >>
rect 415 1491 711 1507
rect 415 1457 444 1491
rect 478 1457 512 1491
rect 546 1457 580 1491
rect 614 1457 648 1491
rect 682 1457 711 1491
rect 415 1438 711 1457
rect 415 370 711 386
rect 415 336 449 370
rect 483 336 517 370
rect 551 336 585 370
rect 619 336 653 370
rect 687 336 711 370
rect 415 320 711 336
<< polycont >>
rect 444 1457 478 1491
rect 512 1457 546 1491
rect 580 1457 614 1491
rect 648 1457 682 1491
rect 449 336 483 370
rect 517 336 551 370
rect 585 336 619 370
rect 653 336 687 370
<< locali >>
rect 68 2794 1058 2828
rect 68 2724 102 2794
rect 68 2678 102 2690
rect 68 2609 102 2616
rect 68 2540 102 2542
rect 68 2502 102 2506
rect 68 2428 102 2437
rect 68 2354 102 2367
rect 68 2280 102 2297
rect 68 2206 102 2227
rect 68 2132 102 2157
rect 68 2058 102 2087
rect 68 1984 102 2017
rect 68 1911 102 1947
rect 68 1841 102 1876
rect 68 1771 102 1802
rect 68 1701 102 1728
rect 68 1631 102 1654
rect 68 1561 102 1580
rect 68 1491 102 1506
rect 68 1421 102 1432
rect 68 1351 102 1358
rect 68 1281 102 1284
rect 68 1244 102 1247
rect 68 1170 102 1177
rect 68 1096 102 1107
rect 68 1022 102 1037
rect 68 948 102 967
rect 68 874 102 897
rect 68 800 102 827
rect 68 726 102 757
rect 68 652 102 687
rect 68 581 102 617
rect 68 511 102 544
rect 68 441 102 470
rect 68 371 102 396
rect 68 301 102 321
rect 254 2607 278 2641
rect 312 2607 351 2641
rect 390 2607 423 2641
rect 466 2607 495 2641
rect 542 2607 567 2641
rect 618 2607 660 2641
rect 694 2607 701 2641
rect 735 2607 736 2641
rect 770 2617 872 2641
rect 770 2607 838 2617
rect 254 2547 288 2607
rect 838 2547 872 2583
rect 254 2478 288 2503
rect 254 2409 288 2430
rect 254 2340 288 2356
rect 254 2271 288 2282
rect 254 2202 288 2208
rect 254 2132 288 2134
rect 254 2094 288 2098
rect 254 2020 288 2028
rect 254 1946 288 1958
rect 254 1872 288 1888
rect 254 1798 288 1818
rect 254 1724 288 1748
rect 254 1650 288 1678
rect 254 1576 288 1608
rect 254 1502 288 1538
rect 254 1432 288 1468
rect 254 1362 288 1394
rect 254 1292 288 1320
rect 254 1222 288 1246
rect 254 1152 288 1172
rect 254 1082 288 1098
rect 254 1012 288 1024
rect 254 942 288 950
rect 254 872 288 876
rect 254 836 288 838
rect 254 762 288 768
rect 254 688 288 698
rect 254 614 288 628
rect 254 540 288 558
rect 254 466 288 488
rect 254 392 288 418
rect 356 2463 390 2503
rect 356 2389 390 2429
rect 356 2315 390 2355
rect 356 2241 390 2281
rect 356 2167 390 2207
rect 356 2093 390 2133
rect 356 2019 390 2059
rect 356 1945 390 1985
rect 356 1871 390 1911
rect 356 1797 390 1837
rect 356 1723 390 1763
rect 356 1649 390 1689
rect 356 1575 390 1615
rect 546 2447 580 2489
rect 546 2371 580 2413
rect 546 2296 580 2337
rect 546 2221 580 2262
rect 546 2146 580 2187
rect 546 2071 580 2112
rect 546 1996 580 2037
rect 546 1921 580 1962
rect 546 1846 580 1887
rect 546 1771 580 1812
rect 546 1696 580 1737
rect 546 1621 580 1662
rect 737 2463 771 2503
rect 737 2389 771 2429
rect 737 2315 771 2355
rect 737 2241 771 2281
rect 737 2167 771 2207
rect 737 2093 771 2133
rect 737 2019 771 2059
rect 737 1945 771 1985
rect 737 1871 771 1911
rect 737 1797 771 1837
rect 737 1723 771 1763
rect 737 1649 771 1689
rect 737 1575 771 1615
rect 356 1501 390 1541
rect 472 1491 506 1511
rect 737 1501 771 1541
rect 356 1427 390 1467
rect 428 1457 444 1491
rect 478 1473 512 1491
rect 506 1457 512 1473
rect 546 1457 580 1491
rect 614 1457 648 1491
rect 682 1457 698 1491
rect 737 1427 771 1467
rect 356 1353 390 1393
rect 356 1279 390 1319
rect 356 1205 390 1245
rect 356 1131 390 1171
rect 356 1057 390 1097
rect 356 983 390 1023
rect 356 909 390 949
rect 356 835 390 875
rect 356 761 390 801
rect 356 687 390 727
rect 356 613 390 653
rect 356 539 390 579
rect 356 465 390 505
rect 546 1326 580 1368
rect 546 1250 580 1292
rect 546 1175 580 1216
rect 546 1100 580 1141
rect 546 1025 580 1066
rect 546 950 580 991
rect 546 875 580 916
rect 546 800 580 841
rect 546 725 580 766
rect 546 650 580 691
rect 546 575 580 616
rect 546 500 580 541
rect 737 1353 771 1393
rect 737 1279 771 1319
rect 737 1205 771 1245
rect 737 1131 771 1171
rect 737 1057 771 1097
rect 737 983 771 1023
rect 737 909 771 949
rect 737 835 771 875
rect 737 761 771 801
rect 737 687 771 727
rect 737 613 771 653
rect 737 539 771 579
rect 737 465 771 505
rect 356 390 390 431
rect 472 370 506 408
rect 737 390 771 431
rect 254 312 288 348
rect 433 336 449 370
rect 506 336 517 370
rect 551 336 585 370
rect 619 336 653 370
rect 687 336 703 370
rect 838 2477 872 2503
rect 838 2407 872 2430
rect 838 2337 872 2356
rect 838 2267 872 2282
rect 838 2197 872 2208
rect 838 2127 872 2134
rect 838 2057 872 2060
rect 838 2020 872 2023
rect 838 1946 872 1953
rect 838 1872 872 1883
rect 838 1798 872 1813
rect 838 1724 872 1743
rect 838 1650 872 1673
rect 838 1576 872 1603
rect 838 1502 872 1533
rect 838 1428 872 1463
rect 838 1357 872 1393
rect 838 1287 872 1320
rect 838 1217 872 1246
rect 838 1147 872 1172
rect 838 1077 872 1098
rect 838 1007 872 1024
rect 838 937 872 950
rect 838 867 872 876
rect 838 797 872 802
rect 838 762 872 763
rect 838 727 872 728
rect 838 688 872 693
rect 838 614 872 624
rect 838 540 872 555
rect 838 466 872 486
rect 838 392 872 417
rect 838 288 872 348
rect 288 278 356 288
rect 254 254 356 278
rect 394 254 432 288
rect 469 254 508 288
rect 544 254 584 288
rect 620 254 660 288
rect 696 254 736 288
rect 772 254 814 288
rect 848 254 872 288
rect 68 231 102 246
rect 68 101 102 171
rect 1024 101 1058 2794
rect 68 67 203 101
rect 237 67 277 101
rect 311 67 351 101
rect 385 67 425 101
rect 459 67 499 101
rect 533 67 573 101
rect 607 67 647 101
rect 681 67 721 101
rect 755 67 796 101
rect 830 67 871 101
rect 905 67 946 101
rect 980 67 1058 101
<< viali >>
rect 68 2690 102 2724
rect 68 2644 102 2650
rect 68 2616 102 2644
rect 68 2575 102 2576
rect 68 2542 102 2575
rect 68 2471 102 2502
rect 68 2468 102 2471
rect 68 2401 102 2428
rect 68 2394 102 2401
rect 68 2331 102 2354
rect 68 2320 102 2331
rect 68 2261 102 2280
rect 68 2246 102 2261
rect 68 2191 102 2206
rect 68 2172 102 2191
rect 68 2121 102 2132
rect 68 2098 102 2121
rect 68 2051 102 2058
rect 68 2024 102 2051
rect 68 1981 102 1984
rect 68 1950 102 1981
rect 68 1877 102 1910
rect 68 1876 102 1877
rect 68 1807 102 1836
rect 68 1802 102 1807
rect 68 1737 102 1762
rect 68 1728 102 1737
rect 68 1667 102 1688
rect 68 1654 102 1667
rect 68 1597 102 1614
rect 68 1580 102 1597
rect 68 1527 102 1540
rect 68 1506 102 1527
rect 68 1457 102 1466
rect 68 1432 102 1457
rect 68 1387 102 1392
rect 68 1358 102 1387
rect 68 1317 102 1318
rect 68 1284 102 1317
rect 68 1211 102 1244
rect 68 1210 102 1211
rect 68 1141 102 1170
rect 68 1136 102 1141
rect 68 1071 102 1096
rect 68 1062 102 1071
rect 68 1001 102 1022
rect 68 988 102 1001
rect 68 931 102 948
rect 68 914 102 931
rect 68 861 102 874
rect 68 840 102 861
rect 68 791 102 800
rect 68 766 102 791
rect 68 721 102 726
rect 68 692 102 721
rect 68 651 102 652
rect 68 618 102 651
rect 68 547 102 578
rect 68 544 102 547
rect 68 477 102 504
rect 68 470 102 477
rect 68 407 102 430
rect 68 396 102 407
rect 68 337 102 355
rect 68 321 102 337
rect 68 267 102 280
rect 68 246 102 267
rect 356 2607 385 2641
rect 385 2607 390 2641
rect 432 2607 457 2641
rect 457 2607 466 2641
rect 508 2607 529 2641
rect 529 2607 542 2641
rect 584 2607 601 2641
rect 601 2607 618 2641
rect 660 2607 694 2641
rect 736 2607 770 2641
rect 254 2513 288 2537
rect 254 2503 288 2513
rect 254 2444 288 2464
rect 254 2430 288 2444
rect 254 2375 288 2390
rect 254 2356 288 2375
rect 254 2306 288 2316
rect 254 2282 288 2306
rect 254 2237 288 2242
rect 254 2208 288 2237
rect 254 2134 288 2168
rect 254 2062 288 2094
rect 254 2060 288 2062
rect 254 1992 288 2020
rect 254 1986 288 1992
rect 254 1922 288 1946
rect 254 1912 288 1922
rect 254 1852 288 1872
rect 254 1838 288 1852
rect 254 1782 288 1798
rect 254 1764 288 1782
rect 254 1712 288 1724
rect 254 1690 288 1712
rect 254 1642 288 1650
rect 254 1616 288 1642
rect 254 1572 288 1576
rect 254 1542 288 1572
rect 254 1468 288 1502
rect 254 1398 288 1428
rect 254 1394 288 1398
rect 254 1328 288 1354
rect 254 1320 288 1328
rect 254 1258 288 1280
rect 254 1246 288 1258
rect 254 1188 288 1206
rect 254 1172 288 1188
rect 254 1118 288 1132
rect 254 1098 288 1118
rect 254 1048 288 1058
rect 254 1024 288 1048
rect 254 978 288 984
rect 254 950 288 978
rect 254 908 288 910
rect 254 876 288 908
rect 254 802 288 836
rect 254 732 288 762
rect 254 728 288 732
rect 254 662 288 688
rect 254 654 288 662
rect 254 592 288 614
rect 254 580 288 592
rect 254 522 288 540
rect 254 506 288 522
rect 254 452 288 466
rect 254 432 288 452
rect 254 382 288 392
rect 254 358 288 382
rect 356 2503 390 2537
rect 356 2429 390 2463
rect 356 2355 390 2389
rect 356 2281 390 2315
rect 356 2207 390 2241
rect 356 2133 390 2167
rect 356 2059 390 2093
rect 356 1985 390 2019
rect 356 1911 390 1945
rect 356 1837 390 1871
rect 356 1763 390 1797
rect 356 1689 390 1723
rect 356 1615 390 1649
rect 546 2489 580 2523
rect 546 2413 580 2447
rect 546 2337 580 2371
rect 546 2262 580 2296
rect 546 2187 580 2221
rect 546 2112 580 2146
rect 546 2037 580 2071
rect 546 1962 580 1996
rect 546 1887 580 1921
rect 546 1812 580 1846
rect 546 1737 580 1771
rect 546 1662 580 1696
rect 546 1587 580 1621
rect 737 2503 771 2537
rect 737 2429 771 2463
rect 737 2355 771 2389
rect 737 2281 771 2315
rect 737 2207 771 2241
rect 737 2133 771 2167
rect 737 2059 771 2093
rect 737 1985 771 2019
rect 737 1911 771 1945
rect 737 1837 771 1871
rect 737 1763 771 1797
rect 737 1689 771 1723
rect 737 1615 771 1649
rect 356 1541 390 1575
rect 356 1467 390 1501
rect 472 1511 506 1545
rect 737 1541 771 1575
rect 472 1457 478 1473
rect 478 1457 506 1473
rect 737 1467 771 1501
rect 472 1439 506 1457
rect 356 1393 390 1427
rect 356 1319 390 1353
rect 356 1245 390 1279
rect 356 1171 390 1205
rect 356 1097 390 1131
rect 356 1023 390 1057
rect 356 949 390 983
rect 356 875 390 909
rect 356 801 390 835
rect 356 727 390 761
rect 356 653 390 687
rect 356 579 390 613
rect 356 505 390 539
rect 546 1368 580 1402
rect 546 1292 580 1326
rect 546 1216 580 1250
rect 546 1141 580 1175
rect 546 1066 580 1100
rect 546 991 580 1025
rect 546 916 580 950
rect 546 841 580 875
rect 546 766 580 800
rect 546 691 580 725
rect 546 616 580 650
rect 546 541 580 575
rect 546 466 580 500
rect 737 1393 771 1427
rect 737 1319 771 1353
rect 737 1245 771 1279
rect 737 1171 771 1205
rect 737 1097 771 1131
rect 737 1023 771 1057
rect 737 949 771 983
rect 737 875 771 909
rect 737 801 771 835
rect 737 727 771 761
rect 737 653 771 687
rect 737 579 771 613
rect 737 505 771 539
rect 356 431 390 465
rect 356 356 390 390
rect 472 408 506 442
rect 737 431 771 465
rect 472 336 483 370
rect 483 336 506 370
rect 737 356 771 390
rect 838 2513 872 2537
rect 838 2503 872 2513
rect 838 2443 872 2464
rect 838 2430 872 2443
rect 838 2373 872 2390
rect 838 2356 872 2373
rect 838 2303 872 2316
rect 838 2282 872 2303
rect 838 2233 872 2242
rect 838 2208 872 2233
rect 838 2163 872 2168
rect 838 2134 872 2163
rect 838 2093 872 2094
rect 838 2060 872 2093
rect 838 1987 872 2020
rect 838 1986 872 1987
rect 838 1917 872 1946
rect 838 1912 872 1917
rect 838 1847 872 1872
rect 838 1838 872 1847
rect 838 1777 872 1798
rect 838 1764 872 1777
rect 838 1707 872 1724
rect 838 1690 872 1707
rect 838 1637 872 1650
rect 838 1616 872 1637
rect 838 1567 872 1576
rect 838 1542 872 1567
rect 838 1497 872 1502
rect 838 1468 872 1497
rect 838 1427 872 1428
rect 838 1394 872 1427
rect 838 1323 872 1354
rect 838 1320 872 1323
rect 838 1253 872 1280
rect 838 1246 872 1253
rect 838 1183 872 1206
rect 838 1172 872 1183
rect 838 1113 872 1132
rect 838 1098 872 1113
rect 838 1043 872 1058
rect 838 1024 872 1043
rect 838 973 872 984
rect 838 950 872 973
rect 838 903 872 910
rect 838 876 872 903
rect 838 833 872 836
rect 838 802 872 833
rect 838 728 872 762
rect 838 658 872 688
rect 838 654 872 658
rect 838 589 872 614
rect 838 580 872 589
rect 838 520 872 540
rect 838 506 872 520
rect 838 451 872 466
rect 838 432 872 451
rect 838 382 872 392
rect 838 358 872 382
rect 356 254 360 288
rect 360 254 390 288
rect 432 254 435 288
rect 435 254 466 288
rect 508 254 510 288
rect 510 254 542 288
rect 584 254 586 288
rect 586 254 618 288
rect 660 254 662 288
rect 662 254 694 288
rect 736 254 738 288
rect 738 254 770 288
rect 68 197 102 205
rect 68 171 102 197
<< metal1 >>
rect 62 2724 108 2834
rect 62 2690 68 2724
rect 102 2690 108 2724
rect 62 2650 108 2690
rect 62 2616 68 2650
rect 102 2616 108 2650
rect 62 2576 108 2616
rect 62 2542 68 2576
rect 102 2542 108 2576
rect 62 2502 108 2542
rect 62 2468 68 2502
rect 102 2468 108 2502
rect 62 2428 108 2468
rect 62 2394 68 2428
rect 102 2394 108 2428
rect 62 2354 108 2394
rect 62 2320 68 2354
rect 102 2320 108 2354
rect 62 2280 108 2320
rect 62 2246 68 2280
rect 102 2246 108 2280
rect 62 2206 108 2246
rect 62 2172 68 2206
rect 102 2172 108 2206
rect 62 2132 108 2172
rect 62 2098 68 2132
rect 102 2098 108 2132
rect 62 2058 108 2098
rect 62 2024 68 2058
rect 102 2024 108 2058
rect 62 1984 108 2024
rect 62 1950 68 1984
rect 102 1950 108 1984
rect 62 1910 108 1950
rect 62 1876 68 1910
rect 102 1876 108 1910
rect 62 1836 108 1876
rect 62 1802 68 1836
rect 102 1802 108 1836
rect 62 1762 108 1802
rect 62 1728 68 1762
rect 102 1728 108 1762
rect 62 1688 108 1728
rect 62 1654 68 1688
rect 102 1654 108 1688
rect 62 1614 108 1654
rect 62 1580 68 1614
rect 102 1580 108 1614
rect 62 1540 108 1580
rect 62 1506 68 1540
rect 102 1506 108 1540
rect 62 1466 108 1506
rect 62 1432 68 1466
rect 102 1432 108 1466
rect 62 1392 108 1432
rect 62 1358 68 1392
rect 102 1358 108 1392
rect 62 1318 108 1358
rect 62 1284 68 1318
rect 102 1284 108 1318
rect 62 1244 108 1284
rect 62 1210 68 1244
rect 102 1210 108 1244
rect 62 1170 108 1210
rect 62 1136 68 1170
rect 102 1136 108 1170
rect 62 1096 108 1136
rect 62 1062 68 1096
rect 102 1062 108 1096
rect 62 1022 108 1062
rect 62 988 68 1022
rect 102 988 108 1022
rect 62 948 108 988
rect 62 914 68 948
rect 102 914 108 948
rect 62 874 108 914
rect 62 840 68 874
rect 102 840 108 874
rect 62 800 108 840
rect 62 766 68 800
rect 102 766 108 800
rect 62 726 108 766
rect 62 692 68 726
rect 102 692 108 726
rect 62 652 108 692
rect 62 618 68 652
rect 102 618 108 652
rect 62 578 108 618
rect 62 544 68 578
rect 102 544 108 578
rect 62 504 108 544
rect 62 470 68 504
rect 102 470 108 504
rect 62 430 108 470
rect 62 396 68 430
rect 102 396 108 430
rect 62 355 108 396
rect 62 321 68 355
rect 102 321 108 355
rect 62 280 108 321
rect 62 246 68 280
rect 102 246 108 280
rect 248 2641 878 2647
rect 248 2607 356 2641
rect 390 2607 432 2641
rect 466 2607 508 2641
rect 542 2607 584 2641
rect 618 2607 660 2641
rect 694 2607 736 2641
rect 770 2607 878 2641
rect 248 2601 878 2607
rect 248 2537 396 2601
tri 396 2565 432 2601 nw
tri 695 2565 731 2601 ne
rect 248 2503 254 2537
rect 288 2503 356 2537
rect 390 2503 396 2537
rect 731 2537 878 2601
rect 248 2464 396 2503
rect 248 2430 254 2464
rect 288 2463 396 2464
rect 288 2430 356 2463
rect 248 2429 356 2430
rect 390 2429 396 2463
rect 248 2390 396 2429
rect 248 2356 254 2390
rect 288 2389 396 2390
rect 288 2356 356 2389
rect 248 2355 356 2356
rect 390 2355 396 2389
rect 248 2316 396 2355
rect 248 2282 254 2316
rect 288 2315 396 2316
rect 288 2282 356 2315
rect 248 2281 356 2282
rect 390 2281 396 2315
rect 248 2242 396 2281
rect 248 2208 254 2242
rect 288 2241 396 2242
rect 288 2208 356 2241
rect 248 2207 356 2208
rect 390 2207 396 2241
rect 248 2168 396 2207
rect 248 2134 254 2168
rect 288 2167 396 2168
rect 288 2134 356 2167
rect 248 2133 356 2134
rect 390 2133 396 2167
rect 248 2094 396 2133
rect 248 2060 254 2094
rect 288 2093 396 2094
rect 288 2060 356 2093
rect 248 2059 356 2060
rect 390 2059 396 2093
rect 248 2020 396 2059
rect 248 1986 254 2020
rect 288 2019 396 2020
rect 288 1986 356 2019
rect 248 1985 356 1986
rect 390 1985 396 2019
rect 248 1946 396 1985
rect 248 1912 254 1946
rect 288 1945 396 1946
rect 288 1912 356 1945
rect 248 1911 356 1912
rect 390 1911 396 1945
rect 248 1872 396 1911
rect 248 1838 254 1872
rect 288 1871 396 1872
rect 288 1838 356 1871
rect 248 1837 356 1838
rect 390 1837 396 1871
rect 248 1798 396 1837
rect 248 1764 254 1798
rect 288 1797 396 1798
rect 288 1764 356 1797
rect 248 1763 356 1764
rect 390 1763 396 1797
rect 248 1724 396 1763
rect 248 1690 254 1724
rect 288 1723 396 1724
rect 288 1690 356 1723
rect 248 1689 356 1690
rect 390 1689 396 1723
rect 248 1650 396 1689
rect 248 1616 254 1650
rect 288 1649 396 1650
rect 288 1616 356 1649
rect 248 1615 356 1616
rect 390 1615 396 1649
rect 248 1576 396 1615
rect 248 1542 254 1576
rect 288 1575 396 1576
rect 288 1542 356 1575
rect 248 1541 356 1542
rect 390 1541 396 1575
rect 248 1502 396 1541
rect 248 1468 254 1502
rect 288 1501 396 1502
rect 288 1468 356 1501
rect 248 1467 356 1468
rect 390 1467 396 1501
rect 248 1428 396 1467
rect 248 1394 254 1428
rect 288 1427 396 1428
rect 288 1394 356 1427
rect 248 1393 356 1394
rect 390 1393 396 1427
rect 248 1354 396 1393
rect 248 1320 254 1354
rect 288 1353 396 1354
rect 288 1320 356 1353
rect 248 1319 356 1320
rect 390 1319 396 1353
rect 248 1280 396 1319
rect 248 1246 254 1280
rect 288 1279 396 1280
rect 288 1246 356 1279
rect 248 1245 356 1246
rect 390 1245 396 1279
rect 248 1206 396 1245
rect 248 1172 254 1206
rect 288 1205 396 1206
rect 288 1172 356 1205
rect 248 1171 356 1172
rect 390 1171 396 1205
rect 248 1132 396 1171
rect 248 1098 254 1132
rect 288 1131 396 1132
rect 288 1098 356 1131
rect 248 1097 356 1098
rect 390 1097 396 1131
rect 248 1058 396 1097
rect 248 1024 254 1058
rect 288 1057 396 1058
rect 288 1024 356 1057
rect 248 1023 356 1024
rect 390 1023 396 1057
rect 248 984 396 1023
rect 248 950 254 984
rect 288 983 396 984
rect 288 950 356 983
rect 248 949 356 950
rect 390 949 396 983
rect 248 910 396 949
rect 248 876 254 910
rect 288 909 396 910
rect 288 876 356 909
rect 248 875 356 876
rect 390 875 396 909
rect 248 836 396 875
rect 248 802 254 836
rect 288 835 396 836
rect 288 802 356 835
rect 248 801 356 802
rect 390 801 396 835
rect 248 762 396 801
rect 248 728 254 762
rect 288 761 396 762
rect 288 728 356 761
rect 248 727 356 728
rect 390 727 396 761
rect 248 688 396 727
rect 248 654 254 688
rect 288 687 396 688
rect 288 654 356 687
rect 248 653 356 654
rect 390 653 396 687
rect 248 614 396 653
rect 248 580 254 614
rect 288 613 396 614
rect 288 580 356 613
rect 248 579 356 580
rect 390 579 396 613
rect 248 540 396 579
rect 248 506 254 540
rect 288 539 396 540
rect 288 506 356 539
rect 248 505 356 506
rect 390 505 396 539
rect 248 466 396 505
rect 248 432 254 466
rect 288 465 396 466
rect 288 432 356 465
rect 248 431 356 432
rect 390 431 396 465
rect 248 392 396 431
rect 248 358 254 392
rect 288 390 396 392
rect 288 358 356 390
rect 248 356 356 358
rect 390 356 396 390
rect 248 324 396 356
rect 466 1545 512 2528
rect 466 1511 472 1545
rect 506 1511 512 1545
rect 466 1473 512 1511
rect 466 1439 472 1473
rect 506 1439 512 1473
rect 466 442 512 1439
rect 540 2523 586 2535
rect 540 2489 546 2523
rect 580 2489 586 2523
rect 540 2447 586 2489
rect 540 2413 546 2447
rect 580 2413 586 2447
rect 540 2371 586 2413
rect 540 2337 546 2371
rect 580 2337 586 2371
rect 540 2296 586 2337
rect 540 2262 546 2296
rect 580 2262 586 2296
rect 540 2221 586 2262
rect 540 2187 546 2221
rect 580 2187 586 2221
rect 540 2146 586 2187
rect 540 2112 546 2146
rect 580 2112 586 2146
rect 540 2071 586 2112
rect 540 2037 546 2071
rect 580 2037 586 2071
rect 540 1996 586 2037
rect 540 1962 546 1996
rect 580 1962 586 1996
rect 540 1921 586 1962
rect 540 1887 546 1921
rect 580 1887 586 1921
rect 540 1846 586 1887
rect 540 1812 546 1846
rect 580 1812 586 1846
rect 540 1771 586 1812
rect 540 1737 546 1771
rect 580 1737 586 1771
rect 540 1696 586 1737
rect 540 1662 546 1696
rect 580 1662 586 1696
rect 540 1621 586 1662
rect 540 1587 546 1621
rect 580 1587 586 1621
rect 540 1402 586 1587
rect 540 1368 546 1402
rect 580 1368 586 1402
rect 540 1326 586 1368
rect 540 1292 546 1326
rect 580 1292 586 1326
rect 540 1250 586 1292
rect 540 1216 546 1250
rect 580 1216 586 1250
rect 540 1175 586 1216
rect 540 1141 546 1175
rect 580 1141 586 1175
rect 540 1100 586 1141
rect 540 1066 546 1100
rect 580 1066 586 1100
rect 540 1025 586 1066
rect 540 991 546 1025
rect 580 991 586 1025
rect 540 950 586 991
rect 540 916 546 950
rect 580 916 586 950
rect 540 875 586 916
rect 540 841 546 875
rect 580 841 586 875
rect 540 800 586 841
rect 540 766 546 800
rect 580 766 586 800
rect 540 725 586 766
rect 540 691 546 725
rect 580 691 586 725
rect 540 650 586 691
rect 540 616 546 650
rect 580 616 586 650
rect 540 575 586 616
rect 540 541 546 575
rect 580 541 586 575
rect 540 500 586 541
rect 540 466 546 500
rect 580 466 586 500
rect 540 454 586 466
rect 731 2503 737 2537
rect 771 2503 838 2537
rect 872 2503 878 2537
rect 731 2464 878 2503
rect 731 2463 838 2464
rect 731 2429 737 2463
rect 771 2430 838 2463
rect 872 2430 878 2464
rect 771 2429 878 2430
rect 731 2390 878 2429
rect 731 2389 838 2390
rect 731 2355 737 2389
rect 771 2356 838 2389
rect 872 2356 878 2390
rect 771 2355 878 2356
rect 731 2316 878 2355
rect 731 2315 838 2316
rect 731 2281 737 2315
rect 771 2282 838 2315
rect 872 2282 878 2316
rect 771 2281 878 2282
rect 731 2242 878 2281
rect 731 2241 838 2242
rect 731 2207 737 2241
rect 771 2208 838 2241
rect 872 2208 878 2242
rect 771 2207 878 2208
rect 731 2168 878 2207
rect 731 2167 838 2168
rect 731 2133 737 2167
rect 771 2134 838 2167
rect 872 2134 878 2168
rect 771 2133 878 2134
rect 731 2094 878 2133
rect 731 2093 838 2094
rect 731 2059 737 2093
rect 771 2060 838 2093
rect 872 2060 878 2094
rect 771 2059 878 2060
rect 731 2020 878 2059
rect 731 2019 838 2020
rect 731 1985 737 2019
rect 771 1986 838 2019
rect 872 1986 878 2020
rect 771 1985 878 1986
rect 731 1946 878 1985
rect 731 1945 838 1946
rect 731 1911 737 1945
rect 771 1912 838 1945
rect 872 1912 878 1946
rect 771 1911 878 1912
rect 731 1872 878 1911
rect 731 1871 838 1872
rect 731 1837 737 1871
rect 771 1838 838 1871
rect 872 1838 878 1872
rect 771 1837 878 1838
rect 731 1798 878 1837
rect 731 1797 838 1798
rect 731 1763 737 1797
rect 771 1764 838 1797
rect 872 1764 878 1798
rect 771 1763 878 1764
rect 731 1724 878 1763
rect 731 1723 838 1724
rect 731 1689 737 1723
rect 771 1690 838 1723
rect 872 1690 878 1724
rect 771 1689 878 1690
rect 731 1650 878 1689
rect 731 1649 838 1650
rect 731 1615 737 1649
rect 771 1616 838 1649
rect 872 1616 878 1650
rect 771 1615 878 1616
rect 731 1576 878 1615
rect 731 1575 838 1576
rect 731 1541 737 1575
rect 771 1542 838 1575
rect 872 1542 878 1576
rect 771 1541 878 1542
rect 731 1502 878 1541
rect 731 1501 838 1502
rect 731 1467 737 1501
rect 771 1468 838 1501
rect 872 1468 878 1502
rect 771 1467 878 1468
rect 731 1428 878 1467
rect 731 1427 838 1428
rect 731 1393 737 1427
rect 771 1394 838 1427
rect 872 1394 878 1428
rect 771 1393 878 1394
rect 731 1354 878 1393
rect 731 1353 838 1354
rect 731 1319 737 1353
rect 771 1320 838 1353
rect 872 1320 878 1354
rect 771 1319 878 1320
rect 731 1280 878 1319
rect 731 1279 838 1280
rect 731 1245 737 1279
rect 771 1246 838 1279
rect 872 1246 878 1280
rect 771 1245 878 1246
rect 731 1206 878 1245
rect 731 1205 838 1206
rect 731 1171 737 1205
rect 771 1172 838 1205
rect 872 1172 878 1206
rect 771 1171 878 1172
rect 731 1132 878 1171
rect 731 1131 838 1132
rect 731 1097 737 1131
rect 771 1098 838 1131
rect 872 1098 878 1132
rect 771 1097 878 1098
rect 731 1058 878 1097
rect 731 1057 838 1058
rect 731 1023 737 1057
rect 771 1024 838 1057
rect 872 1024 878 1058
rect 771 1023 878 1024
rect 731 984 878 1023
rect 731 983 838 984
rect 731 949 737 983
rect 771 950 838 983
rect 872 950 878 984
rect 771 949 878 950
rect 731 910 878 949
rect 731 909 838 910
rect 731 875 737 909
rect 771 876 838 909
rect 872 876 878 910
rect 771 875 878 876
rect 731 836 878 875
rect 731 835 838 836
rect 731 801 737 835
rect 771 802 838 835
rect 872 802 878 836
rect 771 801 878 802
rect 731 762 878 801
rect 731 761 838 762
rect 731 727 737 761
rect 771 728 838 761
rect 872 728 878 762
rect 771 727 878 728
rect 731 688 878 727
rect 731 687 838 688
rect 731 653 737 687
rect 771 654 838 687
rect 872 654 878 688
rect 771 653 878 654
rect 731 614 878 653
rect 731 613 838 614
rect 731 579 737 613
rect 771 580 838 613
rect 872 580 878 614
rect 771 579 878 580
rect 731 540 878 579
rect 731 539 838 540
rect 731 505 737 539
rect 771 506 838 539
rect 872 506 878 540
rect 771 505 878 506
rect 731 466 878 505
rect 731 465 838 466
rect 466 408 472 442
rect 506 408 512 442
rect 466 370 512 408
rect 466 336 472 370
rect 506 336 512 370
tri 396 324 402 330 sw
rect 466 324 512 336
rect 731 431 737 465
rect 771 432 838 465
rect 872 432 878 466
rect 771 431 878 432
rect 731 392 878 431
rect 731 390 838 392
rect 731 356 737 390
rect 771 358 838 390
rect 872 358 878 392
rect 771 356 878 358
tri 725 324 731 330 se
rect 731 324 878 356
rect 248 294 402 324
tri 402 294 432 324 sw
tri 695 294 725 324 se
rect 725 294 878 324
rect 248 288 878 294
rect 248 254 356 288
rect 390 254 432 288
rect 466 254 508 288
rect 542 254 584 288
rect 618 254 660 288
rect 694 254 736 288
rect 770 254 878 288
rect 248 248 878 254
rect 62 205 108 246
rect 62 171 68 205
rect 102 171 108 205
rect 62 159 108 171
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 506 1 0 336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 506 1 0 1439
box 0 0 1 1
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_0
timestamp 1707688321
transform 1 0 415 0 -1 2533
box -79 -26 375 1026
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_1
timestamp 1707688321
transform 1 0 415 0 -1 1412
box -79 -26 375 1026
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 1 428 1 0 1441
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1707688321
transform 0 1 433 1 0 320
box 0 0 1 1
<< labels >>
flabel metal1 s 775 2504 830 2532 7 FreeSans 200 90 0 0 vgnd_io
port 1 nsew
flabel metal1 s 466 2496 512 2528 7 FreeSans 200 90 0 0 pd_h
port 3 nsew
flabel metal1 s 293 2504 348 2532 7 FreeSans 200 90 0 0 vgnd_io
port 1 nsew
flabel metal1 s 74 2799 96 2816 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
<< properties >>
string GDS_END 92015758
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91990352
string path 2.125 3.675 2.125 68.200 
<< end >>
