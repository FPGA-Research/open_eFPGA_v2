magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 112 226
<< nmos >>
rect 0 0 36 200
<< ndiff >>
rect -50 0 0 200
rect 36 0 86 200
<< poly >>
rect 0 200 36 226
rect 0 -26 36 0
<< metal1 >>
rect -51 -16 -5 186
rect 41 -16 87 186
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1707688321
transform 1 0 36 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 64 85 64 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86869862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86869036
<< end >>
