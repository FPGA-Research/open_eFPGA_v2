##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 17:26:08 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO LUT4AB
  CLASS BLOCK ;
  SIZE 210.2200 BY 219.6400 ;
  FOREIGN LUT4AB 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 219.3100 14.1150 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.04805 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.233 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 27.697 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 138.411 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 219.3100 12.7350 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.4864 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 97.3175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.737 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 219.3100 11.3550 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3744 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.7945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 219.3100 10.4350 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.7328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.712 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 219.3100 25.1550 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.9965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.1516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.416 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 219.3100 23.7750 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.7258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.008 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 219.3100 22.3950 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.9136 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 219.3100 21.0150 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.4708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 219.3100 19.6350 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 219.3100 18.2550 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.991 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.027 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 219.3100 16.8750 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.16365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.369 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.3764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 101.805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.152 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 219.3100 15.4950 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.5756 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 219.3100 35.7350 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.3978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.592 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 219.3100 34.3550 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.691 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 192.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 219.3100 33.4350 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.0755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.1035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 219.3100 32.0550 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.86 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.064 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 219.3100 30.6750 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7998 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.2632 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.198 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 219.3100 29.2950 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.867 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.7234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 219.3100 27.9150 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 219.3100 26.5350 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 219.3100 57.3550 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6268 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8368 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.066 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 219.3100 56.4350 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.4928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.3865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.3428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 219.3100 55.0550 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.6057 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.408 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 219.3100 53.6750 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4297 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.5178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 219.3100 52.2950 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.60605 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.713 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.402 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.7156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.46 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 219.3100 50.9150 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.4308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 274.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 219.3100 49.5350 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.9674 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.904 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 219.3100 48.1550 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 219.3100 46.7750 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2386 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.075 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 219.3100 45.3950 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.962 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 219.3100 44.0150 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.6936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.64 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 219.3100 42.6350 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 219.3100 41.2550 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.672 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.2825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.6976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 303.328 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 219.3100 39.8750 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 219.3100 38.4950 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8853 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.5874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.896 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 219.3100 37.1150 219.6400 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.264 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 219.3100 79.4350 219.6400 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.281 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9352 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.0768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.88 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 219.3100 78.0550 219.6400 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.9166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 219.3100 76.6750 219.6400 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9155 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.1826 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 219.3100 75.2950 219.6400 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.401 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 219.3100 73.9150 219.6400 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.8112 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 58.9785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 219.3100 72.5350 219.6400 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1685 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.711 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.2478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 219.3100 71.1550 219.6400 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0425 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.192 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 219.3100 69.7750 219.6400 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.127 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 219.3100 68.3950 219.6400 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.8745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.292 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 219.3100 67.0150 219.6400 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.1505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9792 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.778 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 219.3100 65.6350 219.6400 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9624 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 278.544 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 219.3100 64.2550 219.6400 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 21.5342 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 107.597 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 219.3100 62.8750 219.6400 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.5528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 280.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 219.3100 61.4950 219.6400 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.6428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 169.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 219.3100 60.1150 219.6400 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51045 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.777 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.6365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 219.3100 58.7350 219.6400 ;
    END
  END NN4BEG[0]
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.581 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.3736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 177.2600 219.1550 177.4000 219.6400 ;
    END
  END Co
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.4656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.9975 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0675 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4529 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.431 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 0.0000 14.1150 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.4976 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.3405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 110.415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.8876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.008 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 0.0000 12.7350 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.07 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.0532 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 0.0000 11.3550 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.8688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 245.104 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.0277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.3825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4635 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.6269 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 13.4821 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 65.0263 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 0.0000 25.1550 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.6896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 38.3705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.062 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4549 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.2909 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 0.0000 23.7750 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.7272 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 117.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 41.506 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 221.425 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 0.0000 22.3950 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.1371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.9092 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 211.169 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 0.0000 21.0150 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.3533 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.5955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7488 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.5447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.704 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 8.61845 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 44.2936 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 0.0000 19.6350 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.136 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8292 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.5347 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.345 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.64 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 29.7215 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 150.922 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.8985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.1 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 0.0000 18.2550 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22145 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.437 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.5612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.4084 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 22.3484 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.853 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 0.0000 16.8750 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.4871 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.923 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.70425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.0003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.8305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1376 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.4627 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.6 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 0.0000 35.7350 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.9935 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 79.7965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.8273 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 0.0000 34.3550 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.587 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.336 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 0.0000 33.4350 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.0688 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.2665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 0.0000 32.0550 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9249 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.7116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 0.0000 30.6750 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.178 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.6482 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.672 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 0.0000 29.2950 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.3147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.1936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.64 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 0.0000 27.9150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.4964 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 0.0000 26.5350 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.00148 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.6128 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 0.0000 57.3550 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.33 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 368.921 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.594 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.4116 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.6633 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 0.0000 55.0550 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.47005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.553 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.6044 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.9445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.688 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.62855 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.7481 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 0.0000 53.6750 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.1018 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.68 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.6563 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1624 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.6975 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5455 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.4548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 67.2061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 357.788 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 0.0000 50.9150 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.0714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.9972 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 374.216 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 0.0000 49.5350 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 17.9884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 89.8275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.03 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.6435 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.9138 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 0.0000 48.1550 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.7275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.5398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.4562 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 0.0000 46.7750 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.9475 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10869 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.9899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 0.0000 45.3950 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.1608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.3848 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.037 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 0.0000 44.0150 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 20.7576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 103.674 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.454 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.152 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.83246 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.7677 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 0.0000 42.6350 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.5644 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.088 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 0.0000 41.2550 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.602 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.3478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 191.344 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 0.0000 39.8750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.193 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.885 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 0.0000 38.4950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.9447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.8672 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.84 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 0.0000 37.1150 0.3300 ;
    END
  END N4END[0]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.0092 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 87.2604 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 465.226 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 0.0000 79.4350 0.3300 ;
    END
  END NN4END[15]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.7916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.4726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 73.5896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 394.499 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 0.0000 78.0550 0.3300 ;
    END
  END NN4END[14]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.942 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.5823 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.5232 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 0.0000 76.6750 0.3300 ;
    END
  END NN4END[13]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.06845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 19.829 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 99.071 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 27.002 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 133.779 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.0389226 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 0.0000 75.2950 0.3300 ;
    END
  END NN4END[12]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9911 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.3888 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 37.0986 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.798 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 0.0000 73.9150 0.3300 ;
    END
  END NN4END[11]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.1124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 75.4845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 49.7358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8881 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.713 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END NN4END[10]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.2174 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 279.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.666 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 430.543 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END NN4END[9]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.9656 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.7135 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.116 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.83973 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.804 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 0.0000 69.7750 0.3300 ;
    END
  END NN4END[8]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.7102 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 78.4735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.582 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.792 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.82155 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.7131 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 0.0000 68.3950 0.3300 ;
    END
  END NN4END[7]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.61811 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.6525 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END NN4END[6]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.9975 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.32525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.2316 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 0.0000 65.6350 0.3300 ;
    END
  END NN4END[5]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5148 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4595 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.5728 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.707 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 0.0000 64.2550 0.3300 ;
    END
  END NN4END[4]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.9955 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END NN4END[3]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.5786 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 0.0000 61.4950 0.3300 ;
    END
  END NN4END[2]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.161 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.544 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 0.0000 60.1150 0.3300 ;
    END
  END NN4END[1]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7671 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.8538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 213.024 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 0.0000 58.7350 0.3300 ;
    END
  END NN4END[0]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.069 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.184 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3735 LAYER met4  ;
    ANTENNAMAXAREACAR 45.712 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.999 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.800698 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 177.2600 0.0000 177.4000 0.4850 ;
    END
  END Ci
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.693 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.536 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 84.7600 210.2200 84.9000 ;
    END
  END E1BEG[3]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.534 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.976 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 83.4000 210.2200 83.5400 ;
    END
  END E1BEG[2]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 81.7000 210.2200 81.8400 ;
    END
  END E1BEG[1]
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 80.3400 210.2200 80.4800 ;
    END
  END E1BEG[0]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.757 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 65.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 96.6600 210.2200 96.8000 ;
    END
  END E2BEG[7]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3085 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.371 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.887 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.416 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 94.9600 210.2200 95.1000 ;
    END
  END E2BEG[6]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 45.0621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 241.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 93.6000 210.2200 93.7400 ;
    END
  END E2BEG[5]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.7648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 92.2400 210.2200 92.3800 ;
    END
  END E2BEG[4]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 90.5400 210.2200 90.6800 ;
    END
  END E2BEG[3]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.985 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 89.1800 210.2200 89.3200 ;
    END
  END E2BEG[2]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 87.8200 210.2200 87.9600 ;
    END
  END E2BEG[1]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 86.1200 210.2200 86.2600 ;
    END
  END E2BEG[0]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.009 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.8316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 108.2200 210.2200 108.3600 ;
    END
  END E2BEGb[7]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.9154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 106.8600 210.2200 107.0000 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.034 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 105.5000 210.2200 105.6400 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3921 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.8248 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 103.8000 210.2200 103.9400 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.631 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.6298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 48.848 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 102.4400 210.2200 102.5800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 26.146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 101.0800 210.2200 101.2200 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 99.3800 210.2200 99.5200 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.546 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.569 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.257 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.4928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 136.432 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 98.0200 210.2200 98.1600 ;
    END
  END E2BEGb[0]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 24.658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 131.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 132.0200 210.2200 132.1600 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8834 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.256 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 44.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 237.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 130.3200 210.2200 130.4600 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.4148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.016 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 128.9600 210.2200 129.1000 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.817 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.5258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.608 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 127.6000 210.2200 127.7400 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 125.9000 210.2200 126.0400 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5647 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 124.5400 210.2200 124.6800 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.842 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.7926 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 85.168 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 123.1800 210.2200 123.3200 ;
    END
  END EE4BEG[9]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.144 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 121.4800 210.2200 121.6200 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.9376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.636 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 120.1200 210.2200 120.2600 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.101 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.6532 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 118.7600 210.2200 118.9000 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.789 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.3156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 117.0600 210.2200 117.2000 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.036 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 115.7000 210.2200 115.8400 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 114.3400 210.2200 114.4800 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.0968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.258 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 112.6400 210.2200 112.7800 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 111.2800 210.2200 111.4200 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 109.9200 210.2200 110.0600 ;
    END
  END EE4BEG[0]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.9496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 149.7000 210.2200 149.8400 ;
    END
  END E6BEG[11]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.279 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 247.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.9548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 148.0000 210.2200 148.1400 ;
    END
  END E6BEG[10]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.4652 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.1 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 146.6400 210.2200 146.7800 ;
    END
  END E6BEG[9]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.582 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 145.2800 210.2200 145.4200 ;
    END
  END E6BEG[8]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.276 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 143.5800 210.2200 143.7200 ;
    END
  END E6BEG[7]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.4895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 142.2200 210.2200 142.3600 ;
    END
  END E6BEG[6]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 140.8600 210.2200 141.0000 ;
    END
  END E6BEG[5]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 139.1600 210.2200 139.3000 ;
    END
  END E6BEG[4]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 137.8000 210.2200 137.9400 ;
    END
  END E6BEG[3]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.245 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.367 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.2386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.88 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 136.4400 210.2200 136.5800 ;
    END
  END E6BEG[2]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 134.7400 210.2200 134.8800 ;
    END
  END E6BEG[1]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 133.3800 210.2200 133.5200 ;
    END
  END E6BEG[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.6956 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.3044 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.3393 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 84.7600 0.4850 84.9000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1795 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.8828 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 43.2853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.0736 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 83.4000 0.4850 83.5400 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.5128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 81.7000 0.4850 81.8400 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7046 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.136 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3212 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5935 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.6992 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 80.3400 0.4850 80.4800 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2499 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.851 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.4656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 115.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.0092 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 309.488 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 96.6600 0.4850 96.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.003 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 17.9572 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.402 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 94.9600 0.4850 95.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.344 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.8966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 61.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4829 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 194.245 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 93.6000 0.4850 93.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4525 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.71488 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.1038 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.024 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 31.0971 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.327 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 92.2400 0.4850 92.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2979 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10754 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.4357 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.9828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.712 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.4716 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 51.6774 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 90.5400 0.4850 90.6800 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.73731 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.936 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.8496 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 117.472 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 35.1644 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 184.147 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.153401 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 89.1800 0.4850 89.3200 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.0294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.568 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.9992 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 334.197 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 87.8200 0.4850 87.9600 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6467 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.298 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 86.1200 0.4850 86.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 85.0885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.0869 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.954 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.704 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 108.2200 0.4850 108.3600 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1448 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.9704 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.358 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 106.8600 0.4850 107.0000 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1448 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.2782 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 142.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 105.5000 0.4850 105.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 103.8000 0.4850 103.9400 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4835 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3284 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 102.4400 0.4850 102.5800 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.2898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 199.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.332 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.4726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 46.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 101.0800 0.4850 101.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 39.8158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 99.3800 0.4850 99.5200 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.5685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.9865 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 98.0200 0.4850 98.1600 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 40.234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 215.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.3404 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 35.2968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 188.861 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 132.0200 0.4850 132.1600 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.14182 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 24.169 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 130.3200 0.4850 130.4600 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.92101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 27.1805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 128.9600 0.4850 129.1000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 84.175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9092 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 117.151 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 127.6000 0.4850 127.7400 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.48269 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.9825 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 125.9000 0.4850 126.0400 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.81024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 12.6202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 124.5400 0.4850 124.6800 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.75865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.3623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 123.1800 0.4850 123.3200 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.0168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.444 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 228.649 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 121.4800 0.4850 121.6200 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0713 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.0775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.122 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 267.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 9.24673 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 47.1663 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 120.1200 0.4850 120.2600 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.75 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.397 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 143.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.4793 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.4 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 118.7600 0.4850 118.9000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.219 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.9224 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.664 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8815 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 371.362 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 117.0600 0.4850 117.2000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3549 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.3734 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 21.8641 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.567 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 115.7000 0.4850 115.8400 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.9588 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.5576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 114.3400 0.4850 114.4800 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.4395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 112.6400 0.4850 112.7800 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.3048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.3572 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.12 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 111.2800 0.4850 111.4200 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.688 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.9338 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 109.9200 0.4850 110.0600 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.193 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.048 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1011 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.572 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 149.7000 0.4850 149.8400 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.3017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 86.2295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.098 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 12.5616 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.27 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 148.0000 0.4850 148.1400 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2506 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.092 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.629 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.6936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 31.6729 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 170.768 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 146.6400 0.4850 146.7800 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.136 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 68.5738 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.611 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 145.2800 0.4850 145.4200 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.1274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 157.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.3994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 43.6704 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 233.529 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 143.5800 0.4850 143.7200 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.6604 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 159.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.8274 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.912 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 142.2200 0.4850 142.3600 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.3714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.392 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.6929 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.589 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 140.8600 0.4850 141.0000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.48646 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.0013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 139.1600 0.4850 139.3000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.3864 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 250.675 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 137.8000 0.4850 137.9400 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.8914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.832 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.4807 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 136.4400 0.4850 136.5800 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.2644 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0164 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 134.7400 0.4850 134.8800 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.903 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 106.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.8594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 133.3800 0.4850 133.5200 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.0148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.216 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 0.0000 84.4950 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3687 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.3204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 0.0000 83.1150 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8147 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.9884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.016 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 0.0000 81.7350 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.496 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 0.0000 80.3550 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.1925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.9576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 182.048 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 0.0000 106.1150 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.2012 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.288 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 0.0000 104.7350 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.5714 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 0.0000 103.3550 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.76545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.077 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.9974 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.064 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 0.0000 102.4350 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.5124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.144 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 0.0000 101.0550 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.864 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 0.0000 99.6750 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0894 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 0.0000 98.2950 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.1948 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.8827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 0.0000 96.9150 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 0.0000 95.5350 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 0.0000 94.1550 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.9996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 0.0000 92.7750 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.5928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 0.0000 91.3950 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.33705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.573 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.1368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.6065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.9944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.854 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 0.0000 90.0150 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.1268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.48 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 0.0000 88.6350 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.71 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.4725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.0918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.96 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 0.0000 87.2550 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 0.0000 85.8750 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 13.2237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 65.5935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.2708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.248 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 0.0000 127.7350 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.70425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.4456 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 0.0000 126.3550 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.256 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.8132 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 0.0000 125.4350 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8495 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3859 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.5268 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 243.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 0.0000 124.0550 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.9014 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 315.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 0.0000 122.6750 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2771 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.4232 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 297.472 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 0.0000 121.2950 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.8116 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 53.9805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.796 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 0.0000 119.9150 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 0.0000 118.5350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0628 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 0.0000 117.1550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.5132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.4885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 0.0000 115.7750 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 48.8112 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 262.208 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 0.0000 114.3950 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.0288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.748 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 0.0000 113.0150 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.818 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 0.0000 111.6350 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.188 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 0.0000 110.2550 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 65.1444 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 351.2 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 0.0000 108.8750 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.305 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.76 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.1596 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 289.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 0.0000 107.4950 0.3300 ;
    END
  END S4BEG[0]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.8662 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 193.168 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 0.0000 149.3550 0.3300 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5145 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.0458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.048 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 0.0000 148.4350 0.3300 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.2378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.072 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 0.0000 147.0550 0.3300 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.8984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.536 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 0.0000 145.6750 0.3300 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.2622 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 275.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 0.0000 144.2950 0.3300 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4148 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.9965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7524 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.526 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 0.0000 142.9150 0.3300 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.5678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 296.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 0.0000 141.5350 0.3300 ;
    END
  END SS4BEG[9]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.4152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.664 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 0.0000 140.1550 0.3300 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 0.0000 138.7750 0.3300 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 0.0000 137.3950 0.3300 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 0.0000 136.0150 0.3300 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6287 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.4582 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.992 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 0.0000 134.6350 0.3300 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.29665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.349 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2521 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.437 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.1628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.672 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 0.0000 133.2550 0.3300 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.3894 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 307.488 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 0.0000 131.8750 0.3300 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.23885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.281 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.2048 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 0.0000 130.4950 0.3300 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.0185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 0.0000 129.1150 0.3300 ;
    END
  END SS4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.756 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.7235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.9468 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.6507 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.936 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 219.3100 84.4950 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.01065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5927 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.9528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.552 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 219.3100 83.1150 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.87765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.5263 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 6.1477 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2527 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 219.3100 81.7350 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8825 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.24 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 219.3100 80.3550 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.7936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 287.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 90.8111 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 479.341 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230842 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 219.3100 106.1150 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4275 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1955 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.8087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 298.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.3717 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 415.876 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 219.3100 104.7350 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.4015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.9304 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.3218 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 299.605 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 219.3100 103.3550 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 57.7364 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.403 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 219.3100 102.4350 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2805 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.457 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.5184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 62.2706 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.607 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 219.3100 101.0550 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.078 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.2725 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 59.4373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 316.839 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 219.3100 99.6750 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.99365 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.169 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.2996 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 46.4205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7488 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.1348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.1589 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 370.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 219.3100 98.2950 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9039 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.8168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8006 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 379.122 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 219.3100 96.9150 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7524 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.7085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.792 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 219.3100 95.5350 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8475 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.5463 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 132.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 219.3100 94.1550 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8305 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9587 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.912 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 219.3100 92.7750 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2809 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1542 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 114.704 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 219.3100 91.3950 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6706 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2755 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1408 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.908 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 219.3100 90.0150 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.134 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.7296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.832 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 219.3100 88.6350 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.1301 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.5555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.2618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.2 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 219.3100 87.2550 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.3138 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 1.1304 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.2216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.456 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 219.3100 85.8750 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.8828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 39.3365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3584 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.674 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.37865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 29.4 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 219.3100 127.7350 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.89505 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.053 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8488 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.64929 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.9428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 219.3100 126.3550 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.8452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 54.1485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.7488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.0454 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 426.195 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 219.3100 125.4350 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4864 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.3545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.464 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 30.045 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 219.3100 124.0550 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8484 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.0905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.7313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.7916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 24.9644 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 126.615 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 219.3100 122.6750 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.8316 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 49.0805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2235 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 46.5204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 249.52 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.4341 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.108 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 219.3100 121.2950 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.6556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.294 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.80572 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.938 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 219.3100 119.9150 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5877 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.3276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.688 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 71.7896 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 381.308 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 219.3100 118.5350 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.0738 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 240.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 76.9806 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 406.593 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 219.3100 117.1550 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 22.1976 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 119.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 40.1574 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 215.095 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 219.3100 115.7750 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.5876 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.8605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.4392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.078 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.6707 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 219.3100 114.3950 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.47005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.553 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.2892 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 71.3685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.27152 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.0539 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 219.3100 113.0150 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.8684 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.192 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 219.3100 111.6350 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.28 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.6993 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 72.5095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.1469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9432 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 219.3100 110.2550 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8143 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9468 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.4081 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.72 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 219.3100 108.8750 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8787 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.9504 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.7848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 219.3100 107.4950 219.6400 ;
    END
  END S4END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6492 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 39.6273 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.135 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 219.3100 149.3550 219.6400 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.2758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 60.4189 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 322.9 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 219.3100 148.4350 219.6400 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.47305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 22.0576 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.9 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 219.3100 147.0550 219.6400 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.5233 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.3275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.9446 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 45.9277 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 219.3100 145.6750 219.6400 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.1388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 294.544 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 80.8567 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 430.283 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 219.3100 144.2950 219.6400 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 18.6373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 91.7175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.7096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 10.7549 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 56.1387 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 219.3100 142.9150 219.6400 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 54.8358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 292.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.77 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 419.248 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 219.3100 141.5350 219.6400 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.2048 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.9465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2943 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.3811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 219.3100 140.1550 219.6400 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1208 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.486 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.63946 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.8027 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 219.3100 138.7750 219.6400 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.3364 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 76.6045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.80229 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.6168 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 219.3100 137.3950 219.6400 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.60565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.889 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.6616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.2305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3588 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.69589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.0849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 219.3100 136.0150 219.6400 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.1104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.224 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.65481 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.7205 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 219.3100 134.6350 219.6400 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.9614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.872 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 219.3100 133.2550 219.6400 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.7363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 68.2745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.8706 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.584 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 219.3100 131.8750 219.6400 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5085 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.648 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 219.3100 130.4950 219.6400 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.9545 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 171.36 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 219.3100 129.1150 219.6400 ;
    END
  END SS4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.5676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.5339 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.0365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.1508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.6800 0.4850 12.8200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5062 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 255.248 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 11.3200 0.4850 11.4600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.7654 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112.16 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 9.9600 0.4850 10.1000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.319 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.3858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.01 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.784 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.2 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.5800 0.4850 24.7200 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.21 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.8800 0.4850 23.0200 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.511 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.6986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 138 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 21.5200 0.4850 21.6600 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.931 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.352 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.896 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.1600 0.4850 20.3000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2675 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 154.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.7214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 154.592 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 18.4600 0.4850 18.6000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.2146 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 188.752 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.1000 0.4850 17.2400 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1981 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.6548 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.648 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.1278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.152 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 37.8400 0.4850 37.9800 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.7135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.853 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 36.1400 0.4850 36.2800 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5563 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5025 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.722 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.999 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 34.7800 0.4850 34.9200 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 33.4200 0.4850 33.5600 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 31.7200 0.4850 31.8600 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.657 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 30.3600 0.4850 30.5000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.931 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1306 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 29.0000 0.4850 29.1400 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9903 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.7118 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.6 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.3000 0.4850 27.4400 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.7075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 61.3000 0.4850 61.4400 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 18.9318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.44 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 59.9400 0.4850 60.0800 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.9288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 165.424 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 58.2400 0.4850 58.3800 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 56.8800 0.4850 57.0200 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.818 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 55.5200 0.4850 55.6600 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.773 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.5866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 53.8200 0.4850 53.9600 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.5618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.8 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 52.4600 0.4850 52.6000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.9008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 51.1000 0.4850 51.2400 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 56.5968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 302.32 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 49.4000 0.4850 49.5400 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.807 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.809 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 48.0400 0.4850 48.1800 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.259 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.1386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 46.6800 0.4850 46.8200 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1883 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 43.42 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 232.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.2636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 44.9800 0.4850 45.1200 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6318 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.8 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.952 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 43.6200 0.4850 43.7600 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7141 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.6948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 212.176 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 42.2600 0.4850 42.4000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.459 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.6874 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 40.5600 0.4850 40.7000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9737 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.465 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 39.2000 0.4850 39.3400 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 78.9800 0.4850 79.1200 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.7318 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.04 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 77.6200 0.4850 77.7600 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2456 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.12 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 75.9200 0.4850 76.0600 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 74.5600 0.4850 74.7000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.2426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 295.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 73.2000 0.4850 73.3400 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1581 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6825 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 71.5000 0.4850 71.6400 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 70.1400 0.4850 70.2800 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 17.7496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.522 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 68.7800 0.4850 68.9200 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.444 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.5914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.232 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 67.0800 0.4850 67.2200 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5703 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.9292 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.504 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 65.7200 0.4850 65.8600 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.12 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.632 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 64.3600 0.4850 64.5000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 62.6600 0.4850 62.8000 ;
    END
  END W6BEG[0]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.241 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.4748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 266.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 14.0400 210.2200 14.1800 ;
    END
  END W1END[3]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.7968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 2.088 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.6641 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 12.6800 210.2200 12.8200 ;
    END
  END W1END[2]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2366 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.022 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.692 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.7398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 11.3200 210.2200 11.4600 ;
    END
  END W1END[1]
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5012 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 35.4618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 189.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 9.9600 210.2200 10.1000 ;
    END
  END W1END[0]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.242 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 37.5975 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.456 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 56.8059 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 300.218 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 25.9400 210.2200 26.0800 ;
    END
  END W2MID[7]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 38.8128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 207.472 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 63.7494 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 333.246 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 24.5800 210.2200 24.7200 ;
    END
  END W2MID[6]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.2415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.6715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.4559 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.248 LAYER met3  ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 16.9906 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 85.2983 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 22.8800 210.2200 23.0200 ;
    END
  END W2MID[5]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1575 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5966 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 84.5768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 451.354 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 21.5200 210.2200 21.6600 ;
    END
  END W2MID[4]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.5557 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 18.8632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 101.104 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 20.1600 210.2200 20.3000 ;
    END
  END W2MID[3]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.106 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.711 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.2672 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.274 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 18.4600 210.2200 18.6000 ;
    END
  END W2MID[2]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.2799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.4855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 18.8708 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.3051 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.129832 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 17.1000 210.2200 17.2400 ;
    END
  END W2MID[1]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.4592 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 51.618 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 16.7558 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.7886 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 15.7400 210.2200 15.8800 ;
    END
  END W2MID[0]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.74 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 95.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.9426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.968 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 37.8400 210.2200 37.9800 ;
    END
  END W2END[7]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3314 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.496 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.888 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.1062 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 130.448 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 36.1400 210.2200 36.2800 ;
    END
  END W2END[6]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.293 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.7648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 175.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 34.7800 210.2200 34.9200 ;
    END
  END W2END[5]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3176 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.8182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 33.4200 210.2200 33.5600 ;
    END
  END W2END[4]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.84 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.039 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.0618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.9626 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 75.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 31.7200 210.2200 31.8600 ;
    END
  END W2END[3]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2009 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.699 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1268 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.512 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 30.3600 210.2200 30.5000 ;
    END
  END W2END[2]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.67 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.1304 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.3994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.728 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 29.0000 210.2200 29.1400 ;
    END
  END W2END[1]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8538 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.99 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.85 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.1386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 161.68 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 27.3000 210.2200 27.4400 ;
    END
  END W2END[0]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.566 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.7854 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 33.7682 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 178.156 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 61.3000 210.2200 61.4400 ;
    END
  END WW4END[15]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.73535 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.2458 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 59.9400 210.2200 60.0800 ;
    END
  END WW4END[14]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1457 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.3 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.22 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.457 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 338.481 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 58.2400 210.2200 58.3800 ;
    END
  END WW4END[13]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.83003 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 47.7192 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 56.8800 210.2200 57.0200 ;
    END
  END WW4END[12]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.45185 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.8283 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 55.5200 210.2200 55.6600 ;
    END
  END WW4END[11]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1617 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 41.704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 222.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.4238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8838 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.875 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 53.8200 210.2200 53.9600 ;
    END
  END WW4END[10]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 90.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 24.9131 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 123.117 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 52.4600 210.2200 52.6000 ;
    END
  END WW4END[9]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.48997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.0687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 51.1000 210.2200 51.2400 ;
    END
  END WW4END[8]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.0588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 53.6869 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 283.84 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 49.4000 210.2200 49.5400 ;
    END
  END WW4END[7]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.2101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 75.7715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.5434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 42.8769 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 225.661 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 48.0400 210.2200 48.1800 ;
    END
  END WW4END[6]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.986 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8199 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.268 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 46.6800 210.2200 46.8200 ;
    END
  END WW4END[5]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.651 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.8298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 228.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 66.1234 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 349.923 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 44.9800 210.2200 45.1200 ;
    END
  END WW4END[4]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.266 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.9021 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.688 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 43.6200 210.2200 43.7600 ;
    END
  END WW4END[3]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0477 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7596 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.541 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 111.904 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 42.2600 210.2200 42.4000 ;
    END
  END WW4END[2]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.138 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.8328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 40.5600 210.2200 40.7000 ;
    END
  END WW4END[1]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 31.5148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.104 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 39.2000 210.2200 39.3400 ;
    END
  END WW4END[0]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.901 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.861 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 41.1071 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 220.525 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 78.9800 210.2200 79.1200 ;
    END
  END W6END[11]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 46.5516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 249.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 67.6389 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 358.894 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 77.6200 210.2200 77.7600 ;
    END
  END W6END[10]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.778 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.49024 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.002 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 75.9200 210.2200 76.0600 ;
    END
  END W6END[9]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5345 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 19.282 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 103.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.872 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 63.5222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 333.437 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 74.5600 210.2200 74.7000 ;
    END
  END W6END[8]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.726 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.2064 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 180.864 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 48.3134 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 261.064 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 73.2000 210.2200 73.3400 ;
    END
  END W6END[7]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 44.9987 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 241.515 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 71.5000 210.2200 71.6400 ;
    END
  END W6END[6]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.882 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.68687 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.9535 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 70.1400 210.2200 70.2800 ;
    END
  END W6END[5]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.4078 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 125.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8325 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 244.832 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 68.7800 210.2200 68.9200 ;
    END
  END W6END[4]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.138 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.32835 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.1017 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 67.0800 210.2200 67.2200 ;
    END
  END W6END[3]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.7564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.3463 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.62 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 65.7200 210.2200 65.8600 ;
    END
  END W6END[2]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.457 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.8972 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.8498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 236.208 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 64.3600 210.2200 64.5000 ;
    END
  END W6END[1]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9468 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.7784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.204 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 1.3248 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.8877 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.5156 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 62.6600 210.2200 62.8000 ;
    END
  END W6END[0]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.3906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 51.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 5.65473 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 29.6641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met4 ;
        RECT 88.8600 0.0000 89.1600 0.8000 ;
    END
  END UserCLK
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.2659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.2445 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9915 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.8919 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.646632 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.72 LAYER met3  ;
    ANTENNAGATEAREA 0.9915 LAYER met3  ;
    ANTENNAMAXAREACAR 21.498 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 100.644 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.686975 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.8394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 375.28 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 64.1948 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 332.988 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.842138 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 209.5400 0.4850 209.6800 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.8415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.6736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 63.7308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 344.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 69.8794 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 362.313 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.1566 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 207.8400 0.4850 207.9800 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6796 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.237 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 79.7052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 428.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 77.3028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 403.915 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.910273 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 206.1400 0.4850 206.2800 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.23 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 36.852 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 198.896 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 74.1568 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 393.078 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 204.4400 0.4850 204.5800 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1561 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.9141 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 265.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 62.1352 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.646 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 202.7400 0.4850 202.8800 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.3306 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.795 LAYER met3  ;
    ANTENNAMAXAREACAR 38.1416 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 192.053 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.615723 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.2608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 158.88 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 64.3919 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.808 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 201.0400 0.4850 201.1800 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0585 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met2  ;
    ANTENNAMAXAREACAR 7.69847 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.7852 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.382662 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 8.08748 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 36.5529 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.442053 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.2737 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 156.592 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 47.5344 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 240.446 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.713017 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 199.0000 0.4850 199.1400 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.1195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met2  ;
    ANTENNAMAXAREACAR 18.793 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.3446 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.495326 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAGATEAREA 1.3095 LAYER met3  ;
    ANTENNAMAXAREACAR 19.2565 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.1732 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.525872 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.6416 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 185.696 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 63.3251 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 336.208 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 197.3000 0.4850 197.4400 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9915 LAYER met2  ;
    ANTENNAMAXAREACAR 48.4497 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 235.991 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.686975 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.0837 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.512 LAYER met3  ;
    ANTENNAGATEAREA 1.7865 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6917 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 296.731 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.0127 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.5052 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 100.576 LAYER met4  ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4431 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.99 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 195.6000 0.4850 195.7400 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.666 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.8087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 363.984 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.2175 LAYER met4  ;
    ANTENNAMAXAREACAR 65.4516 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 335.693 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.03082 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 193.9000 0.4850 194.0400 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.1861 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 69.8355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9915 LAYER met2  ;
    ANTENNAMAXAREACAR 43.5096 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 210.94 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.646632 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAGATEAREA 0.9915 LAYER met3  ;
    ANTENNAMAXAREACAR 44.3306 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 215.79 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.686975 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.5585 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.248 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 63.748 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 318.141 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01824 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 192.2000 0.4850 192.3400 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.1019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.1885 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3095 LAYER met2  ;
    ANTENNAMAXAREACAR 38.1985 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 185.413 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.495326 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.5708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.648 LAYER met3  ;
    ANTENNAGATEAREA 2.5815 LAYER met3  ;
    ANTENNAMAXAREACAR 40.3565 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 197.285 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.543168 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.1827 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 81.44 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 45.3206 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.913 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 190.1600 0.4850 190.3000 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9905 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8325 LAYER met2  ;
    ANTENNAMAXAREACAR 62.667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 308.872 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.442073 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAGATEAREA 0.8325 LAYER met3  ;
    ANTENNAMAXAREACAR 62.8959 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 310.63 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.490121 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.3814 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.112 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 73.4832 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 367.558 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 188.4600 0.4850 188.6000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.4508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.56 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8543 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 235.65 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.05878 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 186.7600 0.4850 186.9000 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1491 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.128 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 44.6265 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 241.296 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 53.1585 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.162 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 185.0600 0.4850 185.2000 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.966 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.4543 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 222.496 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 73.2327 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 373.549 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.84653 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 183.3600 0.4850 183.5000 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.399 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.9525 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 56.2596 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 282.58 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 181.3200 0.4850 181.4600 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.84 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.6286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 58.2934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 295.192 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.788679 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 179.6200 0.4850 179.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 55.932 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 300.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 60.7631 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.925 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.06402 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 177.9200 0.4850 178.0600 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0957 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.9752 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 172.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 51.8786 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.945 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.884067 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 176.2200 0.4850 176.3600 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9385 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.1824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5145 LAYER met3  ;
    ANTENNAMAXAREACAR 76.6645 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 399.014 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.775761 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.9252 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.816 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 85.7948 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 448.324 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 174.5200 0.4850 174.6600 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.5324 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 128.735 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 665.059 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 172.4800 0.4850 172.6200 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.6568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.24 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3555 LAYER met3  ;
    ANTENNAMAXAREACAR 53.5936 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.431 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 1.05317 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 69.8577 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 375.392 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 112.034 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 581.2 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.05317 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 170.7800 0.4850 170.9200 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9441 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.8859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 188.384 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.2635 LAYER met3  ;
    ANTENNAMAXAREACAR 51.9561 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 260.909 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.661495 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.9098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 205.008 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 64.351 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.938 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 169.0800 0.4850 169.2200 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.0596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6735 LAYER met3  ;
    ANTENNAMAXAREACAR 70.685 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 361.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.775743 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 48.1776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 259.76 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 109.245 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 578.534 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.72264 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 167.3800 0.4850 167.5200 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2625 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.967 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.3003 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 99.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 60.8865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 304.351 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.00985 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 165.6800 0.4850 165.8200 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.733 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.4223 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 55.6687 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 286.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.03082 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 163.6400 0.4850 163.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5559 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.2094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8007 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 297.073 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 161.9400 0.4850 162.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.8859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.52 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 97.4936 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 504.351 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 62.4135 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 335.68 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 117.9 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 614.104 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.32956 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 160.2400 0.4850 160.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 67.9221 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 366.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 81.9182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.25 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 158.5400 0.4850 158.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.773 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 42.2651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 201.562 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.0468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.52 LAYER met3  ;
    ANTENNAGATEAREA 0.5145 LAYER met3  ;
    ANTENNAMAXAREACAR 67.6234 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 338.627 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.794098 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 41.9055 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.784 LAYER met4  ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 81.3247 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.776 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 156.8400 0.4850 156.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.161 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 47.9706 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 258.656 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0585 LAYER met4  ;
    ANTENNAMAXAREACAR 79.6982 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 409.108 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 155.1400 0.4850 155.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.915 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 209.5400 210.2200 209.6800 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.3215 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 207.8400 210.2200 207.9800 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 206.1400 210.2200 206.2800 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.817 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 204.4400 210.2200 204.5800 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.3022 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.76 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.9508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.208 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 202.7400 210.2200 202.8800 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.237 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.6458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 251.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 201.0400 210.2200 201.1800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.63 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.989 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.176 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1234 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.736 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 199.0000 210.2200 199.1400 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2289 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 42.2968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 226.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 197.3000 210.2200 197.4400 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.736 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.9474 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 195.6000 210.2200 195.7400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4363 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.9555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 193.9000 210.2200 194.0400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.884 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.8144 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 267.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 192.2000 210.2200 192.3400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 39.889 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 213.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 128.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 190.1600 210.2200 190.3000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 188.4600 210.2200 188.6000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2247 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.3954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.52 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 186.7600 210.2200 186.9000 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.682 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 185.0600 210.2200 185.2000 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.6155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.5818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 183.3600 210.2200 183.5000 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2317 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9975 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.645 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.5598 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.456 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 181.3200 210.2200 181.4600 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 122.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.3184 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 173.776 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 179.6200 210.2200 179.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9587 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 59.3635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.1418 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.772 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 177.9200 210.2200 178.0600 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3837 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.5264 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.552 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 176.2200 210.2200 176.3600 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1337 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.4658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.288 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 174.5200 210.2200 174.6600 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.1458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 172.4800 210.2200 172.6200 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7595 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.281 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 124.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.808 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 170.7800 210.2200 170.9200 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 22.222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 169.0800 210.2200 169.2200 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.3405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.5048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.496 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 167.3800 210.2200 167.5200 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.183 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.776 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7614 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 165.6800 210.2200 165.8200 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.4538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.7536 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.96 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 163.6400 210.2200 163.7800 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6973 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 27.904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 149.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.607 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 161.9400 210.2200 162.0800 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.328 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 160.2400 210.2200 160.3800 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8279 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.037 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 158.5400 210.2200 158.6800 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 156.8400 210.2200 156.9800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2387 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 33.029 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.7154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.7350 155.1400 210.2200 155.2800 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.4639 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 146.976 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 40.8166 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 202.384 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 199.3400 0.0000 199.4800 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4231 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.8775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.3325 LAYER met2  ;
    ANTENNAMAXAREACAR 11.9137 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.4781 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 197.5000 0.0000 197.6400 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 34.7655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.113 LAYER met2  ;
    ANTENNAMAXAREACAR 46.5338 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 219.513 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.68248 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAGATEAREA 1.113 LAYER met3  ;
    ANTENNAMAXAREACAR 46.8932 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 221.849 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.718419 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 47.2498 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 223.929 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.807228 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 195.2000 0.0000 195.3400 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1646 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.2097 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.703 LAYER met3  ;
    ANTENNAMAXAREACAR 20.1273 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 92.4769 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.690936 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 20.4268 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 94.1633 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.690936 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 192.9000 0.0000 193.0400 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.1255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 96.7855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9266 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.6672 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.646541 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 190.6000 0.0000 190.7400 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.3481 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 88.3505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met2  ;
    ANTENNAMAXAREACAR 17.3677 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.8194 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.646541 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 188.3000 0.0000 188.4400 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.044 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.643 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 26.3154 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.28 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 57.5709 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.394 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 185.5400 0.0000 185.6800 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.5038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 109.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 34.9184 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.752 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.914087 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 184.1600 0.0000 184.3000 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.393 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.804 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.575 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.0996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 32.3757 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.165 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.774004 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 181.4000 0.0000 181.5400 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9526 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.602 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.5934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 34.1698 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.262 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.669718 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 179.5600 0.0000 179.7000 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.3618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 29.3604 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 144.274 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.975494 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 174.9600 0.0000 175.1000 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9302 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.49 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 38.8422 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.04 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 37.5691 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.026 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.767615 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 172.6600 0.0000 172.8000 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7818 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.748 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 45.2634 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.223 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 210.006 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.772327 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 170.3600 0.0000 170.5000 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.0691 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 141.81 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.3305 LAYER met2  ;
    ANTENNAMAXAREACAR 38.234 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 184.69 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.806524 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.7258 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.808 LAYER met3  ;
    ANTENNAGATEAREA 4.4895 LAYER met3  ;
    ANTENNAMAXAREACAR 39.0639 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 189.325 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.815434 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 40.2292 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 195.629 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.815434 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 168.5200 0.0000 168.6600 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.0132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.41 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 50.0868 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 244.066 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 52.4214 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 257.991 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.637736 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 17.0238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 93.616 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 55.6428 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 275.706 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.01824 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 166.2200 0.0000 166.3600 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.0096 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 224.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 133.334 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 163.9200 0.0000 164.0600 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 32.8329 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 176.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 52.0231 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 266.641 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 161.1600 0.0000 161.3000 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.3308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.568 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8102 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 93.3202 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.65411 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 159.3200 0.0000 159.4600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.3722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 143.388 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.0125 LAYER met2  ;
    ANTENNAMAXAREACAR 22.3768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.034 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.474749 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.416 LAYER met3  ;
    ANTENNAGATEAREA 4.0125 LAYER met3  ;
    ANTENNAMAXAREACAR 22.6081 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 107.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.484718 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.8954 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 203.52 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 37.4738 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 187.317 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 157.0200 0.0000 157.1600 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.947 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.73 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.0378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.672 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 27.9378 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 134.623 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.621428 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 0.0000 155.3200 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2455 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 199.3400 219.1550 199.4800 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.1248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.136 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 197.5000 219.1550 197.6400 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.8114 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.896 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.7494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.3716 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.256 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 194.7400 219.1550 194.8800 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.93 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.528 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 192.9000 219.1550 193.0400 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4294 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.986 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.2068 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 204.24 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 190.6000 219.1550 190.7400 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.3496 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.472 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 188.3000 219.1550 188.4400 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.2495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 186.0000 219.1550 186.1400 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.7643 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.7135 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.1600 219.1550 184.3000 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.243 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.5748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.888 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.4000 219.1550 181.5400 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2403 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0935 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 179.5600 219.1550 179.7000 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 16.5323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 82.4355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 174.9600 219.1550 175.1000 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.6623 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0855 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.6600 219.1550 172.8000 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.8035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 170.3600 219.1550 170.5000 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.1475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 168.5200 219.1550 168.6600 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6123 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.8355 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.2200 219.1550 166.3600 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7811 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6795 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.9200 219.1550 164.0600 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.413 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.803 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.9038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 234.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 161.6200 219.1550 161.7600 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.69 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.9286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 272.56 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 159.3200 219.1550 159.4600 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.9831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 119.69 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 156.5600 219.1550 156.7000 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.652 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.757 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.2648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 327.216 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 155.1800 219.1550 155.3200 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 204.6600 8.4300 ;
        RECT 5.5600 210.5300 204.6600 213.5300 ;
        RECT 5.5600 12.3400 8.5600 12.8200 ;
        RECT 5.5600 17.7800 8.5600 18.2600 ;
        RECT 5.5600 23.2200 8.5600 23.7000 ;
        RECT 5.5600 34.1000 8.5600 34.5800 ;
        RECT 5.5600 28.6600 8.5600 29.1400 ;
        RECT 5.5600 39.5400 8.5600 40.0200 ;
        RECT 5.5600 44.9800 8.5600 45.4600 ;
        RECT 5.5600 50.4200 8.5600 50.9000 ;
        RECT 55.1200 12.3400 56.7200 12.8200 ;
        RECT 55.1200 23.2200 56.7200 23.7000 ;
        RECT 55.1200 17.7800 56.7200 18.2600 ;
        RECT 100.1200 12.3400 101.7200 12.8200 ;
        RECT 100.1200 23.2200 101.7200 23.7000 ;
        RECT 100.1200 17.7800 101.7200 18.2600 ;
        RECT 55.1200 28.6600 56.7200 29.1400 ;
        RECT 55.1200 34.1000 56.7200 34.5800 ;
        RECT 55.1200 39.5400 56.7200 40.0200 ;
        RECT 55.1200 44.9800 56.7200 45.4600 ;
        RECT 55.1200 50.4200 56.7200 50.9000 ;
        RECT 100.1200 28.6600 101.7200 29.1400 ;
        RECT 100.1200 34.1000 101.7200 34.5800 ;
        RECT 100.1200 39.5400 101.7200 40.0200 ;
        RECT 100.1200 44.9800 101.7200 45.4600 ;
        RECT 100.1200 50.4200 101.7200 50.9000 ;
        RECT 5.5600 61.3000 8.5600 61.7800 ;
        RECT 5.5600 55.8600 8.5600 56.3400 ;
        RECT 5.5600 66.7400 8.5600 67.2200 ;
        RECT 5.5600 72.1800 8.5600 72.6600 ;
        RECT 5.5600 77.6200 8.5600 78.1000 ;
        RECT 5.5600 88.5000 8.5600 88.9800 ;
        RECT 5.5600 83.0600 8.5600 83.5400 ;
        RECT 5.5600 93.9400 8.5600 94.4200 ;
        RECT 5.5600 99.3800 8.5600 99.8600 ;
        RECT 5.5600 104.8200 8.5600 105.3000 ;
        RECT 55.1200 55.8600 56.7200 56.3400 ;
        RECT 55.1200 61.3000 56.7200 61.7800 ;
        RECT 55.1200 66.7400 56.7200 67.2200 ;
        RECT 55.1200 72.1800 56.7200 72.6600 ;
        RECT 55.1200 77.6200 56.7200 78.1000 ;
        RECT 100.1200 55.8600 101.7200 56.3400 ;
        RECT 100.1200 61.3000 101.7200 61.7800 ;
        RECT 100.1200 66.7400 101.7200 67.2200 ;
        RECT 100.1200 72.1800 101.7200 72.6600 ;
        RECT 100.1200 77.6200 101.7200 78.1000 ;
        RECT 55.1200 83.0600 56.7200 83.5400 ;
        RECT 55.1200 88.5000 56.7200 88.9800 ;
        RECT 55.1200 93.9400 56.7200 94.4200 ;
        RECT 55.1200 99.3800 56.7200 99.8600 ;
        RECT 55.1200 104.8200 56.7200 105.3000 ;
        RECT 100.1200 83.0600 101.7200 83.5400 ;
        RECT 100.1200 88.5000 101.7200 88.9800 ;
        RECT 100.1200 93.9400 101.7200 94.4200 ;
        RECT 100.1200 99.3800 101.7200 99.8600 ;
        RECT 100.1200 104.8200 101.7200 105.3000 ;
        RECT 145.1200 12.3400 146.7200 12.8200 ;
        RECT 145.1200 17.7800 146.7200 18.2600 ;
        RECT 145.1200 23.2200 146.7200 23.7000 ;
        RECT 145.1200 28.6600 146.7200 29.1400 ;
        RECT 145.1200 34.1000 146.7200 34.5800 ;
        RECT 145.1200 39.5400 146.7200 40.0200 ;
        RECT 145.1200 44.9800 146.7200 45.4600 ;
        RECT 145.1200 50.4200 146.7200 50.9000 ;
        RECT 201.6600 12.3400 204.6600 12.8200 ;
        RECT 190.1200 12.3400 191.7200 12.8200 ;
        RECT 190.1200 17.7800 191.7200 18.2600 ;
        RECT 190.1200 23.2200 191.7200 23.7000 ;
        RECT 201.6600 17.7800 204.6600 18.2600 ;
        RECT 201.6600 23.2200 204.6600 23.7000 ;
        RECT 190.1200 28.6600 191.7200 29.1400 ;
        RECT 190.1200 34.1000 191.7200 34.5800 ;
        RECT 190.1200 39.5400 191.7200 40.0200 ;
        RECT 201.6600 28.6600 204.6600 29.1400 ;
        RECT 201.6600 34.1000 204.6600 34.5800 ;
        RECT 201.6600 39.5400 204.6600 40.0200 ;
        RECT 190.1200 44.9800 191.7200 45.4600 ;
        RECT 190.1200 50.4200 191.7200 50.9000 ;
        RECT 201.6600 44.9800 204.6600 45.4600 ;
        RECT 201.6600 50.4200 204.6600 50.9000 ;
        RECT 145.1200 55.8600 146.7200 56.3400 ;
        RECT 145.1200 61.3000 146.7200 61.7800 ;
        RECT 145.1200 66.7400 146.7200 67.2200 ;
        RECT 145.1200 72.1800 146.7200 72.6600 ;
        RECT 145.1200 77.6200 146.7200 78.1000 ;
        RECT 145.1200 83.0600 146.7200 83.5400 ;
        RECT 145.1200 88.5000 146.7200 88.9800 ;
        RECT 145.1200 93.9400 146.7200 94.4200 ;
        RECT 145.1200 99.3800 146.7200 99.8600 ;
        RECT 145.1200 104.8200 146.7200 105.3000 ;
        RECT 190.1200 55.8600 191.7200 56.3400 ;
        RECT 190.1200 61.3000 191.7200 61.7800 ;
        RECT 190.1200 66.7400 191.7200 67.2200 ;
        RECT 201.6600 55.8600 204.6600 56.3400 ;
        RECT 201.6600 61.3000 204.6600 61.7800 ;
        RECT 201.6600 66.7400 204.6600 67.2200 ;
        RECT 190.1200 72.1800 191.7200 72.6600 ;
        RECT 190.1200 77.6200 191.7200 78.1000 ;
        RECT 201.6600 72.1800 204.6600 72.6600 ;
        RECT 201.6600 77.6200 204.6600 78.1000 ;
        RECT 190.1200 83.0600 191.7200 83.5400 ;
        RECT 190.1200 88.5000 191.7200 88.9800 ;
        RECT 190.1200 93.9400 191.7200 94.4200 ;
        RECT 201.6600 83.0600 204.6600 83.5400 ;
        RECT 201.6600 88.5000 204.6600 88.9800 ;
        RECT 201.6600 93.9400 204.6600 94.4200 ;
        RECT 190.1200 99.3800 191.7200 99.8600 ;
        RECT 190.1200 104.8200 191.7200 105.3000 ;
        RECT 201.6600 99.3800 204.6600 99.8600 ;
        RECT 201.6600 104.8200 204.6600 105.3000 ;
        RECT 5.5600 164.6600 8.5600 165.1400 ;
        RECT 55.1200 164.6600 56.7200 165.1400 ;
        RECT 100.1200 164.6600 101.7200 165.1400 ;
        RECT 5.5600 115.7000 8.5600 116.1800 ;
        RECT 5.5600 110.2600 8.5600 110.7400 ;
        RECT 5.5600 121.1400 8.5600 121.6200 ;
        RECT 5.5600 126.5800 8.5600 127.0600 ;
        RECT 5.5600 132.0200 8.5600 132.5000 ;
        RECT 5.5600 142.9000 8.5600 143.3800 ;
        RECT 5.5600 137.4600 8.5600 137.9400 ;
        RECT 5.5600 148.3400 8.5600 148.8200 ;
        RECT 5.5600 153.7800 8.5600 154.2600 ;
        RECT 5.5600 159.2200 8.5600 159.7000 ;
        RECT 55.1200 110.2600 56.7200 110.7400 ;
        RECT 55.1200 115.7000 56.7200 116.1800 ;
        RECT 55.1200 121.1400 56.7200 121.6200 ;
        RECT 55.1200 126.5800 56.7200 127.0600 ;
        RECT 55.1200 132.0200 56.7200 132.5000 ;
        RECT 100.1200 110.2600 101.7200 110.7400 ;
        RECT 100.1200 115.7000 101.7200 116.1800 ;
        RECT 100.1200 121.1400 101.7200 121.6200 ;
        RECT 100.1200 126.5800 101.7200 127.0600 ;
        RECT 100.1200 132.0200 101.7200 132.5000 ;
        RECT 55.1200 137.4600 56.7200 137.9400 ;
        RECT 55.1200 142.9000 56.7200 143.3800 ;
        RECT 55.1200 148.3400 56.7200 148.8200 ;
        RECT 55.1200 153.7800 56.7200 154.2600 ;
        RECT 55.1200 159.2200 56.7200 159.7000 ;
        RECT 100.1200 137.4600 101.7200 137.9400 ;
        RECT 100.1200 142.9000 101.7200 143.3800 ;
        RECT 100.1200 148.3400 101.7200 148.8200 ;
        RECT 100.1200 153.7800 101.7200 154.2600 ;
        RECT 100.1200 159.2200 101.7200 159.7000 ;
        RECT 5.5600 191.8600 8.5600 192.3400 ;
        RECT 5.5600 175.5400 8.5600 176.0200 ;
        RECT 5.5600 170.1000 8.5600 170.5800 ;
        RECT 5.5600 186.4200 8.5600 186.9000 ;
        RECT 5.5600 180.9800 8.5600 181.4600 ;
        RECT 5.5600 202.7400 8.5600 203.2200 ;
        RECT 5.5600 197.3000 8.5600 197.7800 ;
        RECT 5.5600 208.1800 8.5600 208.6600 ;
        RECT 55.1200 191.8600 56.7200 192.3400 ;
        RECT 100.1200 191.8600 101.7200 192.3400 ;
        RECT 55.1200 170.1000 56.7200 170.5800 ;
        RECT 55.1200 175.5400 56.7200 176.0200 ;
        RECT 55.1200 180.9800 56.7200 181.4600 ;
        RECT 55.1200 186.4200 56.7200 186.9000 ;
        RECT 100.1200 170.1000 101.7200 170.5800 ;
        RECT 100.1200 175.5400 101.7200 176.0200 ;
        RECT 100.1200 180.9800 101.7200 181.4600 ;
        RECT 100.1200 186.4200 101.7200 186.9000 ;
        RECT 55.1200 197.3000 56.7200 197.7800 ;
        RECT 55.1200 202.7400 56.7200 203.2200 ;
        RECT 55.1200 208.1800 56.7200 208.6600 ;
        RECT 100.1200 197.3000 101.7200 197.7800 ;
        RECT 100.1200 202.7400 101.7200 203.2200 ;
        RECT 100.1200 208.1800 101.7200 208.6600 ;
        RECT 201.6600 164.6600 204.6600 165.1400 ;
        RECT 145.1200 164.6600 146.7200 165.1400 ;
        RECT 190.1200 164.6600 191.7200 165.1400 ;
        RECT 145.1200 110.2600 146.7200 110.7400 ;
        RECT 145.1200 115.7000 146.7200 116.1800 ;
        RECT 145.1200 121.1400 146.7200 121.6200 ;
        RECT 145.1200 126.5800 146.7200 127.0600 ;
        RECT 145.1200 132.0200 146.7200 132.5000 ;
        RECT 145.1200 137.4600 146.7200 137.9400 ;
        RECT 145.1200 142.9000 146.7200 143.3800 ;
        RECT 145.1200 148.3400 146.7200 148.8200 ;
        RECT 145.1200 153.7800 146.7200 154.2600 ;
        RECT 145.1200 159.2200 146.7200 159.7000 ;
        RECT 190.1200 110.2600 191.7200 110.7400 ;
        RECT 190.1200 115.7000 191.7200 116.1800 ;
        RECT 190.1200 121.1400 191.7200 121.6200 ;
        RECT 201.6600 110.2600 204.6600 110.7400 ;
        RECT 201.6600 115.7000 204.6600 116.1800 ;
        RECT 201.6600 121.1400 204.6600 121.6200 ;
        RECT 190.1200 126.5800 191.7200 127.0600 ;
        RECT 190.1200 132.0200 191.7200 132.5000 ;
        RECT 201.6600 126.5800 204.6600 127.0600 ;
        RECT 201.6600 132.0200 204.6600 132.5000 ;
        RECT 190.1200 137.4600 191.7200 137.9400 ;
        RECT 190.1200 142.9000 191.7200 143.3800 ;
        RECT 190.1200 148.3400 191.7200 148.8200 ;
        RECT 201.6600 137.4600 204.6600 137.9400 ;
        RECT 201.6600 142.9000 204.6600 143.3800 ;
        RECT 201.6600 148.3400 204.6600 148.8200 ;
        RECT 190.1200 153.7800 191.7200 154.2600 ;
        RECT 190.1200 159.2200 191.7200 159.7000 ;
        RECT 201.6600 153.7800 204.6600 154.2600 ;
        RECT 201.6600 159.2200 204.6600 159.7000 ;
        RECT 145.1200 191.8600 146.7200 192.3400 ;
        RECT 145.1200 175.5400 146.7200 176.0200 ;
        RECT 145.1200 170.1000 146.7200 170.5800 ;
        RECT 145.1200 180.9800 146.7200 181.4600 ;
        RECT 145.1200 186.4200 146.7200 186.9000 ;
        RECT 145.1200 197.3000 146.7200 197.7800 ;
        RECT 145.1200 202.7400 146.7200 203.2200 ;
        RECT 145.1200 208.1800 146.7200 208.6600 ;
        RECT 201.6600 191.8600 204.6600 192.3400 ;
        RECT 190.1200 191.8600 191.7200 192.3400 ;
        RECT 190.1200 170.1000 191.7200 170.5800 ;
        RECT 190.1200 175.5400 191.7200 176.0200 ;
        RECT 201.6600 170.1000 204.6600 170.5800 ;
        RECT 201.6600 175.5400 204.6600 176.0200 ;
        RECT 190.1200 180.9800 191.7200 181.4600 ;
        RECT 190.1200 186.4200 191.7200 186.9000 ;
        RECT 201.6600 180.9800 204.6600 181.4600 ;
        RECT 201.6600 186.4200 204.6600 186.9000 ;
        RECT 190.1200 197.3000 191.7200 197.7800 ;
        RECT 190.1200 202.7400 191.7200 203.2200 ;
        RECT 201.6600 197.3000 204.6600 197.7800 ;
        RECT 201.6600 202.7400 204.6600 203.2200 ;
        RECT 201.6600 208.1800 204.6600 208.6600 ;
        RECT 190.1200 208.1800 191.7200 208.6600 ;
      LAYER met4 ;
        RECT 190.1200 5.4300 191.7200 213.5300 ;
        RECT 145.1200 5.4300 146.7200 213.5300 ;
        RECT 100.1200 5.4300 101.7200 213.5300 ;
        RECT 55.1200 5.4300 56.7200 213.5300 ;
        RECT 201.6600 5.4300 204.6600 213.5300 ;
        RECT 5.5600 5.4300 8.5600 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 1.5600 1.4300 208.6600 4.4300 ;
        RECT 1.5600 214.5300 208.6600 217.5300 ;
        RECT 1.5600 9.6200 4.5600 10.1000 ;
        RECT 13.3200 9.6200 14.9200 10.1000 ;
        RECT 1.5600 15.0600 4.5600 15.5400 ;
        RECT 1.5600 20.5000 4.5600 20.9800 ;
        RECT 1.5600 25.9400 4.5600 26.4200 ;
        RECT 13.3200 15.0600 14.9200 15.5400 ;
        RECT 13.3200 20.5000 14.9200 20.9800 ;
        RECT 13.3200 25.9400 14.9200 26.4200 ;
        RECT 1.5600 31.3800 4.5600 31.8600 ;
        RECT 1.5600 36.8200 4.5600 37.3000 ;
        RECT 13.3200 31.3800 14.9200 31.8600 ;
        RECT 13.3200 36.8200 14.9200 37.3000 ;
        RECT 1.5600 42.2600 4.5600 42.7400 ;
        RECT 1.5600 47.7000 4.5600 48.1800 ;
        RECT 1.5600 53.1400 4.5600 53.6200 ;
        RECT 13.3200 42.2600 14.9200 42.7400 ;
        RECT 13.3200 47.7000 14.9200 48.1800 ;
        RECT 13.3200 53.1400 14.9200 53.6200 ;
        RECT 58.3200 9.6200 59.9200 10.1000 ;
        RECT 58.3200 15.0600 59.9200 15.5400 ;
        RECT 58.3200 20.5000 59.9200 20.9800 ;
        RECT 58.3200 25.9400 59.9200 26.4200 ;
        RECT 103.3200 9.6200 104.9200 10.1000 ;
        RECT 103.3200 15.0600 104.9200 15.5400 ;
        RECT 103.3200 20.5000 104.9200 20.9800 ;
        RECT 103.3200 25.9400 104.9200 26.4200 ;
        RECT 58.3200 31.3800 59.9200 31.8600 ;
        RECT 58.3200 36.8200 59.9200 37.3000 ;
        RECT 58.3200 42.2600 59.9200 42.7400 ;
        RECT 58.3200 47.7000 59.9200 48.1800 ;
        RECT 58.3200 53.1400 59.9200 53.6200 ;
        RECT 103.3200 31.3800 104.9200 31.8600 ;
        RECT 103.3200 36.8200 104.9200 37.3000 ;
        RECT 103.3200 42.2600 104.9200 42.7400 ;
        RECT 103.3200 47.7000 104.9200 48.1800 ;
        RECT 103.3200 53.1400 104.9200 53.6200 ;
        RECT 1.5600 58.5800 4.5600 59.0600 ;
        RECT 1.5600 64.0200 4.5600 64.5000 ;
        RECT 13.3200 58.5800 14.9200 59.0600 ;
        RECT 13.3200 64.0200 14.9200 64.5000 ;
        RECT 1.5600 69.4600 4.5600 69.9400 ;
        RECT 1.5600 74.9000 4.5600 75.3800 ;
        RECT 1.5600 80.3400 4.5600 80.8200 ;
        RECT 13.3200 69.4600 14.9200 69.9400 ;
        RECT 13.3200 74.9000 14.9200 75.3800 ;
        RECT 13.3200 80.3400 14.9200 80.8200 ;
        RECT 1.5600 85.7800 4.5600 86.2600 ;
        RECT 1.5600 91.2200 4.5600 91.7000 ;
        RECT 13.3200 85.7800 14.9200 86.2600 ;
        RECT 13.3200 91.2200 14.9200 91.7000 ;
        RECT 1.5600 96.6600 4.5600 97.1400 ;
        RECT 1.5600 102.1000 4.5600 102.5800 ;
        RECT 1.5600 107.5400 4.5600 108.0200 ;
        RECT 13.3200 96.6600 14.9200 97.1400 ;
        RECT 13.3200 102.1000 14.9200 102.5800 ;
        RECT 13.3200 107.5400 14.9200 108.0200 ;
        RECT 58.3200 58.5800 59.9200 59.0600 ;
        RECT 58.3200 64.0200 59.9200 64.5000 ;
        RECT 58.3200 69.4600 59.9200 69.9400 ;
        RECT 58.3200 74.9000 59.9200 75.3800 ;
        RECT 58.3200 80.3400 59.9200 80.8200 ;
        RECT 103.3200 58.5800 104.9200 59.0600 ;
        RECT 103.3200 64.0200 104.9200 64.5000 ;
        RECT 103.3200 69.4600 104.9200 69.9400 ;
        RECT 103.3200 74.9000 104.9200 75.3800 ;
        RECT 103.3200 80.3400 104.9200 80.8200 ;
        RECT 58.3200 85.7800 59.9200 86.2600 ;
        RECT 58.3200 91.2200 59.9200 91.7000 ;
        RECT 58.3200 96.6600 59.9200 97.1400 ;
        RECT 58.3200 102.1000 59.9200 102.5800 ;
        RECT 58.3200 107.5400 59.9200 108.0200 ;
        RECT 103.3200 85.7800 104.9200 86.2600 ;
        RECT 103.3200 91.2200 104.9200 91.7000 ;
        RECT 103.3200 96.6600 104.9200 97.1400 ;
        RECT 103.3200 102.1000 104.9200 102.5800 ;
        RECT 103.3200 107.5400 104.9200 108.0200 ;
        RECT 148.3200 9.6200 149.9200 10.1000 ;
        RECT 148.3200 15.0600 149.9200 15.5400 ;
        RECT 148.3200 20.5000 149.9200 20.9800 ;
        RECT 148.3200 25.9400 149.9200 26.4200 ;
        RECT 148.3200 31.3800 149.9200 31.8600 ;
        RECT 148.3200 36.8200 149.9200 37.3000 ;
        RECT 148.3200 42.2600 149.9200 42.7400 ;
        RECT 148.3200 47.7000 149.9200 48.1800 ;
        RECT 148.3200 53.1400 149.9200 53.6200 ;
        RECT 205.6600 9.6200 208.6600 10.1000 ;
        RECT 193.3200 9.6200 194.9200 10.1000 ;
        RECT 193.3200 15.0600 194.9200 15.5400 ;
        RECT 193.3200 20.5000 194.9200 20.9800 ;
        RECT 193.3200 25.9400 194.9200 26.4200 ;
        RECT 205.6600 15.0600 208.6600 15.5400 ;
        RECT 205.6600 20.5000 208.6600 20.9800 ;
        RECT 205.6600 25.9400 208.6600 26.4200 ;
        RECT 193.3200 31.3800 194.9200 31.8600 ;
        RECT 193.3200 36.8200 194.9200 37.3000 ;
        RECT 205.6600 31.3800 208.6600 31.8600 ;
        RECT 205.6600 36.8200 208.6600 37.3000 ;
        RECT 193.3200 42.2600 194.9200 42.7400 ;
        RECT 193.3200 47.7000 194.9200 48.1800 ;
        RECT 193.3200 53.1400 194.9200 53.6200 ;
        RECT 205.6600 42.2600 208.6600 42.7400 ;
        RECT 205.6600 47.7000 208.6600 48.1800 ;
        RECT 205.6600 53.1400 208.6600 53.6200 ;
        RECT 148.3200 58.5800 149.9200 59.0600 ;
        RECT 148.3200 64.0200 149.9200 64.5000 ;
        RECT 148.3200 69.4600 149.9200 69.9400 ;
        RECT 148.3200 74.9000 149.9200 75.3800 ;
        RECT 148.3200 80.3400 149.9200 80.8200 ;
        RECT 148.3200 85.7800 149.9200 86.2600 ;
        RECT 148.3200 91.2200 149.9200 91.7000 ;
        RECT 148.3200 96.6600 149.9200 97.1400 ;
        RECT 148.3200 102.1000 149.9200 102.5800 ;
        RECT 148.3200 107.5400 149.9200 108.0200 ;
        RECT 193.3200 58.5800 194.9200 59.0600 ;
        RECT 193.3200 64.0200 194.9200 64.5000 ;
        RECT 205.6600 58.5800 208.6600 59.0600 ;
        RECT 205.6600 64.0200 208.6600 64.5000 ;
        RECT 193.3200 69.4600 194.9200 69.9400 ;
        RECT 193.3200 74.9000 194.9200 75.3800 ;
        RECT 193.3200 80.3400 194.9200 80.8200 ;
        RECT 205.6600 69.4600 208.6600 69.9400 ;
        RECT 205.6600 74.9000 208.6600 75.3800 ;
        RECT 205.6600 80.3400 208.6600 80.8200 ;
        RECT 193.3200 85.7800 194.9200 86.2600 ;
        RECT 193.3200 91.2200 194.9200 91.7000 ;
        RECT 205.6600 85.7800 208.6600 86.2600 ;
        RECT 205.6600 91.2200 208.6600 91.7000 ;
        RECT 193.3200 96.6600 194.9200 97.1400 ;
        RECT 193.3200 102.1000 194.9200 102.5800 ;
        RECT 193.3200 107.5400 194.9200 108.0200 ;
        RECT 205.6600 96.6600 208.6600 97.1400 ;
        RECT 205.6600 102.1000 208.6600 102.5800 ;
        RECT 205.6600 107.5400 208.6600 108.0200 ;
        RECT 1.5600 112.9800 4.5600 113.4600 ;
        RECT 1.5600 118.4200 4.5600 118.9000 ;
        RECT 13.3200 112.9800 14.9200 113.4600 ;
        RECT 13.3200 118.4200 14.9200 118.9000 ;
        RECT 1.5600 123.8600 4.5600 124.3400 ;
        RECT 1.5600 129.3000 4.5600 129.7800 ;
        RECT 1.5600 134.7400 4.5600 135.2200 ;
        RECT 13.3200 123.8600 14.9200 124.3400 ;
        RECT 13.3200 129.3000 14.9200 129.7800 ;
        RECT 13.3200 134.7400 14.9200 135.2200 ;
        RECT 1.5600 140.1800 4.5600 140.6600 ;
        RECT 1.5600 145.6200 4.5600 146.1000 ;
        RECT 13.3200 140.1800 14.9200 140.6600 ;
        RECT 13.3200 145.6200 14.9200 146.1000 ;
        RECT 1.5600 151.0600 4.5600 151.5400 ;
        RECT 1.5600 156.5000 4.5600 156.9800 ;
        RECT 1.5600 161.9400 4.5600 162.4200 ;
        RECT 13.3200 151.0600 14.9200 151.5400 ;
        RECT 13.3200 156.5000 14.9200 156.9800 ;
        RECT 13.3200 161.9400 14.9200 162.4200 ;
        RECT 58.3200 112.9800 59.9200 113.4600 ;
        RECT 58.3200 118.4200 59.9200 118.9000 ;
        RECT 58.3200 123.8600 59.9200 124.3400 ;
        RECT 58.3200 129.3000 59.9200 129.7800 ;
        RECT 58.3200 134.7400 59.9200 135.2200 ;
        RECT 103.3200 112.9800 104.9200 113.4600 ;
        RECT 103.3200 118.4200 104.9200 118.9000 ;
        RECT 103.3200 123.8600 104.9200 124.3400 ;
        RECT 103.3200 129.3000 104.9200 129.7800 ;
        RECT 103.3200 134.7400 104.9200 135.2200 ;
        RECT 58.3200 140.1800 59.9200 140.6600 ;
        RECT 58.3200 145.6200 59.9200 146.1000 ;
        RECT 58.3200 151.0600 59.9200 151.5400 ;
        RECT 58.3200 156.5000 59.9200 156.9800 ;
        RECT 58.3200 161.9400 59.9200 162.4200 ;
        RECT 103.3200 140.1800 104.9200 140.6600 ;
        RECT 103.3200 145.6200 104.9200 146.1000 ;
        RECT 103.3200 151.0600 104.9200 151.5400 ;
        RECT 103.3200 156.5000 104.9200 156.9800 ;
        RECT 103.3200 161.9400 104.9200 162.4200 ;
        RECT 1.5600 178.2600 4.5600 178.7400 ;
        RECT 13.3200 178.2600 14.9200 178.7400 ;
        RECT 1.5600 172.8200 4.5600 173.3000 ;
        RECT 1.5600 167.3800 4.5600 167.8600 ;
        RECT 13.3200 167.3800 14.9200 167.8600 ;
        RECT 13.3200 172.8200 14.9200 173.3000 ;
        RECT 1.5600 189.1400 4.5600 189.6200 ;
        RECT 1.5600 183.7000 4.5600 184.1800 ;
        RECT 13.3200 183.7000 14.9200 184.1800 ;
        RECT 13.3200 189.1400 14.9200 189.6200 ;
        RECT 1.5600 205.4600 4.5600 205.9400 ;
        RECT 13.3200 205.4600 14.9200 205.9400 ;
        RECT 1.5600 200.0200 4.5600 200.5000 ;
        RECT 1.5600 194.5800 4.5600 195.0600 ;
        RECT 13.3200 194.5800 14.9200 195.0600 ;
        RECT 13.3200 200.0200 14.9200 200.5000 ;
        RECT 58.3200 178.2600 59.9200 178.7400 ;
        RECT 58.3200 167.3800 59.9200 167.8600 ;
        RECT 58.3200 172.8200 59.9200 173.3000 ;
        RECT 58.3200 183.7000 59.9200 184.1800 ;
        RECT 58.3200 189.1400 59.9200 189.6200 ;
        RECT 103.3200 178.2600 104.9200 178.7400 ;
        RECT 103.3200 167.3800 104.9200 167.8600 ;
        RECT 103.3200 172.8200 104.9200 173.3000 ;
        RECT 103.3200 183.7000 104.9200 184.1800 ;
        RECT 103.3200 189.1400 104.9200 189.6200 ;
        RECT 58.3200 194.5800 59.9200 195.0600 ;
        RECT 58.3200 200.0200 59.9200 200.5000 ;
        RECT 58.3200 205.4600 59.9200 205.9400 ;
        RECT 103.3200 194.5800 104.9200 195.0600 ;
        RECT 103.3200 200.0200 104.9200 200.5000 ;
        RECT 103.3200 205.4600 104.9200 205.9400 ;
        RECT 148.3200 112.9800 149.9200 113.4600 ;
        RECT 148.3200 118.4200 149.9200 118.9000 ;
        RECT 148.3200 123.8600 149.9200 124.3400 ;
        RECT 148.3200 129.3000 149.9200 129.7800 ;
        RECT 148.3200 134.7400 149.9200 135.2200 ;
        RECT 148.3200 140.1800 149.9200 140.6600 ;
        RECT 148.3200 145.6200 149.9200 146.1000 ;
        RECT 148.3200 151.0600 149.9200 151.5400 ;
        RECT 148.3200 156.5000 149.9200 156.9800 ;
        RECT 148.3200 161.9400 149.9200 162.4200 ;
        RECT 193.3200 112.9800 194.9200 113.4600 ;
        RECT 193.3200 118.4200 194.9200 118.9000 ;
        RECT 205.6600 112.9800 208.6600 113.4600 ;
        RECT 205.6600 118.4200 208.6600 118.9000 ;
        RECT 193.3200 123.8600 194.9200 124.3400 ;
        RECT 193.3200 129.3000 194.9200 129.7800 ;
        RECT 193.3200 134.7400 194.9200 135.2200 ;
        RECT 205.6600 123.8600 208.6600 124.3400 ;
        RECT 205.6600 129.3000 208.6600 129.7800 ;
        RECT 205.6600 134.7400 208.6600 135.2200 ;
        RECT 193.3200 140.1800 194.9200 140.6600 ;
        RECT 193.3200 145.6200 194.9200 146.1000 ;
        RECT 205.6600 140.1800 208.6600 140.6600 ;
        RECT 205.6600 145.6200 208.6600 146.1000 ;
        RECT 193.3200 151.0600 194.9200 151.5400 ;
        RECT 193.3200 156.5000 194.9200 156.9800 ;
        RECT 193.3200 161.9400 194.9200 162.4200 ;
        RECT 205.6600 151.0600 208.6600 151.5400 ;
        RECT 205.6600 156.5000 208.6600 156.9800 ;
        RECT 205.6600 161.9400 208.6600 162.4200 ;
        RECT 148.3200 178.2600 149.9200 178.7400 ;
        RECT 148.3200 167.3800 149.9200 167.8600 ;
        RECT 148.3200 172.8200 149.9200 173.3000 ;
        RECT 148.3200 183.7000 149.9200 184.1800 ;
        RECT 148.3200 189.1400 149.9200 189.6200 ;
        RECT 148.3200 194.5800 149.9200 195.0600 ;
        RECT 148.3200 200.0200 149.9200 200.5000 ;
        RECT 148.3200 205.4600 149.9200 205.9400 ;
        RECT 205.6600 178.2600 208.6600 178.7400 ;
        RECT 193.3200 178.2600 194.9200 178.7400 ;
        RECT 193.3200 167.3800 194.9200 167.8600 ;
        RECT 193.3200 172.8200 194.9200 173.3000 ;
        RECT 205.6600 167.3800 208.6600 167.8600 ;
        RECT 205.6600 172.8200 208.6600 173.3000 ;
        RECT 193.3200 183.7000 194.9200 184.1800 ;
        RECT 193.3200 189.1400 194.9200 189.6200 ;
        RECT 205.6600 183.7000 208.6600 184.1800 ;
        RECT 205.6600 189.1400 208.6600 189.6200 ;
        RECT 205.6600 205.4600 208.6600 205.9400 ;
        RECT 193.3200 205.4600 194.9200 205.9400 ;
        RECT 193.3200 194.5800 194.9200 195.0600 ;
        RECT 193.3200 200.0200 194.9200 200.5000 ;
        RECT 205.6600 194.5800 208.6600 195.0600 ;
        RECT 205.6600 200.0200 208.6600 200.5000 ;
      LAYER met4 ;
        RECT 193.3200 1.4300 194.9200 217.5300 ;
        RECT 148.3200 1.4300 149.9200 217.5300 ;
        RECT 103.3200 1.4300 104.9200 217.5300 ;
        RECT 58.3200 1.4300 59.9200 217.5300 ;
        RECT 13.3200 1.4300 14.9200 217.5300 ;
        RECT 205.6600 1.4300 208.6600 217.5300 ;
        RECT 1.5600 1.4300 4.5600 217.5300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.5250 219.1400 210.2200 219.6400 ;
      RECT 148.6050 219.1400 149.0150 219.6400 ;
      RECT 147.2250 219.1400 148.0950 219.6400 ;
      RECT 145.8450 219.1400 146.7150 219.6400 ;
      RECT 144.4650 219.1400 145.3350 219.6400 ;
      RECT 143.0850 219.1400 143.9550 219.6400 ;
      RECT 141.7050 219.1400 142.5750 219.6400 ;
      RECT 140.3250 219.1400 141.1950 219.6400 ;
      RECT 138.9450 219.1400 139.8150 219.6400 ;
      RECT 137.5650 219.1400 138.4350 219.6400 ;
      RECT 136.1850 219.1400 137.0550 219.6400 ;
      RECT 134.8050 219.1400 135.6750 219.6400 ;
      RECT 133.4250 219.1400 134.2950 219.6400 ;
      RECT 132.0450 219.1400 132.9150 219.6400 ;
      RECT 130.6650 219.1400 131.5350 219.6400 ;
      RECT 129.2850 219.1400 130.1550 219.6400 ;
      RECT 127.9050 219.1400 128.7750 219.6400 ;
      RECT 126.5250 219.1400 127.3950 219.6400 ;
      RECT 125.6050 219.1400 126.0150 219.6400 ;
      RECT 124.2250 219.1400 125.0950 219.6400 ;
      RECT 122.8450 219.1400 123.7150 219.6400 ;
      RECT 121.4650 219.1400 122.3350 219.6400 ;
      RECT 120.0850 219.1400 120.9550 219.6400 ;
      RECT 118.7050 219.1400 119.5750 219.6400 ;
      RECT 117.3250 219.1400 118.1950 219.6400 ;
      RECT 115.9450 219.1400 116.8150 219.6400 ;
      RECT 114.5650 219.1400 115.4350 219.6400 ;
      RECT 113.1850 219.1400 114.0550 219.6400 ;
      RECT 111.8050 219.1400 112.6750 219.6400 ;
      RECT 110.4250 219.1400 111.2950 219.6400 ;
      RECT 109.0450 219.1400 109.9150 219.6400 ;
      RECT 107.6650 219.1400 108.5350 219.6400 ;
      RECT 106.2850 219.1400 107.1550 219.6400 ;
      RECT 104.9050 219.1400 105.7750 219.6400 ;
      RECT 103.5250 219.1400 104.3950 219.6400 ;
      RECT 102.6050 219.1400 103.0150 219.6400 ;
      RECT 101.2250 219.1400 102.0950 219.6400 ;
      RECT 99.8450 219.1400 100.7150 219.6400 ;
      RECT 98.4650 219.1400 99.3350 219.6400 ;
      RECT 97.0850 219.1400 97.9550 219.6400 ;
      RECT 95.7050 219.1400 96.5750 219.6400 ;
      RECT 94.3250 219.1400 95.1950 219.6400 ;
      RECT 92.9450 219.1400 93.8150 219.6400 ;
      RECT 91.5650 219.1400 92.4350 219.6400 ;
      RECT 90.1850 219.1400 91.0550 219.6400 ;
      RECT 88.8050 219.1400 89.6750 219.6400 ;
      RECT 87.4250 219.1400 88.2950 219.6400 ;
      RECT 86.0450 219.1400 86.9150 219.6400 ;
      RECT 84.6650 219.1400 85.5350 219.6400 ;
      RECT 83.2850 219.1400 84.1550 219.6400 ;
      RECT 81.9050 219.1400 82.7750 219.6400 ;
      RECT 80.5250 219.1400 81.3950 219.6400 ;
      RECT 79.6050 219.1400 80.0150 219.6400 ;
      RECT 78.2250 219.1400 79.0950 219.6400 ;
      RECT 76.8450 219.1400 77.7150 219.6400 ;
      RECT 75.4650 219.1400 76.3350 219.6400 ;
      RECT 74.0850 219.1400 74.9550 219.6400 ;
      RECT 72.7050 219.1400 73.5750 219.6400 ;
      RECT 71.3250 219.1400 72.1950 219.6400 ;
      RECT 69.9450 219.1400 70.8150 219.6400 ;
      RECT 68.5650 219.1400 69.4350 219.6400 ;
      RECT 67.1850 219.1400 68.0550 219.6400 ;
      RECT 65.8050 219.1400 66.6750 219.6400 ;
      RECT 64.4250 219.1400 65.2950 219.6400 ;
      RECT 63.0450 219.1400 63.9150 219.6400 ;
      RECT 61.6650 219.1400 62.5350 219.6400 ;
      RECT 60.2850 219.1400 61.1550 219.6400 ;
      RECT 58.9050 219.1400 59.7750 219.6400 ;
      RECT 57.5250 219.1400 58.3950 219.6400 ;
      RECT 56.6050 219.1400 57.0150 219.6400 ;
      RECT 55.2250 219.1400 56.0950 219.6400 ;
      RECT 53.8450 219.1400 54.7150 219.6400 ;
      RECT 52.4650 219.1400 53.3350 219.6400 ;
      RECT 51.0850 219.1400 51.9550 219.6400 ;
      RECT 49.7050 219.1400 50.5750 219.6400 ;
      RECT 48.3250 219.1400 49.1950 219.6400 ;
      RECT 46.9450 219.1400 47.8150 219.6400 ;
      RECT 45.5650 219.1400 46.4350 219.6400 ;
      RECT 44.1850 219.1400 45.0550 219.6400 ;
      RECT 42.8050 219.1400 43.6750 219.6400 ;
      RECT 41.4250 219.1400 42.2950 219.6400 ;
      RECT 40.0450 219.1400 40.9150 219.6400 ;
      RECT 38.6650 219.1400 39.5350 219.6400 ;
      RECT 37.2850 219.1400 38.1550 219.6400 ;
      RECT 35.9050 219.1400 36.7750 219.6400 ;
      RECT 34.5250 219.1400 35.3950 219.6400 ;
      RECT 33.6050 219.1400 34.0150 219.6400 ;
      RECT 32.2250 219.1400 33.0950 219.6400 ;
      RECT 30.8450 219.1400 31.7150 219.6400 ;
      RECT 29.4650 219.1400 30.3350 219.6400 ;
      RECT 28.0850 219.1400 28.9550 219.6400 ;
      RECT 26.7050 219.1400 27.5750 219.6400 ;
      RECT 25.3250 219.1400 26.1950 219.6400 ;
      RECT 23.9450 219.1400 24.8150 219.6400 ;
      RECT 22.5650 219.1400 23.4350 219.6400 ;
      RECT 21.1850 219.1400 22.0550 219.6400 ;
      RECT 19.8050 219.1400 20.6750 219.6400 ;
      RECT 18.4250 219.1400 19.2950 219.6400 ;
      RECT 17.0450 219.1400 17.9150 219.6400 ;
      RECT 15.6650 219.1400 16.5350 219.6400 ;
      RECT 14.2850 219.1400 15.1550 219.6400 ;
      RECT 12.9050 219.1400 13.7750 219.6400 ;
      RECT 11.5250 219.1400 12.3950 219.6400 ;
      RECT 10.6050 219.1400 11.0150 219.6400 ;
      RECT 0.0000 219.1400 10.0950 219.6400 ;
      RECT 0.0000 0.5000 210.2200 219.1400 ;
      RECT 149.5250 0.0000 210.2200 0.5000 ;
      RECT 148.6050 0.0000 149.0150 0.5000 ;
      RECT 147.2250 0.0000 148.0950 0.5000 ;
      RECT 145.8450 0.0000 146.7150 0.5000 ;
      RECT 144.4650 0.0000 145.3350 0.5000 ;
      RECT 143.0850 0.0000 143.9550 0.5000 ;
      RECT 141.7050 0.0000 142.5750 0.5000 ;
      RECT 140.3250 0.0000 141.1950 0.5000 ;
      RECT 138.9450 0.0000 139.8150 0.5000 ;
      RECT 137.5650 0.0000 138.4350 0.5000 ;
      RECT 136.1850 0.0000 137.0550 0.5000 ;
      RECT 134.8050 0.0000 135.6750 0.5000 ;
      RECT 133.4250 0.0000 134.2950 0.5000 ;
      RECT 132.0450 0.0000 132.9150 0.5000 ;
      RECT 130.6650 0.0000 131.5350 0.5000 ;
      RECT 129.2850 0.0000 130.1550 0.5000 ;
      RECT 127.9050 0.0000 128.7750 0.5000 ;
      RECT 126.5250 0.0000 127.3950 0.5000 ;
      RECT 125.6050 0.0000 126.0150 0.5000 ;
      RECT 124.2250 0.0000 125.0950 0.5000 ;
      RECT 122.8450 0.0000 123.7150 0.5000 ;
      RECT 121.4650 0.0000 122.3350 0.5000 ;
      RECT 120.0850 0.0000 120.9550 0.5000 ;
      RECT 118.7050 0.0000 119.5750 0.5000 ;
      RECT 117.3250 0.0000 118.1950 0.5000 ;
      RECT 115.9450 0.0000 116.8150 0.5000 ;
      RECT 114.5650 0.0000 115.4350 0.5000 ;
      RECT 113.1850 0.0000 114.0550 0.5000 ;
      RECT 111.8050 0.0000 112.6750 0.5000 ;
      RECT 110.4250 0.0000 111.2950 0.5000 ;
      RECT 109.0450 0.0000 109.9150 0.5000 ;
      RECT 107.6650 0.0000 108.5350 0.5000 ;
      RECT 106.2850 0.0000 107.1550 0.5000 ;
      RECT 104.9050 0.0000 105.7750 0.5000 ;
      RECT 103.5250 0.0000 104.3950 0.5000 ;
      RECT 102.6050 0.0000 103.0150 0.5000 ;
      RECT 101.2250 0.0000 102.0950 0.5000 ;
      RECT 99.8450 0.0000 100.7150 0.5000 ;
      RECT 98.4650 0.0000 99.3350 0.5000 ;
      RECT 97.0850 0.0000 97.9550 0.5000 ;
      RECT 95.7050 0.0000 96.5750 0.5000 ;
      RECT 94.3250 0.0000 95.1950 0.5000 ;
      RECT 92.9450 0.0000 93.8150 0.5000 ;
      RECT 91.5650 0.0000 92.4350 0.5000 ;
      RECT 90.1850 0.0000 91.0550 0.5000 ;
      RECT 88.8050 0.0000 89.6750 0.5000 ;
      RECT 87.4250 0.0000 88.2950 0.5000 ;
      RECT 86.0450 0.0000 86.9150 0.5000 ;
      RECT 84.6650 0.0000 85.5350 0.5000 ;
      RECT 83.2850 0.0000 84.1550 0.5000 ;
      RECT 81.9050 0.0000 82.7750 0.5000 ;
      RECT 80.5250 0.0000 81.3950 0.5000 ;
      RECT 79.6050 0.0000 80.0150 0.5000 ;
      RECT 78.2250 0.0000 79.0950 0.5000 ;
      RECT 76.8450 0.0000 77.7150 0.5000 ;
      RECT 75.4650 0.0000 76.3350 0.5000 ;
      RECT 74.0850 0.0000 74.9550 0.5000 ;
      RECT 72.7050 0.0000 73.5750 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 69.9450 0.0000 70.8150 0.5000 ;
      RECT 68.5650 0.0000 69.4350 0.5000 ;
      RECT 67.1850 0.0000 68.0550 0.5000 ;
      RECT 65.8050 0.0000 66.6750 0.5000 ;
      RECT 64.4250 0.0000 65.2950 0.5000 ;
      RECT 63.0450 0.0000 63.9150 0.5000 ;
      RECT 61.6650 0.0000 62.5350 0.5000 ;
      RECT 60.2850 0.0000 61.1550 0.5000 ;
      RECT 58.9050 0.0000 59.7750 0.5000 ;
      RECT 57.5250 0.0000 58.3950 0.5000 ;
      RECT 56.6050 0.0000 57.0150 0.5000 ;
      RECT 55.2250 0.0000 56.0950 0.5000 ;
      RECT 53.8450 0.0000 54.7150 0.5000 ;
      RECT 52.4650 0.0000 53.3350 0.5000 ;
      RECT 51.0850 0.0000 51.9550 0.5000 ;
      RECT 49.7050 0.0000 50.5750 0.5000 ;
      RECT 48.3250 0.0000 49.1950 0.5000 ;
      RECT 46.9450 0.0000 47.8150 0.5000 ;
      RECT 45.5650 0.0000 46.4350 0.5000 ;
      RECT 44.1850 0.0000 45.0550 0.5000 ;
      RECT 42.8050 0.0000 43.6750 0.5000 ;
      RECT 41.4250 0.0000 42.2950 0.5000 ;
      RECT 40.0450 0.0000 40.9150 0.5000 ;
      RECT 38.6650 0.0000 39.5350 0.5000 ;
      RECT 37.2850 0.0000 38.1550 0.5000 ;
      RECT 35.9050 0.0000 36.7750 0.5000 ;
      RECT 34.5250 0.0000 35.3950 0.5000 ;
      RECT 33.6050 0.0000 34.0150 0.5000 ;
      RECT 32.2250 0.0000 33.0950 0.5000 ;
      RECT 30.8450 0.0000 31.7150 0.5000 ;
      RECT 29.4650 0.0000 30.3350 0.5000 ;
      RECT 28.0850 0.0000 28.9550 0.5000 ;
      RECT 26.7050 0.0000 27.5750 0.5000 ;
      RECT 25.3250 0.0000 26.1950 0.5000 ;
      RECT 23.9450 0.0000 24.8150 0.5000 ;
      RECT 22.5650 0.0000 23.4350 0.5000 ;
      RECT 21.1850 0.0000 22.0550 0.5000 ;
      RECT 19.8050 0.0000 20.6750 0.5000 ;
      RECT 18.4250 0.0000 19.2950 0.5000 ;
      RECT 17.0450 0.0000 17.9150 0.5000 ;
      RECT 15.6650 0.0000 16.5350 0.5000 ;
      RECT 14.2850 0.0000 15.1550 0.5000 ;
      RECT 12.9050 0.0000 13.7750 0.5000 ;
      RECT 11.5250 0.0000 12.3950 0.5000 ;
      RECT 10.6050 0.0000 11.0150 0.5000 ;
      RECT 0.0000 0.0000 10.0950 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 210.2200 219.6400 ;
    LAYER met2 ;
      RECT 199.6200 219.0150 210.2200 219.6400 ;
      RECT 197.7800 219.0150 199.2000 219.6400 ;
      RECT 195.0200 219.0150 197.3600 219.6400 ;
      RECT 193.1800 219.0150 194.6000 219.6400 ;
      RECT 190.8800 219.0150 192.7600 219.6400 ;
      RECT 188.5800 219.0150 190.4600 219.6400 ;
      RECT 186.2800 219.0150 188.1600 219.6400 ;
      RECT 184.4400 219.0150 185.8600 219.6400 ;
      RECT 181.6800 219.0150 184.0200 219.6400 ;
      RECT 179.8400 219.0150 181.2600 219.6400 ;
      RECT 177.5400 219.0150 179.4200 219.6400 ;
      RECT 175.2400 219.0150 177.1200 219.6400 ;
      RECT 172.9400 219.0150 174.8200 219.6400 ;
      RECT 170.6400 219.0150 172.5200 219.6400 ;
      RECT 168.8000 219.0150 170.2200 219.6400 ;
      RECT 166.5000 219.0150 168.3800 219.6400 ;
      RECT 164.2000 219.0150 166.0800 219.6400 ;
      RECT 161.9000 219.0150 163.7800 219.6400 ;
      RECT 159.6000 219.0150 161.4800 219.6400 ;
      RECT 156.8400 219.0150 159.1800 219.6400 ;
      RECT 155.4600 219.0150 156.4200 219.6400 ;
      RECT 0.0000 219.0150 155.0400 219.6400 ;
      RECT 0.0000 209.8200 210.2200 219.0150 ;
      RECT 0.6250 209.4000 209.5950 209.8200 ;
      RECT 0.0000 208.1200 210.2200 209.4000 ;
      RECT 0.6250 207.7000 209.5950 208.1200 ;
      RECT 0.0000 206.4200 210.2200 207.7000 ;
      RECT 0.6250 206.0000 209.5950 206.4200 ;
      RECT 0.0000 204.7200 210.2200 206.0000 ;
      RECT 0.6250 204.3000 209.5950 204.7200 ;
      RECT 0.0000 203.0200 210.2200 204.3000 ;
      RECT 0.6250 202.6000 209.5950 203.0200 ;
      RECT 0.0000 201.3200 210.2200 202.6000 ;
      RECT 0.6250 200.9000 209.5950 201.3200 ;
      RECT 0.0000 199.2800 210.2200 200.9000 ;
      RECT 0.6250 198.8600 209.5950 199.2800 ;
      RECT 0.0000 197.5800 210.2200 198.8600 ;
      RECT 0.6250 197.1600 209.5950 197.5800 ;
      RECT 0.0000 195.8800 210.2200 197.1600 ;
      RECT 0.6250 195.4600 209.5950 195.8800 ;
      RECT 0.0000 194.1800 210.2200 195.4600 ;
      RECT 0.6250 193.7600 209.5950 194.1800 ;
      RECT 0.0000 192.4800 210.2200 193.7600 ;
      RECT 0.6250 192.0600 209.5950 192.4800 ;
      RECT 0.0000 190.4400 210.2200 192.0600 ;
      RECT 0.6250 190.0200 209.5950 190.4400 ;
      RECT 0.0000 188.7400 210.2200 190.0200 ;
      RECT 0.6250 188.3200 209.5950 188.7400 ;
      RECT 0.0000 187.0400 210.2200 188.3200 ;
      RECT 0.6250 186.6200 209.5950 187.0400 ;
      RECT 0.0000 185.3400 210.2200 186.6200 ;
      RECT 0.6250 184.9200 209.5950 185.3400 ;
      RECT 0.0000 183.6400 210.2200 184.9200 ;
      RECT 0.6250 183.2200 209.5950 183.6400 ;
      RECT 0.0000 181.6000 210.2200 183.2200 ;
      RECT 0.6250 181.1800 209.5950 181.6000 ;
      RECT 0.0000 179.9000 210.2200 181.1800 ;
      RECT 0.6250 179.4800 209.5950 179.9000 ;
      RECT 0.0000 178.2000 210.2200 179.4800 ;
      RECT 0.6250 177.7800 209.5950 178.2000 ;
      RECT 0.0000 176.5000 210.2200 177.7800 ;
      RECT 0.6250 176.0800 209.5950 176.5000 ;
      RECT 0.0000 174.8000 210.2200 176.0800 ;
      RECT 0.6250 174.3800 209.5950 174.8000 ;
      RECT 0.0000 172.7600 210.2200 174.3800 ;
      RECT 0.6250 172.3400 209.5950 172.7600 ;
      RECT 0.0000 171.0600 210.2200 172.3400 ;
      RECT 0.6250 170.6400 209.5950 171.0600 ;
      RECT 0.0000 169.3600 210.2200 170.6400 ;
      RECT 0.6250 168.9400 209.5950 169.3600 ;
      RECT 0.0000 167.6600 210.2200 168.9400 ;
      RECT 0.6250 167.2400 209.5950 167.6600 ;
      RECT 0.0000 165.9600 210.2200 167.2400 ;
      RECT 0.6250 165.5400 209.5950 165.9600 ;
      RECT 0.0000 163.9200 210.2200 165.5400 ;
      RECT 0.6250 163.5000 209.5950 163.9200 ;
      RECT 0.0000 162.2200 210.2200 163.5000 ;
      RECT 0.6250 161.8000 209.5950 162.2200 ;
      RECT 0.0000 160.5200 210.2200 161.8000 ;
      RECT 0.6250 160.1000 209.5950 160.5200 ;
      RECT 0.0000 158.8200 210.2200 160.1000 ;
      RECT 0.6250 158.4000 209.5950 158.8200 ;
      RECT 0.0000 157.1200 210.2200 158.4000 ;
      RECT 0.6250 156.7000 209.5950 157.1200 ;
      RECT 0.0000 155.4200 210.2200 156.7000 ;
      RECT 0.6250 155.0000 209.5950 155.4200 ;
      RECT 0.0000 149.9800 210.2200 155.0000 ;
      RECT 0.6250 149.5600 209.5950 149.9800 ;
      RECT 0.0000 148.2800 210.2200 149.5600 ;
      RECT 0.6250 147.8600 209.5950 148.2800 ;
      RECT 0.0000 146.9200 210.2200 147.8600 ;
      RECT 0.6250 146.5000 209.5950 146.9200 ;
      RECT 0.0000 145.5600 210.2200 146.5000 ;
      RECT 0.6250 145.1400 209.5950 145.5600 ;
      RECT 0.0000 143.8600 210.2200 145.1400 ;
      RECT 0.6250 143.4400 209.5950 143.8600 ;
      RECT 0.0000 142.5000 210.2200 143.4400 ;
      RECT 0.6250 142.0800 209.5950 142.5000 ;
      RECT 0.0000 141.1400 210.2200 142.0800 ;
      RECT 0.6250 140.7200 209.5950 141.1400 ;
      RECT 0.0000 139.4400 210.2200 140.7200 ;
      RECT 0.6250 139.0200 209.5950 139.4400 ;
      RECT 0.0000 138.0800 210.2200 139.0200 ;
      RECT 0.6250 137.6600 209.5950 138.0800 ;
      RECT 0.0000 136.7200 210.2200 137.6600 ;
      RECT 0.6250 136.3000 209.5950 136.7200 ;
      RECT 0.0000 135.0200 210.2200 136.3000 ;
      RECT 0.6250 134.6000 209.5950 135.0200 ;
      RECT 0.0000 133.6600 210.2200 134.6000 ;
      RECT 0.6250 133.2400 209.5950 133.6600 ;
      RECT 0.0000 132.3000 210.2200 133.2400 ;
      RECT 0.6250 131.8800 209.5950 132.3000 ;
      RECT 0.0000 130.6000 210.2200 131.8800 ;
      RECT 0.6250 130.1800 209.5950 130.6000 ;
      RECT 0.0000 129.2400 210.2200 130.1800 ;
      RECT 0.6250 128.8200 209.5950 129.2400 ;
      RECT 0.0000 127.8800 210.2200 128.8200 ;
      RECT 0.6250 127.4600 209.5950 127.8800 ;
      RECT 0.0000 126.1800 210.2200 127.4600 ;
      RECT 0.6250 125.7600 209.5950 126.1800 ;
      RECT 0.0000 124.8200 210.2200 125.7600 ;
      RECT 0.6250 124.4000 209.5950 124.8200 ;
      RECT 0.0000 123.4600 210.2200 124.4000 ;
      RECT 0.6250 123.0400 209.5950 123.4600 ;
      RECT 0.0000 121.7600 210.2200 123.0400 ;
      RECT 0.6250 121.3400 209.5950 121.7600 ;
      RECT 0.0000 120.4000 210.2200 121.3400 ;
      RECT 0.6250 119.9800 209.5950 120.4000 ;
      RECT 0.0000 119.0400 210.2200 119.9800 ;
      RECT 0.6250 118.6200 209.5950 119.0400 ;
      RECT 0.0000 117.3400 210.2200 118.6200 ;
      RECT 0.6250 116.9200 209.5950 117.3400 ;
      RECT 0.0000 115.9800 210.2200 116.9200 ;
      RECT 0.6250 115.5600 209.5950 115.9800 ;
      RECT 0.0000 114.6200 210.2200 115.5600 ;
      RECT 0.6250 114.2000 209.5950 114.6200 ;
      RECT 0.0000 112.9200 210.2200 114.2000 ;
      RECT 0.6250 112.5000 209.5950 112.9200 ;
      RECT 0.0000 111.5600 210.2200 112.5000 ;
      RECT 0.6250 111.1400 209.5950 111.5600 ;
      RECT 0.0000 110.2000 210.2200 111.1400 ;
      RECT 0.6250 109.7800 209.5950 110.2000 ;
      RECT 0.0000 108.5000 210.2200 109.7800 ;
      RECT 0.6250 108.0800 209.5950 108.5000 ;
      RECT 0.0000 107.1400 210.2200 108.0800 ;
      RECT 0.6250 106.7200 209.5950 107.1400 ;
      RECT 0.0000 105.7800 210.2200 106.7200 ;
      RECT 0.6250 105.3600 209.5950 105.7800 ;
      RECT 0.0000 104.0800 210.2200 105.3600 ;
      RECT 0.6250 103.6600 209.5950 104.0800 ;
      RECT 0.0000 102.7200 210.2200 103.6600 ;
      RECT 0.6250 102.3000 209.5950 102.7200 ;
      RECT 0.0000 101.3600 210.2200 102.3000 ;
      RECT 0.6250 100.9400 209.5950 101.3600 ;
      RECT 0.0000 99.6600 210.2200 100.9400 ;
      RECT 0.6250 99.2400 209.5950 99.6600 ;
      RECT 0.0000 98.3000 210.2200 99.2400 ;
      RECT 0.6250 97.8800 209.5950 98.3000 ;
      RECT 0.0000 96.9400 210.2200 97.8800 ;
      RECT 0.6250 96.5200 209.5950 96.9400 ;
      RECT 0.0000 95.2400 210.2200 96.5200 ;
      RECT 0.6250 94.8200 209.5950 95.2400 ;
      RECT 0.0000 93.8800 210.2200 94.8200 ;
      RECT 0.6250 93.4600 209.5950 93.8800 ;
      RECT 0.0000 92.5200 210.2200 93.4600 ;
      RECT 0.6250 92.1000 209.5950 92.5200 ;
      RECT 0.0000 90.8200 210.2200 92.1000 ;
      RECT 0.6250 90.4000 209.5950 90.8200 ;
      RECT 0.0000 89.4600 210.2200 90.4000 ;
      RECT 0.6250 89.0400 209.5950 89.4600 ;
      RECT 0.0000 88.1000 210.2200 89.0400 ;
      RECT 0.6250 87.6800 209.5950 88.1000 ;
      RECT 0.0000 86.4000 210.2200 87.6800 ;
      RECT 0.6250 85.9800 209.5950 86.4000 ;
      RECT 0.0000 85.0400 210.2200 85.9800 ;
      RECT 0.6250 84.6200 209.5950 85.0400 ;
      RECT 0.0000 83.6800 210.2200 84.6200 ;
      RECT 0.6250 83.2600 209.5950 83.6800 ;
      RECT 0.0000 81.9800 210.2200 83.2600 ;
      RECT 0.6250 81.5600 209.5950 81.9800 ;
      RECT 0.0000 80.6200 210.2200 81.5600 ;
      RECT 0.6250 80.2000 209.5950 80.6200 ;
      RECT 0.0000 79.2600 210.2200 80.2000 ;
      RECT 0.6250 78.8400 209.5950 79.2600 ;
      RECT 0.0000 77.9000 210.2200 78.8400 ;
      RECT 0.6250 77.4800 209.5950 77.9000 ;
      RECT 0.0000 76.2000 210.2200 77.4800 ;
      RECT 0.6250 75.7800 209.5950 76.2000 ;
      RECT 0.0000 74.8400 210.2200 75.7800 ;
      RECT 0.6250 74.4200 209.5950 74.8400 ;
      RECT 0.0000 73.4800 210.2200 74.4200 ;
      RECT 0.6250 73.0600 209.5950 73.4800 ;
      RECT 0.0000 71.7800 210.2200 73.0600 ;
      RECT 0.6250 71.3600 209.5950 71.7800 ;
      RECT 0.0000 70.4200 210.2200 71.3600 ;
      RECT 0.6250 70.0000 209.5950 70.4200 ;
      RECT 0.0000 69.0600 210.2200 70.0000 ;
      RECT 0.6250 68.6400 209.5950 69.0600 ;
      RECT 0.0000 67.3600 210.2200 68.6400 ;
      RECT 0.6250 66.9400 209.5950 67.3600 ;
      RECT 0.0000 66.0000 210.2200 66.9400 ;
      RECT 0.6250 65.5800 209.5950 66.0000 ;
      RECT 0.0000 64.6400 210.2200 65.5800 ;
      RECT 0.6250 64.2200 209.5950 64.6400 ;
      RECT 0.0000 62.9400 210.2200 64.2200 ;
      RECT 0.6250 62.5200 209.5950 62.9400 ;
      RECT 0.0000 61.5800 210.2200 62.5200 ;
      RECT 0.6250 61.1600 209.5950 61.5800 ;
      RECT 0.0000 60.2200 210.2200 61.1600 ;
      RECT 0.6250 59.8000 209.5950 60.2200 ;
      RECT 0.0000 58.5200 210.2200 59.8000 ;
      RECT 0.6250 58.1000 209.5950 58.5200 ;
      RECT 0.0000 57.1600 210.2200 58.1000 ;
      RECT 0.6250 56.7400 209.5950 57.1600 ;
      RECT 0.0000 55.8000 210.2200 56.7400 ;
      RECT 0.6250 55.3800 209.5950 55.8000 ;
      RECT 0.0000 54.1000 210.2200 55.3800 ;
      RECT 0.6250 53.6800 209.5950 54.1000 ;
      RECT 0.0000 52.7400 210.2200 53.6800 ;
      RECT 0.6250 52.3200 209.5950 52.7400 ;
      RECT 0.0000 51.3800 210.2200 52.3200 ;
      RECT 0.6250 50.9600 209.5950 51.3800 ;
      RECT 0.0000 49.6800 210.2200 50.9600 ;
      RECT 0.6250 49.2600 209.5950 49.6800 ;
      RECT 0.0000 48.3200 210.2200 49.2600 ;
      RECT 0.6250 47.9000 209.5950 48.3200 ;
      RECT 0.0000 46.9600 210.2200 47.9000 ;
      RECT 0.6250 46.5400 209.5950 46.9600 ;
      RECT 0.0000 45.2600 210.2200 46.5400 ;
      RECT 0.6250 44.8400 209.5950 45.2600 ;
      RECT 0.0000 43.9000 210.2200 44.8400 ;
      RECT 0.6250 43.4800 209.5950 43.9000 ;
      RECT 0.0000 42.5400 210.2200 43.4800 ;
      RECT 0.6250 42.1200 209.5950 42.5400 ;
      RECT 0.0000 40.8400 210.2200 42.1200 ;
      RECT 0.6250 40.4200 209.5950 40.8400 ;
      RECT 0.0000 39.4800 210.2200 40.4200 ;
      RECT 0.6250 39.0600 209.5950 39.4800 ;
      RECT 0.0000 38.1200 210.2200 39.0600 ;
      RECT 0.6250 37.7000 209.5950 38.1200 ;
      RECT 0.0000 36.4200 210.2200 37.7000 ;
      RECT 0.6250 36.0000 209.5950 36.4200 ;
      RECT 0.0000 35.0600 210.2200 36.0000 ;
      RECT 0.6250 34.6400 209.5950 35.0600 ;
      RECT 0.0000 33.7000 210.2200 34.6400 ;
      RECT 0.6250 33.2800 209.5950 33.7000 ;
      RECT 0.0000 32.0000 210.2200 33.2800 ;
      RECT 0.6250 31.5800 209.5950 32.0000 ;
      RECT 0.0000 30.6400 210.2200 31.5800 ;
      RECT 0.6250 30.2200 209.5950 30.6400 ;
      RECT 0.0000 29.2800 210.2200 30.2200 ;
      RECT 0.6250 28.8600 209.5950 29.2800 ;
      RECT 0.0000 27.5800 210.2200 28.8600 ;
      RECT 0.6250 27.1600 209.5950 27.5800 ;
      RECT 0.0000 26.2200 210.2200 27.1600 ;
      RECT 0.6250 25.8000 209.5950 26.2200 ;
      RECT 0.0000 24.8600 210.2200 25.8000 ;
      RECT 0.6250 24.4400 209.5950 24.8600 ;
      RECT 0.0000 23.1600 210.2200 24.4400 ;
      RECT 0.6250 22.7400 209.5950 23.1600 ;
      RECT 0.0000 21.8000 210.2200 22.7400 ;
      RECT 0.6250 21.3800 209.5950 21.8000 ;
      RECT 0.0000 20.4400 210.2200 21.3800 ;
      RECT 0.6250 20.0200 209.5950 20.4400 ;
      RECT 0.0000 18.7400 210.2200 20.0200 ;
      RECT 0.6250 18.3200 209.5950 18.7400 ;
      RECT 0.0000 17.3800 210.2200 18.3200 ;
      RECT 0.6250 16.9600 209.5950 17.3800 ;
      RECT 0.0000 16.0200 210.2200 16.9600 ;
      RECT 0.6250 15.6000 209.5950 16.0200 ;
      RECT 0.0000 14.3200 210.2200 15.6000 ;
      RECT 0.6250 13.9000 209.5950 14.3200 ;
      RECT 0.0000 12.9600 210.2200 13.9000 ;
      RECT 0.6250 12.5400 209.5950 12.9600 ;
      RECT 0.0000 11.6000 210.2200 12.5400 ;
      RECT 0.6250 11.1800 209.5950 11.6000 ;
      RECT 0.0000 10.2400 210.2200 11.1800 ;
      RECT 0.6250 9.8200 209.5950 10.2400 ;
      RECT 0.0000 0.6250 210.2200 9.8200 ;
      RECT 199.6200 0.0000 210.2200 0.6250 ;
      RECT 197.7800 0.0000 199.2000 0.6250 ;
      RECT 195.4800 0.0000 197.3600 0.6250 ;
      RECT 193.1800 0.0000 195.0600 0.6250 ;
      RECT 190.8800 0.0000 192.7600 0.6250 ;
      RECT 188.5800 0.0000 190.4600 0.6250 ;
      RECT 185.8200 0.0000 188.1600 0.6250 ;
      RECT 184.4400 0.0000 185.4000 0.6250 ;
      RECT 181.6800 0.0000 184.0200 0.6250 ;
      RECT 179.8400 0.0000 181.2600 0.6250 ;
      RECT 177.5400 0.0000 179.4200 0.6250 ;
      RECT 175.2400 0.0000 177.1200 0.6250 ;
      RECT 172.9400 0.0000 174.8200 0.6250 ;
      RECT 170.6400 0.0000 172.5200 0.6250 ;
      RECT 168.8000 0.0000 170.2200 0.6250 ;
      RECT 166.5000 0.0000 168.3800 0.6250 ;
      RECT 164.2000 0.0000 166.0800 0.6250 ;
      RECT 161.4400 0.0000 163.7800 0.6250 ;
      RECT 159.6000 0.0000 161.0200 0.6250 ;
      RECT 157.3000 0.0000 159.1800 0.6250 ;
      RECT 155.4600 0.0000 156.8800 0.6250 ;
      RECT 0.0000 0.0000 155.0400 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 217.8300 210.2200 219.6400 ;
      RECT 208.9600 214.2300 210.2200 217.8300 ;
      RECT 0.0000 214.2300 1.2600 217.8300 ;
      RECT 0.0000 213.8300 210.2200 214.2300 ;
      RECT 204.9600 210.2300 210.2200 213.8300 ;
      RECT 0.0000 210.2300 5.2600 213.8300 ;
      RECT 0.0000 208.9600 210.2200 210.2300 ;
      RECT 204.9600 207.8800 210.2200 208.9600 ;
      RECT 192.0200 207.8800 201.3600 208.9600 ;
      RECT 147.0200 207.8800 189.8200 208.9600 ;
      RECT 102.0200 207.8800 144.8200 208.9600 ;
      RECT 57.0200 207.8800 99.8200 208.9600 ;
      RECT 8.8600 207.8800 54.8200 208.9600 ;
      RECT 0.0000 207.8800 5.2600 208.9600 ;
      RECT 0.0000 206.2400 210.2200 207.8800 ;
      RECT 208.9600 205.1600 210.2200 206.2400 ;
      RECT 195.2200 205.1600 205.3600 206.2400 ;
      RECT 150.2200 205.1600 193.0200 206.2400 ;
      RECT 105.2200 205.1600 148.0200 206.2400 ;
      RECT 60.2200 205.1600 103.0200 206.2400 ;
      RECT 15.2200 205.1600 58.0200 206.2400 ;
      RECT 4.8600 205.1600 13.0200 206.2400 ;
      RECT 0.0000 205.1600 1.2600 206.2400 ;
      RECT 0.0000 203.5200 210.2200 205.1600 ;
      RECT 204.9600 202.4400 210.2200 203.5200 ;
      RECT 192.0200 202.4400 201.3600 203.5200 ;
      RECT 147.0200 202.4400 189.8200 203.5200 ;
      RECT 102.0200 202.4400 144.8200 203.5200 ;
      RECT 57.0200 202.4400 99.8200 203.5200 ;
      RECT 8.8600 202.4400 54.8200 203.5200 ;
      RECT 0.0000 202.4400 5.2600 203.5200 ;
      RECT 0.0000 200.8000 210.2200 202.4400 ;
      RECT 208.9600 199.7200 210.2200 200.8000 ;
      RECT 195.2200 199.7200 205.3600 200.8000 ;
      RECT 150.2200 199.7200 193.0200 200.8000 ;
      RECT 105.2200 199.7200 148.0200 200.8000 ;
      RECT 60.2200 199.7200 103.0200 200.8000 ;
      RECT 15.2200 199.7200 58.0200 200.8000 ;
      RECT 4.8600 199.7200 13.0200 200.8000 ;
      RECT 0.0000 199.7200 1.2600 200.8000 ;
      RECT 0.0000 198.0800 210.2200 199.7200 ;
      RECT 204.9600 197.0000 210.2200 198.0800 ;
      RECT 192.0200 197.0000 201.3600 198.0800 ;
      RECT 147.0200 197.0000 189.8200 198.0800 ;
      RECT 102.0200 197.0000 144.8200 198.0800 ;
      RECT 57.0200 197.0000 99.8200 198.0800 ;
      RECT 8.8600 197.0000 54.8200 198.0800 ;
      RECT 0.0000 197.0000 5.2600 198.0800 ;
      RECT 0.0000 195.3600 210.2200 197.0000 ;
      RECT 208.9600 194.2800 210.2200 195.3600 ;
      RECT 195.2200 194.2800 205.3600 195.3600 ;
      RECT 150.2200 194.2800 193.0200 195.3600 ;
      RECT 105.2200 194.2800 148.0200 195.3600 ;
      RECT 60.2200 194.2800 103.0200 195.3600 ;
      RECT 15.2200 194.2800 58.0200 195.3600 ;
      RECT 4.8600 194.2800 13.0200 195.3600 ;
      RECT 0.0000 194.2800 1.2600 195.3600 ;
      RECT 0.0000 192.6400 210.2200 194.2800 ;
      RECT 204.9600 191.5600 210.2200 192.6400 ;
      RECT 192.0200 191.5600 201.3600 192.6400 ;
      RECT 147.0200 191.5600 189.8200 192.6400 ;
      RECT 102.0200 191.5600 144.8200 192.6400 ;
      RECT 57.0200 191.5600 99.8200 192.6400 ;
      RECT 8.8600 191.5600 54.8200 192.6400 ;
      RECT 0.0000 191.5600 5.2600 192.6400 ;
      RECT 0.0000 189.9200 210.2200 191.5600 ;
      RECT 208.9600 188.8400 210.2200 189.9200 ;
      RECT 195.2200 188.8400 205.3600 189.9200 ;
      RECT 150.2200 188.8400 193.0200 189.9200 ;
      RECT 105.2200 188.8400 148.0200 189.9200 ;
      RECT 60.2200 188.8400 103.0200 189.9200 ;
      RECT 15.2200 188.8400 58.0200 189.9200 ;
      RECT 4.8600 188.8400 13.0200 189.9200 ;
      RECT 0.0000 188.8400 1.2600 189.9200 ;
      RECT 0.0000 187.2000 210.2200 188.8400 ;
      RECT 204.9600 186.1200 210.2200 187.2000 ;
      RECT 192.0200 186.1200 201.3600 187.2000 ;
      RECT 147.0200 186.1200 189.8200 187.2000 ;
      RECT 102.0200 186.1200 144.8200 187.2000 ;
      RECT 57.0200 186.1200 99.8200 187.2000 ;
      RECT 8.8600 186.1200 54.8200 187.2000 ;
      RECT 0.0000 186.1200 5.2600 187.2000 ;
      RECT 0.0000 184.4800 210.2200 186.1200 ;
      RECT 208.9600 183.4000 210.2200 184.4800 ;
      RECT 195.2200 183.4000 205.3600 184.4800 ;
      RECT 150.2200 183.4000 193.0200 184.4800 ;
      RECT 105.2200 183.4000 148.0200 184.4800 ;
      RECT 60.2200 183.4000 103.0200 184.4800 ;
      RECT 15.2200 183.4000 58.0200 184.4800 ;
      RECT 4.8600 183.4000 13.0200 184.4800 ;
      RECT 0.0000 183.4000 1.2600 184.4800 ;
      RECT 0.0000 181.7600 210.2200 183.4000 ;
      RECT 204.9600 180.6800 210.2200 181.7600 ;
      RECT 192.0200 180.6800 201.3600 181.7600 ;
      RECT 147.0200 180.6800 189.8200 181.7600 ;
      RECT 102.0200 180.6800 144.8200 181.7600 ;
      RECT 57.0200 180.6800 99.8200 181.7600 ;
      RECT 8.8600 180.6800 54.8200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 181.7600 ;
      RECT 0.0000 179.0400 210.2200 180.6800 ;
      RECT 208.9600 177.9600 210.2200 179.0400 ;
      RECT 195.2200 177.9600 205.3600 179.0400 ;
      RECT 150.2200 177.9600 193.0200 179.0400 ;
      RECT 105.2200 177.9600 148.0200 179.0400 ;
      RECT 60.2200 177.9600 103.0200 179.0400 ;
      RECT 15.2200 177.9600 58.0200 179.0400 ;
      RECT 4.8600 177.9600 13.0200 179.0400 ;
      RECT 0.0000 177.9600 1.2600 179.0400 ;
      RECT 0.0000 176.3200 210.2200 177.9600 ;
      RECT 204.9600 175.2400 210.2200 176.3200 ;
      RECT 192.0200 175.2400 201.3600 176.3200 ;
      RECT 147.0200 175.2400 189.8200 176.3200 ;
      RECT 102.0200 175.2400 144.8200 176.3200 ;
      RECT 57.0200 175.2400 99.8200 176.3200 ;
      RECT 8.8600 175.2400 54.8200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 176.3200 ;
      RECT 0.0000 173.6000 210.2200 175.2400 ;
      RECT 208.9600 172.5200 210.2200 173.6000 ;
      RECT 195.2200 172.5200 205.3600 173.6000 ;
      RECT 150.2200 172.5200 193.0200 173.6000 ;
      RECT 105.2200 172.5200 148.0200 173.6000 ;
      RECT 60.2200 172.5200 103.0200 173.6000 ;
      RECT 15.2200 172.5200 58.0200 173.6000 ;
      RECT 4.8600 172.5200 13.0200 173.6000 ;
      RECT 0.0000 172.5200 1.2600 173.6000 ;
      RECT 0.0000 170.8800 210.2200 172.5200 ;
      RECT 204.9600 169.8000 210.2200 170.8800 ;
      RECT 192.0200 169.8000 201.3600 170.8800 ;
      RECT 147.0200 169.8000 189.8200 170.8800 ;
      RECT 102.0200 169.8000 144.8200 170.8800 ;
      RECT 57.0200 169.8000 99.8200 170.8800 ;
      RECT 8.8600 169.8000 54.8200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.8800 ;
      RECT 0.0000 168.1600 210.2200 169.8000 ;
      RECT 208.9600 167.0800 210.2200 168.1600 ;
      RECT 195.2200 167.0800 205.3600 168.1600 ;
      RECT 150.2200 167.0800 193.0200 168.1600 ;
      RECT 105.2200 167.0800 148.0200 168.1600 ;
      RECT 60.2200 167.0800 103.0200 168.1600 ;
      RECT 15.2200 167.0800 58.0200 168.1600 ;
      RECT 4.8600 167.0800 13.0200 168.1600 ;
      RECT 0.0000 167.0800 1.2600 168.1600 ;
      RECT 0.0000 165.4400 210.2200 167.0800 ;
      RECT 204.9600 164.3600 210.2200 165.4400 ;
      RECT 192.0200 164.3600 201.3600 165.4400 ;
      RECT 147.0200 164.3600 189.8200 165.4400 ;
      RECT 102.0200 164.3600 144.8200 165.4400 ;
      RECT 57.0200 164.3600 99.8200 165.4400 ;
      RECT 8.8600 164.3600 54.8200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.4400 ;
      RECT 0.0000 162.7200 210.2200 164.3600 ;
      RECT 208.9600 161.6400 210.2200 162.7200 ;
      RECT 195.2200 161.6400 205.3600 162.7200 ;
      RECT 150.2200 161.6400 193.0200 162.7200 ;
      RECT 105.2200 161.6400 148.0200 162.7200 ;
      RECT 60.2200 161.6400 103.0200 162.7200 ;
      RECT 15.2200 161.6400 58.0200 162.7200 ;
      RECT 4.8600 161.6400 13.0200 162.7200 ;
      RECT 0.0000 161.6400 1.2600 162.7200 ;
      RECT 0.0000 160.0000 210.2200 161.6400 ;
      RECT 204.9600 158.9200 210.2200 160.0000 ;
      RECT 192.0200 158.9200 201.3600 160.0000 ;
      RECT 147.0200 158.9200 189.8200 160.0000 ;
      RECT 102.0200 158.9200 144.8200 160.0000 ;
      RECT 57.0200 158.9200 99.8200 160.0000 ;
      RECT 8.8600 158.9200 54.8200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 160.0000 ;
      RECT 0.0000 157.2800 210.2200 158.9200 ;
      RECT 208.9600 156.2000 210.2200 157.2800 ;
      RECT 195.2200 156.2000 205.3600 157.2800 ;
      RECT 150.2200 156.2000 193.0200 157.2800 ;
      RECT 105.2200 156.2000 148.0200 157.2800 ;
      RECT 60.2200 156.2000 103.0200 157.2800 ;
      RECT 15.2200 156.2000 58.0200 157.2800 ;
      RECT 4.8600 156.2000 13.0200 157.2800 ;
      RECT 0.0000 156.2000 1.2600 157.2800 ;
      RECT 0.0000 154.5600 210.2200 156.2000 ;
      RECT 204.9600 153.4800 210.2200 154.5600 ;
      RECT 192.0200 153.4800 201.3600 154.5600 ;
      RECT 147.0200 153.4800 189.8200 154.5600 ;
      RECT 102.0200 153.4800 144.8200 154.5600 ;
      RECT 57.0200 153.4800 99.8200 154.5600 ;
      RECT 8.8600 153.4800 54.8200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 210.2200 153.4800 ;
      RECT 208.9600 150.7600 210.2200 151.8400 ;
      RECT 195.2200 150.7600 205.3600 151.8400 ;
      RECT 150.2200 150.7600 193.0200 151.8400 ;
      RECT 105.2200 150.7600 148.0200 151.8400 ;
      RECT 60.2200 150.7600 103.0200 151.8400 ;
      RECT 15.2200 150.7600 58.0200 151.8400 ;
      RECT 4.8600 150.7600 13.0200 151.8400 ;
      RECT 0.0000 150.7600 1.2600 151.8400 ;
      RECT 0.0000 149.1200 210.2200 150.7600 ;
      RECT 204.9600 148.0400 210.2200 149.1200 ;
      RECT 192.0200 148.0400 201.3600 149.1200 ;
      RECT 147.0200 148.0400 189.8200 149.1200 ;
      RECT 102.0200 148.0400 144.8200 149.1200 ;
      RECT 57.0200 148.0400 99.8200 149.1200 ;
      RECT 8.8600 148.0400 54.8200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 210.2200 148.0400 ;
      RECT 208.9600 145.3200 210.2200 146.4000 ;
      RECT 195.2200 145.3200 205.3600 146.4000 ;
      RECT 150.2200 145.3200 193.0200 146.4000 ;
      RECT 105.2200 145.3200 148.0200 146.4000 ;
      RECT 60.2200 145.3200 103.0200 146.4000 ;
      RECT 15.2200 145.3200 58.0200 146.4000 ;
      RECT 4.8600 145.3200 13.0200 146.4000 ;
      RECT 0.0000 145.3200 1.2600 146.4000 ;
      RECT 0.0000 143.6800 210.2200 145.3200 ;
      RECT 204.9600 142.6000 210.2200 143.6800 ;
      RECT 192.0200 142.6000 201.3600 143.6800 ;
      RECT 147.0200 142.6000 189.8200 143.6800 ;
      RECT 102.0200 142.6000 144.8200 143.6800 ;
      RECT 57.0200 142.6000 99.8200 143.6800 ;
      RECT 8.8600 142.6000 54.8200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 210.2200 142.6000 ;
      RECT 208.9600 139.8800 210.2200 140.9600 ;
      RECT 195.2200 139.8800 205.3600 140.9600 ;
      RECT 150.2200 139.8800 193.0200 140.9600 ;
      RECT 105.2200 139.8800 148.0200 140.9600 ;
      RECT 60.2200 139.8800 103.0200 140.9600 ;
      RECT 15.2200 139.8800 58.0200 140.9600 ;
      RECT 4.8600 139.8800 13.0200 140.9600 ;
      RECT 0.0000 139.8800 1.2600 140.9600 ;
      RECT 0.0000 138.2400 210.2200 139.8800 ;
      RECT 204.9600 137.1600 210.2200 138.2400 ;
      RECT 192.0200 137.1600 201.3600 138.2400 ;
      RECT 147.0200 137.1600 189.8200 138.2400 ;
      RECT 102.0200 137.1600 144.8200 138.2400 ;
      RECT 57.0200 137.1600 99.8200 138.2400 ;
      RECT 8.8600 137.1600 54.8200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 210.2200 137.1600 ;
      RECT 208.9600 134.4400 210.2200 135.5200 ;
      RECT 195.2200 134.4400 205.3600 135.5200 ;
      RECT 150.2200 134.4400 193.0200 135.5200 ;
      RECT 105.2200 134.4400 148.0200 135.5200 ;
      RECT 60.2200 134.4400 103.0200 135.5200 ;
      RECT 15.2200 134.4400 58.0200 135.5200 ;
      RECT 4.8600 134.4400 13.0200 135.5200 ;
      RECT 0.0000 134.4400 1.2600 135.5200 ;
      RECT 0.0000 132.8000 210.2200 134.4400 ;
      RECT 204.9600 131.7200 210.2200 132.8000 ;
      RECT 192.0200 131.7200 201.3600 132.8000 ;
      RECT 147.0200 131.7200 189.8200 132.8000 ;
      RECT 102.0200 131.7200 144.8200 132.8000 ;
      RECT 57.0200 131.7200 99.8200 132.8000 ;
      RECT 8.8600 131.7200 54.8200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 210.2200 131.7200 ;
      RECT 208.9600 129.0000 210.2200 130.0800 ;
      RECT 195.2200 129.0000 205.3600 130.0800 ;
      RECT 150.2200 129.0000 193.0200 130.0800 ;
      RECT 105.2200 129.0000 148.0200 130.0800 ;
      RECT 60.2200 129.0000 103.0200 130.0800 ;
      RECT 15.2200 129.0000 58.0200 130.0800 ;
      RECT 4.8600 129.0000 13.0200 130.0800 ;
      RECT 0.0000 129.0000 1.2600 130.0800 ;
      RECT 0.0000 127.3600 210.2200 129.0000 ;
      RECT 204.9600 126.2800 210.2200 127.3600 ;
      RECT 192.0200 126.2800 201.3600 127.3600 ;
      RECT 147.0200 126.2800 189.8200 127.3600 ;
      RECT 102.0200 126.2800 144.8200 127.3600 ;
      RECT 57.0200 126.2800 99.8200 127.3600 ;
      RECT 8.8600 126.2800 54.8200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 210.2200 126.2800 ;
      RECT 208.9600 123.5600 210.2200 124.6400 ;
      RECT 195.2200 123.5600 205.3600 124.6400 ;
      RECT 150.2200 123.5600 193.0200 124.6400 ;
      RECT 105.2200 123.5600 148.0200 124.6400 ;
      RECT 60.2200 123.5600 103.0200 124.6400 ;
      RECT 15.2200 123.5600 58.0200 124.6400 ;
      RECT 4.8600 123.5600 13.0200 124.6400 ;
      RECT 0.0000 123.5600 1.2600 124.6400 ;
      RECT 0.0000 121.9200 210.2200 123.5600 ;
      RECT 204.9600 120.8400 210.2200 121.9200 ;
      RECT 192.0200 120.8400 201.3600 121.9200 ;
      RECT 147.0200 120.8400 189.8200 121.9200 ;
      RECT 102.0200 120.8400 144.8200 121.9200 ;
      RECT 57.0200 120.8400 99.8200 121.9200 ;
      RECT 8.8600 120.8400 54.8200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 210.2200 120.8400 ;
      RECT 208.9600 118.1200 210.2200 119.2000 ;
      RECT 195.2200 118.1200 205.3600 119.2000 ;
      RECT 150.2200 118.1200 193.0200 119.2000 ;
      RECT 105.2200 118.1200 148.0200 119.2000 ;
      RECT 60.2200 118.1200 103.0200 119.2000 ;
      RECT 15.2200 118.1200 58.0200 119.2000 ;
      RECT 4.8600 118.1200 13.0200 119.2000 ;
      RECT 0.0000 118.1200 1.2600 119.2000 ;
      RECT 0.0000 116.4800 210.2200 118.1200 ;
      RECT 204.9600 115.4000 210.2200 116.4800 ;
      RECT 192.0200 115.4000 201.3600 116.4800 ;
      RECT 147.0200 115.4000 189.8200 116.4800 ;
      RECT 102.0200 115.4000 144.8200 116.4800 ;
      RECT 57.0200 115.4000 99.8200 116.4800 ;
      RECT 8.8600 115.4000 54.8200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 210.2200 115.4000 ;
      RECT 208.9600 112.6800 210.2200 113.7600 ;
      RECT 195.2200 112.6800 205.3600 113.7600 ;
      RECT 150.2200 112.6800 193.0200 113.7600 ;
      RECT 105.2200 112.6800 148.0200 113.7600 ;
      RECT 60.2200 112.6800 103.0200 113.7600 ;
      RECT 15.2200 112.6800 58.0200 113.7600 ;
      RECT 4.8600 112.6800 13.0200 113.7600 ;
      RECT 0.0000 112.6800 1.2600 113.7600 ;
      RECT 0.0000 111.0400 210.2200 112.6800 ;
      RECT 204.9600 109.9600 210.2200 111.0400 ;
      RECT 192.0200 109.9600 201.3600 111.0400 ;
      RECT 147.0200 109.9600 189.8200 111.0400 ;
      RECT 102.0200 109.9600 144.8200 111.0400 ;
      RECT 57.0200 109.9600 99.8200 111.0400 ;
      RECT 8.8600 109.9600 54.8200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 210.2200 109.9600 ;
      RECT 208.9600 107.2400 210.2200 108.3200 ;
      RECT 195.2200 107.2400 205.3600 108.3200 ;
      RECT 150.2200 107.2400 193.0200 108.3200 ;
      RECT 105.2200 107.2400 148.0200 108.3200 ;
      RECT 60.2200 107.2400 103.0200 108.3200 ;
      RECT 15.2200 107.2400 58.0200 108.3200 ;
      RECT 4.8600 107.2400 13.0200 108.3200 ;
      RECT 0.0000 107.2400 1.2600 108.3200 ;
      RECT 0.0000 105.6000 210.2200 107.2400 ;
      RECT 204.9600 104.5200 210.2200 105.6000 ;
      RECT 192.0200 104.5200 201.3600 105.6000 ;
      RECT 147.0200 104.5200 189.8200 105.6000 ;
      RECT 102.0200 104.5200 144.8200 105.6000 ;
      RECT 57.0200 104.5200 99.8200 105.6000 ;
      RECT 8.8600 104.5200 54.8200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 210.2200 104.5200 ;
      RECT 208.9600 101.8000 210.2200 102.8800 ;
      RECT 195.2200 101.8000 205.3600 102.8800 ;
      RECT 150.2200 101.8000 193.0200 102.8800 ;
      RECT 105.2200 101.8000 148.0200 102.8800 ;
      RECT 60.2200 101.8000 103.0200 102.8800 ;
      RECT 15.2200 101.8000 58.0200 102.8800 ;
      RECT 4.8600 101.8000 13.0200 102.8800 ;
      RECT 0.0000 101.8000 1.2600 102.8800 ;
      RECT 0.0000 100.1600 210.2200 101.8000 ;
      RECT 204.9600 99.0800 210.2200 100.1600 ;
      RECT 192.0200 99.0800 201.3600 100.1600 ;
      RECT 147.0200 99.0800 189.8200 100.1600 ;
      RECT 102.0200 99.0800 144.8200 100.1600 ;
      RECT 57.0200 99.0800 99.8200 100.1600 ;
      RECT 8.8600 99.0800 54.8200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 210.2200 99.0800 ;
      RECT 208.9600 96.3600 210.2200 97.4400 ;
      RECT 195.2200 96.3600 205.3600 97.4400 ;
      RECT 150.2200 96.3600 193.0200 97.4400 ;
      RECT 105.2200 96.3600 148.0200 97.4400 ;
      RECT 60.2200 96.3600 103.0200 97.4400 ;
      RECT 15.2200 96.3600 58.0200 97.4400 ;
      RECT 4.8600 96.3600 13.0200 97.4400 ;
      RECT 0.0000 96.3600 1.2600 97.4400 ;
      RECT 0.0000 94.7200 210.2200 96.3600 ;
      RECT 204.9600 93.6400 210.2200 94.7200 ;
      RECT 192.0200 93.6400 201.3600 94.7200 ;
      RECT 147.0200 93.6400 189.8200 94.7200 ;
      RECT 102.0200 93.6400 144.8200 94.7200 ;
      RECT 57.0200 93.6400 99.8200 94.7200 ;
      RECT 8.8600 93.6400 54.8200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 210.2200 93.6400 ;
      RECT 208.9600 90.9200 210.2200 92.0000 ;
      RECT 195.2200 90.9200 205.3600 92.0000 ;
      RECT 150.2200 90.9200 193.0200 92.0000 ;
      RECT 105.2200 90.9200 148.0200 92.0000 ;
      RECT 60.2200 90.9200 103.0200 92.0000 ;
      RECT 15.2200 90.9200 58.0200 92.0000 ;
      RECT 4.8600 90.9200 13.0200 92.0000 ;
      RECT 0.0000 90.9200 1.2600 92.0000 ;
      RECT 0.0000 89.2800 210.2200 90.9200 ;
      RECT 204.9600 88.2000 210.2200 89.2800 ;
      RECT 192.0200 88.2000 201.3600 89.2800 ;
      RECT 147.0200 88.2000 189.8200 89.2800 ;
      RECT 102.0200 88.2000 144.8200 89.2800 ;
      RECT 57.0200 88.2000 99.8200 89.2800 ;
      RECT 8.8600 88.2000 54.8200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 210.2200 88.2000 ;
      RECT 208.9600 85.4800 210.2200 86.5600 ;
      RECT 195.2200 85.4800 205.3600 86.5600 ;
      RECT 150.2200 85.4800 193.0200 86.5600 ;
      RECT 105.2200 85.4800 148.0200 86.5600 ;
      RECT 60.2200 85.4800 103.0200 86.5600 ;
      RECT 15.2200 85.4800 58.0200 86.5600 ;
      RECT 4.8600 85.4800 13.0200 86.5600 ;
      RECT 0.0000 85.4800 1.2600 86.5600 ;
      RECT 0.0000 83.8400 210.2200 85.4800 ;
      RECT 204.9600 82.7600 210.2200 83.8400 ;
      RECT 192.0200 82.7600 201.3600 83.8400 ;
      RECT 147.0200 82.7600 189.8200 83.8400 ;
      RECT 102.0200 82.7600 144.8200 83.8400 ;
      RECT 57.0200 82.7600 99.8200 83.8400 ;
      RECT 8.8600 82.7600 54.8200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 210.2200 82.7600 ;
      RECT 208.9600 80.0400 210.2200 81.1200 ;
      RECT 195.2200 80.0400 205.3600 81.1200 ;
      RECT 150.2200 80.0400 193.0200 81.1200 ;
      RECT 105.2200 80.0400 148.0200 81.1200 ;
      RECT 60.2200 80.0400 103.0200 81.1200 ;
      RECT 15.2200 80.0400 58.0200 81.1200 ;
      RECT 4.8600 80.0400 13.0200 81.1200 ;
      RECT 0.0000 80.0400 1.2600 81.1200 ;
      RECT 0.0000 78.4000 210.2200 80.0400 ;
      RECT 204.9600 77.3200 210.2200 78.4000 ;
      RECT 192.0200 77.3200 201.3600 78.4000 ;
      RECT 147.0200 77.3200 189.8200 78.4000 ;
      RECT 102.0200 77.3200 144.8200 78.4000 ;
      RECT 57.0200 77.3200 99.8200 78.4000 ;
      RECT 8.8600 77.3200 54.8200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 210.2200 77.3200 ;
      RECT 208.9600 74.6000 210.2200 75.6800 ;
      RECT 195.2200 74.6000 205.3600 75.6800 ;
      RECT 150.2200 74.6000 193.0200 75.6800 ;
      RECT 105.2200 74.6000 148.0200 75.6800 ;
      RECT 60.2200 74.6000 103.0200 75.6800 ;
      RECT 15.2200 74.6000 58.0200 75.6800 ;
      RECT 4.8600 74.6000 13.0200 75.6800 ;
      RECT 0.0000 74.6000 1.2600 75.6800 ;
      RECT 0.0000 72.9600 210.2200 74.6000 ;
      RECT 204.9600 71.8800 210.2200 72.9600 ;
      RECT 192.0200 71.8800 201.3600 72.9600 ;
      RECT 147.0200 71.8800 189.8200 72.9600 ;
      RECT 102.0200 71.8800 144.8200 72.9600 ;
      RECT 57.0200 71.8800 99.8200 72.9600 ;
      RECT 8.8600 71.8800 54.8200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 210.2200 71.8800 ;
      RECT 208.9600 69.1600 210.2200 70.2400 ;
      RECT 195.2200 69.1600 205.3600 70.2400 ;
      RECT 150.2200 69.1600 193.0200 70.2400 ;
      RECT 105.2200 69.1600 148.0200 70.2400 ;
      RECT 60.2200 69.1600 103.0200 70.2400 ;
      RECT 15.2200 69.1600 58.0200 70.2400 ;
      RECT 4.8600 69.1600 13.0200 70.2400 ;
      RECT 0.0000 69.1600 1.2600 70.2400 ;
      RECT 0.0000 67.5200 210.2200 69.1600 ;
      RECT 204.9600 66.4400 210.2200 67.5200 ;
      RECT 192.0200 66.4400 201.3600 67.5200 ;
      RECT 147.0200 66.4400 189.8200 67.5200 ;
      RECT 102.0200 66.4400 144.8200 67.5200 ;
      RECT 57.0200 66.4400 99.8200 67.5200 ;
      RECT 8.8600 66.4400 54.8200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 210.2200 66.4400 ;
      RECT 208.9600 63.7200 210.2200 64.8000 ;
      RECT 195.2200 63.7200 205.3600 64.8000 ;
      RECT 150.2200 63.7200 193.0200 64.8000 ;
      RECT 105.2200 63.7200 148.0200 64.8000 ;
      RECT 60.2200 63.7200 103.0200 64.8000 ;
      RECT 15.2200 63.7200 58.0200 64.8000 ;
      RECT 4.8600 63.7200 13.0200 64.8000 ;
      RECT 0.0000 63.7200 1.2600 64.8000 ;
      RECT 0.0000 62.0800 210.2200 63.7200 ;
      RECT 204.9600 61.0000 210.2200 62.0800 ;
      RECT 192.0200 61.0000 201.3600 62.0800 ;
      RECT 147.0200 61.0000 189.8200 62.0800 ;
      RECT 102.0200 61.0000 144.8200 62.0800 ;
      RECT 57.0200 61.0000 99.8200 62.0800 ;
      RECT 8.8600 61.0000 54.8200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 210.2200 61.0000 ;
      RECT 208.9600 58.2800 210.2200 59.3600 ;
      RECT 195.2200 58.2800 205.3600 59.3600 ;
      RECT 150.2200 58.2800 193.0200 59.3600 ;
      RECT 105.2200 58.2800 148.0200 59.3600 ;
      RECT 60.2200 58.2800 103.0200 59.3600 ;
      RECT 15.2200 58.2800 58.0200 59.3600 ;
      RECT 4.8600 58.2800 13.0200 59.3600 ;
      RECT 0.0000 58.2800 1.2600 59.3600 ;
      RECT 0.0000 56.6400 210.2200 58.2800 ;
      RECT 204.9600 55.5600 210.2200 56.6400 ;
      RECT 192.0200 55.5600 201.3600 56.6400 ;
      RECT 147.0200 55.5600 189.8200 56.6400 ;
      RECT 102.0200 55.5600 144.8200 56.6400 ;
      RECT 57.0200 55.5600 99.8200 56.6400 ;
      RECT 8.8600 55.5600 54.8200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 210.2200 55.5600 ;
      RECT 208.9600 52.8400 210.2200 53.9200 ;
      RECT 195.2200 52.8400 205.3600 53.9200 ;
      RECT 150.2200 52.8400 193.0200 53.9200 ;
      RECT 105.2200 52.8400 148.0200 53.9200 ;
      RECT 60.2200 52.8400 103.0200 53.9200 ;
      RECT 15.2200 52.8400 58.0200 53.9200 ;
      RECT 4.8600 52.8400 13.0200 53.9200 ;
      RECT 0.0000 52.8400 1.2600 53.9200 ;
      RECT 0.0000 51.2000 210.2200 52.8400 ;
      RECT 204.9600 50.1200 210.2200 51.2000 ;
      RECT 192.0200 50.1200 201.3600 51.2000 ;
      RECT 147.0200 50.1200 189.8200 51.2000 ;
      RECT 102.0200 50.1200 144.8200 51.2000 ;
      RECT 57.0200 50.1200 99.8200 51.2000 ;
      RECT 8.8600 50.1200 54.8200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 210.2200 50.1200 ;
      RECT 208.9600 47.4000 210.2200 48.4800 ;
      RECT 195.2200 47.4000 205.3600 48.4800 ;
      RECT 150.2200 47.4000 193.0200 48.4800 ;
      RECT 105.2200 47.4000 148.0200 48.4800 ;
      RECT 60.2200 47.4000 103.0200 48.4800 ;
      RECT 15.2200 47.4000 58.0200 48.4800 ;
      RECT 4.8600 47.4000 13.0200 48.4800 ;
      RECT 0.0000 47.4000 1.2600 48.4800 ;
      RECT 0.0000 45.7600 210.2200 47.4000 ;
      RECT 204.9600 44.6800 210.2200 45.7600 ;
      RECT 192.0200 44.6800 201.3600 45.7600 ;
      RECT 147.0200 44.6800 189.8200 45.7600 ;
      RECT 102.0200 44.6800 144.8200 45.7600 ;
      RECT 57.0200 44.6800 99.8200 45.7600 ;
      RECT 8.8600 44.6800 54.8200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 210.2200 44.6800 ;
      RECT 208.9600 41.9600 210.2200 43.0400 ;
      RECT 195.2200 41.9600 205.3600 43.0400 ;
      RECT 150.2200 41.9600 193.0200 43.0400 ;
      RECT 105.2200 41.9600 148.0200 43.0400 ;
      RECT 60.2200 41.9600 103.0200 43.0400 ;
      RECT 15.2200 41.9600 58.0200 43.0400 ;
      RECT 4.8600 41.9600 13.0200 43.0400 ;
      RECT 0.0000 41.9600 1.2600 43.0400 ;
      RECT 0.0000 40.3200 210.2200 41.9600 ;
      RECT 204.9600 39.2400 210.2200 40.3200 ;
      RECT 192.0200 39.2400 201.3600 40.3200 ;
      RECT 147.0200 39.2400 189.8200 40.3200 ;
      RECT 102.0200 39.2400 144.8200 40.3200 ;
      RECT 57.0200 39.2400 99.8200 40.3200 ;
      RECT 8.8600 39.2400 54.8200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 210.2200 39.2400 ;
      RECT 208.9600 36.5200 210.2200 37.6000 ;
      RECT 195.2200 36.5200 205.3600 37.6000 ;
      RECT 150.2200 36.5200 193.0200 37.6000 ;
      RECT 105.2200 36.5200 148.0200 37.6000 ;
      RECT 60.2200 36.5200 103.0200 37.6000 ;
      RECT 15.2200 36.5200 58.0200 37.6000 ;
      RECT 4.8600 36.5200 13.0200 37.6000 ;
      RECT 0.0000 36.5200 1.2600 37.6000 ;
      RECT 0.0000 34.8800 210.2200 36.5200 ;
      RECT 204.9600 33.8000 210.2200 34.8800 ;
      RECT 192.0200 33.8000 201.3600 34.8800 ;
      RECT 147.0200 33.8000 189.8200 34.8800 ;
      RECT 102.0200 33.8000 144.8200 34.8800 ;
      RECT 57.0200 33.8000 99.8200 34.8800 ;
      RECT 8.8600 33.8000 54.8200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 210.2200 33.8000 ;
      RECT 208.9600 31.0800 210.2200 32.1600 ;
      RECT 195.2200 31.0800 205.3600 32.1600 ;
      RECT 150.2200 31.0800 193.0200 32.1600 ;
      RECT 105.2200 31.0800 148.0200 32.1600 ;
      RECT 60.2200 31.0800 103.0200 32.1600 ;
      RECT 15.2200 31.0800 58.0200 32.1600 ;
      RECT 4.8600 31.0800 13.0200 32.1600 ;
      RECT 0.0000 31.0800 1.2600 32.1600 ;
      RECT 0.0000 29.4400 210.2200 31.0800 ;
      RECT 204.9600 28.3600 210.2200 29.4400 ;
      RECT 192.0200 28.3600 201.3600 29.4400 ;
      RECT 147.0200 28.3600 189.8200 29.4400 ;
      RECT 102.0200 28.3600 144.8200 29.4400 ;
      RECT 57.0200 28.3600 99.8200 29.4400 ;
      RECT 8.8600 28.3600 54.8200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 210.2200 28.3600 ;
      RECT 208.9600 25.6400 210.2200 26.7200 ;
      RECT 195.2200 25.6400 205.3600 26.7200 ;
      RECT 150.2200 25.6400 193.0200 26.7200 ;
      RECT 105.2200 25.6400 148.0200 26.7200 ;
      RECT 60.2200 25.6400 103.0200 26.7200 ;
      RECT 15.2200 25.6400 58.0200 26.7200 ;
      RECT 4.8600 25.6400 13.0200 26.7200 ;
      RECT 0.0000 25.6400 1.2600 26.7200 ;
      RECT 0.0000 24.0000 210.2200 25.6400 ;
      RECT 204.9600 22.9200 210.2200 24.0000 ;
      RECT 192.0200 22.9200 201.3600 24.0000 ;
      RECT 147.0200 22.9200 189.8200 24.0000 ;
      RECT 102.0200 22.9200 144.8200 24.0000 ;
      RECT 57.0200 22.9200 99.8200 24.0000 ;
      RECT 8.8600 22.9200 54.8200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 210.2200 22.9200 ;
      RECT 208.9600 20.2000 210.2200 21.2800 ;
      RECT 195.2200 20.2000 205.3600 21.2800 ;
      RECT 150.2200 20.2000 193.0200 21.2800 ;
      RECT 105.2200 20.2000 148.0200 21.2800 ;
      RECT 60.2200 20.2000 103.0200 21.2800 ;
      RECT 15.2200 20.2000 58.0200 21.2800 ;
      RECT 4.8600 20.2000 13.0200 21.2800 ;
      RECT 0.0000 20.2000 1.2600 21.2800 ;
      RECT 0.0000 18.5600 210.2200 20.2000 ;
      RECT 204.9600 17.4800 210.2200 18.5600 ;
      RECT 192.0200 17.4800 201.3600 18.5600 ;
      RECT 147.0200 17.4800 189.8200 18.5600 ;
      RECT 102.0200 17.4800 144.8200 18.5600 ;
      RECT 57.0200 17.4800 99.8200 18.5600 ;
      RECT 8.8600 17.4800 54.8200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 210.2200 17.4800 ;
      RECT 208.9600 14.7600 210.2200 15.8400 ;
      RECT 195.2200 14.7600 205.3600 15.8400 ;
      RECT 150.2200 14.7600 193.0200 15.8400 ;
      RECT 105.2200 14.7600 148.0200 15.8400 ;
      RECT 60.2200 14.7600 103.0200 15.8400 ;
      RECT 15.2200 14.7600 58.0200 15.8400 ;
      RECT 4.8600 14.7600 13.0200 15.8400 ;
      RECT 0.0000 14.7600 1.2600 15.8400 ;
      RECT 0.0000 13.1200 210.2200 14.7600 ;
      RECT 204.9600 12.0400 210.2200 13.1200 ;
      RECT 192.0200 12.0400 201.3600 13.1200 ;
      RECT 147.0200 12.0400 189.8200 13.1200 ;
      RECT 102.0200 12.0400 144.8200 13.1200 ;
      RECT 57.0200 12.0400 99.8200 13.1200 ;
      RECT 8.8600 12.0400 54.8200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 210.2200 12.0400 ;
      RECT 208.9600 9.3200 210.2200 10.4000 ;
      RECT 195.2200 9.3200 205.3600 10.4000 ;
      RECT 150.2200 9.3200 193.0200 10.4000 ;
      RECT 105.2200 9.3200 148.0200 10.4000 ;
      RECT 60.2200 9.3200 103.0200 10.4000 ;
      RECT 15.2200 9.3200 58.0200 10.4000 ;
      RECT 4.8600 9.3200 13.0200 10.4000 ;
      RECT 0.0000 9.3200 1.2600 10.4000 ;
      RECT 0.0000 8.7300 210.2200 9.3200 ;
      RECT 204.9600 5.1300 210.2200 8.7300 ;
      RECT 0.0000 5.1300 5.2600 8.7300 ;
      RECT 0.0000 4.7300 210.2200 5.1300 ;
      RECT 208.9600 1.1300 210.2200 4.7300 ;
      RECT 0.0000 1.1300 1.2600 4.7300 ;
      RECT 0.0000 0.0000 210.2200 1.1300 ;
    LAYER met4 ;
      RECT 0.0000 217.8300 210.2200 219.6400 ;
      RECT 195.2200 213.8300 205.3600 217.8300 ;
      RECT 150.2200 213.8300 193.0200 217.8300 ;
      RECT 105.2200 213.8300 148.0200 217.8300 ;
      RECT 60.2200 213.8300 103.0200 217.8300 ;
      RECT 15.2200 213.8300 58.0200 217.8300 ;
      RECT 4.8600 213.8300 13.0200 217.8300 ;
      RECT 204.9600 5.1300 205.3600 213.8300 ;
      RECT 195.2200 5.1300 201.3600 213.8300 ;
      RECT 192.0200 5.1300 193.0200 213.8300 ;
      RECT 150.2200 5.1300 189.8200 213.8300 ;
      RECT 147.0200 5.1300 148.0200 213.8300 ;
      RECT 105.2200 5.1300 144.8200 213.8300 ;
      RECT 102.0200 5.1300 103.0200 213.8300 ;
      RECT 60.2200 5.1300 99.8200 213.8300 ;
      RECT 57.0200 5.1300 58.0200 213.8300 ;
      RECT 15.2200 5.1300 54.8200 213.8300 ;
      RECT 8.8600 5.1300 13.0200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 208.9600 1.1300 210.2200 217.8300 ;
      RECT 195.2200 1.1300 205.3600 5.1300 ;
      RECT 150.2200 1.1300 193.0200 5.1300 ;
      RECT 105.2200 1.1300 148.0200 5.1300 ;
      RECT 60.2200 1.1300 103.0200 5.1300 ;
      RECT 15.2200 1.1300 58.0200 5.1300 ;
      RECT 4.8600 1.1300 13.0200 5.1300 ;
      RECT 0.0000 1.1300 1.2600 217.8300 ;
      RECT 0.0000 1.1000 210.2200 1.1300 ;
      RECT 89.4600 0.0000 210.2200 1.1000 ;
      RECT 0.0000 0.0000 88.5600 1.1000 ;
  END
END LUT4AB

END LIBRARY
