magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 12748 3012 20068 4144
<< mvnsubdiff >>
rect 12814 4035 12852 4078
rect 12814 4001 12816 4035
rect 12850 4001 12852 4035
rect 13610 4035 13648 4078
rect 12814 3967 12852 4001
rect 12814 3933 12816 3967
rect 12850 3933 12852 3967
rect 12814 3899 12852 3933
rect 12814 3865 12816 3899
rect 12850 3865 12852 3899
rect 12814 3831 12852 3865
rect 12814 3797 12816 3831
rect 12850 3797 12852 3831
rect 12814 3763 12852 3797
rect 12814 3729 12816 3763
rect 12850 3729 12852 3763
rect 13610 4001 13612 4035
rect 13646 4001 13648 4035
rect 13610 3967 13648 4001
rect 13610 3933 13612 3967
rect 13646 3933 13648 3967
rect 13610 3899 13648 3933
rect 13610 3865 13612 3899
rect 13646 3865 13648 3899
rect 13610 3831 13648 3865
rect 13610 3797 13612 3831
rect 13646 3797 13648 3831
rect 13610 3763 13648 3797
rect 12814 3695 12852 3729
rect 13610 3729 13612 3763
rect 13646 3729 13648 3763
rect 12814 3661 12816 3695
rect 12850 3661 12852 3695
rect 12814 3627 12852 3661
rect 12814 3593 12816 3627
rect 12850 3593 12852 3627
rect 12814 3559 12852 3593
rect 12814 3525 12816 3559
rect 12850 3525 12852 3559
rect 12814 3491 12852 3525
rect 12814 3457 12816 3491
rect 12850 3457 12852 3491
rect 12814 3423 12852 3457
rect 12814 3389 12816 3423
rect 12850 3389 12852 3423
rect 12814 3355 12852 3389
rect 12814 3321 12816 3355
rect 12850 3321 12852 3355
rect 12814 3287 12852 3321
rect 12814 3253 12816 3287
rect 12850 3253 12852 3287
rect 12814 3219 12852 3253
rect 12814 3185 12816 3219
rect 12850 3185 12852 3219
rect 12814 3151 12852 3185
rect 12814 3117 12816 3151
rect 12850 3117 12852 3151
rect 12814 3078 12852 3117
rect 13610 3695 13648 3729
rect 13610 3661 13612 3695
rect 13646 3661 13648 3695
rect 13610 3627 13648 3661
rect 13610 3593 13612 3627
rect 13646 3593 13648 3627
rect 13610 3559 13648 3593
rect 13610 3525 13612 3559
rect 13646 3525 13648 3559
rect 13610 3491 13648 3525
rect 13610 3457 13612 3491
rect 13646 3457 13648 3491
rect 13610 3423 13648 3457
rect 13610 3389 13612 3423
rect 13646 3389 13648 3423
rect 13610 3355 13648 3389
rect 13610 3321 13612 3355
rect 13646 3321 13648 3355
rect 13610 3287 13648 3321
rect 13610 3253 13612 3287
rect 13646 3253 13648 3287
rect 13610 3219 13648 3253
rect 13610 3185 13612 3219
rect 13646 3185 13648 3219
rect 13610 3151 13648 3185
rect 13610 3117 13612 3151
rect 13646 3117 13648 3151
rect 13610 3078 13648 3117
rect 15210 4035 15248 4078
rect 15210 4001 15212 4035
rect 15246 4001 15248 4035
rect 15210 3967 15248 4001
rect 15210 3933 15212 3967
rect 15246 3933 15248 3967
rect 15210 3899 15248 3933
rect 15210 3865 15212 3899
rect 15246 3865 15248 3899
rect 15210 3831 15248 3865
rect 15210 3797 15212 3831
rect 15246 3797 15248 3831
rect 15210 3763 15248 3797
rect 15210 3729 15212 3763
rect 15246 3729 15248 3763
rect 15210 3695 15248 3729
rect 15210 3661 15212 3695
rect 15246 3661 15248 3695
rect 15210 3627 15248 3661
rect 15210 3593 15212 3627
rect 15246 3593 15248 3627
rect 15210 3559 15248 3593
rect 15210 3525 15212 3559
rect 15246 3525 15248 3559
rect 15210 3491 15248 3525
rect 15210 3457 15212 3491
rect 15246 3457 15248 3491
rect 15210 3423 15248 3457
rect 15210 3389 15212 3423
rect 15246 3389 15248 3423
rect 15210 3355 15248 3389
rect 15210 3321 15212 3355
rect 15246 3321 15248 3355
rect 15210 3287 15248 3321
rect 15210 3253 15212 3287
rect 15246 3253 15248 3287
rect 15210 3219 15248 3253
rect 15210 3185 15212 3219
rect 15246 3185 15248 3219
rect 15210 3151 15248 3185
rect 15210 3117 15212 3151
rect 15246 3117 15248 3151
rect 15210 3078 15248 3117
rect 16654 4035 16692 4078
rect 16654 4001 16656 4035
rect 16690 4001 16692 4035
rect 16654 3967 16692 4001
rect 16654 3933 16656 3967
rect 16690 3933 16692 3967
rect 16654 3899 16692 3933
rect 16654 3865 16656 3899
rect 16690 3865 16692 3899
rect 16654 3831 16692 3865
rect 16654 3797 16656 3831
rect 16690 3797 16692 3831
rect 16654 3763 16692 3797
rect 16654 3729 16656 3763
rect 16690 3729 16692 3763
rect 16654 3695 16692 3729
rect 16654 3661 16656 3695
rect 16690 3661 16692 3695
rect 16654 3627 16692 3661
rect 16654 3593 16656 3627
rect 16690 3593 16692 3627
rect 16654 3559 16692 3593
rect 16654 3525 16656 3559
rect 16690 3525 16692 3559
rect 16654 3491 16692 3525
rect 16654 3457 16656 3491
rect 16690 3457 16692 3491
rect 16654 3423 16692 3457
rect 16654 3389 16656 3423
rect 16690 3389 16692 3423
rect 16654 3355 16692 3389
rect 16654 3321 16656 3355
rect 16690 3321 16692 3355
rect 16654 3287 16692 3321
rect 16654 3253 16656 3287
rect 16690 3253 16692 3287
rect 16654 3219 16692 3253
rect 16654 3185 16656 3219
rect 16690 3185 16692 3219
rect 16654 3151 16692 3185
rect 16654 3117 16656 3151
rect 16690 3117 16692 3151
rect 16654 3078 16692 3117
rect 18098 4035 18136 4078
rect 18098 4001 18100 4035
rect 18134 4001 18136 4035
rect 18098 3967 18136 4001
rect 18098 3933 18100 3967
rect 18134 3933 18136 3967
rect 18098 3899 18136 3933
rect 18098 3865 18100 3899
rect 18134 3865 18136 3899
rect 18098 3831 18136 3865
rect 18098 3797 18100 3831
rect 18134 3797 18136 3831
rect 18098 3763 18136 3797
rect 18098 3729 18100 3763
rect 18134 3729 18136 3763
rect 18098 3695 18136 3729
rect 18098 3661 18100 3695
rect 18134 3661 18136 3695
rect 18098 3627 18136 3661
rect 18098 3593 18100 3627
rect 18134 3593 18136 3627
rect 18098 3559 18136 3593
rect 18098 3525 18100 3559
rect 18134 3525 18136 3559
rect 18098 3491 18136 3525
rect 18098 3457 18100 3491
rect 18134 3457 18136 3491
rect 18098 3423 18136 3457
rect 18098 3389 18100 3423
rect 18134 3389 18136 3423
rect 18098 3355 18136 3389
rect 18098 3321 18100 3355
rect 18134 3321 18136 3355
rect 18098 3287 18136 3321
rect 18098 3253 18100 3287
rect 18134 3253 18136 3287
rect 18098 3219 18136 3253
rect 18098 3185 18100 3219
rect 18134 3185 18136 3219
rect 18098 3151 18136 3185
rect 18098 3117 18100 3151
rect 18134 3117 18136 3151
rect 18098 3078 18136 3117
rect 19964 4035 20002 4078
rect 19964 4001 19966 4035
rect 20000 4001 20002 4035
rect 19964 3967 20002 4001
rect 19964 3933 19966 3967
rect 20000 3933 20002 3967
rect 19964 3899 20002 3933
rect 19964 3865 19966 3899
rect 20000 3865 20002 3899
rect 19964 3831 20002 3865
rect 19964 3797 19966 3831
rect 20000 3797 20002 3831
rect 19964 3763 20002 3797
rect 19964 3729 19966 3763
rect 20000 3729 20002 3763
rect 19964 3695 20002 3729
rect 19964 3661 19966 3695
rect 20000 3661 20002 3695
rect 19964 3627 20002 3661
rect 19964 3593 19966 3627
rect 20000 3593 20002 3627
rect 19964 3559 20002 3593
rect 19964 3525 19966 3559
rect 20000 3525 20002 3559
rect 19964 3491 20002 3525
rect 19964 3457 19966 3491
rect 20000 3457 20002 3491
rect 19964 3423 20002 3457
rect 19964 3389 19966 3423
rect 20000 3389 20002 3423
rect 19964 3355 20002 3389
rect 19964 3321 19966 3355
rect 20000 3321 20002 3355
rect 19964 3287 20002 3321
rect 19964 3253 19966 3287
rect 20000 3253 20002 3287
rect 19964 3219 20002 3253
rect 19964 3185 19966 3219
rect 20000 3185 20002 3219
rect 19964 3151 20002 3185
rect 19964 3117 19966 3151
rect 20000 3117 20002 3151
rect 19964 3078 20002 3117
<< mvnsubdiffcont >>
rect 12816 4001 12850 4035
rect 12816 3933 12850 3967
rect 12816 3865 12850 3899
rect 12816 3797 12850 3831
rect 12816 3729 12850 3763
rect 13612 4001 13646 4035
rect 13612 3933 13646 3967
rect 13612 3865 13646 3899
rect 13612 3797 13646 3831
rect 13612 3729 13646 3763
rect 12816 3661 12850 3695
rect 12816 3593 12850 3627
rect 12816 3525 12850 3559
rect 12816 3457 12850 3491
rect 12816 3389 12850 3423
rect 12816 3321 12850 3355
rect 12816 3253 12850 3287
rect 12816 3185 12850 3219
rect 12816 3117 12850 3151
rect 13612 3661 13646 3695
rect 13612 3593 13646 3627
rect 13612 3525 13646 3559
rect 13612 3457 13646 3491
rect 13612 3389 13646 3423
rect 13612 3321 13646 3355
rect 13612 3253 13646 3287
rect 13612 3185 13646 3219
rect 13612 3117 13646 3151
rect 15212 4001 15246 4035
rect 15212 3933 15246 3967
rect 15212 3865 15246 3899
rect 15212 3797 15246 3831
rect 15212 3729 15246 3763
rect 15212 3661 15246 3695
rect 15212 3593 15246 3627
rect 15212 3525 15246 3559
rect 15212 3457 15246 3491
rect 15212 3389 15246 3423
rect 15212 3321 15246 3355
rect 15212 3253 15246 3287
rect 15212 3185 15246 3219
rect 15212 3117 15246 3151
rect 16656 4001 16690 4035
rect 16656 3933 16690 3967
rect 16656 3865 16690 3899
rect 16656 3797 16690 3831
rect 16656 3729 16690 3763
rect 16656 3661 16690 3695
rect 16656 3593 16690 3627
rect 16656 3525 16690 3559
rect 16656 3457 16690 3491
rect 16656 3389 16690 3423
rect 16656 3321 16690 3355
rect 16656 3253 16690 3287
rect 16656 3185 16690 3219
rect 16656 3117 16690 3151
rect 18100 4001 18134 4035
rect 18100 3933 18134 3967
rect 18100 3865 18134 3899
rect 18100 3797 18134 3831
rect 18100 3729 18134 3763
rect 18100 3661 18134 3695
rect 18100 3593 18134 3627
rect 18100 3525 18134 3559
rect 18100 3457 18134 3491
rect 18100 3389 18134 3423
rect 18100 3321 18134 3355
rect 18100 3253 18134 3287
rect 18100 3185 18134 3219
rect 18100 3117 18134 3151
rect 19966 4001 20000 4035
rect 19966 3933 20000 3967
rect 19966 3865 20000 3899
rect 19966 3797 20000 3831
rect 19966 3729 20000 3763
rect 19966 3661 20000 3695
rect 19966 3593 20000 3627
rect 19966 3525 20000 3559
rect 19966 3457 20000 3491
rect 19966 3389 20000 3423
rect 19966 3321 20000 3355
rect 19966 3253 20000 3287
rect 19966 3185 20000 3219
rect 19966 3117 20000 3151
<< poly >>
rect 12159 5655 12293 5671
rect 12159 5621 12175 5655
rect 12209 5621 12243 5655
rect 12277 5621 12293 5655
rect 12159 5599 12293 5621
rect 13432 4788 13504 4804
rect 11368 4770 11434 4786
rect 11368 4736 11384 4770
rect 11418 4736 11434 4770
rect 11368 4702 11434 4736
rect 11368 4668 11384 4702
rect 11418 4668 11434 4702
rect 13432 4754 13454 4788
rect 13488 4754 13504 4788
rect 13432 4720 13504 4754
rect 13432 4686 13454 4720
rect 13488 4686 13504 4720
rect 13432 4670 13504 4686
rect 11368 4652 11434 4668
rect 12770 4593 12904 4609
rect 12770 4559 12786 4593
rect 12820 4559 12854 4593
rect 12888 4559 12904 4593
rect 12093 4537 12293 4547
rect 12770 4537 12904 4559
rect 13122 4593 13256 4609
rect 13122 4559 13138 4593
rect 13172 4559 13206 4593
rect 13240 4559 13256 4593
rect 13122 4537 13256 4559
rect 11581 4213 12549 4285
rect 12605 4263 12739 4285
rect 12605 4229 12621 4263
rect 12655 4229 12689 4263
rect 12723 4229 12739 4263
rect 12605 4213 12739 4229
rect 12957 4263 13091 4285
rect 12957 4229 12973 4263
rect 13007 4229 13041 4263
rect 13075 4229 13091 4263
rect 12957 4213 13091 4229
rect 13295 4263 13429 4285
rect 17679 4282 19279 4354
rect 13295 4229 13311 4263
rect 13345 4229 13379 4263
rect 13413 4229 13429 4263
rect 13295 4171 13429 4229
rect 13155 4155 13503 4171
rect 13155 4121 13171 4155
rect 13205 4121 13239 4155
rect 13273 4121 13307 4155
rect 13341 4121 13503 4155
rect 13155 4099 13503 4121
rect 19583 4160 19857 4176
rect 19583 4126 19599 4160
rect 19633 4126 19667 4160
rect 19701 4126 19735 4160
rect 19769 4126 19803 4160
rect 19837 4126 19857 4160
rect 19583 4104 19857 4126
rect 12336 3225 12408 4025
rect 12544 3225 12552 4025
rect 13016 4009 13088 4025
rect 13016 3975 13038 4009
rect 13072 3975 13088 4009
rect 13016 3941 13088 3975
rect 13016 3907 13038 3941
rect 13072 3907 13088 3941
rect 13016 3873 13088 3907
rect 13016 3839 13038 3873
rect 13072 3839 13088 3873
rect 13016 3805 13088 3839
rect 13016 3771 13038 3805
rect 13072 3771 13088 3805
rect 13016 3755 13088 3771
rect 13244 3789 13378 3805
rect 13244 3755 13260 3789
rect 13294 3755 13328 3789
rect 13362 3755 13378 3789
rect 13244 3739 13378 3755
rect 13261 3704 13361 3739
rect 13068 3030 13202 3052
rect 13068 2996 13084 3030
rect 13118 2996 13152 3030
rect 13186 2996 13202 3030
rect 13068 2980 13202 2996
rect 13420 3030 13554 3052
rect 13420 2996 13436 3030
rect 13470 2996 13504 3030
rect 13538 2996 13554 3030
rect 13420 2980 13554 2996
rect 13721 3030 13855 3052
rect 13721 2996 13737 3030
rect 13771 2996 13805 3030
rect 13839 2996 13855 3030
rect 13721 2980 13855 2996
rect 13911 2980 15103 3052
rect 15355 2980 16547 3052
rect 16799 2980 17991 3052
rect 18244 2980 18811 3052
rect 18868 2980 19435 3052
<< polycont >>
rect 12175 5621 12209 5655
rect 12243 5621 12277 5655
rect 11384 4736 11418 4770
rect 11384 4668 11418 4702
rect 13454 4754 13488 4788
rect 13454 4686 13488 4720
rect 12786 4559 12820 4593
rect 12854 4559 12888 4593
rect 13138 4559 13172 4593
rect 13206 4559 13240 4593
rect 12621 4229 12655 4263
rect 12689 4229 12723 4263
rect 12973 4229 13007 4263
rect 13041 4229 13075 4263
rect 13311 4229 13345 4263
rect 13379 4229 13413 4263
rect 13171 4121 13205 4155
rect 13239 4121 13273 4155
rect 13307 4121 13341 4155
rect 19599 4126 19633 4160
rect 19667 4126 19701 4160
rect 19735 4126 19769 4160
rect 19803 4126 19837 4160
rect 13038 3975 13072 4009
rect 13038 3907 13072 3941
rect 13038 3839 13072 3873
rect 13038 3771 13072 3805
rect 13260 3755 13294 3789
rect 13328 3755 13362 3789
rect 13084 2996 13118 3030
rect 13152 2996 13186 3030
rect 13436 2996 13470 3030
rect 13504 2996 13538 3030
rect 13737 2996 13771 3030
rect 13805 2996 13839 3030
<< locali >>
rect 12159 5621 12175 5655
rect 12209 5621 12243 5655
rect 12277 5621 12293 5655
rect 12304 5369 12338 5407
rect 12304 5297 12338 5335
rect 12296 4845 12841 4851
rect 12875 4845 12913 4879
rect 12947 4845 12985 4879
rect 13019 4845 13352 4851
rect 12296 4815 13352 4845
rect 11384 4770 11418 4786
rect 11572 4771 11610 4805
rect 11644 4771 11682 4805
rect 11716 4771 11754 4805
rect 11788 4771 11826 4805
rect 11860 4771 11898 4805
rect 11932 4771 11970 4805
rect 13420 4788 13458 4805
rect 13420 4771 13454 4788
rect 11384 4702 11418 4736
rect 13454 4720 13488 4754
rect 11418 4668 11522 4673
rect 11384 4639 11522 4668
rect 11572 4629 11610 4663
rect 11644 4629 11682 4663
rect 11716 4629 11754 4663
rect 11788 4629 11826 4663
rect 11860 4629 11898 4663
rect 11932 4629 11970 4663
rect 12090 4553 12128 4587
rect 11752 4391 11790 4425
rect 12266 4387 12304 4421
rect 11582 4313 11620 4347
rect 12048 4313 12086 4347
rect 12372 4229 12430 4673
rect 13454 4670 13488 4686
rect 12664 4571 12702 4605
rect 11590 4155 12430 4229
rect 12464 4307 12488 4341
rect 12522 4307 12560 4341
rect 12630 4307 12736 4571
rect 12770 4559 12786 4593
rect 12822 4559 12854 4593
rect 12894 4559 12904 4593
rect 12874 4313 12912 4347
rect 12980 4307 13088 4639
rect 13188 4593 13226 4602
rect 13122 4559 13138 4593
rect 13188 4568 13206 4593
rect 13260 4568 13298 4602
rect 13172 4559 13206 4568
rect 13240 4559 13256 4568
rect 13264 4313 13302 4347
rect 12464 4036 12530 4307
rect 12605 4229 12621 4263
rect 12655 4229 12689 4263
rect 12723 4229 12973 4263
rect 13007 4229 13041 4263
rect 13075 4229 13311 4263
rect 13345 4229 13379 4263
rect 13413 4229 13429 4263
rect 13148 4189 13412 4229
rect 13463 4195 13497 4509
rect 13024 4155 13062 4189
rect 13096 4155 13108 4189
rect 12602 4036 12640 4070
rect 12816 4035 12850 4070
rect 12816 3967 12850 4001
rect 12884 4013 12990 4070
rect 12918 3979 12956 4013
rect 13038 4009 13108 4155
rect 13182 4155 13220 4189
rect 13254 4155 13412 4189
rect 13148 4121 13171 4155
rect 13205 4121 13239 4155
rect 13273 4121 13307 4155
rect 13341 4121 13412 4155
rect 13446 4189 13497 4195
rect 13446 4155 13475 4189
rect 13509 4155 13547 4189
rect 13446 4141 13497 4155
rect 13446 4087 13480 4141
rect 12816 3899 12850 3933
rect 12816 3831 12850 3865
rect 13072 3975 13108 4009
rect 13038 3941 13108 3975
rect 13072 3907 13108 3941
rect 13038 3873 13108 3907
rect 13072 3839 13108 3873
rect 12816 3763 12850 3797
rect 12816 3695 12850 3729
rect 12816 3627 12850 3661
rect 12816 3559 12850 3593
rect 12816 3491 12850 3525
rect 12333 3395 12371 3429
rect 12816 3423 12850 3457
rect 12816 3355 12850 3389
rect 12816 3287 12850 3321
rect 12816 3219 12850 3253
rect 12522 3180 12600 3214
rect 12816 3151 12850 3185
rect 12888 3180 12994 3828
rect 13038 3805 13108 3839
rect 13072 3771 13108 3805
rect 13038 3140 13108 3771
rect 13192 3816 13226 4077
rect 13358 4053 13480 4087
rect 13358 4014 13392 4053
rect 13612 4035 13646 4051
rect 13320 3942 13358 3976
rect 13612 3967 13646 4001
rect 15212 4035 15246 4070
rect 16656 4035 16690 4070
rect 13612 3899 13646 3933
rect 13192 3744 13226 3782
rect 13192 3672 13226 3710
rect 13192 3631 13226 3638
rect 13260 3789 13362 3805
rect 13294 3755 13328 3789
rect 13260 3592 13362 3755
rect 13514 3669 13548 3875
rect 13710 3902 13744 3940
rect 15212 3967 15246 4001
rect 15212 3899 15246 3933
rect 13612 3831 13646 3865
rect 15212 3831 15246 3865
rect 13612 3763 13646 3797
rect 13612 3695 13646 3729
rect 13514 3616 13548 3638
rect 13612 3627 13646 3661
rect 13866 3744 13900 3782
rect 13866 3672 13900 3710
rect 14178 3744 14212 3782
rect 14178 3672 14212 3710
rect 14490 3744 14524 3782
rect 14490 3672 14524 3710
rect 14802 3744 14836 3782
rect 14802 3672 14836 3710
rect 15212 3763 15246 3797
rect 15212 3695 15246 3729
rect 13221 3558 13362 3592
rect 13187 3520 13362 3558
rect 13221 3486 13362 3520
rect 13612 3559 13646 3593
rect 13612 3491 13646 3525
rect 13612 3423 13646 3457
rect 13612 3355 13646 3389
rect 13612 3287 13646 3321
rect 13612 3219 13646 3253
rect 13612 3151 13646 3185
rect 12816 3082 12850 3117
rect 15212 3627 15246 3661
rect 15212 3559 15246 3593
rect 15212 3491 15246 3525
rect 15212 3423 15246 3457
rect 15212 3355 15246 3389
rect 15212 3287 15246 3321
rect 15212 3219 15246 3253
rect 15212 3151 15246 3185
rect 13612 3082 13646 3117
rect 14022 3066 14056 3132
rect 14334 3066 14368 3132
rect 14646 3066 14680 3132
rect 14958 3066 14992 3132
rect 15212 3082 15246 3117
rect 15305 3592 15339 4024
rect 16656 3967 16690 4001
rect 16656 3899 16690 3933
rect 15466 3862 15504 3896
rect 15778 3862 15816 3896
rect 16090 3862 16128 3896
rect 16402 3862 16440 3896
rect 16656 3831 16690 3865
rect 17634 3816 17724 4258
rect 18100 4035 18134 4070
rect 19290 4024 19324 4194
rect 19583 4155 19591 4189
rect 19625 4160 19663 4189
rect 19697 4160 19735 4189
rect 19769 4160 19807 4189
rect 19633 4155 19663 4160
rect 19583 4126 19599 4155
rect 19633 4126 19667 4155
rect 19701 4126 19735 4160
rect 19769 4126 19803 4160
rect 19841 4155 19853 4189
rect 19837 4126 19853 4155
rect 19966 4035 20000 4070
rect 18100 3967 18134 4001
rect 18100 3899 18134 3933
rect 18100 3831 18134 3865
rect 16656 3763 16690 3797
rect 16656 3695 16690 3729
rect 16656 3627 16690 3661
rect 17066 3744 17100 3782
rect 17066 3672 17100 3710
rect 17378 3744 17412 3782
rect 17378 3672 17412 3710
rect 17634 3638 17640 3816
rect 18100 3763 18134 3797
rect 18100 3695 18134 3729
rect 15305 3558 15311 3592
rect 15345 3558 15383 3592
rect 15623 3558 15661 3592
rect 15935 3558 15973 3592
rect 16247 3558 16285 3592
rect 16521 3558 16559 3592
rect 16656 3559 16690 3593
rect 13068 2996 13084 3064
rect 13118 3030 13156 3064
rect 13190 3030 13202 3064
rect 13438 3030 13476 3064
rect 13510 3030 13554 3064
rect 13118 2996 13152 3030
rect 13186 2996 13202 3030
rect 13420 2996 13436 3030
rect 13470 2996 13504 3030
rect 13538 2996 13554 3030
rect 13721 3030 13855 3066
rect 13721 2996 13737 3030
rect 13771 2996 13805 3030
rect 13839 2996 13855 3030
rect 13928 3032 15082 3066
rect 15305 3032 15339 3558
rect 16911 3558 16949 3592
rect 17222 3558 17260 3592
rect 17528 3558 17566 3592
rect 16656 3491 16690 3525
rect 16656 3423 16690 3457
rect 16656 3355 16690 3389
rect 16656 3287 16690 3321
rect 16656 3219 16690 3253
rect 16656 3151 16690 3185
rect 15466 3066 15500 3132
rect 15778 3066 15812 3132
rect 16090 3066 16124 3132
rect 16402 3066 16436 3132
rect 17634 3132 17724 3638
rect 18100 3627 18134 3661
rect 17846 3558 17884 3592
rect 18100 3559 18134 3593
rect 18833 3592 18867 4024
rect 19966 3967 20000 4001
rect 19966 3899 20000 3933
rect 19830 3862 19868 3896
rect 19966 3831 20000 3865
rect 19712 3744 19746 3782
rect 19712 3672 19746 3710
rect 19966 3763 20000 3782
rect 19966 3695 20000 3710
rect 19966 3627 20000 3638
rect 18232 3558 18270 3592
rect 18510 3558 18548 3592
rect 18822 3558 18860 3592
rect 19134 3558 19172 3592
rect 19408 3558 19446 3592
rect 19966 3559 20000 3593
rect 18100 3491 18134 3525
rect 18100 3423 18134 3457
rect 18354 3422 18392 3456
rect 18665 3422 18703 3456
rect 18100 3355 18134 3389
rect 18100 3287 18134 3321
rect 18100 3219 18134 3253
rect 18100 3151 18134 3185
rect 16656 3082 16690 3117
rect 18100 3082 18134 3117
rect 13928 2996 15339 3032
rect 15373 3030 16527 3066
rect 16817 2996 17971 3060
rect 18354 3030 18388 3132
rect 18666 3030 18700 3132
rect 18833 3030 18867 3558
rect 19966 3491 20000 3525
rect 19966 3423 20000 3457
rect 18978 3336 19016 3370
rect 19289 3336 19327 3370
rect 19590 3336 19628 3370
rect 19966 3355 20000 3389
rect 19966 3287 20000 3321
rect 19966 3219 20000 3253
rect 19966 3151 20000 3185
rect 19134 3030 19168 3132
rect 19446 3030 19480 3132
rect 19966 3082 20000 3117
rect 18833 2996 18890 3030
rect 19423 2996 19480 3030
<< viali >>
rect 12304 5407 12338 5441
rect 12304 5335 12338 5369
rect 12304 5263 12338 5297
rect 12296 4851 12402 4957
rect 12841 4845 12875 4879
rect 12913 4845 12947 4879
rect 12985 4845 13019 4879
rect 11538 4771 11572 4805
rect 11610 4771 11644 4805
rect 11682 4771 11716 4805
rect 11754 4771 11788 4805
rect 11826 4771 11860 4805
rect 11898 4771 11932 4805
rect 11970 4771 12004 4805
rect 13386 4771 13420 4805
rect 13458 4788 13492 4805
rect 13458 4771 13488 4788
rect 13488 4771 13492 4788
rect 11538 4629 11572 4663
rect 11610 4629 11644 4663
rect 11682 4629 11716 4663
rect 11754 4629 11788 4663
rect 11826 4629 11860 4663
rect 11898 4629 11932 4663
rect 11970 4629 12004 4663
rect 12056 4553 12090 4587
rect 12128 4553 12162 4587
rect 11718 4391 11752 4425
rect 11790 4391 11824 4425
rect 12232 4387 12266 4421
rect 12304 4387 12338 4421
rect 11548 4313 11582 4347
rect 11620 4313 11654 4347
rect 12014 4313 12048 4347
rect 12086 4313 12120 4347
rect 12630 4571 12664 4605
rect 12702 4571 12736 4605
rect 12488 4307 12522 4341
rect 12560 4307 12594 4341
rect 12788 4559 12820 4593
rect 12820 4559 12822 4593
rect 12860 4559 12888 4593
rect 12888 4559 12894 4593
rect 12840 4313 12874 4347
rect 12912 4313 12946 4347
rect 13154 4593 13188 4602
rect 13226 4593 13260 4602
rect 13154 4568 13172 4593
rect 13172 4568 13188 4593
rect 13226 4568 13240 4593
rect 13240 4568 13260 4593
rect 13298 4568 13332 4602
rect 13230 4313 13264 4347
rect 13302 4313 13336 4347
rect 12990 4155 13024 4189
rect 13062 4155 13096 4189
rect 12568 4036 12602 4070
rect 12640 4036 12674 4070
rect 12884 3979 12918 4013
rect 12956 3979 12990 4013
rect 13148 4155 13182 4189
rect 13220 4155 13254 4189
rect 13475 4155 13509 4189
rect 13547 4155 13581 4189
rect 12299 3395 12333 3429
rect 12371 3395 12405 3429
rect 13286 3942 13320 3976
rect 13358 3942 13392 3976
rect 13192 3782 13226 3816
rect 13192 3710 13226 3744
rect 13192 3638 13226 3672
rect 13710 3940 13744 3974
rect 13710 3868 13744 3902
rect 13866 3782 13900 3816
rect 13866 3710 13900 3744
rect 13866 3638 13900 3672
rect 14178 3782 14212 3816
rect 14178 3710 14212 3744
rect 14178 3638 14212 3672
rect 14490 3782 14524 3816
rect 14490 3710 14524 3744
rect 14490 3638 14524 3672
rect 14802 3782 14836 3816
rect 14802 3710 14836 3744
rect 14802 3638 14836 3672
rect 13187 3558 13221 3592
rect 13187 3486 13221 3520
rect 15432 3862 15466 3896
rect 15504 3862 15538 3896
rect 15744 3862 15778 3896
rect 15816 3862 15850 3896
rect 16056 3862 16090 3896
rect 16128 3862 16162 3896
rect 16368 3862 16402 3896
rect 16440 3862 16474 3896
rect 19591 4160 19625 4189
rect 19663 4160 19697 4189
rect 19735 4160 19769 4189
rect 19807 4160 19841 4189
rect 19591 4155 19599 4160
rect 19599 4155 19625 4160
rect 19663 4155 19667 4160
rect 19667 4155 19697 4160
rect 19735 4155 19769 4160
rect 19807 4155 19837 4160
rect 19837 4155 19841 4160
rect 17066 3782 17100 3816
rect 17066 3710 17100 3744
rect 17066 3638 17100 3672
rect 17378 3782 17412 3816
rect 17378 3710 17412 3744
rect 17378 3638 17412 3672
rect 17640 3638 17746 3816
rect 15311 3558 15345 3592
rect 15383 3558 15417 3592
rect 15589 3558 15623 3592
rect 15661 3558 15695 3592
rect 15901 3558 15935 3592
rect 15973 3558 16007 3592
rect 16213 3558 16247 3592
rect 16285 3558 16319 3592
rect 16487 3558 16521 3592
rect 16559 3558 16593 3592
rect 13084 3030 13118 3064
rect 13156 3030 13190 3064
rect 13404 3030 13438 3064
rect 13476 3030 13510 3064
rect 16877 3558 16911 3592
rect 16949 3558 16983 3592
rect 17188 3558 17222 3592
rect 17260 3558 17294 3592
rect 17494 3558 17528 3592
rect 17566 3558 17600 3592
rect 17812 3558 17846 3592
rect 17884 3558 17918 3592
rect 19796 3862 19830 3896
rect 19868 3862 19902 3896
rect 19712 3782 19746 3816
rect 19712 3710 19746 3744
rect 19712 3638 19746 3672
rect 19966 3797 20000 3816
rect 19966 3782 20000 3797
rect 19966 3729 20000 3744
rect 19966 3710 20000 3729
rect 19966 3661 20000 3672
rect 19966 3638 20000 3661
rect 18198 3558 18232 3592
rect 18270 3558 18304 3592
rect 18476 3558 18510 3592
rect 18548 3558 18582 3592
rect 18788 3558 18822 3592
rect 18860 3558 18894 3592
rect 19100 3558 19134 3592
rect 19172 3558 19206 3592
rect 19374 3558 19408 3592
rect 19446 3558 19480 3592
rect 18320 3422 18354 3456
rect 18392 3422 18426 3456
rect 18631 3422 18665 3456
rect 18703 3422 18737 3456
rect 18944 3336 18978 3370
rect 19016 3336 19050 3370
rect 19255 3336 19289 3370
rect 19327 3336 19361 3370
rect 19556 3336 19590 3370
rect 19628 3336 19662 3370
<< metal1 >>
rect 11364 5441 13508 5453
rect 11364 5407 12304 5441
rect 12338 5407 13508 5441
rect 11364 5369 13508 5407
rect 11364 5335 12304 5369
rect 12338 5335 13508 5369
rect 11364 5297 13508 5335
rect 11364 5263 12304 5297
rect 12338 5263 13508 5297
rect 11364 5251 13508 5263
rect 11364 4957 13508 4969
rect 11364 4851 12296 4957
rect 12402 4879 13508 4957
rect 12402 4851 12841 4879
rect 11364 4845 12841 4851
rect 12875 4845 12913 4879
rect 12947 4845 12985 4879
rect 13019 4845 13508 4879
rect 11364 4839 13508 4845
rect 11523 4805 13504 4811
rect 11523 4771 11538 4805
rect 11572 4771 11610 4805
rect 11644 4771 11682 4805
rect 11716 4771 11754 4805
rect 11788 4771 11826 4805
rect 11860 4771 11898 4805
rect 11932 4771 11970 4805
rect 12004 4771 13386 4805
rect 13420 4771 13458 4805
rect 13492 4771 13504 4805
rect 11523 4765 13504 4771
rect 11523 4740 12023 4765
tri 12023 4740 12048 4765 nw
tri 12593 4740 12618 4765 ne
rect 11524 4738 12022 4739
rect 11524 4701 12022 4702
rect 11523 4675 12023 4700
tri 12023 4675 12048 4700 sw
rect 11523 4623 11529 4675
rect 11581 4623 11593 4675
rect 11645 4663 12258 4675
rect 11645 4629 11682 4663
rect 11716 4629 11754 4663
rect 11788 4629 11826 4663
rect 11860 4629 11898 4663
rect 11932 4629 11970 4663
rect 12004 4629 12258 4663
rect 11645 4623 12258 4629
rect 12618 4605 12748 4765
tri 12748 4740 12773 4765 nw
rect 11612 4543 11618 4595
rect 11670 4543 11682 4595
rect 11734 4587 12174 4595
rect 11734 4553 12056 4587
rect 12090 4553 12128 4587
rect 12162 4553 12174 4587
rect 12618 4571 12630 4605
rect 12664 4571 12702 4605
rect 12736 4571 12748 4605
rect 12618 4565 12748 4571
rect 12776 4636 13508 4682
rect 12776 4623 12918 4636
tri 12918 4623 12931 4636 nw
rect 12776 4593 12906 4623
tri 12906 4611 12918 4623 nw
rect 12776 4559 12788 4593
rect 12822 4559 12860 4593
rect 12894 4559 12906 4593
rect 12776 4553 12906 4559
rect 13142 4602 13222 4608
rect 13142 4568 13154 4602
rect 13188 4568 13222 4602
rect 13142 4556 13222 4568
rect 13274 4556 13286 4608
rect 13338 4556 13344 4608
rect 11734 4543 12174 4553
rect 11706 4425 11839 4433
rect 11841 4432 11877 4433
rect 11706 4391 11718 4425
rect 11752 4391 11790 4425
rect 11824 4391 11839 4425
rect 11706 4381 11839 4391
rect 11840 4382 11878 4432
rect 11879 4421 12478 4433
rect 11879 4387 12232 4421
rect 12266 4387 12304 4421
rect 12338 4387 12478 4421
rect 11841 4381 11877 4382
rect 11879 4381 12478 4387
rect 12530 4381 12542 4433
rect 12594 4381 12600 4433
rect 11364 4347 20068 4353
rect 11364 4313 11548 4347
rect 11582 4313 11620 4347
rect 11654 4313 12014 4347
rect 12048 4313 12086 4347
rect 12120 4341 12840 4347
rect 12120 4313 12488 4341
rect 11364 4307 12488 4313
rect 12522 4307 12560 4341
rect 12594 4313 12840 4341
rect 12874 4313 12912 4347
rect 12946 4313 13230 4347
rect 13264 4313 13302 4347
rect 13336 4313 20068 4347
rect 12594 4307 20068 4313
rect 11364 4223 20068 4307
rect 11589 4189 13108 4195
rect 11589 4155 12990 4189
rect 13024 4155 13062 4189
rect 13096 4155 13108 4189
rect 11589 4149 13108 4155
tri 12531 4124 12556 4149 ne
rect 12556 4143 12705 4149
tri 12705 4143 12711 4149 nw
rect 13136 4143 13142 4195
rect 13194 4143 13206 4195
rect 13258 4143 13266 4195
rect 13463 4189 19854 4195
rect 13463 4155 13475 4189
rect 13509 4155 13547 4189
rect 13581 4155 19591 4189
rect 19625 4155 19663 4189
rect 19697 4155 19735 4189
rect 19769 4155 19807 4189
rect 19841 4155 19854 4189
rect 13463 4149 19854 4155
rect 12556 4124 12686 4143
tri 12686 4124 12705 4143 nw
rect 12557 4122 12685 4123
rect 12556 4086 12686 4122
rect 12557 4085 12685 4086
rect 12556 4070 12686 4084
rect 12556 4036 12568 4070
rect 12602 4036 12640 4070
rect 12674 4036 12686 4070
rect 12556 4030 12686 4036
rect 12872 4013 13002 4025
rect 12872 3979 12884 4013
rect 12918 3979 12956 4013
rect 12990 3979 13002 4013
rect 12872 3973 13002 3979
rect 12873 3971 13001 3972
rect 12872 3935 13002 3971
rect 13274 3976 13404 3982
rect 13274 3942 13286 3976
rect 13320 3942 13358 3976
rect 13392 3942 13404 3976
rect 13274 3936 13404 3942
rect 13704 3974 13750 3986
rect 13704 3940 13710 3974
rect 13744 3940 13750 3974
rect 12873 3934 13001 3935
tri 12847 3908 12872 3933 se
rect 12872 3908 13002 3933
tri 13002 3908 13027 3933 sw
tri 13679 3908 13704 3933 se
rect 13704 3908 13750 3940
tri 13750 3908 13775 3933 sw
rect 11428 3856 12478 3908
rect 12530 3856 12542 3908
rect 12594 3902 19963 3908
rect 12594 3868 13710 3902
rect 13744 3896 19963 3902
rect 13744 3868 15432 3896
rect 12594 3862 15432 3868
rect 15466 3862 15504 3896
rect 15538 3862 15744 3896
rect 15778 3862 15816 3896
rect 15850 3862 16056 3896
rect 16090 3862 16128 3896
rect 16162 3862 16368 3896
rect 16402 3862 16440 3896
rect 16474 3862 19796 3896
rect 19830 3862 19868 3896
rect 19902 3862 19963 3896
rect 12594 3856 19963 3862
rect 11364 3816 20068 3828
rect 11364 3782 13192 3816
rect 13226 3782 13866 3816
rect 13900 3782 14178 3816
rect 14212 3782 14490 3816
rect 14524 3782 14802 3816
rect 14836 3782 17066 3816
rect 17100 3782 17378 3816
rect 17412 3782 17640 3816
rect 11364 3744 17640 3782
rect 11364 3710 13192 3744
rect 13226 3710 13866 3744
rect 13900 3710 14178 3744
rect 14212 3710 14490 3744
rect 14524 3710 14802 3744
rect 14836 3710 17066 3744
rect 17100 3710 17378 3744
rect 17412 3710 17640 3744
rect 11364 3672 17640 3710
rect 11364 3638 13192 3672
rect 13226 3638 13866 3672
rect 13900 3638 14178 3672
rect 14212 3638 14490 3672
rect 14524 3638 14802 3672
rect 14836 3638 17066 3672
rect 17100 3638 17378 3672
rect 17412 3638 17640 3672
rect 17746 3782 19712 3816
rect 19746 3782 19966 3816
rect 20000 3782 20068 3816
rect 17746 3744 20068 3782
rect 17746 3710 19712 3744
rect 19746 3710 19966 3744
rect 20000 3710 20068 3744
rect 17746 3672 20068 3710
rect 17746 3638 19712 3672
rect 19746 3638 19966 3672
rect 20000 3638 20068 3672
rect 11364 3626 20068 3638
rect 11523 3546 11529 3598
rect 11581 3546 11593 3598
rect 11645 3592 13250 3598
rect 11645 3558 13187 3592
rect 13221 3558 13250 3592
rect 11645 3546 13250 3558
tri 13104 3520 13130 3546 ne
rect 13130 3520 13250 3546
tri 13130 3518 13132 3520 ne
rect 13132 3518 13187 3520
rect 11612 3466 11618 3518
rect 11670 3466 11682 3518
rect 11734 3516 13092 3518
tri 13092 3516 13094 3518 sw
tri 13132 3516 13134 3518 ne
rect 13134 3516 13187 3518
rect 11734 3486 13094 3516
tri 13094 3486 13124 3516 sw
tri 13134 3486 13164 3516 ne
rect 13164 3486 13187 3516
rect 13221 3486 13250 3520
rect 11734 3482 13124 3486
tri 13124 3482 13128 3486 sw
tri 13164 3482 13168 3486 ne
rect 13168 3482 13250 3486
rect 11734 3480 13128 3482
tri 13128 3480 13130 3482 sw
tri 13168 3480 13170 3482 ne
rect 13170 3480 13250 3482
rect 11734 3470 13130 3480
tri 13130 3470 13140 3480 sw
tri 13170 3470 13180 3480 ne
rect 13180 3470 13250 3480
rect 13251 3471 13252 3597
rect 13288 3471 13289 3597
rect 13290 3592 13344 3598
rect 13290 3540 13292 3592
rect 15299 3592 16796 3598
rect 16798 3597 16834 3598
rect 15299 3558 15311 3592
rect 15345 3558 15383 3592
rect 15417 3558 15589 3592
rect 15623 3558 15661 3592
rect 15695 3558 15901 3592
rect 15935 3558 15973 3592
rect 16007 3558 16213 3592
rect 16247 3558 16285 3592
rect 16319 3558 16487 3592
rect 16521 3558 16559 3592
rect 16593 3558 16796 3592
rect 15299 3552 16796 3558
rect 16797 3553 16835 3597
rect 16836 3592 17930 3598
rect 16836 3558 16877 3592
rect 16911 3558 16949 3592
rect 16983 3558 17188 3592
rect 17222 3558 17260 3592
rect 17294 3558 17494 3592
rect 17528 3558 17566 3592
rect 17600 3558 17812 3592
rect 17846 3558 17884 3592
rect 17918 3558 17930 3592
rect 16798 3552 16834 3553
rect 16836 3552 17930 3558
rect 18186 3592 19492 3598
rect 18186 3558 18198 3592
rect 18232 3558 18270 3592
rect 18304 3558 18476 3592
rect 18510 3558 18548 3592
rect 18582 3558 18788 3592
rect 18822 3558 18860 3592
rect 18894 3558 19100 3592
rect 19134 3558 19172 3592
rect 19206 3558 19374 3592
rect 19408 3558 19446 3592
rect 19480 3558 19492 3592
rect 18186 3552 19492 3558
rect 13290 3528 13344 3540
rect 13290 3476 13292 3528
rect 13290 3470 13344 3476
rect 11734 3466 13140 3470
tri 13140 3466 13144 3470 sw
tri 13070 3456 13080 3466 ne
rect 13080 3462 13144 3466
tri 13144 3462 13148 3466 sw
rect 13080 3456 13148 3462
tri 13148 3456 13154 3462 sw
tri 13474 3456 13480 3462 se
rect 13480 3456 18749 3462
tri 13080 3442 13094 3456 ne
rect 13094 3442 13154 3456
tri 13154 3442 13168 3456 sw
tri 13460 3442 13474 3456 se
rect 13474 3442 18320 3456
tri 13094 3438 13098 3442 ne
rect 13098 3438 18320 3442
rect 11523 3386 11529 3438
rect 11581 3386 11593 3438
rect 11645 3386 11680 3438
rect 11682 3437 11718 3438
rect 11681 3387 11719 3437
rect 11720 3429 12417 3438
tri 13098 3435 13101 3438 ne
rect 13101 3435 18320 3438
rect 11720 3395 12299 3429
rect 12333 3395 12371 3429
rect 12405 3395 12417 3429
tri 13101 3422 13114 3435 ne
rect 13114 3422 18320 3435
rect 18354 3422 18392 3456
rect 18426 3422 18631 3456
rect 18665 3422 18703 3456
rect 18737 3422 18749 3456
tri 13114 3416 13120 3422 ne
rect 13120 3416 18749 3422
rect 11682 3386 11718 3387
rect 11720 3386 12417 3395
tri 13120 3390 13146 3416 ne
rect 13146 3410 18749 3416
rect 13146 3390 13482 3410
tri 13482 3390 13502 3410 nw
rect 17238 3330 17736 3382
rect 17788 3330 17800 3382
rect 17852 3370 19674 3382
rect 17852 3336 18944 3370
rect 18978 3336 19016 3370
rect 19050 3336 19255 3370
rect 19289 3336 19327 3370
rect 19361 3336 19556 3370
rect 19590 3336 19628 3370
rect 19662 3336 19674 3370
rect 17852 3330 19674 3336
rect 11364 3100 20068 3302
rect 13068 3064 13142 3072
rect 13068 3030 13084 3064
rect 13118 3030 13142 3064
rect 13068 3020 13142 3030
rect 13194 3020 13206 3072
rect 13258 3020 13264 3072
rect 13292 3020 13298 3072
rect 13350 3020 13362 3072
rect 13414 3064 13554 3072
rect 13438 3030 13476 3064
rect 13510 3030 13554 3064
rect 13414 3020 13554 3030
rect 15077 3026 15352 3072
rect 15353 3027 15354 3071
rect 15390 3027 15391 3071
rect 15392 3026 15444 3072
rect 16818 3020 17736 3072
rect 17788 3020 17800 3072
rect 17852 3020 17956 3072
<< rmetal1 >>
rect 11523 4739 12023 4740
rect 11523 4738 11524 4739
rect 12022 4738 12023 4739
rect 11523 4701 11524 4702
rect 12022 4701 12023 4702
rect 11523 4700 12023 4701
rect 11839 4432 11841 4433
rect 11877 4432 11879 4433
rect 11839 4382 11840 4432
rect 11878 4382 11879 4432
rect 11839 4381 11841 4382
rect 11877 4381 11879 4382
rect 12556 4123 12686 4124
rect 12556 4122 12557 4123
rect 12685 4122 12686 4123
rect 12556 4085 12557 4086
rect 12685 4085 12686 4086
rect 12556 4084 12686 4085
rect 12872 3972 13002 3973
rect 12872 3971 12873 3972
rect 13001 3971 13002 3972
rect 12872 3934 12873 3935
rect 13001 3934 13002 3935
rect 12872 3933 13002 3934
rect 13250 3597 13252 3598
rect 13250 3471 13251 3597
rect 13250 3470 13252 3471
rect 13288 3597 13290 3598
rect 13289 3471 13290 3597
rect 16796 3597 16798 3598
rect 16834 3597 16836 3598
rect 16796 3553 16797 3597
rect 16835 3553 16836 3597
rect 16796 3552 16798 3553
rect 16834 3552 16836 3553
rect 13288 3470 13290 3471
rect 11680 3437 11682 3438
rect 11718 3437 11720 3438
rect 11680 3387 11681 3437
rect 11719 3387 11720 3437
rect 11680 3386 11682 3387
rect 11718 3386 11720 3387
rect 15352 3071 15354 3072
rect 15352 3027 15353 3071
rect 15352 3026 15354 3027
rect 15390 3071 15392 3072
rect 15391 3027 15392 3071
rect 15390 3026 15392 3027
<< via1 >>
rect 11529 4663 11581 4675
rect 11529 4629 11538 4663
rect 11538 4629 11572 4663
rect 11572 4629 11581 4663
rect 11529 4623 11581 4629
rect 11593 4663 11645 4675
rect 11593 4629 11610 4663
rect 11610 4629 11644 4663
rect 11644 4629 11645 4663
rect 11593 4623 11645 4629
rect 11618 4543 11670 4595
rect 11682 4543 11734 4595
rect 13222 4602 13274 4608
rect 13222 4568 13226 4602
rect 13226 4568 13260 4602
rect 13260 4568 13274 4602
rect 13222 4556 13274 4568
rect 13286 4602 13338 4608
rect 13286 4568 13298 4602
rect 13298 4568 13332 4602
rect 13332 4568 13338 4602
rect 13286 4556 13338 4568
rect 12478 4381 12530 4433
rect 12542 4381 12594 4433
rect 13142 4189 13194 4195
rect 13142 4155 13148 4189
rect 13148 4155 13182 4189
rect 13182 4155 13194 4189
rect 13142 4143 13194 4155
rect 13206 4189 13258 4195
rect 13206 4155 13220 4189
rect 13220 4155 13254 4189
rect 13254 4155 13258 4189
rect 13206 4143 13258 4155
rect 12478 3856 12530 3908
rect 12542 3856 12594 3908
rect 11529 3546 11581 3598
rect 11593 3546 11645 3598
rect 11618 3466 11670 3518
rect 11682 3466 11734 3518
rect 13292 3540 13344 3592
rect 13292 3476 13344 3528
rect 11529 3386 11581 3438
rect 11593 3386 11645 3438
rect 17736 3330 17788 3382
rect 17800 3330 17852 3382
rect 13142 3064 13194 3072
rect 13142 3030 13156 3064
rect 13156 3030 13190 3064
rect 13190 3030 13194 3064
rect 13142 3020 13194 3030
rect 13206 3020 13258 3072
rect 13298 3020 13350 3072
rect 13362 3064 13414 3072
rect 13362 3030 13404 3064
rect 13404 3030 13414 3064
rect 13362 3020 13414 3030
rect 17736 3020 17788 3072
rect 17800 3020 17852 3072
<< metal2 >>
rect 11523 4623 11529 4675
rect 11581 4623 11593 4675
rect 11645 4623 11651 4675
rect 11523 4608 11585 4623
tri 11585 4608 11600 4623 nw
rect 11523 3598 11575 4608
tri 11575 4598 11585 4608 nw
rect 11612 4543 11618 4595
rect 11670 4543 11682 4595
rect 11734 4543 11740 4595
rect 13216 4556 13222 4608
rect 13274 4556 13286 4608
rect 13338 4556 13344 4608
tri 13267 4543 13280 4556 ne
rect 13280 4543 13344 4556
tri 11663 4531 11675 4543 ne
rect 11675 4531 11740 4543
tri 13280 4531 13292 4543 ne
tri 11675 4518 11688 4531 ne
tri 11575 3598 11600 3623 sw
rect 11523 3546 11529 3598
rect 11581 3546 11593 3598
rect 11645 3546 11651 3598
rect 11523 3540 11594 3546
tri 11594 3540 11600 3546 nw
tri 11685 3540 11688 3543 se
rect 11688 3540 11740 4531
rect 12472 4381 12478 4433
rect 12530 4381 12542 4433
rect 12594 4381 12600 4433
rect 12472 3908 12524 4381
tri 12524 4356 12549 4381 nw
rect 13136 4143 13142 4195
rect 13194 4143 13206 4195
rect 13258 4143 13264 4195
tri 12524 3908 12549 3933 sw
rect 12472 3856 12478 3908
rect 12530 3856 12542 3908
rect 12594 3856 12600 3908
rect 11523 3528 11582 3540
tri 11582 3528 11594 3540 nw
tri 11673 3528 11685 3540 se
rect 11685 3528 11740 3540
rect 11523 3438 11575 3528
tri 11575 3521 11582 3528 nw
tri 11666 3521 11673 3528 se
rect 11673 3521 11740 3528
tri 11663 3518 11666 3521 se
rect 11666 3518 11740 3521
rect 11612 3466 11618 3518
rect 11670 3466 11682 3518
rect 11734 3466 11740 3518
tri 11575 3438 11600 3463 sw
rect 11523 3386 11529 3438
rect 11581 3386 11593 3438
rect 11645 3386 11651 3438
rect 13136 3072 13188 4143
tri 13188 4118 13213 4143 nw
rect 13292 3592 13344 4543
rect 13292 3528 13344 3540
tri 13188 3072 13213 3097 sw
rect 13292 3072 13344 3476
rect 17730 3330 17736 3382
rect 17788 3330 17800 3382
rect 17852 3330 17858 3382
tri 13344 3072 13369 3097 sw
rect 17730 3072 17858 3330
rect 13136 3020 13142 3072
rect 13194 3020 13206 3072
rect 13258 3020 13264 3072
rect 13292 3020 13298 3072
rect 13350 3020 13362 3072
rect 13414 3020 13420 3072
rect 17730 3020 17736 3072
rect 17788 3020 17800 3072
rect 17852 3020 17858 3072
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 13221 0 -1 3592
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 12894 0 1 4559
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 13510 0 1 3030
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 12736 0 1 4571
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 12674 0 1 4036
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 12990 0 -1 4013
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 13392 0 -1 3976
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 1 13710 1 0 3868
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 1 0 13386 0 -1 4805
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 1 0 13084 0 -1 3064
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 12299 0 -1 3429
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 12840 0 1 4313
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 13230 0 1 4313
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 12488 0 1 4307
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 11548 0 1 4313
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 12014 0 1 4313
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 18788 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 19100 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 19374 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 18476 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 18198 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 18944 0 1 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 19255 0 1 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 18320 0 1 3422
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 18631 0 1 3422
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 19556 0 1 3336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 15311 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 15589 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 1 0 16487 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 1 0 16213 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1707688321
transform 1 0 15901 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1707688321
transform 1 0 17188 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1707688321
transform 1 0 16877 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1707688321
transform 1 0 17812 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1707688321
transform 1 0 17494 0 1 3558
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1707688321
transform 1 0 13148 0 1 4155
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1707688321
transform 1 0 13475 0 1 4155
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1707688321
transform 1 0 12056 0 1 4553
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1707688321
transform 1 0 19796 0 1 3862
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1707688321
transform 1 0 15432 0 1 3862
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1707688321
transform 1 0 15744 0 1 3862
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1707688321
transform 1 0 16056 0 1 3862
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1707688321
transform 1 0 16368 0 1 3862
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1707688321
transform 1 0 12232 0 1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1707688321
transform 1 0 11718 0 1 4391
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1707688321
transform 1 0 12990 0 1 4155
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1707688321
transform 0 -1 12402 1 0 4851
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 17412 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 17100 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 14524 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 -1 14212 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 -1 14836 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 13900 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 12338 -1 0 5441
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 13226 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1707688321
transform -1 0 13332 0 1 4568
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1707688321
transform 0 -1 19746 1 0 3638
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1707688321
transform 0 -1 20000 1 0 3638
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_11
timestamp 1707688321
transform 1 0 12841 0 1 4845
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform 1 0 11623 0 1 4155
box -12 -6 766 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 1 0 19591 0 1 4155
box 0 0 1 1
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_0
timestamp 1707688321
transform 0 -1 12994 -1 0 3816
box -12 -6 190 184
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_1
timestamp 1707688321
transform 0 1 17956 -1 0 3816
box -12 -6 190 184
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_2
timestamp 1707688321
transform 0 1 15068 -1 0 3816
box -12 -6 190 184
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_3
timestamp 1707688321
transform 0 1 16657 -1 0 3816
box -12 -6 190 184
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_4
timestamp 1707688321
transform 0 1 13498 1 0 3638
box -12 -6 190 184
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1707688321
transform 0 1 17640 -1 0 3816
box 0 0 1 1
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform -1 0 17944 0 1 3026
box -12 -6 1126 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_1
timestamp 1707688321
transform -1 0 16515 0 1 3032
box -12 -6 1126 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_2
timestamp 1707688321
transform 1 0 13951 0 1 3032
box -12 -6 1126 40
use L1M1_CDNS_52468879185336  L1M1_CDNS_52468879185336_0
timestamp 1707688321
transform 1 0 17719 0 1 4304
box -12 -6 1558 40
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1707688321
transform 1 0 11538 0 1 4771
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_1
timestamp 1707688321
transform 1 0 11538 0 1 4629
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 1 13292 -1 0 3598
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 12600 0 1 3856
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 17858 0 1 3020
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform -1 0 11651 0 1 3386
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform -1 0 13264 0 1 4143
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform -1 0 13264 0 1 3020
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform -1 0 11740 0 1 4543
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform -1 0 11740 0 1 3466
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform -1 0 12600 0 1 4381
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform -1 0 13344 0 1 4556
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform -1 0 11651 0 1 3546
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform -1 0 11651 0 1 4623
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform 1 0 17730 0 1 3330
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform 1 0 13292 0 1 3020
box 0 0 1 1
use nfet_CDNS_52468879185342  nfet_CDNS_52468879185342_0
timestamp 1707688321
transform -1 0 13253 0 1 4311
box -79 -26 199 226
use nfet_CDNS_52468879185342  nfet_CDNS_52468879185342_1
timestamp 1707688321
transform 1 0 12605 0 1 4311
box -79 -26 199 226
use nfet_CDNS_52468879185342  nfet_CDNS_52468879185342_2
timestamp 1707688321
transform 1 0 12957 0 1 4311
box -79 -26 199 226
use nfet_CDNS_52468879185342  nfet_CDNS_52468879185342_3
timestamp 1707688321
transform 1 0 13309 0 1 4311
box -79 -26 199 226
use nfet_CDNS_52468879185343  nfet_CDNS_52468879185343_0
timestamp 1707688321
transform 0 1 12406 -1 0 4804
box -79 -26 199 1026
use nfet_CDNS_52468879185343  nfet_CDNS_52468879185343_1
timestamp 1707688321
transform -1 0 12293 0 1 4573
box -79 -26 199 1026
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_0
timestamp 1707688321
transform 0 -1 12060 -1 0 4784
box -79 -26 179 626
use nfet_CDNS_52468879185345  nfet_CDNS_52468879185345_0
timestamp 1707688321
transform 1 0 11581 0 1 4311
box -79 -26 535 226
use nfet_CDNS_52468879185346  nfet_CDNS_52468879185346_0
timestamp 1707688321
transform -1 0 12901 0 1 4311
box -79 -26 199 226
use nfet_CDNS_52468879185347  nfet_CDNS_52468879185347_0
timestamp 1707688321
transform 1 0 12093 0 1 4311
box -79 -26 535 226
use nfet_CDNS_52468879185348  nfet_CDNS_52468879185348_0
timestamp 1707688321
transform 0 -1 12662 1 0 3225
box -79 -26 879 110
use nfet_CDNS_52468879185350  nfet_CDNS_52468879185350_0
timestamp 1707688321
transform 0 -1 12518 -1 0 4025
box -79 -26 879 110
use pfet_CDNS_52468879185351  pfet_CDNS_52468879185351_0
timestamp 1707688321
transform -1 0 17991 0 -1 4078
box -119 -66 1311 1066
use pfet_CDNS_52468879185351  pfet_CDNS_52468879185351_1
timestamp 1707688321
transform 1 0 15355 0 -1 4078
box -119 -66 1311 1066
use pfet_CDNS_52468879185351  pfet_CDNS_52468879185351_2
timestamp 1707688321
transform 1 0 13911 0 -1 4078
box -119 -66 1311 1066
use pfet_CDNS_52468879185352  pfet_CDNS_52468879185352_0
timestamp 1707688321
transform -1 0 13855 0 -1 4078
box -119 -66 219 1066
use pfet_CDNS_52468879185352  pfet_CDNS_52468879185352_1
timestamp 1707688321
transform -1 0 19701 0 -1 4078
box -119 -66 219 1066
use pfet_CDNS_52468879185352  pfet_CDNS_52468879185352_2
timestamp 1707688321
transform 1 0 19757 0 -1 4078
box -119 -66 219 1066
use pfet_CDNS_52468879185353  pfet_CDNS_52468879185353_0
timestamp 1707688321
transform 0 -1 12990 1 0 3225
box -119 -66 919 150
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_0
timestamp 1707688321
transform 1 0 18243 0 -1 4078
box -119 -66 687 1066
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_1
timestamp 1707688321
transform 1 0 18867 0 -1 4078
box -119 -66 687 1066
use pfet_CDNS_52468879185356  pfet_CDNS_52468879185356_0
timestamp 1707688321
transform -1 0 13503 0 -1 4073
box -119 -66 375 266
use pfet_CDNS_52468879185357  pfet_CDNS_52468879185357_0
timestamp 1707688321
transform 1 0 17679 0 -1 4256
box -119 -66 1719 150
use pfet_CDNS_52468879185358  pfet_CDNS_52468879185358_0
timestamp 1707688321
transform 1 0 13119 0 -1 3678
box -119 -66 216 666
use pfet_CDNS_52468879185359  pfet_CDNS_52468879185359_0
timestamp 1707688321
transform 1 0 13261 0 -1 3678
box -116 -66 216 666
use pfet_CDNS_52468879185360  pfet_CDNS_52468879185360_0
timestamp 1707688321
transform 1 0 13403 0 -1 3678
box -116 -66 219 666
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 1 0 13244 0 1 3739
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 13429 -1 0 4279
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 -1 13855 -1 0 3046
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 -1 13202 -1 0 3046
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 -1 13091 -1 0 4279
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 -1 12739 -1 0 4279
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 1 13420 -1 0 3046
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 -1 13256 1 0 4543
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 -1 12904 1 0 4543
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 0 -1 12293 1 0 5605
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1707688321
transform 1 0 11368 0 -1 4786
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1707688321
transform 1 0 13438 0 -1 4804
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 -1 13357 1 0 4105
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 1 19583 1 0 4110
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1707688321
transform 1 0 13022 0 -1 4025
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1707688321
transform -1 0 12402 0 1 3252
box 0 0 66 746
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 -1 19423 -1 0 3046
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1707688321
transform 0 -1 18799 -1 0 3046
box 0 0 66 542
use PYL1_CDNS_52468879185330  PYL1_CDNS_52468879185330_0
timestamp 1707688321
transform 0 -1 19265 -1 0 4354
box 0 0 66 1562
use PYL1_CDNS_52468879185331  PYL1_CDNS_52468879185331_0
timestamp 1707688321
transform 0 -1 17971 -1 0 3046
box 0 0 66 1154
use PYL1_CDNS_52468879185331  PYL1_CDNS_52468879185331_1
timestamp 1707688321
transform 0 -1 16527 -1 0 3046
box 0 0 66 1154
use PYL1_CDNS_52468879185331  PYL1_CDNS_52468879185331_2
timestamp 1707688321
transform 0 -1 15082 -1 0 3046
box 0 0 66 1154
use PYL1_CDNS_52468879185332  PYL1_CDNS_52468879185332_0
timestamp 1707688321
transform 0 1 11590 -1 0 4279
box 0 0 66 814
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_0
timestamp 1707688321
transform -1 0 15444 0 1 3026
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851416  sky130_fd_io__sio_tk_em1o_CDNS_524688791851416_0
timestamp 1707688321
transform 0 -1 12023 -1 0 4792
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851417  sky130_fd_io__sio_tk_em1o_CDNS_524688791851417_0
timestamp 1707688321
transform -1 0 13342 0 1 3470
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1707688321
transform 1 0 11628 0 1 3386
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1707688321
transform 1 0 11787 0 1 4381
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_0
timestamp 1707688321
transform 1 0 16744 0 1 3552
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851418  sky130_fd_io__sio_tk_em1s_CDNS_524688791851418_0
timestamp 1707688321
transform 0 -1 13002 1 0 3881
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851418  sky130_fd_io__sio_tk_em1s_CDNS_524688791851418_1
timestamp 1707688321
transform 0 -1 12686 1 0 4032
box 0 0 1 1
<< labels >>
flabel comment s 12105 3483 12105 3483 0 FreeSans 300 180 0 0 net157 of I31
flabel comment s 12082 3895 12082 3895 0 FreeSans 300 0 0 0 pbias
flabel comment s 15965 3895 15965 3895 0 FreeSans 300 0 0 0 pbias
flabel comment s 18462 3871 18462 3871 0 FreeSans 300 180 0 0 pbias
flabel comment s 13061 3380 13061 3380 0 FreeSans 300 90 0 0 bias_g
flabel comment s 16136 3566 16136 3566 0 FreeSans 300 180 0 0 pbias1
flabel comment s 18593 3455 18593 3455 0 FreeSans 300 0 0 0 net157
flabel comment s 19225 3369 19225 3369 0 FreeSans 300 0 0 0 2vtp
flabel comment s 19076 3586 19076 3586 0 FreeSans 300 0 0 0 net161
flabel comment s 19723 4170 19723 4170 0 FreeSans 300 0 0 0 drvlo_i_h
flabel comment s 19133 2989 19133 2989 0 FreeSans 300 0 0 0 net161 gt & dr tied
flabel comment s 18516 2989 18516 2989 0 FreeSans 300 0 0 0 net157 gt & dr tied
flabel comment s 17404 2982 17404 2982 0 FreeSans 300 0 0 0 2vtp
flabel comment s 15914 2974 15914 2974 0 FreeSans 300 180 0 0 pbias
flabel comment s 14349 2974 14349 2974 0 FreeSans 300 180 0 0 pbias1
flabel comment s 13319 3721 13319 3721 0 FreeSans 300 180 0 0 n<0>
flabel comment s 12838 4609 12838 4609 0 FreeSans 300 0 0 0 pden_h_n
flabel comment s 13205 4614 13205 4614 0 FreeSans 300 0 0 0 en_h_n
flabel comment s 13067 4540 13067 4540 0 FreeSans 300 270 0 0 bias_g
flabel comment s 12749 4500 12749 4500 0 FreeSans 300 180 0 0 n<1>
flabel comment s 12201 4397 12201 4397 0 FreeSans 300 180 0 0 pbias
flabel comment s 11805 4403 11805 4403 0 FreeSans 300 180 0 0 m1 opt to pbias
flabel comment s 12114 4991 12114 4991 0 FreeSans 300 90 0 0 net157 of I31
flabel comment s 12221 5593 12221 5593 0 FreeSans 300 0 0 0 bias_g
flabel comment s 11491 4653 11491 4653 0 FreeSans 300 180 0 0 n<0>
flabel comment s 11514 4821 11514 4821 0 FreeSans 300 180 0 0 n<1>
flabel comment s 12740 3563 12740 3563 0 FreeSans 300 180 0 0 n<0>
flabel comment s 13500 4753 13500 4753 0 FreeSans 300 90 0 0 n<1>
flabel comment s 13765 4162 13765 4162 0 FreeSans 300 180 0 0 drvlo_i_h
flabel comment s 13215 4218 13215 4218 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 12922 4076 12922 4076 0 FreeSans 300 0 0 0 m1 opt to pbias
flabel comment s 12950 3166 12950 3166 0 FreeSans 300 0 0 0 vcc_io
flabel comment s 11940 4227 11940 4227 0 FreeSans 300 0 0 0 bias_g
flabel comment s 12545 4128 12545 4128 0 FreeSans 300 0 0 0 m1 opt to bias_g
flabel comment s 13078 3951 13078 3951 0 FreeSans 300 90 0 0 bias_g
flabel comment s 19328 4220 19328 4220 0 FreeSans 300 90 0 0 2vtp
flabel comment s 17627 4233 17627 4233 0 FreeSans 300 90 0 0 vcc_io
flabel comment s 18487 4363 18487 4363 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 13808 3895 13808 3895 0 FreeSans 300 0 0 0 pbias
flabel metal1 s 12352 3401 12386 3435 7 FreeSans 300 180 0 0 pd_h
port 1 nsew
flabel metal1 s 13475 4636 13508 4682 3 FreeSans 300 0 0 0 pden_h_n
port 2 nsew
flabel metal1 s 13510 3020 13554 3072 3 FreeSans 300 0 0 0 en_h_n
port 3 nsew
flabel metal1 s 13068 3020 13113 3072 8 FreeSans 300 0 0 0 drvlo_h_n
port 7 nsew
flabel metal1 s 19927 3856 19963 3908 8 FreeSans 300 180 0 0 pbias
port 4 nsew
flabel metal1 s 11428 3856 11464 3908 3 FreeSans 300 180 0 0 pbias
port 4 nsew
flabel metal1 s 11364 3626 11400 3828 3 FreeSans 300 180 0 0 vcc_io
port 5 nsew
flabel metal1 s 11364 3100 11400 3302 3 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 20032 3100 20068 3302 7 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 13475 4839 13508 4969 7 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 13475 5251 13508 5453 7 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 11364 4839 11400 4969 3 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 11364 5251 11400 5453 3 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 20032 3626 20068 3828 7 FreeSans 300 180 0 0 vcc_io
port 5 nsew
flabel metal1 s 20032 4223 20068 4353 7 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel metal1 s 11364 4223 11400 4353 3 FreeSans 300 180 0 0 vgnd_io
port 6 nsew
flabel locali s 13805 2996 13855 3030 7 FreeSans 300 0 0 0 en_h
port 8 nsew
<< properties >>
string GDS_END 87921296
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87892196
<< end >>
