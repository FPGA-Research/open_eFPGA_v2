magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 37 41 311 203
rect 37 17 63 41
rect 29 -17 63 17
<< locali >>
rect 29 199 120 333
rect 162 150 247 491
rect 162 63 289 150
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 45 525 348 527
rect 45 367 111 525
rect 288 291 348 525
rect 59 17 125 149
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 29 199 120 333 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 368 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 3 nsew ground bidirectional
rlabel pwell s 37 17 63 41 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 37 41 311 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 162 63 289 150 6 Y
port 6 nsew signal output
rlabel locali s 162 150 247 491 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3339856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3336266
<< end >>
