magic
tech sky130B
timestamp 1707688321
<< poly >>
rect 0 1623 33 1631
rect 0 1606 8 1623
rect 25 1606 33 1623
rect 0 1589 33 1606
rect 0 1572 8 1589
rect 25 1572 33 1589
rect 0 1555 33 1572
rect 0 1538 8 1555
rect 25 1538 33 1555
rect 0 1521 33 1538
rect 0 1504 8 1521
rect 25 1504 33 1521
rect 0 1487 33 1504
rect 0 1470 8 1487
rect 25 1470 33 1487
rect 0 1453 33 1470
rect 0 1436 8 1453
rect 25 1436 33 1453
rect 0 1419 33 1436
rect 0 1402 8 1419
rect 25 1402 33 1419
rect 0 1385 33 1402
rect 0 1368 8 1385
rect 25 1368 33 1385
rect 0 1351 33 1368
rect 0 1334 8 1351
rect 25 1334 33 1351
rect 0 1317 33 1334
rect 0 1300 8 1317
rect 25 1300 33 1317
rect 0 1283 33 1300
rect 0 1266 8 1283
rect 25 1266 33 1283
rect 0 1249 33 1266
rect 0 1232 8 1249
rect 25 1232 33 1249
rect 0 1215 33 1232
rect 0 1198 8 1215
rect 25 1198 33 1215
rect 0 1181 33 1198
rect 0 1164 8 1181
rect 25 1164 33 1181
rect 0 1147 33 1164
rect 0 1130 8 1147
rect 25 1130 33 1147
rect 0 1113 33 1130
rect 0 1096 8 1113
rect 25 1096 33 1113
rect 0 1079 33 1096
rect 0 1062 8 1079
rect 25 1062 33 1079
rect 0 1045 33 1062
rect 0 1028 8 1045
rect 25 1028 33 1045
rect 0 1011 33 1028
rect 0 994 8 1011
rect 25 994 33 1011
rect 0 977 33 994
rect 0 960 8 977
rect 25 960 33 977
rect 0 943 33 960
rect 0 926 8 943
rect 25 926 33 943
rect 0 909 33 926
rect 0 892 8 909
rect 25 892 33 909
rect 0 875 33 892
rect 0 858 8 875
rect 25 858 33 875
rect 0 841 33 858
rect 0 824 8 841
rect 25 824 33 841
rect 0 807 33 824
rect 0 790 8 807
rect 25 790 33 807
rect 0 773 33 790
rect 0 756 8 773
rect 25 756 33 773
rect 0 739 33 756
rect 0 722 8 739
rect 25 722 33 739
rect 0 705 33 722
rect 0 688 8 705
rect 25 688 33 705
rect 0 671 33 688
rect 0 654 8 671
rect 25 654 33 671
rect 0 637 33 654
rect 0 620 8 637
rect 25 620 33 637
rect 0 603 33 620
rect 0 586 8 603
rect 25 586 33 603
rect 0 569 33 586
rect 0 552 8 569
rect 25 552 33 569
rect 0 535 33 552
rect 0 518 8 535
rect 25 518 33 535
rect 0 501 33 518
rect 0 484 8 501
rect 25 484 33 501
rect 0 467 33 484
rect 0 450 8 467
rect 25 450 33 467
rect 0 433 33 450
rect 0 416 8 433
rect 25 416 33 433
rect 0 399 33 416
rect 0 382 8 399
rect 25 382 33 399
rect 0 365 33 382
rect 0 348 8 365
rect 25 348 33 365
rect 0 331 33 348
rect 0 314 8 331
rect 25 314 33 331
rect 0 297 33 314
rect 0 280 8 297
rect 25 280 33 297
rect 0 263 33 280
rect 0 246 8 263
rect 25 246 33 263
rect 0 229 33 246
rect 0 212 8 229
rect 25 212 33 229
rect 0 195 33 212
rect 0 178 8 195
rect 25 178 33 195
rect 0 161 33 178
rect 0 144 8 161
rect 25 144 33 161
rect 0 127 33 144
rect 0 110 8 127
rect 25 110 33 127
rect 0 93 33 110
rect 0 76 8 93
rect 25 76 33 93
rect 0 59 33 76
rect 0 42 8 59
rect 25 42 33 59
rect 0 25 33 42
rect 0 8 8 25
rect 25 8 33 25
rect 0 0 33 8
<< polycont >>
rect 8 1606 25 1623
rect 8 1572 25 1589
rect 8 1538 25 1555
rect 8 1504 25 1521
rect 8 1470 25 1487
rect 8 1436 25 1453
rect 8 1402 25 1419
rect 8 1368 25 1385
rect 8 1334 25 1351
rect 8 1300 25 1317
rect 8 1266 25 1283
rect 8 1232 25 1249
rect 8 1198 25 1215
rect 8 1164 25 1181
rect 8 1130 25 1147
rect 8 1096 25 1113
rect 8 1062 25 1079
rect 8 1028 25 1045
rect 8 994 25 1011
rect 8 960 25 977
rect 8 926 25 943
rect 8 892 25 909
rect 8 858 25 875
rect 8 824 25 841
rect 8 790 25 807
rect 8 756 25 773
rect 8 722 25 739
rect 8 688 25 705
rect 8 654 25 671
rect 8 620 25 637
rect 8 586 25 603
rect 8 552 25 569
rect 8 518 25 535
rect 8 484 25 501
rect 8 450 25 467
rect 8 416 25 433
rect 8 382 25 399
rect 8 348 25 365
rect 8 314 25 331
rect 8 280 25 297
rect 8 246 25 263
rect 8 212 25 229
rect 8 178 25 195
rect 8 144 25 161
rect 8 110 25 127
rect 8 76 25 93
rect 8 42 25 59
rect 8 8 25 25
<< locali >>
rect 8 1623 25 1631
rect 8 1589 25 1606
rect 8 1555 25 1572
rect 8 1521 25 1538
rect 8 1487 25 1504
rect 8 1453 25 1470
rect 8 1419 25 1436
rect 8 1385 25 1402
rect 8 1351 25 1368
rect 8 1317 25 1334
rect 8 1283 25 1300
rect 8 1249 25 1266
rect 8 1215 25 1232
rect 8 1181 25 1198
rect 8 1147 25 1164
rect 8 1113 25 1130
rect 8 1079 25 1096
rect 8 1045 25 1062
rect 8 1011 25 1028
rect 8 977 25 994
rect 8 943 25 960
rect 8 909 25 926
rect 8 875 25 892
rect 8 841 25 858
rect 8 807 25 824
rect 8 773 25 790
rect 8 739 25 756
rect 8 705 25 722
rect 8 671 25 688
rect 8 637 25 654
rect 8 603 25 620
rect 8 569 25 586
rect 8 535 25 552
rect 8 501 25 518
rect 8 467 25 484
rect 8 433 25 450
rect 8 399 25 416
rect 8 365 25 382
rect 8 331 25 348
rect 8 297 25 314
rect 8 263 25 280
rect 8 229 25 246
rect 8 195 25 212
rect 8 161 25 178
rect 8 127 25 144
rect 8 93 25 110
rect 8 59 25 76
rect 8 25 25 42
rect 8 0 25 8
<< properties >>
string GDS_END 88596418
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88593150
<< end >>
