magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 1946
rect 61 0 64 1946
<< via1 >>
rect 3 0 61 1946
<< metal2 >>
rect 0 0 3 1946
rect 61 0 64 1946
<< properties >>
string GDS_END 89707108
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89699168
<< end >>
