magic
tech sky130B
timestamp 1707688321
<< pwell >>
rect -13 -13 54 1618
<< psubdiff >>
rect 0 1593 41 1605
rect 0 1576 12 1593
rect 29 1576 41 1593
rect 0 1559 41 1576
rect 0 1542 12 1559
rect 29 1542 41 1559
rect 0 1525 41 1542
rect 0 1508 12 1525
rect 29 1508 41 1525
rect 0 1491 41 1508
rect 0 1474 12 1491
rect 29 1474 41 1491
rect 0 1457 41 1474
rect 0 1440 12 1457
rect 29 1440 41 1457
rect 0 1423 41 1440
rect 0 1406 12 1423
rect 29 1406 41 1423
rect 0 1389 41 1406
rect 0 1372 12 1389
rect 29 1372 41 1389
rect 0 1355 41 1372
rect 0 1338 12 1355
rect 29 1338 41 1355
rect 0 1321 41 1338
rect 0 1304 12 1321
rect 29 1304 41 1321
rect 0 1287 41 1304
rect 0 1270 12 1287
rect 29 1270 41 1287
rect 0 1253 41 1270
rect 0 1236 12 1253
rect 29 1236 41 1253
rect 0 1219 41 1236
rect 0 1202 12 1219
rect 29 1202 41 1219
rect 0 1185 41 1202
rect 0 1168 12 1185
rect 29 1168 41 1185
rect 0 1151 41 1168
rect 0 1134 12 1151
rect 29 1134 41 1151
rect 0 1117 41 1134
rect 0 1100 12 1117
rect 29 1100 41 1117
rect 0 1083 41 1100
rect 0 1066 12 1083
rect 29 1066 41 1083
rect 0 1049 41 1066
rect 0 1032 12 1049
rect 29 1032 41 1049
rect 0 1015 41 1032
rect 0 998 12 1015
rect 29 998 41 1015
rect 0 981 41 998
rect 0 964 12 981
rect 29 964 41 981
rect 0 947 41 964
rect 0 930 12 947
rect 29 930 41 947
rect 0 913 41 930
rect 0 896 12 913
rect 29 896 41 913
rect 0 879 41 896
rect 0 862 12 879
rect 29 862 41 879
rect 0 845 41 862
rect 0 828 12 845
rect 29 828 41 845
rect 0 811 41 828
rect 0 794 12 811
rect 29 794 41 811
rect 0 777 41 794
rect 0 760 12 777
rect 29 760 41 777
rect 0 743 41 760
rect 0 726 12 743
rect 29 726 41 743
rect 0 709 41 726
rect 0 692 12 709
rect 29 692 41 709
rect 0 675 41 692
rect 0 658 12 675
rect 29 658 41 675
rect 0 641 41 658
rect 0 624 12 641
rect 29 624 41 641
rect 0 607 41 624
rect 0 590 12 607
rect 29 590 41 607
rect 0 573 41 590
rect 0 556 12 573
rect 29 556 41 573
rect 0 539 41 556
rect 0 522 12 539
rect 29 522 41 539
rect 0 505 41 522
rect 0 488 12 505
rect 29 488 41 505
rect 0 471 41 488
rect 0 454 12 471
rect 29 454 41 471
rect 0 437 41 454
rect 0 420 12 437
rect 29 420 41 437
rect 0 403 41 420
rect 0 386 12 403
rect 29 386 41 403
rect 0 369 41 386
rect 0 352 12 369
rect 29 352 41 369
rect 0 335 41 352
rect 0 318 12 335
rect 29 318 41 335
rect 0 301 41 318
rect 0 284 12 301
rect 29 284 41 301
rect 0 267 41 284
rect 0 250 12 267
rect 29 250 41 267
rect 0 233 41 250
rect 0 216 12 233
rect 29 216 41 233
rect 0 199 41 216
rect 0 182 12 199
rect 29 182 41 199
rect 0 165 41 182
rect 0 148 12 165
rect 29 148 41 165
rect 0 131 41 148
rect 0 114 12 131
rect 29 114 41 131
rect 0 97 41 114
rect 0 80 12 97
rect 29 80 41 97
rect 0 63 41 80
rect 0 46 12 63
rect 29 46 41 63
rect 0 29 41 46
rect 0 12 12 29
rect 29 12 41 29
rect 0 0 41 12
<< psubdiffcont >>
rect 12 1576 29 1593
rect 12 1542 29 1559
rect 12 1508 29 1525
rect 12 1474 29 1491
rect 12 1440 29 1457
rect 12 1406 29 1423
rect 12 1372 29 1389
rect 12 1338 29 1355
rect 12 1304 29 1321
rect 12 1270 29 1287
rect 12 1236 29 1253
rect 12 1202 29 1219
rect 12 1168 29 1185
rect 12 1134 29 1151
rect 12 1100 29 1117
rect 12 1066 29 1083
rect 12 1032 29 1049
rect 12 998 29 1015
rect 12 964 29 981
rect 12 930 29 947
rect 12 896 29 913
rect 12 862 29 879
rect 12 828 29 845
rect 12 794 29 811
rect 12 760 29 777
rect 12 726 29 743
rect 12 692 29 709
rect 12 658 29 675
rect 12 624 29 641
rect 12 590 29 607
rect 12 556 29 573
rect 12 522 29 539
rect 12 488 29 505
rect 12 454 29 471
rect 12 420 29 437
rect 12 386 29 403
rect 12 352 29 369
rect 12 318 29 335
rect 12 284 29 301
rect 12 250 29 267
rect 12 216 29 233
rect 12 182 29 199
rect 12 148 29 165
rect 12 114 29 131
rect 12 80 29 97
rect 12 46 29 63
rect 12 12 29 29
<< locali >>
rect 12 1593 29 1601
rect 12 1559 29 1576
rect 12 1525 29 1542
rect 12 1491 29 1508
rect 12 1457 29 1474
rect 12 1423 29 1440
rect 12 1389 29 1406
rect 12 1355 29 1372
rect 12 1321 29 1338
rect 12 1287 29 1304
rect 12 1253 29 1270
rect 12 1219 29 1236
rect 12 1185 29 1202
rect 12 1151 29 1168
rect 12 1117 29 1134
rect 12 1083 29 1100
rect 12 1049 29 1066
rect 12 1015 29 1032
rect 12 981 29 998
rect 12 947 29 964
rect 12 913 29 930
rect 12 879 29 896
rect 12 845 29 862
rect 12 811 29 828
rect 12 777 29 794
rect 12 743 29 760
rect 12 709 29 726
rect 12 675 29 692
rect 12 641 29 658
rect 12 607 29 624
rect 12 573 29 590
rect 12 539 29 556
rect 12 505 29 522
rect 12 471 29 488
rect 12 437 29 454
rect 12 403 29 420
rect 12 369 29 386
rect 12 335 29 352
rect 12 301 29 318
rect 12 267 29 284
rect 12 233 29 250
rect 12 199 29 216
rect 12 165 29 182
rect 12 131 29 148
rect 12 97 29 114
rect 12 63 29 80
rect 12 29 29 46
rect 12 4 29 12
<< properties >>
string GDS_END 42949400
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42946196
<< end >>
