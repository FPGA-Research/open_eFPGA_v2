magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 1640 839 3459 1311
rect -175 -753 3459 839
<< nwell >>
rect 1294 3005 1589 3047
rect 1264 2873 1619 3005
rect 1294 2831 1589 2873
rect 760 2511 1589 2831
rect 2141 2531 2263 3243
rect 1560 1161 3539 1391
rect 0 1105 3539 1161
rect 0 681 1846 1105
rect 3253 -217 3539 1105
<< nsubdiff >>
rect 1640 1231 1679 1265
rect 1713 1231 1747 1265
rect 1781 1231 1815 1265
rect 1849 1231 1883 1265
rect 1917 1231 1951 1265
rect 1985 1231 2019 1265
rect 2053 1231 2087 1265
rect 2121 1231 2155 1265
rect 2189 1231 2223 1265
rect 2257 1231 2291 1265
rect 2325 1231 2359 1265
rect 2393 1231 2427 1265
rect 2461 1231 2495 1265
rect 2529 1231 2563 1265
rect 2597 1231 2631 1265
rect 2665 1231 2699 1265
rect 2733 1231 2767 1265
rect 2801 1231 2835 1265
rect 2869 1231 2903 1265
rect 2937 1231 2971 1265
rect 3005 1231 3039 1265
rect 3073 1231 3107 1265
rect 3141 1231 3175 1265
rect 3209 1231 3243 1265
rect 3277 1231 3311 1265
rect 3345 1231 3413 1265
rect 3379 1143 3413 1231
rect 3379 1075 3413 1109
rect 3379 1007 3413 1041
rect 3379 939 3413 973
rect 3379 871 3413 905
rect 3379 803 3413 837
rect 3379 735 3413 769
rect 3379 667 3413 701
rect 3379 599 3413 633
rect 3379 531 3413 565
rect 3379 463 3413 497
rect 3379 395 3413 429
rect 3379 327 3413 361
rect 3379 259 3413 293
rect 3379 191 3413 225
rect 3379 123 3413 157
rect 3379 55 3413 89
rect 3379 -13 3413 21
rect 3379 -81 3413 -47
rect 3379 -149 3413 -115
rect 3379 -217 3413 -183
<< mvnsubdiff >>
rect 2177 3094 2227 3171
rect 2177 3060 2185 3094
rect 2219 3060 2227 3094
rect 2177 3026 2227 3060
rect 2177 2992 2185 3026
rect 2219 2992 2227 3026
rect 1300 2956 1583 2969
rect 1300 2922 1324 2956
rect 1358 2922 1392 2956
rect 1426 2922 1460 2956
rect 1494 2922 1583 2956
rect 1300 2909 1583 2922
rect 2177 2958 2227 2992
rect 2177 2924 2185 2958
rect 2219 2924 2227 2958
rect 2177 2890 2227 2924
rect 2177 2856 2185 2890
rect 2219 2856 2227 2890
rect 2177 2822 2227 2856
rect 2177 2788 2185 2822
rect 2219 2788 2227 2822
rect 2177 2754 2227 2788
rect 2177 2720 2185 2754
rect 2219 2720 2227 2754
rect 2177 2686 2227 2720
rect 2177 2652 2185 2686
rect 2219 2652 2227 2686
rect 2177 2603 2227 2652
<< nsubdiffcont >>
rect 2185 3060 2219 3094
rect 2185 2992 2219 3026
rect 2185 2924 2219 2958
rect 2185 2856 2219 2890
rect 2185 2788 2219 2822
rect 2185 2720 2219 2754
rect 2185 2652 2219 2686
rect 1679 1231 1713 1265
rect 1747 1231 1781 1265
rect 1815 1231 1849 1265
rect 1883 1231 1917 1265
rect 1951 1231 1985 1265
rect 2019 1231 2053 1265
rect 2087 1231 2121 1265
rect 2155 1231 2189 1265
rect 2223 1231 2257 1265
rect 2291 1231 2325 1265
rect 2359 1231 2393 1265
rect 2427 1231 2461 1265
rect 2495 1231 2529 1265
rect 2563 1231 2597 1265
rect 2631 1231 2665 1265
rect 2699 1231 2733 1265
rect 2767 1231 2801 1265
rect 2835 1231 2869 1265
rect 2903 1231 2937 1265
rect 2971 1231 3005 1265
rect 3039 1231 3073 1265
rect 3107 1231 3141 1265
rect 3175 1231 3209 1265
rect 3243 1231 3277 1265
rect 3311 1231 3345 1265
rect 3379 1109 3413 1143
rect 3379 1041 3413 1075
rect 3379 973 3413 1007
rect 3379 905 3413 939
rect 3379 837 3413 871
rect 3379 769 3413 803
rect 3379 701 3413 735
rect 3379 633 3413 667
rect 3379 565 3413 599
rect 3379 497 3413 531
rect 3379 429 3413 463
rect 3379 361 3413 395
rect 3379 293 3413 327
rect 3379 225 3413 259
rect 3379 157 3413 191
rect 3379 89 3413 123
rect 3379 21 3413 55
rect 3379 -47 3413 -13
rect 3379 -115 3413 -81
rect 3379 -183 3413 -149
<< mvnsubdiffcont >>
rect 1324 2922 1358 2956
rect 1392 2922 1426 2956
rect 1460 2922 1494 2956
<< poly >>
rect 865 3063 999 3079
rect 865 3029 881 3063
rect 915 3029 949 3063
rect 983 3029 999 3063
rect 865 3013 999 3029
rect 1055 2849 1189 2865
rect 1055 2815 1071 2849
rect 1105 2815 1139 2849
rect 1173 2815 1189 2849
rect 1055 2799 1189 2815
rect 1708 2529 2004 2545
rect 1708 2495 1724 2529
rect 1758 2495 1801 2529
rect 1835 2495 1878 2529
rect 1912 2495 1954 2529
rect 1988 2495 2004 2529
rect 1708 2479 2004 2495
rect 2404 2529 2700 2545
rect 2404 2495 2420 2529
rect 2454 2495 2496 2529
rect 2530 2495 2573 2529
rect 2607 2495 2650 2529
rect 2684 2495 2700 2529
rect 2404 2479 2700 2495
rect 2251 1077 2547 1093
rect 2251 1043 2267 1077
rect 2301 1043 2344 1077
rect 2378 1043 2421 1077
rect 2455 1043 2497 1077
rect 2531 1043 2547 1077
rect 2251 1027 2547 1043
rect 2603 1077 2899 1093
rect 2603 1043 2619 1077
rect 2653 1043 2696 1077
rect 2730 1043 2773 1077
rect 2807 1043 2849 1077
rect 2883 1043 2899 1077
rect 2603 1027 2899 1043
rect 119 847 415 863
rect 119 813 135 847
rect 169 813 212 847
rect 246 813 289 847
rect 323 813 365 847
rect 399 813 415 847
rect 119 797 415 813
rect 815 847 1111 863
rect 815 813 831 847
rect 865 813 907 847
rect 941 813 984 847
rect 1018 813 1061 847
rect 1095 813 1111 847
rect 815 797 1111 813
rect 295 576 415 797
rect 958 576 1078 797
rect 1331 677 1465 693
rect 1331 643 1347 677
rect 1381 643 1415 677
rect 1449 643 1465 677
rect 1331 627 1465 643
rect 1738 677 1872 693
rect 1738 643 1754 677
rect 1788 643 1822 677
rect 1856 643 1872 677
rect 1738 627 1872 643
<< polycont >>
rect 881 3029 915 3063
rect 949 3029 983 3063
rect 1071 2815 1105 2849
rect 1139 2815 1173 2849
rect 1724 2495 1758 2529
rect 1801 2495 1835 2529
rect 1878 2495 1912 2529
rect 1954 2495 1988 2529
rect 2420 2495 2454 2529
rect 2496 2495 2530 2529
rect 2573 2495 2607 2529
rect 2650 2495 2684 2529
rect 2267 1043 2301 1077
rect 2344 1043 2378 1077
rect 2421 1043 2455 1077
rect 2497 1043 2531 1077
rect 2619 1043 2653 1077
rect 2696 1043 2730 1077
rect 2773 1043 2807 1077
rect 2849 1043 2883 1077
rect 135 813 169 847
rect 212 813 246 847
rect 289 813 323 847
rect 365 813 399 847
rect 831 813 865 847
rect 907 813 941 847
rect 984 813 1018 847
rect 1061 813 1095 847
rect 1347 643 1381 677
rect 1415 643 1449 677
rect 1754 643 1788 677
rect 1822 643 1856 677
<< locali >>
rect 2117 3136 2291 3181
rect 865 3069 1255 3099
rect 865 3035 866 3069
rect 900 3063 938 3069
rect 972 3063 1255 3069
rect 915 3035 938 3063
rect 865 3029 881 3035
rect 915 3029 949 3035
rect 983 3029 1255 3063
rect 803 2942 894 2959
rect 803 2908 819 2942
rect 853 2908 894 2942
rect 803 2870 894 2908
rect 1010 2920 1044 2958
rect 1148 2893 1255 3029
rect 1663 3064 1697 3102
rect 1663 2992 1697 3030
rect 1300 2956 1583 2969
rect 1358 2922 1383 2956
rect 1426 2922 1460 2956
rect 1500 2922 1549 2956
rect 1300 2909 1583 2922
rect 1663 2920 1697 2958
rect 2049 3102 2101 3136
rect 2135 3102 2187 3136
rect 2221 3102 2273 3136
rect 2307 3102 2359 3136
rect 2015 3064 2393 3102
rect 2049 3030 2101 3064
rect 2135 3030 2187 3064
rect 2221 3030 2273 3064
rect 2307 3030 2359 3064
rect 2015 2992 2393 3030
rect 2049 2958 2101 2992
rect 2135 2958 2187 2992
rect 2221 2958 2273 2992
rect 2307 2958 2359 2992
rect 2015 2920 2393 2958
rect 2049 2886 2101 2920
rect 2135 2886 2187 2920
rect 2221 2886 2273 2920
rect 2307 2886 2359 2920
rect 2711 3064 2745 3102
rect 2711 2992 2745 3030
rect 2711 2920 2745 2958
rect 803 2836 819 2870
rect 853 2849 894 2870
rect 853 2836 1071 2849
rect 803 2815 1071 2836
rect 1105 2815 1139 2849
rect 1173 2815 1189 2849
rect 1839 2673 1873 2711
rect 2117 2627 2291 2886
rect 2535 2673 2569 2711
rect 2177 2603 2227 2627
rect 1698 2495 1724 2529
rect 1770 2495 1801 2529
rect 1835 2495 1878 2529
rect 1912 2495 1954 2529
rect 1988 2495 2004 2529
rect 2397 2495 2420 2529
rect 2469 2495 2496 2529
rect 2530 2495 2573 2529
rect 2607 2495 2650 2529
rect 2684 2495 2700 2529
rect 11 1542 74 1576
rect 108 1542 127 1576
rect 11 1504 127 1542
rect 11 1470 74 1504
rect 108 1470 127 1504
rect 11 1432 127 1470
rect 11 1398 74 1432
rect 108 1398 127 1432
rect 11 1360 127 1398
rect 11 1326 74 1360
rect 108 1326 127 1360
rect 11 897 127 1326
rect 460 1542 512 1576
rect 546 1542 598 1576
rect 632 1542 684 1576
rect 718 1542 770 1576
rect 426 1504 804 1542
rect 460 1470 512 1504
rect 546 1470 598 1504
rect 632 1470 684 1504
rect 718 1470 770 1504
rect 426 1432 804 1470
rect 460 1398 512 1432
rect 546 1398 598 1432
rect 632 1398 684 1432
rect 718 1398 770 1432
rect 426 1360 804 1398
rect 460 1326 512 1360
rect 546 1326 598 1360
rect 632 1326 684 1360
rect 718 1326 770 1360
rect 250 958 284 996
rect 426 897 804 1326
rect 1074 1542 1122 1576
rect 1156 1542 1190 1576
rect 1074 1504 1190 1542
rect 1074 1470 1122 1504
rect 1156 1470 1190 1504
rect 1074 1432 1190 1470
rect 1074 1398 1122 1432
rect 1156 1398 1190 1432
rect 1074 1360 1190 1398
rect 1074 1326 1122 1360
rect 1156 1326 1190 1360
rect 1074 1265 1190 1326
rect 1074 1231 1679 1265
rect 1713 1231 1747 1265
rect 1781 1231 1815 1265
rect 1849 1231 1883 1265
rect 1917 1231 1951 1265
rect 1985 1231 2019 1265
rect 2053 1231 2087 1265
rect 2121 1231 2155 1265
rect 2189 1231 2223 1265
rect 2257 1231 2291 1265
rect 2325 1231 2359 1265
rect 2393 1231 2427 1265
rect 2461 1231 2495 1265
rect 2529 1231 2563 1265
rect 2597 1231 2631 1265
rect 2665 1231 2699 1265
rect 2733 1231 2767 1265
rect 2801 1231 2835 1265
rect 2869 1231 2903 1265
rect 2937 1231 2971 1265
rect 3005 1231 3039 1265
rect 3073 1231 3107 1265
rect 3141 1231 3175 1265
rect 3209 1231 3243 1265
rect 3277 1231 3311 1265
rect 3345 1231 3413 1265
rect 946 958 980 996
rect 1074 897 1190 1231
rect 1310 1136 1348 1170
rect 1382 1136 2899 1152
rect 1276 1115 2899 1136
rect 2603 1077 2899 1115
rect 1329 1043 1367 1077
rect 1401 1043 2267 1077
rect 2301 1043 2344 1077
rect 2378 1043 2421 1077
rect 2455 1043 2497 1077
rect 2531 1043 2547 1077
rect 2603 1043 2619 1077
rect 2653 1043 2696 1077
rect 2730 1043 2773 1077
rect 2807 1043 2849 1077
rect 2883 1043 2899 1077
rect 3379 1143 3413 1231
rect 3379 1075 3413 1109
rect 3379 1007 3413 1041
rect 3379 939 3413 973
rect 3379 871 3413 905
rect 129 813 135 847
rect 201 813 212 847
rect 246 813 289 847
rect 323 813 365 847
rect 399 813 415 847
rect 801 813 831 847
rect 873 813 907 847
rect 941 813 984 847
rect 1018 813 1061 847
rect 1095 813 1111 847
rect 2383 769 2417 811
rect 2383 693 2417 735
rect 1331 643 1345 677
rect 1381 643 1415 677
rect 1451 643 1465 677
rect 1738 643 1750 677
rect 1788 643 1822 677
rect 1856 643 1872 677
rect 2383 617 2417 659
rect 250 523 284 561
rect 426 282 947 542
rect 1089 461 1123 499
rect 1292 461 1326 499
rect 1570 282 1630 545
rect 2383 541 2417 583
rect 2735 766 2769 811
rect 2735 687 2769 732
rect 2735 607 2769 653
rect 3379 803 3413 837
rect 3379 735 3413 769
rect 3379 667 3413 701
rect 3379 599 3413 633
rect 1874 461 1908 499
rect 2383 464 2417 507
rect 3379 531 3413 565
rect 3379 463 3413 497
rect 1874 389 1908 427
rect 3379 395 3413 429
rect 3379 327 3413 361
rect 460 248 536 282
rect 570 248 803 282
rect 837 248 913 282
rect 426 210 947 248
rect 460 176 536 210
rect 570 176 803 210
rect 837 176 913 210
rect 426 138 947 176
rect 460 104 536 138
rect 570 104 803 138
rect 837 104 913 138
rect 426 66 947 104
rect 460 32 536 66
rect 570 32 803 66
rect 837 32 913 66
rect 1468 248 1469 282
rect 1503 248 1545 282
rect 1579 248 1621 282
rect 1655 248 1697 282
rect 1731 248 1732 282
rect 1468 210 1732 248
rect 1468 176 1469 210
rect 1503 176 1545 210
rect 1579 176 1621 210
rect 1655 176 1697 210
rect 1731 176 1732 210
rect 1468 138 1732 176
rect 1468 104 1469 138
rect 1503 104 1545 138
rect 1579 104 1621 138
rect 1655 104 1697 138
rect 1731 104 1732 138
rect 1468 66 1732 104
rect 1468 32 1469 66
rect 1503 32 1545 66
rect 1579 32 1621 66
rect 1655 32 1697 66
rect 1731 32 1732 66
rect 2207 210 2241 248
rect 2207 138 2241 176
rect 2207 66 2241 104
rect 2559 210 2593 248
rect 2559 138 2593 176
rect 2559 66 2593 104
rect 2911 210 2945 248
rect 2911 138 2945 176
rect 2911 66 2945 104
rect 3379 259 3413 293
rect 3379 191 3413 225
rect 3379 123 3413 157
rect 3379 55 3413 89
rect 426 26 947 32
rect 3379 -13 3413 21
rect 3379 -81 3413 -47
rect 3379 -149 3413 -115
rect 3379 -217 3413 -183
<< viali >>
rect 1663 3102 1697 3136
rect 866 3063 900 3069
rect 938 3063 972 3069
rect 866 3035 881 3063
rect 881 3035 900 3063
rect 938 3035 949 3063
rect 949 3035 972 3063
rect 819 2908 853 2942
rect 1010 2958 1044 2992
rect 1010 2886 1044 2920
rect 1663 3030 1697 3064
rect 1300 2922 1324 2956
rect 1324 2922 1334 2956
rect 1383 2922 1392 2956
rect 1392 2922 1417 2956
rect 1466 2922 1494 2956
rect 1494 2922 1500 2956
rect 1549 2922 1583 2956
rect 1663 2958 1697 2992
rect 1663 2886 1697 2920
rect 2015 3102 2049 3136
rect 2101 3102 2135 3136
rect 2187 3102 2221 3136
rect 2273 3102 2307 3136
rect 2359 3102 2393 3136
rect 2015 3030 2049 3064
rect 2101 3030 2135 3064
rect 2187 3030 2221 3064
rect 2273 3030 2307 3064
rect 2359 3030 2393 3064
rect 2015 2958 2049 2992
rect 2101 2958 2135 2992
rect 2187 2958 2221 2992
rect 2273 2958 2307 2992
rect 2359 2958 2393 2992
rect 2015 2886 2049 2920
rect 2101 2886 2135 2920
rect 2187 2886 2221 2920
rect 2273 2886 2307 2920
rect 2359 2886 2393 2920
rect 2711 3102 2745 3136
rect 2711 3030 2745 3064
rect 2711 2958 2745 2992
rect 2711 2886 2745 2920
rect 819 2836 853 2870
rect 1839 2711 1873 2745
rect 1839 2639 1873 2673
rect 2535 2711 2569 2745
rect 2535 2639 2569 2673
rect 1664 2495 1698 2529
rect 1736 2495 1758 2529
rect 1758 2495 1770 2529
rect 2363 2495 2397 2529
rect 2435 2495 2454 2529
rect 2454 2495 2469 2529
rect 74 1542 108 1576
rect 74 1470 108 1504
rect 74 1398 108 1432
rect 74 1326 108 1360
rect 426 1542 460 1576
rect 512 1542 546 1576
rect 598 1542 632 1576
rect 684 1542 718 1576
rect 770 1542 804 1576
rect 426 1470 460 1504
rect 512 1470 546 1504
rect 598 1470 632 1504
rect 684 1470 718 1504
rect 770 1470 804 1504
rect 426 1398 460 1432
rect 512 1398 546 1432
rect 598 1398 632 1432
rect 684 1398 718 1432
rect 770 1398 804 1432
rect 426 1326 460 1360
rect 512 1326 546 1360
rect 598 1326 632 1360
rect 684 1326 718 1360
rect 770 1326 804 1360
rect 250 996 284 1030
rect 250 924 284 958
rect 1122 1542 1156 1576
rect 1122 1470 1156 1504
rect 1122 1398 1156 1432
rect 1122 1326 1156 1360
rect 946 996 980 1030
rect 946 924 980 958
rect 1276 1136 1310 1170
rect 1348 1136 1382 1170
rect 1295 1043 1329 1077
rect 1367 1043 1401 1077
rect 95 813 129 847
rect 167 813 169 847
rect 169 813 201 847
rect 767 813 801 847
rect 839 813 865 847
rect 865 813 873 847
rect 2383 811 2417 845
rect 2383 735 2417 769
rect 1345 643 1347 677
rect 1347 643 1379 677
rect 1417 643 1449 677
rect 1449 643 1451 677
rect 1750 643 1754 677
rect 1754 643 1784 677
rect 1822 643 1856 677
rect 2383 659 2417 693
rect 250 561 284 595
rect 2383 583 2417 617
rect 250 489 284 523
rect 1089 499 1123 533
rect 1089 427 1123 461
rect 1292 499 1326 533
rect 1292 427 1326 461
rect 2735 811 2769 845
rect 2735 732 2769 766
rect 2735 653 2769 687
rect 2735 573 2769 607
rect 1874 499 1908 533
rect 1874 427 1908 461
rect 2383 507 2417 541
rect 2383 430 2417 464
rect 1874 355 1908 389
rect 426 248 460 282
rect 536 248 570 282
rect 803 248 837 282
rect 913 248 947 282
rect 426 176 460 210
rect 536 176 570 210
rect 803 176 837 210
rect 913 176 947 210
rect 426 104 460 138
rect 536 104 570 138
rect 803 104 837 138
rect 913 104 947 138
rect 426 32 460 66
rect 536 32 570 66
rect 803 32 837 66
rect 913 32 947 66
rect 1469 248 1503 282
rect 1545 248 1579 282
rect 1621 248 1655 282
rect 1697 248 1731 282
rect 1469 176 1503 210
rect 1545 176 1579 210
rect 1621 176 1655 210
rect 1697 176 1731 210
rect 1469 104 1503 138
rect 1545 104 1579 138
rect 1621 104 1655 138
rect 1697 104 1731 138
rect 1469 32 1503 66
rect 1545 32 1579 66
rect 1621 32 1655 66
rect 1697 32 1731 66
rect 2207 248 2241 282
rect 2207 176 2241 210
rect 2207 104 2241 138
rect 2207 32 2241 66
rect 2559 248 2593 282
rect 2559 176 2593 210
rect 2559 104 2593 138
rect 2559 32 2593 66
rect 2911 248 2945 282
rect 2911 176 2945 210
rect 2911 104 2945 138
rect 2911 32 2945 66
<< metal1 >>
rect 1657 3136 2751 3148
rect 1657 3102 1663 3136
rect 1697 3102 2015 3136
rect 2049 3102 2101 3136
rect 2135 3102 2187 3136
rect 2221 3102 2273 3136
rect 2307 3102 2359 3136
rect 2393 3102 2711 3136
rect 2745 3102 2751 3136
rect 854 3069 984 3075
rect 854 3035 866 3069
rect 900 3035 938 3069
rect 972 3035 984 3069
rect 854 3029 984 3035
rect 1657 3064 2751 3102
rect 1657 3030 1663 3064
rect 1697 3030 2015 3064
rect 2049 3030 2101 3064
rect 2135 3030 2187 3064
rect 2221 3030 2273 3064
rect 2307 3030 2359 3064
rect 2393 3030 2711 3064
rect 2745 3030 2751 3064
rect 813 2942 859 2954
rect 813 2908 819 2942
rect 853 2908 859 2942
rect 813 2870 859 2908
rect 813 2836 819 2870
rect 853 2836 859 2870
rect 813 2789 859 2836
rect 926 2832 972 3029
rect 1657 3004 2751 3030
rect 1004 2992 2751 3004
rect 1004 2958 1010 2992
rect 1044 2958 1663 2992
rect 1697 2958 2015 2992
rect 2049 2958 2101 2992
rect 2135 2958 2187 2992
rect 2221 2958 2273 2992
rect 2307 2958 2359 2992
rect 2393 2958 2711 2992
rect 2745 2958 2751 2992
rect 1004 2956 2751 2958
rect 1004 2922 1300 2956
rect 1334 2922 1383 2956
rect 1417 2922 1466 2956
rect 1500 2922 1549 2956
rect 1583 2922 2751 2956
rect 1004 2920 2751 2922
rect 1004 2886 1010 2920
rect 1044 2886 1663 2920
rect 1697 2886 2015 2920
rect 2049 2886 2101 2920
rect 2135 2886 2187 2920
rect 2221 2886 2273 2920
rect 2307 2886 2359 2920
rect 2393 2886 2711 2920
rect 2745 2886 2751 2920
rect 1004 2874 2751 2886
tri 926 2824 934 2832 ne
rect 934 2824 972 2832
tri 972 2824 1000 2852 sw
tri 934 2819 939 2824 ne
rect 939 2819 1000 2824
tri 1000 2819 1005 2824 sw
tri 939 2809 949 2819 ne
rect 949 2809 1414 2819
tri 1414 2809 1424 2819 sw
tri 813 2765 837 2789 ne
rect 837 2765 859 2789
tri 859 2765 903 2809 sw
tri 949 2803 955 2809 ne
rect 955 2803 1424 2809
tri 1424 2803 1430 2809 sw
tri 955 2786 972 2803 ne
rect 972 2786 1430 2803
tri 972 2773 985 2786 ne
rect 985 2773 1430 2786
tri 1394 2765 1402 2773 ne
rect 1402 2765 1430 2773
tri 1430 2765 1468 2803 sw
tri 837 2745 857 2765 ne
rect 857 2745 903 2765
tri 903 2745 923 2765 sw
tri 1402 2745 1422 2765 ne
rect 1422 2745 1468 2765
tri 1468 2745 1488 2765 sw
rect 1833 2745 1879 2757
tri 857 2743 859 2745 ne
rect 859 2743 923 2745
tri 859 2711 891 2743 ne
rect 891 2711 923 2743
tri 923 2711 957 2745 sw
tri 1422 2737 1430 2745 ne
rect 1430 2737 1488 2745
tri 1488 2737 1496 2745 sw
tri 1430 2711 1456 2737 ne
rect 1456 2711 1496 2737
tri 1496 2711 1522 2737 sw
rect 1833 2711 1839 2745
rect 1873 2711 1879 2745
tri 891 2699 903 2711 ne
rect 903 2699 957 2711
tri 957 2699 969 2711 sw
tri 1456 2699 1468 2711 ne
rect 1468 2699 1522 2711
tri 1522 2699 1534 2711 sw
tri 903 2673 929 2699 ne
rect 929 2673 1338 2699
tri 1338 2673 1364 2699 sw
tri 1468 2673 1494 2699 ne
rect 1494 2673 1534 2699
tri 1534 2673 1560 2699 sw
rect 1833 2673 1879 2711
tri 929 2653 949 2673 ne
rect 949 2653 1364 2673
tri 1318 2645 1326 2653 ne
rect 1326 2645 1364 2653
tri 1364 2645 1392 2673 sw
tri 1494 2671 1496 2673 ne
rect 1496 2671 1560 2673
tri 1560 2671 1562 2673 sw
tri 1496 2651 1516 2671 ne
tri 1326 2639 1332 2645 ne
rect 1332 2639 1392 2645
tri 1392 2639 1398 2645 sw
tri 1332 2633 1338 2639 ne
rect 1338 2633 1398 2639
tri 1338 2579 1392 2633 ne
rect 1392 2627 1398 2633
tri 1398 2627 1410 2639 sw
rect 1392 2579 1410 2627
tri 1410 2579 1458 2627 sw
tri 1392 2559 1412 2579 ne
tri 1386 1739 1412 1765 se
rect 1412 1739 1458 2579
rect 1330 1687 1336 1739
rect 1388 1687 1400 1739
rect 1452 1687 1458 1739
rect 1516 2535 1562 2671
rect 1833 2639 1839 2673
rect 1873 2639 1879 2673
tri 1562 2535 1596 2569 sw
rect 1516 2529 1782 2535
rect 1516 2495 1664 2529
rect 1698 2495 1736 2529
rect 1770 2495 1782 2529
rect 1516 2489 1782 2495
rect 1516 2483 1582 2489
tri 1582 2483 1588 2489 nw
rect 1516 2477 1576 2483
tri 1576 2477 1582 2483 nw
rect 1516 2475 1574 2477
tri 1574 2475 1576 2477 nw
rect 1516 2469 1568 2475
tri 1568 2469 1574 2475 nw
rect 1516 1874 1562 2469
tri 1562 2463 1568 2469 nw
tri 1562 1874 1569 1881 sw
rect 1516 1867 1569 1874
tri 1569 1867 1576 1874 sw
rect 1516 1862 1576 1867
tri 1576 1862 1581 1867 sw
rect 1516 1855 1581 1862
tri 1581 1855 1588 1862 sw
rect 1516 1803 1522 1855
rect 1574 1803 1586 1855
rect 1638 1803 1644 1855
rect 1516 1796 1581 1803
tri 1581 1796 1588 1803 nw
rect 1516 1791 1576 1796
tri 1576 1791 1581 1796 nw
rect 1516 1784 1569 1791
tri 1569 1784 1576 1791 nw
rect 68 1576 1162 1588
rect 68 1542 74 1576
rect 108 1542 426 1576
rect 460 1542 512 1576
rect 546 1542 598 1576
rect 632 1542 684 1576
rect 718 1542 770 1576
rect 804 1542 1122 1576
rect 1156 1542 1162 1576
rect 68 1504 1162 1542
rect 68 1470 74 1504
rect 108 1470 426 1504
rect 460 1470 512 1504
rect 546 1470 598 1504
rect 632 1470 684 1504
rect 718 1470 770 1504
rect 804 1470 1122 1504
rect 1156 1470 1162 1504
rect 68 1432 1162 1470
rect 68 1398 74 1432
rect 108 1398 426 1432
rect 460 1398 512 1432
rect 546 1398 598 1432
rect 632 1398 684 1432
rect 718 1398 770 1432
rect 804 1398 1122 1432
rect 1156 1398 1162 1432
rect 68 1360 1162 1398
rect 68 1326 74 1360
rect 108 1326 426 1360
rect 460 1326 512 1360
rect 546 1326 598 1360
rect 632 1326 684 1360
rect 718 1326 770 1360
rect 804 1326 1122 1360
rect 1156 1326 1162 1360
rect 68 1314 1162 1326
tri 868 1170 874 1176 se
rect 874 1170 1394 1176
tri 834 1136 868 1170 se
rect 868 1136 1276 1170
rect 1310 1136 1348 1170
rect 1382 1136 1394 1170
tri 829 1131 834 1136 se
rect 834 1131 1394 1136
rect 829 1130 1394 1131
rect 244 1030 290 1042
rect 244 996 250 1030
rect 284 996 290 1030
rect 244 958 290 996
rect 244 924 250 958
rect 284 924 290 958
rect 244 869 290 924
tri 828 878 829 879 se
rect 829 878 875 1130
tri 875 1081 924 1130 nw
tri 978 1081 980 1083 se
rect 980 1081 1413 1083
tri 974 1077 978 1081 se
rect 978 1077 1413 1081
tri 290 869 299 878 sw
tri 819 869 828 878 se
rect 828 869 875 878
rect 244 853 299 869
tri 299 853 315 869 sw
tri 813 863 819 869 se
rect 819 863 875 869
tri 940 1043 974 1077 se
rect 974 1043 1295 1077
rect 1329 1043 1367 1077
rect 1401 1043 1413 1077
rect 940 1037 1413 1043
rect 940 1030 986 1037
rect 940 996 946 1030
rect 980 996 986 1030
tri 986 1009 1014 1037 nw
rect 940 958 986 996
rect 940 924 946 958
rect 980 924 986 958
tri 803 853 813 863 se
rect 813 853 875 863
tri 875 853 885 863 sw
rect 83 847 213 853
rect 83 813 95 847
rect 129 813 167 847
rect 201 813 213 847
rect 83 807 213 813
rect 244 847 885 853
rect 244 813 767 847
rect 801 813 839 847
rect 873 813 885 847
rect 244 807 885 813
rect 244 595 290 807
tri 290 781 316 807 nw
rect 940 705 986 924
tri 1478 876 1516 914 se
rect 1516 894 1562 1784
tri 1562 1777 1569 1784 nw
tri 1767 942 1833 1008 se
rect 1833 988 1879 2639
rect 2529 2745 2575 2757
rect 2529 2711 2535 2745
rect 2569 2711 2575 2745
rect 2529 2673 2575 2711
rect 2529 2639 2535 2673
rect 2569 2639 2575 2673
tri 2120 2529 2126 2535 se
rect 2126 2529 2481 2535
tri 2086 2495 2120 2529 se
rect 2120 2495 2363 2529
rect 2397 2495 2435 2529
rect 2469 2495 2481 2529
tri 2060 2469 2086 2495 se
rect 2086 2489 2481 2495
rect 2086 2469 2126 2489
tri 2126 2469 2146 2489 nw
tri 2042 2451 2060 2469 se
rect 2060 2451 2108 2469
tri 2108 2451 2126 2469 nw
tri 2035 1758 2042 1765 se
rect 2042 1758 2088 2451
tri 2088 2431 2108 2451 nw
tri 2463 2310 2529 2376 se
rect 2529 2356 2575 2639
tri 2529 2310 2575 2356 nw
tri 2458 2305 2463 2310 se
rect 2463 2305 2524 2310
tri 2524 2305 2529 2310 nw
tri 2196 2239 2262 2305 se
rect 2262 2259 2478 2305
tri 2478 2259 2524 2305 nw
tri 2262 2239 2282 2259 nw
tri 2028 1751 2035 1758 se
rect 2035 1751 2088 1758
tri 2023 1746 2028 1751 se
rect 2028 1746 2088 1751
tri 2016 1739 2023 1746 se
rect 2023 1739 2088 1746
rect 1959 1687 1965 1739
rect 2017 1687 2029 1739
rect 2081 1687 2088 1739
tri 2016 1680 2023 1687 ne
rect 2023 1680 2088 1687
tri 2023 1675 2028 1680 ne
rect 2028 1675 2088 1680
tri 2028 1668 2035 1675 ne
rect 2035 1668 2088 1675
tri 2035 1661 2042 1668 ne
tri 1833 942 1879 988 nw
tri 1976 950 2042 1016 se
rect 2042 996 2088 1668
tri 2042 950 2088 996 nw
tri 2154 2197 2196 2239 se
rect 2196 2197 2220 2239
tri 2220 2197 2262 2239 nw
tri 1968 942 1976 950 se
rect 1516 876 1544 894
tri 1544 876 1562 894 nw
tri 1701 876 1767 942 se
tri 1767 876 1833 942 nw
tri 1910 884 1968 942 se
rect 1968 884 1976 942
tri 1976 884 2042 950 nw
tri 1902 876 1910 884 se
rect 1910 876 1937 884
tri 1450 848 1478 876 se
rect 1478 848 1516 876
tri 1516 848 1544 876 nw
tri 1673 848 1701 876 se
rect 1701 848 1736 876
tri 1447 845 1450 848 se
rect 1450 845 1513 848
tri 1513 845 1516 848 nw
tri 1670 845 1673 848 se
rect 1673 845 1736 848
tri 1736 845 1767 876 nw
tri 1871 845 1902 876 se
rect 1902 845 1937 876
tri 1937 845 1976 884 nw
tri 1417 815 1447 845 se
rect 1447 815 1483 845
tri 1483 815 1513 845 nw
tri 1640 815 1670 845 se
rect 1670 815 1702 845
rect 1417 811 1479 815
tri 1479 811 1483 815 nw
tri 1636 811 1640 815 se
rect 1640 811 1702 815
tri 1702 811 1736 845 nw
tri 1844 818 1871 845 se
rect 1871 818 1910 845
tri 1910 818 1937 845 nw
tri 1837 811 1844 818 se
rect 1844 811 1903 818
tri 1903 811 1910 818 nw
rect 1417 810 1478 811
tri 1478 810 1479 811 nw
tri 1635 810 1636 811 se
rect 1636 810 1701 811
tri 1701 810 1702 811 nw
tri 1836 810 1837 811 se
rect 1837 810 1888 811
tri 986 705 1011 730 sw
tri 1413 705 1417 709 se
rect 1417 705 1463 810
tri 1463 795 1478 810 nw
tri 1620 795 1635 810 se
rect 1635 795 1675 810
tri 1609 784 1620 795 se
rect 1620 784 1675 795
tri 1675 784 1701 810 nw
tri 1822 796 1836 810 se
rect 1836 796 1888 810
tri 1888 796 1903 811 nw
rect 1822 784 1876 796
tri 1876 784 1888 796 nw
rect 940 693 1011 705
tri 1011 693 1023 705 sw
tri 1409 701 1413 705 se
rect 1413 701 1463 705
tri 1405 697 1409 701 se
rect 1409 697 1463 701
tri 1401 693 1405 697 se
rect 1405 693 1463 697
rect 940 685 1023 693
tri 1023 685 1031 693 sw
tri 1397 689 1401 693 se
rect 1401 689 1463 693
tri 1393 685 1397 689 se
rect 1397 685 1463 689
rect 940 639 1129 685
tri 1391 683 1393 685 se
rect 1393 683 1463 685
tri 1038 617 1060 639 ne
rect 1060 617 1129 639
rect 1333 677 1463 683
rect 1333 643 1345 677
rect 1379 643 1417 677
rect 1451 643 1463 677
rect 1333 637 1463 643
tri 1605 780 1609 784 se
rect 1609 780 1671 784
tri 1671 780 1675 784 nw
rect 1822 780 1872 784
tri 1872 780 1876 784 nw
tri 2150 780 2154 784 se
rect 2154 780 2200 2197
tri 2200 2177 2220 2197 nw
rect 2445 1803 2451 1855
rect 2503 1803 2515 1855
rect 2567 1803 2573 1855
tri 2501 1796 2508 1803 ne
rect 2508 1796 2573 1803
tri 2508 1791 2513 1796 ne
rect 2513 1791 2573 1796
tri 2513 1784 2520 1791 ne
rect 2520 1784 2573 1791
tri 2520 1777 2527 1784 ne
rect 2295 1687 2301 1739
rect 2353 1687 2365 1739
rect 2417 1687 2423 1739
tri 2351 1680 2358 1687 ne
rect 2358 1680 2423 1687
tri 2358 1675 2363 1680 ne
rect 2363 1675 2423 1680
tri 2363 1668 2370 1675 ne
rect 2370 1668 2423 1675
tri 2370 1661 2377 1668 ne
rect 1605 769 1660 780
tri 1660 769 1671 780 nw
tri 1060 601 1076 617 ne
rect 1076 601 1129 617
tri 526 599 528 601 ne
rect 528 599 530 601
tri 576 599 578 601 nw
tri 1076 599 1078 601 ne
rect 1078 599 1129 601
tri 528 597 530 599 ne
tri 1078 597 1080 599 ne
rect 1080 597 1129 599
rect 244 561 250 595
rect 284 561 290 595
tri 1080 594 1083 597 ne
rect 244 523 290 561
rect 244 489 250 523
rect 284 489 290 523
rect 244 477 290 489
rect 1083 533 1129 597
tri 1597 583 1605 591 se
rect 1605 583 1651 769
tri 1651 760 1660 769 nw
tri 1813 700 1822 709 se
rect 1822 700 1868 780
tri 1868 776 1872 780 nw
tri 2146 776 2150 780 se
rect 2150 776 2200 780
tri 2139 769 2146 776 se
rect 2146 769 2200 776
tri 2105 735 2139 769 se
rect 2139 764 2200 769
rect 2139 735 2171 764
tri 2171 735 2200 764 nw
rect 2377 845 2423 1668
rect 2527 1201 2573 1784
tri 2573 1201 2577 1205 sw
rect 2527 1185 2577 1201
tri 2527 1135 2577 1185 ne
tri 2577 1135 2643 1201 sw
tri 2577 1069 2643 1135 ne
tri 2643 1069 2709 1135 sw
tri 2643 1003 2709 1069 ne
tri 2709 1003 2775 1069 sw
tri 2709 983 2729 1003 ne
rect 2377 811 2383 845
rect 2417 811 2423 845
rect 2377 769 2423 811
rect 2377 735 2383 769
rect 2417 735 2423 769
tri 2102 732 2105 735 se
rect 2105 732 2168 735
tri 2168 732 2171 735 nw
tri 2088 718 2102 732 se
rect 2102 718 2154 732
tri 2154 718 2168 732 nw
tri 1806 693 1813 700 se
rect 1813 693 1868 700
tri 2063 693 2088 718 se
rect 2088 693 2129 718
tri 2129 693 2154 718 nw
rect 2377 693 2423 735
tri 1805 692 1806 693 se
rect 1806 692 1868 693
tri 1796 683 1805 692 se
rect 1805 683 1868 692
tri 2053 683 2063 693 se
rect 2063 683 2095 693
rect 1738 677 1868 683
rect 1738 643 1750 677
rect 1784 643 1822 677
rect 1856 643 1868 677
tri 2029 659 2053 683 se
rect 2053 659 2095 683
tri 2095 659 2129 693 nw
rect 2377 659 2383 693
rect 2417 659 2423 693
tri 2023 653 2029 659 se
rect 2029 653 2089 659
tri 2089 653 2095 659 nw
tri 2022 652 2023 653 se
rect 2023 652 2088 653
tri 2088 652 2089 653 nw
rect 1738 637 1868 643
tri 2007 637 2022 652 se
rect 2022 637 2070 652
tri 1596 582 1597 583 se
rect 1597 582 1651 583
tri 2004 634 2007 637 se
rect 2007 634 2070 637
tri 2070 634 2088 652 nw
rect 2004 617 2053 634
tri 2053 617 2070 634 nw
rect 2377 617 2423 659
tri 1587 573 1596 582 se
rect 1596 573 1651 582
tri 1995 573 2004 582 se
rect 2004 573 2050 617
tri 2050 614 2053 617 nw
tri 1559 545 1587 573 se
rect 1587 571 1651 573
rect 1587 545 1625 571
tri 1625 545 1651 571 nw
tri 1967 545 1995 573 se
rect 1995 545 2050 573
rect 1083 499 1089 533
rect 1123 499 1129 533
rect 1083 461 1129 499
tri 153 427 154 428 sw
rect 1083 427 1089 461
rect 1123 427 1129 461
rect 153 415 154 427
tri 154 415 166 427 sw
rect 1083 415 1129 427
rect 1286 541 1621 545
tri 1621 541 1625 545 nw
rect 1286 533 1613 541
tri 1613 533 1621 541 nw
rect 1868 533 2050 545
rect 1286 499 1292 533
rect 1326 499 1579 533
tri 1579 499 1613 533 nw
rect 1868 499 1874 533
rect 1908 499 2050 533
rect 1286 464 1342 499
tri 1342 464 1377 499 nw
rect 1868 471 2050 499
rect 2377 583 2383 617
rect 2417 583 2423 617
rect 2377 541 2423 583
rect 2729 845 2775 1003
rect 2729 811 2735 845
rect 2769 811 2775 845
rect 2729 766 2775 811
rect 2729 732 2735 766
rect 2769 732 2775 766
rect 2729 687 2775 732
rect 2729 653 2735 687
rect 2769 653 2775 687
rect 2729 607 2775 653
rect 2729 573 2735 607
rect 2769 573 2775 607
rect 2729 561 2775 573
rect 2377 507 2383 541
rect 2417 507 2423 541
tri 2050 471 2056 477 sw
rect 1868 465 2056 471
rect 1286 461 1339 464
tri 1339 461 1342 464 nw
rect 1868 461 2004 465
rect 1286 427 1292 461
rect 1326 427 1332 461
tri 1332 454 1339 461 nw
rect 1286 415 1332 427
rect 1868 427 1874 461
rect 1908 427 2004 461
rect 153 402 166 415
tri 166 402 179 415 sw
rect 1868 413 2004 427
rect 2377 464 2423 507
rect 2377 430 2383 464
rect 2417 430 2423 464
rect 2377 418 2423 430
rect 1868 401 2056 413
rect 1868 389 2004 401
rect 1868 355 1874 389
rect 1908 355 2004 389
rect 1868 349 2004 355
rect 1868 343 2056 349
rect 420 282 3418 294
rect 420 248 426 282
rect 460 248 536 282
rect 570 248 803 282
rect 837 248 913 282
rect 947 248 1469 282
rect 1503 248 1545 282
rect 1579 248 1621 282
rect 1655 248 1697 282
rect 1731 248 2207 282
rect 2241 248 2559 282
rect 2593 248 2911 282
rect 2945 248 3418 282
rect 420 210 3418 248
rect 420 176 426 210
rect 460 176 536 210
rect 570 176 803 210
rect 837 176 913 210
rect 947 176 1469 210
rect 1503 176 1545 210
rect 1579 176 1621 210
rect 1655 176 1697 210
rect 1731 176 2207 210
rect 2241 176 2559 210
rect 2593 176 2911 210
rect 2945 176 3418 210
rect 420 138 3418 176
rect 420 104 426 138
rect 460 104 536 138
rect 570 104 803 138
rect 837 104 913 138
rect 947 104 1469 138
rect 1503 104 1545 138
rect 1579 104 1621 138
rect 1655 104 1697 138
rect 1731 104 2207 138
rect 2241 104 2559 138
rect 2593 104 2911 138
rect 2945 104 3418 138
rect 420 66 3418 104
rect 420 32 426 66
rect 460 32 536 66
rect 570 32 803 66
rect 837 32 913 66
rect 947 32 1469 66
rect 1503 32 1545 66
rect 1579 32 1621 66
rect 1655 32 1697 66
rect 1731 32 2207 66
rect 2241 32 2559 66
rect 2593 32 2911 66
rect 2945 32 3418 66
rect 420 20 3418 32
rect 1922 -125 1928 -73
rect 1980 -125 1992 -73
rect 2044 -125 2050 -73
<< via1 >>
rect 1336 1687 1388 1739
rect 1400 1687 1452 1739
rect 1522 1803 1574 1855
rect 1586 1803 1638 1855
rect 1965 1687 2017 1739
rect 2029 1687 2081 1739
rect 2451 1803 2503 1855
rect 2515 1803 2567 1855
rect 2301 1687 2353 1739
rect 2365 1687 2417 1739
rect 2004 413 2056 465
rect 2004 349 2056 401
rect 1928 -125 1980 -73
rect 1992 -125 2044 -73
<< metal2 >>
rect 1516 1803 1522 1855
rect 1574 1803 1586 1855
rect 1638 1803 2451 1855
rect 2503 1803 2515 1855
rect 2567 1803 2573 1855
rect 1330 1687 1336 1739
rect 1388 1687 1400 1739
rect 1452 1687 1965 1739
rect 2017 1687 2029 1739
rect 2081 1687 2301 1739
rect 2353 1687 2365 1739
rect 2417 1687 2423 1739
rect 2004 465 2056 471
rect 2004 401 2056 413
rect 2004 343 2056 349
rect 2004 -73 2050 343
rect 1922 -125 1928 -73
rect 1980 -125 1992 -73
rect 2044 -125 2050 -73
use nfet_CDNS_52468879185919  nfet_CDNS_52468879185919_0
timestamp 1707688321
transform 1 0 2604 0 1 -5
box -79 -32 522 1032
use nfet_CDNS_52468879185921  nfet_CDNS_52468879185921_0
timestamp 1707688321
transform 1 0 2252 0 1 -5
box -79 -32 375 1032
use nfet_CDNS_52468879185922  nfet_CDNS_52468879185922_0
timestamp 1707688321
transform -1 0 1863 0 1 -5
box -79 -32 346 632
use nfet_CDNS_52468879185922  nfet_CDNS_52468879185922_1
timestamp 1707688321
transform 1 0 1337 0 1 -5
box -79 -32 346 632
use nfet_CDNS_52468879185928  nfet_CDNS_52468879185928_0
timestamp 1707688321
transform -1 0 1078 0 1 344
box -79 -32 346 232
use nfet_CDNS_52468879185928  nfet_CDNS_52468879185928_1
timestamp 1707688321
transform 1 0 295 0 1 344
box -79 -32 346 232
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_0
timestamp 1707688321
transform -1 0 999 0 1 2897
box -119 -66 239 150
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_1
timestamp 1707688321
transform 1 0 1055 0 1 2897
box -119 -66 239 150
use pfet_CDNS_52468879185920  pfet_CDNS_52468879185920_0
timestamp 1707688321
transform -1 0 2700 0 -1 3177
box -119 -66 562 666
use pfet_CDNS_52468879185920  pfet_CDNS_52468879185920_1
timestamp 1707688321
transform 1 0 1708 0 -1 3177
box -119 -66 562 666
use pfet_CDNS_52468879185926  pfet_CDNS_52468879185926_0
timestamp 1707688321
transform -1 0 1111 0 -1 1095
box -119 -66 562 266
use pfet_CDNS_52468879185926  pfet_CDNS_52468879185926_1
timestamp 1707688321
transform 1 0 119 0 -1 1095
box -119 -66 562 266
<< labels >>
flabel metal1 s 2183 2979 2319 3100 0 FreeSans 200 0 0 0 vswitch
port 1 nsew
flabel metal1 s 1223 123 1294 209 0 FreeSans 200 0 0 0 vssio_q
port 2 nsew
flabel metal1 s 520 1394 678 1504 0 FreeSans 200 0 0 0 vddio_q
port 3 nsew
flabel metal1 s 105 818 184 845 0 FreeSans 200 0 0 0 in_h
port 4 nsew
<< properties >>
string GDS_END 80564636
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80535304
string path 84.900 -5.425 84.900 31.200 41.000 31.200 
<< end >>
