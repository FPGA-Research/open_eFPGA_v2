magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 0 1022 3324
<< mvnsubdiff >>
rect 66 3224 90 3258
rect 124 3224 164 3258
rect 198 3224 237 3258
rect 271 3224 310 3258
rect 344 3224 383 3258
rect 417 3224 597 3258
rect 631 3224 667 3258
rect 701 3224 736 3258
rect 770 3224 805 3258
rect 839 3224 956 3258
rect 66 3164 100 3224
rect 66 3095 100 3130
rect 66 3026 100 3061
rect 66 2957 100 2992
rect 66 2888 100 2923
rect 66 2819 100 2854
rect 66 2750 100 2785
rect 66 2681 100 2716
rect 66 2612 100 2647
rect 66 2543 100 2578
rect 66 2474 100 2509
rect 66 2405 100 2440
rect 66 2336 100 2371
rect 66 2267 100 2302
rect 66 2198 100 2233
rect 66 2129 100 2164
rect 66 2060 100 2095
rect 66 1991 100 2026
rect 66 1922 100 1957
rect 66 1853 100 1888
rect 66 1784 100 1819
rect 66 1715 100 1750
rect 66 1646 100 1681
rect 66 1577 100 1612
rect 66 1508 100 1543
rect 66 1439 100 1474
rect 66 1370 100 1405
rect 66 1301 100 1336
rect 66 1232 100 1267
rect 66 1163 100 1198
rect 66 1094 100 1129
rect 66 1025 100 1060
rect 66 956 100 991
rect 66 887 100 922
rect 66 818 100 853
rect 66 749 100 784
rect 66 680 100 715
rect 66 611 100 646
rect 66 542 100 577
rect 66 473 100 508
rect 66 404 100 439
rect 66 334 100 370
rect 66 264 100 300
rect 66 194 100 230
rect 66 124 100 160
rect 922 100 956 3224
rect 100 90 168 100
rect 66 66 168 90
rect 202 66 241 100
rect 275 66 314 100
rect 348 66 387 100
rect 421 66 461 100
rect 495 66 535 100
rect 569 66 609 100
rect 643 66 683 100
rect 717 66 757 100
rect 791 66 831 100
rect 865 66 956 100
<< mvnsubdiffcont >>
rect 90 3224 124 3258
rect 164 3224 198 3258
rect 237 3224 271 3258
rect 310 3224 344 3258
rect 383 3224 417 3258
rect 597 3224 631 3258
rect 667 3224 701 3258
rect 736 3224 770 3258
rect 805 3224 839 3258
rect 66 3130 100 3164
rect 66 3061 100 3095
rect 66 2992 100 3026
rect 66 2923 100 2957
rect 66 2854 100 2888
rect 66 2785 100 2819
rect 66 2716 100 2750
rect 66 2647 100 2681
rect 66 2578 100 2612
rect 66 2509 100 2543
rect 66 2440 100 2474
rect 66 2371 100 2405
rect 66 2302 100 2336
rect 66 2233 100 2267
rect 66 2164 100 2198
rect 66 2095 100 2129
rect 66 2026 100 2060
rect 66 1957 100 1991
rect 66 1888 100 1922
rect 66 1819 100 1853
rect 66 1750 100 1784
rect 66 1681 100 1715
rect 66 1612 100 1646
rect 66 1543 100 1577
rect 66 1474 100 1508
rect 66 1405 100 1439
rect 66 1336 100 1370
rect 66 1267 100 1301
rect 66 1198 100 1232
rect 66 1129 100 1163
rect 66 1060 100 1094
rect 66 991 100 1025
rect 66 922 100 956
rect 66 853 100 887
rect 66 784 100 818
rect 66 715 100 749
rect 66 646 100 680
rect 66 577 100 611
rect 66 508 100 542
rect 66 439 100 473
rect 66 370 100 404
rect 66 300 100 334
rect 66 230 100 264
rect 66 160 100 194
rect 66 90 100 124
rect 168 66 202 100
rect 241 66 275 100
rect 314 66 348 100
rect 387 66 421 100
rect 461 66 495 100
rect 535 66 569 100
rect 609 66 643 100
rect 683 66 717 100
rect 757 66 791 100
rect 831 66 865 100
<< poly >>
rect 227 1646 327 1724
rect 383 1646 483 1724
rect 539 1646 639 1724
rect 695 1646 795 1724
rect 227 122 327 194
rect 383 122 483 194
rect 539 122 639 194
rect 695 122 795 194
<< locali >>
rect 66 3224 90 3258
rect 124 3224 164 3258
rect 198 3224 237 3258
rect 271 3224 310 3258
rect 344 3224 383 3258
rect 417 3224 597 3258
rect 631 3224 667 3258
rect 701 3224 736 3258
rect 770 3224 805 3258
rect 839 3224 956 3258
rect 66 3164 100 3224
rect 66 3095 100 3130
rect 66 3026 100 3061
rect 66 2957 100 2992
rect 66 2888 100 2923
rect 66 2819 100 2854
rect 66 2750 100 2785
rect 66 2681 100 2716
rect 66 2612 100 2647
rect 66 2543 100 2578
rect 66 2474 100 2509
rect 66 2405 100 2440
rect 66 2336 100 2371
rect 66 2267 100 2302
rect 66 2198 100 2233
rect 66 2129 100 2164
rect 66 2060 100 2095
rect 66 1991 100 2026
rect 66 1922 100 1957
rect 182 2982 216 3021
rect 182 2909 216 2948
rect 494 2982 528 3021
rect 494 2909 528 2948
rect 182 2836 216 2875
rect 182 2763 216 2802
rect 182 2690 216 2729
rect 182 2617 216 2656
rect 182 2545 216 2583
rect 182 2473 216 2511
rect 182 2401 216 2439
rect 182 2329 216 2367
rect 182 2257 216 2295
rect 182 2185 216 2223
rect 182 2113 216 2151
rect 182 2041 216 2079
rect 182 1969 216 2007
rect 338 2818 372 2857
rect 338 2745 372 2784
rect 338 2672 372 2711
rect 338 2599 372 2638
rect 338 2526 372 2565
rect 338 2453 372 2492
rect 338 2380 372 2419
rect 338 2307 372 2346
rect 338 2234 372 2273
rect 338 2161 372 2200
rect 338 2089 372 2127
rect 338 2017 372 2055
rect 338 1945 372 1983
rect 66 1853 100 1888
rect 66 1784 100 1819
rect 806 3039 840 3082
rect 806 2962 840 3005
rect 494 2836 528 2875
rect 494 2763 528 2802
rect 494 2690 528 2729
rect 494 2617 528 2656
rect 494 2545 528 2583
rect 494 2473 528 2511
rect 494 2401 528 2439
rect 494 2329 528 2367
rect 494 2257 528 2295
rect 494 2185 528 2223
rect 494 2113 528 2151
rect 494 2041 528 2079
rect 494 1969 528 2007
rect 650 2818 684 2857
rect 650 2745 684 2784
rect 650 2672 684 2711
rect 650 2599 684 2638
rect 650 2526 684 2565
rect 650 2453 684 2492
rect 650 2380 684 2419
rect 650 2307 684 2346
rect 650 2234 684 2273
rect 650 2161 684 2200
rect 650 2089 684 2127
rect 650 2017 684 2055
rect 650 1945 684 1983
rect 338 1873 372 1911
rect 338 1801 372 1839
rect 806 2885 840 2928
rect 806 2808 840 2851
rect 806 2731 840 2774
rect 806 2654 840 2697
rect 806 2577 840 2620
rect 806 2501 840 2543
rect 806 2425 840 2467
rect 806 2349 840 2391
rect 806 2273 840 2315
rect 806 2197 840 2239
rect 806 2121 840 2163
rect 806 2045 840 2087
rect 806 1969 840 2011
rect 650 1873 684 1911
rect 650 1801 684 1839
rect 66 1715 100 1750
rect 66 1646 100 1681
rect 240 1650 782 1702
rect 240 1616 251 1650
rect 285 1616 334 1650
rect 368 1616 417 1650
rect 451 1616 500 1650
rect 534 1616 583 1650
rect 617 1616 666 1650
rect 700 1616 748 1650
rect 66 1577 100 1612
rect 66 1508 100 1543
rect 66 1439 100 1474
rect 66 1370 100 1405
rect 66 1301 100 1336
rect 66 1232 100 1267
rect 66 1163 100 1198
rect 66 1094 100 1129
rect 66 1025 100 1060
rect 66 956 100 991
rect 66 887 100 922
rect 66 818 100 853
rect 66 749 100 784
rect 66 680 100 715
rect 66 611 100 646
rect 66 542 100 577
rect 66 473 100 508
rect 66 404 100 439
rect 66 334 100 370
rect 66 264 100 300
rect 182 1303 216 1341
rect 182 1231 216 1269
rect 182 1159 216 1197
rect 182 1087 216 1125
rect 182 1015 216 1053
rect 182 943 216 981
rect 182 871 216 909
rect 182 799 216 837
rect 182 727 216 765
rect 182 654 216 693
rect 182 581 216 620
rect 182 508 216 547
rect 182 435 216 474
rect 182 362 216 401
rect 182 289 216 328
rect 66 194 100 230
rect 66 124 100 160
rect 250 138 304 1616
rect 338 1497 372 1536
rect 338 1424 372 1463
rect 338 1351 372 1390
rect 338 1278 372 1317
rect 338 1206 372 1244
rect 338 1134 372 1172
rect 338 1062 372 1100
rect 338 990 372 1028
rect 338 918 372 956
rect 338 846 372 884
rect 338 774 372 812
rect 338 702 372 740
rect 338 630 372 668
rect 338 558 372 596
rect 338 486 372 524
rect 406 138 460 1616
rect 494 1303 528 1341
rect 494 1231 528 1269
rect 494 1159 528 1197
rect 494 1087 528 1125
rect 494 1015 528 1053
rect 494 943 528 981
rect 494 871 528 909
rect 494 799 528 837
rect 494 727 528 765
rect 494 654 528 693
rect 494 581 528 620
rect 494 508 528 547
rect 494 435 528 474
rect 494 362 528 401
rect 494 289 528 328
rect 562 138 616 1616
rect 650 1497 684 1536
rect 650 1424 684 1463
rect 650 1351 684 1390
rect 650 1278 684 1317
rect 650 1206 684 1244
rect 650 1134 684 1172
rect 650 1062 684 1100
rect 650 990 684 1028
rect 650 918 684 956
rect 650 846 684 884
rect 650 774 684 812
rect 650 702 684 740
rect 650 630 684 668
rect 650 558 684 596
rect 650 486 684 524
rect 718 138 772 1616
rect 806 1303 840 1341
rect 806 1231 840 1269
rect 806 1159 840 1197
rect 806 1087 840 1125
rect 806 1015 840 1053
rect 806 943 840 981
rect 806 871 840 909
rect 806 799 840 837
rect 806 727 840 765
rect 806 654 840 693
rect 806 581 840 620
rect 806 508 840 547
rect 806 435 840 474
rect 806 362 840 401
rect 806 289 840 328
rect 922 100 956 3224
rect 100 90 168 100
rect 66 66 168 90
rect 202 66 241 100
rect 275 66 314 100
rect 348 66 387 100
rect 421 66 461 100
rect 495 66 535 100
rect 569 66 609 100
rect 643 66 683 100
rect 717 66 757 100
rect 791 66 831 100
rect 865 66 956 100
<< viali >>
rect 806 3082 840 3116
rect 182 3021 216 3055
rect 182 2948 216 2982
rect 182 2875 216 2909
rect 494 3021 528 3055
rect 494 2948 528 2982
rect 182 2802 216 2836
rect 182 2729 216 2763
rect 182 2656 216 2690
rect 182 2583 216 2617
rect 182 2511 216 2545
rect 182 2439 216 2473
rect 182 2367 216 2401
rect 182 2295 216 2329
rect 182 2223 216 2257
rect 182 2151 216 2185
rect 182 2079 216 2113
rect 182 2007 216 2041
rect 182 1935 216 1969
rect 338 2857 372 2891
rect 338 2784 372 2818
rect 338 2711 372 2745
rect 338 2638 372 2672
rect 338 2565 372 2599
rect 338 2492 372 2526
rect 338 2419 372 2453
rect 338 2346 372 2380
rect 338 2273 372 2307
rect 338 2200 372 2234
rect 338 2127 372 2161
rect 338 2055 372 2089
rect 338 1983 372 2017
rect 338 1911 372 1945
rect 494 2875 528 2909
rect 806 3005 840 3039
rect 806 2928 840 2962
rect 494 2802 528 2836
rect 494 2729 528 2763
rect 494 2656 528 2690
rect 494 2583 528 2617
rect 494 2511 528 2545
rect 494 2439 528 2473
rect 494 2367 528 2401
rect 494 2295 528 2329
rect 494 2223 528 2257
rect 494 2151 528 2185
rect 494 2079 528 2113
rect 494 2007 528 2041
rect 494 1935 528 1969
rect 650 2857 684 2891
rect 650 2784 684 2818
rect 650 2711 684 2745
rect 650 2638 684 2672
rect 650 2565 684 2599
rect 650 2492 684 2526
rect 650 2419 684 2453
rect 650 2346 684 2380
rect 650 2273 684 2307
rect 650 2200 684 2234
rect 650 2127 684 2161
rect 650 2055 684 2089
rect 650 1983 684 2017
rect 338 1839 372 1873
rect 338 1767 372 1801
rect 650 1911 684 1945
rect 806 2851 840 2885
rect 806 2774 840 2808
rect 806 2697 840 2731
rect 806 2620 840 2654
rect 806 2543 840 2577
rect 806 2467 840 2501
rect 806 2391 840 2425
rect 806 2315 840 2349
rect 806 2239 840 2273
rect 806 2163 840 2197
rect 806 2087 840 2121
rect 806 2011 840 2045
rect 806 1935 840 1969
rect 650 1839 684 1873
rect 650 1767 684 1801
rect 251 1616 285 1650
rect 334 1616 368 1650
rect 417 1616 451 1650
rect 500 1616 534 1650
rect 583 1616 617 1650
rect 666 1616 700 1650
rect 748 1616 782 1650
rect 182 1341 216 1375
rect 182 1269 216 1303
rect 182 1197 216 1231
rect 182 1125 216 1159
rect 182 1053 216 1087
rect 182 981 216 1015
rect 182 909 216 943
rect 182 837 216 871
rect 182 765 216 799
rect 182 693 216 727
rect 182 620 216 654
rect 182 547 216 581
rect 182 474 216 508
rect 182 401 216 435
rect 182 328 216 362
rect 182 255 216 289
rect 338 1536 372 1570
rect 338 1463 372 1497
rect 338 1390 372 1424
rect 338 1317 372 1351
rect 338 1244 372 1278
rect 338 1172 372 1206
rect 338 1100 372 1134
rect 338 1028 372 1062
rect 338 956 372 990
rect 338 884 372 918
rect 338 812 372 846
rect 338 740 372 774
rect 338 668 372 702
rect 338 596 372 630
rect 338 524 372 558
rect 338 452 372 486
rect 494 1341 528 1375
rect 494 1269 528 1303
rect 494 1197 528 1231
rect 494 1125 528 1159
rect 494 1053 528 1087
rect 494 981 528 1015
rect 494 909 528 943
rect 494 837 528 871
rect 494 765 528 799
rect 494 693 528 727
rect 494 620 528 654
rect 494 547 528 581
rect 494 474 528 508
rect 494 401 528 435
rect 494 328 528 362
rect 494 255 528 289
rect 650 1536 684 1570
rect 650 1463 684 1497
rect 650 1390 684 1424
rect 650 1317 684 1351
rect 650 1244 684 1278
rect 650 1172 684 1206
rect 650 1100 684 1134
rect 650 1028 684 1062
rect 650 956 684 990
rect 650 884 684 918
rect 650 812 684 846
rect 650 740 684 774
rect 650 668 684 702
rect 650 596 684 630
rect 650 524 684 558
rect 650 452 684 486
rect 806 1341 840 1375
rect 806 1269 840 1303
rect 806 1197 840 1231
rect 806 1125 840 1159
rect 806 1053 840 1087
rect 806 981 840 1015
rect 806 909 840 943
rect 806 837 840 871
rect 806 765 840 799
rect 806 693 840 727
rect 806 620 840 654
rect 806 547 840 581
rect 806 474 840 508
rect 806 401 840 435
rect 806 328 840 362
rect 806 255 840 289
<< metal1 >>
rect 176 3116 846 3128
rect 176 3082 806 3116
rect 840 3082 846 3116
rect 176 3055 846 3082
rect 176 3021 182 3055
rect 216 3021 494 3055
rect 528 3039 846 3055
rect 528 3021 806 3039
rect 176 3005 806 3021
rect 840 3005 846 3039
rect 176 2982 846 3005
rect 176 2948 182 2982
rect 216 2959 494 2982
rect 216 2948 236 2959
tri 236 2948 247 2959 nw
tri 463 2948 474 2959 ne
rect 474 2948 494 2959
rect 528 2962 846 2982
rect 528 2959 806 2962
rect 528 2948 534 2959
rect 176 2909 222 2948
tri 222 2934 236 2948 nw
tri 474 2934 488 2948 ne
rect 176 2875 182 2909
rect 216 2875 222 2909
rect 488 2909 534 2948
tri 534 2934 559 2959 nw
tri 775 2934 800 2959 ne
rect 176 2836 222 2875
rect 176 2802 182 2836
rect 216 2802 222 2836
rect 176 2763 222 2802
rect 176 2729 182 2763
rect 216 2729 222 2763
rect 176 2690 222 2729
rect 176 2656 182 2690
rect 216 2656 222 2690
rect 176 2617 222 2656
rect 176 2583 182 2617
rect 216 2583 222 2617
rect 176 2545 222 2583
rect 176 2511 182 2545
rect 216 2511 222 2545
rect 176 2473 222 2511
rect 176 2439 182 2473
rect 216 2439 222 2473
rect 176 2401 222 2439
rect 176 2367 182 2401
rect 216 2367 222 2401
rect 176 2329 222 2367
rect 176 2295 182 2329
rect 216 2295 222 2329
rect 176 2257 222 2295
rect 176 2223 182 2257
rect 216 2223 222 2257
rect 176 2185 222 2223
rect 176 2151 182 2185
rect 216 2151 222 2185
rect 176 2113 222 2151
rect 176 2079 182 2113
rect 216 2079 222 2113
rect 176 2041 222 2079
rect 176 2007 182 2041
rect 216 2007 222 2041
rect 176 1969 222 2007
rect 176 1935 182 1969
rect 216 1935 222 1969
rect 176 1923 222 1935
rect 332 2891 378 2903
rect 332 2857 338 2891
rect 372 2857 378 2891
rect 332 2818 378 2857
rect 332 2784 338 2818
rect 372 2784 378 2818
rect 332 2745 378 2784
rect 332 2711 338 2745
rect 372 2711 378 2745
rect 332 2672 378 2711
rect 332 2638 338 2672
rect 372 2638 378 2672
rect 332 2599 378 2638
rect 332 2565 338 2599
rect 372 2565 378 2599
rect 332 2526 378 2565
rect 332 2492 338 2526
rect 372 2492 378 2526
rect 332 2453 378 2492
rect 332 2419 338 2453
rect 372 2419 378 2453
rect 332 2380 378 2419
rect 332 2346 338 2380
rect 372 2346 378 2380
rect 332 2307 378 2346
rect 332 2273 338 2307
rect 372 2273 378 2307
rect 332 2234 378 2273
rect 332 2200 338 2234
rect 372 2200 378 2234
rect 332 2161 378 2200
rect 332 2127 338 2161
rect 372 2127 378 2161
rect 332 2089 378 2127
rect 332 2055 338 2089
rect 372 2055 378 2089
rect 332 2017 378 2055
rect 332 1983 338 2017
rect 372 1983 378 2017
rect 332 1945 378 1983
rect 332 1911 338 1945
rect 372 1911 378 1945
rect 488 2875 494 2909
rect 528 2875 534 2909
rect 800 2928 806 2959
rect 840 2928 846 2962
rect 488 2836 534 2875
rect 488 2802 494 2836
rect 528 2802 534 2836
rect 488 2763 534 2802
rect 488 2729 494 2763
rect 528 2729 534 2763
rect 488 2690 534 2729
rect 488 2656 494 2690
rect 528 2656 534 2690
rect 488 2617 534 2656
rect 488 2583 494 2617
rect 528 2583 534 2617
rect 488 2545 534 2583
rect 488 2511 494 2545
rect 528 2511 534 2545
rect 488 2473 534 2511
rect 488 2439 494 2473
rect 528 2439 534 2473
rect 488 2401 534 2439
rect 488 2367 494 2401
rect 528 2367 534 2401
rect 488 2329 534 2367
rect 488 2295 494 2329
rect 528 2295 534 2329
rect 488 2257 534 2295
rect 488 2223 494 2257
rect 528 2223 534 2257
rect 488 2185 534 2223
rect 488 2151 494 2185
rect 528 2151 534 2185
rect 488 2113 534 2151
rect 488 2079 494 2113
rect 528 2079 534 2113
rect 488 2041 534 2079
rect 488 2007 494 2041
rect 528 2007 534 2041
rect 488 1969 534 2007
rect 488 1935 494 1969
rect 528 1935 534 1969
rect 488 1923 534 1935
rect 644 2891 690 2903
rect 644 2857 650 2891
rect 684 2857 690 2891
rect 644 2818 690 2857
rect 644 2784 650 2818
rect 684 2784 690 2818
rect 644 2745 690 2784
rect 644 2711 650 2745
rect 684 2711 690 2745
rect 644 2672 690 2711
rect 644 2638 650 2672
rect 684 2638 690 2672
rect 644 2599 690 2638
rect 644 2565 650 2599
rect 684 2565 690 2599
rect 644 2526 690 2565
rect 644 2492 650 2526
rect 684 2492 690 2526
rect 644 2453 690 2492
rect 644 2419 650 2453
rect 684 2419 690 2453
rect 644 2380 690 2419
rect 644 2346 650 2380
rect 684 2346 690 2380
rect 644 2307 690 2346
rect 644 2273 650 2307
rect 684 2273 690 2307
rect 644 2234 690 2273
rect 644 2200 650 2234
rect 684 2200 690 2234
rect 644 2161 690 2200
rect 644 2127 650 2161
rect 684 2127 690 2161
rect 644 2089 690 2127
rect 644 2055 650 2089
rect 684 2055 690 2089
rect 644 2017 690 2055
rect 644 1983 650 2017
rect 684 1983 690 2017
rect 644 1945 690 1983
tri 307 1885 332 1910 se
rect 332 1885 378 1911
rect 644 1911 650 1945
rect 684 1911 690 1945
rect 800 2885 846 2928
rect 800 2851 806 2885
rect 840 2851 846 2885
rect 800 2808 846 2851
rect 800 2774 806 2808
rect 840 2774 846 2808
rect 800 2731 846 2774
rect 800 2697 806 2731
rect 840 2697 846 2731
rect 800 2654 846 2697
rect 800 2620 806 2654
rect 840 2620 846 2654
rect 800 2577 846 2620
rect 800 2543 806 2577
rect 840 2543 846 2577
rect 800 2501 846 2543
rect 800 2467 806 2501
rect 840 2467 846 2501
rect 800 2425 846 2467
rect 800 2391 806 2425
rect 840 2391 846 2425
rect 800 2349 846 2391
rect 800 2315 806 2349
rect 840 2315 846 2349
rect 800 2273 846 2315
rect 800 2239 806 2273
rect 840 2239 846 2273
rect 800 2197 846 2239
rect 800 2163 806 2197
rect 840 2163 846 2197
rect 800 2121 846 2163
rect 800 2087 806 2121
rect 840 2087 846 2121
rect 800 2045 846 2087
rect 800 2011 806 2045
rect 840 2011 846 2045
rect 800 1969 846 2011
rect 800 1935 806 1969
rect 840 1935 846 1969
rect 800 1923 846 1935
tri 378 1885 403 1910 sw
tri 619 1885 644 1910 se
rect 644 1885 690 1911
rect 147 1873 690 1885
rect 147 1839 338 1873
rect 372 1839 650 1873
rect 684 1839 690 1873
rect 147 1801 690 1839
rect 147 1767 338 1801
rect 372 1767 650 1801
rect 684 1767 690 1801
rect 147 1755 690 1767
rect 147 1582 202 1755
tri 202 1730 227 1755 nw
rect 239 1650 794 1656
rect 239 1616 251 1650
rect 285 1616 334 1650
rect 368 1616 417 1650
rect 451 1616 500 1650
rect 534 1616 583 1650
rect 617 1616 666 1650
rect 700 1616 748 1650
rect 782 1616 794 1650
rect 239 1610 794 1616
tri 202 1582 227 1607 sw
rect 147 1570 690 1582
rect 147 1536 338 1570
rect 372 1536 650 1570
rect 684 1536 690 1570
rect 147 1497 690 1536
rect 147 1463 338 1497
rect 372 1463 650 1497
rect 684 1463 690 1497
rect 147 1452 690 1463
tri 307 1427 332 1452 ne
rect 332 1424 378 1452
tri 378 1427 403 1452 nw
tri 619 1427 644 1452 ne
rect 332 1390 338 1424
rect 372 1390 378 1424
rect 176 1375 222 1387
rect 176 1341 182 1375
rect 216 1341 222 1375
rect 176 1303 222 1341
rect 176 1269 182 1303
rect 216 1269 222 1303
rect 176 1231 222 1269
rect 176 1197 182 1231
rect 216 1197 222 1231
rect 176 1159 222 1197
rect 176 1125 182 1159
rect 216 1125 222 1159
rect 176 1087 222 1125
rect 176 1053 182 1087
rect 216 1053 222 1087
rect 176 1015 222 1053
rect 176 981 182 1015
rect 216 981 222 1015
rect 176 943 222 981
rect 176 909 182 943
rect 216 909 222 943
rect 176 871 222 909
rect 176 837 182 871
rect 216 837 222 871
rect 176 799 222 837
rect 176 765 182 799
rect 216 765 222 799
rect 176 727 222 765
rect 176 693 182 727
rect 216 693 222 727
rect 176 654 222 693
rect 176 620 182 654
rect 216 620 222 654
rect 176 581 222 620
rect 176 547 182 581
rect 216 547 222 581
rect 176 508 222 547
rect 176 474 182 508
rect 216 474 222 508
rect 176 435 222 474
rect 332 1351 378 1390
rect 644 1424 690 1452
rect 644 1390 650 1424
rect 684 1390 690 1424
rect 332 1317 338 1351
rect 372 1317 378 1351
rect 332 1278 378 1317
rect 332 1244 338 1278
rect 372 1244 378 1278
rect 332 1206 378 1244
rect 332 1172 338 1206
rect 372 1172 378 1206
rect 332 1134 378 1172
rect 332 1100 338 1134
rect 372 1100 378 1134
rect 332 1062 378 1100
rect 332 1028 338 1062
rect 372 1028 378 1062
rect 332 990 378 1028
rect 332 956 338 990
rect 372 956 378 990
rect 332 918 378 956
rect 332 884 338 918
rect 372 884 378 918
rect 332 846 378 884
rect 332 812 338 846
rect 372 812 378 846
rect 332 774 378 812
rect 332 740 338 774
rect 372 740 378 774
rect 332 702 378 740
rect 332 668 338 702
rect 372 668 378 702
rect 332 630 378 668
rect 332 596 338 630
rect 372 596 378 630
rect 332 558 378 596
rect 332 524 338 558
rect 372 524 378 558
rect 332 486 378 524
rect 332 452 338 486
rect 372 452 378 486
rect 332 440 378 452
rect 488 1375 534 1387
rect 488 1341 494 1375
rect 528 1341 534 1375
rect 488 1303 534 1341
rect 488 1269 494 1303
rect 528 1269 534 1303
rect 488 1231 534 1269
rect 488 1197 494 1231
rect 528 1197 534 1231
rect 488 1159 534 1197
rect 488 1125 494 1159
rect 528 1125 534 1159
rect 488 1087 534 1125
rect 488 1053 494 1087
rect 528 1053 534 1087
rect 488 1015 534 1053
rect 488 981 494 1015
rect 528 981 534 1015
rect 488 943 534 981
rect 488 909 494 943
rect 528 909 534 943
rect 488 871 534 909
rect 488 837 494 871
rect 528 837 534 871
rect 488 799 534 837
rect 488 765 494 799
rect 528 765 534 799
rect 488 727 534 765
rect 488 693 494 727
rect 528 693 534 727
rect 488 654 534 693
rect 488 620 494 654
rect 528 620 534 654
rect 488 581 534 620
rect 488 547 494 581
rect 528 547 534 581
rect 488 508 534 547
rect 488 474 494 508
rect 528 474 534 508
tri 222 435 224 437 sw
tri 486 435 488 437 se
rect 488 435 534 474
rect 644 1351 690 1390
rect 644 1317 650 1351
rect 684 1317 690 1351
rect 644 1278 690 1317
rect 644 1244 650 1278
rect 684 1244 690 1278
rect 644 1206 690 1244
rect 644 1172 650 1206
rect 684 1172 690 1206
rect 644 1134 690 1172
rect 644 1100 650 1134
rect 684 1100 690 1134
rect 644 1062 690 1100
rect 644 1028 650 1062
rect 684 1028 690 1062
rect 644 990 690 1028
rect 644 956 650 990
rect 684 956 690 990
rect 644 918 690 956
rect 644 884 650 918
rect 684 884 690 918
rect 644 846 690 884
rect 644 812 650 846
rect 684 812 690 846
rect 644 774 690 812
rect 644 740 650 774
rect 684 740 690 774
rect 644 702 690 740
rect 644 668 650 702
rect 684 668 690 702
rect 644 630 690 668
rect 644 596 650 630
rect 684 596 690 630
rect 644 558 690 596
rect 644 524 650 558
rect 684 524 690 558
rect 644 486 690 524
rect 644 452 650 486
rect 684 452 690 486
rect 644 440 690 452
rect 800 1375 846 1387
rect 800 1341 806 1375
rect 840 1341 846 1375
rect 800 1303 846 1341
rect 800 1269 806 1303
rect 840 1269 846 1303
rect 800 1231 846 1269
rect 800 1197 806 1231
rect 840 1197 846 1231
rect 800 1159 846 1197
rect 800 1125 806 1159
rect 840 1125 846 1159
rect 800 1087 846 1125
rect 800 1053 806 1087
rect 840 1053 846 1087
rect 800 1015 846 1053
rect 800 981 806 1015
rect 840 981 846 1015
rect 800 943 846 981
rect 800 909 806 943
rect 840 909 846 943
rect 800 871 846 909
rect 800 837 806 871
rect 840 837 846 871
rect 800 799 846 837
rect 800 765 806 799
rect 840 765 846 799
rect 800 727 846 765
rect 800 693 806 727
rect 840 693 846 727
rect 800 654 846 693
rect 800 620 806 654
rect 840 620 846 654
rect 800 581 846 620
rect 800 547 806 581
rect 840 547 846 581
rect 800 508 846 547
rect 800 474 806 508
rect 840 474 846 508
tri 534 435 536 437 sw
tri 798 435 800 437 se
rect 800 435 846 474
rect 176 401 182 435
rect 216 412 224 435
tri 224 412 247 435 sw
tri 463 412 486 435 se
rect 486 412 494 435
rect 216 401 494 412
rect 528 412 536 435
tri 536 412 559 435 sw
tri 775 412 798 435 se
rect 798 412 806 435
rect 528 401 806 412
rect 840 401 846 435
rect 176 362 846 401
rect 176 328 182 362
rect 216 328 494 362
rect 528 328 806 362
rect 840 328 846 362
rect 176 289 846 328
rect 176 255 182 289
rect 216 255 494 289
rect 528 255 806 289
rect 840 255 846 289
rect 176 243 846 255
use pfet_CDNS_524688791851506  pfet_CDNS_524688791851506_0
timestamp 1707688321
transform 1 0 227 0 1 220
box -119 -66 687 1466
use pfet_CDNS_524688791851506  pfet_CDNS_524688791851506_1
timestamp 1707688321
transform 1 0 227 0 1 1750
box -119 -66 687 1466
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 1 240 1 0 1652
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1707688321
transform 0 1 240 1 0 122
box 0 0 66 542
<< labels >>
flabel comment s 455 1756 455 1756 0 FreeSans 4000 90 0 0 vpb_drvr
flabel metal1 s 348 3006 641 3078 0 FreeSans 200 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 368 275 626 363 0 FreeSans 200 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 298 1489 558 1541 0 FreeSans 200 0 0 0 pad
port 2 nsew
<< properties >>
string GDS_END 90856168
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90837526
string path 13.675 81.025 23.475 81.025 23.475 2.075 2.075 2.075 2.075 81.025 11.675 81.025 
<< end >>
