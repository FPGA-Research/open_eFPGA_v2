magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 9073 31184 9199 33647
rect 9743 27456 14485 34842
rect 9743 26324 12512 27456
rect 173 16896 2252 17326
rect 173 9911 4863 16896
rect 173 385 6231 9911
rect 4863 190 6231 385
<< nwell >>
rect 9663 34636 14565 34922
rect 9663 33647 9949 34636
rect 8993 31184 9279 33647
rect 9855 33581 9949 33647
rect 9663 26530 9949 31310
rect 14279 27662 14565 34636
rect 12306 27376 14565 27662
rect 12306 26530 12592 27376
rect 9663 26244 12592 26530
rect 63 16976 2337 17411
rect 63 16951 370 16976
rect 744 16951 4973 16976
rect 63 16806 4973 16951
rect 63 12216 233 16806
rect 2433 12216 2603 16806
rect 4803 12216 4973 16806
rect 63 12046 4973 12216
rect 63 9801 575 12046
rect 2433 9801 2603 12046
rect 4461 9991 4973 12046
rect 4461 9801 6311 9991
rect 63 9631 6311 9801
rect 63 470 453 9631
rect 5951 470 6311 9631
rect 63 300 6311 470
rect 4583 110 6311 300
<< pwell >>
rect 10014 34486 14219 34572
rect 10014 32320 10100 34486
rect 14133 32320 14219 34486
rect 10014 32234 14219 32320
rect 10014 30069 10100 32234
rect 14133 30069 14219 32234
rect 10014 29983 14219 30069
rect 10014 27815 10100 29983
rect 14133 27815 14219 29983
rect 10014 27729 14219 27815
rect 635 9861 723 11986
rect 2285 9861 2373 11986
rect 2663 9861 2751 11986
rect 4313 9861 4401 11986
rect 5033 15752 5710 15840
rect 5033 15000 5121 15752
rect 5622 15000 5710 15752
rect 5033 14885 5710 15000
rect 5033 14655 6365 14885
rect 5033 13788 5555 14655
rect 5033 10281 5121 13788
rect 6277 10281 6365 14655
rect 5033 10051 6365 10281
rect 513 9483 5891 9571
rect 513 7314 601 9483
rect 3330 7314 3418 9483
rect 5803 7314 5891 9483
rect 513 7226 993 7314
rect 1211 7226 1849 7314
rect 2067 7226 2705 7314
rect 2923 7226 3825 7314
rect 4043 7226 4481 7314
rect 4699 7226 4937 7314
rect 5155 7226 5393 7314
rect 5611 7226 5891 7314
rect 513 5094 601 7226
rect 3330 5094 3418 7226
rect 5803 5094 5891 7226
rect 513 5006 993 5094
rect 1211 5006 1849 5094
rect 2067 5006 2705 5094
rect 2923 5006 3825 5094
rect 4043 5006 4481 5094
rect 4699 5006 4937 5094
rect 5155 5006 5393 5094
rect 5611 5006 5891 5094
rect 513 2875 601 5006
rect 3330 2875 3418 5006
rect 5803 2875 5891 5006
rect 513 2787 993 2875
rect 1211 2787 1849 2875
rect 2067 2787 2705 2875
rect 2923 2787 3825 2875
rect 4043 2787 4481 2875
rect 4699 2787 4937 2875
rect 5155 2787 5393 2875
rect 5611 2787 5891 2875
rect 513 618 601 2787
rect 3330 618 3418 2787
rect 5803 618 5891 2787
rect 513 530 5891 618
<< mvndiff >>
rect 5169 14741 5249 14749
rect 5169 14707 5192 14741
rect 5226 14707 5249 14741
rect 5169 14681 5249 14707
rect 5309 13874 5389 14749
rect 5309 13840 5332 13874
rect 5366 13840 5389 13874
rect 5309 13814 5389 13840
rect 5449 13874 5529 14749
rect 5589 14741 5669 14749
rect 5589 14707 5612 14741
rect 5646 14707 5669 14741
rect 5589 14681 5669 14707
rect 5729 14741 5809 14749
rect 5729 14707 5752 14741
rect 5786 14707 5809 14741
rect 5729 14681 5809 14707
rect 5869 14741 5949 14749
rect 5869 14707 5892 14741
rect 5926 14707 5949 14741
rect 5869 14681 5949 14707
rect 6009 14741 6089 14749
rect 6009 14707 6032 14741
rect 6066 14707 6089 14741
rect 6009 14681 6089 14707
rect 6149 14741 6229 14749
rect 6149 14707 6172 14741
rect 6206 14707 6229 14741
rect 6149 14681 6229 14707
rect 5449 13840 5472 13874
rect 5506 13840 5529 13874
rect 5449 13814 5529 13840
rect 5169 10229 5249 10255
rect 5169 10195 5192 10229
rect 5226 10195 5249 10229
rect 5169 10187 5249 10195
rect 5309 10229 5389 10255
rect 5309 10195 5332 10229
rect 5366 10195 5389 10229
rect 5309 10187 5389 10195
rect 5449 10229 5529 10255
rect 5449 10195 5472 10229
rect 5506 10195 5529 10229
rect 5449 10187 5529 10195
rect 5589 10229 5669 10255
rect 5589 10195 5612 10229
rect 5646 10195 5669 10229
rect 5589 10187 5669 10195
rect 5729 10229 5809 10255
rect 5729 10195 5752 10229
rect 5786 10195 5809 10229
rect 5729 10187 5809 10195
rect 5869 10229 5949 10255
rect 5869 10195 5892 10229
rect 5926 10195 5949 10229
rect 5869 10187 5949 10195
rect 6009 10229 6089 10255
rect 6009 10195 6032 10229
rect 6066 10195 6089 10229
rect 6009 10187 6089 10195
rect 6149 10229 6229 10255
rect 6149 10195 6172 10229
rect 6206 10195 6229 10229
rect 6149 10187 6229 10195
<< mvndiffc >>
rect 5192 14707 5226 14741
rect 5332 13840 5366 13874
rect 5612 14707 5646 14741
rect 5752 14707 5786 14741
rect 5892 14707 5926 14741
rect 6032 14707 6066 14741
rect 6172 14707 6206 14741
rect 5472 13840 5506 13874
rect 5192 10195 5226 10229
rect 5332 10195 5366 10229
rect 5472 10195 5506 10229
rect 5612 10195 5646 10229
rect 5752 10195 5786 10229
rect 5892 10195 5926 10229
rect 6032 10195 6066 10229
rect 6172 10195 6206 10229
<< psubdiff >>
rect 10040 34512 10147 34546
rect 10181 34512 10215 34546
rect 10249 34512 10283 34546
rect 10317 34512 10351 34546
rect 10385 34512 10419 34546
rect 10453 34512 10487 34546
rect 10521 34512 10555 34546
rect 10589 34512 10623 34546
rect 10657 34512 10691 34546
rect 10725 34512 10759 34546
rect 10793 34512 10827 34546
rect 10861 34512 10895 34546
rect 10929 34512 10963 34546
rect 10997 34512 11031 34546
rect 11065 34512 11099 34546
rect 11133 34512 11167 34546
rect 11201 34512 11235 34546
rect 11269 34512 11303 34546
rect 11337 34512 11371 34546
rect 11405 34512 11439 34546
rect 11473 34512 11507 34546
rect 11541 34512 11575 34546
rect 11609 34512 11643 34546
rect 11677 34512 11711 34546
rect 11745 34512 11779 34546
rect 11813 34512 11847 34546
rect 11881 34512 11915 34546
rect 11949 34512 11983 34546
rect 12017 34512 12051 34546
rect 12085 34512 12119 34546
rect 12153 34512 12187 34546
rect 12221 34512 12255 34546
rect 12289 34512 12323 34546
rect 12357 34512 12391 34546
rect 12425 34512 12459 34546
rect 12493 34512 12527 34546
rect 12561 34512 12595 34546
rect 12629 34512 12663 34546
rect 12697 34512 12731 34546
rect 12765 34512 12799 34546
rect 12833 34512 12867 34546
rect 12901 34512 12935 34546
rect 12969 34512 13003 34546
rect 13037 34512 13071 34546
rect 13105 34512 13139 34546
rect 13173 34512 13207 34546
rect 13241 34512 13275 34546
rect 13309 34512 13343 34546
rect 13377 34512 13411 34546
rect 13445 34512 13479 34546
rect 13513 34512 13547 34546
rect 13581 34512 13615 34546
rect 13649 34512 13683 34546
rect 13717 34512 13751 34546
rect 13785 34512 13819 34546
rect 13853 34512 13887 34546
rect 13921 34512 13955 34546
rect 13989 34512 14023 34546
rect 14057 34512 14091 34546
rect 14125 34512 14193 34546
rect 10040 34478 10074 34512
rect 10040 34410 10074 34444
rect 10040 34342 10074 34376
rect 10040 34274 10074 34308
rect 10040 34206 10074 34240
rect 10040 34138 10074 34172
rect 10040 34070 10074 34104
rect 10040 34002 10074 34036
rect 10040 33934 10074 33968
rect 10040 33866 10074 33900
rect 10040 33798 10074 33832
rect 10040 33730 10074 33764
rect 10040 33662 10074 33696
rect 10040 33594 10074 33628
rect 10040 33526 10074 33560
rect 10040 33458 10074 33492
rect 10040 33390 10074 33424
rect 10040 33322 10074 33356
rect 10040 33254 10074 33288
rect 10040 33186 10074 33220
rect 10040 33118 10074 33152
rect 10040 33050 10074 33084
rect 10040 32982 10074 33016
rect 10040 32914 10074 32948
rect 10040 32846 10074 32880
rect 10040 32778 10074 32812
rect 10040 32710 10074 32744
rect 10040 32642 10074 32676
rect 10040 32574 10074 32608
rect 10040 32506 10074 32540
rect 10040 32438 10074 32472
rect 10040 32370 10074 32404
rect 10040 32302 10074 32336
rect 14159 34385 14193 34512
rect 14159 34317 14193 34351
rect 14159 34249 14193 34283
rect 14159 34181 14193 34215
rect 14159 34113 14193 34147
rect 14159 34045 14193 34079
rect 14159 33977 14193 34011
rect 14159 33909 14193 33943
rect 14159 33841 14193 33875
rect 14159 33773 14193 33807
rect 14159 33705 14193 33739
rect 14159 33637 14193 33671
rect 14159 33569 14193 33603
rect 14159 33501 14193 33535
rect 14159 33433 14193 33467
rect 14159 33365 14193 33399
rect 14159 33297 14193 33331
rect 14159 33229 14193 33263
rect 14159 33161 14193 33195
rect 14159 33093 14193 33127
rect 14159 33025 14193 33059
rect 14159 32957 14193 32991
rect 14159 32889 14193 32923
rect 14159 32821 14193 32855
rect 14159 32753 14193 32787
rect 14159 32685 14193 32719
rect 14159 32617 14193 32651
rect 14159 32549 14193 32583
rect 14159 32481 14193 32515
rect 14159 32413 14193 32447
rect 14159 32345 14193 32379
rect 14159 32294 14193 32311
rect 10074 32268 10108 32294
rect 10040 32260 10108 32268
rect 10142 32260 10193 32294
rect 10227 32260 10278 32294
rect 10312 32260 10363 32294
rect 10397 32260 10448 32294
rect 10482 32260 10533 32294
rect 10567 32260 10618 32294
rect 10652 32260 10703 32294
rect 10737 32260 10788 32294
rect 10822 32260 10873 32294
rect 10907 32260 10958 32294
rect 10992 32260 11043 32294
rect 11077 32260 11128 32294
rect 11162 32260 11213 32294
rect 11247 32260 11298 32294
rect 11332 32260 11383 32294
rect 11417 32260 11468 32294
rect 11502 32260 11553 32294
rect 11587 32260 11638 32294
rect 11672 32260 11723 32294
rect 11757 32260 11808 32294
rect 11842 32260 11893 32294
rect 11927 32260 11978 32294
rect 12012 32260 12063 32294
rect 12097 32260 12148 32294
rect 12182 32260 12233 32294
rect 12267 32260 12318 32294
rect 12352 32260 12403 32294
rect 12437 32260 12488 32294
rect 12522 32260 12573 32294
rect 12607 32260 12658 32294
rect 12692 32260 12743 32294
rect 12777 32260 12828 32294
rect 12862 32260 12913 32294
rect 12947 32260 12998 32294
rect 13032 32260 13083 32294
rect 13117 32260 13167 32294
rect 13201 32260 13251 32294
rect 13285 32260 13335 32294
rect 13369 32260 13419 32294
rect 13453 32260 13503 32294
rect 13537 32260 13587 32294
rect 13621 32260 13671 32294
rect 13705 32260 13755 32294
rect 13789 32260 13839 32294
rect 13873 32260 13923 32294
rect 13957 32260 14007 32294
rect 14041 32260 14091 32294
rect 14125 32277 14193 32294
rect 14125 32260 14159 32277
rect 10040 32234 10074 32260
rect 10040 32166 10074 32200
rect 14159 32209 14193 32243
rect 10040 32098 10074 32132
rect 10040 32030 10074 32064
rect 10040 31962 10074 31996
rect 10040 31894 10074 31928
rect 10040 31826 10074 31860
rect 10040 31758 10074 31792
rect 10040 31690 10074 31724
rect 10040 31622 10074 31656
rect 10040 31554 10074 31588
rect 10040 31486 10074 31520
rect 10040 31418 10074 31452
rect 10040 31350 10074 31384
rect 10040 31282 10074 31316
rect 10040 31214 10074 31248
rect 10040 31146 10074 31180
rect 10040 31078 10074 31112
rect 10040 31010 10074 31044
rect 10040 30942 10074 30976
rect 10040 30874 10074 30908
rect 10040 30806 10074 30840
rect 10040 30738 10074 30772
rect 10040 30670 10074 30704
rect 10040 30602 10074 30636
rect 10040 30534 10074 30568
rect 10040 30466 10074 30500
rect 10040 30398 10074 30432
rect 10040 30330 10074 30364
rect 10040 30262 10074 30296
rect 10040 30194 10074 30228
rect 10040 30126 10074 30160
rect 10040 30058 10074 30092
rect 14159 32141 14193 32175
rect 14159 32073 14193 32107
rect 14159 32005 14193 32039
rect 14159 31937 14193 31971
rect 14159 31869 14193 31903
rect 14159 31801 14193 31835
rect 14159 31733 14193 31767
rect 14159 31665 14193 31699
rect 14159 31597 14193 31631
rect 14159 31529 14193 31563
rect 14159 31461 14193 31495
rect 14159 31393 14193 31427
rect 14159 31325 14193 31359
rect 14159 31257 14193 31291
rect 14159 31189 14193 31223
rect 14159 31121 14193 31155
rect 14159 31053 14193 31087
rect 14159 30985 14193 31019
rect 14159 30917 14193 30951
rect 14159 30849 14193 30883
rect 14159 30781 14193 30815
rect 14159 30713 14193 30747
rect 14159 30645 14193 30679
rect 14159 30577 14193 30611
rect 14159 30509 14193 30543
rect 14159 30441 14193 30475
rect 14159 30373 14193 30407
rect 14159 30305 14193 30339
rect 14159 30237 14193 30271
rect 14159 30169 14193 30203
rect 14159 30101 14193 30135
rect 14159 30043 14193 30067
rect 10074 30024 10108 30043
rect 10040 30009 10108 30024
rect 10142 30009 10193 30043
rect 10227 30009 10278 30043
rect 10312 30009 10363 30043
rect 10397 30009 10448 30043
rect 10482 30009 10533 30043
rect 10567 30009 10618 30043
rect 10652 30009 10703 30043
rect 10737 30009 10788 30043
rect 10822 30009 10873 30043
rect 10907 30009 10958 30043
rect 10992 30009 11043 30043
rect 11077 30009 11128 30043
rect 11162 30009 11213 30043
rect 11247 30009 11298 30043
rect 11332 30009 11383 30043
rect 11417 30009 11468 30043
rect 11502 30009 11553 30043
rect 11587 30009 11638 30043
rect 11672 30009 11723 30043
rect 11757 30009 11808 30043
rect 11842 30009 11893 30043
rect 11927 30009 11978 30043
rect 12012 30009 12063 30043
rect 12097 30009 12148 30043
rect 12182 30009 12233 30043
rect 12267 30009 12318 30043
rect 12352 30009 12403 30043
rect 12437 30009 12488 30043
rect 12522 30009 12573 30043
rect 12607 30009 12658 30043
rect 12692 30009 12743 30043
rect 12777 30009 12828 30043
rect 12862 30009 12913 30043
rect 12947 30009 12998 30043
rect 13032 30009 13083 30043
rect 13117 30009 13167 30043
rect 13201 30009 13251 30043
rect 13285 30009 13335 30043
rect 13369 30009 13419 30043
rect 13453 30009 13503 30043
rect 13537 30009 13587 30043
rect 13621 30009 13671 30043
rect 13705 30009 13755 30043
rect 13789 30009 13839 30043
rect 13873 30009 13923 30043
rect 13957 30009 14007 30043
rect 14041 30009 14091 30043
rect 14125 30033 14193 30043
rect 14125 30009 14159 30033
rect 10040 29990 10074 30009
rect 10040 29922 10074 29956
rect 14159 29965 14193 29999
rect 10040 29854 10074 29888
rect 10040 29786 10074 29820
rect 10040 29718 10074 29752
rect 10040 29650 10074 29684
rect 10040 29582 10074 29616
rect 10040 29514 10074 29548
rect 10040 29446 10074 29480
rect 10040 29378 10074 29412
rect 10040 29310 10074 29344
rect 10040 29242 10074 29276
rect 10040 29174 10074 29208
rect 10040 29106 10074 29140
rect 10040 29038 10074 29072
rect 10040 28970 10074 29004
rect 10040 28902 10074 28936
rect 10040 28834 10074 28868
rect 10040 28766 10074 28800
rect 10040 28698 10074 28732
rect 10040 28630 10074 28664
rect 10040 28562 10074 28596
rect 10040 28494 10074 28528
rect 10040 28426 10074 28460
rect 10040 28358 10074 28392
rect 10040 28290 10074 28324
rect 10040 28222 10074 28256
rect 10040 28154 10074 28188
rect 10040 28086 10074 28120
rect 10040 28018 10074 28052
rect 10040 27950 10074 27984
rect 10040 27882 10074 27916
rect 10040 27789 10074 27848
rect 14159 29897 14193 29931
rect 14159 29829 14193 29863
rect 14159 29761 14193 29795
rect 14159 29693 14193 29727
rect 14159 29625 14193 29659
rect 14159 29557 14193 29591
rect 14159 29489 14193 29523
rect 14159 29421 14193 29455
rect 14159 29353 14193 29387
rect 14159 29285 14193 29319
rect 14159 29217 14193 29251
rect 14159 29149 14193 29183
rect 14159 29081 14193 29115
rect 14159 29013 14193 29047
rect 14159 28945 14193 28979
rect 14159 28877 14193 28911
rect 14159 28809 14193 28843
rect 14159 28741 14193 28775
rect 14159 28673 14193 28707
rect 14159 28605 14193 28639
rect 14159 28537 14193 28571
rect 14159 28469 14193 28503
rect 14159 28401 14193 28435
rect 14159 28333 14193 28367
rect 14159 28265 14193 28299
rect 14159 28197 14193 28231
rect 14159 28129 14193 28163
rect 14159 28061 14193 28095
rect 14159 27993 14193 28027
rect 14159 27925 14193 27959
rect 14159 27857 14193 27891
rect 14159 27789 14193 27823
rect 10040 27755 10108 27789
rect 10142 27755 10176 27789
rect 10210 27755 10244 27789
rect 10278 27755 10312 27789
rect 10346 27755 10380 27789
rect 10414 27755 10448 27789
rect 10482 27755 10516 27789
rect 10550 27755 10584 27789
rect 10618 27755 10652 27789
rect 10686 27755 10720 27789
rect 10754 27755 10788 27789
rect 10822 27755 10856 27789
rect 10890 27755 10924 27789
rect 10958 27755 10992 27789
rect 11026 27755 11060 27789
rect 11094 27755 11128 27789
rect 11162 27755 11196 27789
rect 11230 27755 11264 27789
rect 11298 27755 11332 27789
rect 11366 27755 11400 27789
rect 11434 27755 11468 27789
rect 11502 27755 11536 27789
rect 11570 27755 11604 27789
rect 11638 27755 11672 27789
rect 11706 27755 11740 27789
rect 11774 27755 11808 27789
rect 11842 27755 11876 27789
rect 11910 27755 11944 27789
rect 11978 27755 12012 27789
rect 12046 27755 12080 27789
rect 12114 27755 12148 27789
rect 12182 27755 12216 27789
rect 12250 27755 12284 27789
rect 12318 27755 12352 27789
rect 12386 27755 12420 27789
rect 12454 27755 12488 27789
rect 12522 27755 12556 27789
rect 12590 27755 12624 27789
rect 12658 27755 12692 27789
rect 12726 27755 12760 27789
rect 12794 27755 12828 27789
rect 12862 27755 12896 27789
rect 12930 27755 12964 27789
rect 12998 27755 13032 27789
rect 13066 27755 13100 27789
rect 13134 27755 13168 27789
rect 13202 27755 13236 27789
rect 13270 27755 13304 27789
rect 13338 27755 13372 27789
rect 13406 27755 13440 27789
rect 13474 27755 13508 27789
rect 13542 27755 13576 27789
rect 13610 27755 13644 27789
rect 13678 27755 13712 27789
rect 13746 27755 13780 27789
rect 13814 27755 13848 27789
rect 13882 27755 13916 27789
rect 13950 27755 13984 27789
rect 14018 27755 14052 27789
rect 14086 27755 14193 27789
<< nsubdiff >>
rect 9789 34762 9917 34796
rect 9951 34762 9985 34796
rect 10019 34762 10053 34796
rect 10087 34762 10121 34796
rect 10155 34762 10189 34796
rect 10223 34762 10257 34796
rect 10291 34762 10325 34796
rect 10359 34762 10393 34796
rect 10427 34762 10461 34796
rect 10495 34762 10529 34796
rect 10563 34762 10597 34796
rect 10631 34762 10665 34796
rect 10699 34762 10733 34796
rect 10767 34762 10801 34796
rect 10835 34762 10869 34796
rect 10903 34762 10937 34796
rect 10971 34762 11005 34796
rect 11039 34762 11073 34796
rect 11107 34762 11141 34796
rect 11175 34762 11209 34796
rect 11243 34762 11277 34796
rect 11311 34762 11345 34796
rect 11379 34762 11413 34796
rect 11447 34762 11481 34796
rect 11515 34762 11549 34796
rect 11583 34762 11617 34796
rect 11651 34762 11685 34796
rect 11719 34762 11753 34796
rect 11787 34762 11821 34796
rect 11855 34762 11889 34796
rect 11923 34762 11957 34796
rect 11991 34762 12025 34796
rect 12059 34762 12093 34796
rect 12127 34762 12161 34796
rect 12195 34762 12229 34796
rect 12263 34762 12297 34796
rect 12331 34762 12365 34796
rect 12399 34762 12433 34796
rect 12467 34762 12501 34796
rect 12535 34762 12569 34796
rect 12603 34762 12637 34796
rect 12671 34762 12705 34796
rect 12739 34762 12773 34796
rect 12807 34762 12841 34796
rect 12875 34762 12909 34796
rect 12943 34762 12977 34796
rect 13011 34762 13045 34796
rect 13079 34762 13113 34796
rect 13147 34762 13181 34796
rect 13215 34762 13249 34796
rect 13283 34762 13317 34796
rect 13351 34762 13385 34796
rect 13419 34762 13453 34796
rect 13487 34762 13521 34796
rect 13555 34762 13589 34796
rect 13623 34762 13657 34796
rect 13691 34762 13725 34796
rect 13759 34762 13793 34796
rect 13827 34762 13861 34796
rect 13895 34762 13929 34796
rect 13963 34762 13997 34796
rect 14031 34762 14065 34796
rect 14099 34762 14133 34796
rect 14167 34762 14201 34796
rect 14235 34762 14269 34796
rect 14303 34762 14337 34796
rect 14371 34762 14439 34796
rect 9789 34728 9823 34762
rect 9789 34660 9823 34694
rect 9789 34592 9823 34626
rect 9789 34524 9823 34558
rect 14405 34704 14439 34762
rect 9789 34456 9823 34490
rect 9789 34388 9823 34422
rect 9789 34320 9823 34354
rect 9789 34252 9823 34286
rect 9789 34184 9823 34218
rect 9789 34116 9823 34150
rect 9789 34048 9823 34082
rect 9789 33980 9823 34014
rect 9789 33912 9823 33946
rect 9789 33844 9823 33878
rect 9789 33776 9823 33810
rect 9789 33647 9823 33742
rect 9119 33613 9153 33647
rect 9119 33545 9153 33579
rect 9119 33477 9153 33511
rect 9119 33409 9153 33443
rect 9119 33341 9153 33375
rect 9119 33273 9153 33307
rect 9119 33205 9153 33239
rect 9119 33137 9153 33171
rect 9119 33069 9153 33103
rect 9119 33001 9153 33035
rect 9119 32933 9153 32967
rect 9119 32865 9153 32899
rect 9119 32797 9153 32831
rect 9119 32729 9153 32763
rect 9119 32661 9153 32695
rect 9119 32593 9153 32627
rect 9119 32525 9153 32559
rect 9119 32457 9153 32491
rect 9119 32389 9153 32423
rect 9119 32321 9153 32355
rect 9119 32253 9153 32287
rect 9119 32185 9153 32219
rect 9119 32117 9153 32151
rect 9119 32049 9153 32083
rect 9119 31981 9153 32015
rect 9119 31913 9153 31947
rect 9119 31845 9153 31879
rect 9119 31777 9153 31811
rect 9119 31709 9153 31743
rect 9119 31641 9153 31675
rect 9119 31573 9153 31607
rect 9119 31505 9153 31539
rect 9119 31437 9153 31471
rect 9119 31369 9153 31403
rect 9119 31301 9153 31335
rect 9119 31184 9153 31267
rect 9789 31150 9823 31184
rect 9789 31082 9823 31116
rect 9789 31014 9823 31048
rect 9789 30946 9823 30980
rect 9789 30878 9823 30912
rect 9789 30810 9823 30844
rect 9789 30742 9823 30776
rect 9789 30674 9823 30708
rect 9789 30606 9823 30640
rect 9789 30538 9823 30572
rect 9789 30470 9823 30504
rect 9789 30402 9823 30436
rect 9789 30334 9823 30368
rect 9789 30266 9823 30300
rect 9789 30198 9823 30232
rect 9789 30130 9823 30164
rect 9789 30062 9823 30096
rect 9789 29994 9823 30028
rect 9789 29926 9823 29960
rect 9789 29858 9823 29892
rect 9789 29790 9823 29824
rect 9789 29722 9823 29756
rect 9789 29654 9823 29688
rect 9789 29586 9823 29620
rect 9789 29518 9823 29552
rect 9789 29450 9823 29484
rect 9789 29382 9823 29416
rect 9789 29314 9823 29348
rect 9789 29246 9823 29280
rect 9789 29178 9823 29212
rect 9789 29110 9823 29144
rect 9789 29042 9823 29076
rect 9789 28974 9823 29008
rect 9789 28906 9823 28940
rect 9789 28838 9823 28872
rect 9789 28770 9823 28804
rect 9789 28702 9823 28736
rect 9789 28634 9823 28668
rect 9789 28566 9823 28600
rect 9789 28498 9823 28532
rect 9789 28430 9823 28464
rect 9789 28362 9823 28396
rect 9789 28294 9823 28328
rect 9789 28226 9823 28260
rect 9789 28158 9823 28192
rect 9789 28090 9823 28124
rect 9789 28022 9823 28056
rect 9789 27954 9823 27988
rect 9789 27886 9823 27920
rect 9789 27818 9823 27852
rect 9789 27750 9823 27784
rect 14405 34540 14439 34670
rect 14405 34472 14439 34506
rect 14405 34404 14439 34438
rect 14405 34336 14439 34370
rect 14405 34268 14439 34302
rect 14405 34200 14439 34234
rect 14405 34132 14439 34166
rect 14405 34064 14439 34098
rect 14405 33996 14439 34030
rect 14405 33928 14439 33962
rect 14405 33860 14439 33894
rect 14405 33792 14439 33826
rect 14405 33724 14439 33758
rect 14405 33656 14439 33690
rect 14405 33588 14439 33622
rect 14405 33520 14439 33554
rect 14405 33452 14439 33486
rect 14405 33384 14439 33418
rect 14405 33316 14439 33350
rect 14405 33248 14439 33282
rect 14405 33180 14439 33214
rect 14405 33112 14439 33146
rect 14405 33044 14439 33078
rect 14405 32976 14439 33010
rect 14405 32908 14439 32942
rect 14405 32840 14439 32874
rect 14405 32772 14439 32806
rect 14405 32704 14439 32738
rect 14405 32636 14439 32670
rect 14405 32568 14439 32602
rect 14405 32500 14439 32534
rect 14405 32432 14439 32466
rect 14405 32364 14439 32398
rect 14405 32296 14439 32330
rect 14405 32228 14439 32262
rect 14405 32160 14439 32194
rect 14405 32092 14439 32126
rect 14405 32024 14439 32058
rect 14405 31956 14439 31990
rect 14405 31888 14439 31922
rect 14405 31820 14439 31854
rect 14405 31752 14439 31786
rect 14405 31684 14439 31718
rect 14405 31616 14439 31650
rect 14405 31548 14439 31582
rect 14405 31480 14439 31514
rect 14405 31412 14439 31446
rect 14405 31344 14439 31378
rect 14405 31276 14439 31310
rect 14405 31208 14439 31242
rect 14405 31140 14439 31174
rect 14405 31072 14439 31106
rect 14405 31004 14439 31038
rect 14405 30936 14439 30970
rect 14405 30868 14439 30902
rect 14405 30800 14439 30834
rect 14405 30732 14439 30766
rect 14405 30664 14439 30698
rect 14405 30596 14439 30630
rect 14405 30528 14439 30562
rect 14405 30460 14439 30494
rect 14405 30392 14439 30426
rect 14405 30324 14439 30358
rect 14405 30256 14439 30290
rect 14405 30188 14439 30222
rect 14405 30120 14439 30154
rect 14405 30052 14439 30086
rect 14405 29984 14439 30018
rect 14405 29916 14439 29950
rect 14405 29848 14439 29882
rect 14405 29780 14439 29814
rect 14405 29712 14439 29746
rect 14405 29644 14439 29678
rect 14405 29576 14439 29610
rect 14405 29508 14439 29542
rect 14405 29440 14439 29474
rect 14405 29372 14439 29406
rect 14405 29304 14439 29338
rect 14405 29236 14439 29270
rect 14405 29168 14439 29202
rect 14405 29100 14439 29134
rect 14405 29032 14439 29066
rect 14405 28964 14439 28998
rect 14405 28896 14439 28930
rect 14405 28828 14439 28862
rect 14405 28760 14439 28794
rect 14405 28692 14439 28726
rect 14405 28624 14439 28658
rect 14405 28556 14439 28590
rect 14405 28488 14439 28522
rect 14405 28420 14439 28454
rect 14405 28352 14439 28386
rect 14405 28284 14439 28318
rect 14405 28216 14439 28250
rect 14405 28148 14439 28182
rect 14405 28080 14439 28114
rect 14405 28012 14439 28046
rect 14405 27944 14439 27978
rect 14405 27876 14439 27910
rect 14405 27808 14439 27842
rect 9789 27682 9823 27716
rect 9789 27614 9823 27648
rect 9789 27546 9823 27580
rect 14405 27740 14439 27774
rect 14405 27672 14439 27706
rect 14405 27604 14439 27638
rect 14405 27536 14439 27570
rect 9789 27478 9823 27512
rect 12432 27502 12500 27536
rect 12534 27502 12568 27536
rect 12602 27502 12636 27536
rect 12670 27502 12704 27536
rect 12738 27502 12772 27536
rect 12806 27502 12840 27536
rect 12874 27502 12908 27536
rect 12942 27502 12976 27536
rect 13010 27502 13044 27536
rect 13078 27502 13112 27536
rect 13146 27502 13180 27536
rect 13214 27502 13248 27536
rect 13282 27502 13316 27536
rect 13350 27502 13384 27536
rect 13418 27502 13452 27536
rect 13486 27502 13520 27536
rect 13554 27502 13588 27536
rect 13622 27502 13656 27536
rect 13690 27502 13724 27536
rect 13758 27502 13792 27536
rect 13826 27502 13860 27536
rect 13894 27502 13928 27536
rect 13962 27502 13996 27536
rect 14030 27502 14064 27536
rect 14098 27502 14132 27536
rect 14166 27502 14200 27536
rect 14234 27502 14268 27536
rect 14302 27502 14336 27536
rect 14370 27502 14439 27536
rect 9789 27410 9823 27444
rect 9789 27342 9823 27376
rect 9789 27274 9823 27308
rect 9789 27206 9823 27240
rect 9789 27138 9823 27172
rect 9789 27070 9823 27104
rect 9789 27002 9823 27036
rect 9789 26934 9823 26968
rect 9789 26866 9823 26900
rect 9789 26798 9823 26832
rect 9789 26730 9823 26764
rect 9789 26662 9823 26696
rect 12432 27424 12466 27502
rect 12432 27356 12466 27390
rect 12432 27288 12466 27322
rect 12432 27220 12466 27254
rect 12432 27152 12466 27186
rect 12432 27084 12466 27118
rect 12432 27016 12466 27050
rect 12432 26948 12466 26982
rect 12432 26880 12466 26914
rect 12432 26812 12466 26846
rect 12432 26744 12466 26778
rect 12432 26676 12466 26710
rect 9789 26594 9823 26628
rect 9789 26526 9823 26560
rect 9789 26404 9823 26492
rect 12432 26608 12466 26642
rect 12432 26540 12466 26574
rect 12432 26472 12466 26506
rect 12432 26404 12466 26438
rect 9789 26370 9857 26404
rect 9891 26370 9925 26404
rect 9959 26370 9993 26404
rect 10027 26370 10061 26404
rect 10095 26370 10129 26404
rect 10163 26370 10197 26404
rect 10231 26370 10265 26404
rect 10299 26370 10333 26404
rect 10367 26370 10401 26404
rect 10435 26370 10469 26404
rect 10503 26370 10537 26404
rect 10571 26370 10605 26404
rect 10639 26370 10673 26404
rect 10707 26370 10741 26404
rect 10775 26370 10809 26404
rect 10843 26370 10877 26404
rect 10911 26370 10945 26404
rect 10979 26370 11013 26404
rect 11047 26370 11081 26404
rect 11115 26370 11149 26404
rect 11183 26370 11217 26404
rect 11251 26370 11285 26404
rect 11319 26370 11353 26404
rect 11387 26370 11421 26404
rect 11455 26370 11489 26404
rect 11523 26370 11557 26404
rect 11591 26370 11625 26404
rect 11659 26370 11693 26404
rect 11727 26370 11761 26404
rect 11795 26370 11829 26404
rect 11863 26370 11897 26404
rect 11931 26370 11965 26404
rect 11999 26370 12033 26404
rect 12067 26370 12101 26404
rect 12135 26370 12169 26404
rect 12203 26370 12237 26404
rect 12271 26370 12305 26404
rect 12339 26370 12466 26404
<< mvpsubdiff >>
rect 5059 15813 5684 15814
rect 5059 15780 5140 15813
rect 5059 15746 5060 15780
rect 5094 15779 5140 15780
rect 5174 15779 5208 15813
rect 5242 15779 5276 15813
rect 5310 15779 5344 15813
rect 5378 15779 5412 15813
rect 5446 15779 5480 15813
rect 5514 15779 5548 15813
rect 5582 15779 5616 15813
rect 5650 15779 5684 15813
rect 5094 15778 5684 15779
rect 5094 15746 5095 15778
rect 5059 15712 5095 15746
rect 5059 15678 5060 15712
rect 5094 15678 5095 15712
rect 5059 15644 5095 15678
rect 5648 15686 5684 15778
rect 5059 15610 5060 15644
rect 5094 15610 5095 15644
rect 5059 15576 5095 15610
rect 5059 15542 5060 15576
rect 5094 15542 5095 15576
rect 5059 15508 5095 15542
rect 5059 15474 5060 15508
rect 5094 15474 5095 15508
rect 5059 15440 5095 15474
rect 5059 15406 5060 15440
rect 5094 15406 5095 15440
rect 5059 15372 5095 15406
rect 5059 15338 5060 15372
rect 5094 15338 5095 15372
rect 5059 15304 5095 15338
rect 5059 15270 5060 15304
rect 5094 15270 5095 15304
rect 5059 15236 5095 15270
rect 5059 15202 5060 15236
rect 5094 15202 5095 15236
rect 5059 15168 5095 15202
rect 5059 15134 5060 15168
rect 5094 15134 5095 15168
rect 5059 15100 5095 15134
rect 5059 15066 5060 15100
rect 5094 15066 5095 15100
rect 5059 14974 5095 15066
rect 5648 15652 5649 15686
rect 5683 15652 5684 15686
rect 5648 15618 5684 15652
rect 5648 15584 5649 15618
rect 5683 15584 5684 15618
rect 5648 15550 5684 15584
rect 5648 15516 5649 15550
rect 5683 15516 5684 15550
rect 5648 15482 5684 15516
rect 5648 15448 5649 15482
rect 5683 15448 5684 15482
rect 5648 15414 5684 15448
rect 5648 15380 5649 15414
rect 5683 15380 5684 15414
rect 5648 15346 5684 15380
rect 5648 15312 5649 15346
rect 5683 15312 5684 15346
rect 5648 15278 5684 15312
rect 5648 15244 5649 15278
rect 5683 15244 5684 15278
rect 5648 15210 5684 15244
rect 5648 15176 5649 15210
rect 5683 15176 5684 15210
rect 5648 15142 5684 15176
rect 5648 15108 5649 15142
rect 5683 15108 5684 15142
rect 5648 15074 5684 15108
rect 5648 15040 5649 15074
rect 5683 15040 5684 15074
rect 5648 15006 5684 15040
rect 5648 14974 5649 15006
rect 5059 14973 5649 14974
rect 5059 14939 5093 14973
rect 5127 14939 5161 14973
rect 5195 14939 5229 14973
rect 5263 14939 5297 14973
rect 5331 14939 5365 14973
rect 5399 14939 5433 14973
rect 5467 14939 5501 14973
rect 5535 14939 5569 14973
rect 5603 14972 5649 14973
rect 5683 14972 5684 15006
rect 5603 14939 5684 14972
rect 5059 14938 5684 14939
rect 5059 14858 6339 14859
rect 5059 14824 5093 14858
rect 5127 14824 5161 14858
rect 5195 14824 5229 14858
rect 5263 14824 5297 14858
rect 5331 14824 5365 14858
rect 5399 14824 5433 14858
rect 5467 14824 5501 14858
rect 5535 14824 5569 14858
rect 5603 14824 5637 14858
rect 5671 14824 5705 14858
rect 5739 14824 5773 14858
rect 5807 14824 5841 14858
rect 5875 14824 5909 14858
rect 5943 14824 5977 14858
rect 6011 14824 6045 14858
rect 6079 14824 6113 14858
rect 6147 14824 6181 14858
rect 6215 14825 6339 14858
rect 6215 14824 6304 14825
rect 5059 14823 6304 14824
rect 5059 14769 5095 14823
rect 5059 14735 5060 14769
rect 5094 14735 5095 14769
rect 6303 14791 6304 14823
rect 6338 14791 6339 14825
rect 6303 14757 6339 14791
rect 5059 14701 5095 14735
rect 5059 14667 5060 14701
rect 5094 14667 5095 14701
rect 5059 14633 5095 14667
rect 5059 14599 5060 14633
rect 5094 14599 5095 14633
rect 5059 14565 5095 14599
rect 5059 14531 5060 14565
rect 5094 14531 5095 14565
rect 5059 14497 5095 14531
rect 5059 14463 5060 14497
rect 5094 14463 5095 14497
rect 5059 14429 5095 14463
rect 5059 14395 5060 14429
rect 5094 14395 5095 14429
rect 5059 14361 5095 14395
rect 5059 14327 5060 14361
rect 5094 14327 5095 14361
rect 5059 14293 5095 14327
rect 5059 14259 5060 14293
rect 5094 14259 5095 14293
rect 5059 14225 5095 14259
rect 5059 14191 5060 14225
rect 5094 14191 5095 14225
rect 5059 14157 5095 14191
rect 5059 14123 5060 14157
rect 5094 14123 5095 14157
rect 5059 14089 5095 14123
rect 5059 14055 5060 14089
rect 5094 14055 5095 14089
rect 5059 14021 5095 14055
rect 5059 13987 5060 14021
rect 5094 13987 5095 14021
rect 5059 13953 5095 13987
rect 5059 13919 5060 13953
rect 5094 13919 5095 13953
rect 5059 13885 5095 13919
rect 5059 13851 5060 13885
rect 5094 13851 5095 13885
rect 5059 13817 5095 13851
rect 5059 13783 5060 13817
rect 5094 13783 5095 13817
rect 6303 14723 6304 14757
rect 6338 14723 6339 14757
rect 6303 14689 6339 14723
rect 6303 14655 6304 14689
rect 6338 14655 6339 14689
rect 6303 14621 6339 14655
rect 6303 14587 6304 14621
rect 6338 14587 6339 14621
rect 6303 14553 6339 14587
rect 6303 14519 6304 14553
rect 6338 14519 6339 14553
rect 6303 14485 6339 14519
rect 6303 14451 6304 14485
rect 6338 14451 6339 14485
rect 6303 14417 6339 14451
rect 6303 14383 6304 14417
rect 6338 14383 6339 14417
rect 6303 14349 6339 14383
rect 6303 14315 6304 14349
rect 6338 14315 6339 14349
rect 6303 14281 6339 14315
rect 6303 14247 6304 14281
rect 6338 14247 6339 14281
rect 6303 14213 6339 14247
rect 6303 14179 6304 14213
rect 6338 14179 6339 14213
rect 6303 14145 6339 14179
rect 6303 14111 6304 14145
rect 6338 14111 6339 14145
rect 6303 14077 6339 14111
rect 6303 14043 6304 14077
rect 6338 14043 6339 14077
rect 6303 14009 6339 14043
rect 6303 13975 6304 14009
rect 6338 13975 6339 14009
rect 6303 13941 6339 13975
rect 6303 13907 6304 13941
rect 6338 13907 6339 13941
rect 6303 13873 6339 13907
rect 6303 13839 6304 13873
rect 6338 13839 6339 13873
rect 5059 13749 5095 13783
rect 5059 13715 5060 13749
rect 5094 13715 5095 13749
rect 5059 13681 5095 13715
rect 5059 13647 5060 13681
rect 5094 13647 5095 13681
rect 5059 13613 5095 13647
rect 5059 13579 5060 13613
rect 5094 13579 5095 13613
rect 5059 13545 5095 13579
rect 5059 13511 5060 13545
rect 5094 13511 5095 13545
rect 5059 13477 5095 13511
rect 5059 13443 5060 13477
rect 5094 13443 5095 13477
rect 5059 13409 5095 13443
rect 5059 13375 5060 13409
rect 5094 13375 5095 13409
rect 5059 13341 5095 13375
rect 5059 13307 5060 13341
rect 5094 13307 5095 13341
rect 5059 13273 5095 13307
rect 5059 13239 5060 13273
rect 5094 13239 5095 13273
rect 5059 13205 5095 13239
rect 5059 13171 5060 13205
rect 5094 13171 5095 13205
rect 5059 13137 5095 13171
rect 5059 13103 5060 13137
rect 5094 13103 5095 13137
rect 5059 13069 5095 13103
rect 5059 13035 5060 13069
rect 5094 13035 5095 13069
rect 5059 13001 5095 13035
rect 5059 12967 5060 13001
rect 5094 12967 5095 13001
rect 5059 12933 5095 12967
rect 5059 12899 5060 12933
rect 5094 12899 5095 12933
rect 5059 12865 5095 12899
rect 5059 12831 5060 12865
rect 5094 12831 5095 12865
rect 5059 12797 5095 12831
rect 5059 12763 5060 12797
rect 5094 12763 5095 12797
rect 5059 12729 5095 12763
rect 5059 12695 5060 12729
rect 5094 12695 5095 12729
rect 5059 12661 5095 12695
rect 5059 12627 5060 12661
rect 5094 12627 5095 12661
rect 5059 12593 5095 12627
rect 5059 12559 5060 12593
rect 5094 12559 5095 12593
rect 5059 12525 5095 12559
rect 5059 12491 5060 12525
rect 5094 12491 5095 12525
rect 5059 12457 5095 12491
rect 5059 12423 5060 12457
rect 5094 12423 5095 12457
rect 5059 12389 5095 12423
rect 5059 12355 5060 12389
rect 5094 12355 5095 12389
rect 5059 12321 5095 12355
rect 5059 12287 5060 12321
rect 5094 12287 5095 12321
rect 5059 12253 5095 12287
rect 5059 12219 5060 12253
rect 5094 12219 5095 12253
rect 5059 12185 5095 12219
rect 5059 12151 5060 12185
rect 5094 12151 5095 12185
rect 5059 12117 5095 12151
rect 661 11926 697 11960
rect 661 11892 662 11926
rect 696 11892 697 11926
rect 661 11858 697 11892
rect 661 11824 662 11858
rect 696 11824 697 11858
rect 661 11790 697 11824
rect 661 11756 662 11790
rect 696 11756 697 11790
rect 661 11722 697 11756
rect 661 11688 662 11722
rect 696 11688 697 11722
rect 661 11654 697 11688
rect 661 11620 662 11654
rect 696 11620 697 11654
rect 661 11586 697 11620
rect 661 11552 662 11586
rect 696 11552 697 11586
rect 661 11518 697 11552
rect 661 11484 662 11518
rect 696 11484 697 11518
rect 661 11450 697 11484
rect 661 11416 662 11450
rect 696 11416 697 11450
rect 661 11382 697 11416
rect 661 11348 662 11382
rect 696 11348 697 11382
rect 661 11314 697 11348
rect 661 11280 662 11314
rect 696 11280 697 11314
rect 661 11246 697 11280
rect 661 11212 662 11246
rect 696 11212 697 11246
rect 661 11178 697 11212
rect 661 11144 662 11178
rect 696 11144 697 11178
rect 661 11110 697 11144
rect 661 11076 662 11110
rect 696 11076 697 11110
rect 661 11042 697 11076
rect 661 11008 662 11042
rect 696 11008 697 11042
rect 661 10974 697 11008
rect 661 10940 662 10974
rect 696 10940 697 10974
rect 661 10906 697 10940
rect 661 10872 662 10906
rect 696 10872 697 10906
rect 661 10838 697 10872
rect 661 10804 662 10838
rect 696 10804 697 10838
rect 661 10770 697 10804
rect 661 10736 662 10770
rect 696 10736 697 10770
rect 661 10702 697 10736
rect 661 10668 662 10702
rect 696 10668 697 10702
rect 661 10634 697 10668
rect 661 10600 662 10634
rect 696 10600 697 10634
rect 661 10566 697 10600
rect 661 10532 662 10566
rect 696 10532 697 10566
rect 661 10498 697 10532
rect 661 10464 662 10498
rect 696 10464 697 10498
rect 661 10430 697 10464
rect 661 10396 662 10430
rect 696 10396 697 10430
rect 661 10362 697 10396
rect 661 10328 662 10362
rect 696 10328 697 10362
rect 661 10294 697 10328
rect 661 10260 662 10294
rect 696 10260 697 10294
rect 661 10226 697 10260
rect 661 10192 662 10226
rect 696 10192 697 10226
rect 661 10158 697 10192
rect 661 10124 662 10158
rect 696 10124 697 10158
rect 661 10090 697 10124
rect 661 10056 662 10090
rect 696 10056 697 10090
rect 661 10022 697 10056
rect 661 9988 662 10022
rect 696 9988 697 10022
rect 661 9887 697 9988
rect 2311 11859 2347 11960
rect 2311 11825 2312 11859
rect 2346 11825 2347 11859
rect 2311 11791 2347 11825
rect 2311 11757 2312 11791
rect 2346 11757 2347 11791
rect 2311 11723 2347 11757
rect 2311 11689 2312 11723
rect 2346 11689 2347 11723
rect 2311 11655 2347 11689
rect 2311 11621 2312 11655
rect 2346 11621 2347 11655
rect 2311 11587 2347 11621
rect 2311 11553 2312 11587
rect 2346 11553 2347 11587
rect 2311 11519 2347 11553
rect 2311 11485 2312 11519
rect 2346 11485 2347 11519
rect 2311 11451 2347 11485
rect 2311 11417 2312 11451
rect 2346 11417 2347 11451
rect 2311 11383 2347 11417
rect 2311 11349 2312 11383
rect 2346 11349 2347 11383
rect 2311 11315 2347 11349
rect 2311 11281 2312 11315
rect 2346 11281 2347 11315
rect 2311 11247 2347 11281
rect 2311 11213 2312 11247
rect 2346 11213 2347 11247
rect 2311 11179 2347 11213
rect 2311 11145 2312 11179
rect 2346 11145 2347 11179
rect 2311 11111 2347 11145
rect 2311 11077 2312 11111
rect 2346 11077 2347 11111
rect 2311 11043 2347 11077
rect 2311 11009 2312 11043
rect 2346 11009 2347 11043
rect 2311 10975 2347 11009
rect 2311 10941 2312 10975
rect 2346 10941 2347 10975
rect 2311 10907 2347 10941
rect 2311 10873 2312 10907
rect 2346 10873 2347 10907
rect 2311 10839 2347 10873
rect 2311 10805 2312 10839
rect 2346 10805 2347 10839
rect 2311 10771 2347 10805
rect 2311 10737 2312 10771
rect 2346 10737 2347 10771
rect 2311 10703 2347 10737
rect 2311 10669 2312 10703
rect 2346 10669 2347 10703
rect 2311 10635 2347 10669
rect 2311 10601 2312 10635
rect 2346 10601 2347 10635
rect 2311 10567 2347 10601
rect 2311 10533 2312 10567
rect 2346 10533 2347 10567
rect 2311 10499 2347 10533
rect 2311 10465 2312 10499
rect 2346 10465 2347 10499
rect 2311 10431 2347 10465
rect 2311 10397 2312 10431
rect 2346 10397 2347 10431
rect 2311 10363 2347 10397
rect 2311 10329 2312 10363
rect 2346 10329 2347 10363
rect 2311 10295 2347 10329
rect 2311 10261 2312 10295
rect 2346 10261 2347 10295
rect 2311 10227 2347 10261
rect 2311 10193 2312 10227
rect 2346 10193 2347 10227
rect 2311 10159 2347 10193
rect 2311 10125 2312 10159
rect 2346 10125 2347 10159
rect 2311 10091 2347 10125
rect 2311 10057 2312 10091
rect 2346 10057 2347 10091
rect 2311 10023 2347 10057
rect 2311 9989 2312 10023
rect 2346 9989 2347 10023
rect 2311 9955 2347 9989
rect 2311 9921 2312 9955
rect 2346 9921 2347 9955
rect 2311 9887 2347 9921
rect 2689 11926 2725 11960
rect 2689 11892 2690 11926
rect 2724 11892 2725 11926
rect 2689 11858 2725 11892
rect 2689 11824 2690 11858
rect 2724 11824 2725 11858
rect 2689 11790 2725 11824
rect 2689 11756 2690 11790
rect 2724 11756 2725 11790
rect 2689 11722 2725 11756
rect 2689 11688 2690 11722
rect 2724 11688 2725 11722
rect 2689 11654 2725 11688
rect 2689 11620 2690 11654
rect 2724 11620 2725 11654
rect 2689 11586 2725 11620
rect 2689 11552 2690 11586
rect 2724 11552 2725 11586
rect 2689 11518 2725 11552
rect 2689 11484 2690 11518
rect 2724 11484 2725 11518
rect 2689 11450 2725 11484
rect 2689 11416 2690 11450
rect 2724 11416 2725 11450
rect 2689 11382 2725 11416
rect 2689 11348 2690 11382
rect 2724 11348 2725 11382
rect 2689 11314 2725 11348
rect 2689 11280 2690 11314
rect 2724 11280 2725 11314
rect 2689 11246 2725 11280
rect 2689 11212 2690 11246
rect 2724 11212 2725 11246
rect 2689 11178 2725 11212
rect 2689 11144 2690 11178
rect 2724 11144 2725 11178
rect 2689 11110 2725 11144
rect 2689 11076 2690 11110
rect 2724 11076 2725 11110
rect 2689 11042 2725 11076
rect 2689 11008 2690 11042
rect 2724 11008 2725 11042
rect 2689 10974 2725 11008
rect 2689 10940 2690 10974
rect 2724 10940 2725 10974
rect 2689 10906 2725 10940
rect 2689 10872 2690 10906
rect 2724 10872 2725 10906
rect 2689 10838 2725 10872
rect 2689 10804 2690 10838
rect 2724 10804 2725 10838
rect 2689 10770 2725 10804
rect 2689 10736 2690 10770
rect 2724 10736 2725 10770
rect 2689 10702 2725 10736
rect 2689 10668 2690 10702
rect 2724 10668 2725 10702
rect 2689 10634 2725 10668
rect 2689 10600 2690 10634
rect 2724 10600 2725 10634
rect 2689 10566 2725 10600
rect 2689 10532 2690 10566
rect 2724 10532 2725 10566
rect 2689 10498 2725 10532
rect 2689 10464 2690 10498
rect 2724 10464 2725 10498
rect 2689 10430 2725 10464
rect 2689 10396 2690 10430
rect 2724 10396 2725 10430
rect 2689 10362 2725 10396
rect 2689 10328 2690 10362
rect 2724 10328 2725 10362
rect 2689 10294 2725 10328
rect 2689 10260 2690 10294
rect 2724 10260 2725 10294
rect 2689 10226 2725 10260
rect 2689 10192 2690 10226
rect 2724 10192 2725 10226
rect 2689 10158 2725 10192
rect 2689 10124 2690 10158
rect 2724 10124 2725 10158
rect 2689 10090 2725 10124
rect 2689 10056 2690 10090
rect 2724 10056 2725 10090
rect 2689 10022 2725 10056
rect 2689 9988 2690 10022
rect 2724 9988 2725 10022
rect 2689 9887 2725 9988
rect 4339 11859 4375 11960
rect 4339 11825 4340 11859
rect 4374 11825 4375 11859
rect 4339 11791 4375 11825
rect 4339 11757 4340 11791
rect 4374 11757 4375 11791
rect 4339 11723 4375 11757
rect 4339 11689 4340 11723
rect 4374 11689 4375 11723
rect 4339 11655 4375 11689
rect 4339 11621 4340 11655
rect 4374 11621 4375 11655
rect 4339 11587 4375 11621
rect 4339 11553 4340 11587
rect 4374 11553 4375 11587
rect 4339 11519 4375 11553
rect 4339 11485 4340 11519
rect 4374 11485 4375 11519
rect 4339 11451 4375 11485
rect 4339 11417 4340 11451
rect 4374 11417 4375 11451
rect 4339 11383 4375 11417
rect 4339 11349 4340 11383
rect 4374 11349 4375 11383
rect 4339 11315 4375 11349
rect 4339 11281 4340 11315
rect 4374 11281 4375 11315
rect 4339 11247 4375 11281
rect 4339 11213 4340 11247
rect 4374 11213 4375 11247
rect 4339 11179 4375 11213
rect 4339 11145 4340 11179
rect 4374 11145 4375 11179
rect 4339 11111 4375 11145
rect 4339 11077 4340 11111
rect 4374 11077 4375 11111
rect 4339 11043 4375 11077
rect 4339 11009 4340 11043
rect 4374 11009 4375 11043
rect 4339 10975 4375 11009
rect 4339 10941 4340 10975
rect 4374 10941 4375 10975
rect 4339 10907 4375 10941
rect 4339 10873 4340 10907
rect 4374 10873 4375 10907
rect 4339 10839 4375 10873
rect 4339 10805 4340 10839
rect 4374 10805 4375 10839
rect 4339 10771 4375 10805
rect 4339 10737 4340 10771
rect 4374 10737 4375 10771
rect 4339 10703 4375 10737
rect 4339 10669 4340 10703
rect 4374 10669 4375 10703
rect 4339 10635 4375 10669
rect 4339 10601 4340 10635
rect 4374 10601 4375 10635
rect 4339 10567 4375 10601
rect 4339 10533 4340 10567
rect 4374 10533 4375 10567
rect 4339 10499 4375 10533
rect 4339 10465 4340 10499
rect 4374 10465 4375 10499
rect 4339 10431 4375 10465
rect 4339 10397 4340 10431
rect 4374 10397 4375 10431
rect 4339 10363 4375 10397
rect 4339 10329 4340 10363
rect 4374 10329 4375 10363
rect 4339 10295 4375 10329
rect 4339 10261 4340 10295
rect 4374 10261 4375 10295
rect 4339 10227 4375 10261
rect 4339 10193 4340 10227
rect 4374 10193 4375 10227
rect 4339 10159 4375 10193
rect 4339 10125 4340 10159
rect 4374 10125 4375 10159
rect 4339 10091 4375 10125
rect 4339 10057 4340 10091
rect 4374 10057 4375 10091
rect 4339 10023 4375 10057
rect 4339 9989 4340 10023
rect 4374 9989 4375 10023
rect 4339 9955 4375 9989
rect 4339 9921 4340 9955
rect 4374 9921 4375 9955
rect 4339 9887 4375 9921
rect 5059 12083 5060 12117
rect 5094 12083 5095 12117
rect 5059 12049 5095 12083
rect 5059 12015 5060 12049
rect 5094 12015 5095 12049
rect 5059 11981 5095 12015
rect 5059 11947 5060 11981
rect 5094 11947 5095 11981
rect 5059 11913 5095 11947
rect 5059 11879 5060 11913
rect 5094 11879 5095 11913
rect 5059 11845 5095 11879
rect 5059 11811 5060 11845
rect 5094 11811 5095 11845
rect 5059 11777 5095 11811
rect 5059 11743 5060 11777
rect 5094 11743 5095 11777
rect 5059 11709 5095 11743
rect 5059 11675 5060 11709
rect 5094 11675 5095 11709
rect 5059 11641 5095 11675
rect 5059 11607 5060 11641
rect 5094 11607 5095 11641
rect 5059 11573 5095 11607
rect 5059 11539 5060 11573
rect 5094 11539 5095 11573
rect 5059 11505 5095 11539
rect 5059 11471 5060 11505
rect 5094 11471 5095 11505
rect 5059 11437 5095 11471
rect 5059 11403 5060 11437
rect 5094 11403 5095 11437
rect 5059 11369 5095 11403
rect 5059 11335 5060 11369
rect 5094 11335 5095 11369
rect 5059 11301 5095 11335
rect 5059 11267 5060 11301
rect 5094 11267 5095 11301
rect 5059 11233 5095 11267
rect 5059 11199 5060 11233
rect 5094 11199 5095 11233
rect 5059 11165 5095 11199
rect 5059 11131 5060 11165
rect 5094 11131 5095 11165
rect 5059 11097 5095 11131
rect 5059 11063 5060 11097
rect 5094 11063 5095 11097
rect 5059 11029 5095 11063
rect 5059 10995 5060 11029
rect 5094 10995 5095 11029
rect 5059 10961 5095 10995
rect 5059 10927 5060 10961
rect 5094 10927 5095 10961
rect 5059 10893 5095 10927
rect 5059 10859 5060 10893
rect 5094 10859 5095 10893
rect 5059 10825 5095 10859
rect 5059 10791 5060 10825
rect 5094 10791 5095 10825
rect 5059 10757 5095 10791
rect 5059 10723 5060 10757
rect 5094 10723 5095 10757
rect 5059 10689 5095 10723
rect 5059 10655 5060 10689
rect 5094 10655 5095 10689
rect 5059 10621 5095 10655
rect 5059 10587 5060 10621
rect 5094 10587 5095 10621
rect 5059 10553 5095 10587
rect 5059 10519 5060 10553
rect 5094 10519 5095 10553
rect 5059 10485 5095 10519
rect 5059 10451 5060 10485
rect 5094 10451 5095 10485
rect 5059 10417 5095 10451
rect 5059 10383 5060 10417
rect 5094 10383 5095 10417
rect 5059 10349 5095 10383
rect 5059 10315 5060 10349
rect 5094 10315 5095 10349
rect 5059 10281 5095 10315
rect 5059 10247 5060 10281
rect 5094 10247 5095 10281
rect 6303 13805 6339 13839
rect 6303 13771 6304 13805
rect 6338 13771 6339 13805
rect 6303 13737 6339 13771
rect 6303 13703 6304 13737
rect 6338 13703 6339 13737
rect 6303 13669 6339 13703
rect 6303 13635 6304 13669
rect 6338 13635 6339 13669
rect 6303 13601 6339 13635
rect 6303 13567 6304 13601
rect 6338 13567 6339 13601
rect 6303 13533 6339 13567
rect 6303 13499 6304 13533
rect 6338 13499 6339 13533
rect 6303 13465 6339 13499
rect 6303 13431 6304 13465
rect 6338 13431 6339 13465
rect 6303 13397 6339 13431
rect 6303 13363 6304 13397
rect 6338 13363 6339 13397
rect 6303 13329 6339 13363
rect 6303 13295 6304 13329
rect 6338 13295 6339 13329
rect 6303 13261 6339 13295
rect 6303 13227 6304 13261
rect 6338 13227 6339 13261
rect 6303 13193 6339 13227
rect 6303 13159 6304 13193
rect 6338 13159 6339 13193
rect 6303 13125 6339 13159
rect 6303 13091 6304 13125
rect 6338 13091 6339 13125
rect 6303 13057 6339 13091
rect 6303 13023 6304 13057
rect 6338 13023 6339 13057
rect 6303 12989 6339 13023
rect 6303 12955 6304 12989
rect 6338 12955 6339 12989
rect 6303 12921 6339 12955
rect 6303 12887 6304 12921
rect 6338 12887 6339 12921
rect 6303 12853 6339 12887
rect 6303 12819 6304 12853
rect 6338 12819 6339 12853
rect 6303 12785 6339 12819
rect 6303 12751 6304 12785
rect 6338 12751 6339 12785
rect 6303 12717 6339 12751
rect 6303 12683 6304 12717
rect 6338 12683 6339 12717
rect 6303 12649 6339 12683
rect 6303 12615 6304 12649
rect 6338 12615 6339 12649
rect 6303 12581 6339 12615
rect 6303 12547 6304 12581
rect 6338 12547 6339 12581
rect 6303 12513 6339 12547
rect 6303 12479 6304 12513
rect 6338 12479 6339 12513
rect 6303 12445 6339 12479
rect 6303 12411 6304 12445
rect 6338 12411 6339 12445
rect 6303 12377 6339 12411
rect 6303 12343 6304 12377
rect 6338 12343 6339 12377
rect 6303 12309 6339 12343
rect 6303 12275 6304 12309
rect 6338 12275 6339 12309
rect 6303 12241 6339 12275
rect 6303 12207 6304 12241
rect 6338 12207 6339 12241
rect 6303 12173 6339 12207
rect 6303 12139 6304 12173
rect 6338 12139 6339 12173
rect 6303 12105 6339 12139
rect 6303 12071 6304 12105
rect 6338 12071 6339 12105
rect 6303 12037 6339 12071
rect 6303 12003 6304 12037
rect 6338 12003 6339 12037
rect 6303 11969 6339 12003
rect 6303 11935 6304 11969
rect 6338 11935 6339 11969
rect 6303 11901 6339 11935
rect 6303 11867 6304 11901
rect 6338 11867 6339 11901
rect 6303 11833 6339 11867
rect 6303 11799 6304 11833
rect 6338 11799 6339 11833
rect 6303 11765 6339 11799
rect 6303 11731 6304 11765
rect 6338 11731 6339 11765
rect 6303 11697 6339 11731
rect 6303 11663 6304 11697
rect 6338 11663 6339 11697
rect 6303 11629 6339 11663
rect 6303 11595 6304 11629
rect 6338 11595 6339 11629
rect 6303 11561 6339 11595
rect 6303 11527 6304 11561
rect 6338 11527 6339 11561
rect 6303 11493 6339 11527
rect 6303 11459 6304 11493
rect 6338 11459 6339 11493
rect 6303 11425 6339 11459
rect 6303 11391 6304 11425
rect 6338 11391 6339 11425
rect 6303 11357 6339 11391
rect 6303 11323 6304 11357
rect 6338 11323 6339 11357
rect 6303 11289 6339 11323
rect 6303 11255 6304 11289
rect 6338 11255 6339 11289
rect 6303 11221 6339 11255
rect 6303 11187 6304 11221
rect 6338 11187 6339 11221
rect 6303 11153 6339 11187
rect 6303 11119 6304 11153
rect 6338 11119 6339 11153
rect 6303 11085 6339 11119
rect 6303 11051 6304 11085
rect 6338 11051 6339 11085
rect 6303 10972 6339 11051
rect 6303 10938 6304 10972
rect 6338 10938 6339 10972
rect 6303 10904 6339 10938
rect 6303 10870 6304 10904
rect 6338 10870 6339 10904
rect 6303 10836 6339 10870
rect 6303 10802 6304 10836
rect 6338 10802 6339 10836
rect 6303 10768 6339 10802
rect 6303 10734 6304 10768
rect 6338 10734 6339 10768
rect 6303 10700 6339 10734
rect 6303 10666 6304 10700
rect 6338 10666 6339 10700
rect 6303 10632 6339 10666
rect 6303 10598 6304 10632
rect 6338 10598 6339 10632
rect 6303 10564 6339 10598
rect 6303 10530 6304 10564
rect 6338 10530 6339 10564
rect 6303 10496 6339 10530
rect 6303 10462 6304 10496
rect 6338 10462 6339 10496
rect 6303 10428 6339 10462
rect 6303 10394 6304 10428
rect 6338 10394 6339 10428
rect 6303 10360 6339 10394
rect 6303 10326 6304 10360
rect 6338 10326 6339 10360
rect 6303 10292 6339 10326
rect 6303 10258 6304 10292
rect 6338 10258 6339 10292
rect 5059 10213 5095 10247
rect 5059 10179 5060 10213
rect 5094 10179 5095 10213
rect 6303 10224 6339 10258
rect 6303 10190 6304 10224
rect 6338 10190 6339 10224
rect 5059 10145 5095 10179
rect 5059 10111 5060 10145
rect 5094 10113 5095 10145
rect 6303 10113 6339 10190
rect 5094 10112 6339 10113
rect 5094 10111 5183 10112
rect 5059 10078 5183 10111
rect 5217 10078 5251 10112
rect 5285 10078 5319 10112
rect 5353 10078 5387 10112
rect 5421 10078 5455 10112
rect 5489 10078 5523 10112
rect 5557 10078 5591 10112
rect 5625 10078 5659 10112
rect 5693 10078 5727 10112
rect 5761 10078 5795 10112
rect 5829 10078 5863 10112
rect 5897 10078 5931 10112
rect 5965 10078 5999 10112
rect 6033 10078 6067 10112
rect 6101 10078 6135 10112
rect 6169 10078 6203 10112
rect 6237 10078 6271 10112
rect 6305 10078 6339 10112
rect 5059 10077 6339 10078
rect 539 9544 5865 9545
rect 539 9511 632 9544
rect 539 9477 540 9511
rect 574 9510 632 9511
rect 666 9510 700 9544
rect 734 9510 768 9544
rect 802 9510 836 9544
rect 870 9510 904 9544
rect 938 9510 972 9544
rect 1006 9510 1040 9544
rect 1074 9510 1108 9544
rect 1142 9510 1176 9544
rect 1210 9510 1244 9544
rect 1278 9510 1312 9544
rect 1346 9510 1380 9544
rect 1414 9510 1448 9544
rect 1482 9510 1516 9544
rect 1550 9510 1584 9544
rect 1618 9510 1652 9544
rect 1686 9510 1720 9544
rect 1754 9510 1788 9544
rect 1822 9510 1856 9544
rect 1890 9510 1924 9544
rect 1958 9510 1992 9544
rect 2026 9510 2060 9544
rect 2094 9510 2128 9544
rect 2162 9510 2196 9544
rect 2230 9510 2264 9544
rect 2298 9510 2332 9544
rect 2366 9510 2400 9544
rect 2434 9510 2468 9544
rect 2502 9510 2576 9544
rect 2610 9510 2644 9544
rect 2678 9510 2712 9544
rect 2746 9510 2780 9544
rect 2814 9510 2848 9544
rect 2882 9510 2916 9544
rect 2950 9510 2984 9544
rect 3018 9510 3052 9544
rect 3086 9510 3120 9544
rect 3154 9510 3188 9544
rect 3222 9510 3256 9544
rect 3290 9510 3324 9544
rect 3358 9510 3426 9544
rect 3460 9510 3494 9544
rect 3528 9510 3562 9544
rect 3596 9510 3630 9544
rect 3664 9510 3698 9544
rect 3732 9510 3766 9544
rect 3800 9510 3834 9544
rect 3868 9510 3902 9544
rect 3936 9510 3970 9544
rect 4004 9510 4038 9544
rect 4072 9510 4106 9544
rect 4140 9510 4174 9544
rect 4208 9510 4242 9544
rect 4276 9510 4310 9544
rect 4344 9510 4378 9544
rect 4412 9510 4446 9544
rect 4480 9510 4514 9544
rect 4548 9510 4582 9544
rect 4616 9510 4650 9544
rect 4684 9510 4718 9544
rect 4752 9510 4786 9544
rect 4820 9510 4854 9544
rect 4888 9510 4922 9544
rect 4956 9510 4990 9544
rect 5024 9510 5058 9544
rect 5092 9510 5126 9544
rect 5160 9510 5194 9544
rect 5228 9510 5262 9544
rect 5296 9510 5330 9544
rect 5364 9510 5398 9544
rect 5432 9510 5466 9544
rect 5500 9510 5534 9544
rect 5568 9510 5602 9544
rect 5636 9510 5670 9544
rect 5704 9510 5738 9544
rect 5772 9510 5865 9544
rect 574 9509 5865 9510
rect 574 9477 575 9509
rect 539 9443 575 9477
rect 539 9409 540 9443
rect 574 9409 575 9443
rect 539 9375 575 9409
rect 539 9341 540 9375
rect 574 9341 575 9375
rect 539 9307 575 9341
rect 539 9273 540 9307
rect 574 9273 575 9307
rect 539 9239 575 9273
rect 539 9205 540 9239
rect 574 9205 575 9239
rect 539 9171 575 9205
rect 539 9137 540 9171
rect 574 9137 575 9171
rect 539 9103 575 9137
rect 539 9069 540 9103
rect 574 9069 575 9103
rect 539 9035 575 9069
rect 539 9001 540 9035
rect 574 9001 575 9035
rect 539 8967 575 9001
rect 539 8933 540 8967
rect 574 8933 575 8967
rect 539 8899 575 8933
rect 539 8865 540 8899
rect 574 8865 575 8899
rect 539 8831 575 8865
rect 539 8797 540 8831
rect 574 8797 575 8831
rect 539 8763 575 8797
rect 539 8729 540 8763
rect 574 8729 575 8763
rect 539 8695 575 8729
rect 539 8661 540 8695
rect 574 8661 575 8695
rect 539 8627 575 8661
rect 539 8593 540 8627
rect 574 8593 575 8627
rect 539 8559 575 8593
rect 539 8525 540 8559
rect 574 8525 575 8559
rect 539 8491 575 8525
rect 539 8457 540 8491
rect 574 8457 575 8491
rect 539 8423 575 8457
rect 539 8389 540 8423
rect 574 8389 575 8423
rect 539 8355 575 8389
rect 539 8321 540 8355
rect 574 8321 575 8355
rect 539 8287 575 8321
rect 539 8253 540 8287
rect 574 8253 575 8287
rect 539 8219 575 8253
rect 539 8185 540 8219
rect 574 8185 575 8219
rect 539 8151 575 8185
rect 539 8117 540 8151
rect 574 8117 575 8151
rect 539 8083 575 8117
rect 539 8049 540 8083
rect 574 8049 575 8083
rect 539 8015 575 8049
rect 539 7981 540 8015
rect 574 7981 575 8015
rect 539 7947 575 7981
rect 539 7913 540 7947
rect 574 7913 575 7947
rect 539 7879 575 7913
rect 539 7845 540 7879
rect 574 7845 575 7879
rect 539 7811 575 7845
rect 539 7777 540 7811
rect 574 7777 575 7811
rect 539 7743 575 7777
rect 539 7709 540 7743
rect 574 7709 575 7743
rect 539 7675 575 7709
rect 539 7641 540 7675
rect 574 7641 575 7675
rect 539 7607 575 7641
rect 539 7573 540 7607
rect 574 7573 575 7607
rect 539 7539 575 7573
rect 539 7505 540 7539
rect 574 7505 575 7539
rect 539 7471 575 7505
rect 539 7437 540 7471
rect 574 7437 575 7471
rect 539 7403 575 7437
rect 539 7369 540 7403
rect 574 7369 575 7403
rect 539 7288 575 7369
rect 3356 9396 3392 9509
rect 5829 9475 5865 9509
rect 5829 9441 5830 9475
rect 5864 9441 5865 9475
rect 5829 9407 5865 9441
rect 3356 9362 3357 9396
rect 3391 9362 3392 9396
rect 3356 9328 3392 9362
rect 3356 9294 3357 9328
rect 3391 9294 3392 9328
rect 3356 9260 3392 9294
rect 3356 9226 3357 9260
rect 3391 9226 3392 9260
rect 3356 9192 3392 9226
rect 3356 9158 3357 9192
rect 3391 9158 3392 9192
rect 3356 9124 3392 9158
rect 3356 9090 3357 9124
rect 3391 9090 3392 9124
rect 3356 9056 3392 9090
rect 3356 9022 3357 9056
rect 3391 9022 3392 9056
rect 3356 8988 3392 9022
rect 3356 8954 3357 8988
rect 3391 8954 3392 8988
rect 3356 8920 3392 8954
rect 3356 8886 3357 8920
rect 3391 8886 3392 8920
rect 3356 8852 3392 8886
rect 3356 8818 3357 8852
rect 3391 8818 3392 8852
rect 3356 8784 3392 8818
rect 3356 8750 3357 8784
rect 3391 8750 3392 8784
rect 3356 8716 3392 8750
rect 3356 8682 3357 8716
rect 3391 8682 3392 8716
rect 3356 8648 3392 8682
rect 3356 8614 3357 8648
rect 3391 8614 3392 8648
rect 3356 8580 3392 8614
rect 3356 8546 3357 8580
rect 3391 8546 3392 8580
rect 3356 8512 3392 8546
rect 3356 8478 3357 8512
rect 3391 8478 3392 8512
rect 3356 8444 3392 8478
rect 3356 8410 3357 8444
rect 3391 8410 3392 8444
rect 3356 8376 3392 8410
rect 3356 8342 3357 8376
rect 3391 8342 3392 8376
rect 3356 8308 3392 8342
rect 3356 8274 3357 8308
rect 3391 8274 3392 8308
rect 3356 8240 3392 8274
rect 3356 8206 3357 8240
rect 3391 8206 3392 8240
rect 3356 8172 3392 8206
rect 3356 8138 3357 8172
rect 3391 8138 3392 8172
rect 3356 8104 3392 8138
rect 3356 8070 3357 8104
rect 3391 8070 3392 8104
rect 3356 8036 3392 8070
rect 3356 8002 3357 8036
rect 3391 8002 3392 8036
rect 3356 7968 3392 8002
rect 3356 7934 3357 7968
rect 3391 7934 3392 7968
rect 3356 7900 3392 7934
rect 3356 7866 3357 7900
rect 3391 7866 3392 7900
rect 3356 7832 3392 7866
rect 3356 7798 3357 7832
rect 3391 7798 3392 7832
rect 3356 7764 3392 7798
rect 3356 7730 3357 7764
rect 3391 7730 3392 7764
rect 3356 7696 3392 7730
rect 3356 7662 3357 7696
rect 3391 7662 3392 7696
rect 3356 7628 3392 7662
rect 3356 7594 3357 7628
rect 3391 7594 3392 7628
rect 3356 7560 3392 7594
rect 3356 7526 3357 7560
rect 3391 7526 3392 7560
rect 3356 7492 3392 7526
rect 3356 7458 3357 7492
rect 3391 7458 3392 7492
rect 3356 7424 3392 7458
rect 3356 7390 3357 7424
rect 3391 7390 3392 7424
rect 3356 7356 3392 7390
rect 3356 7322 3357 7356
rect 3391 7322 3392 7356
rect 5829 9373 5830 9407
rect 5864 9373 5865 9407
rect 5829 9339 5865 9373
rect 5829 9305 5830 9339
rect 5864 9305 5865 9339
rect 5829 9271 5865 9305
rect 5829 9237 5830 9271
rect 5864 9237 5865 9271
rect 5829 9203 5865 9237
rect 5829 9169 5830 9203
rect 5864 9169 5865 9203
rect 5829 9135 5865 9169
rect 5829 9101 5830 9135
rect 5864 9101 5865 9135
rect 5829 9067 5865 9101
rect 5829 9033 5830 9067
rect 5864 9033 5865 9067
rect 5829 8999 5865 9033
rect 5829 8965 5830 8999
rect 5864 8965 5865 8999
rect 5829 8931 5865 8965
rect 5829 8897 5830 8931
rect 5864 8897 5865 8931
rect 5829 8863 5865 8897
rect 5829 8829 5830 8863
rect 5864 8829 5865 8863
rect 5829 8795 5865 8829
rect 5829 8761 5830 8795
rect 5864 8761 5865 8795
rect 5829 8727 5865 8761
rect 5829 8693 5830 8727
rect 5864 8693 5865 8727
rect 5829 8659 5865 8693
rect 5829 8625 5830 8659
rect 5864 8625 5865 8659
rect 5829 8591 5865 8625
rect 5829 8557 5830 8591
rect 5864 8557 5865 8591
rect 5829 8523 5865 8557
rect 5829 8489 5830 8523
rect 5864 8489 5865 8523
rect 5829 8455 5865 8489
rect 5829 8421 5830 8455
rect 5864 8421 5865 8455
rect 5829 8387 5865 8421
rect 5829 8353 5830 8387
rect 5864 8353 5865 8387
rect 5829 8319 5865 8353
rect 5829 8285 5830 8319
rect 5864 8285 5865 8319
rect 5829 8251 5865 8285
rect 5829 8217 5830 8251
rect 5864 8217 5865 8251
rect 5829 8183 5865 8217
rect 5829 8149 5830 8183
rect 5864 8149 5865 8183
rect 5829 8115 5865 8149
rect 5829 8081 5830 8115
rect 5864 8081 5865 8115
rect 5829 8047 5865 8081
rect 5829 8013 5830 8047
rect 5864 8013 5865 8047
rect 5829 7979 5865 8013
rect 5829 7945 5830 7979
rect 5864 7945 5865 7979
rect 5829 7911 5865 7945
rect 5829 7877 5830 7911
rect 5864 7877 5865 7911
rect 5829 7843 5865 7877
rect 5829 7809 5830 7843
rect 5864 7809 5865 7843
rect 5829 7775 5865 7809
rect 5829 7741 5830 7775
rect 5864 7741 5865 7775
rect 5829 7707 5865 7741
rect 5829 7673 5830 7707
rect 5864 7673 5865 7707
rect 5829 7639 5865 7673
rect 5829 7605 5830 7639
rect 5864 7605 5865 7639
rect 5829 7571 5865 7605
rect 5829 7537 5830 7571
rect 5864 7537 5865 7571
rect 5829 7503 5865 7537
rect 5829 7469 5830 7503
rect 5864 7469 5865 7503
rect 5829 7435 5865 7469
rect 5829 7401 5830 7435
rect 5864 7401 5865 7435
rect 5829 7367 5865 7401
rect 539 7287 967 7288
rect 539 7253 657 7287
rect 691 7253 741 7287
rect 775 7253 825 7287
rect 859 7253 909 7287
rect 943 7253 967 7287
rect 539 7252 967 7253
rect 1237 7287 1823 7288
rect 1237 7253 1261 7287
rect 1295 7253 1345 7287
rect 1379 7253 1429 7287
rect 1463 7253 1513 7287
rect 1547 7253 1597 7287
rect 1631 7253 1681 7287
rect 1715 7253 1765 7287
rect 1799 7253 1823 7287
rect 1237 7252 1823 7253
rect 2093 7287 2679 7288
rect 2093 7253 2117 7287
rect 2151 7253 2201 7287
rect 2235 7253 2285 7287
rect 2319 7253 2369 7287
rect 2403 7253 2453 7287
rect 2487 7253 2537 7287
rect 2571 7253 2621 7287
rect 2655 7253 2679 7287
rect 2093 7252 2679 7253
rect 3356 7288 3392 7322
rect 5829 7333 5830 7367
rect 5864 7333 5865 7367
rect 2949 7287 3357 7288
rect 2949 7253 2973 7287
rect 3007 7253 3057 7287
rect 3091 7253 3141 7287
rect 3175 7253 3225 7287
rect 3259 7254 3357 7287
rect 3391 7287 3799 7288
rect 3391 7254 3489 7287
rect 3259 7253 3489 7254
rect 3523 7253 3573 7287
rect 3607 7253 3657 7287
rect 3691 7253 3741 7287
rect 3775 7253 3799 7287
rect 2949 7252 3799 7253
rect 4069 7287 4455 7288
rect 4069 7253 4093 7287
rect 4127 7253 4177 7287
rect 4211 7253 4261 7287
rect 4295 7253 4345 7287
rect 4379 7253 4455 7287
rect 4069 7252 4455 7253
rect 4725 7287 4911 7288
rect 4725 7253 4801 7287
rect 4835 7253 4911 7287
rect 4725 7252 4911 7253
rect 5181 7287 5367 7288
rect 5181 7253 5257 7287
rect 5291 7253 5367 7287
rect 5181 7252 5367 7253
rect 5829 7299 5865 7333
rect 5829 7288 5830 7299
rect 5637 7287 5830 7288
rect 5637 7253 5713 7287
rect 5747 7265 5830 7287
rect 5864 7265 5865 7299
rect 5747 7253 5865 7265
rect 5637 7252 5865 7253
rect 539 7251 575 7252
rect 539 7217 540 7251
rect 574 7217 575 7251
rect 539 7183 575 7217
rect 3356 7220 3392 7252
rect 539 7149 540 7183
rect 574 7149 575 7183
rect 539 7115 575 7149
rect 539 7081 540 7115
rect 574 7081 575 7115
rect 539 7047 575 7081
rect 539 7013 540 7047
rect 574 7013 575 7047
rect 539 6979 575 7013
rect 539 6945 540 6979
rect 574 6945 575 6979
rect 539 6911 575 6945
rect 539 6877 540 6911
rect 574 6877 575 6911
rect 539 6843 575 6877
rect 539 6809 540 6843
rect 574 6809 575 6843
rect 539 6775 575 6809
rect 539 6741 540 6775
rect 574 6741 575 6775
rect 539 6707 575 6741
rect 539 6673 540 6707
rect 574 6673 575 6707
rect 539 6639 575 6673
rect 539 6605 540 6639
rect 574 6605 575 6639
rect 539 6571 575 6605
rect 539 6537 540 6571
rect 574 6537 575 6571
rect 539 6503 575 6537
rect 539 6469 540 6503
rect 574 6469 575 6503
rect 539 6435 575 6469
rect 539 6401 540 6435
rect 574 6401 575 6435
rect 539 6367 575 6401
rect 539 6333 540 6367
rect 574 6333 575 6367
rect 539 6299 575 6333
rect 539 6265 540 6299
rect 574 6265 575 6299
rect 539 6231 575 6265
rect 539 6197 540 6231
rect 574 6197 575 6231
rect 539 6163 575 6197
rect 539 6129 540 6163
rect 574 6129 575 6163
rect 539 6095 575 6129
rect 539 6061 540 6095
rect 574 6061 575 6095
rect 539 6027 575 6061
rect 539 5993 540 6027
rect 574 5993 575 6027
rect 539 5959 575 5993
rect 539 5925 540 5959
rect 574 5925 575 5959
rect 539 5891 575 5925
rect 539 5857 540 5891
rect 574 5857 575 5891
rect 539 5823 575 5857
rect 539 5789 540 5823
rect 574 5789 575 5823
rect 539 5755 575 5789
rect 539 5721 540 5755
rect 574 5721 575 5755
rect 539 5687 575 5721
rect 539 5653 540 5687
rect 574 5653 575 5687
rect 539 5619 575 5653
rect 539 5585 540 5619
rect 574 5585 575 5619
rect 539 5551 575 5585
rect 539 5517 540 5551
rect 574 5517 575 5551
rect 539 5483 575 5517
rect 539 5449 540 5483
rect 574 5449 575 5483
rect 539 5415 575 5449
rect 539 5381 540 5415
rect 574 5381 575 5415
rect 539 5347 575 5381
rect 539 5313 540 5347
rect 574 5313 575 5347
rect 539 5279 575 5313
rect 539 5245 540 5279
rect 574 5245 575 5279
rect 539 5211 575 5245
rect 539 5177 540 5211
rect 574 5177 575 5211
rect 539 5068 575 5177
rect 3356 7186 3357 7220
rect 3391 7186 3392 7220
rect 5829 7231 5865 7252
rect 5829 7197 5830 7231
rect 5864 7197 5865 7231
rect 3356 7152 3392 7186
rect 3356 7118 3357 7152
rect 3391 7118 3392 7152
rect 3356 7084 3392 7118
rect 3356 7050 3357 7084
rect 3391 7050 3392 7084
rect 3356 7016 3392 7050
rect 3356 6982 3357 7016
rect 3391 6982 3392 7016
rect 3356 6948 3392 6982
rect 3356 6914 3357 6948
rect 3391 6914 3392 6948
rect 3356 6880 3392 6914
rect 3356 6846 3357 6880
rect 3391 6846 3392 6880
rect 3356 6812 3392 6846
rect 3356 6778 3357 6812
rect 3391 6778 3392 6812
rect 3356 6744 3392 6778
rect 3356 6710 3357 6744
rect 3391 6710 3392 6744
rect 3356 6676 3392 6710
rect 3356 6642 3357 6676
rect 3391 6642 3392 6676
rect 3356 6608 3392 6642
rect 3356 6574 3357 6608
rect 3391 6574 3392 6608
rect 3356 6540 3392 6574
rect 3356 6506 3357 6540
rect 3391 6506 3392 6540
rect 3356 6472 3392 6506
rect 3356 6438 3357 6472
rect 3391 6438 3392 6472
rect 3356 6404 3392 6438
rect 3356 6370 3357 6404
rect 3391 6370 3392 6404
rect 3356 6336 3392 6370
rect 3356 6302 3357 6336
rect 3391 6302 3392 6336
rect 3356 6268 3392 6302
rect 3356 6234 3357 6268
rect 3391 6234 3392 6268
rect 3356 6200 3392 6234
rect 3356 6166 3357 6200
rect 3391 6166 3392 6200
rect 3356 6132 3392 6166
rect 3356 6098 3357 6132
rect 3391 6098 3392 6132
rect 3356 6064 3392 6098
rect 3356 6030 3357 6064
rect 3391 6030 3392 6064
rect 3356 5996 3392 6030
rect 3356 5962 3357 5996
rect 3391 5962 3392 5996
rect 3356 5928 3392 5962
rect 3356 5894 3357 5928
rect 3391 5894 3392 5928
rect 3356 5860 3392 5894
rect 3356 5826 3357 5860
rect 3391 5826 3392 5860
rect 3356 5792 3392 5826
rect 3356 5758 3357 5792
rect 3391 5758 3392 5792
rect 3356 5724 3392 5758
rect 3356 5690 3357 5724
rect 3391 5690 3392 5724
rect 3356 5656 3392 5690
rect 3356 5622 3357 5656
rect 3391 5622 3392 5656
rect 3356 5588 3392 5622
rect 3356 5554 3357 5588
rect 3391 5554 3392 5588
rect 3356 5520 3392 5554
rect 3356 5486 3357 5520
rect 3391 5486 3392 5520
rect 3356 5452 3392 5486
rect 3356 5418 3357 5452
rect 3391 5418 3392 5452
rect 3356 5384 3392 5418
rect 3356 5350 3357 5384
rect 3391 5350 3392 5384
rect 3356 5316 3392 5350
rect 3356 5282 3357 5316
rect 3391 5282 3392 5316
rect 3356 5248 3392 5282
rect 3356 5214 3357 5248
rect 3391 5214 3392 5248
rect 3356 5180 3392 5214
rect 3356 5146 3357 5180
rect 3391 5146 3392 5180
rect 3356 5112 3392 5146
rect 5829 7163 5865 7197
rect 5829 7129 5830 7163
rect 5864 7129 5865 7163
rect 5829 7095 5865 7129
rect 5829 7061 5830 7095
rect 5864 7061 5865 7095
rect 5829 7027 5865 7061
rect 5829 6993 5830 7027
rect 5864 6993 5865 7027
rect 5829 6959 5865 6993
rect 5829 6925 5830 6959
rect 5864 6925 5865 6959
rect 5829 6891 5865 6925
rect 5829 6857 5830 6891
rect 5864 6857 5865 6891
rect 5829 6823 5865 6857
rect 5829 6789 5830 6823
rect 5864 6789 5865 6823
rect 5829 6755 5865 6789
rect 5829 6721 5830 6755
rect 5864 6721 5865 6755
rect 5829 6687 5865 6721
rect 5829 6653 5830 6687
rect 5864 6653 5865 6687
rect 5829 6619 5865 6653
rect 5829 6585 5830 6619
rect 5864 6585 5865 6619
rect 5829 6551 5865 6585
rect 5829 6517 5830 6551
rect 5864 6517 5865 6551
rect 5829 6483 5865 6517
rect 5829 6449 5830 6483
rect 5864 6449 5865 6483
rect 5829 6415 5865 6449
rect 5829 6381 5830 6415
rect 5864 6381 5865 6415
rect 5829 6347 5865 6381
rect 5829 6313 5830 6347
rect 5864 6313 5865 6347
rect 5829 6279 5865 6313
rect 5829 6245 5830 6279
rect 5864 6245 5865 6279
rect 5829 6211 5865 6245
rect 5829 6177 5830 6211
rect 5864 6177 5865 6211
rect 5829 6143 5865 6177
rect 5829 6109 5830 6143
rect 5864 6109 5865 6143
rect 5829 6075 5865 6109
rect 5829 6041 5830 6075
rect 5864 6041 5865 6075
rect 5829 6007 5865 6041
rect 5829 5973 5830 6007
rect 5864 5973 5865 6007
rect 5829 5939 5865 5973
rect 5829 5905 5830 5939
rect 5864 5905 5865 5939
rect 5829 5871 5865 5905
rect 5829 5837 5830 5871
rect 5864 5837 5865 5871
rect 5829 5803 5865 5837
rect 5829 5769 5830 5803
rect 5864 5769 5865 5803
rect 5829 5735 5865 5769
rect 5829 5701 5830 5735
rect 5864 5701 5865 5735
rect 5829 5667 5865 5701
rect 5829 5633 5830 5667
rect 5864 5633 5865 5667
rect 5829 5599 5865 5633
rect 5829 5565 5830 5599
rect 5864 5565 5865 5599
rect 5829 5531 5865 5565
rect 5829 5497 5830 5531
rect 5864 5497 5865 5531
rect 5829 5463 5865 5497
rect 5829 5429 5830 5463
rect 5864 5429 5865 5463
rect 5829 5395 5865 5429
rect 5829 5361 5830 5395
rect 5864 5361 5865 5395
rect 5829 5327 5865 5361
rect 5829 5293 5830 5327
rect 5864 5293 5865 5327
rect 5829 5259 5865 5293
rect 5829 5225 5830 5259
rect 5864 5225 5865 5259
rect 5829 5191 5865 5225
rect 5829 5157 5830 5191
rect 5864 5157 5865 5191
rect 539 5067 967 5068
rect 539 5048 657 5067
rect 539 5014 540 5048
rect 574 5033 657 5048
rect 691 5033 741 5067
rect 775 5033 825 5067
rect 859 5033 909 5067
rect 943 5033 967 5067
rect 574 5032 967 5033
rect 1237 5067 1823 5068
rect 1237 5033 1261 5067
rect 1295 5033 1345 5067
rect 1379 5033 1429 5067
rect 1463 5033 1513 5067
rect 1547 5033 1597 5067
rect 1631 5033 1681 5067
rect 1715 5033 1765 5067
rect 1799 5033 1823 5067
rect 1237 5032 1823 5033
rect 2093 5067 2679 5068
rect 2093 5033 2117 5067
rect 2151 5033 2201 5067
rect 2235 5033 2285 5067
rect 2319 5033 2369 5067
rect 2403 5033 2453 5067
rect 2487 5033 2537 5067
rect 2571 5033 2621 5067
rect 2655 5033 2679 5067
rect 2093 5032 2679 5033
rect 3356 5078 3357 5112
rect 3391 5078 3392 5112
rect 5829 5123 5865 5157
rect 5829 5089 5830 5123
rect 5864 5089 5865 5123
rect 3356 5068 3392 5078
rect 2949 5067 3799 5068
rect 2949 5033 2973 5067
rect 3007 5033 3057 5067
rect 3091 5033 3141 5067
rect 3175 5033 3225 5067
rect 3259 5044 3489 5067
rect 3259 5033 3357 5044
rect 2949 5032 3357 5033
rect 574 5014 575 5032
rect 539 4980 575 5014
rect 539 4946 540 4980
rect 574 4946 575 4980
rect 3356 5010 3357 5032
rect 3391 5033 3489 5044
rect 3523 5033 3573 5067
rect 3607 5033 3657 5067
rect 3691 5033 3741 5067
rect 3775 5033 3799 5067
rect 3391 5032 3799 5033
rect 4069 5067 4455 5068
rect 4069 5033 4093 5067
rect 4127 5033 4177 5067
rect 4211 5033 4261 5067
rect 4295 5033 4345 5067
rect 4379 5033 4455 5067
rect 4069 5032 4455 5033
rect 4725 5067 4911 5068
rect 4725 5033 4801 5067
rect 4835 5033 4911 5067
rect 4725 5032 4911 5033
rect 5181 5067 5367 5068
rect 5181 5033 5257 5067
rect 5291 5033 5367 5067
rect 5181 5032 5367 5033
rect 5829 5068 5865 5089
rect 5637 5067 5865 5068
rect 5637 5033 5713 5067
rect 5747 5055 5865 5067
rect 5747 5033 5830 5055
rect 5637 5032 5830 5033
rect 3391 5010 3392 5032
rect 5829 5021 5830 5032
rect 5864 5021 5865 5055
rect 3356 4976 3392 5010
rect 539 4912 575 4946
rect 539 4878 540 4912
rect 574 4878 575 4912
rect 539 4844 575 4878
rect 539 4810 540 4844
rect 574 4810 575 4844
rect 539 4776 575 4810
rect 539 4742 540 4776
rect 574 4742 575 4776
rect 539 4708 575 4742
rect 539 4674 540 4708
rect 574 4674 575 4708
rect 539 4640 575 4674
rect 539 4606 540 4640
rect 574 4606 575 4640
rect 539 4572 575 4606
rect 539 4538 540 4572
rect 574 4538 575 4572
rect 539 4504 575 4538
rect 539 4470 540 4504
rect 574 4470 575 4504
rect 539 4436 575 4470
rect 539 4402 540 4436
rect 574 4402 575 4436
rect 539 4368 575 4402
rect 539 4334 540 4368
rect 574 4334 575 4368
rect 539 4300 575 4334
rect 539 4266 540 4300
rect 574 4266 575 4300
rect 539 4232 575 4266
rect 539 4198 540 4232
rect 574 4198 575 4232
rect 539 4164 575 4198
rect 539 4130 540 4164
rect 574 4130 575 4164
rect 539 4096 575 4130
rect 539 4062 540 4096
rect 574 4062 575 4096
rect 539 4028 575 4062
rect 539 3994 540 4028
rect 574 3994 575 4028
rect 539 3960 575 3994
rect 539 3926 540 3960
rect 574 3926 575 3960
rect 539 3892 575 3926
rect 539 3858 540 3892
rect 574 3858 575 3892
rect 539 3824 575 3858
rect 539 3790 540 3824
rect 574 3790 575 3824
rect 539 3756 575 3790
rect 539 3722 540 3756
rect 574 3722 575 3756
rect 539 3688 575 3722
rect 539 3654 540 3688
rect 574 3654 575 3688
rect 539 3620 575 3654
rect 539 3586 540 3620
rect 574 3586 575 3620
rect 539 3552 575 3586
rect 539 3518 540 3552
rect 574 3518 575 3552
rect 539 3484 575 3518
rect 539 3450 540 3484
rect 574 3450 575 3484
rect 539 3416 575 3450
rect 539 3382 540 3416
rect 574 3382 575 3416
rect 539 3348 575 3382
rect 539 3314 540 3348
rect 574 3314 575 3348
rect 539 3280 575 3314
rect 539 3246 540 3280
rect 574 3246 575 3280
rect 539 3212 575 3246
rect 539 3178 540 3212
rect 574 3178 575 3212
rect 539 3144 575 3178
rect 539 3110 540 3144
rect 574 3110 575 3144
rect 539 3076 575 3110
rect 539 3042 540 3076
rect 574 3042 575 3076
rect 539 3008 575 3042
rect 539 2974 540 3008
rect 574 2974 575 3008
rect 539 2940 575 2974
rect 539 2906 540 2940
rect 574 2906 575 2940
rect 3356 4942 3357 4976
rect 3391 4942 3392 4976
rect 5829 4987 5865 5021
rect 3356 4908 3392 4942
rect 3356 4874 3357 4908
rect 3391 4874 3392 4908
rect 3356 4840 3392 4874
rect 3356 4806 3357 4840
rect 3391 4806 3392 4840
rect 3356 4772 3392 4806
rect 3356 4738 3357 4772
rect 3391 4738 3392 4772
rect 3356 4704 3392 4738
rect 3356 4670 3357 4704
rect 3391 4670 3392 4704
rect 3356 4636 3392 4670
rect 3356 4602 3357 4636
rect 3391 4602 3392 4636
rect 3356 4568 3392 4602
rect 3356 4534 3357 4568
rect 3391 4534 3392 4568
rect 3356 4500 3392 4534
rect 3356 4466 3357 4500
rect 3391 4466 3392 4500
rect 3356 4432 3392 4466
rect 3356 4398 3357 4432
rect 3391 4398 3392 4432
rect 3356 4364 3392 4398
rect 3356 4330 3357 4364
rect 3391 4330 3392 4364
rect 3356 4296 3392 4330
rect 3356 4262 3357 4296
rect 3391 4262 3392 4296
rect 3356 4228 3392 4262
rect 3356 4194 3357 4228
rect 3391 4194 3392 4228
rect 3356 4160 3392 4194
rect 3356 4126 3357 4160
rect 3391 4126 3392 4160
rect 3356 4092 3392 4126
rect 3356 4058 3357 4092
rect 3391 4058 3392 4092
rect 3356 4024 3392 4058
rect 3356 3990 3357 4024
rect 3391 3990 3392 4024
rect 3356 3956 3392 3990
rect 3356 3922 3357 3956
rect 3391 3922 3392 3956
rect 3356 3888 3392 3922
rect 3356 3854 3357 3888
rect 3391 3854 3392 3888
rect 3356 3820 3392 3854
rect 3356 3786 3357 3820
rect 3391 3786 3392 3820
rect 3356 3752 3392 3786
rect 3356 3718 3357 3752
rect 3391 3718 3392 3752
rect 3356 3684 3392 3718
rect 3356 3650 3357 3684
rect 3391 3650 3392 3684
rect 3356 3616 3392 3650
rect 3356 3582 3357 3616
rect 3391 3582 3392 3616
rect 3356 3548 3392 3582
rect 3356 3514 3357 3548
rect 3391 3514 3392 3548
rect 3356 3480 3392 3514
rect 3356 3446 3357 3480
rect 3391 3446 3392 3480
rect 3356 3412 3392 3446
rect 3356 3378 3357 3412
rect 3391 3378 3392 3412
rect 3356 3344 3392 3378
rect 3356 3310 3357 3344
rect 3391 3310 3392 3344
rect 3356 3276 3392 3310
rect 3356 3242 3357 3276
rect 3391 3242 3392 3276
rect 3356 3208 3392 3242
rect 3356 3174 3357 3208
rect 3391 3174 3392 3208
rect 3356 3140 3392 3174
rect 3356 3106 3357 3140
rect 3391 3106 3392 3140
rect 3356 3072 3392 3106
rect 3356 3038 3357 3072
rect 3391 3038 3392 3072
rect 3356 3004 3392 3038
rect 3356 2970 3357 3004
rect 3391 2970 3392 3004
rect 3356 2936 3392 2970
rect 539 2872 575 2906
rect 539 2838 540 2872
rect 574 2849 575 2872
rect 3356 2902 3357 2936
rect 3391 2902 3392 2936
rect 5829 4953 5830 4987
rect 5864 4953 5865 4987
rect 5829 4919 5865 4953
rect 5829 4885 5830 4919
rect 5864 4885 5865 4919
rect 5829 4851 5865 4885
rect 5829 4817 5830 4851
rect 5864 4817 5865 4851
rect 5829 4783 5865 4817
rect 5829 4749 5830 4783
rect 5864 4749 5865 4783
rect 5829 4715 5865 4749
rect 5829 4681 5830 4715
rect 5864 4681 5865 4715
rect 5829 4647 5865 4681
rect 5829 4613 5830 4647
rect 5864 4613 5865 4647
rect 5829 4579 5865 4613
rect 5829 4545 5830 4579
rect 5864 4545 5865 4579
rect 5829 4511 5865 4545
rect 5829 4477 5830 4511
rect 5864 4477 5865 4511
rect 5829 4443 5865 4477
rect 5829 4409 5830 4443
rect 5864 4409 5865 4443
rect 5829 4375 5865 4409
rect 5829 4341 5830 4375
rect 5864 4341 5865 4375
rect 5829 4307 5865 4341
rect 5829 4273 5830 4307
rect 5864 4273 5865 4307
rect 5829 4239 5865 4273
rect 5829 4205 5830 4239
rect 5864 4205 5865 4239
rect 5829 4171 5865 4205
rect 5829 4137 5830 4171
rect 5864 4137 5865 4171
rect 5829 4103 5865 4137
rect 5829 4069 5830 4103
rect 5864 4069 5865 4103
rect 5829 4035 5865 4069
rect 5829 4001 5830 4035
rect 5864 4001 5865 4035
rect 5829 3967 5865 4001
rect 5829 3933 5830 3967
rect 5864 3933 5865 3967
rect 5829 3899 5865 3933
rect 5829 3865 5830 3899
rect 5864 3865 5865 3899
rect 5829 3831 5865 3865
rect 5829 3797 5830 3831
rect 5864 3797 5865 3831
rect 5829 3763 5865 3797
rect 5829 3729 5830 3763
rect 5864 3729 5865 3763
rect 5829 3695 5865 3729
rect 5829 3661 5830 3695
rect 5864 3661 5865 3695
rect 5829 3627 5865 3661
rect 5829 3593 5830 3627
rect 5864 3593 5865 3627
rect 5829 3559 5865 3593
rect 5829 3525 5830 3559
rect 5864 3525 5865 3559
rect 5829 3491 5865 3525
rect 5829 3457 5830 3491
rect 5864 3457 5865 3491
rect 5829 3423 5865 3457
rect 5829 3389 5830 3423
rect 5864 3389 5865 3423
rect 5829 3355 5865 3389
rect 5829 3321 5830 3355
rect 5864 3321 5865 3355
rect 5829 3287 5865 3321
rect 5829 3253 5830 3287
rect 5864 3253 5865 3287
rect 5829 3219 5865 3253
rect 5829 3185 5830 3219
rect 5864 3185 5865 3219
rect 5829 3151 5865 3185
rect 5829 3117 5830 3151
rect 5864 3117 5865 3151
rect 5829 3083 5865 3117
rect 5829 3049 5830 3083
rect 5864 3049 5865 3083
rect 5829 3015 5865 3049
rect 5829 2981 5830 3015
rect 5864 2981 5865 3015
rect 5829 2947 5865 2981
rect 5829 2913 5830 2947
rect 5864 2913 5865 2947
rect 574 2848 967 2849
rect 574 2838 657 2848
rect 539 2814 657 2838
rect 691 2814 741 2848
rect 775 2814 825 2848
rect 859 2814 909 2848
rect 943 2814 967 2848
rect 539 2813 967 2814
rect 1237 2848 1823 2849
rect 1237 2814 1261 2848
rect 1295 2814 1345 2848
rect 1379 2814 1429 2848
rect 1463 2814 1513 2848
rect 1547 2814 1597 2848
rect 1631 2814 1681 2848
rect 1715 2814 1765 2848
rect 1799 2814 1823 2848
rect 1237 2813 1823 2814
rect 2093 2848 2679 2849
rect 2093 2814 2117 2848
rect 2151 2814 2201 2848
rect 2235 2814 2285 2848
rect 2319 2814 2369 2848
rect 2403 2814 2453 2848
rect 2487 2814 2537 2848
rect 2571 2814 2621 2848
rect 2655 2814 2679 2848
rect 2093 2813 2679 2814
rect 3356 2868 3392 2902
rect 5829 2879 5865 2913
rect 3356 2849 3357 2868
rect 2949 2848 3357 2849
rect 2949 2814 2973 2848
rect 3007 2814 3057 2848
rect 3091 2814 3141 2848
rect 3175 2814 3225 2848
rect 3259 2834 3357 2848
rect 3391 2849 3392 2868
rect 3391 2848 3799 2849
rect 3391 2834 3489 2848
rect 3259 2814 3489 2834
rect 3523 2814 3573 2848
rect 3607 2814 3657 2848
rect 3691 2814 3741 2848
rect 3775 2814 3799 2848
rect 2949 2813 3799 2814
rect 4069 2848 4455 2849
rect 4069 2814 4093 2848
rect 4127 2814 4177 2848
rect 4211 2814 4261 2848
rect 4295 2814 4345 2848
rect 4379 2814 4455 2848
rect 4069 2813 4455 2814
rect 4725 2848 4911 2849
rect 4725 2814 4801 2848
rect 4835 2814 4911 2848
rect 4725 2813 4911 2814
rect 5181 2848 5367 2849
rect 5181 2814 5257 2848
rect 5291 2814 5367 2848
rect 5181 2813 5367 2814
rect 5829 2849 5830 2879
rect 5637 2848 5830 2849
rect 5637 2814 5713 2848
rect 5747 2845 5830 2848
rect 5864 2845 5865 2879
rect 5747 2814 5865 2845
rect 5637 2813 5865 2814
rect 539 2804 575 2813
rect 539 2770 540 2804
rect 574 2770 575 2804
rect 3356 2800 3392 2813
rect 539 2736 575 2770
rect 3356 2766 3357 2800
rect 3391 2766 3392 2800
rect 5829 2811 5865 2813
rect 539 2702 540 2736
rect 574 2702 575 2736
rect 539 2584 575 2702
rect 539 2550 540 2584
rect 574 2550 575 2584
rect 539 2516 575 2550
rect 539 2482 540 2516
rect 574 2482 575 2516
rect 539 2448 575 2482
rect 539 2414 540 2448
rect 574 2414 575 2448
rect 539 2380 575 2414
rect 539 2346 540 2380
rect 574 2346 575 2380
rect 539 2312 575 2346
rect 539 2278 540 2312
rect 574 2278 575 2312
rect 539 2244 575 2278
rect 539 2210 540 2244
rect 574 2210 575 2244
rect 539 2176 575 2210
rect 539 2142 540 2176
rect 574 2142 575 2176
rect 539 2108 575 2142
rect 539 2074 540 2108
rect 574 2074 575 2108
rect 539 2040 575 2074
rect 539 2006 540 2040
rect 574 2006 575 2040
rect 539 1972 575 2006
rect 539 1938 540 1972
rect 574 1938 575 1972
rect 539 1904 575 1938
rect 539 1870 540 1904
rect 574 1870 575 1904
rect 539 1836 575 1870
rect 539 1802 540 1836
rect 574 1802 575 1836
rect 539 1768 575 1802
rect 539 1734 540 1768
rect 574 1734 575 1768
rect 539 1700 575 1734
rect 539 1666 540 1700
rect 574 1666 575 1700
rect 539 1632 575 1666
rect 539 1598 540 1632
rect 574 1598 575 1632
rect 539 1564 575 1598
rect 539 1530 540 1564
rect 574 1530 575 1564
rect 539 1496 575 1530
rect 539 1462 540 1496
rect 574 1462 575 1496
rect 539 1428 575 1462
rect 539 1394 540 1428
rect 574 1394 575 1428
rect 539 1360 575 1394
rect 539 1326 540 1360
rect 574 1326 575 1360
rect 539 1292 575 1326
rect 539 1258 540 1292
rect 574 1258 575 1292
rect 539 1224 575 1258
rect 539 1190 540 1224
rect 574 1190 575 1224
rect 539 1156 575 1190
rect 539 1122 540 1156
rect 574 1122 575 1156
rect 539 1088 575 1122
rect 539 1054 540 1088
rect 574 1054 575 1088
rect 539 1020 575 1054
rect 539 986 540 1020
rect 574 986 575 1020
rect 539 952 575 986
rect 539 918 540 952
rect 574 918 575 952
rect 539 884 575 918
rect 539 850 540 884
rect 574 850 575 884
rect 539 816 575 850
rect 539 782 540 816
rect 574 782 575 816
rect 539 748 575 782
rect 539 714 540 748
rect 574 714 575 748
rect 539 592 575 714
rect 3356 2732 3392 2766
rect 5829 2777 5830 2811
rect 5864 2777 5865 2811
rect 3356 2698 3357 2732
rect 3391 2698 3392 2732
rect 3356 2664 3392 2698
rect 3356 2630 3357 2664
rect 3391 2630 3392 2664
rect 3356 2596 3392 2630
rect 3356 2562 3357 2596
rect 3391 2562 3392 2596
rect 3356 2528 3392 2562
rect 3356 2494 3357 2528
rect 3391 2494 3392 2528
rect 3356 2460 3392 2494
rect 3356 2426 3357 2460
rect 3391 2426 3392 2460
rect 3356 2392 3392 2426
rect 3356 2358 3357 2392
rect 3391 2358 3392 2392
rect 3356 2324 3392 2358
rect 3356 2290 3357 2324
rect 3391 2290 3392 2324
rect 3356 2256 3392 2290
rect 3356 2222 3357 2256
rect 3391 2222 3392 2256
rect 3356 2188 3392 2222
rect 3356 2154 3357 2188
rect 3391 2154 3392 2188
rect 3356 2120 3392 2154
rect 3356 2086 3357 2120
rect 3391 2086 3392 2120
rect 3356 2052 3392 2086
rect 3356 2018 3357 2052
rect 3391 2018 3392 2052
rect 3356 1984 3392 2018
rect 3356 1950 3357 1984
rect 3391 1950 3392 1984
rect 3356 1916 3392 1950
rect 3356 1882 3357 1916
rect 3391 1882 3392 1916
rect 3356 1848 3392 1882
rect 3356 1814 3357 1848
rect 3391 1814 3392 1848
rect 3356 1780 3392 1814
rect 3356 1746 3357 1780
rect 3391 1746 3392 1780
rect 3356 1712 3392 1746
rect 3356 1678 3357 1712
rect 3391 1678 3392 1712
rect 3356 1644 3392 1678
rect 3356 1610 3357 1644
rect 3391 1610 3392 1644
rect 3356 1576 3392 1610
rect 3356 1542 3357 1576
rect 3391 1542 3392 1576
rect 3356 1508 3392 1542
rect 3356 1474 3357 1508
rect 3391 1474 3392 1508
rect 3356 1440 3392 1474
rect 3356 1406 3357 1440
rect 3391 1406 3392 1440
rect 3356 1372 3392 1406
rect 3356 1338 3357 1372
rect 3391 1338 3392 1372
rect 3356 1304 3392 1338
rect 3356 1270 3357 1304
rect 3391 1270 3392 1304
rect 3356 1236 3392 1270
rect 3356 1202 3357 1236
rect 3391 1202 3392 1236
rect 3356 1168 3392 1202
rect 3356 1134 3357 1168
rect 3391 1134 3392 1168
rect 3356 1100 3392 1134
rect 3356 1066 3357 1100
rect 3391 1066 3392 1100
rect 3356 1032 3392 1066
rect 3356 998 3357 1032
rect 3391 998 3392 1032
rect 3356 964 3392 998
rect 3356 930 3357 964
rect 3391 930 3392 964
rect 3356 896 3392 930
rect 3356 862 3357 896
rect 3391 862 3392 896
rect 3356 828 3392 862
rect 3356 794 3357 828
rect 3391 794 3392 828
rect 3356 760 3392 794
rect 3356 726 3357 760
rect 3391 726 3392 760
rect 3356 692 3392 726
rect 5829 2743 5865 2777
rect 5829 2709 5830 2743
rect 5864 2709 5865 2743
rect 5829 2675 5865 2709
rect 5829 2641 5830 2675
rect 5864 2641 5865 2675
rect 5829 2607 5865 2641
rect 5829 2573 5830 2607
rect 5864 2573 5865 2607
rect 5829 2539 5865 2573
rect 5829 2505 5830 2539
rect 5864 2505 5865 2539
rect 5829 2471 5865 2505
rect 5829 2437 5830 2471
rect 5864 2437 5865 2471
rect 5829 2403 5865 2437
rect 5829 2369 5830 2403
rect 5864 2369 5865 2403
rect 5829 2335 5865 2369
rect 5829 2301 5830 2335
rect 5864 2301 5865 2335
rect 5829 2267 5865 2301
rect 5829 2233 5830 2267
rect 5864 2233 5865 2267
rect 5829 2199 5865 2233
rect 5829 2165 5830 2199
rect 5864 2165 5865 2199
rect 5829 2131 5865 2165
rect 5829 2097 5830 2131
rect 5864 2097 5865 2131
rect 5829 2063 5865 2097
rect 5829 2029 5830 2063
rect 5864 2029 5865 2063
rect 5829 1995 5865 2029
rect 5829 1961 5830 1995
rect 5864 1961 5865 1995
rect 5829 1927 5865 1961
rect 5829 1893 5830 1927
rect 5864 1893 5865 1927
rect 5829 1859 5865 1893
rect 5829 1825 5830 1859
rect 5864 1825 5865 1859
rect 5829 1791 5865 1825
rect 5829 1757 5830 1791
rect 5864 1757 5865 1791
rect 5829 1723 5865 1757
rect 5829 1689 5830 1723
rect 5864 1689 5865 1723
rect 5829 1655 5865 1689
rect 5829 1621 5830 1655
rect 5864 1621 5865 1655
rect 5829 1587 5865 1621
rect 5829 1553 5830 1587
rect 5864 1553 5865 1587
rect 5829 1519 5865 1553
rect 5829 1485 5830 1519
rect 5864 1485 5865 1519
rect 5829 1451 5865 1485
rect 5829 1417 5830 1451
rect 5864 1417 5865 1451
rect 5829 1383 5865 1417
rect 5829 1349 5830 1383
rect 5864 1349 5865 1383
rect 5829 1315 5865 1349
rect 5829 1281 5830 1315
rect 5864 1281 5865 1315
rect 5829 1247 5865 1281
rect 5829 1213 5830 1247
rect 5864 1213 5865 1247
rect 5829 1179 5865 1213
rect 5829 1145 5830 1179
rect 5864 1145 5865 1179
rect 5829 1111 5865 1145
rect 5829 1077 5830 1111
rect 5864 1077 5865 1111
rect 5829 1043 5865 1077
rect 5829 1009 5830 1043
rect 5864 1009 5865 1043
rect 5829 975 5865 1009
rect 5829 941 5830 975
rect 5864 941 5865 975
rect 5829 907 5865 941
rect 5829 873 5830 907
rect 5864 873 5865 907
rect 5829 839 5865 873
rect 5829 805 5830 839
rect 5864 805 5865 839
rect 5829 771 5865 805
rect 5829 737 5830 771
rect 5864 737 5865 771
rect 5829 703 5865 737
rect 3356 658 3357 692
rect 3391 658 3392 692
rect 3356 624 3392 658
rect 5829 669 5830 703
rect 5864 669 5865 703
rect 3356 592 3357 624
rect 539 591 3357 592
rect 539 557 573 591
rect 607 557 641 591
rect 675 557 709 591
rect 743 557 777 591
rect 811 557 845 591
rect 879 557 913 591
rect 947 557 1253 591
rect 1287 557 1321 591
rect 1355 557 1389 591
rect 1423 557 1457 591
rect 1491 557 1525 591
rect 1559 557 1593 591
rect 1627 557 1661 591
rect 1695 557 1729 591
rect 1763 557 1797 591
rect 1831 557 1865 591
rect 1899 557 2205 591
rect 2239 557 2273 591
rect 2307 557 2341 591
rect 2375 557 2409 591
rect 2443 557 2559 591
rect 2593 557 2627 591
rect 2661 557 2695 591
rect 2729 557 2763 591
rect 2797 557 2831 591
rect 2865 557 3152 591
rect 3186 557 3220 591
rect 3254 557 3288 591
rect 3322 590 3357 591
rect 3391 592 3392 624
rect 5829 592 5865 669
rect 3391 591 5865 592
rect 3391 590 3426 591
rect 3322 557 3426 590
rect 3460 557 3494 591
rect 3528 557 3562 591
rect 3596 557 3630 591
rect 3664 557 3979 591
rect 4013 557 4047 591
rect 4081 557 4115 591
rect 4149 557 4183 591
rect 4217 557 4251 591
rect 4285 557 4319 591
rect 4353 557 4639 591
rect 4673 557 4707 591
rect 4741 557 4775 591
rect 4809 557 5109 591
rect 5143 557 5177 591
rect 5211 557 5457 591
rect 5491 557 5525 591
rect 5559 557 5593 591
rect 5627 557 5661 591
rect 5695 557 5729 591
rect 5763 557 5797 591
rect 5831 557 5865 591
rect 539 556 5865 557
<< mvnsubdiff >>
rect 130 17343 2270 17344
rect 130 17309 176 17343
rect 210 17309 244 17343
rect 278 17309 312 17343
rect 346 17309 380 17343
rect 414 17309 448 17343
rect 482 17309 516 17343
rect 550 17309 584 17343
rect 618 17309 652 17343
rect 686 17309 720 17343
rect 754 17309 788 17343
rect 822 17309 856 17343
rect 890 17309 924 17343
rect 958 17309 992 17343
rect 1026 17309 1060 17343
rect 1094 17309 1128 17343
rect 1162 17309 1196 17343
rect 1230 17309 1264 17343
rect 1298 17309 1332 17343
rect 1366 17309 1400 17343
rect 1434 17309 1468 17343
rect 1502 17309 1536 17343
rect 1570 17309 1604 17343
rect 1638 17309 1672 17343
rect 1706 17309 1740 17343
rect 1774 17309 1808 17343
rect 1842 17309 1876 17343
rect 1910 17309 1944 17343
rect 1978 17309 2012 17343
rect 2046 17309 2080 17343
rect 2114 17309 2148 17343
rect 2182 17309 2270 17343
rect 130 17308 2270 17309
rect 130 16913 166 17308
rect 2234 17249 2270 17308
rect 2234 17215 2235 17249
rect 2269 17215 2270 17249
rect 2234 17181 2270 17215
rect 2234 17147 2235 17181
rect 2269 17147 2270 17181
rect 2234 17113 2270 17147
rect 2234 17079 2235 17113
rect 2269 17079 2270 17113
rect 2234 17045 2270 17079
rect 2234 17011 2235 17045
rect 2269 17011 2270 17045
rect 2234 16977 2270 17011
rect 2234 16943 2235 16977
rect 2269 16943 2270 16977
rect 2234 16913 2270 16943
rect 130 16909 2270 16913
rect 130 16908 4906 16909
rect 130 16874 234 16908
rect 268 16874 302 16908
rect 336 16874 714 16908
rect 748 16874 836 16908
rect 870 16874 904 16908
rect 938 16874 972 16908
rect 1006 16874 1040 16908
rect 1074 16874 1108 16908
rect 1142 16874 1176 16908
rect 1210 16874 1244 16908
rect 1278 16874 1312 16908
rect 1346 16874 1380 16908
rect 1414 16874 1448 16908
rect 1482 16874 1516 16908
rect 1550 16874 1584 16908
rect 1618 16874 1652 16908
rect 1686 16874 1720 16908
rect 1754 16874 1788 16908
rect 1822 16874 1856 16908
rect 1890 16874 1924 16908
rect 1958 16874 1992 16908
rect 2026 16874 2060 16908
rect 2094 16874 2128 16908
rect 2162 16874 2196 16908
rect 2230 16874 2264 16908
rect 2298 16874 2332 16908
rect 2366 16874 2400 16908
rect 2434 16874 2468 16908
rect 2502 16874 2570 16908
rect 2604 16874 2638 16908
rect 2672 16874 2706 16908
rect 2740 16874 2774 16908
rect 2808 16874 2842 16908
rect 2876 16874 2910 16908
rect 2944 16874 2978 16908
rect 3012 16874 3046 16908
rect 3080 16874 3114 16908
rect 3148 16874 3182 16908
rect 3216 16874 3250 16908
rect 3284 16874 3318 16908
rect 3352 16874 3386 16908
rect 3420 16874 3454 16908
rect 3488 16874 3522 16908
rect 3556 16874 3590 16908
rect 3624 16874 3658 16908
rect 3692 16874 3726 16908
rect 3760 16874 3794 16908
rect 3828 16874 3862 16908
rect 3896 16874 3930 16908
rect 3964 16874 3998 16908
rect 4032 16874 4066 16908
rect 4100 16874 4134 16908
rect 4168 16874 4202 16908
rect 4236 16874 4270 16908
rect 4304 16874 4338 16908
rect 4372 16874 4406 16908
rect 4440 16874 4474 16908
rect 4508 16874 4542 16908
rect 4576 16874 4610 16908
rect 4644 16874 4678 16908
rect 4712 16874 4746 16908
rect 4780 16875 4906 16908
rect 4780 16874 4871 16875
rect 130 16873 4871 16874
rect 130 12149 166 16873
rect 2500 16805 2536 16873
rect 4870 16841 4871 16873
rect 4905 16841 4906 16875
rect 2500 16771 2501 16805
rect 2535 16771 2536 16805
rect 2500 16737 2536 16771
rect 4870 16807 4906 16841
rect 4870 16773 4871 16807
rect 4905 16773 4906 16807
rect 2500 16703 2501 16737
rect 2535 16703 2536 16737
rect 2500 16669 2536 16703
rect 2500 16635 2501 16669
rect 2535 16635 2536 16669
rect 2500 16601 2536 16635
rect 2500 16567 2501 16601
rect 2535 16567 2536 16601
rect 2500 16533 2536 16567
rect 2500 16499 2501 16533
rect 2535 16499 2536 16533
rect 2500 16465 2536 16499
rect 2500 16431 2501 16465
rect 2535 16431 2536 16465
rect 2500 16397 2536 16431
rect 2500 16363 2501 16397
rect 2535 16363 2536 16397
rect 2500 16329 2536 16363
rect 2500 16295 2501 16329
rect 2535 16295 2536 16329
rect 2500 16261 2536 16295
rect 2500 16227 2501 16261
rect 2535 16227 2536 16261
rect 2500 16193 2536 16227
rect 2500 16159 2501 16193
rect 2535 16159 2536 16193
rect 2500 16125 2536 16159
rect 2500 16091 2501 16125
rect 2535 16091 2536 16125
rect 2500 16057 2536 16091
rect 2500 16023 2501 16057
rect 2535 16023 2536 16057
rect 2500 15989 2536 16023
rect 2500 15955 2501 15989
rect 2535 15955 2536 15989
rect 2500 15921 2536 15955
rect 2500 15887 2501 15921
rect 2535 15887 2536 15921
rect 2500 15853 2536 15887
rect 2500 15819 2501 15853
rect 2535 15819 2536 15853
rect 2500 15785 2536 15819
rect 2500 15751 2501 15785
rect 2535 15751 2536 15785
rect 2500 15717 2536 15751
rect 2500 15683 2501 15717
rect 2535 15683 2536 15717
rect 2500 15649 2536 15683
rect 2500 15615 2501 15649
rect 2535 15615 2536 15649
rect 2500 15581 2536 15615
rect 2500 15547 2501 15581
rect 2535 15547 2536 15581
rect 2500 15513 2536 15547
rect 2500 15479 2501 15513
rect 2535 15479 2536 15513
rect 2500 15445 2536 15479
rect 2500 15411 2501 15445
rect 2535 15411 2536 15445
rect 2500 15377 2536 15411
rect 2500 15343 2501 15377
rect 2535 15343 2536 15377
rect 2500 15309 2536 15343
rect 4870 16739 4906 16773
rect 4870 16705 4871 16739
rect 4905 16705 4906 16739
rect 4870 16671 4906 16705
rect 4870 16637 4871 16671
rect 4905 16637 4906 16671
rect 4870 16603 4906 16637
rect 4870 16569 4871 16603
rect 4905 16569 4906 16603
rect 4870 16535 4906 16569
rect 4870 16501 4871 16535
rect 4905 16501 4906 16535
rect 4870 16467 4906 16501
rect 4870 16433 4871 16467
rect 4905 16433 4906 16467
rect 4870 16399 4906 16433
rect 4870 16365 4871 16399
rect 4905 16365 4906 16399
rect 4870 16331 4906 16365
rect 4870 16297 4871 16331
rect 4905 16297 4906 16331
rect 4870 16263 4906 16297
rect 4870 16229 4871 16263
rect 4905 16229 4906 16263
rect 4870 16195 4906 16229
rect 4870 16161 4871 16195
rect 4905 16161 4906 16195
rect 4870 16127 4906 16161
rect 4870 16093 4871 16127
rect 4905 16093 4906 16127
rect 4870 16059 4906 16093
rect 4870 16025 4871 16059
rect 4905 16025 4906 16059
rect 4870 15991 4906 16025
rect 4870 15957 4871 15991
rect 4905 15957 4906 15991
rect 4870 15923 4906 15957
rect 4870 15889 4871 15923
rect 4905 15889 4906 15923
rect 4870 15855 4906 15889
rect 4870 15821 4871 15855
rect 4905 15821 4906 15855
rect 4870 15787 4906 15821
rect 4870 15753 4871 15787
rect 4905 15753 4906 15787
rect 4870 15719 4906 15753
rect 4870 15685 4871 15719
rect 4905 15685 4906 15719
rect 4870 15651 4906 15685
rect 4870 15617 4871 15651
rect 4905 15617 4906 15651
rect 4870 15583 4906 15617
rect 4870 15549 4871 15583
rect 4905 15549 4906 15583
rect 4870 15515 4906 15549
rect 4870 15481 4871 15515
rect 4905 15481 4906 15515
rect 4870 15447 4906 15481
rect 4870 15413 4871 15447
rect 4905 15413 4906 15447
rect 4870 15379 4906 15413
rect 4870 15345 4871 15379
rect 4905 15345 4906 15379
rect 2500 15275 2501 15309
rect 2535 15275 2536 15309
rect 2500 15241 2536 15275
rect 2500 15207 2501 15241
rect 2535 15207 2536 15241
rect 4870 15311 4906 15345
rect 4870 15277 4871 15311
rect 4905 15277 4906 15311
rect 4870 15243 4906 15277
rect 2500 15173 2536 15207
rect 2500 15139 2501 15173
rect 2535 15139 2536 15173
rect 2500 15105 2536 15139
rect 2500 15071 2501 15105
rect 2535 15071 2536 15105
rect 2500 15037 2536 15071
rect 2500 15003 2501 15037
rect 2535 15003 2536 15037
rect 2500 14969 2536 15003
rect 2500 14935 2501 14969
rect 2535 14935 2536 14969
rect 2500 14901 2536 14935
rect 2500 14867 2501 14901
rect 2535 14867 2536 14901
rect 2500 14833 2536 14867
rect 2500 14799 2501 14833
rect 2535 14799 2536 14833
rect 2500 14765 2536 14799
rect 2500 14731 2501 14765
rect 2535 14731 2536 14765
rect 2500 14697 2536 14731
rect 2500 14663 2501 14697
rect 2535 14663 2536 14697
rect 2500 14629 2536 14663
rect 2500 14595 2501 14629
rect 2535 14595 2536 14629
rect 2500 14561 2536 14595
rect 2500 14527 2501 14561
rect 2535 14527 2536 14561
rect 2500 14493 2536 14527
rect 2500 14459 2501 14493
rect 2535 14459 2536 14493
rect 2500 14425 2536 14459
rect 2500 14391 2501 14425
rect 2535 14391 2536 14425
rect 2500 14357 2536 14391
rect 2500 14323 2501 14357
rect 2535 14323 2536 14357
rect 2500 14289 2536 14323
rect 2500 14255 2501 14289
rect 2535 14255 2536 14289
rect 2500 14221 2536 14255
rect 2500 14187 2501 14221
rect 2535 14187 2536 14221
rect 2500 14153 2536 14187
rect 2500 14119 2501 14153
rect 2535 14119 2536 14153
rect 2500 14085 2536 14119
rect 2500 14051 2501 14085
rect 2535 14051 2536 14085
rect 2500 14017 2536 14051
rect 2500 13983 2501 14017
rect 2535 13983 2536 14017
rect 2500 13949 2536 13983
rect 2500 13915 2501 13949
rect 2535 13915 2536 13949
rect 2500 13881 2536 13915
rect 2500 13847 2501 13881
rect 2535 13847 2536 13881
rect 2500 13813 2536 13847
rect 2500 13779 2501 13813
rect 2535 13779 2536 13813
rect 4870 15209 4871 15243
rect 4905 15209 4906 15243
rect 4870 15175 4906 15209
rect 4870 15141 4871 15175
rect 4905 15141 4906 15175
rect 4870 15107 4906 15141
rect 4870 15073 4871 15107
rect 4905 15073 4906 15107
rect 4870 15039 4906 15073
rect 4870 15005 4871 15039
rect 4905 15005 4906 15039
rect 4870 14971 4906 15005
rect 4870 14937 4871 14971
rect 4905 14937 4906 14971
rect 4870 14903 4906 14937
rect 4870 14869 4871 14903
rect 4905 14869 4906 14903
rect 4870 14835 4906 14869
rect 4870 14801 4871 14835
rect 4905 14801 4906 14835
rect 4870 14767 4906 14801
rect 4870 14733 4871 14767
rect 4905 14733 4906 14767
rect 4870 14699 4906 14733
rect 4870 14665 4871 14699
rect 4905 14665 4906 14699
rect 4870 14631 4906 14665
rect 4870 14597 4871 14631
rect 4905 14597 4906 14631
rect 4870 14563 4906 14597
rect 4870 14529 4871 14563
rect 4905 14529 4906 14563
rect 4870 14495 4906 14529
rect 4870 14461 4871 14495
rect 4905 14461 4906 14495
rect 4870 14427 4906 14461
rect 4870 14393 4871 14427
rect 4905 14393 4906 14427
rect 4870 14359 4906 14393
rect 4870 14325 4871 14359
rect 4905 14325 4906 14359
rect 4870 14291 4906 14325
rect 4870 14257 4871 14291
rect 4905 14257 4906 14291
rect 4870 14223 4906 14257
rect 4870 14189 4871 14223
rect 4905 14189 4906 14223
rect 4870 14155 4906 14189
rect 4870 14121 4871 14155
rect 4905 14121 4906 14155
rect 4870 14087 4906 14121
rect 4870 14053 4871 14087
rect 4905 14053 4906 14087
rect 4870 14019 4906 14053
rect 4870 13985 4871 14019
rect 4905 13985 4906 14019
rect 4870 13951 4906 13985
rect 4870 13917 4871 13951
rect 4905 13917 4906 13951
rect 4870 13883 4906 13917
rect 4870 13849 4871 13883
rect 4905 13849 4906 13883
rect 4870 13815 4906 13849
rect 2500 13745 2536 13779
rect 2500 13711 2501 13745
rect 2535 13711 2536 13745
rect 2500 13677 2536 13711
rect 4870 13781 4871 13815
rect 4905 13781 4906 13815
rect 4870 13747 4906 13781
rect 4870 13713 4871 13747
rect 4905 13713 4906 13747
rect 2500 13643 2501 13677
rect 2535 13643 2536 13677
rect 2500 13609 2536 13643
rect 2500 13575 2501 13609
rect 2535 13575 2536 13609
rect 2500 13541 2536 13575
rect 2500 13507 2501 13541
rect 2535 13507 2536 13541
rect 2500 13473 2536 13507
rect 2500 13439 2501 13473
rect 2535 13439 2536 13473
rect 2500 13405 2536 13439
rect 2500 13371 2501 13405
rect 2535 13371 2536 13405
rect 2500 13337 2536 13371
rect 2500 13303 2501 13337
rect 2535 13303 2536 13337
rect 2500 13269 2536 13303
rect 2500 13235 2501 13269
rect 2535 13235 2536 13269
rect 2500 13201 2536 13235
rect 2500 13167 2501 13201
rect 2535 13167 2536 13201
rect 2500 13133 2536 13167
rect 2500 13099 2501 13133
rect 2535 13099 2536 13133
rect 2500 13065 2536 13099
rect 2500 13031 2501 13065
rect 2535 13031 2536 13065
rect 2500 12997 2536 13031
rect 2500 12963 2501 12997
rect 2535 12963 2536 12997
rect 2500 12929 2536 12963
rect 2500 12895 2501 12929
rect 2535 12895 2536 12929
rect 2500 12861 2536 12895
rect 2500 12827 2501 12861
rect 2535 12827 2536 12861
rect 2500 12793 2536 12827
rect 2500 12759 2501 12793
rect 2535 12759 2536 12793
rect 2500 12725 2536 12759
rect 2500 12691 2501 12725
rect 2535 12691 2536 12725
rect 2500 12657 2536 12691
rect 2500 12623 2501 12657
rect 2535 12623 2536 12657
rect 2500 12589 2536 12623
rect 2500 12555 2501 12589
rect 2535 12555 2536 12589
rect 2500 12521 2536 12555
rect 2500 12487 2501 12521
rect 2535 12487 2536 12521
rect 2500 12453 2536 12487
rect 2500 12419 2501 12453
rect 2535 12419 2536 12453
rect 2500 12385 2536 12419
rect 2500 12351 2501 12385
rect 2535 12351 2536 12385
rect 2500 12317 2536 12351
rect 2500 12283 2501 12317
rect 2535 12283 2536 12317
rect 2500 12249 2536 12283
rect 4870 13679 4906 13713
rect 4870 13645 4871 13679
rect 4905 13645 4906 13679
rect 4870 13611 4906 13645
rect 4870 13577 4871 13611
rect 4905 13577 4906 13611
rect 4870 13543 4906 13577
rect 4870 13509 4871 13543
rect 4905 13509 4906 13543
rect 4870 13475 4906 13509
rect 4870 13441 4871 13475
rect 4905 13441 4906 13475
rect 4870 13407 4906 13441
rect 4870 13373 4871 13407
rect 4905 13373 4906 13407
rect 4870 13339 4906 13373
rect 4870 13305 4871 13339
rect 4905 13305 4906 13339
rect 4870 13271 4906 13305
rect 4870 13237 4871 13271
rect 4905 13237 4906 13271
rect 4870 13203 4906 13237
rect 4870 13169 4871 13203
rect 4905 13169 4906 13203
rect 4870 13135 4906 13169
rect 4870 13101 4871 13135
rect 4905 13101 4906 13135
rect 4870 13067 4906 13101
rect 4870 13033 4871 13067
rect 4905 13033 4906 13067
rect 4870 12999 4906 13033
rect 4870 12965 4871 12999
rect 4905 12965 4906 12999
rect 4870 12931 4906 12965
rect 4870 12897 4871 12931
rect 4905 12897 4906 12931
rect 4870 12863 4906 12897
rect 4870 12829 4871 12863
rect 4905 12829 4906 12863
rect 4870 12795 4906 12829
rect 4870 12761 4871 12795
rect 4905 12761 4906 12795
rect 4870 12727 4906 12761
rect 4870 12693 4871 12727
rect 4905 12693 4906 12727
rect 4870 12659 4906 12693
rect 4870 12625 4871 12659
rect 4905 12625 4906 12659
rect 4870 12591 4906 12625
rect 4870 12557 4871 12591
rect 4905 12557 4906 12591
rect 4870 12523 4906 12557
rect 4870 12489 4871 12523
rect 4905 12489 4906 12523
rect 4870 12455 4906 12489
rect 4870 12421 4871 12455
rect 4905 12421 4906 12455
rect 4870 12387 4906 12421
rect 4870 12353 4871 12387
rect 4905 12353 4906 12387
rect 4870 12319 4906 12353
rect 4870 12285 4871 12319
rect 4905 12285 4906 12319
rect 2500 12215 2501 12249
rect 2535 12215 2536 12249
rect 2500 12181 2536 12215
rect 2500 12149 2501 12181
rect 130 12148 2501 12149
rect 130 12114 291 12148
rect 325 12114 359 12148
rect 393 12114 427 12148
rect 461 12114 495 12148
rect 529 12114 563 12148
rect 597 12114 631 12148
rect 665 12114 699 12148
rect 733 12114 767 12148
rect 801 12114 835 12148
rect 869 12114 903 12148
rect 937 12114 971 12148
rect 1005 12114 1039 12148
rect 1073 12114 1107 12148
rect 1141 12114 1175 12148
rect 1209 12114 1243 12148
rect 1277 12114 1311 12148
rect 1345 12114 1379 12148
rect 1413 12114 1447 12148
rect 1481 12114 1515 12148
rect 1549 12114 1583 12148
rect 1617 12114 1651 12148
rect 1685 12114 1719 12148
rect 1753 12114 1787 12148
rect 1821 12114 1855 12148
rect 1889 12114 1923 12148
rect 1957 12114 1991 12148
rect 2025 12114 2059 12148
rect 2093 12114 2127 12148
rect 2161 12114 2195 12148
rect 2229 12114 2263 12148
rect 2297 12114 2331 12148
rect 2365 12114 2399 12148
rect 2433 12147 2501 12148
rect 2535 12149 2536 12181
rect 4870 12182 4906 12285
rect 4870 12149 4871 12182
rect 2535 12148 4871 12149
rect 4905 12148 4906 12182
rect 2535 12147 2596 12148
rect 2433 12114 2596 12147
rect 2630 12114 2664 12148
rect 2698 12114 2732 12148
rect 2766 12114 2800 12148
rect 2834 12114 2868 12148
rect 2902 12114 2936 12148
rect 2970 12114 3004 12148
rect 3038 12114 3072 12148
rect 3106 12114 3140 12148
rect 3174 12114 3208 12148
rect 3242 12114 3276 12148
rect 3310 12114 3344 12148
rect 3378 12114 3412 12148
rect 3446 12114 3480 12148
rect 3514 12114 3548 12148
rect 3582 12114 3616 12148
rect 3650 12114 3684 12148
rect 3718 12114 3752 12148
rect 3786 12114 3820 12148
rect 3854 12114 3888 12148
rect 3922 12114 3956 12148
rect 3990 12114 4024 12148
rect 4058 12114 4092 12148
rect 4126 12114 4160 12148
rect 4194 12114 4228 12148
rect 4262 12114 4296 12148
rect 4330 12114 4364 12148
rect 4398 12114 4432 12148
rect 4466 12114 4500 12148
rect 4534 12114 4568 12148
rect 4602 12114 4636 12148
rect 4670 12114 4704 12148
rect 4738 12114 4772 12148
rect 4806 12114 4906 12148
rect 130 12113 4906 12114
rect 350 12079 507 12113
rect 350 12045 351 12079
rect 385 12045 472 12079
rect 506 12045 507 12079
rect 350 12011 507 12045
rect 2500 12078 2536 12113
rect 2500 12044 2501 12078
rect 2535 12044 2536 12078
rect 350 11977 351 12011
rect 385 11977 472 12011
rect 506 11977 507 12011
rect 350 11943 507 11977
rect 350 11909 351 11943
rect 385 11909 472 11943
rect 506 11909 507 11943
rect 350 11875 507 11909
rect 350 11841 351 11875
rect 385 11841 472 11875
rect 506 11841 507 11875
rect 350 11807 507 11841
rect 350 11773 351 11807
rect 385 11773 472 11807
rect 506 11773 507 11807
rect 350 11739 507 11773
rect 350 11705 351 11739
rect 385 11705 472 11739
rect 506 11705 507 11739
rect 350 11671 507 11705
rect 350 11637 351 11671
rect 385 11637 472 11671
rect 506 11637 507 11671
rect 350 11603 507 11637
rect 350 11569 351 11603
rect 385 11569 472 11603
rect 506 11569 507 11603
rect 350 11535 507 11569
rect 350 11501 351 11535
rect 385 11501 472 11535
rect 506 11501 507 11535
rect 350 11467 507 11501
rect 350 11433 351 11467
rect 385 11433 472 11467
rect 506 11433 507 11467
rect 350 11399 507 11433
rect 350 11365 351 11399
rect 385 11365 472 11399
rect 506 11365 507 11399
rect 350 11331 507 11365
rect 350 11297 351 11331
rect 385 11297 472 11331
rect 506 11297 507 11331
rect 350 11263 507 11297
rect 350 11229 351 11263
rect 385 11229 472 11263
rect 506 11229 507 11263
rect 350 11195 507 11229
rect 350 11161 351 11195
rect 385 11161 472 11195
rect 506 11161 507 11195
rect 350 11127 507 11161
rect 350 11093 351 11127
rect 385 11093 472 11127
rect 506 11093 507 11127
rect 350 11059 507 11093
rect 350 11025 351 11059
rect 385 11025 472 11059
rect 506 11025 507 11059
rect 350 10991 507 11025
rect 350 10957 351 10991
rect 385 10957 472 10991
rect 506 10957 507 10991
rect 350 10923 507 10957
rect 350 10889 351 10923
rect 385 10889 472 10923
rect 506 10889 507 10923
rect 350 10855 507 10889
rect 350 10821 351 10855
rect 385 10821 472 10855
rect 506 10821 507 10855
rect 350 10787 507 10821
rect 350 10753 351 10787
rect 385 10753 472 10787
rect 506 10753 507 10787
rect 350 10719 507 10753
rect 350 10685 351 10719
rect 385 10685 472 10719
rect 506 10685 507 10719
rect 350 10651 507 10685
rect 350 10617 351 10651
rect 385 10617 472 10651
rect 506 10617 507 10651
rect 350 10583 507 10617
rect 350 10549 351 10583
rect 385 10549 472 10583
rect 506 10549 507 10583
rect 350 10515 507 10549
rect 350 10481 351 10515
rect 385 10481 472 10515
rect 506 10481 507 10515
rect 350 10447 507 10481
rect 350 10413 351 10447
rect 385 10413 472 10447
rect 506 10413 507 10447
rect 350 10379 507 10413
rect 350 10345 351 10379
rect 385 10345 472 10379
rect 506 10345 507 10379
rect 350 10311 507 10345
rect 350 10277 351 10311
rect 385 10277 472 10311
rect 506 10277 507 10311
rect 350 10243 507 10277
rect 350 10209 351 10243
rect 385 10209 472 10243
rect 506 10209 507 10243
rect 350 10175 507 10209
rect 350 10141 351 10175
rect 385 10141 472 10175
rect 506 10141 507 10175
rect 350 10107 507 10141
rect 350 10073 351 10107
rect 385 10073 472 10107
rect 506 10073 507 10107
rect 350 10039 507 10073
rect 350 10005 351 10039
rect 385 10005 472 10039
rect 506 10005 507 10039
rect 350 9971 507 10005
rect 350 9937 351 9971
rect 385 9937 472 9971
rect 506 9937 507 9971
rect 350 9903 507 9937
rect 350 9869 351 9903
rect 385 9869 472 9903
rect 506 9869 507 9903
rect 2500 12010 2536 12044
rect 4528 12079 4686 12113
rect 4528 12045 4529 12079
rect 4563 12078 4686 12079
rect 4563 12045 4651 12078
rect 4528 12044 4651 12045
rect 4685 12044 4686 12078
rect 2500 11976 2501 12010
rect 2535 11976 2536 12010
rect 350 9835 507 9869
rect 350 9801 351 9835
rect 385 9801 472 9835
rect 506 9801 507 9835
rect 2500 11942 2536 11976
rect 2500 11908 2501 11942
rect 2535 11908 2536 11942
rect 2500 11874 2536 11908
rect 2500 11840 2501 11874
rect 2535 11840 2536 11874
rect 2500 11806 2536 11840
rect 2500 11772 2501 11806
rect 2535 11772 2536 11806
rect 2500 11738 2536 11772
rect 2500 11704 2501 11738
rect 2535 11704 2536 11738
rect 2500 11670 2536 11704
rect 2500 11636 2501 11670
rect 2535 11636 2536 11670
rect 2500 11602 2536 11636
rect 2500 11568 2501 11602
rect 2535 11568 2536 11602
rect 2500 11534 2536 11568
rect 2500 11500 2501 11534
rect 2535 11500 2536 11534
rect 2500 11466 2536 11500
rect 2500 11432 2501 11466
rect 2535 11432 2536 11466
rect 2500 11398 2536 11432
rect 2500 11364 2501 11398
rect 2535 11364 2536 11398
rect 2500 11330 2536 11364
rect 2500 11296 2501 11330
rect 2535 11296 2536 11330
rect 2500 11262 2536 11296
rect 2500 11228 2501 11262
rect 2535 11228 2536 11262
rect 2500 11194 2536 11228
rect 2500 11160 2501 11194
rect 2535 11160 2536 11194
rect 2500 11126 2536 11160
rect 2500 11092 2501 11126
rect 2535 11092 2536 11126
rect 2500 11058 2536 11092
rect 2500 11024 2501 11058
rect 2535 11024 2536 11058
rect 2500 10990 2536 11024
rect 2500 10956 2501 10990
rect 2535 10956 2536 10990
rect 2500 10922 2536 10956
rect 2500 10888 2501 10922
rect 2535 10888 2536 10922
rect 2500 10854 2536 10888
rect 2500 10820 2501 10854
rect 2535 10820 2536 10854
rect 2500 10786 2536 10820
rect 2500 10752 2501 10786
rect 2535 10752 2536 10786
rect 2500 10718 2536 10752
rect 2500 10684 2501 10718
rect 2535 10684 2536 10718
rect 2500 10650 2536 10684
rect 2500 10616 2501 10650
rect 2535 10616 2536 10650
rect 2500 10582 2536 10616
rect 2500 10548 2501 10582
rect 2535 10548 2536 10582
rect 2500 10514 2536 10548
rect 2500 10480 2501 10514
rect 2535 10480 2536 10514
rect 2500 10446 2536 10480
rect 2500 10412 2501 10446
rect 2535 10412 2536 10446
rect 2500 10378 2536 10412
rect 2500 10344 2501 10378
rect 2535 10344 2536 10378
rect 2500 10310 2536 10344
rect 2500 10276 2501 10310
rect 2535 10276 2536 10310
rect 2500 10242 2536 10276
rect 2500 10208 2501 10242
rect 2535 10208 2536 10242
rect 2500 10174 2536 10208
rect 2500 10140 2501 10174
rect 2535 10140 2536 10174
rect 2500 10106 2536 10140
rect 2500 10072 2501 10106
rect 2535 10072 2536 10106
rect 2500 10038 2536 10072
rect 2500 10004 2501 10038
rect 2535 10004 2536 10038
rect 2500 9970 2536 10004
rect 2500 9936 2501 9970
rect 2535 9936 2536 9970
rect 2500 9902 2536 9936
rect 2500 9868 2501 9902
rect 2535 9868 2536 9902
rect 4528 12011 4686 12044
rect 4528 11977 4529 12011
rect 4563 12010 4686 12011
rect 4563 11977 4651 12010
rect 4528 11976 4651 11977
rect 4685 11976 4686 12010
rect 2500 9834 2536 9868
rect 350 9767 507 9801
rect 350 9733 351 9767
rect 385 9733 472 9767
rect 506 9734 507 9767
rect 2500 9800 2501 9834
rect 2535 9800 2536 9834
rect 4528 11943 4686 11976
rect 4528 11909 4529 11943
rect 4563 11942 4686 11943
rect 4563 11909 4651 11942
rect 4528 11908 4651 11909
rect 4685 11908 4686 11942
rect 4528 11875 4686 11908
rect 4528 11841 4529 11875
rect 4563 11874 4686 11875
rect 4563 11841 4651 11874
rect 4528 11840 4651 11841
rect 4685 11840 4686 11874
rect 4528 11807 4686 11840
rect 4528 11773 4529 11807
rect 4563 11806 4686 11807
rect 4563 11773 4651 11806
rect 4528 11772 4651 11773
rect 4685 11772 4686 11806
rect 4528 11739 4686 11772
rect 4528 11705 4529 11739
rect 4563 11738 4686 11739
rect 4563 11705 4651 11738
rect 4528 11704 4651 11705
rect 4685 11704 4686 11738
rect 4528 11671 4686 11704
rect 4528 11637 4529 11671
rect 4563 11670 4686 11671
rect 4563 11637 4651 11670
rect 4528 11636 4651 11637
rect 4685 11636 4686 11670
rect 4528 11603 4686 11636
rect 4528 11569 4529 11603
rect 4563 11602 4686 11603
rect 4563 11569 4651 11602
rect 4528 11568 4651 11569
rect 4685 11568 4686 11602
rect 4528 11535 4686 11568
rect 4528 11501 4529 11535
rect 4563 11534 4686 11535
rect 4563 11501 4651 11534
rect 4528 11500 4651 11501
rect 4685 11500 4686 11534
rect 4528 11467 4686 11500
rect 4528 11433 4529 11467
rect 4563 11466 4686 11467
rect 4563 11433 4651 11466
rect 4528 11432 4651 11433
rect 4685 11432 4686 11466
rect 4528 11399 4686 11432
rect 4528 11365 4529 11399
rect 4563 11398 4686 11399
rect 4563 11365 4651 11398
rect 4528 11364 4651 11365
rect 4685 11364 4686 11398
rect 4528 11331 4686 11364
rect 4528 11297 4529 11331
rect 4563 11330 4686 11331
rect 4563 11297 4651 11330
rect 4528 11296 4651 11297
rect 4685 11296 4686 11330
rect 4528 11263 4686 11296
rect 4528 11229 4529 11263
rect 4563 11262 4686 11263
rect 4563 11229 4651 11262
rect 4528 11228 4651 11229
rect 4685 11228 4686 11262
rect 4528 11195 4686 11228
rect 4528 11161 4529 11195
rect 4563 11194 4686 11195
rect 4563 11161 4651 11194
rect 4528 11160 4651 11161
rect 4685 11160 4686 11194
rect 4528 11127 4686 11160
rect 4528 11093 4529 11127
rect 4563 11126 4686 11127
rect 4563 11093 4651 11126
rect 4528 11092 4651 11093
rect 4685 11092 4686 11126
rect 4528 11059 4686 11092
rect 4528 11025 4529 11059
rect 4563 11058 4686 11059
rect 4563 11025 4651 11058
rect 4528 11024 4651 11025
rect 4685 11024 4686 11058
rect 4528 10991 4686 11024
rect 4528 10957 4529 10991
rect 4563 10990 4686 10991
rect 4563 10957 4651 10990
rect 4528 10956 4651 10957
rect 4685 10956 4686 10990
rect 4528 10923 4686 10956
rect 4528 10889 4529 10923
rect 4563 10922 4686 10923
rect 4563 10889 4651 10922
rect 4528 10888 4651 10889
rect 4685 10888 4686 10922
rect 4528 10855 4686 10888
rect 4528 10821 4529 10855
rect 4563 10854 4686 10855
rect 4563 10821 4651 10854
rect 4528 10820 4651 10821
rect 4685 10820 4686 10854
rect 4528 10787 4686 10820
rect 4528 10753 4529 10787
rect 4563 10786 4686 10787
rect 4563 10753 4651 10786
rect 4528 10752 4651 10753
rect 4685 10752 4686 10786
rect 4528 10719 4686 10752
rect 4528 10685 4529 10719
rect 4563 10718 4686 10719
rect 4563 10685 4651 10718
rect 4528 10684 4651 10685
rect 4685 10684 4686 10718
rect 4528 10651 4686 10684
rect 4528 10617 4529 10651
rect 4563 10650 4686 10651
rect 4563 10617 4651 10650
rect 4528 10616 4651 10617
rect 4685 10616 4686 10650
rect 4528 10583 4686 10616
rect 4528 10549 4529 10583
rect 4563 10582 4686 10583
rect 4563 10549 4651 10582
rect 4528 10548 4651 10549
rect 4685 10548 4686 10582
rect 4528 10515 4686 10548
rect 4528 10481 4529 10515
rect 4563 10514 4686 10515
rect 4563 10481 4651 10514
rect 4528 10480 4651 10481
rect 4685 10480 4686 10514
rect 4528 10447 4686 10480
rect 4528 10413 4529 10447
rect 4563 10446 4686 10447
rect 4563 10413 4651 10446
rect 4528 10412 4651 10413
rect 4685 10412 4686 10446
rect 4528 10379 4686 10412
rect 4528 10345 4529 10379
rect 4563 10378 4686 10379
rect 4563 10345 4651 10378
rect 4528 10344 4651 10345
rect 4685 10344 4686 10378
rect 4528 10311 4686 10344
rect 4528 10277 4529 10311
rect 4563 10310 4686 10311
rect 4563 10277 4651 10310
rect 4528 10276 4651 10277
rect 4685 10276 4686 10310
rect 4528 10243 4686 10276
rect 4528 10209 4529 10243
rect 4563 10242 4686 10243
rect 4563 10209 4651 10242
rect 4528 10208 4651 10209
rect 4685 10208 4686 10242
rect 4528 10175 4686 10208
rect 4528 10141 4529 10175
rect 4563 10174 4686 10175
rect 4563 10141 4651 10174
rect 4528 10140 4651 10141
rect 4685 10140 4686 10174
rect 4528 10107 4686 10140
rect 4528 10073 4529 10107
rect 4563 10106 4686 10107
rect 4563 10073 4651 10106
rect 4528 10072 4651 10073
rect 4685 10072 4686 10106
rect 4528 10039 4686 10072
rect 4528 10005 4529 10039
rect 4563 10038 4686 10039
rect 4563 10005 4651 10038
rect 4528 10004 4651 10005
rect 4685 10004 4686 10038
rect 4528 9971 4686 10004
rect 4528 9937 4529 9971
rect 4563 9970 4686 9971
rect 4563 9937 4651 9970
rect 4528 9936 4651 9937
rect 4685 9936 4686 9970
rect 4528 9903 4686 9936
rect 4528 9869 4529 9903
rect 4563 9902 4686 9903
rect 4563 9869 4651 9902
rect 4528 9868 4651 9869
rect 4685 9868 4686 9902
rect 4528 9835 4686 9868
rect 2500 9766 2536 9800
rect 2500 9734 2501 9766
rect 506 9733 2501 9734
rect 350 9699 710 9733
rect 744 9699 778 9733
rect 812 9699 846 9733
rect 880 9699 914 9733
rect 948 9699 982 9733
rect 1016 9699 1050 9733
rect 1084 9699 1118 9733
rect 1152 9699 1186 9733
rect 1220 9699 1254 9733
rect 1288 9699 1322 9733
rect 1356 9699 1390 9733
rect 1424 9699 1458 9733
rect 1492 9699 1526 9733
rect 1560 9699 1594 9733
rect 1628 9699 1662 9733
rect 1696 9699 1730 9733
rect 1764 9699 1798 9733
rect 1832 9699 1866 9733
rect 1900 9699 1934 9733
rect 1968 9699 2002 9733
rect 2036 9699 2070 9733
rect 2104 9699 2138 9733
rect 2172 9699 2206 9733
rect 2240 9699 2274 9733
rect 2308 9732 2501 9733
rect 2535 9734 2536 9766
rect 4528 9801 4529 9835
rect 4563 9834 4686 9835
rect 4563 9801 4651 9834
rect 4528 9800 4651 9801
rect 4685 9800 4686 9834
rect 4528 9767 4686 9800
rect 4528 9734 4529 9767
rect 2535 9733 4529 9734
rect 4563 9766 4686 9767
rect 4563 9733 4651 9766
rect 2535 9732 2728 9733
rect 2308 9699 2728 9732
rect 2762 9699 2796 9733
rect 2830 9699 2864 9733
rect 2898 9699 2932 9733
rect 2966 9699 3000 9733
rect 3034 9699 3068 9733
rect 3102 9699 3136 9733
rect 3170 9699 3204 9733
rect 3238 9699 3272 9733
rect 3306 9699 3340 9733
rect 3374 9699 3408 9733
rect 3442 9699 3476 9733
rect 3510 9699 3544 9733
rect 3578 9699 3612 9733
rect 3646 9699 3680 9733
rect 3714 9699 3748 9733
rect 3782 9699 3816 9733
rect 3850 9699 3884 9733
rect 3918 9699 3952 9733
rect 3986 9699 4020 9733
rect 4054 9699 4088 9733
rect 4122 9699 4156 9733
rect 4190 9699 4224 9733
rect 4258 9699 4292 9733
rect 4326 9732 4651 9733
rect 4685 9734 4686 9766
rect 4685 9733 6054 9734
rect 4685 9732 4762 9733
rect 4326 9699 4762 9732
rect 4796 9699 4830 9733
rect 4864 9699 4898 9733
rect 4932 9699 4966 9733
rect 5000 9699 5034 9733
rect 5068 9699 5102 9733
rect 5136 9699 5170 9733
rect 5204 9699 5238 9733
rect 5272 9699 5306 9733
rect 5340 9699 5374 9733
rect 5408 9699 5442 9733
rect 5476 9699 5510 9733
rect 5544 9699 5578 9733
rect 5612 9699 5646 9733
rect 5680 9699 5714 9733
rect 5748 9699 5782 9733
rect 5816 9699 5850 9733
rect 5884 9699 5918 9733
rect 5952 9699 5986 9733
rect 6020 9699 6054 9733
rect 350 9665 351 9699
rect 385 9698 6054 9699
rect 385 9665 386 9698
rect 350 9631 386 9665
rect 350 9597 351 9631
rect 385 9597 386 9631
rect 350 9563 386 9597
rect 350 9529 351 9563
rect 385 9529 386 9563
rect 6018 9650 6054 9698
rect 6018 9616 6019 9650
rect 6053 9616 6054 9650
rect 6018 9582 6054 9616
rect 6018 9548 6019 9582
rect 6053 9548 6054 9582
rect 350 9495 386 9529
rect 350 9461 351 9495
rect 385 9461 386 9495
rect 350 9427 386 9461
rect 350 9393 351 9427
rect 385 9393 386 9427
rect 350 9359 386 9393
rect 350 9325 351 9359
rect 385 9325 386 9359
rect 350 9291 386 9325
rect 350 9257 351 9291
rect 385 9257 386 9291
rect 350 9223 386 9257
rect 350 9189 351 9223
rect 385 9189 386 9223
rect 350 9155 386 9189
rect 350 9121 351 9155
rect 385 9121 386 9155
rect 350 9087 386 9121
rect 350 9053 351 9087
rect 385 9053 386 9087
rect 350 9019 386 9053
rect 350 8985 351 9019
rect 385 8985 386 9019
rect 350 8951 386 8985
rect 350 8917 351 8951
rect 385 8917 386 8951
rect 350 8883 386 8917
rect 350 8849 351 8883
rect 385 8849 386 8883
rect 350 8815 386 8849
rect 350 8781 351 8815
rect 385 8781 386 8815
rect 350 8747 386 8781
rect 350 8713 351 8747
rect 385 8713 386 8747
rect 350 8679 386 8713
rect 350 8645 351 8679
rect 385 8645 386 8679
rect 350 8611 386 8645
rect 350 8577 351 8611
rect 385 8577 386 8611
rect 350 8543 386 8577
rect 350 8509 351 8543
rect 385 8509 386 8543
rect 350 8475 386 8509
rect 350 8441 351 8475
rect 385 8441 386 8475
rect 350 8407 386 8441
rect 350 8373 351 8407
rect 385 8373 386 8407
rect 350 8339 386 8373
rect 350 8305 351 8339
rect 385 8305 386 8339
rect 350 8271 386 8305
rect 350 8237 351 8271
rect 385 8237 386 8271
rect 350 8203 386 8237
rect 350 8169 351 8203
rect 385 8169 386 8203
rect 350 8135 386 8169
rect 350 8101 351 8135
rect 385 8101 386 8135
rect 350 8067 386 8101
rect 350 8033 351 8067
rect 385 8033 386 8067
rect 350 7999 386 8033
rect 350 7965 351 7999
rect 385 7965 386 7999
rect 350 7931 386 7965
rect 350 7897 351 7931
rect 385 7897 386 7931
rect 350 7863 386 7897
rect 350 7829 351 7863
rect 385 7829 386 7863
rect 350 7795 386 7829
rect 350 7761 351 7795
rect 385 7761 386 7795
rect 350 7727 386 7761
rect 350 7693 351 7727
rect 385 7693 386 7727
rect 350 7659 386 7693
rect 350 7625 351 7659
rect 385 7625 386 7659
rect 350 7591 386 7625
rect 350 7557 351 7591
rect 385 7557 386 7591
rect 350 7523 386 7557
rect 350 7489 351 7523
rect 385 7489 386 7523
rect 350 7455 386 7489
rect 350 7421 351 7455
rect 385 7421 386 7455
rect 350 7387 386 7421
rect 350 7353 351 7387
rect 385 7353 386 7387
rect 350 7319 386 7353
rect 350 7285 351 7319
rect 385 7285 386 7319
rect 350 7251 386 7285
rect 350 7217 351 7251
rect 385 7217 386 7251
rect 350 7183 386 7217
rect 350 7149 351 7183
rect 385 7149 386 7183
rect 350 7115 386 7149
rect 350 7081 351 7115
rect 385 7081 386 7115
rect 350 7047 386 7081
rect 350 7013 351 7047
rect 385 7013 386 7047
rect 350 6979 386 7013
rect 350 6945 351 6979
rect 385 6945 386 6979
rect 350 6911 386 6945
rect 350 6877 351 6911
rect 385 6877 386 6911
rect 350 6843 386 6877
rect 350 6809 351 6843
rect 385 6809 386 6843
rect 350 6775 386 6809
rect 350 6741 351 6775
rect 385 6741 386 6775
rect 350 6707 386 6741
rect 350 6673 351 6707
rect 385 6673 386 6707
rect 350 6639 386 6673
rect 350 6605 351 6639
rect 385 6605 386 6639
rect 350 6571 386 6605
rect 350 6537 351 6571
rect 385 6537 386 6571
rect 350 6503 386 6537
rect 350 6469 351 6503
rect 385 6469 386 6503
rect 350 6435 386 6469
rect 350 6401 351 6435
rect 385 6401 386 6435
rect 350 6367 386 6401
rect 350 6333 351 6367
rect 385 6333 386 6367
rect 350 6299 386 6333
rect 350 6265 351 6299
rect 385 6265 386 6299
rect 350 6231 386 6265
rect 350 6197 351 6231
rect 385 6197 386 6231
rect 350 6163 386 6197
rect 350 6129 351 6163
rect 385 6129 386 6163
rect 350 6095 386 6129
rect 350 6061 351 6095
rect 385 6061 386 6095
rect 350 6027 386 6061
rect 350 5993 351 6027
rect 385 5993 386 6027
rect 350 5959 386 5993
rect 350 5925 351 5959
rect 385 5925 386 5959
rect 350 5891 386 5925
rect 350 5857 351 5891
rect 385 5857 386 5891
rect 350 5823 386 5857
rect 350 5789 351 5823
rect 385 5789 386 5823
rect 350 5755 386 5789
rect 350 5721 351 5755
rect 385 5721 386 5755
rect 350 5687 386 5721
rect 350 5653 351 5687
rect 385 5653 386 5687
rect 350 5619 386 5653
rect 350 5585 351 5619
rect 385 5585 386 5619
rect 350 5551 386 5585
rect 350 5517 351 5551
rect 385 5517 386 5551
rect 350 5483 386 5517
rect 350 5449 351 5483
rect 385 5449 386 5483
rect 350 5415 386 5449
rect 350 5381 351 5415
rect 385 5381 386 5415
rect 350 5347 386 5381
rect 350 5313 351 5347
rect 385 5313 386 5347
rect 350 5279 386 5313
rect 350 5245 351 5279
rect 385 5245 386 5279
rect 350 5211 386 5245
rect 350 5177 351 5211
rect 385 5177 386 5211
rect 350 5143 386 5177
rect 350 5109 351 5143
rect 385 5109 386 5143
rect 350 5075 386 5109
rect 350 5041 351 5075
rect 385 5041 386 5075
rect 350 5007 386 5041
rect 350 4973 351 5007
rect 385 4973 386 5007
rect 350 4939 386 4973
rect 350 4905 351 4939
rect 385 4905 386 4939
rect 350 4871 386 4905
rect 350 4837 351 4871
rect 385 4837 386 4871
rect 350 4803 386 4837
rect 350 4769 351 4803
rect 385 4769 386 4803
rect 350 4735 386 4769
rect 350 4701 351 4735
rect 385 4701 386 4735
rect 350 4667 386 4701
rect 350 4633 351 4667
rect 385 4633 386 4667
rect 350 4599 386 4633
rect 350 4565 351 4599
rect 385 4565 386 4599
rect 350 4531 386 4565
rect 350 4497 351 4531
rect 385 4497 386 4531
rect 350 4463 386 4497
rect 350 4429 351 4463
rect 385 4429 386 4463
rect 350 4395 386 4429
rect 350 4361 351 4395
rect 385 4361 386 4395
rect 350 4327 386 4361
rect 350 4293 351 4327
rect 385 4293 386 4327
rect 350 4259 386 4293
rect 350 4225 351 4259
rect 385 4225 386 4259
rect 350 4191 386 4225
rect 350 4157 351 4191
rect 385 4157 386 4191
rect 350 4123 386 4157
rect 350 4089 351 4123
rect 385 4089 386 4123
rect 350 4055 386 4089
rect 350 4021 351 4055
rect 385 4021 386 4055
rect 350 3987 386 4021
rect 350 3953 351 3987
rect 385 3953 386 3987
rect 350 3919 386 3953
rect 350 3885 351 3919
rect 385 3885 386 3919
rect 350 3851 386 3885
rect 350 3817 351 3851
rect 385 3817 386 3851
rect 350 3783 386 3817
rect 350 3749 351 3783
rect 385 3749 386 3783
rect 350 3715 386 3749
rect 350 3681 351 3715
rect 385 3681 386 3715
rect 350 3647 386 3681
rect 350 3613 351 3647
rect 385 3613 386 3647
rect 350 3579 386 3613
rect 350 3545 351 3579
rect 385 3545 386 3579
rect 350 3511 386 3545
rect 350 3477 351 3511
rect 385 3477 386 3511
rect 350 3443 386 3477
rect 350 3409 351 3443
rect 385 3409 386 3443
rect 350 3375 386 3409
rect 350 3341 351 3375
rect 385 3341 386 3375
rect 350 3307 386 3341
rect 350 3273 351 3307
rect 385 3273 386 3307
rect 350 3239 386 3273
rect 350 3205 351 3239
rect 385 3205 386 3239
rect 350 3171 386 3205
rect 350 3137 351 3171
rect 385 3137 386 3171
rect 350 3103 386 3137
rect 350 3069 351 3103
rect 385 3069 386 3103
rect 350 3035 386 3069
rect 350 3001 351 3035
rect 385 3001 386 3035
rect 350 2967 386 3001
rect 350 2933 351 2967
rect 385 2933 386 2967
rect 350 2899 386 2933
rect 350 2865 351 2899
rect 385 2865 386 2899
rect 350 2831 386 2865
rect 350 2797 351 2831
rect 385 2797 386 2831
rect 350 2763 386 2797
rect 350 2729 351 2763
rect 385 2729 386 2763
rect 350 2695 386 2729
rect 350 2661 351 2695
rect 385 2661 386 2695
rect 350 2627 386 2661
rect 350 2593 351 2627
rect 385 2593 386 2627
rect 350 2559 386 2593
rect 350 2525 351 2559
rect 385 2525 386 2559
rect 350 2491 386 2525
rect 350 2457 351 2491
rect 385 2457 386 2491
rect 350 2423 386 2457
rect 350 2389 351 2423
rect 385 2389 386 2423
rect 350 2355 386 2389
rect 350 2321 351 2355
rect 385 2321 386 2355
rect 350 2287 386 2321
rect 350 2253 351 2287
rect 385 2253 386 2287
rect 350 2219 386 2253
rect 350 2185 351 2219
rect 385 2185 386 2219
rect 350 2151 386 2185
rect 350 2117 351 2151
rect 385 2117 386 2151
rect 350 2083 386 2117
rect 350 2049 351 2083
rect 385 2049 386 2083
rect 350 2015 386 2049
rect 350 1981 351 2015
rect 385 1981 386 2015
rect 350 1947 386 1981
rect 350 1913 351 1947
rect 385 1913 386 1947
rect 350 1879 386 1913
rect 350 1845 351 1879
rect 385 1845 386 1879
rect 350 1811 386 1845
rect 350 1777 351 1811
rect 385 1777 386 1811
rect 350 1743 386 1777
rect 350 1709 351 1743
rect 385 1709 386 1743
rect 350 1675 386 1709
rect 350 1641 351 1675
rect 385 1641 386 1675
rect 350 1607 386 1641
rect 350 1573 351 1607
rect 385 1573 386 1607
rect 350 1539 386 1573
rect 350 1505 351 1539
rect 385 1505 386 1539
rect 350 1471 386 1505
rect 350 1437 351 1471
rect 385 1437 386 1471
rect 350 1403 386 1437
rect 350 1369 351 1403
rect 385 1369 386 1403
rect 350 1335 386 1369
rect 350 1301 351 1335
rect 385 1301 386 1335
rect 350 1267 386 1301
rect 350 1233 351 1267
rect 385 1233 386 1267
rect 350 1199 386 1233
rect 350 1165 351 1199
rect 385 1165 386 1199
rect 350 1131 386 1165
rect 350 1097 351 1131
rect 385 1097 386 1131
rect 350 1063 386 1097
rect 350 1029 351 1063
rect 385 1029 386 1063
rect 350 995 386 1029
rect 350 961 351 995
rect 385 961 386 995
rect 350 927 386 961
rect 350 893 351 927
rect 385 893 386 927
rect 350 859 386 893
rect 350 825 351 859
rect 385 825 386 859
rect 350 791 386 825
rect 350 757 351 791
rect 385 757 386 791
rect 350 723 386 757
rect 350 689 351 723
rect 385 689 386 723
rect 350 655 386 689
rect 350 621 351 655
rect 385 621 386 655
rect 350 587 386 621
rect 350 553 351 587
rect 385 553 386 587
rect 6018 9514 6054 9548
rect 6018 9480 6019 9514
rect 6053 9480 6054 9514
rect 6018 9446 6054 9480
rect 6018 9412 6019 9446
rect 6053 9412 6054 9446
rect 6018 9378 6054 9412
rect 6018 9344 6019 9378
rect 6053 9344 6054 9378
rect 6018 9310 6054 9344
rect 6018 9276 6019 9310
rect 6053 9276 6054 9310
rect 6018 9242 6054 9276
rect 6018 9208 6019 9242
rect 6053 9208 6054 9242
rect 6018 9174 6054 9208
rect 6018 9140 6019 9174
rect 6053 9140 6054 9174
rect 6018 9106 6054 9140
rect 6018 9072 6019 9106
rect 6053 9072 6054 9106
rect 6018 9038 6054 9072
rect 6018 9004 6019 9038
rect 6053 9004 6054 9038
rect 6018 8970 6054 9004
rect 6018 8936 6019 8970
rect 6053 8936 6054 8970
rect 6018 8902 6054 8936
rect 6018 8868 6019 8902
rect 6053 8868 6054 8902
rect 6018 8834 6054 8868
rect 6018 8800 6019 8834
rect 6053 8800 6054 8834
rect 6018 8766 6054 8800
rect 6018 8732 6019 8766
rect 6053 8732 6054 8766
rect 6018 8698 6054 8732
rect 6018 8664 6019 8698
rect 6053 8664 6054 8698
rect 6018 8630 6054 8664
rect 6018 8596 6019 8630
rect 6053 8596 6054 8630
rect 6018 8562 6054 8596
rect 6018 8528 6019 8562
rect 6053 8528 6054 8562
rect 6018 8494 6054 8528
rect 6018 8460 6019 8494
rect 6053 8460 6054 8494
rect 6018 8426 6054 8460
rect 6018 8392 6019 8426
rect 6053 8392 6054 8426
rect 6018 8358 6054 8392
rect 6018 8324 6019 8358
rect 6053 8324 6054 8358
rect 6018 8290 6054 8324
rect 6018 8256 6019 8290
rect 6053 8256 6054 8290
rect 6018 8222 6054 8256
rect 6018 8188 6019 8222
rect 6053 8188 6054 8222
rect 6018 8154 6054 8188
rect 6018 8120 6019 8154
rect 6053 8120 6054 8154
rect 6018 8086 6054 8120
rect 6018 8052 6019 8086
rect 6053 8052 6054 8086
rect 6018 8018 6054 8052
rect 6018 7984 6019 8018
rect 6053 7984 6054 8018
rect 6018 7950 6054 7984
rect 6018 7916 6019 7950
rect 6053 7916 6054 7950
rect 6018 7882 6054 7916
rect 6018 7848 6019 7882
rect 6053 7848 6054 7882
rect 6018 7814 6054 7848
rect 6018 7780 6019 7814
rect 6053 7780 6054 7814
rect 6018 7746 6054 7780
rect 6018 7712 6019 7746
rect 6053 7712 6054 7746
rect 6018 7678 6054 7712
rect 6018 7644 6019 7678
rect 6053 7644 6054 7678
rect 6018 7610 6054 7644
rect 6018 7576 6019 7610
rect 6053 7576 6054 7610
rect 6018 7542 6054 7576
rect 6018 7508 6019 7542
rect 6053 7508 6054 7542
rect 6018 7474 6054 7508
rect 6018 7440 6019 7474
rect 6053 7440 6054 7474
rect 6018 7406 6054 7440
rect 6018 7372 6019 7406
rect 6053 7372 6054 7406
rect 6018 7338 6054 7372
rect 6018 7304 6019 7338
rect 6053 7304 6054 7338
rect 6018 7270 6054 7304
rect 6018 7236 6019 7270
rect 6053 7236 6054 7270
rect 6018 7202 6054 7236
rect 6018 7168 6019 7202
rect 6053 7168 6054 7202
rect 6018 7134 6054 7168
rect 6018 7100 6019 7134
rect 6053 7100 6054 7134
rect 6018 7066 6054 7100
rect 6018 7032 6019 7066
rect 6053 7032 6054 7066
rect 6018 6998 6054 7032
rect 6018 6964 6019 6998
rect 6053 6964 6054 6998
rect 6018 6930 6054 6964
rect 6018 6896 6019 6930
rect 6053 6896 6054 6930
rect 6018 6862 6054 6896
rect 6018 6828 6019 6862
rect 6053 6828 6054 6862
rect 6018 6794 6054 6828
rect 6018 6760 6019 6794
rect 6053 6760 6054 6794
rect 6018 6726 6054 6760
rect 6018 6692 6019 6726
rect 6053 6692 6054 6726
rect 6018 6658 6054 6692
rect 6018 6624 6019 6658
rect 6053 6624 6054 6658
rect 6018 6590 6054 6624
rect 6018 6556 6019 6590
rect 6053 6556 6054 6590
rect 6018 6522 6054 6556
rect 6018 6488 6019 6522
rect 6053 6488 6054 6522
rect 6018 6454 6054 6488
rect 6018 6420 6019 6454
rect 6053 6420 6054 6454
rect 6018 6386 6054 6420
rect 6018 6352 6019 6386
rect 6053 6352 6054 6386
rect 6018 6318 6054 6352
rect 6018 6284 6019 6318
rect 6053 6284 6054 6318
rect 6018 6250 6054 6284
rect 6018 6216 6019 6250
rect 6053 6216 6054 6250
rect 6018 6182 6054 6216
rect 6018 6148 6019 6182
rect 6053 6148 6054 6182
rect 6018 6114 6054 6148
rect 6018 6080 6019 6114
rect 6053 6080 6054 6114
rect 6018 6046 6054 6080
rect 6018 6012 6019 6046
rect 6053 6012 6054 6046
rect 6018 5978 6054 6012
rect 6018 5944 6019 5978
rect 6053 5944 6054 5978
rect 6018 5910 6054 5944
rect 6018 5876 6019 5910
rect 6053 5876 6054 5910
rect 6018 5842 6054 5876
rect 6018 5808 6019 5842
rect 6053 5808 6054 5842
rect 6018 5774 6054 5808
rect 6018 5740 6019 5774
rect 6053 5740 6054 5774
rect 6018 5706 6054 5740
rect 6018 5672 6019 5706
rect 6053 5672 6054 5706
rect 6018 5638 6054 5672
rect 6018 5604 6019 5638
rect 6053 5604 6054 5638
rect 6018 5570 6054 5604
rect 6018 5536 6019 5570
rect 6053 5536 6054 5570
rect 6018 5502 6054 5536
rect 6018 5468 6019 5502
rect 6053 5468 6054 5502
rect 6018 5434 6054 5468
rect 6018 5400 6019 5434
rect 6053 5400 6054 5434
rect 6018 5366 6054 5400
rect 6018 5332 6019 5366
rect 6053 5332 6054 5366
rect 6018 5298 6054 5332
rect 6018 5264 6019 5298
rect 6053 5264 6054 5298
rect 6018 5230 6054 5264
rect 6018 5196 6019 5230
rect 6053 5196 6054 5230
rect 6018 5162 6054 5196
rect 6018 5128 6019 5162
rect 6053 5128 6054 5162
rect 6018 5094 6054 5128
rect 6018 5060 6019 5094
rect 6053 5060 6054 5094
rect 6018 5026 6054 5060
rect 6018 4992 6019 5026
rect 6053 4992 6054 5026
rect 6018 4958 6054 4992
rect 6018 4924 6019 4958
rect 6053 4924 6054 4958
rect 6018 4890 6054 4924
rect 6018 4856 6019 4890
rect 6053 4856 6054 4890
rect 6018 4822 6054 4856
rect 6018 4788 6019 4822
rect 6053 4788 6054 4822
rect 6018 4754 6054 4788
rect 6018 4720 6019 4754
rect 6053 4720 6054 4754
rect 6018 4686 6054 4720
rect 6018 4652 6019 4686
rect 6053 4652 6054 4686
rect 6018 4618 6054 4652
rect 6018 4584 6019 4618
rect 6053 4584 6054 4618
rect 6018 4550 6054 4584
rect 6018 4516 6019 4550
rect 6053 4516 6054 4550
rect 6018 4482 6054 4516
rect 6018 4448 6019 4482
rect 6053 4448 6054 4482
rect 6018 4414 6054 4448
rect 6018 4380 6019 4414
rect 6053 4380 6054 4414
rect 6018 4346 6054 4380
rect 6018 4312 6019 4346
rect 6053 4312 6054 4346
rect 6018 4278 6054 4312
rect 6018 4244 6019 4278
rect 6053 4244 6054 4278
rect 6018 4210 6054 4244
rect 6018 4176 6019 4210
rect 6053 4176 6054 4210
rect 6018 4142 6054 4176
rect 6018 4108 6019 4142
rect 6053 4108 6054 4142
rect 6018 4074 6054 4108
rect 6018 4040 6019 4074
rect 6053 4040 6054 4074
rect 6018 4006 6054 4040
rect 6018 3972 6019 4006
rect 6053 3972 6054 4006
rect 6018 3938 6054 3972
rect 6018 3904 6019 3938
rect 6053 3904 6054 3938
rect 6018 3870 6054 3904
rect 6018 3836 6019 3870
rect 6053 3836 6054 3870
rect 6018 3802 6054 3836
rect 6018 3768 6019 3802
rect 6053 3768 6054 3802
rect 6018 3734 6054 3768
rect 6018 3700 6019 3734
rect 6053 3700 6054 3734
rect 6018 3666 6054 3700
rect 6018 3632 6019 3666
rect 6053 3632 6054 3666
rect 6018 3598 6054 3632
rect 6018 3564 6019 3598
rect 6053 3564 6054 3598
rect 6018 3530 6054 3564
rect 6018 3496 6019 3530
rect 6053 3496 6054 3530
rect 6018 3462 6054 3496
rect 6018 3428 6019 3462
rect 6053 3428 6054 3462
rect 6018 3394 6054 3428
rect 6018 3360 6019 3394
rect 6053 3360 6054 3394
rect 6018 3326 6054 3360
rect 6018 3292 6019 3326
rect 6053 3292 6054 3326
rect 6018 3258 6054 3292
rect 6018 3224 6019 3258
rect 6053 3224 6054 3258
rect 6018 3190 6054 3224
rect 6018 3156 6019 3190
rect 6053 3156 6054 3190
rect 6018 3122 6054 3156
rect 6018 3088 6019 3122
rect 6053 3088 6054 3122
rect 6018 3054 6054 3088
rect 6018 3020 6019 3054
rect 6053 3020 6054 3054
rect 6018 2986 6054 3020
rect 6018 2952 6019 2986
rect 6053 2952 6054 2986
rect 6018 2918 6054 2952
rect 6018 2884 6019 2918
rect 6053 2884 6054 2918
rect 6018 2850 6054 2884
rect 6018 2816 6019 2850
rect 6053 2816 6054 2850
rect 6018 2782 6054 2816
rect 6018 2748 6019 2782
rect 6053 2748 6054 2782
rect 6018 2714 6054 2748
rect 6018 2680 6019 2714
rect 6053 2680 6054 2714
rect 6018 2646 6054 2680
rect 6018 2612 6019 2646
rect 6053 2612 6054 2646
rect 6018 2578 6054 2612
rect 6018 2544 6019 2578
rect 6053 2544 6054 2578
rect 6018 2510 6054 2544
rect 6018 2476 6019 2510
rect 6053 2476 6054 2510
rect 6018 2442 6054 2476
rect 6018 2408 6019 2442
rect 6053 2408 6054 2442
rect 6018 2374 6054 2408
rect 6018 2340 6019 2374
rect 6053 2340 6054 2374
rect 6018 2306 6054 2340
rect 6018 2272 6019 2306
rect 6053 2272 6054 2306
rect 6018 2238 6054 2272
rect 6018 2204 6019 2238
rect 6053 2204 6054 2238
rect 6018 2170 6054 2204
rect 6018 2136 6019 2170
rect 6053 2136 6054 2170
rect 6018 2102 6054 2136
rect 6018 2068 6019 2102
rect 6053 2068 6054 2102
rect 6018 2034 6054 2068
rect 6018 2000 6019 2034
rect 6053 2000 6054 2034
rect 6018 1966 6054 2000
rect 6018 1932 6019 1966
rect 6053 1932 6054 1966
rect 6018 1898 6054 1932
rect 6018 1864 6019 1898
rect 6053 1864 6054 1898
rect 6018 1830 6054 1864
rect 6018 1796 6019 1830
rect 6053 1796 6054 1830
rect 6018 1762 6054 1796
rect 6018 1728 6019 1762
rect 6053 1728 6054 1762
rect 6018 1694 6054 1728
rect 6018 1660 6019 1694
rect 6053 1660 6054 1694
rect 6018 1626 6054 1660
rect 6018 1592 6019 1626
rect 6053 1592 6054 1626
rect 6018 1558 6054 1592
rect 6018 1524 6019 1558
rect 6053 1524 6054 1558
rect 6018 1490 6054 1524
rect 6018 1456 6019 1490
rect 6053 1456 6054 1490
rect 6018 1422 6054 1456
rect 6018 1388 6019 1422
rect 6053 1388 6054 1422
rect 6018 1354 6054 1388
rect 6018 1320 6019 1354
rect 6053 1320 6054 1354
rect 6018 1286 6054 1320
rect 6018 1252 6019 1286
rect 6053 1252 6054 1286
rect 6018 1218 6054 1252
rect 6018 1184 6019 1218
rect 6053 1184 6054 1218
rect 6018 1150 6054 1184
rect 6018 1116 6019 1150
rect 6053 1116 6054 1150
rect 6018 1082 6054 1116
rect 6018 1048 6019 1082
rect 6053 1048 6054 1082
rect 6018 1014 6054 1048
rect 6018 980 6019 1014
rect 6053 980 6054 1014
rect 6018 946 6054 980
rect 6018 912 6019 946
rect 6053 912 6054 946
rect 6018 878 6054 912
rect 6018 844 6019 878
rect 6053 844 6054 878
rect 6018 810 6054 844
rect 6018 776 6019 810
rect 6053 776 6054 810
rect 6018 742 6054 776
rect 6018 708 6019 742
rect 6053 708 6054 742
rect 6018 674 6054 708
rect 6018 640 6019 674
rect 6053 640 6054 674
rect 6018 606 6054 640
rect 6018 572 6019 606
rect 6053 572 6054 606
rect 350 403 386 553
rect 6018 538 6054 572
rect 6018 504 6019 538
rect 6053 504 6054 538
rect 6018 435 6054 504
rect 6018 403 6019 435
rect 350 402 6019 403
rect 350 368 384 402
rect 418 368 452 402
rect 486 368 520 402
rect 554 368 588 402
rect 622 368 656 402
rect 690 368 724 402
rect 758 368 792 402
rect 826 368 860 402
rect 894 368 928 402
rect 962 368 996 402
rect 1030 368 1064 402
rect 1098 368 1132 402
rect 1166 368 1200 402
rect 1234 368 1268 402
rect 1302 368 1336 402
rect 1370 368 1404 402
rect 1438 368 1472 402
rect 1506 368 1540 402
rect 1574 368 1608 402
rect 1642 368 1676 402
rect 1710 368 1744 402
rect 1778 368 1812 402
rect 1846 368 1880 402
rect 1914 368 1948 402
rect 1982 368 2016 402
rect 2050 368 2084 402
rect 2118 368 2152 402
rect 2186 368 2220 402
rect 2254 368 2288 402
rect 2322 368 2356 402
rect 2390 368 2424 402
rect 2458 368 2492 402
rect 2526 368 2560 402
rect 2594 368 2628 402
rect 2662 368 2696 402
rect 2730 368 2764 402
rect 2798 368 2832 402
rect 2866 368 2900 402
rect 2934 368 2968 402
rect 3002 368 3036 402
rect 3070 368 3104 402
rect 3138 368 3172 402
rect 3206 368 3240 402
rect 3274 368 3308 402
rect 3342 368 3376 402
rect 3410 368 3444 402
rect 3478 368 3512 402
rect 3546 368 3580 402
rect 3614 368 3648 402
rect 3682 368 3716 402
rect 3750 368 3784 402
rect 3818 368 3852 402
rect 3886 368 3920 402
rect 3954 368 3988 402
rect 4022 368 4056 402
rect 4090 368 4124 402
rect 4158 368 4192 402
rect 4226 368 4260 402
rect 4294 368 4328 402
rect 4362 368 4396 402
rect 4430 368 4464 402
rect 4498 368 4532 402
rect 4566 368 4600 402
rect 4634 368 4668 402
rect 4702 368 4736 402
rect 4770 368 4804 402
rect 4838 368 4872 402
rect 4906 368 4940 402
rect 4974 368 5008 402
rect 5042 368 5076 402
rect 5110 368 5144 402
rect 5178 368 5212 402
rect 5246 368 5280 402
rect 5314 368 5348 402
rect 5382 368 5416 402
rect 5450 368 5484 402
rect 5518 368 5552 402
rect 5586 368 5620 402
rect 5654 368 5688 402
rect 5722 368 5756 402
rect 5790 368 5824 402
rect 5858 368 5892 402
rect 5926 401 6019 402
rect 6053 401 6054 435
rect 5926 368 6054 401
rect 350 367 6054 368
<< psubdiffcont >>
rect 10147 34512 10181 34546
rect 10215 34512 10249 34546
rect 10283 34512 10317 34546
rect 10351 34512 10385 34546
rect 10419 34512 10453 34546
rect 10487 34512 10521 34546
rect 10555 34512 10589 34546
rect 10623 34512 10657 34546
rect 10691 34512 10725 34546
rect 10759 34512 10793 34546
rect 10827 34512 10861 34546
rect 10895 34512 10929 34546
rect 10963 34512 10997 34546
rect 11031 34512 11065 34546
rect 11099 34512 11133 34546
rect 11167 34512 11201 34546
rect 11235 34512 11269 34546
rect 11303 34512 11337 34546
rect 11371 34512 11405 34546
rect 11439 34512 11473 34546
rect 11507 34512 11541 34546
rect 11575 34512 11609 34546
rect 11643 34512 11677 34546
rect 11711 34512 11745 34546
rect 11779 34512 11813 34546
rect 11847 34512 11881 34546
rect 11915 34512 11949 34546
rect 11983 34512 12017 34546
rect 12051 34512 12085 34546
rect 12119 34512 12153 34546
rect 12187 34512 12221 34546
rect 12255 34512 12289 34546
rect 12323 34512 12357 34546
rect 12391 34512 12425 34546
rect 12459 34512 12493 34546
rect 12527 34512 12561 34546
rect 12595 34512 12629 34546
rect 12663 34512 12697 34546
rect 12731 34512 12765 34546
rect 12799 34512 12833 34546
rect 12867 34512 12901 34546
rect 12935 34512 12969 34546
rect 13003 34512 13037 34546
rect 13071 34512 13105 34546
rect 13139 34512 13173 34546
rect 13207 34512 13241 34546
rect 13275 34512 13309 34546
rect 13343 34512 13377 34546
rect 13411 34512 13445 34546
rect 13479 34512 13513 34546
rect 13547 34512 13581 34546
rect 13615 34512 13649 34546
rect 13683 34512 13717 34546
rect 13751 34512 13785 34546
rect 13819 34512 13853 34546
rect 13887 34512 13921 34546
rect 13955 34512 13989 34546
rect 14023 34512 14057 34546
rect 14091 34512 14125 34546
rect 10040 34444 10074 34478
rect 10040 34376 10074 34410
rect 10040 34308 10074 34342
rect 10040 34240 10074 34274
rect 10040 34172 10074 34206
rect 10040 34104 10074 34138
rect 10040 34036 10074 34070
rect 10040 33968 10074 34002
rect 10040 33900 10074 33934
rect 10040 33832 10074 33866
rect 10040 33764 10074 33798
rect 10040 33696 10074 33730
rect 10040 33628 10074 33662
rect 10040 33560 10074 33594
rect 10040 33492 10074 33526
rect 10040 33424 10074 33458
rect 10040 33356 10074 33390
rect 10040 33288 10074 33322
rect 10040 33220 10074 33254
rect 10040 33152 10074 33186
rect 10040 33084 10074 33118
rect 10040 33016 10074 33050
rect 10040 32948 10074 32982
rect 10040 32880 10074 32914
rect 10040 32812 10074 32846
rect 10040 32744 10074 32778
rect 10040 32676 10074 32710
rect 10040 32608 10074 32642
rect 10040 32540 10074 32574
rect 10040 32472 10074 32506
rect 10040 32404 10074 32438
rect 10040 32336 10074 32370
rect 10040 32268 10074 32302
rect 14159 34351 14193 34385
rect 14159 34283 14193 34317
rect 14159 34215 14193 34249
rect 14159 34147 14193 34181
rect 14159 34079 14193 34113
rect 14159 34011 14193 34045
rect 14159 33943 14193 33977
rect 14159 33875 14193 33909
rect 14159 33807 14193 33841
rect 14159 33739 14193 33773
rect 14159 33671 14193 33705
rect 14159 33603 14193 33637
rect 14159 33535 14193 33569
rect 14159 33467 14193 33501
rect 14159 33399 14193 33433
rect 14159 33331 14193 33365
rect 14159 33263 14193 33297
rect 14159 33195 14193 33229
rect 14159 33127 14193 33161
rect 14159 33059 14193 33093
rect 14159 32991 14193 33025
rect 14159 32923 14193 32957
rect 14159 32855 14193 32889
rect 14159 32787 14193 32821
rect 14159 32719 14193 32753
rect 14159 32651 14193 32685
rect 14159 32583 14193 32617
rect 14159 32515 14193 32549
rect 14159 32447 14193 32481
rect 14159 32379 14193 32413
rect 14159 32311 14193 32345
rect 10108 32260 10142 32294
rect 10193 32260 10227 32294
rect 10278 32260 10312 32294
rect 10363 32260 10397 32294
rect 10448 32260 10482 32294
rect 10533 32260 10567 32294
rect 10618 32260 10652 32294
rect 10703 32260 10737 32294
rect 10788 32260 10822 32294
rect 10873 32260 10907 32294
rect 10958 32260 10992 32294
rect 11043 32260 11077 32294
rect 11128 32260 11162 32294
rect 11213 32260 11247 32294
rect 11298 32260 11332 32294
rect 11383 32260 11417 32294
rect 11468 32260 11502 32294
rect 11553 32260 11587 32294
rect 11638 32260 11672 32294
rect 11723 32260 11757 32294
rect 11808 32260 11842 32294
rect 11893 32260 11927 32294
rect 11978 32260 12012 32294
rect 12063 32260 12097 32294
rect 12148 32260 12182 32294
rect 12233 32260 12267 32294
rect 12318 32260 12352 32294
rect 12403 32260 12437 32294
rect 12488 32260 12522 32294
rect 12573 32260 12607 32294
rect 12658 32260 12692 32294
rect 12743 32260 12777 32294
rect 12828 32260 12862 32294
rect 12913 32260 12947 32294
rect 12998 32260 13032 32294
rect 13083 32260 13117 32294
rect 13167 32260 13201 32294
rect 13251 32260 13285 32294
rect 13335 32260 13369 32294
rect 13419 32260 13453 32294
rect 13503 32260 13537 32294
rect 13587 32260 13621 32294
rect 13671 32260 13705 32294
rect 13755 32260 13789 32294
rect 13839 32260 13873 32294
rect 13923 32260 13957 32294
rect 14007 32260 14041 32294
rect 14091 32260 14125 32294
rect 10040 32200 10074 32234
rect 14159 32243 14193 32277
rect 10040 32132 10074 32166
rect 14159 32175 14193 32209
rect 10040 32064 10074 32098
rect 10040 31996 10074 32030
rect 10040 31928 10074 31962
rect 10040 31860 10074 31894
rect 10040 31792 10074 31826
rect 10040 31724 10074 31758
rect 10040 31656 10074 31690
rect 10040 31588 10074 31622
rect 10040 31520 10074 31554
rect 10040 31452 10074 31486
rect 10040 31384 10074 31418
rect 10040 31316 10074 31350
rect 10040 31248 10074 31282
rect 10040 31180 10074 31214
rect 10040 31112 10074 31146
rect 10040 31044 10074 31078
rect 10040 30976 10074 31010
rect 10040 30908 10074 30942
rect 10040 30840 10074 30874
rect 10040 30772 10074 30806
rect 10040 30704 10074 30738
rect 10040 30636 10074 30670
rect 10040 30568 10074 30602
rect 10040 30500 10074 30534
rect 10040 30432 10074 30466
rect 10040 30364 10074 30398
rect 10040 30296 10074 30330
rect 10040 30228 10074 30262
rect 10040 30160 10074 30194
rect 10040 30092 10074 30126
rect 10040 30024 10074 30058
rect 14159 32107 14193 32141
rect 14159 32039 14193 32073
rect 14159 31971 14193 32005
rect 14159 31903 14193 31937
rect 14159 31835 14193 31869
rect 14159 31767 14193 31801
rect 14159 31699 14193 31733
rect 14159 31631 14193 31665
rect 14159 31563 14193 31597
rect 14159 31495 14193 31529
rect 14159 31427 14193 31461
rect 14159 31359 14193 31393
rect 14159 31291 14193 31325
rect 14159 31223 14193 31257
rect 14159 31155 14193 31189
rect 14159 31087 14193 31121
rect 14159 31019 14193 31053
rect 14159 30951 14193 30985
rect 14159 30883 14193 30917
rect 14159 30815 14193 30849
rect 14159 30747 14193 30781
rect 14159 30679 14193 30713
rect 14159 30611 14193 30645
rect 14159 30543 14193 30577
rect 14159 30475 14193 30509
rect 14159 30407 14193 30441
rect 14159 30339 14193 30373
rect 14159 30271 14193 30305
rect 14159 30203 14193 30237
rect 14159 30135 14193 30169
rect 14159 30067 14193 30101
rect 10108 30009 10142 30043
rect 10193 30009 10227 30043
rect 10278 30009 10312 30043
rect 10363 30009 10397 30043
rect 10448 30009 10482 30043
rect 10533 30009 10567 30043
rect 10618 30009 10652 30043
rect 10703 30009 10737 30043
rect 10788 30009 10822 30043
rect 10873 30009 10907 30043
rect 10958 30009 10992 30043
rect 11043 30009 11077 30043
rect 11128 30009 11162 30043
rect 11213 30009 11247 30043
rect 11298 30009 11332 30043
rect 11383 30009 11417 30043
rect 11468 30009 11502 30043
rect 11553 30009 11587 30043
rect 11638 30009 11672 30043
rect 11723 30009 11757 30043
rect 11808 30009 11842 30043
rect 11893 30009 11927 30043
rect 11978 30009 12012 30043
rect 12063 30009 12097 30043
rect 12148 30009 12182 30043
rect 12233 30009 12267 30043
rect 12318 30009 12352 30043
rect 12403 30009 12437 30043
rect 12488 30009 12522 30043
rect 12573 30009 12607 30043
rect 12658 30009 12692 30043
rect 12743 30009 12777 30043
rect 12828 30009 12862 30043
rect 12913 30009 12947 30043
rect 12998 30009 13032 30043
rect 13083 30009 13117 30043
rect 13167 30009 13201 30043
rect 13251 30009 13285 30043
rect 13335 30009 13369 30043
rect 13419 30009 13453 30043
rect 13503 30009 13537 30043
rect 13587 30009 13621 30043
rect 13671 30009 13705 30043
rect 13755 30009 13789 30043
rect 13839 30009 13873 30043
rect 13923 30009 13957 30043
rect 14007 30009 14041 30043
rect 14091 30009 14125 30043
rect 10040 29956 10074 29990
rect 14159 29999 14193 30033
rect 10040 29888 10074 29922
rect 14159 29931 14193 29965
rect 10040 29820 10074 29854
rect 10040 29752 10074 29786
rect 10040 29684 10074 29718
rect 10040 29616 10074 29650
rect 10040 29548 10074 29582
rect 10040 29480 10074 29514
rect 10040 29412 10074 29446
rect 10040 29344 10074 29378
rect 10040 29276 10074 29310
rect 10040 29208 10074 29242
rect 10040 29140 10074 29174
rect 10040 29072 10074 29106
rect 10040 29004 10074 29038
rect 10040 28936 10074 28970
rect 10040 28868 10074 28902
rect 10040 28800 10074 28834
rect 10040 28732 10074 28766
rect 10040 28664 10074 28698
rect 10040 28596 10074 28630
rect 10040 28528 10074 28562
rect 10040 28460 10074 28494
rect 10040 28392 10074 28426
rect 10040 28324 10074 28358
rect 10040 28256 10074 28290
rect 10040 28188 10074 28222
rect 10040 28120 10074 28154
rect 10040 28052 10074 28086
rect 10040 27984 10074 28018
rect 10040 27916 10074 27950
rect 10040 27848 10074 27882
rect 14159 29863 14193 29897
rect 14159 29795 14193 29829
rect 14159 29727 14193 29761
rect 14159 29659 14193 29693
rect 14159 29591 14193 29625
rect 14159 29523 14193 29557
rect 14159 29455 14193 29489
rect 14159 29387 14193 29421
rect 14159 29319 14193 29353
rect 14159 29251 14193 29285
rect 14159 29183 14193 29217
rect 14159 29115 14193 29149
rect 14159 29047 14193 29081
rect 14159 28979 14193 29013
rect 14159 28911 14193 28945
rect 14159 28843 14193 28877
rect 14159 28775 14193 28809
rect 14159 28707 14193 28741
rect 14159 28639 14193 28673
rect 14159 28571 14193 28605
rect 14159 28503 14193 28537
rect 14159 28435 14193 28469
rect 14159 28367 14193 28401
rect 14159 28299 14193 28333
rect 14159 28231 14193 28265
rect 14159 28163 14193 28197
rect 14159 28095 14193 28129
rect 14159 28027 14193 28061
rect 14159 27959 14193 27993
rect 14159 27891 14193 27925
rect 14159 27823 14193 27857
rect 10108 27755 10142 27789
rect 10176 27755 10210 27789
rect 10244 27755 10278 27789
rect 10312 27755 10346 27789
rect 10380 27755 10414 27789
rect 10448 27755 10482 27789
rect 10516 27755 10550 27789
rect 10584 27755 10618 27789
rect 10652 27755 10686 27789
rect 10720 27755 10754 27789
rect 10788 27755 10822 27789
rect 10856 27755 10890 27789
rect 10924 27755 10958 27789
rect 10992 27755 11026 27789
rect 11060 27755 11094 27789
rect 11128 27755 11162 27789
rect 11196 27755 11230 27789
rect 11264 27755 11298 27789
rect 11332 27755 11366 27789
rect 11400 27755 11434 27789
rect 11468 27755 11502 27789
rect 11536 27755 11570 27789
rect 11604 27755 11638 27789
rect 11672 27755 11706 27789
rect 11740 27755 11774 27789
rect 11808 27755 11842 27789
rect 11876 27755 11910 27789
rect 11944 27755 11978 27789
rect 12012 27755 12046 27789
rect 12080 27755 12114 27789
rect 12148 27755 12182 27789
rect 12216 27755 12250 27789
rect 12284 27755 12318 27789
rect 12352 27755 12386 27789
rect 12420 27755 12454 27789
rect 12488 27755 12522 27789
rect 12556 27755 12590 27789
rect 12624 27755 12658 27789
rect 12692 27755 12726 27789
rect 12760 27755 12794 27789
rect 12828 27755 12862 27789
rect 12896 27755 12930 27789
rect 12964 27755 12998 27789
rect 13032 27755 13066 27789
rect 13100 27755 13134 27789
rect 13168 27755 13202 27789
rect 13236 27755 13270 27789
rect 13304 27755 13338 27789
rect 13372 27755 13406 27789
rect 13440 27755 13474 27789
rect 13508 27755 13542 27789
rect 13576 27755 13610 27789
rect 13644 27755 13678 27789
rect 13712 27755 13746 27789
rect 13780 27755 13814 27789
rect 13848 27755 13882 27789
rect 13916 27755 13950 27789
rect 13984 27755 14018 27789
rect 14052 27755 14086 27789
<< nsubdiffcont >>
rect 9917 34762 9951 34796
rect 9985 34762 10019 34796
rect 10053 34762 10087 34796
rect 10121 34762 10155 34796
rect 10189 34762 10223 34796
rect 10257 34762 10291 34796
rect 10325 34762 10359 34796
rect 10393 34762 10427 34796
rect 10461 34762 10495 34796
rect 10529 34762 10563 34796
rect 10597 34762 10631 34796
rect 10665 34762 10699 34796
rect 10733 34762 10767 34796
rect 10801 34762 10835 34796
rect 10869 34762 10903 34796
rect 10937 34762 10971 34796
rect 11005 34762 11039 34796
rect 11073 34762 11107 34796
rect 11141 34762 11175 34796
rect 11209 34762 11243 34796
rect 11277 34762 11311 34796
rect 11345 34762 11379 34796
rect 11413 34762 11447 34796
rect 11481 34762 11515 34796
rect 11549 34762 11583 34796
rect 11617 34762 11651 34796
rect 11685 34762 11719 34796
rect 11753 34762 11787 34796
rect 11821 34762 11855 34796
rect 11889 34762 11923 34796
rect 11957 34762 11991 34796
rect 12025 34762 12059 34796
rect 12093 34762 12127 34796
rect 12161 34762 12195 34796
rect 12229 34762 12263 34796
rect 12297 34762 12331 34796
rect 12365 34762 12399 34796
rect 12433 34762 12467 34796
rect 12501 34762 12535 34796
rect 12569 34762 12603 34796
rect 12637 34762 12671 34796
rect 12705 34762 12739 34796
rect 12773 34762 12807 34796
rect 12841 34762 12875 34796
rect 12909 34762 12943 34796
rect 12977 34762 13011 34796
rect 13045 34762 13079 34796
rect 13113 34762 13147 34796
rect 13181 34762 13215 34796
rect 13249 34762 13283 34796
rect 13317 34762 13351 34796
rect 13385 34762 13419 34796
rect 13453 34762 13487 34796
rect 13521 34762 13555 34796
rect 13589 34762 13623 34796
rect 13657 34762 13691 34796
rect 13725 34762 13759 34796
rect 13793 34762 13827 34796
rect 13861 34762 13895 34796
rect 13929 34762 13963 34796
rect 13997 34762 14031 34796
rect 14065 34762 14099 34796
rect 14133 34762 14167 34796
rect 14201 34762 14235 34796
rect 14269 34762 14303 34796
rect 14337 34762 14371 34796
rect 9789 34694 9823 34728
rect 9789 34626 9823 34660
rect 9789 34558 9823 34592
rect 14405 34670 14439 34704
rect 9789 34490 9823 34524
rect 9789 34422 9823 34456
rect 9789 34354 9823 34388
rect 9789 34286 9823 34320
rect 9789 34218 9823 34252
rect 9789 34150 9823 34184
rect 9789 34082 9823 34116
rect 9789 34014 9823 34048
rect 9789 33946 9823 33980
rect 9789 33878 9823 33912
rect 9789 33810 9823 33844
rect 9789 33742 9823 33776
rect 9119 33579 9153 33613
rect 9119 33511 9153 33545
rect 9119 33443 9153 33477
rect 9119 33375 9153 33409
rect 9119 33307 9153 33341
rect 9119 33239 9153 33273
rect 9119 33171 9153 33205
rect 9119 33103 9153 33137
rect 9119 33035 9153 33069
rect 9119 32967 9153 33001
rect 9119 32899 9153 32933
rect 9119 32831 9153 32865
rect 9119 32763 9153 32797
rect 9119 32695 9153 32729
rect 9119 32627 9153 32661
rect 9119 32559 9153 32593
rect 9119 32491 9153 32525
rect 9119 32423 9153 32457
rect 9119 32355 9153 32389
rect 9119 32287 9153 32321
rect 9119 32219 9153 32253
rect 9119 32151 9153 32185
rect 9119 32083 9153 32117
rect 9119 32015 9153 32049
rect 9119 31947 9153 31981
rect 9119 31879 9153 31913
rect 9119 31811 9153 31845
rect 9119 31743 9153 31777
rect 9119 31675 9153 31709
rect 9119 31607 9153 31641
rect 9119 31539 9153 31573
rect 9119 31471 9153 31505
rect 9119 31403 9153 31437
rect 9119 31335 9153 31369
rect 9119 31267 9153 31301
rect 9789 31116 9823 31150
rect 9789 31048 9823 31082
rect 9789 30980 9823 31014
rect 9789 30912 9823 30946
rect 9789 30844 9823 30878
rect 9789 30776 9823 30810
rect 9789 30708 9823 30742
rect 9789 30640 9823 30674
rect 9789 30572 9823 30606
rect 9789 30504 9823 30538
rect 9789 30436 9823 30470
rect 9789 30368 9823 30402
rect 9789 30300 9823 30334
rect 9789 30232 9823 30266
rect 9789 30164 9823 30198
rect 9789 30096 9823 30130
rect 9789 30028 9823 30062
rect 9789 29960 9823 29994
rect 9789 29892 9823 29926
rect 9789 29824 9823 29858
rect 9789 29756 9823 29790
rect 9789 29688 9823 29722
rect 9789 29620 9823 29654
rect 9789 29552 9823 29586
rect 9789 29484 9823 29518
rect 9789 29416 9823 29450
rect 9789 29348 9823 29382
rect 9789 29280 9823 29314
rect 9789 29212 9823 29246
rect 9789 29144 9823 29178
rect 9789 29076 9823 29110
rect 9789 29008 9823 29042
rect 9789 28940 9823 28974
rect 9789 28872 9823 28906
rect 9789 28804 9823 28838
rect 9789 28736 9823 28770
rect 9789 28668 9823 28702
rect 9789 28600 9823 28634
rect 9789 28532 9823 28566
rect 9789 28464 9823 28498
rect 9789 28396 9823 28430
rect 9789 28328 9823 28362
rect 9789 28260 9823 28294
rect 9789 28192 9823 28226
rect 9789 28124 9823 28158
rect 9789 28056 9823 28090
rect 9789 27988 9823 28022
rect 9789 27920 9823 27954
rect 9789 27852 9823 27886
rect 9789 27784 9823 27818
rect 14405 34506 14439 34540
rect 14405 34438 14439 34472
rect 14405 34370 14439 34404
rect 14405 34302 14439 34336
rect 14405 34234 14439 34268
rect 14405 34166 14439 34200
rect 14405 34098 14439 34132
rect 14405 34030 14439 34064
rect 14405 33962 14439 33996
rect 14405 33894 14439 33928
rect 14405 33826 14439 33860
rect 14405 33758 14439 33792
rect 14405 33690 14439 33724
rect 14405 33622 14439 33656
rect 14405 33554 14439 33588
rect 14405 33486 14439 33520
rect 14405 33418 14439 33452
rect 14405 33350 14439 33384
rect 14405 33282 14439 33316
rect 14405 33214 14439 33248
rect 14405 33146 14439 33180
rect 14405 33078 14439 33112
rect 14405 33010 14439 33044
rect 14405 32942 14439 32976
rect 14405 32874 14439 32908
rect 14405 32806 14439 32840
rect 14405 32738 14439 32772
rect 14405 32670 14439 32704
rect 14405 32602 14439 32636
rect 14405 32534 14439 32568
rect 14405 32466 14439 32500
rect 14405 32398 14439 32432
rect 14405 32330 14439 32364
rect 14405 32262 14439 32296
rect 14405 32194 14439 32228
rect 14405 32126 14439 32160
rect 14405 32058 14439 32092
rect 14405 31990 14439 32024
rect 14405 31922 14439 31956
rect 14405 31854 14439 31888
rect 14405 31786 14439 31820
rect 14405 31718 14439 31752
rect 14405 31650 14439 31684
rect 14405 31582 14439 31616
rect 14405 31514 14439 31548
rect 14405 31446 14439 31480
rect 14405 31378 14439 31412
rect 14405 31310 14439 31344
rect 14405 31242 14439 31276
rect 14405 31174 14439 31208
rect 14405 31106 14439 31140
rect 14405 31038 14439 31072
rect 14405 30970 14439 31004
rect 14405 30902 14439 30936
rect 14405 30834 14439 30868
rect 14405 30766 14439 30800
rect 14405 30698 14439 30732
rect 14405 30630 14439 30664
rect 14405 30562 14439 30596
rect 14405 30494 14439 30528
rect 14405 30426 14439 30460
rect 14405 30358 14439 30392
rect 14405 30290 14439 30324
rect 14405 30222 14439 30256
rect 14405 30154 14439 30188
rect 14405 30086 14439 30120
rect 14405 30018 14439 30052
rect 14405 29950 14439 29984
rect 14405 29882 14439 29916
rect 14405 29814 14439 29848
rect 14405 29746 14439 29780
rect 14405 29678 14439 29712
rect 14405 29610 14439 29644
rect 14405 29542 14439 29576
rect 14405 29474 14439 29508
rect 14405 29406 14439 29440
rect 14405 29338 14439 29372
rect 14405 29270 14439 29304
rect 14405 29202 14439 29236
rect 14405 29134 14439 29168
rect 14405 29066 14439 29100
rect 14405 28998 14439 29032
rect 14405 28930 14439 28964
rect 14405 28862 14439 28896
rect 14405 28794 14439 28828
rect 14405 28726 14439 28760
rect 14405 28658 14439 28692
rect 14405 28590 14439 28624
rect 14405 28522 14439 28556
rect 14405 28454 14439 28488
rect 14405 28386 14439 28420
rect 14405 28318 14439 28352
rect 14405 28250 14439 28284
rect 14405 28182 14439 28216
rect 14405 28114 14439 28148
rect 14405 28046 14439 28080
rect 14405 27978 14439 28012
rect 14405 27910 14439 27944
rect 14405 27842 14439 27876
rect 14405 27774 14439 27808
rect 9789 27716 9823 27750
rect 9789 27648 9823 27682
rect 9789 27580 9823 27614
rect 9789 27512 9823 27546
rect 14405 27706 14439 27740
rect 14405 27638 14439 27672
rect 14405 27570 14439 27604
rect 9789 27444 9823 27478
rect 12500 27502 12534 27536
rect 12568 27502 12602 27536
rect 12636 27502 12670 27536
rect 12704 27502 12738 27536
rect 12772 27502 12806 27536
rect 12840 27502 12874 27536
rect 12908 27502 12942 27536
rect 12976 27502 13010 27536
rect 13044 27502 13078 27536
rect 13112 27502 13146 27536
rect 13180 27502 13214 27536
rect 13248 27502 13282 27536
rect 13316 27502 13350 27536
rect 13384 27502 13418 27536
rect 13452 27502 13486 27536
rect 13520 27502 13554 27536
rect 13588 27502 13622 27536
rect 13656 27502 13690 27536
rect 13724 27502 13758 27536
rect 13792 27502 13826 27536
rect 13860 27502 13894 27536
rect 13928 27502 13962 27536
rect 13996 27502 14030 27536
rect 14064 27502 14098 27536
rect 14132 27502 14166 27536
rect 14200 27502 14234 27536
rect 14268 27502 14302 27536
rect 14336 27502 14370 27536
rect 9789 27376 9823 27410
rect 9789 27308 9823 27342
rect 9789 27240 9823 27274
rect 9789 27172 9823 27206
rect 9789 27104 9823 27138
rect 9789 27036 9823 27070
rect 9789 26968 9823 27002
rect 9789 26900 9823 26934
rect 9789 26832 9823 26866
rect 9789 26764 9823 26798
rect 9789 26696 9823 26730
rect 12432 27390 12466 27424
rect 12432 27322 12466 27356
rect 12432 27254 12466 27288
rect 12432 27186 12466 27220
rect 12432 27118 12466 27152
rect 12432 27050 12466 27084
rect 12432 26982 12466 27016
rect 12432 26914 12466 26948
rect 12432 26846 12466 26880
rect 12432 26778 12466 26812
rect 12432 26710 12466 26744
rect 9789 26628 9823 26662
rect 9789 26560 9823 26594
rect 9789 26492 9823 26526
rect 12432 26642 12466 26676
rect 12432 26574 12466 26608
rect 12432 26506 12466 26540
rect 12432 26438 12466 26472
rect 9857 26370 9891 26404
rect 9925 26370 9959 26404
rect 9993 26370 10027 26404
rect 10061 26370 10095 26404
rect 10129 26370 10163 26404
rect 10197 26370 10231 26404
rect 10265 26370 10299 26404
rect 10333 26370 10367 26404
rect 10401 26370 10435 26404
rect 10469 26370 10503 26404
rect 10537 26370 10571 26404
rect 10605 26370 10639 26404
rect 10673 26370 10707 26404
rect 10741 26370 10775 26404
rect 10809 26370 10843 26404
rect 10877 26370 10911 26404
rect 10945 26370 10979 26404
rect 11013 26370 11047 26404
rect 11081 26370 11115 26404
rect 11149 26370 11183 26404
rect 11217 26370 11251 26404
rect 11285 26370 11319 26404
rect 11353 26370 11387 26404
rect 11421 26370 11455 26404
rect 11489 26370 11523 26404
rect 11557 26370 11591 26404
rect 11625 26370 11659 26404
rect 11693 26370 11727 26404
rect 11761 26370 11795 26404
rect 11829 26370 11863 26404
rect 11897 26370 11931 26404
rect 11965 26370 11999 26404
rect 12033 26370 12067 26404
rect 12101 26370 12135 26404
rect 12169 26370 12203 26404
rect 12237 26370 12271 26404
rect 12305 26370 12339 26404
<< mvpsubdiffcont >>
rect 5060 15746 5094 15780
rect 5140 15779 5174 15813
rect 5208 15779 5242 15813
rect 5276 15779 5310 15813
rect 5344 15779 5378 15813
rect 5412 15779 5446 15813
rect 5480 15779 5514 15813
rect 5548 15779 5582 15813
rect 5616 15779 5650 15813
rect 5060 15678 5094 15712
rect 5060 15610 5094 15644
rect 5060 15542 5094 15576
rect 5060 15474 5094 15508
rect 5060 15406 5094 15440
rect 5060 15338 5094 15372
rect 5060 15270 5094 15304
rect 5060 15202 5094 15236
rect 5060 15134 5094 15168
rect 5060 15066 5094 15100
rect 5649 15652 5683 15686
rect 5649 15584 5683 15618
rect 5649 15516 5683 15550
rect 5649 15448 5683 15482
rect 5649 15380 5683 15414
rect 5649 15312 5683 15346
rect 5649 15244 5683 15278
rect 5649 15176 5683 15210
rect 5649 15108 5683 15142
rect 5649 15040 5683 15074
rect 5093 14939 5127 14973
rect 5161 14939 5195 14973
rect 5229 14939 5263 14973
rect 5297 14939 5331 14973
rect 5365 14939 5399 14973
rect 5433 14939 5467 14973
rect 5501 14939 5535 14973
rect 5569 14939 5603 14973
rect 5649 14972 5683 15006
rect 5093 14824 5127 14858
rect 5161 14824 5195 14858
rect 5229 14824 5263 14858
rect 5297 14824 5331 14858
rect 5365 14824 5399 14858
rect 5433 14824 5467 14858
rect 5501 14824 5535 14858
rect 5569 14824 5603 14858
rect 5637 14824 5671 14858
rect 5705 14824 5739 14858
rect 5773 14824 5807 14858
rect 5841 14824 5875 14858
rect 5909 14824 5943 14858
rect 5977 14824 6011 14858
rect 6045 14824 6079 14858
rect 6113 14824 6147 14858
rect 6181 14824 6215 14858
rect 5060 14735 5094 14769
rect 6304 14791 6338 14825
rect 5060 14667 5094 14701
rect 5060 14599 5094 14633
rect 5060 14531 5094 14565
rect 5060 14463 5094 14497
rect 5060 14395 5094 14429
rect 5060 14327 5094 14361
rect 5060 14259 5094 14293
rect 5060 14191 5094 14225
rect 5060 14123 5094 14157
rect 5060 14055 5094 14089
rect 5060 13987 5094 14021
rect 5060 13919 5094 13953
rect 5060 13851 5094 13885
rect 5060 13783 5094 13817
rect 6304 14723 6338 14757
rect 6304 14655 6338 14689
rect 6304 14587 6338 14621
rect 6304 14519 6338 14553
rect 6304 14451 6338 14485
rect 6304 14383 6338 14417
rect 6304 14315 6338 14349
rect 6304 14247 6338 14281
rect 6304 14179 6338 14213
rect 6304 14111 6338 14145
rect 6304 14043 6338 14077
rect 6304 13975 6338 14009
rect 6304 13907 6338 13941
rect 6304 13839 6338 13873
rect 5060 13715 5094 13749
rect 5060 13647 5094 13681
rect 5060 13579 5094 13613
rect 5060 13511 5094 13545
rect 5060 13443 5094 13477
rect 5060 13375 5094 13409
rect 5060 13307 5094 13341
rect 5060 13239 5094 13273
rect 5060 13171 5094 13205
rect 5060 13103 5094 13137
rect 5060 13035 5094 13069
rect 5060 12967 5094 13001
rect 5060 12899 5094 12933
rect 5060 12831 5094 12865
rect 5060 12763 5094 12797
rect 5060 12695 5094 12729
rect 5060 12627 5094 12661
rect 5060 12559 5094 12593
rect 5060 12491 5094 12525
rect 5060 12423 5094 12457
rect 5060 12355 5094 12389
rect 5060 12287 5094 12321
rect 5060 12219 5094 12253
rect 5060 12151 5094 12185
rect 662 11892 696 11926
rect 662 11824 696 11858
rect 662 11756 696 11790
rect 662 11688 696 11722
rect 662 11620 696 11654
rect 662 11552 696 11586
rect 662 11484 696 11518
rect 662 11416 696 11450
rect 662 11348 696 11382
rect 662 11280 696 11314
rect 662 11212 696 11246
rect 662 11144 696 11178
rect 662 11076 696 11110
rect 662 11008 696 11042
rect 662 10940 696 10974
rect 662 10872 696 10906
rect 662 10804 696 10838
rect 662 10736 696 10770
rect 662 10668 696 10702
rect 662 10600 696 10634
rect 662 10532 696 10566
rect 662 10464 696 10498
rect 662 10396 696 10430
rect 662 10328 696 10362
rect 662 10260 696 10294
rect 662 10192 696 10226
rect 662 10124 696 10158
rect 662 10056 696 10090
rect 662 9988 696 10022
rect 2312 11825 2346 11859
rect 2312 11757 2346 11791
rect 2312 11689 2346 11723
rect 2312 11621 2346 11655
rect 2312 11553 2346 11587
rect 2312 11485 2346 11519
rect 2312 11417 2346 11451
rect 2312 11349 2346 11383
rect 2312 11281 2346 11315
rect 2312 11213 2346 11247
rect 2312 11145 2346 11179
rect 2312 11077 2346 11111
rect 2312 11009 2346 11043
rect 2312 10941 2346 10975
rect 2312 10873 2346 10907
rect 2312 10805 2346 10839
rect 2312 10737 2346 10771
rect 2312 10669 2346 10703
rect 2312 10601 2346 10635
rect 2312 10533 2346 10567
rect 2312 10465 2346 10499
rect 2312 10397 2346 10431
rect 2312 10329 2346 10363
rect 2312 10261 2346 10295
rect 2312 10193 2346 10227
rect 2312 10125 2346 10159
rect 2312 10057 2346 10091
rect 2312 9989 2346 10023
rect 2312 9921 2346 9955
rect 2690 11892 2724 11926
rect 2690 11824 2724 11858
rect 2690 11756 2724 11790
rect 2690 11688 2724 11722
rect 2690 11620 2724 11654
rect 2690 11552 2724 11586
rect 2690 11484 2724 11518
rect 2690 11416 2724 11450
rect 2690 11348 2724 11382
rect 2690 11280 2724 11314
rect 2690 11212 2724 11246
rect 2690 11144 2724 11178
rect 2690 11076 2724 11110
rect 2690 11008 2724 11042
rect 2690 10940 2724 10974
rect 2690 10872 2724 10906
rect 2690 10804 2724 10838
rect 2690 10736 2724 10770
rect 2690 10668 2724 10702
rect 2690 10600 2724 10634
rect 2690 10532 2724 10566
rect 2690 10464 2724 10498
rect 2690 10396 2724 10430
rect 2690 10328 2724 10362
rect 2690 10260 2724 10294
rect 2690 10192 2724 10226
rect 2690 10124 2724 10158
rect 2690 10056 2724 10090
rect 2690 9988 2724 10022
rect 4340 11825 4374 11859
rect 4340 11757 4374 11791
rect 4340 11689 4374 11723
rect 4340 11621 4374 11655
rect 4340 11553 4374 11587
rect 4340 11485 4374 11519
rect 4340 11417 4374 11451
rect 4340 11349 4374 11383
rect 4340 11281 4374 11315
rect 4340 11213 4374 11247
rect 4340 11145 4374 11179
rect 4340 11077 4374 11111
rect 4340 11009 4374 11043
rect 4340 10941 4374 10975
rect 4340 10873 4374 10907
rect 4340 10805 4374 10839
rect 4340 10737 4374 10771
rect 4340 10669 4374 10703
rect 4340 10601 4374 10635
rect 4340 10533 4374 10567
rect 4340 10465 4374 10499
rect 4340 10397 4374 10431
rect 4340 10329 4374 10363
rect 4340 10261 4374 10295
rect 4340 10193 4374 10227
rect 4340 10125 4374 10159
rect 4340 10057 4374 10091
rect 4340 9989 4374 10023
rect 4340 9921 4374 9955
rect 5060 12083 5094 12117
rect 5060 12015 5094 12049
rect 5060 11947 5094 11981
rect 5060 11879 5094 11913
rect 5060 11811 5094 11845
rect 5060 11743 5094 11777
rect 5060 11675 5094 11709
rect 5060 11607 5094 11641
rect 5060 11539 5094 11573
rect 5060 11471 5094 11505
rect 5060 11403 5094 11437
rect 5060 11335 5094 11369
rect 5060 11267 5094 11301
rect 5060 11199 5094 11233
rect 5060 11131 5094 11165
rect 5060 11063 5094 11097
rect 5060 10995 5094 11029
rect 5060 10927 5094 10961
rect 5060 10859 5094 10893
rect 5060 10791 5094 10825
rect 5060 10723 5094 10757
rect 5060 10655 5094 10689
rect 5060 10587 5094 10621
rect 5060 10519 5094 10553
rect 5060 10451 5094 10485
rect 5060 10383 5094 10417
rect 5060 10315 5094 10349
rect 5060 10247 5094 10281
rect 6304 13771 6338 13805
rect 6304 13703 6338 13737
rect 6304 13635 6338 13669
rect 6304 13567 6338 13601
rect 6304 13499 6338 13533
rect 6304 13431 6338 13465
rect 6304 13363 6338 13397
rect 6304 13295 6338 13329
rect 6304 13227 6338 13261
rect 6304 13159 6338 13193
rect 6304 13091 6338 13125
rect 6304 13023 6338 13057
rect 6304 12955 6338 12989
rect 6304 12887 6338 12921
rect 6304 12819 6338 12853
rect 6304 12751 6338 12785
rect 6304 12683 6338 12717
rect 6304 12615 6338 12649
rect 6304 12547 6338 12581
rect 6304 12479 6338 12513
rect 6304 12411 6338 12445
rect 6304 12343 6338 12377
rect 6304 12275 6338 12309
rect 6304 12207 6338 12241
rect 6304 12139 6338 12173
rect 6304 12071 6338 12105
rect 6304 12003 6338 12037
rect 6304 11935 6338 11969
rect 6304 11867 6338 11901
rect 6304 11799 6338 11833
rect 6304 11731 6338 11765
rect 6304 11663 6338 11697
rect 6304 11595 6338 11629
rect 6304 11527 6338 11561
rect 6304 11459 6338 11493
rect 6304 11391 6338 11425
rect 6304 11323 6338 11357
rect 6304 11255 6338 11289
rect 6304 11187 6338 11221
rect 6304 11119 6338 11153
rect 6304 11051 6338 11085
rect 6304 10938 6338 10972
rect 6304 10870 6338 10904
rect 6304 10802 6338 10836
rect 6304 10734 6338 10768
rect 6304 10666 6338 10700
rect 6304 10598 6338 10632
rect 6304 10530 6338 10564
rect 6304 10462 6338 10496
rect 6304 10394 6338 10428
rect 6304 10326 6338 10360
rect 6304 10258 6338 10292
rect 5060 10179 5094 10213
rect 6304 10190 6338 10224
rect 5060 10111 5094 10145
rect 5183 10078 5217 10112
rect 5251 10078 5285 10112
rect 5319 10078 5353 10112
rect 5387 10078 5421 10112
rect 5455 10078 5489 10112
rect 5523 10078 5557 10112
rect 5591 10078 5625 10112
rect 5659 10078 5693 10112
rect 5727 10078 5761 10112
rect 5795 10078 5829 10112
rect 5863 10078 5897 10112
rect 5931 10078 5965 10112
rect 5999 10078 6033 10112
rect 6067 10078 6101 10112
rect 6135 10078 6169 10112
rect 6203 10078 6237 10112
rect 6271 10078 6305 10112
rect 540 9477 574 9511
rect 632 9510 666 9544
rect 700 9510 734 9544
rect 768 9510 802 9544
rect 836 9510 870 9544
rect 904 9510 938 9544
rect 972 9510 1006 9544
rect 1040 9510 1074 9544
rect 1108 9510 1142 9544
rect 1176 9510 1210 9544
rect 1244 9510 1278 9544
rect 1312 9510 1346 9544
rect 1380 9510 1414 9544
rect 1448 9510 1482 9544
rect 1516 9510 1550 9544
rect 1584 9510 1618 9544
rect 1652 9510 1686 9544
rect 1720 9510 1754 9544
rect 1788 9510 1822 9544
rect 1856 9510 1890 9544
rect 1924 9510 1958 9544
rect 1992 9510 2026 9544
rect 2060 9510 2094 9544
rect 2128 9510 2162 9544
rect 2196 9510 2230 9544
rect 2264 9510 2298 9544
rect 2332 9510 2366 9544
rect 2400 9510 2434 9544
rect 2468 9510 2502 9544
rect 2576 9510 2610 9544
rect 2644 9510 2678 9544
rect 2712 9510 2746 9544
rect 2780 9510 2814 9544
rect 2848 9510 2882 9544
rect 2916 9510 2950 9544
rect 2984 9510 3018 9544
rect 3052 9510 3086 9544
rect 3120 9510 3154 9544
rect 3188 9510 3222 9544
rect 3256 9510 3290 9544
rect 3324 9510 3358 9544
rect 3426 9510 3460 9544
rect 3494 9510 3528 9544
rect 3562 9510 3596 9544
rect 3630 9510 3664 9544
rect 3698 9510 3732 9544
rect 3766 9510 3800 9544
rect 3834 9510 3868 9544
rect 3902 9510 3936 9544
rect 3970 9510 4004 9544
rect 4038 9510 4072 9544
rect 4106 9510 4140 9544
rect 4174 9510 4208 9544
rect 4242 9510 4276 9544
rect 4310 9510 4344 9544
rect 4378 9510 4412 9544
rect 4446 9510 4480 9544
rect 4514 9510 4548 9544
rect 4582 9510 4616 9544
rect 4650 9510 4684 9544
rect 4718 9510 4752 9544
rect 4786 9510 4820 9544
rect 4854 9510 4888 9544
rect 4922 9510 4956 9544
rect 4990 9510 5024 9544
rect 5058 9510 5092 9544
rect 5126 9510 5160 9544
rect 5194 9510 5228 9544
rect 5262 9510 5296 9544
rect 5330 9510 5364 9544
rect 5398 9510 5432 9544
rect 5466 9510 5500 9544
rect 5534 9510 5568 9544
rect 5602 9510 5636 9544
rect 5670 9510 5704 9544
rect 5738 9510 5772 9544
rect 540 9409 574 9443
rect 540 9341 574 9375
rect 540 9273 574 9307
rect 540 9205 574 9239
rect 540 9137 574 9171
rect 540 9069 574 9103
rect 540 9001 574 9035
rect 540 8933 574 8967
rect 540 8865 574 8899
rect 540 8797 574 8831
rect 540 8729 574 8763
rect 540 8661 574 8695
rect 540 8593 574 8627
rect 540 8525 574 8559
rect 540 8457 574 8491
rect 540 8389 574 8423
rect 540 8321 574 8355
rect 540 8253 574 8287
rect 540 8185 574 8219
rect 540 8117 574 8151
rect 540 8049 574 8083
rect 540 7981 574 8015
rect 540 7913 574 7947
rect 540 7845 574 7879
rect 540 7777 574 7811
rect 540 7709 574 7743
rect 540 7641 574 7675
rect 540 7573 574 7607
rect 540 7505 574 7539
rect 540 7437 574 7471
rect 540 7369 574 7403
rect 5830 9441 5864 9475
rect 3357 9362 3391 9396
rect 3357 9294 3391 9328
rect 3357 9226 3391 9260
rect 3357 9158 3391 9192
rect 3357 9090 3391 9124
rect 3357 9022 3391 9056
rect 3357 8954 3391 8988
rect 3357 8886 3391 8920
rect 3357 8818 3391 8852
rect 3357 8750 3391 8784
rect 3357 8682 3391 8716
rect 3357 8614 3391 8648
rect 3357 8546 3391 8580
rect 3357 8478 3391 8512
rect 3357 8410 3391 8444
rect 3357 8342 3391 8376
rect 3357 8274 3391 8308
rect 3357 8206 3391 8240
rect 3357 8138 3391 8172
rect 3357 8070 3391 8104
rect 3357 8002 3391 8036
rect 3357 7934 3391 7968
rect 3357 7866 3391 7900
rect 3357 7798 3391 7832
rect 3357 7730 3391 7764
rect 3357 7662 3391 7696
rect 3357 7594 3391 7628
rect 3357 7526 3391 7560
rect 3357 7458 3391 7492
rect 3357 7390 3391 7424
rect 3357 7322 3391 7356
rect 5830 9373 5864 9407
rect 5830 9305 5864 9339
rect 5830 9237 5864 9271
rect 5830 9169 5864 9203
rect 5830 9101 5864 9135
rect 5830 9033 5864 9067
rect 5830 8965 5864 8999
rect 5830 8897 5864 8931
rect 5830 8829 5864 8863
rect 5830 8761 5864 8795
rect 5830 8693 5864 8727
rect 5830 8625 5864 8659
rect 5830 8557 5864 8591
rect 5830 8489 5864 8523
rect 5830 8421 5864 8455
rect 5830 8353 5864 8387
rect 5830 8285 5864 8319
rect 5830 8217 5864 8251
rect 5830 8149 5864 8183
rect 5830 8081 5864 8115
rect 5830 8013 5864 8047
rect 5830 7945 5864 7979
rect 5830 7877 5864 7911
rect 5830 7809 5864 7843
rect 5830 7741 5864 7775
rect 5830 7673 5864 7707
rect 5830 7605 5864 7639
rect 5830 7537 5864 7571
rect 5830 7469 5864 7503
rect 5830 7401 5864 7435
rect 657 7253 691 7287
rect 741 7253 775 7287
rect 825 7253 859 7287
rect 909 7253 943 7287
rect 1261 7253 1295 7287
rect 1345 7253 1379 7287
rect 1429 7253 1463 7287
rect 1513 7253 1547 7287
rect 1597 7253 1631 7287
rect 1681 7253 1715 7287
rect 1765 7253 1799 7287
rect 2117 7253 2151 7287
rect 2201 7253 2235 7287
rect 2285 7253 2319 7287
rect 2369 7253 2403 7287
rect 2453 7253 2487 7287
rect 2537 7253 2571 7287
rect 2621 7253 2655 7287
rect 5830 7333 5864 7367
rect 2973 7253 3007 7287
rect 3057 7253 3091 7287
rect 3141 7253 3175 7287
rect 3225 7253 3259 7287
rect 3357 7254 3391 7288
rect 3489 7253 3523 7287
rect 3573 7253 3607 7287
rect 3657 7253 3691 7287
rect 3741 7253 3775 7287
rect 4093 7253 4127 7287
rect 4177 7253 4211 7287
rect 4261 7253 4295 7287
rect 4345 7253 4379 7287
rect 4801 7253 4835 7287
rect 5257 7253 5291 7287
rect 5713 7253 5747 7287
rect 5830 7265 5864 7299
rect 540 7217 574 7251
rect 540 7149 574 7183
rect 540 7081 574 7115
rect 540 7013 574 7047
rect 540 6945 574 6979
rect 540 6877 574 6911
rect 540 6809 574 6843
rect 540 6741 574 6775
rect 540 6673 574 6707
rect 540 6605 574 6639
rect 540 6537 574 6571
rect 540 6469 574 6503
rect 540 6401 574 6435
rect 540 6333 574 6367
rect 540 6265 574 6299
rect 540 6197 574 6231
rect 540 6129 574 6163
rect 540 6061 574 6095
rect 540 5993 574 6027
rect 540 5925 574 5959
rect 540 5857 574 5891
rect 540 5789 574 5823
rect 540 5721 574 5755
rect 540 5653 574 5687
rect 540 5585 574 5619
rect 540 5517 574 5551
rect 540 5449 574 5483
rect 540 5381 574 5415
rect 540 5313 574 5347
rect 540 5245 574 5279
rect 540 5177 574 5211
rect 3357 7186 3391 7220
rect 5830 7197 5864 7231
rect 3357 7118 3391 7152
rect 3357 7050 3391 7084
rect 3357 6982 3391 7016
rect 3357 6914 3391 6948
rect 3357 6846 3391 6880
rect 3357 6778 3391 6812
rect 3357 6710 3391 6744
rect 3357 6642 3391 6676
rect 3357 6574 3391 6608
rect 3357 6506 3391 6540
rect 3357 6438 3391 6472
rect 3357 6370 3391 6404
rect 3357 6302 3391 6336
rect 3357 6234 3391 6268
rect 3357 6166 3391 6200
rect 3357 6098 3391 6132
rect 3357 6030 3391 6064
rect 3357 5962 3391 5996
rect 3357 5894 3391 5928
rect 3357 5826 3391 5860
rect 3357 5758 3391 5792
rect 3357 5690 3391 5724
rect 3357 5622 3391 5656
rect 3357 5554 3391 5588
rect 3357 5486 3391 5520
rect 3357 5418 3391 5452
rect 3357 5350 3391 5384
rect 3357 5282 3391 5316
rect 3357 5214 3391 5248
rect 3357 5146 3391 5180
rect 5830 7129 5864 7163
rect 5830 7061 5864 7095
rect 5830 6993 5864 7027
rect 5830 6925 5864 6959
rect 5830 6857 5864 6891
rect 5830 6789 5864 6823
rect 5830 6721 5864 6755
rect 5830 6653 5864 6687
rect 5830 6585 5864 6619
rect 5830 6517 5864 6551
rect 5830 6449 5864 6483
rect 5830 6381 5864 6415
rect 5830 6313 5864 6347
rect 5830 6245 5864 6279
rect 5830 6177 5864 6211
rect 5830 6109 5864 6143
rect 5830 6041 5864 6075
rect 5830 5973 5864 6007
rect 5830 5905 5864 5939
rect 5830 5837 5864 5871
rect 5830 5769 5864 5803
rect 5830 5701 5864 5735
rect 5830 5633 5864 5667
rect 5830 5565 5864 5599
rect 5830 5497 5864 5531
rect 5830 5429 5864 5463
rect 5830 5361 5864 5395
rect 5830 5293 5864 5327
rect 5830 5225 5864 5259
rect 5830 5157 5864 5191
rect 540 5014 574 5048
rect 657 5033 691 5067
rect 741 5033 775 5067
rect 825 5033 859 5067
rect 909 5033 943 5067
rect 1261 5033 1295 5067
rect 1345 5033 1379 5067
rect 1429 5033 1463 5067
rect 1513 5033 1547 5067
rect 1597 5033 1631 5067
rect 1681 5033 1715 5067
rect 1765 5033 1799 5067
rect 2117 5033 2151 5067
rect 2201 5033 2235 5067
rect 2285 5033 2319 5067
rect 2369 5033 2403 5067
rect 2453 5033 2487 5067
rect 2537 5033 2571 5067
rect 2621 5033 2655 5067
rect 3357 5078 3391 5112
rect 5830 5089 5864 5123
rect 2973 5033 3007 5067
rect 3057 5033 3091 5067
rect 3141 5033 3175 5067
rect 3225 5033 3259 5067
rect 540 4946 574 4980
rect 3357 5010 3391 5044
rect 3489 5033 3523 5067
rect 3573 5033 3607 5067
rect 3657 5033 3691 5067
rect 3741 5033 3775 5067
rect 4093 5033 4127 5067
rect 4177 5033 4211 5067
rect 4261 5033 4295 5067
rect 4345 5033 4379 5067
rect 4801 5033 4835 5067
rect 5257 5033 5291 5067
rect 5713 5033 5747 5067
rect 5830 5021 5864 5055
rect 540 4878 574 4912
rect 540 4810 574 4844
rect 540 4742 574 4776
rect 540 4674 574 4708
rect 540 4606 574 4640
rect 540 4538 574 4572
rect 540 4470 574 4504
rect 540 4402 574 4436
rect 540 4334 574 4368
rect 540 4266 574 4300
rect 540 4198 574 4232
rect 540 4130 574 4164
rect 540 4062 574 4096
rect 540 3994 574 4028
rect 540 3926 574 3960
rect 540 3858 574 3892
rect 540 3790 574 3824
rect 540 3722 574 3756
rect 540 3654 574 3688
rect 540 3586 574 3620
rect 540 3518 574 3552
rect 540 3450 574 3484
rect 540 3382 574 3416
rect 540 3314 574 3348
rect 540 3246 574 3280
rect 540 3178 574 3212
rect 540 3110 574 3144
rect 540 3042 574 3076
rect 540 2974 574 3008
rect 540 2906 574 2940
rect 3357 4942 3391 4976
rect 3357 4874 3391 4908
rect 3357 4806 3391 4840
rect 3357 4738 3391 4772
rect 3357 4670 3391 4704
rect 3357 4602 3391 4636
rect 3357 4534 3391 4568
rect 3357 4466 3391 4500
rect 3357 4398 3391 4432
rect 3357 4330 3391 4364
rect 3357 4262 3391 4296
rect 3357 4194 3391 4228
rect 3357 4126 3391 4160
rect 3357 4058 3391 4092
rect 3357 3990 3391 4024
rect 3357 3922 3391 3956
rect 3357 3854 3391 3888
rect 3357 3786 3391 3820
rect 3357 3718 3391 3752
rect 3357 3650 3391 3684
rect 3357 3582 3391 3616
rect 3357 3514 3391 3548
rect 3357 3446 3391 3480
rect 3357 3378 3391 3412
rect 3357 3310 3391 3344
rect 3357 3242 3391 3276
rect 3357 3174 3391 3208
rect 3357 3106 3391 3140
rect 3357 3038 3391 3072
rect 3357 2970 3391 3004
rect 540 2838 574 2872
rect 3357 2902 3391 2936
rect 5830 4953 5864 4987
rect 5830 4885 5864 4919
rect 5830 4817 5864 4851
rect 5830 4749 5864 4783
rect 5830 4681 5864 4715
rect 5830 4613 5864 4647
rect 5830 4545 5864 4579
rect 5830 4477 5864 4511
rect 5830 4409 5864 4443
rect 5830 4341 5864 4375
rect 5830 4273 5864 4307
rect 5830 4205 5864 4239
rect 5830 4137 5864 4171
rect 5830 4069 5864 4103
rect 5830 4001 5864 4035
rect 5830 3933 5864 3967
rect 5830 3865 5864 3899
rect 5830 3797 5864 3831
rect 5830 3729 5864 3763
rect 5830 3661 5864 3695
rect 5830 3593 5864 3627
rect 5830 3525 5864 3559
rect 5830 3457 5864 3491
rect 5830 3389 5864 3423
rect 5830 3321 5864 3355
rect 5830 3253 5864 3287
rect 5830 3185 5864 3219
rect 5830 3117 5864 3151
rect 5830 3049 5864 3083
rect 5830 2981 5864 3015
rect 5830 2913 5864 2947
rect 657 2814 691 2848
rect 741 2814 775 2848
rect 825 2814 859 2848
rect 909 2814 943 2848
rect 1261 2814 1295 2848
rect 1345 2814 1379 2848
rect 1429 2814 1463 2848
rect 1513 2814 1547 2848
rect 1597 2814 1631 2848
rect 1681 2814 1715 2848
rect 1765 2814 1799 2848
rect 2117 2814 2151 2848
rect 2201 2814 2235 2848
rect 2285 2814 2319 2848
rect 2369 2814 2403 2848
rect 2453 2814 2487 2848
rect 2537 2814 2571 2848
rect 2621 2814 2655 2848
rect 2973 2814 3007 2848
rect 3057 2814 3091 2848
rect 3141 2814 3175 2848
rect 3225 2814 3259 2848
rect 3357 2834 3391 2868
rect 3489 2814 3523 2848
rect 3573 2814 3607 2848
rect 3657 2814 3691 2848
rect 3741 2814 3775 2848
rect 4093 2814 4127 2848
rect 4177 2814 4211 2848
rect 4261 2814 4295 2848
rect 4345 2814 4379 2848
rect 4801 2814 4835 2848
rect 5257 2814 5291 2848
rect 5713 2814 5747 2848
rect 5830 2845 5864 2879
rect 540 2770 574 2804
rect 3357 2766 3391 2800
rect 540 2702 574 2736
rect 540 2550 574 2584
rect 540 2482 574 2516
rect 540 2414 574 2448
rect 540 2346 574 2380
rect 540 2278 574 2312
rect 540 2210 574 2244
rect 540 2142 574 2176
rect 540 2074 574 2108
rect 540 2006 574 2040
rect 540 1938 574 1972
rect 540 1870 574 1904
rect 540 1802 574 1836
rect 540 1734 574 1768
rect 540 1666 574 1700
rect 540 1598 574 1632
rect 540 1530 574 1564
rect 540 1462 574 1496
rect 540 1394 574 1428
rect 540 1326 574 1360
rect 540 1258 574 1292
rect 540 1190 574 1224
rect 540 1122 574 1156
rect 540 1054 574 1088
rect 540 986 574 1020
rect 540 918 574 952
rect 540 850 574 884
rect 540 782 574 816
rect 540 714 574 748
rect 5830 2777 5864 2811
rect 3357 2698 3391 2732
rect 3357 2630 3391 2664
rect 3357 2562 3391 2596
rect 3357 2494 3391 2528
rect 3357 2426 3391 2460
rect 3357 2358 3391 2392
rect 3357 2290 3391 2324
rect 3357 2222 3391 2256
rect 3357 2154 3391 2188
rect 3357 2086 3391 2120
rect 3357 2018 3391 2052
rect 3357 1950 3391 1984
rect 3357 1882 3391 1916
rect 3357 1814 3391 1848
rect 3357 1746 3391 1780
rect 3357 1678 3391 1712
rect 3357 1610 3391 1644
rect 3357 1542 3391 1576
rect 3357 1474 3391 1508
rect 3357 1406 3391 1440
rect 3357 1338 3391 1372
rect 3357 1270 3391 1304
rect 3357 1202 3391 1236
rect 3357 1134 3391 1168
rect 3357 1066 3391 1100
rect 3357 998 3391 1032
rect 3357 930 3391 964
rect 3357 862 3391 896
rect 3357 794 3391 828
rect 3357 726 3391 760
rect 5830 2709 5864 2743
rect 5830 2641 5864 2675
rect 5830 2573 5864 2607
rect 5830 2505 5864 2539
rect 5830 2437 5864 2471
rect 5830 2369 5864 2403
rect 5830 2301 5864 2335
rect 5830 2233 5864 2267
rect 5830 2165 5864 2199
rect 5830 2097 5864 2131
rect 5830 2029 5864 2063
rect 5830 1961 5864 1995
rect 5830 1893 5864 1927
rect 5830 1825 5864 1859
rect 5830 1757 5864 1791
rect 5830 1689 5864 1723
rect 5830 1621 5864 1655
rect 5830 1553 5864 1587
rect 5830 1485 5864 1519
rect 5830 1417 5864 1451
rect 5830 1349 5864 1383
rect 5830 1281 5864 1315
rect 5830 1213 5864 1247
rect 5830 1145 5864 1179
rect 5830 1077 5864 1111
rect 5830 1009 5864 1043
rect 5830 941 5864 975
rect 5830 873 5864 907
rect 5830 805 5864 839
rect 5830 737 5864 771
rect 3357 658 3391 692
rect 5830 669 5864 703
rect 573 557 607 591
rect 641 557 675 591
rect 709 557 743 591
rect 777 557 811 591
rect 845 557 879 591
rect 913 557 947 591
rect 1253 557 1287 591
rect 1321 557 1355 591
rect 1389 557 1423 591
rect 1457 557 1491 591
rect 1525 557 1559 591
rect 1593 557 1627 591
rect 1661 557 1695 591
rect 1729 557 1763 591
rect 1797 557 1831 591
rect 1865 557 1899 591
rect 2205 557 2239 591
rect 2273 557 2307 591
rect 2341 557 2375 591
rect 2409 557 2443 591
rect 2559 557 2593 591
rect 2627 557 2661 591
rect 2695 557 2729 591
rect 2763 557 2797 591
rect 2831 557 2865 591
rect 3152 557 3186 591
rect 3220 557 3254 591
rect 3288 557 3322 591
rect 3357 590 3391 624
rect 3426 557 3460 591
rect 3494 557 3528 591
rect 3562 557 3596 591
rect 3630 557 3664 591
rect 3979 557 4013 591
rect 4047 557 4081 591
rect 4115 557 4149 591
rect 4183 557 4217 591
rect 4251 557 4285 591
rect 4319 557 4353 591
rect 4639 557 4673 591
rect 4707 557 4741 591
rect 4775 557 4809 591
rect 5109 557 5143 591
rect 5177 557 5211 591
rect 5457 557 5491 591
rect 5525 557 5559 591
rect 5593 557 5627 591
rect 5661 557 5695 591
rect 5729 557 5763 591
rect 5797 557 5831 591
<< mvnsubdiffcont >>
rect 176 17309 210 17343
rect 244 17309 278 17343
rect 312 17309 346 17343
rect 380 17309 414 17343
rect 448 17309 482 17343
rect 516 17309 550 17343
rect 584 17309 618 17343
rect 652 17309 686 17343
rect 720 17309 754 17343
rect 788 17309 822 17343
rect 856 17309 890 17343
rect 924 17309 958 17343
rect 992 17309 1026 17343
rect 1060 17309 1094 17343
rect 1128 17309 1162 17343
rect 1196 17309 1230 17343
rect 1264 17309 1298 17343
rect 1332 17309 1366 17343
rect 1400 17309 1434 17343
rect 1468 17309 1502 17343
rect 1536 17309 1570 17343
rect 1604 17309 1638 17343
rect 1672 17309 1706 17343
rect 1740 17309 1774 17343
rect 1808 17309 1842 17343
rect 1876 17309 1910 17343
rect 1944 17309 1978 17343
rect 2012 17309 2046 17343
rect 2080 17309 2114 17343
rect 2148 17309 2182 17343
rect 2235 17215 2269 17249
rect 2235 17147 2269 17181
rect 2235 17079 2269 17113
rect 2235 17011 2269 17045
rect 2235 16943 2269 16977
rect 234 16874 268 16908
rect 302 16874 336 16908
rect 714 16874 748 16908
rect 836 16874 870 16908
rect 904 16874 938 16908
rect 972 16874 1006 16908
rect 1040 16874 1074 16908
rect 1108 16874 1142 16908
rect 1176 16874 1210 16908
rect 1244 16874 1278 16908
rect 1312 16874 1346 16908
rect 1380 16874 1414 16908
rect 1448 16874 1482 16908
rect 1516 16874 1550 16908
rect 1584 16874 1618 16908
rect 1652 16874 1686 16908
rect 1720 16874 1754 16908
rect 1788 16874 1822 16908
rect 1856 16874 1890 16908
rect 1924 16874 1958 16908
rect 1992 16874 2026 16908
rect 2060 16874 2094 16908
rect 2128 16874 2162 16908
rect 2196 16874 2230 16908
rect 2264 16874 2298 16908
rect 2332 16874 2366 16908
rect 2400 16874 2434 16908
rect 2468 16874 2502 16908
rect 2570 16874 2604 16908
rect 2638 16874 2672 16908
rect 2706 16874 2740 16908
rect 2774 16874 2808 16908
rect 2842 16874 2876 16908
rect 2910 16874 2944 16908
rect 2978 16874 3012 16908
rect 3046 16874 3080 16908
rect 3114 16874 3148 16908
rect 3182 16874 3216 16908
rect 3250 16874 3284 16908
rect 3318 16874 3352 16908
rect 3386 16874 3420 16908
rect 3454 16874 3488 16908
rect 3522 16874 3556 16908
rect 3590 16874 3624 16908
rect 3658 16874 3692 16908
rect 3726 16874 3760 16908
rect 3794 16874 3828 16908
rect 3862 16874 3896 16908
rect 3930 16874 3964 16908
rect 3998 16874 4032 16908
rect 4066 16874 4100 16908
rect 4134 16874 4168 16908
rect 4202 16874 4236 16908
rect 4270 16874 4304 16908
rect 4338 16874 4372 16908
rect 4406 16874 4440 16908
rect 4474 16874 4508 16908
rect 4542 16874 4576 16908
rect 4610 16874 4644 16908
rect 4678 16874 4712 16908
rect 4746 16874 4780 16908
rect 4871 16841 4905 16875
rect 2501 16771 2535 16805
rect 4871 16773 4905 16807
rect 2501 16703 2535 16737
rect 2501 16635 2535 16669
rect 2501 16567 2535 16601
rect 2501 16499 2535 16533
rect 2501 16431 2535 16465
rect 2501 16363 2535 16397
rect 2501 16295 2535 16329
rect 2501 16227 2535 16261
rect 2501 16159 2535 16193
rect 2501 16091 2535 16125
rect 2501 16023 2535 16057
rect 2501 15955 2535 15989
rect 2501 15887 2535 15921
rect 2501 15819 2535 15853
rect 2501 15751 2535 15785
rect 2501 15683 2535 15717
rect 2501 15615 2535 15649
rect 2501 15547 2535 15581
rect 2501 15479 2535 15513
rect 2501 15411 2535 15445
rect 2501 15343 2535 15377
rect 4871 16705 4905 16739
rect 4871 16637 4905 16671
rect 4871 16569 4905 16603
rect 4871 16501 4905 16535
rect 4871 16433 4905 16467
rect 4871 16365 4905 16399
rect 4871 16297 4905 16331
rect 4871 16229 4905 16263
rect 4871 16161 4905 16195
rect 4871 16093 4905 16127
rect 4871 16025 4905 16059
rect 4871 15957 4905 15991
rect 4871 15889 4905 15923
rect 4871 15821 4905 15855
rect 4871 15753 4905 15787
rect 4871 15685 4905 15719
rect 4871 15617 4905 15651
rect 4871 15549 4905 15583
rect 4871 15481 4905 15515
rect 4871 15413 4905 15447
rect 4871 15345 4905 15379
rect 2501 15275 2535 15309
rect 2501 15207 2535 15241
rect 4871 15277 4905 15311
rect 2501 15139 2535 15173
rect 2501 15071 2535 15105
rect 2501 15003 2535 15037
rect 2501 14935 2535 14969
rect 2501 14867 2535 14901
rect 2501 14799 2535 14833
rect 2501 14731 2535 14765
rect 2501 14663 2535 14697
rect 2501 14595 2535 14629
rect 2501 14527 2535 14561
rect 2501 14459 2535 14493
rect 2501 14391 2535 14425
rect 2501 14323 2535 14357
rect 2501 14255 2535 14289
rect 2501 14187 2535 14221
rect 2501 14119 2535 14153
rect 2501 14051 2535 14085
rect 2501 13983 2535 14017
rect 2501 13915 2535 13949
rect 2501 13847 2535 13881
rect 2501 13779 2535 13813
rect 4871 15209 4905 15243
rect 4871 15141 4905 15175
rect 4871 15073 4905 15107
rect 4871 15005 4905 15039
rect 4871 14937 4905 14971
rect 4871 14869 4905 14903
rect 4871 14801 4905 14835
rect 4871 14733 4905 14767
rect 4871 14665 4905 14699
rect 4871 14597 4905 14631
rect 4871 14529 4905 14563
rect 4871 14461 4905 14495
rect 4871 14393 4905 14427
rect 4871 14325 4905 14359
rect 4871 14257 4905 14291
rect 4871 14189 4905 14223
rect 4871 14121 4905 14155
rect 4871 14053 4905 14087
rect 4871 13985 4905 14019
rect 4871 13917 4905 13951
rect 4871 13849 4905 13883
rect 2501 13711 2535 13745
rect 4871 13781 4905 13815
rect 4871 13713 4905 13747
rect 2501 13643 2535 13677
rect 2501 13575 2535 13609
rect 2501 13507 2535 13541
rect 2501 13439 2535 13473
rect 2501 13371 2535 13405
rect 2501 13303 2535 13337
rect 2501 13235 2535 13269
rect 2501 13167 2535 13201
rect 2501 13099 2535 13133
rect 2501 13031 2535 13065
rect 2501 12963 2535 12997
rect 2501 12895 2535 12929
rect 2501 12827 2535 12861
rect 2501 12759 2535 12793
rect 2501 12691 2535 12725
rect 2501 12623 2535 12657
rect 2501 12555 2535 12589
rect 2501 12487 2535 12521
rect 2501 12419 2535 12453
rect 2501 12351 2535 12385
rect 2501 12283 2535 12317
rect 4871 13645 4905 13679
rect 4871 13577 4905 13611
rect 4871 13509 4905 13543
rect 4871 13441 4905 13475
rect 4871 13373 4905 13407
rect 4871 13305 4905 13339
rect 4871 13237 4905 13271
rect 4871 13169 4905 13203
rect 4871 13101 4905 13135
rect 4871 13033 4905 13067
rect 4871 12965 4905 12999
rect 4871 12897 4905 12931
rect 4871 12829 4905 12863
rect 4871 12761 4905 12795
rect 4871 12693 4905 12727
rect 4871 12625 4905 12659
rect 4871 12557 4905 12591
rect 4871 12489 4905 12523
rect 4871 12421 4905 12455
rect 4871 12353 4905 12387
rect 4871 12285 4905 12319
rect 2501 12215 2535 12249
rect 291 12114 325 12148
rect 359 12114 393 12148
rect 427 12114 461 12148
rect 495 12114 529 12148
rect 563 12114 597 12148
rect 631 12114 665 12148
rect 699 12114 733 12148
rect 767 12114 801 12148
rect 835 12114 869 12148
rect 903 12114 937 12148
rect 971 12114 1005 12148
rect 1039 12114 1073 12148
rect 1107 12114 1141 12148
rect 1175 12114 1209 12148
rect 1243 12114 1277 12148
rect 1311 12114 1345 12148
rect 1379 12114 1413 12148
rect 1447 12114 1481 12148
rect 1515 12114 1549 12148
rect 1583 12114 1617 12148
rect 1651 12114 1685 12148
rect 1719 12114 1753 12148
rect 1787 12114 1821 12148
rect 1855 12114 1889 12148
rect 1923 12114 1957 12148
rect 1991 12114 2025 12148
rect 2059 12114 2093 12148
rect 2127 12114 2161 12148
rect 2195 12114 2229 12148
rect 2263 12114 2297 12148
rect 2331 12114 2365 12148
rect 2399 12114 2433 12148
rect 2501 12147 2535 12181
rect 4871 12148 4905 12182
rect 2596 12114 2630 12148
rect 2664 12114 2698 12148
rect 2732 12114 2766 12148
rect 2800 12114 2834 12148
rect 2868 12114 2902 12148
rect 2936 12114 2970 12148
rect 3004 12114 3038 12148
rect 3072 12114 3106 12148
rect 3140 12114 3174 12148
rect 3208 12114 3242 12148
rect 3276 12114 3310 12148
rect 3344 12114 3378 12148
rect 3412 12114 3446 12148
rect 3480 12114 3514 12148
rect 3548 12114 3582 12148
rect 3616 12114 3650 12148
rect 3684 12114 3718 12148
rect 3752 12114 3786 12148
rect 3820 12114 3854 12148
rect 3888 12114 3922 12148
rect 3956 12114 3990 12148
rect 4024 12114 4058 12148
rect 4092 12114 4126 12148
rect 4160 12114 4194 12148
rect 4228 12114 4262 12148
rect 4296 12114 4330 12148
rect 4364 12114 4398 12148
rect 4432 12114 4466 12148
rect 4500 12114 4534 12148
rect 4568 12114 4602 12148
rect 4636 12114 4670 12148
rect 4704 12114 4738 12148
rect 4772 12114 4806 12148
rect 351 12045 385 12079
rect 472 12045 506 12079
rect 2501 12044 2535 12078
rect 351 11977 385 12011
rect 472 11977 506 12011
rect 351 11909 385 11943
rect 472 11909 506 11943
rect 351 11841 385 11875
rect 472 11841 506 11875
rect 351 11773 385 11807
rect 472 11773 506 11807
rect 351 11705 385 11739
rect 472 11705 506 11739
rect 351 11637 385 11671
rect 472 11637 506 11671
rect 351 11569 385 11603
rect 472 11569 506 11603
rect 351 11501 385 11535
rect 472 11501 506 11535
rect 351 11433 385 11467
rect 472 11433 506 11467
rect 351 11365 385 11399
rect 472 11365 506 11399
rect 351 11297 385 11331
rect 472 11297 506 11331
rect 351 11229 385 11263
rect 472 11229 506 11263
rect 351 11161 385 11195
rect 472 11161 506 11195
rect 351 11093 385 11127
rect 472 11093 506 11127
rect 351 11025 385 11059
rect 472 11025 506 11059
rect 351 10957 385 10991
rect 472 10957 506 10991
rect 351 10889 385 10923
rect 472 10889 506 10923
rect 351 10821 385 10855
rect 472 10821 506 10855
rect 351 10753 385 10787
rect 472 10753 506 10787
rect 351 10685 385 10719
rect 472 10685 506 10719
rect 351 10617 385 10651
rect 472 10617 506 10651
rect 351 10549 385 10583
rect 472 10549 506 10583
rect 351 10481 385 10515
rect 472 10481 506 10515
rect 351 10413 385 10447
rect 472 10413 506 10447
rect 351 10345 385 10379
rect 472 10345 506 10379
rect 351 10277 385 10311
rect 472 10277 506 10311
rect 351 10209 385 10243
rect 472 10209 506 10243
rect 351 10141 385 10175
rect 472 10141 506 10175
rect 351 10073 385 10107
rect 472 10073 506 10107
rect 351 10005 385 10039
rect 472 10005 506 10039
rect 351 9937 385 9971
rect 472 9937 506 9971
rect 351 9869 385 9903
rect 472 9869 506 9903
rect 4529 12045 4563 12079
rect 4651 12044 4685 12078
rect 2501 11976 2535 12010
rect 351 9801 385 9835
rect 472 9801 506 9835
rect 2501 11908 2535 11942
rect 2501 11840 2535 11874
rect 2501 11772 2535 11806
rect 2501 11704 2535 11738
rect 2501 11636 2535 11670
rect 2501 11568 2535 11602
rect 2501 11500 2535 11534
rect 2501 11432 2535 11466
rect 2501 11364 2535 11398
rect 2501 11296 2535 11330
rect 2501 11228 2535 11262
rect 2501 11160 2535 11194
rect 2501 11092 2535 11126
rect 2501 11024 2535 11058
rect 2501 10956 2535 10990
rect 2501 10888 2535 10922
rect 2501 10820 2535 10854
rect 2501 10752 2535 10786
rect 2501 10684 2535 10718
rect 2501 10616 2535 10650
rect 2501 10548 2535 10582
rect 2501 10480 2535 10514
rect 2501 10412 2535 10446
rect 2501 10344 2535 10378
rect 2501 10276 2535 10310
rect 2501 10208 2535 10242
rect 2501 10140 2535 10174
rect 2501 10072 2535 10106
rect 2501 10004 2535 10038
rect 2501 9936 2535 9970
rect 2501 9868 2535 9902
rect 4529 11977 4563 12011
rect 4651 11976 4685 12010
rect 351 9733 385 9767
rect 472 9733 506 9767
rect 2501 9800 2535 9834
rect 4529 11909 4563 11943
rect 4651 11908 4685 11942
rect 4529 11841 4563 11875
rect 4651 11840 4685 11874
rect 4529 11773 4563 11807
rect 4651 11772 4685 11806
rect 4529 11705 4563 11739
rect 4651 11704 4685 11738
rect 4529 11637 4563 11671
rect 4651 11636 4685 11670
rect 4529 11569 4563 11603
rect 4651 11568 4685 11602
rect 4529 11501 4563 11535
rect 4651 11500 4685 11534
rect 4529 11433 4563 11467
rect 4651 11432 4685 11466
rect 4529 11365 4563 11399
rect 4651 11364 4685 11398
rect 4529 11297 4563 11331
rect 4651 11296 4685 11330
rect 4529 11229 4563 11263
rect 4651 11228 4685 11262
rect 4529 11161 4563 11195
rect 4651 11160 4685 11194
rect 4529 11093 4563 11127
rect 4651 11092 4685 11126
rect 4529 11025 4563 11059
rect 4651 11024 4685 11058
rect 4529 10957 4563 10991
rect 4651 10956 4685 10990
rect 4529 10889 4563 10923
rect 4651 10888 4685 10922
rect 4529 10821 4563 10855
rect 4651 10820 4685 10854
rect 4529 10753 4563 10787
rect 4651 10752 4685 10786
rect 4529 10685 4563 10719
rect 4651 10684 4685 10718
rect 4529 10617 4563 10651
rect 4651 10616 4685 10650
rect 4529 10549 4563 10583
rect 4651 10548 4685 10582
rect 4529 10481 4563 10515
rect 4651 10480 4685 10514
rect 4529 10413 4563 10447
rect 4651 10412 4685 10446
rect 4529 10345 4563 10379
rect 4651 10344 4685 10378
rect 4529 10277 4563 10311
rect 4651 10276 4685 10310
rect 4529 10209 4563 10243
rect 4651 10208 4685 10242
rect 4529 10141 4563 10175
rect 4651 10140 4685 10174
rect 4529 10073 4563 10107
rect 4651 10072 4685 10106
rect 4529 10005 4563 10039
rect 4651 10004 4685 10038
rect 4529 9937 4563 9971
rect 4651 9936 4685 9970
rect 4529 9869 4563 9903
rect 4651 9868 4685 9902
rect 710 9699 744 9733
rect 778 9699 812 9733
rect 846 9699 880 9733
rect 914 9699 948 9733
rect 982 9699 1016 9733
rect 1050 9699 1084 9733
rect 1118 9699 1152 9733
rect 1186 9699 1220 9733
rect 1254 9699 1288 9733
rect 1322 9699 1356 9733
rect 1390 9699 1424 9733
rect 1458 9699 1492 9733
rect 1526 9699 1560 9733
rect 1594 9699 1628 9733
rect 1662 9699 1696 9733
rect 1730 9699 1764 9733
rect 1798 9699 1832 9733
rect 1866 9699 1900 9733
rect 1934 9699 1968 9733
rect 2002 9699 2036 9733
rect 2070 9699 2104 9733
rect 2138 9699 2172 9733
rect 2206 9699 2240 9733
rect 2274 9699 2308 9733
rect 2501 9732 2535 9766
rect 4529 9801 4563 9835
rect 4651 9800 4685 9834
rect 4529 9733 4563 9767
rect 2728 9699 2762 9733
rect 2796 9699 2830 9733
rect 2864 9699 2898 9733
rect 2932 9699 2966 9733
rect 3000 9699 3034 9733
rect 3068 9699 3102 9733
rect 3136 9699 3170 9733
rect 3204 9699 3238 9733
rect 3272 9699 3306 9733
rect 3340 9699 3374 9733
rect 3408 9699 3442 9733
rect 3476 9699 3510 9733
rect 3544 9699 3578 9733
rect 3612 9699 3646 9733
rect 3680 9699 3714 9733
rect 3748 9699 3782 9733
rect 3816 9699 3850 9733
rect 3884 9699 3918 9733
rect 3952 9699 3986 9733
rect 4020 9699 4054 9733
rect 4088 9699 4122 9733
rect 4156 9699 4190 9733
rect 4224 9699 4258 9733
rect 4292 9699 4326 9733
rect 4651 9732 4685 9766
rect 4762 9699 4796 9733
rect 4830 9699 4864 9733
rect 4898 9699 4932 9733
rect 4966 9699 5000 9733
rect 5034 9699 5068 9733
rect 5102 9699 5136 9733
rect 5170 9699 5204 9733
rect 5238 9699 5272 9733
rect 5306 9699 5340 9733
rect 5374 9699 5408 9733
rect 5442 9699 5476 9733
rect 5510 9699 5544 9733
rect 5578 9699 5612 9733
rect 5646 9699 5680 9733
rect 5714 9699 5748 9733
rect 5782 9699 5816 9733
rect 5850 9699 5884 9733
rect 5918 9699 5952 9733
rect 5986 9699 6020 9733
rect 351 9665 385 9699
rect 351 9597 385 9631
rect 351 9529 385 9563
rect 6019 9616 6053 9650
rect 6019 9548 6053 9582
rect 351 9461 385 9495
rect 351 9393 385 9427
rect 351 9325 385 9359
rect 351 9257 385 9291
rect 351 9189 385 9223
rect 351 9121 385 9155
rect 351 9053 385 9087
rect 351 8985 385 9019
rect 351 8917 385 8951
rect 351 8849 385 8883
rect 351 8781 385 8815
rect 351 8713 385 8747
rect 351 8645 385 8679
rect 351 8577 385 8611
rect 351 8509 385 8543
rect 351 8441 385 8475
rect 351 8373 385 8407
rect 351 8305 385 8339
rect 351 8237 385 8271
rect 351 8169 385 8203
rect 351 8101 385 8135
rect 351 8033 385 8067
rect 351 7965 385 7999
rect 351 7897 385 7931
rect 351 7829 385 7863
rect 351 7761 385 7795
rect 351 7693 385 7727
rect 351 7625 385 7659
rect 351 7557 385 7591
rect 351 7489 385 7523
rect 351 7421 385 7455
rect 351 7353 385 7387
rect 351 7285 385 7319
rect 351 7217 385 7251
rect 351 7149 385 7183
rect 351 7081 385 7115
rect 351 7013 385 7047
rect 351 6945 385 6979
rect 351 6877 385 6911
rect 351 6809 385 6843
rect 351 6741 385 6775
rect 351 6673 385 6707
rect 351 6605 385 6639
rect 351 6537 385 6571
rect 351 6469 385 6503
rect 351 6401 385 6435
rect 351 6333 385 6367
rect 351 6265 385 6299
rect 351 6197 385 6231
rect 351 6129 385 6163
rect 351 6061 385 6095
rect 351 5993 385 6027
rect 351 5925 385 5959
rect 351 5857 385 5891
rect 351 5789 385 5823
rect 351 5721 385 5755
rect 351 5653 385 5687
rect 351 5585 385 5619
rect 351 5517 385 5551
rect 351 5449 385 5483
rect 351 5381 385 5415
rect 351 5313 385 5347
rect 351 5245 385 5279
rect 351 5177 385 5211
rect 351 5109 385 5143
rect 351 5041 385 5075
rect 351 4973 385 5007
rect 351 4905 385 4939
rect 351 4837 385 4871
rect 351 4769 385 4803
rect 351 4701 385 4735
rect 351 4633 385 4667
rect 351 4565 385 4599
rect 351 4497 385 4531
rect 351 4429 385 4463
rect 351 4361 385 4395
rect 351 4293 385 4327
rect 351 4225 385 4259
rect 351 4157 385 4191
rect 351 4089 385 4123
rect 351 4021 385 4055
rect 351 3953 385 3987
rect 351 3885 385 3919
rect 351 3817 385 3851
rect 351 3749 385 3783
rect 351 3681 385 3715
rect 351 3613 385 3647
rect 351 3545 385 3579
rect 351 3477 385 3511
rect 351 3409 385 3443
rect 351 3341 385 3375
rect 351 3273 385 3307
rect 351 3205 385 3239
rect 351 3137 385 3171
rect 351 3069 385 3103
rect 351 3001 385 3035
rect 351 2933 385 2967
rect 351 2865 385 2899
rect 351 2797 385 2831
rect 351 2729 385 2763
rect 351 2661 385 2695
rect 351 2593 385 2627
rect 351 2525 385 2559
rect 351 2457 385 2491
rect 351 2389 385 2423
rect 351 2321 385 2355
rect 351 2253 385 2287
rect 351 2185 385 2219
rect 351 2117 385 2151
rect 351 2049 385 2083
rect 351 1981 385 2015
rect 351 1913 385 1947
rect 351 1845 385 1879
rect 351 1777 385 1811
rect 351 1709 385 1743
rect 351 1641 385 1675
rect 351 1573 385 1607
rect 351 1505 385 1539
rect 351 1437 385 1471
rect 351 1369 385 1403
rect 351 1301 385 1335
rect 351 1233 385 1267
rect 351 1165 385 1199
rect 351 1097 385 1131
rect 351 1029 385 1063
rect 351 961 385 995
rect 351 893 385 927
rect 351 825 385 859
rect 351 757 385 791
rect 351 689 385 723
rect 351 621 385 655
rect 351 553 385 587
rect 6019 9480 6053 9514
rect 6019 9412 6053 9446
rect 6019 9344 6053 9378
rect 6019 9276 6053 9310
rect 6019 9208 6053 9242
rect 6019 9140 6053 9174
rect 6019 9072 6053 9106
rect 6019 9004 6053 9038
rect 6019 8936 6053 8970
rect 6019 8868 6053 8902
rect 6019 8800 6053 8834
rect 6019 8732 6053 8766
rect 6019 8664 6053 8698
rect 6019 8596 6053 8630
rect 6019 8528 6053 8562
rect 6019 8460 6053 8494
rect 6019 8392 6053 8426
rect 6019 8324 6053 8358
rect 6019 8256 6053 8290
rect 6019 8188 6053 8222
rect 6019 8120 6053 8154
rect 6019 8052 6053 8086
rect 6019 7984 6053 8018
rect 6019 7916 6053 7950
rect 6019 7848 6053 7882
rect 6019 7780 6053 7814
rect 6019 7712 6053 7746
rect 6019 7644 6053 7678
rect 6019 7576 6053 7610
rect 6019 7508 6053 7542
rect 6019 7440 6053 7474
rect 6019 7372 6053 7406
rect 6019 7304 6053 7338
rect 6019 7236 6053 7270
rect 6019 7168 6053 7202
rect 6019 7100 6053 7134
rect 6019 7032 6053 7066
rect 6019 6964 6053 6998
rect 6019 6896 6053 6930
rect 6019 6828 6053 6862
rect 6019 6760 6053 6794
rect 6019 6692 6053 6726
rect 6019 6624 6053 6658
rect 6019 6556 6053 6590
rect 6019 6488 6053 6522
rect 6019 6420 6053 6454
rect 6019 6352 6053 6386
rect 6019 6284 6053 6318
rect 6019 6216 6053 6250
rect 6019 6148 6053 6182
rect 6019 6080 6053 6114
rect 6019 6012 6053 6046
rect 6019 5944 6053 5978
rect 6019 5876 6053 5910
rect 6019 5808 6053 5842
rect 6019 5740 6053 5774
rect 6019 5672 6053 5706
rect 6019 5604 6053 5638
rect 6019 5536 6053 5570
rect 6019 5468 6053 5502
rect 6019 5400 6053 5434
rect 6019 5332 6053 5366
rect 6019 5264 6053 5298
rect 6019 5196 6053 5230
rect 6019 5128 6053 5162
rect 6019 5060 6053 5094
rect 6019 4992 6053 5026
rect 6019 4924 6053 4958
rect 6019 4856 6053 4890
rect 6019 4788 6053 4822
rect 6019 4720 6053 4754
rect 6019 4652 6053 4686
rect 6019 4584 6053 4618
rect 6019 4516 6053 4550
rect 6019 4448 6053 4482
rect 6019 4380 6053 4414
rect 6019 4312 6053 4346
rect 6019 4244 6053 4278
rect 6019 4176 6053 4210
rect 6019 4108 6053 4142
rect 6019 4040 6053 4074
rect 6019 3972 6053 4006
rect 6019 3904 6053 3938
rect 6019 3836 6053 3870
rect 6019 3768 6053 3802
rect 6019 3700 6053 3734
rect 6019 3632 6053 3666
rect 6019 3564 6053 3598
rect 6019 3496 6053 3530
rect 6019 3428 6053 3462
rect 6019 3360 6053 3394
rect 6019 3292 6053 3326
rect 6019 3224 6053 3258
rect 6019 3156 6053 3190
rect 6019 3088 6053 3122
rect 6019 3020 6053 3054
rect 6019 2952 6053 2986
rect 6019 2884 6053 2918
rect 6019 2816 6053 2850
rect 6019 2748 6053 2782
rect 6019 2680 6053 2714
rect 6019 2612 6053 2646
rect 6019 2544 6053 2578
rect 6019 2476 6053 2510
rect 6019 2408 6053 2442
rect 6019 2340 6053 2374
rect 6019 2272 6053 2306
rect 6019 2204 6053 2238
rect 6019 2136 6053 2170
rect 6019 2068 6053 2102
rect 6019 2000 6053 2034
rect 6019 1932 6053 1966
rect 6019 1864 6053 1898
rect 6019 1796 6053 1830
rect 6019 1728 6053 1762
rect 6019 1660 6053 1694
rect 6019 1592 6053 1626
rect 6019 1524 6053 1558
rect 6019 1456 6053 1490
rect 6019 1388 6053 1422
rect 6019 1320 6053 1354
rect 6019 1252 6053 1286
rect 6019 1184 6053 1218
rect 6019 1116 6053 1150
rect 6019 1048 6053 1082
rect 6019 980 6053 1014
rect 6019 912 6053 946
rect 6019 844 6053 878
rect 6019 776 6053 810
rect 6019 708 6053 742
rect 6019 640 6053 674
rect 6019 572 6053 606
rect 6019 504 6053 538
rect 384 368 418 402
rect 452 368 486 402
rect 520 368 554 402
rect 588 368 622 402
rect 656 368 690 402
rect 724 368 758 402
rect 792 368 826 402
rect 860 368 894 402
rect 928 368 962 402
rect 996 368 1030 402
rect 1064 368 1098 402
rect 1132 368 1166 402
rect 1200 368 1234 402
rect 1268 368 1302 402
rect 1336 368 1370 402
rect 1404 368 1438 402
rect 1472 368 1506 402
rect 1540 368 1574 402
rect 1608 368 1642 402
rect 1676 368 1710 402
rect 1744 368 1778 402
rect 1812 368 1846 402
rect 1880 368 1914 402
rect 1948 368 1982 402
rect 2016 368 2050 402
rect 2084 368 2118 402
rect 2152 368 2186 402
rect 2220 368 2254 402
rect 2288 368 2322 402
rect 2356 368 2390 402
rect 2424 368 2458 402
rect 2492 368 2526 402
rect 2560 368 2594 402
rect 2628 368 2662 402
rect 2696 368 2730 402
rect 2764 368 2798 402
rect 2832 368 2866 402
rect 2900 368 2934 402
rect 2968 368 3002 402
rect 3036 368 3070 402
rect 3104 368 3138 402
rect 3172 368 3206 402
rect 3240 368 3274 402
rect 3308 368 3342 402
rect 3376 368 3410 402
rect 3444 368 3478 402
rect 3512 368 3546 402
rect 3580 368 3614 402
rect 3648 368 3682 402
rect 3716 368 3750 402
rect 3784 368 3818 402
rect 3852 368 3886 402
rect 3920 368 3954 402
rect 3988 368 4022 402
rect 4056 368 4090 402
rect 4124 368 4158 402
rect 4192 368 4226 402
rect 4260 368 4294 402
rect 4328 368 4362 402
rect 4396 368 4430 402
rect 4464 368 4498 402
rect 4532 368 4566 402
rect 4600 368 4634 402
rect 4668 368 4702 402
rect 4736 368 4770 402
rect 4804 368 4838 402
rect 4872 368 4906 402
rect 4940 368 4974 402
rect 5008 368 5042 402
rect 5076 368 5110 402
rect 5144 368 5178 402
rect 5212 368 5246 402
rect 5280 368 5314 402
rect 5348 368 5382 402
rect 5416 368 5450 402
rect 5484 368 5518 402
rect 5552 368 5586 402
rect 5620 368 5654 402
rect 5688 368 5722 402
rect 5756 368 5790 402
rect 5824 368 5858 402
rect 5892 368 5926 402
rect 6019 401 6053 435
<< poly >>
rect 10207 34454 11007 34470
rect 10207 34420 10223 34454
rect 10257 34420 10297 34454
rect 10331 34420 10371 34454
rect 10405 34420 10445 34454
rect 10479 34420 10519 34454
rect 10553 34420 10592 34454
rect 10626 34420 10665 34454
rect 10699 34420 10738 34454
rect 10772 34420 10811 34454
rect 10845 34420 10884 34454
rect 10918 34420 10957 34454
rect 10991 34420 11007 34454
rect 10207 34404 11007 34420
rect 11063 34454 14031 34470
rect 11063 34420 11079 34454
rect 11113 34420 11148 34454
rect 11182 34420 11217 34454
rect 11251 34420 11286 34454
rect 11320 34420 11355 34454
rect 11389 34420 11424 34454
rect 11458 34420 11493 34454
rect 11527 34420 11562 34454
rect 11596 34420 11631 34454
rect 11665 34420 11700 34454
rect 11734 34420 11769 34454
rect 11803 34420 11838 34454
rect 11872 34420 11907 34454
rect 11941 34420 11976 34454
rect 12010 34420 12045 34454
rect 12079 34420 12114 34454
rect 12148 34420 12183 34454
rect 12217 34420 12252 34454
rect 12286 34420 12321 34454
rect 12355 34420 12390 34454
rect 12424 34420 12459 34454
rect 12493 34420 12528 34454
rect 12562 34420 12597 34454
rect 12631 34420 12666 34454
rect 12700 34420 12735 34454
rect 12769 34420 12804 34454
rect 12838 34420 12873 34454
rect 12907 34420 12942 34454
rect 12976 34420 13011 34454
rect 13045 34420 13080 34454
rect 13114 34420 13149 34454
rect 13183 34420 13218 34454
rect 13252 34420 13287 34454
rect 13321 34420 13356 34454
rect 13390 34420 13425 34454
rect 13459 34420 13494 34454
rect 13528 34420 13563 34454
rect 13597 34420 13632 34454
rect 13666 34420 13701 34454
rect 13735 34420 13771 34454
rect 13805 34420 13841 34454
rect 13875 34420 13911 34454
rect 13945 34420 13981 34454
rect 14015 34420 14031 34454
rect 11063 34404 14031 34420
rect 10207 32202 11007 32218
rect 10207 32168 10223 32202
rect 10257 32168 10297 32202
rect 10331 32168 10371 32202
rect 10405 32168 10445 32202
rect 10479 32168 10519 32202
rect 10553 32168 10592 32202
rect 10626 32168 10665 32202
rect 10699 32168 10738 32202
rect 10772 32168 10811 32202
rect 10845 32168 10884 32202
rect 10918 32168 10957 32202
rect 10991 32168 11007 32202
rect 10207 32152 11007 32168
rect 11063 32202 14031 32218
rect 11063 32168 11079 32202
rect 11113 32168 11148 32202
rect 11182 32168 11217 32202
rect 11251 32168 11286 32202
rect 11320 32168 11355 32202
rect 11389 32168 11424 32202
rect 11458 32168 11493 32202
rect 11527 32168 11562 32202
rect 11596 32168 11631 32202
rect 11665 32168 11700 32202
rect 11734 32168 11769 32202
rect 11803 32168 11838 32202
rect 11872 32168 11907 32202
rect 11941 32168 11976 32202
rect 12010 32168 12045 32202
rect 12079 32168 12114 32202
rect 12148 32168 12183 32202
rect 12217 32168 12252 32202
rect 12286 32168 12321 32202
rect 12355 32168 12390 32202
rect 12424 32168 12459 32202
rect 12493 32168 12528 32202
rect 12562 32168 12597 32202
rect 12631 32168 12666 32202
rect 12700 32168 12735 32202
rect 12769 32168 12804 32202
rect 12838 32168 12873 32202
rect 12907 32168 12942 32202
rect 12976 32168 13011 32202
rect 13045 32168 13080 32202
rect 13114 32168 13149 32202
rect 13183 32168 13218 32202
rect 13252 32168 13287 32202
rect 13321 32168 13356 32202
rect 13390 32168 13425 32202
rect 13459 32168 13494 32202
rect 13528 32168 13563 32202
rect 13597 32168 13632 32202
rect 13666 32168 13701 32202
rect 13735 32168 13771 32202
rect 13805 32168 13841 32202
rect 13875 32168 13911 32202
rect 13945 32168 13981 32202
rect 14015 32168 14031 32202
rect 11063 32152 14031 32168
rect 9431 31435 9831 31451
rect 9431 31401 9447 31435
rect 9481 31401 9531 31435
rect 9565 31401 9615 31435
rect 9649 31401 9698 31435
rect 9732 31401 9781 31435
rect 9815 31401 9831 31435
rect 9431 31385 9831 31401
rect 10207 29953 11007 29969
rect 10207 29919 10223 29953
rect 10257 29919 10297 29953
rect 10331 29919 10371 29953
rect 10405 29919 10445 29953
rect 10479 29919 10519 29953
rect 10553 29919 10592 29953
rect 10626 29919 10665 29953
rect 10699 29919 10738 29953
rect 10772 29919 10811 29953
rect 10845 29919 10884 29953
rect 10918 29919 10957 29953
rect 10991 29919 11007 29953
rect 10207 29903 11007 29919
rect 11063 29953 14031 29969
rect 11063 29919 11079 29953
rect 11113 29919 11148 29953
rect 11182 29919 11217 29953
rect 11251 29919 11286 29953
rect 11320 29919 11355 29953
rect 11389 29919 11424 29953
rect 11458 29919 11493 29953
rect 11527 29919 11562 29953
rect 11596 29919 11631 29953
rect 11665 29919 11700 29953
rect 11734 29919 11769 29953
rect 11803 29919 11838 29953
rect 11872 29919 11907 29953
rect 11941 29919 11976 29953
rect 12010 29919 12045 29953
rect 12079 29919 12114 29953
rect 12148 29919 12183 29953
rect 12217 29919 12252 29953
rect 12286 29919 12321 29953
rect 12355 29919 12390 29953
rect 12424 29919 12459 29953
rect 12493 29919 12528 29953
rect 12562 29919 12597 29953
rect 12631 29919 12666 29953
rect 12700 29919 12735 29953
rect 12769 29919 12804 29953
rect 12838 29919 12873 29953
rect 12907 29919 12942 29953
rect 12976 29919 13011 29953
rect 13045 29919 13080 29953
rect 13114 29919 13149 29953
rect 13183 29919 13218 29953
rect 13252 29919 13287 29953
rect 13321 29919 13356 29953
rect 13390 29919 13425 29953
rect 13459 29919 13494 29953
rect 13528 29919 13563 29953
rect 13597 29919 13632 29953
rect 13666 29919 13701 29953
rect 13735 29919 13771 29953
rect 13805 29919 13841 29953
rect 13875 29919 13911 29953
rect 13945 29919 13981 29953
rect 14015 29919 14031 29953
rect 11063 29903 14031 29919
rect 10089 27455 10155 27471
rect 10089 27421 10105 27455
rect 10139 27421 10155 27455
rect 10089 27382 10155 27421
rect 10089 27348 10105 27382
rect 10139 27348 10155 27382
rect 10089 27309 10155 27348
rect 10089 27275 10105 27309
rect 10139 27275 10155 27309
rect 10089 27236 10155 27275
rect 10089 27202 10105 27236
rect 10139 27202 10155 27236
rect 10089 27163 10155 27202
rect 10089 27129 10105 27163
rect 10139 27129 10155 27163
rect 10089 27090 10155 27129
rect 10089 27056 10105 27090
rect 10139 27056 10155 27090
rect 10089 27017 10155 27056
rect 10089 26983 10105 27017
rect 10139 26983 10155 27017
rect 10089 26943 10155 26983
rect 10089 26909 10105 26943
rect 10139 26909 10155 26943
rect 10089 26869 10155 26909
rect 10089 26835 10105 26869
rect 10139 26835 10155 26869
rect 10089 26795 10155 26835
rect 10089 26761 10105 26795
rect 10139 26761 10155 26795
rect 10089 26721 10155 26761
rect 10089 26687 10105 26721
rect 10139 26687 10155 26721
rect 10089 26671 10155 26687
rect 293 17219 306 17285
rect 848 17219 861 17285
rect 293 17213 393 17219
rect 449 17213 549 17219
rect 605 17213 705 17219
rect 761 17213 861 17219
rect 236 16823 393 16839
rect 236 16789 252 16823
rect 286 16789 320 16823
rect 354 16789 393 16823
rect 236 16773 393 16789
rect 293 16767 393 16773
rect 449 16823 849 16839
rect 449 16789 496 16823
rect 530 16789 564 16823
rect 598 16789 632 16823
rect 666 16789 700 16823
rect 734 16789 768 16823
rect 802 16789 849 16823
rect 449 16767 849 16789
rect 905 16823 1305 16839
rect 905 16789 952 16823
rect 986 16789 1020 16823
rect 1054 16789 1088 16823
rect 1122 16789 1156 16823
rect 1190 16789 1224 16823
rect 1258 16789 1305 16823
rect 905 16767 1305 16789
rect 1361 16823 1761 16839
rect 1361 16789 1408 16823
rect 1442 16789 1476 16823
rect 1510 16789 1544 16823
rect 1578 16789 1612 16823
rect 1646 16789 1680 16823
rect 1714 16789 1761 16823
rect 1361 16767 1761 16789
rect 1817 16823 2217 16839
rect 1817 16789 1864 16823
rect 1898 16789 1932 16823
rect 1966 16789 2000 16823
rect 2034 16789 2068 16823
rect 2102 16789 2136 16823
rect 2170 16789 2217 16823
rect 1817 16767 2217 16789
rect 2273 16823 2407 16839
rect 2273 16789 2289 16823
rect 2323 16789 2357 16823
rect 2391 16789 2407 16823
rect 2273 16773 2407 16789
rect 2273 16767 2373 16773
rect 2629 16823 2763 16839
rect 2629 16789 2645 16823
rect 2679 16789 2713 16823
rect 2747 16789 2763 16823
rect 2629 16773 2763 16789
rect 2663 16767 2763 16773
rect 2819 16823 3219 16839
rect 2819 16789 2866 16823
rect 2900 16789 2934 16823
rect 2968 16789 3002 16823
rect 3036 16789 3070 16823
rect 3104 16789 3138 16823
rect 3172 16789 3219 16823
rect 2819 16767 3219 16789
rect 3275 16823 3675 16839
rect 3275 16789 3322 16823
rect 3356 16789 3390 16823
rect 3424 16789 3458 16823
rect 3492 16789 3526 16823
rect 3560 16789 3594 16823
rect 3628 16789 3675 16823
rect 3275 16767 3675 16789
rect 3731 16823 4131 16839
rect 3731 16789 3778 16823
rect 3812 16789 3846 16823
rect 3880 16789 3914 16823
rect 3948 16789 3982 16823
rect 4016 16789 4050 16823
rect 4084 16789 4131 16823
rect 3731 16767 4131 16789
rect 4187 16823 4587 16839
rect 4187 16789 4234 16823
rect 4268 16789 4302 16823
rect 4336 16789 4370 16823
rect 4404 16789 4438 16823
rect 4472 16789 4506 16823
rect 4540 16789 4587 16823
rect 4187 16767 4587 16789
rect 4643 16823 4777 16839
rect 4643 16789 4659 16823
rect 4693 16789 4727 16823
rect 4761 16789 4777 16823
rect 4643 16773 4777 16789
rect 4643 16767 4743 16773
rect 293 15309 393 15315
rect 259 15293 393 15309
rect 259 15259 275 15293
rect 309 15259 343 15293
rect 377 15259 393 15293
rect 259 15243 393 15259
rect 293 15237 393 15243
rect 2273 15309 2373 15315
rect 2663 15309 2763 15315
rect 2273 15293 2407 15309
rect 2273 15259 2289 15293
rect 2323 15259 2357 15293
rect 2391 15259 2407 15293
rect 2273 15243 2407 15259
rect 2273 15237 2373 15243
rect 2629 15293 2763 15309
rect 2629 15259 2645 15293
rect 2679 15259 2713 15293
rect 2747 15259 2763 15293
rect 2629 15243 2763 15259
rect 2663 15237 2763 15243
rect 4643 15309 4743 15315
rect 4643 15293 4777 15309
rect 4643 15259 4659 15293
rect 4693 15259 4727 15293
rect 4761 15259 4777 15293
rect 4643 15243 4777 15259
rect 4643 15237 4743 15243
rect 293 13779 393 13785
rect 259 13763 393 13779
rect 259 13729 275 13763
rect 309 13729 343 13763
rect 377 13729 393 13763
rect 259 13713 393 13729
rect 293 13707 393 13713
rect 449 13763 849 13785
rect 449 13729 496 13763
rect 530 13729 564 13763
rect 598 13729 632 13763
rect 666 13729 700 13763
rect 734 13729 768 13763
rect 802 13729 849 13763
rect 449 13707 849 13729
rect 905 13763 1305 13785
rect 905 13729 952 13763
rect 986 13729 1020 13763
rect 1054 13729 1088 13763
rect 1122 13729 1156 13763
rect 1190 13729 1224 13763
rect 1258 13729 1305 13763
rect 905 13707 1305 13729
rect 1361 13763 1761 13785
rect 1361 13729 1408 13763
rect 1442 13729 1476 13763
rect 1510 13729 1544 13763
rect 1578 13729 1612 13763
rect 1646 13729 1680 13763
rect 1714 13729 1761 13763
rect 1361 13707 1761 13729
rect 1817 13763 2217 13785
rect 1817 13729 1864 13763
rect 1898 13729 1932 13763
rect 1966 13729 2000 13763
rect 2034 13729 2068 13763
rect 2102 13729 2136 13763
rect 2170 13729 2217 13763
rect 1817 13707 2217 13729
rect 2273 13779 2373 13785
rect 5225 15730 5521 15746
rect 5225 15696 5254 15730
rect 5288 15696 5322 15730
rect 5356 15696 5390 15730
rect 5424 15696 5458 15730
rect 5492 15696 5521 15730
rect 5225 15680 5521 15696
rect 5225 15674 5345 15680
rect 5401 15674 5521 15680
rect 2663 13779 2763 13785
rect 2273 13763 2407 13779
rect 2273 13729 2289 13763
rect 2323 13729 2357 13763
rect 2391 13729 2407 13763
rect 2273 13713 2407 13729
rect 2273 13707 2373 13713
rect 2629 13763 2763 13779
rect 2629 13729 2645 13763
rect 2679 13729 2713 13763
rect 2747 13729 2763 13763
rect 2629 13713 2763 13729
rect 2663 13707 2763 13713
rect 2819 13763 3219 13785
rect 2819 13729 2866 13763
rect 2900 13729 2934 13763
rect 2968 13729 3002 13763
rect 3036 13729 3070 13763
rect 3104 13729 3138 13763
rect 3172 13729 3219 13763
rect 2819 13707 3219 13729
rect 3275 13763 3675 13785
rect 3275 13729 3322 13763
rect 3356 13729 3390 13763
rect 3424 13729 3458 13763
rect 3492 13729 3526 13763
rect 3560 13729 3594 13763
rect 3628 13729 3675 13763
rect 3275 13707 3675 13729
rect 3731 13763 4131 13785
rect 3731 13729 3778 13763
rect 3812 13729 3846 13763
rect 3880 13729 3914 13763
rect 3948 13729 3982 13763
rect 4016 13729 4050 13763
rect 4084 13729 4131 13763
rect 3731 13707 4131 13729
rect 4187 13763 4587 13785
rect 4187 13729 4234 13763
rect 4268 13729 4302 13763
rect 4336 13729 4370 13763
rect 4404 13729 4438 13763
rect 4472 13729 4506 13763
rect 4540 13729 4587 13763
rect 4187 13707 4587 13729
rect 4643 13779 4743 13785
rect 4643 13763 4777 13779
rect 4643 13729 4659 13763
rect 4693 13729 4727 13763
rect 4761 13729 4777 13763
rect 4643 13713 4777 13729
rect 4643 13707 4743 13713
rect 293 12249 393 12255
rect 259 12233 393 12249
rect 259 12199 275 12233
rect 309 12199 343 12233
rect 377 12199 393 12233
rect 259 12183 393 12199
rect 449 12233 849 12255
rect 449 12199 496 12233
rect 530 12199 564 12233
rect 598 12199 632 12233
rect 666 12199 700 12233
rect 734 12199 768 12233
rect 802 12199 849 12233
rect 449 12183 849 12199
rect 905 12233 1305 12255
rect 905 12199 952 12233
rect 986 12199 1020 12233
rect 1054 12199 1088 12233
rect 1122 12199 1156 12233
rect 1190 12199 1224 12233
rect 1258 12199 1305 12233
rect 905 12183 1305 12199
rect 1361 12233 1761 12255
rect 1361 12199 1408 12233
rect 1442 12199 1476 12233
rect 1510 12199 1544 12233
rect 1578 12199 1612 12233
rect 1646 12199 1680 12233
rect 1714 12199 1761 12233
rect 1361 12183 1761 12199
rect 1817 12233 2217 12255
rect 1817 12199 1864 12233
rect 1898 12199 1932 12233
rect 1966 12199 2000 12233
rect 2034 12199 2068 12233
rect 2102 12199 2136 12233
rect 2170 12199 2217 12233
rect 1817 12183 2217 12199
rect 2273 12249 2373 12255
rect 2663 12249 2763 12255
rect 2273 12233 2407 12249
rect 2273 12199 2289 12233
rect 2323 12199 2357 12233
rect 2391 12199 2407 12233
rect 2273 12183 2407 12199
rect 2629 12233 2763 12249
rect 2629 12199 2645 12233
rect 2679 12199 2713 12233
rect 2747 12199 2763 12233
rect 2629 12183 2763 12199
rect 2819 12233 3219 12255
rect 2819 12199 2866 12233
rect 2900 12199 2934 12233
rect 2968 12199 3002 12233
rect 3036 12199 3070 12233
rect 3104 12199 3138 12233
rect 3172 12199 3219 12233
rect 2819 12183 3219 12199
rect 3275 12233 3675 12255
rect 3275 12199 3322 12233
rect 3356 12199 3390 12233
rect 3424 12199 3458 12233
rect 3492 12199 3526 12233
rect 3560 12199 3594 12233
rect 3628 12199 3675 12233
rect 3275 12183 3675 12199
rect 3731 12233 4131 12255
rect 3731 12199 3778 12233
rect 3812 12199 3846 12233
rect 3880 12199 3914 12233
rect 3948 12199 3982 12233
rect 4016 12199 4050 12233
rect 4084 12199 4131 12233
rect 3731 12183 4131 12199
rect 4187 12233 4587 12255
rect 4187 12199 4234 12233
rect 4268 12199 4302 12233
rect 4336 12199 4370 12233
rect 4404 12199 4438 12233
rect 4472 12199 4506 12233
rect 4540 12199 4587 12233
rect 4187 12183 4587 12199
rect 4643 12249 4743 12255
rect 4643 12233 4777 12249
rect 4643 12199 4659 12233
rect 4693 12199 4727 12233
rect 4761 12199 4777 12233
rect 4643 12183 4777 12199
rect 824 12005 1004 12021
rect 824 11971 863 12005
rect 897 11971 931 12005
rect 965 11971 1004 12005
rect 824 11949 1004 11971
rect 1060 12005 1240 12021
rect 1060 11971 1099 12005
rect 1133 11971 1167 12005
rect 1201 11971 1240 12005
rect 1060 11949 1240 11971
rect 1296 12005 1476 12021
rect 1296 11971 1335 12005
rect 1369 11971 1403 12005
rect 1437 11971 1476 12005
rect 1296 11949 1476 11971
rect 1532 12005 1712 12021
rect 1532 11971 1571 12005
rect 1605 11971 1639 12005
rect 1673 11971 1712 12005
rect 1532 11949 1712 11971
rect 1768 12005 1948 12021
rect 1768 11971 1807 12005
rect 1841 11971 1875 12005
rect 1909 11971 1948 12005
rect 1768 11949 1948 11971
rect 2004 12005 2184 12021
rect 2004 11971 2043 12005
rect 2077 11971 2111 12005
rect 2145 11971 2184 12005
rect 2004 11949 2184 11971
rect 824 9875 1004 9897
rect 824 9841 863 9875
rect 897 9841 931 9875
rect 965 9841 1004 9875
rect 824 9825 1004 9841
rect 1060 9875 1240 9897
rect 1060 9841 1099 9875
rect 1133 9841 1167 9875
rect 1201 9841 1240 9875
rect 1060 9825 1240 9841
rect 1296 9875 1476 9897
rect 1296 9841 1335 9875
rect 1369 9841 1403 9875
rect 1437 9841 1476 9875
rect 1296 9825 1476 9841
rect 1532 9875 1712 9897
rect 1532 9841 1571 9875
rect 1605 9841 1639 9875
rect 1673 9841 1712 9875
rect 1532 9825 1712 9841
rect 1768 9875 1948 9897
rect 1768 9841 1807 9875
rect 1841 9841 1875 9875
rect 1909 9841 1948 9875
rect 1768 9825 1948 9841
rect 2004 9875 2184 9897
rect 2852 12005 3032 12021
rect 2852 11971 2891 12005
rect 2925 11971 2959 12005
rect 2993 11971 3032 12005
rect 2004 9841 2043 9875
rect 2077 9841 2111 9875
rect 2145 9841 2184 9875
rect 2004 9825 2184 9841
rect 2852 11949 3032 11971
rect 3088 12005 3268 12021
rect 3088 11971 3127 12005
rect 3161 11971 3195 12005
rect 3229 11971 3268 12005
rect 3088 11949 3268 11971
rect 3324 12005 3504 12021
rect 3324 11971 3363 12005
rect 3397 11971 3431 12005
rect 3465 11971 3504 12005
rect 3324 11949 3504 11971
rect 3560 12005 3740 12021
rect 3560 11971 3599 12005
rect 3633 11971 3667 12005
rect 3701 11971 3740 12005
rect 3560 11949 3740 11971
rect 3796 12005 3976 12021
rect 3796 11971 3835 12005
rect 3869 11971 3903 12005
rect 3937 11971 3976 12005
rect 3796 11949 3976 11971
rect 4032 12005 4212 12021
rect 4032 11971 4071 12005
rect 4105 11971 4139 12005
rect 4173 11971 4212 12005
rect 4032 11949 4212 11971
rect 2852 9875 3032 9897
rect 2852 9841 2891 9875
rect 2925 9841 2959 9875
rect 2993 9841 3032 9875
rect 2852 9825 3032 9841
rect 3088 9875 3268 9897
rect 3088 9841 3127 9875
rect 3161 9841 3195 9875
rect 3229 9841 3268 9875
rect 3088 9825 3268 9841
rect 3324 9875 3504 9897
rect 3324 9841 3363 9875
rect 3397 9841 3431 9875
rect 3465 9841 3504 9875
rect 3324 9825 3504 9841
rect 3560 9875 3740 9897
rect 3560 9841 3599 9875
rect 3633 9841 3667 9875
rect 3701 9841 3740 9875
rect 3560 9825 3740 9841
rect 3796 9875 3976 9897
rect 3796 9841 3835 9875
rect 3869 9841 3903 9875
rect 3937 9841 3976 9875
rect 3796 9825 3976 9841
rect 4032 9875 4212 9897
rect 4032 9841 4071 9875
rect 4105 9841 4139 9875
rect 4173 9841 4212 9875
rect 4032 9825 4212 9841
rect 702 9403 1502 9475
rect 1558 9403 2358 9475
rect 2414 9403 3214 9475
rect 3534 9403 4334 9475
rect 4390 9459 4790 9475
rect 4390 9425 4437 9459
rect 4471 9425 4505 9459
rect 4539 9425 4573 9459
rect 4607 9425 4641 9459
rect 4675 9425 4709 9459
rect 4743 9425 4790 9459
rect 4390 9403 4790 9425
rect 4846 9459 5246 9475
rect 4846 9425 4893 9459
rect 4927 9425 4961 9459
rect 4995 9425 5029 9459
rect 5063 9425 5097 9459
rect 5131 9425 5165 9459
rect 5199 9425 5246 9459
rect 4846 9403 5246 9425
rect 5302 9459 5702 9475
rect 5302 9425 5349 9459
rect 5383 9425 5417 9459
rect 5451 9425 5485 9459
rect 5519 9425 5553 9459
rect 5587 9425 5621 9459
rect 5655 9425 5702 9459
rect 5302 9403 5702 9425
rect 702 7308 1502 7351
rect 1558 7308 2358 7351
rect 2414 7308 3214 7351
rect 1001 7286 1203 7308
rect 1001 7252 1017 7286
rect 1051 7252 1085 7286
rect 1119 7252 1153 7286
rect 1187 7252 1203 7286
rect 1857 7286 2059 7308
rect 1857 7252 1873 7286
rect 1907 7252 1941 7286
rect 1975 7252 2009 7286
rect 2043 7252 2059 7286
rect 2713 7286 2915 7308
rect 3534 7308 4334 7351
rect 4390 7308 4790 7351
rect 4846 7308 5246 7351
rect 5302 7308 5702 7351
rect 2713 7252 2729 7286
rect 2763 7252 2797 7286
rect 2831 7252 2865 7286
rect 2899 7252 2915 7286
rect 3833 7286 4035 7308
rect 3833 7252 3849 7286
rect 3883 7252 3917 7286
rect 3951 7252 3985 7286
rect 4019 7252 4035 7286
rect 4489 7286 4691 7308
rect 4489 7252 4505 7286
rect 4539 7252 4573 7286
rect 4607 7252 4641 7286
rect 4675 7252 4691 7286
rect 4945 7286 5147 7308
rect 4945 7252 4961 7286
rect 4995 7252 5029 7286
rect 5063 7252 5097 7286
rect 5131 7252 5147 7286
rect 5401 7286 5603 7308
rect 5401 7252 5417 7286
rect 5451 7252 5485 7286
rect 5519 7252 5553 7286
rect 5587 7252 5603 7286
rect 1001 7232 1203 7252
rect 1857 7232 2059 7252
rect 2713 7232 2915 7252
rect 702 7189 1502 7232
rect 1558 7189 2358 7232
rect 2414 7189 3214 7232
rect 3833 7232 4035 7252
rect 4489 7232 4691 7252
rect 4945 7232 5147 7252
rect 5401 7232 5603 7252
rect 3534 7189 4334 7232
rect 4390 7189 4790 7232
rect 4846 7189 5246 7232
rect 5302 7189 5702 7232
rect 702 5088 1502 5137
rect 1558 5088 2358 5137
rect 2414 5088 3214 5137
rect 1001 5066 1203 5088
rect 1001 5032 1017 5066
rect 1051 5032 1085 5066
rect 1119 5032 1153 5066
rect 1187 5032 1203 5066
rect 1857 5066 2059 5088
rect 1857 5032 1873 5066
rect 1907 5032 1941 5066
rect 1975 5032 2009 5066
rect 2043 5032 2059 5066
rect 2713 5066 2915 5088
rect 3534 5088 4334 5137
rect 4390 5088 4790 5137
rect 4846 5088 5246 5137
rect 5302 5088 5702 5137
rect 2713 5032 2729 5066
rect 2763 5032 2797 5066
rect 2831 5032 2865 5066
rect 2899 5032 2915 5066
rect 1001 5012 1203 5032
rect 1857 5012 2059 5032
rect 2713 5012 2915 5032
rect 702 4964 1502 5012
rect 1558 4964 2358 5012
rect 2414 4964 3214 5012
rect 3833 5066 4035 5088
rect 3833 5032 3849 5066
rect 3883 5032 3917 5066
rect 3951 5032 3985 5066
rect 4019 5032 4035 5066
rect 4489 5066 4691 5088
rect 4489 5032 4505 5066
rect 4539 5032 4573 5066
rect 4607 5032 4641 5066
rect 4675 5032 4691 5066
rect 4945 5066 5147 5088
rect 4945 5032 4961 5066
rect 4995 5032 5029 5066
rect 5063 5032 5097 5066
rect 5131 5032 5147 5066
rect 5401 5066 5603 5088
rect 5401 5032 5417 5066
rect 5451 5032 5485 5066
rect 5519 5032 5553 5066
rect 5587 5032 5603 5066
rect 3833 5012 4035 5032
rect 4489 5012 4691 5032
rect 4945 5012 5147 5032
rect 5401 5012 5603 5032
rect 3534 4964 4334 5012
rect 4390 4964 4790 5012
rect 4846 4964 5246 5012
rect 5302 4964 5702 5012
rect 702 2869 1502 2912
rect 1558 2869 2358 2912
rect 2414 2869 3214 2912
rect 1001 2847 1203 2869
rect 1001 2813 1017 2847
rect 1051 2813 1085 2847
rect 1119 2813 1153 2847
rect 1187 2813 1203 2847
rect 1857 2847 2059 2869
rect 1857 2813 1873 2847
rect 1907 2813 1941 2847
rect 1975 2813 2009 2847
rect 2043 2813 2059 2847
rect 2713 2847 2915 2869
rect 3534 2869 4334 2912
rect 4390 2869 4790 2912
rect 4846 2869 5246 2912
rect 5302 2869 5702 2912
rect 2713 2813 2729 2847
rect 2763 2813 2797 2847
rect 2831 2813 2865 2847
rect 2899 2813 2915 2847
rect 3833 2847 4035 2869
rect 3833 2813 3849 2847
rect 3883 2813 3917 2847
rect 3951 2813 3985 2847
rect 4019 2813 4035 2847
rect 4489 2847 4691 2869
rect 4489 2813 4505 2847
rect 4539 2813 4573 2847
rect 4607 2813 4641 2847
rect 4675 2813 4691 2847
rect 4945 2847 5147 2869
rect 4945 2813 4961 2847
rect 4995 2813 5029 2847
rect 5063 2813 5097 2847
rect 5131 2813 5147 2847
rect 5401 2847 5603 2869
rect 5401 2813 5417 2847
rect 5451 2813 5485 2847
rect 5519 2813 5553 2847
rect 5587 2813 5603 2847
rect 1001 2793 1203 2813
rect 1857 2793 2059 2813
rect 2713 2793 2915 2813
rect 702 2750 1502 2793
rect 1558 2750 2358 2793
rect 2414 2750 3214 2793
rect 3833 2793 4035 2813
rect 4489 2793 4691 2813
rect 4945 2793 5147 2813
rect 5401 2793 5603 2813
rect 3534 2750 4334 2793
rect 4390 2750 4790 2793
rect 4846 2750 5246 2793
rect 5302 2750 5702 2793
rect 702 626 1502 698
rect 1558 626 2358 698
rect 2414 626 3214 698
rect 3534 626 4334 698
rect 4390 676 4790 698
rect 4390 642 4437 676
rect 4471 642 4505 676
rect 4539 642 4573 676
rect 4607 642 4641 676
rect 4675 642 4709 676
rect 4743 642 4790 676
rect 4390 626 4790 642
rect 4846 676 5246 698
rect 4846 642 4893 676
rect 4927 642 4961 676
rect 4995 642 5029 676
rect 5063 642 5097 676
rect 5131 642 5165 676
rect 5199 642 5246 676
rect 4846 626 5246 642
rect 5302 676 5702 698
rect 5302 642 5349 676
rect 5383 642 5417 676
rect 5451 642 5485 676
rect 5519 642 5553 676
rect 5587 642 5621 676
rect 5655 642 5702 676
rect 5302 626 5702 642
<< polycont >>
rect 10223 34420 10257 34454
rect 10297 34420 10331 34454
rect 10371 34420 10405 34454
rect 10445 34420 10479 34454
rect 10519 34420 10553 34454
rect 10592 34420 10626 34454
rect 10665 34420 10699 34454
rect 10738 34420 10772 34454
rect 10811 34420 10845 34454
rect 10884 34420 10918 34454
rect 10957 34420 10991 34454
rect 11079 34420 11113 34454
rect 11148 34420 11182 34454
rect 11217 34420 11251 34454
rect 11286 34420 11320 34454
rect 11355 34420 11389 34454
rect 11424 34420 11458 34454
rect 11493 34420 11527 34454
rect 11562 34420 11596 34454
rect 11631 34420 11665 34454
rect 11700 34420 11734 34454
rect 11769 34420 11803 34454
rect 11838 34420 11872 34454
rect 11907 34420 11941 34454
rect 11976 34420 12010 34454
rect 12045 34420 12079 34454
rect 12114 34420 12148 34454
rect 12183 34420 12217 34454
rect 12252 34420 12286 34454
rect 12321 34420 12355 34454
rect 12390 34420 12424 34454
rect 12459 34420 12493 34454
rect 12528 34420 12562 34454
rect 12597 34420 12631 34454
rect 12666 34420 12700 34454
rect 12735 34420 12769 34454
rect 12804 34420 12838 34454
rect 12873 34420 12907 34454
rect 12942 34420 12976 34454
rect 13011 34420 13045 34454
rect 13080 34420 13114 34454
rect 13149 34420 13183 34454
rect 13218 34420 13252 34454
rect 13287 34420 13321 34454
rect 13356 34420 13390 34454
rect 13425 34420 13459 34454
rect 13494 34420 13528 34454
rect 13563 34420 13597 34454
rect 13632 34420 13666 34454
rect 13701 34420 13735 34454
rect 13771 34420 13805 34454
rect 13841 34420 13875 34454
rect 13911 34420 13945 34454
rect 13981 34420 14015 34454
rect 10223 32168 10257 32202
rect 10297 32168 10331 32202
rect 10371 32168 10405 32202
rect 10445 32168 10479 32202
rect 10519 32168 10553 32202
rect 10592 32168 10626 32202
rect 10665 32168 10699 32202
rect 10738 32168 10772 32202
rect 10811 32168 10845 32202
rect 10884 32168 10918 32202
rect 10957 32168 10991 32202
rect 11079 32168 11113 32202
rect 11148 32168 11182 32202
rect 11217 32168 11251 32202
rect 11286 32168 11320 32202
rect 11355 32168 11389 32202
rect 11424 32168 11458 32202
rect 11493 32168 11527 32202
rect 11562 32168 11596 32202
rect 11631 32168 11665 32202
rect 11700 32168 11734 32202
rect 11769 32168 11803 32202
rect 11838 32168 11872 32202
rect 11907 32168 11941 32202
rect 11976 32168 12010 32202
rect 12045 32168 12079 32202
rect 12114 32168 12148 32202
rect 12183 32168 12217 32202
rect 12252 32168 12286 32202
rect 12321 32168 12355 32202
rect 12390 32168 12424 32202
rect 12459 32168 12493 32202
rect 12528 32168 12562 32202
rect 12597 32168 12631 32202
rect 12666 32168 12700 32202
rect 12735 32168 12769 32202
rect 12804 32168 12838 32202
rect 12873 32168 12907 32202
rect 12942 32168 12976 32202
rect 13011 32168 13045 32202
rect 13080 32168 13114 32202
rect 13149 32168 13183 32202
rect 13218 32168 13252 32202
rect 13287 32168 13321 32202
rect 13356 32168 13390 32202
rect 13425 32168 13459 32202
rect 13494 32168 13528 32202
rect 13563 32168 13597 32202
rect 13632 32168 13666 32202
rect 13701 32168 13735 32202
rect 13771 32168 13805 32202
rect 13841 32168 13875 32202
rect 13911 32168 13945 32202
rect 13981 32168 14015 32202
rect 9447 31401 9481 31435
rect 9531 31401 9565 31435
rect 9615 31401 9649 31435
rect 9698 31401 9732 31435
rect 9781 31401 9815 31435
rect 10223 29919 10257 29953
rect 10297 29919 10331 29953
rect 10371 29919 10405 29953
rect 10445 29919 10479 29953
rect 10519 29919 10553 29953
rect 10592 29919 10626 29953
rect 10665 29919 10699 29953
rect 10738 29919 10772 29953
rect 10811 29919 10845 29953
rect 10884 29919 10918 29953
rect 10957 29919 10991 29953
rect 11079 29919 11113 29953
rect 11148 29919 11182 29953
rect 11217 29919 11251 29953
rect 11286 29919 11320 29953
rect 11355 29919 11389 29953
rect 11424 29919 11458 29953
rect 11493 29919 11527 29953
rect 11562 29919 11596 29953
rect 11631 29919 11665 29953
rect 11700 29919 11734 29953
rect 11769 29919 11803 29953
rect 11838 29919 11872 29953
rect 11907 29919 11941 29953
rect 11976 29919 12010 29953
rect 12045 29919 12079 29953
rect 12114 29919 12148 29953
rect 12183 29919 12217 29953
rect 12252 29919 12286 29953
rect 12321 29919 12355 29953
rect 12390 29919 12424 29953
rect 12459 29919 12493 29953
rect 12528 29919 12562 29953
rect 12597 29919 12631 29953
rect 12666 29919 12700 29953
rect 12735 29919 12769 29953
rect 12804 29919 12838 29953
rect 12873 29919 12907 29953
rect 12942 29919 12976 29953
rect 13011 29919 13045 29953
rect 13080 29919 13114 29953
rect 13149 29919 13183 29953
rect 13218 29919 13252 29953
rect 13287 29919 13321 29953
rect 13356 29919 13390 29953
rect 13425 29919 13459 29953
rect 13494 29919 13528 29953
rect 13563 29919 13597 29953
rect 13632 29919 13666 29953
rect 13701 29919 13735 29953
rect 13771 29919 13805 29953
rect 13841 29919 13875 29953
rect 13911 29919 13945 29953
rect 13981 29919 14015 29953
rect 10105 27421 10139 27455
rect 10105 27348 10139 27382
rect 10105 27275 10139 27309
rect 10105 27202 10139 27236
rect 10105 27129 10139 27163
rect 10105 27056 10139 27090
rect 10105 26983 10139 27017
rect 10105 26909 10139 26943
rect 10105 26835 10139 26869
rect 10105 26761 10139 26795
rect 10105 26687 10139 26721
rect 252 16789 286 16823
rect 320 16789 354 16823
rect 496 16789 530 16823
rect 564 16789 598 16823
rect 632 16789 666 16823
rect 700 16789 734 16823
rect 768 16789 802 16823
rect 952 16789 986 16823
rect 1020 16789 1054 16823
rect 1088 16789 1122 16823
rect 1156 16789 1190 16823
rect 1224 16789 1258 16823
rect 1408 16789 1442 16823
rect 1476 16789 1510 16823
rect 1544 16789 1578 16823
rect 1612 16789 1646 16823
rect 1680 16789 1714 16823
rect 1864 16789 1898 16823
rect 1932 16789 1966 16823
rect 2000 16789 2034 16823
rect 2068 16789 2102 16823
rect 2136 16789 2170 16823
rect 2289 16789 2323 16823
rect 2357 16789 2391 16823
rect 2645 16789 2679 16823
rect 2713 16789 2747 16823
rect 2866 16789 2900 16823
rect 2934 16789 2968 16823
rect 3002 16789 3036 16823
rect 3070 16789 3104 16823
rect 3138 16789 3172 16823
rect 3322 16789 3356 16823
rect 3390 16789 3424 16823
rect 3458 16789 3492 16823
rect 3526 16789 3560 16823
rect 3594 16789 3628 16823
rect 3778 16789 3812 16823
rect 3846 16789 3880 16823
rect 3914 16789 3948 16823
rect 3982 16789 4016 16823
rect 4050 16789 4084 16823
rect 4234 16789 4268 16823
rect 4302 16789 4336 16823
rect 4370 16789 4404 16823
rect 4438 16789 4472 16823
rect 4506 16789 4540 16823
rect 4659 16789 4693 16823
rect 4727 16789 4761 16823
rect 275 15259 309 15293
rect 343 15259 377 15293
rect 2289 15259 2323 15293
rect 2357 15259 2391 15293
rect 2645 15259 2679 15293
rect 2713 15259 2747 15293
rect 4659 15259 4693 15293
rect 4727 15259 4761 15293
rect 275 13729 309 13763
rect 343 13729 377 13763
rect 496 13729 530 13763
rect 564 13729 598 13763
rect 632 13729 666 13763
rect 700 13729 734 13763
rect 768 13729 802 13763
rect 952 13729 986 13763
rect 1020 13729 1054 13763
rect 1088 13729 1122 13763
rect 1156 13729 1190 13763
rect 1224 13729 1258 13763
rect 1408 13729 1442 13763
rect 1476 13729 1510 13763
rect 1544 13729 1578 13763
rect 1612 13729 1646 13763
rect 1680 13729 1714 13763
rect 1864 13729 1898 13763
rect 1932 13729 1966 13763
rect 2000 13729 2034 13763
rect 2068 13729 2102 13763
rect 2136 13729 2170 13763
rect 5254 15696 5288 15730
rect 5322 15696 5356 15730
rect 5390 15696 5424 15730
rect 5458 15696 5492 15730
rect 2289 13729 2323 13763
rect 2357 13729 2391 13763
rect 2645 13729 2679 13763
rect 2713 13729 2747 13763
rect 2866 13729 2900 13763
rect 2934 13729 2968 13763
rect 3002 13729 3036 13763
rect 3070 13729 3104 13763
rect 3138 13729 3172 13763
rect 3322 13729 3356 13763
rect 3390 13729 3424 13763
rect 3458 13729 3492 13763
rect 3526 13729 3560 13763
rect 3594 13729 3628 13763
rect 3778 13729 3812 13763
rect 3846 13729 3880 13763
rect 3914 13729 3948 13763
rect 3982 13729 4016 13763
rect 4050 13729 4084 13763
rect 4234 13729 4268 13763
rect 4302 13729 4336 13763
rect 4370 13729 4404 13763
rect 4438 13729 4472 13763
rect 4506 13729 4540 13763
rect 4659 13729 4693 13763
rect 4727 13729 4761 13763
rect 275 12199 309 12233
rect 343 12199 377 12233
rect 496 12199 530 12233
rect 564 12199 598 12233
rect 632 12199 666 12233
rect 700 12199 734 12233
rect 768 12199 802 12233
rect 952 12199 986 12233
rect 1020 12199 1054 12233
rect 1088 12199 1122 12233
rect 1156 12199 1190 12233
rect 1224 12199 1258 12233
rect 1408 12199 1442 12233
rect 1476 12199 1510 12233
rect 1544 12199 1578 12233
rect 1612 12199 1646 12233
rect 1680 12199 1714 12233
rect 1864 12199 1898 12233
rect 1932 12199 1966 12233
rect 2000 12199 2034 12233
rect 2068 12199 2102 12233
rect 2136 12199 2170 12233
rect 2289 12199 2323 12233
rect 2357 12199 2391 12233
rect 2645 12199 2679 12233
rect 2713 12199 2747 12233
rect 2866 12199 2900 12233
rect 2934 12199 2968 12233
rect 3002 12199 3036 12233
rect 3070 12199 3104 12233
rect 3138 12199 3172 12233
rect 3322 12199 3356 12233
rect 3390 12199 3424 12233
rect 3458 12199 3492 12233
rect 3526 12199 3560 12233
rect 3594 12199 3628 12233
rect 3778 12199 3812 12233
rect 3846 12199 3880 12233
rect 3914 12199 3948 12233
rect 3982 12199 4016 12233
rect 4050 12199 4084 12233
rect 4234 12199 4268 12233
rect 4302 12199 4336 12233
rect 4370 12199 4404 12233
rect 4438 12199 4472 12233
rect 4506 12199 4540 12233
rect 4659 12199 4693 12233
rect 4727 12199 4761 12233
rect 863 11971 897 12005
rect 931 11971 965 12005
rect 1099 11971 1133 12005
rect 1167 11971 1201 12005
rect 1335 11971 1369 12005
rect 1403 11971 1437 12005
rect 1571 11971 1605 12005
rect 1639 11971 1673 12005
rect 1807 11971 1841 12005
rect 1875 11971 1909 12005
rect 2043 11971 2077 12005
rect 2111 11971 2145 12005
rect 863 9841 897 9875
rect 931 9841 965 9875
rect 1099 9841 1133 9875
rect 1167 9841 1201 9875
rect 1335 9841 1369 9875
rect 1403 9841 1437 9875
rect 1571 9841 1605 9875
rect 1639 9841 1673 9875
rect 1807 9841 1841 9875
rect 1875 9841 1909 9875
rect 2891 11971 2925 12005
rect 2959 11971 2993 12005
rect 2043 9841 2077 9875
rect 2111 9841 2145 9875
rect 3127 11971 3161 12005
rect 3195 11971 3229 12005
rect 3363 11971 3397 12005
rect 3431 11971 3465 12005
rect 3599 11971 3633 12005
rect 3667 11971 3701 12005
rect 3835 11971 3869 12005
rect 3903 11971 3937 12005
rect 4071 11971 4105 12005
rect 4139 11971 4173 12005
rect 2891 9841 2925 9875
rect 2959 9841 2993 9875
rect 3127 9841 3161 9875
rect 3195 9841 3229 9875
rect 3363 9841 3397 9875
rect 3431 9841 3465 9875
rect 3599 9841 3633 9875
rect 3667 9841 3701 9875
rect 3835 9841 3869 9875
rect 3903 9841 3937 9875
rect 4071 9841 4105 9875
rect 4139 9841 4173 9875
rect 4437 9425 4471 9459
rect 4505 9425 4539 9459
rect 4573 9425 4607 9459
rect 4641 9425 4675 9459
rect 4709 9425 4743 9459
rect 4893 9425 4927 9459
rect 4961 9425 4995 9459
rect 5029 9425 5063 9459
rect 5097 9425 5131 9459
rect 5165 9425 5199 9459
rect 5349 9425 5383 9459
rect 5417 9425 5451 9459
rect 5485 9425 5519 9459
rect 5553 9425 5587 9459
rect 5621 9425 5655 9459
rect 1017 7252 1051 7286
rect 1085 7252 1119 7286
rect 1153 7252 1187 7286
rect 1873 7252 1907 7286
rect 1941 7252 1975 7286
rect 2009 7252 2043 7286
rect 2729 7252 2763 7286
rect 2797 7252 2831 7286
rect 2865 7252 2899 7286
rect 3849 7252 3883 7286
rect 3917 7252 3951 7286
rect 3985 7252 4019 7286
rect 4505 7252 4539 7286
rect 4573 7252 4607 7286
rect 4641 7252 4675 7286
rect 4961 7252 4995 7286
rect 5029 7252 5063 7286
rect 5097 7252 5131 7286
rect 5417 7252 5451 7286
rect 5485 7252 5519 7286
rect 5553 7252 5587 7286
rect 1017 5032 1051 5066
rect 1085 5032 1119 5066
rect 1153 5032 1187 5066
rect 1873 5032 1907 5066
rect 1941 5032 1975 5066
rect 2009 5032 2043 5066
rect 2729 5032 2763 5066
rect 2797 5032 2831 5066
rect 2865 5032 2899 5066
rect 3849 5032 3883 5066
rect 3917 5032 3951 5066
rect 3985 5032 4019 5066
rect 4505 5032 4539 5066
rect 4573 5032 4607 5066
rect 4641 5032 4675 5066
rect 4961 5032 4995 5066
rect 5029 5032 5063 5066
rect 5097 5032 5131 5066
rect 5417 5032 5451 5066
rect 5485 5032 5519 5066
rect 5553 5032 5587 5066
rect 1017 2813 1051 2847
rect 1085 2813 1119 2847
rect 1153 2813 1187 2847
rect 1873 2813 1907 2847
rect 1941 2813 1975 2847
rect 2009 2813 2043 2847
rect 2729 2813 2763 2847
rect 2797 2813 2831 2847
rect 2865 2813 2899 2847
rect 3849 2813 3883 2847
rect 3917 2813 3951 2847
rect 3985 2813 4019 2847
rect 4505 2813 4539 2847
rect 4573 2813 4607 2847
rect 4641 2813 4675 2847
rect 4961 2813 4995 2847
rect 5029 2813 5063 2847
rect 5097 2813 5131 2847
rect 5417 2813 5451 2847
rect 5485 2813 5519 2847
rect 5553 2813 5587 2847
rect 4437 642 4471 676
rect 4505 642 4539 676
rect 4573 642 4607 676
rect 4641 642 4675 676
rect 4709 642 4743 676
rect 4893 642 4927 676
rect 4961 642 4995 676
rect 5029 642 5063 676
rect 5097 642 5131 676
rect 5165 642 5199 676
rect 5349 642 5383 676
rect 5417 642 5451 676
rect 5485 642 5519 676
rect 5553 642 5587 676
rect 5621 642 5655 676
<< locali >>
rect 9783 34796 14445 34802
rect 9783 34762 9795 34796
rect 9829 34762 9867 34796
rect 9901 34762 9917 34796
rect 9973 34762 9985 34796
rect 10045 34762 10053 34796
rect 10117 34762 10121 34796
rect 10223 34762 10227 34796
rect 10291 34762 10299 34796
rect 10359 34762 10371 34796
rect 10427 34762 10443 34796
rect 10495 34762 10515 34796
rect 10563 34762 10587 34796
rect 10631 34762 10659 34796
rect 10699 34762 10731 34796
rect 10767 34762 10801 34796
rect 10837 34762 10869 34796
rect 10909 34762 10937 34796
rect 10981 34762 11005 34796
rect 11053 34762 11073 34796
rect 11125 34762 11141 34796
rect 11197 34762 11209 34796
rect 11269 34762 11277 34796
rect 11341 34762 11345 34796
rect 11447 34762 11451 34796
rect 11515 34762 11523 34796
rect 11583 34762 11595 34796
rect 11651 34762 11667 34796
rect 11719 34762 11739 34796
rect 11787 34762 11811 34796
rect 11855 34762 11883 34796
rect 11923 34762 11955 34796
rect 11991 34762 12025 34796
rect 12061 34762 12093 34796
rect 12133 34762 12161 34796
rect 12205 34762 12229 34796
rect 12277 34762 12297 34796
rect 12349 34762 12365 34796
rect 12421 34762 12433 34796
rect 12493 34762 12501 34796
rect 12565 34762 12569 34796
rect 12671 34762 12675 34796
rect 12739 34762 12747 34796
rect 12807 34762 12819 34796
rect 12875 34762 12891 34796
rect 12943 34762 12963 34796
rect 13011 34762 13035 34796
rect 13079 34762 13107 34796
rect 13147 34762 13179 34796
rect 13215 34762 13249 34796
rect 13285 34762 13317 34796
rect 13357 34762 13385 34796
rect 13429 34762 13453 34796
rect 13501 34762 13521 34796
rect 13573 34762 13589 34796
rect 13645 34762 13657 34796
rect 13717 34762 13725 34796
rect 13789 34762 13793 34796
rect 13895 34762 13899 34796
rect 13963 34762 13971 34796
rect 14031 34762 14043 34796
rect 14099 34762 14115 34796
rect 14167 34762 14187 34796
rect 14235 34762 14259 34796
rect 14303 34762 14331 34796
rect 14371 34790 14445 34796
rect 14371 34762 14405 34790
rect 9783 34756 14405 34762
rect 14439 34756 14445 34790
rect 9783 34728 9829 34756
rect 9783 34674 9789 34728
rect 9823 34674 9829 34728
rect 9783 34660 9829 34674
rect 9783 34602 9789 34660
rect 9823 34602 9829 34660
rect 9783 34592 9829 34602
rect 9783 34530 9789 34592
rect 9823 34530 9829 34592
rect 14399 34718 14445 34756
rect 14399 34670 14405 34718
rect 14439 34670 14445 34718
rect 14399 34646 14445 34670
rect 14399 34612 14405 34646
rect 14439 34612 14445 34646
rect 14399 34574 14445 34612
rect 9783 34524 9829 34530
rect 9783 34458 9789 34524
rect 9823 34458 9829 34524
rect 9783 34456 9829 34458
rect 9783 34422 9789 34456
rect 9823 34422 9829 34456
rect 9783 34420 9829 34422
rect 9783 34354 9789 34420
rect 9823 34354 9829 34420
rect 9783 34348 9829 34354
rect 9783 34286 9789 34348
rect 9823 34286 9829 34348
rect 9783 34276 9829 34286
rect 9783 34230 9789 34276
rect 9823 34230 9829 34276
rect 10034 34546 14199 34552
rect 10034 34512 10046 34546
rect 10080 34512 10118 34546
rect 10181 34512 10190 34546
rect 10249 34512 10262 34546
rect 10317 34512 10334 34546
rect 10385 34512 10406 34546
rect 10453 34512 10478 34546
rect 10521 34512 10550 34546
rect 10589 34512 10622 34546
rect 10657 34512 10691 34546
rect 10728 34512 10759 34546
rect 10800 34512 10827 34546
rect 10872 34512 10895 34546
rect 10944 34512 10963 34546
rect 11016 34512 11031 34546
rect 11088 34512 11099 34546
rect 11160 34512 11167 34546
rect 11232 34512 11235 34546
rect 11269 34512 11270 34546
rect 11337 34512 11342 34546
rect 11405 34512 11414 34546
rect 11473 34512 11486 34546
rect 11541 34512 11558 34546
rect 11609 34512 11630 34546
rect 11677 34512 11702 34546
rect 11745 34512 11774 34546
rect 11813 34512 11846 34546
rect 11881 34512 11915 34546
rect 11952 34512 11983 34546
rect 12024 34512 12051 34546
rect 12096 34512 12119 34546
rect 12168 34512 12187 34546
rect 12240 34512 12255 34546
rect 12312 34512 12323 34546
rect 12384 34512 12391 34546
rect 12456 34512 12459 34546
rect 12493 34512 12494 34546
rect 12561 34512 12566 34546
rect 12629 34512 12638 34546
rect 12697 34512 12710 34546
rect 12765 34512 12782 34546
rect 12833 34512 12854 34546
rect 12901 34512 12926 34546
rect 12969 34512 12998 34546
rect 13037 34512 13070 34546
rect 13105 34512 13139 34546
rect 13176 34512 13207 34546
rect 13248 34512 13275 34546
rect 13320 34512 13343 34546
rect 13392 34512 13411 34546
rect 13464 34512 13479 34546
rect 13536 34512 13547 34546
rect 13608 34512 13615 34546
rect 13680 34512 13683 34546
rect 13717 34512 13718 34546
rect 13785 34512 13790 34546
rect 13853 34512 13862 34546
rect 13921 34512 13934 34546
rect 13989 34512 14006 34546
rect 14057 34512 14078 34546
rect 14125 34540 14199 34546
rect 14125 34512 14159 34540
rect 10034 34506 14159 34512
rect 14193 34506 14199 34540
rect 10034 34478 10080 34506
rect 10034 34444 10040 34478
rect 10074 34444 10080 34478
rect 14153 34468 14199 34506
rect 10034 34420 10080 34444
rect 10207 34420 10219 34454
rect 10257 34420 10292 34454
rect 10331 34420 10365 34454
rect 10405 34420 10438 34454
rect 10479 34420 10510 34454
rect 10553 34420 10582 34454
rect 10626 34420 10665 34454
rect 10699 34420 10738 34454
rect 10772 34420 10811 34454
rect 10845 34420 10884 34454
rect 10918 34420 10957 34454
rect 10991 34420 11007 34454
rect 11063 34420 11079 34454
rect 11139 34420 11148 34454
rect 11212 34420 11217 34454
rect 11285 34420 11286 34454
rect 11320 34420 11324 34454
rect 11389 34420 11397 34454
rect 11458 34420 11470 34454
rect 11527 34420 11543 34454
rect 11596 34420 11616 34454
rect 11665 34420 11689 34454
rect 11734 34420 11762 34454
rect 11803 34420 11835 34454
rect 11872 34420 11907 34454
rect 11942 34420 11976 34454
rect 12015 34420 12045 34454
rect 12088 34420 12114 34454
rect 12161 34420 12183 34454
rect 12234 34420 12252 34454
rect 12307 34420 12321 34454
rect 12380 34420 12390 34454
rect 12453 34420 12459 34454
rect 12526 34420 12528 34454
rect 12562 34420 12565 34454
rect 12631 34420 12638 34454
rect 12700 34420 12711 34454
rect 12769 34420 12784 34454
rect 12838 34420 12857 34454
rect 12907 34420 12930 34454
rect 12976 34420 13003 34454
rect 13045 34420 13076 34454
rect 13114 34420 13149 34454
rect 13183 34420 13218 34454
rect 13256 34420 13287 34454
rect 13329 34420 13356 34454
rect 13402 34420 13425 34454
rect 13475 34420 13494 34454
rect 13548 34420 13563 34454
rect 13621 34420 13632 34454
rect 13694 34420 13701 34454
rect 13767 34420 13771 34454
rect 13805 34420 13806 34454
rect 13840 34420 13841 34454
rect 13875 34420 13880 34454
rect 13945 34420 13981 34454
rect 14015 34420 14031 34454
rect 14153 34434 14159 34468
rect 14193 34434 14199 34468
rect 10034 34376 10040 34420
rect 10074 34376 10080 34420
rect 10034 34348 10080 34376
rect 10034 34308 10040 34348
rect 10074 34308 10080 34348
rect 10034 34276 10080 34308
rect 10034 34240 10040 34276
rect 10074 34240 10080 34276
rect 10034 34230 10080 34240
rect 14153 34396 14199 34434
rect 14153 34351 14159 34396
rect 14193 34351 14199 34396
rect 14153 34324 14199 34351
rect 14153 34283 14159 34324
rect 14193 34283 14199 34324
rect 14153 34252 14199 34283
rect 9789 34184 9823 34218
rect 9789 34116 9823 34150
rect 9789 34048 9823 34082
rect 9789 33980 9823 34014
rect 9789 33912 9823 33946
rect 9789 33844 9823 33878
rect 9789 33776 9823 33810
rect 9789 33647 9823 33742
rect 10040 34206 10074 34230
rect 10040 34138 10074 34172
rect 10040 34070 10074 34104
rect 10040 34002 10074 34036
rect 10040 33934 10074 33968
rect 10040 33866 10074 33900
rect 10040 33798 10074 33832
rect 10040 33730 10074 33764
rect 10040 33662 10074 33696
rect 9119 33613 9153 33647
rect 9119 33545 9153 33579
rect 9119 33477 9153 33511
rect 10034 33628 10040 33656
rect 14153 34215 14159 34252
rect 14193 34215 14199 34252
rect 14153 34181 14199 34215
rect 14153 34146 14159 34181
rect 14193 34146 14199 34181
rect 14153 34113 14199 34146
rect 14153 34074 14159 34113
rect 14193 34074 14199 34113
rect 14153 34045 14199 34074
rect 14153 34002 14159 34045
rect 14193 34002 14199 34045
rect 14153 33977 14199 34002
rect 14153 33930 14159 33977
rect 14193 33930 14199 33977
rect 14153 33909 14199 33930
rect 14153 33858 14159 33909
rect 14193 33858 14199 33909
rect 14153 33841 14199 33858
rect 14153 33786 14159 33841
rect 14193 33786 14199 33841
rect 14153 33773 14199 33786
rect 14153 33714 14159 33773
rect 14193 33714 14199 33773
rect 14153 33705 14199 33714
rect 10074 33628 10080 33656
rect 10034 33596 10080 33628
rect 10034 33560 10040 33596
rect 10074 33560 10080 33596
rect 14153 33642 14159 33705
rect 14193 33642 14199 33705
rect 14153 33637 14199 33642
rect 14153 33570 14159 33637
rect 14193 33570 14199 33637
rect 14153 33569 14199 33570
rect 10034 33526 10080 33560
rect 10034 33490 10040 33526
rect 10074 33490 10080 33526
rect 9119 33409 9153 33443
rect 9119 33341 9153 33375
rect 9119 33273 9153 33307
rect 9119 33205 9153 33239
rect 9119 33137 9153 33171
rect 9119 33069 9153 33103
rect 9119 33001 9153 33035
rect 9119 32933 9153 32967
rect 9119 32865 9153 32899
rect 9119 32797 9153 32831
rect 9119 32729 9153 32763
rect 9119 32661 9153 32695
rect 9119 32593 9153 32627
rect 9119 32525 9153 32559
rect 9119 32457 9153 32491
rect 9420 33453 9842 33487
rect 9420 33414 9876 33453
rect 9420 33380 9842 33414
rect 9420 33341 9876 33380
rect 9420 33307 9842 33341
rect 9420 33267 9876 33307
rect 9420 33233 9842 33267
rect 9420 33193 9876 33233
rect 9420 32467 9842 33193
rect 10034 33458 10080 33490
rect 10034 33418 10040 33458
rect 10074 33418 10080 33458
rect 10034 33390 10080 33418
rect 10034 33346 10040 33390
rect 10074 33346 10080 33390
rect 10034 33322 10080 33346
rect 10034 33274 10040 33322
rect 10074 33274 10080 33322
rect 10034 33254 10080 33274
rect 10034 33202 10040 33254
rect 10074 33202 10080 33254
rect 10034 33186 10080 33202
rect 10034 33130 10040 33186
rect 10074 33130 10080 33186
rect 10162 33492 10196 33533
rect 10162 33417 10196 33458
rect 10162 33342 10196 33383
rect 10162 33267 10196 33308
rect 10162 33193 10196 33233
rect 11018 33492 11052 33533
rect 11018 33417 11052 33458
rect 11018 33342 11052 33383
rect 11018 33267 11052 33308
rect 11018 33193 11052 33233
rect 11874 33492 11908 33533
rect 11874 33417 11908 33458
rect 11874 33342 11908 33383
rect 11874 33267 11908 33308
rect 11874 33193 11908 33233
rect 12730 33492 12764 33533
rect 12730 33417 12764 33458
rect 12730 33342 12764 33383
rect 12730 33267 12764 33308
rect 12730 33193 12764 33233
rect 13586 33492 13620 33533
rect 13586 33417 13620 33458
rect 13586 33342 13620 33383
rect 13586 33267 13620 33308
rect 13586 33193 13620 33233
rect 14042 33492 14076 33533
rect 14042 33417 14076 33458
rect 14042 33342 14076 33383
rect 14042 33267 14076 33308
rect 14042 33193 14076 33233
rect 14153 33535 14159 33569
rect 14193 33535 14199 33569
rect 14153 33532 14199 33535
rect 14153 33467 14159 33532
rect 14193 33467 14199 33532
rect 14153 33452 14199 33467
rect 14153 33399 14159 33452
rect 14193 33399 14199 33452
rect 14153 33380 14199 33399
rect 14153 33331 14159 33380
rect 14193 33331 14199 33380
rect 14153 33308 14199 33331
rect 14153 33263 14159 33308
rect 14193 33263 14199 33308
rect 14153 33236 14199 33263
rect 14153 33195 14159 33236
rect 14193 33195 14199 33236
rect 14153 33164 14199 33195
rect 10034 33118 10080 33130
rect 10034 33058 10040 33118
rect 10074 33058 10080 33118
rect 10034 33050 10080 33058
rect 10034 32986 10040 33050
rect 10074 32986 10080 33050
rect 10034 32982 10080 32986
rect 10034 32880 10040 32982
rect 10074 32880 10080 32982
rect 10034 32876 10080 32880
rect 10034 32812 10040 32876
rect 10074 32812 10080 32876
rect 10034 32804 10080 32812
rect 10034 32744 10040 32804
rect 10074 32744 10080 32804
rect 10034 32732 10080 32744
rect 10034 32676 10040 32732
rect 10074 32676 10080 32732
rect 10034 32660 10080 32676
rect 10034 32608 10040 32660
rect 10074 32608 10080 32660
rect 10034 32588 10080 32608
rect 10034 32540 10040 32588
rect 10074 32540 10080 32588
rect 10034 32516 10080 32540
rect 10034 32472 10040 32516
rect 10074 32472 10080 32516
rect 9119 32389 9153 32423
rect 9119 32321 9153 32355
rect 9119 32253 9153 32287
rect 10034 32444 10080 32472
rect 10034 32404 10040 32444
rect 10074 32404 10080 32444
rect 10034 32372 10080 32404
rect 10034 32336 10040 32372
rect 10074 32336 10080 32372
rect 10034 32302 10080 32336
rect 10034 32266 10040 32302
rect 10074 32300 10080 32302
rect 14153 33127 14159 33164
rect 14193 33127 14199 33164
rect 14153 33093 14199 33127
rect 14153 33058 14159 33093
rect 14193 33058 14199 33093
rect 14153 33025 14199 33058
rect 14153 32986 14159 33025
rect 14193 32986 14199 33025
rect 14153 32957 14199 32986
rect 14153 32914 14159 32957
rect 14193 32914 14199 32957
rect 14153 32889 14199 32914
rect 14153 32842 14159 32889
rect 14193 32842 14199 32889
rect 14153 32821 14199 32842
rect 14153 32770 14159 32821
rect 14193 32770 14199 32821
rect 14153 32753 14199 32770
rect 14153 32698 14159 32753
rect 14193 32698 14199 32753
rect 14153 32685 14199 32698
rect 14153 32626 14159 32685
rect 14193 32626 14199 32685
rect 14153 32617 14199 32626
rect 14153 32554 14159 32617
rect 14193 32554 14199 32617
rect 14153 32549 14199 32554
rect 14153 32482 14159 32549
rect 14193 32482 14199 32549
rect 14153 32481 14199 32482
rect 14153 32447 14159 32481
rect 14193 32447 14199 32481
rect 14153 32444 14199 32447
rect 14153 32379 14159 32444
rect 14193 32379 14199 32444
rect 14153 32372 14199 32379
rect 14153 32311 14159 32372
rect 14193 32311 14199 32372
rect 14153 32300 14199 32311
rect 10074 32294 14159 32300
rect 10074 32266 10108 32294
rect 10034 32260 10108 32266
rect 10146 32260 10185 32294
rect 10227 32260 10258 32294
rect 10312 32260 10331 32294
rect 10397 32260 10404 32294
rect 10438 32260 10448 32294
rect 10511 32260 10533 32294
rect 10584 32260 10618 32294
rect 10657 32260 10696 32294
rect 10737 32260 10769 32294
rect 10822 32260 10842 32294
rect 10907 32260 10915 32294
rect 10949 32260 10958 32294
rect 11022 32260 11043 32294
rect 11095 32260 11128 32294
rect 11168 32260 11207 32294
rect 11247 32260 11279 32294
rect 11332 32260 11351 32294
rect 11417 32260 11423 32294
rect 11457 32260 11468 32294
rect 11529 32260 11553 32294
rect 11601 32260 11638 32294
rect 11673 32260 11711 32294
rect 11757 32260 11783 32294
rect 11842 32260 11855 32294
rect 11889 32260 11893 32294
rect 11961 32260 11978 32294
rect 12033 32260 12063 32294
rect 12105 32260 12143 32294
rect 12182 32260 12215 32294
rect 12267 32260 12287 32294
rect 12352 32260 12359 32294
rect 12393 32260 12403 32294
rect 12465 32260 12488 32294
rect 12537 32260 12573 32294
rect 12609 32260 12647 32294
rect 12692 32260 12719 32294
rect 12777 32260 12791 32294
rect 12825 32260 12828 32294
rect 12862 32260 12863 32294
rect 12897 32260 12913 32294
rect 12969 32260 12998 32294
rect 13041 32260 13079 32294
rect 13117 32260 13151 32294
rect 13201 32260 13223 32294
rect 13285 32260 13295 32294
rect 13329 32260 13335 32294
rect 13401 32260 13419 32294
rect 13473 32260 13503 32294
rect 13545 32260 13583 32294
rect 13621 32260 13655 32294
rect 13705 32260 13727 32294
rect 13789 32260 13799 32294
rect 13833 32260 13839 32294
rect 13905 32260 13923 32294
rect 13977 32260 14007 32294
rect 14049 32260 14087 32294
rect 14125 32260 14159 32294
rect 10034 32254 14159 32260
rect 9119 32185 9153 32219
rect 10040 32234 10074 32254
rect 9119 32117 9153 32151
rect 9119 32049 9153 32083
rect 9119 31981 9153 32015
rect 9119 31913 9153 31947
rect 9119 31845 9153 31879
rect 9119 31777 9153 31811
rect 9119 31709 9153 31743
rect 9119 31641 9153 31675
rect 9119 31573 9153 31607
rect 9119 31505 9153 31539
rect 9119 31437 9153 31471
rect 9568 32168 9611 32202
rect 9645 32168 9688 32202
rect 9534 31435 9722 32168
rect 14153 32243 14159 32254
rect 14193 32243 14199 32300
rect 14153 32228 14199 32243
rect 10040 32166 10074 32200
rect 10207 32168 10219 32202
rect 10257 32168 10297 32202
rect 10338 32168 10371 32202
rect 10423 32168 10445 32202
rect 10508 32168 10519 32202
rect 10553 32168 10559 32202
rect 10626 32168 10643 32202
rect 10699 32168 10738 32202
rect 10772 32168 10811 32202
rect 10845 32168 10884 32202
rect 10918 32168 10957 32202
rect 10991 32168 11007 32202
rect 11063 32168 11079 32202
rect 11139 32168 11148 32202
rect 11212 32168 11217 32202
rect 11285 32168 11286 32202
rect 11320 32168 11324 32202
rect 11389 32168 11397 32202
rect 11458 32168 11470 32202
rect 11527 32168 11543 32202
rect 11596 32168 11616 32202
rect 11665 32168 11689 32202
rect 11734 32168 11762 32202
rect 11803 32168 11835 32202
rect 11872 32168 11907 32202
rect 11942 32168 11976 32202
rect 12015 32168 12045 32202
rect 12088 32168 12114 32202
rect 12161 32168 12183 32202
rect 12234 32168 12252 32202
rect 12307 32168 12321 32202
rect 12380 32168 12390 32202
rect 12453 32168 12459 32202
rect 12526 32168 12528 32202
rect 12562 32168 12565 32202
rect 12631 32168 12638 32202
rect 12700 32168 12711 32202
rect 12769 32168 12784 32202
rect 12838 32168 12857 32202
rect 12907 32168 12930 32202
rect 12976 32168 13003 32202
rect 13045 32168 13076 32202
rect 13114 32168 13149 32202
rect 13183 32168 13218 32202
rect 13256 32168 13287 32202
rect 13329 32168 13356 32202
rect 13402 32168 13425 32202
rect 13475 32168 13494 32202
rect 13548 32168 13563 32202
rect 13621 32168 13632 32202
rect 13694 32168 13701 32202
rect 13767 32168 13771 32202
rect 13805 32168 13806 32202
rect 13840 32168 13841 32202
rect 13875 32168 13880 32202
rect 13945 32168 13981 32202
rect 14015 32168 14031 32202
rect 14153 32175 14159 32228
rect 14193 32175 14199 32228
rect 10040 32098 10074 32132
rect 10040 32030 10074 32064
rect 10040 31962 10074 31996
rect 10040 31894 10074 31928
rect 10040 31826 10074 31860
rect 10040 31758 10074 31792
rect 10040 31690 10074 31724
rect 10040 31622 10074 31656
rect 10034 31588 10040 31621
rect 14153 32156 14199 32175
rect 14153 32107 14159 32156
rect 14193 32107 14199 32156
rect 14153 32084 14199 32107
rect 14153 32039 14159 32084
rect 14193 32039 14199 32084
rect 14153 32012 14199 32039
rect 14153 31971 14159 32012
rect 14193 31971 14199 32012
rect 14153 31940 14199 31971
rect 14153 31903 14159 31940
rect 14193 31903 14199 31940
rect 14153 31869 14199 31903
rect 14153 31834 14159 31869
rect 14193 31834 14199 31869
rect 14153 31801 14199 31834
rect 14153 31762 14159 31801
rect 14193 31762 14199 31801
rect 14153 31733 14199 31762
rect 14153 31690 14159 31733
rect 14193 31690 14199 31733
rect 14153 31665 14199 31690
rect 10074 31588 10080 31621
rect 10034 31578 10080 31588
rect 10034 31520 10040 31578
rect 10074 31520 10080 31578
rect 10034 31506 10080 31520
rect 10034 31452 10040 31506
rect 10074 31452 10080 31506
rect 9119 31369 9153 31403
rect 9431 31401 9447 31435
rect 9481 31401 9531 31435
rect 9565 31401 9615 31435
rect 9649 31401 9698 31435
rect 9732 31401 9781 31435
rect 9815 31401 9831 31435
rect 10034 31434 10080 31452
rect 9119 31301 9153 31335
rect 9119 31184 9153 31267
rect 10034 31384 10040 31434
rect 10074 31384 10080 31434
rect 10034 31362 10080 31384
rect 10034 31316 10040 31362
rect 10074 31316 10080 31362
rect 10034 31290 10080 31316
rect 10034 31248 10040 31290
rect 10074 31248 10080 31290
rect 14153 31618 14159 31665
rect 14193 31618 14199 31665
rect 14153 31597 14199 31618
rect 14153 31546 14159 31597
rect 14193 31546 14199 31597
rect 14153 31529 14199 31546
rect 14153 31474 14159 31529
rect 14193 31474 14199 31529
rect 14153 31461 14199 31474
rect 14153 31402 14159 31461
rect 14193 31402 14199 31461
rect 14153 31393 14199 31402
rect 14153 31330 14159 31393
rect 14193 31330 14199 31393
rect 14153 31325 14199 31330
rect 10034 31218 10080 31248
rect 9783 31150 9829 31184
rect 9783 31112 9789 31150
rect 9823 31112 9829 31150
rect 9783 31082 9829 31112
rect 9783 31040 9789 31082
rect 9823 31040 9829 31082
rect 9783 31014 9829 31040
rect 9783 30968 9789 31014
rect 9823 30968 9829 31014
rect 9783 30946 9829 30968
rect 9783 30896 9789 30946
rect 9823 30896 9829 30946
rect 9783 30878 9829 30896
rect 9783 30824 9789 30878
rect 9823 30824 9829 30878
rect 9783 30812 9829 30824
rect 10034 31180 10040 31218
rect 10074 31180 10080 31218
rect 10034 31146 10080 31180
rect 10034 31112 10040 31146
rect 10074 31112 10080 31146
rect 10034 31078 10080 31112
rect 10034 31040 10040 31078
rect 10074 31040 10080 31078
rect 10034 31010 10080 31040
rect 10034 30968 10040 31010
rect 10074 30968 10080 31010
rect 10034 30942 10080 30968
rect 10034 30896 10040 30942
rect 10074 30896 10080 30942
rect 10034 30874 10080 30896
rect 10162 31207 10196 31248
rect 10162 31132 10196 31173
rect 10162 31057 10196 31098
rect 10162 30982 10196 31023
rect 10162 30908 10196 30948
rect 11018 31207 11052 31248
rect 11018 31132 11052 31173
rect 11018 31057 11052 31098
rect 11018 30982 11052 31023
rect 11018 30908 11052 30948
rect 11874 31207 11908 31248
rect 11874 31132 11908 31173
rect 11874 31057 11908 31098
rect 11874 30982 11908 31023
rect 11874 30908 11908 30948
rect 12730 31207 12764 31248
rect 12730 31132 12764 31173
rect 12730 31057 12764 31098
rect 12730 30982 12764 31023
rect 12730 30908 12764 30948
rect 13586 31207 13620 31248
rect 13586 31132 13620 31173
rect 13586 31057 13620 31098
rect 13586 30982 13620 31023
rect 13586 30908 13620 30948
rect 14042 31207 14076 31248
rect 14042 31132 14076 31173
rect 14042 31057 14076 31098
rect 14042 30982 14076 31023
rect 14042 30908 14076 30948
rect 14153 31258 14159 31325
rect 14193 31258 14199 31325
rect 14153 31257 14199 31258
rect 14153 31223 14159 31257
rect 14193 31223 14199 31257
rect 14153 31220 14199 31223
rect 14153 31155 14159 31220
rect 14193 31155 14199 31220
rect 14153 31148 14199 31155
rect 14153 31087 14159 31148
rect 14193 31087 14199 31148
rect 14153 31076 14199 31087
rect 14153 31019 14159 31076
rect 14193 31019 14199 31076
rect 14153 31004 14199 31019
rect 14153 30951 14159 31004
rect 14193 30951 14199 31004
rect 14153 30932 14199 30951
rect 14153 30883 14159 30932
rect 14193 30883 14199 30932
rect 10034 30824 10040 30874
rect 10074 30824 10080 30874
rect 10034 30812 10080 30824
rect 14153 30860 14199 30883
rect 14153 30815 14159 30860
rect 14193 30815 14199 30860
rect 9789 30810 9823 30812
rect 9789 30742 9823 30776
rect 9789 30674 9823 30708
rect 9789 30606 9823 30640
rect 9789 30538 9823 30572
rect 9789 30470 9823 30504
rect 9789 30402 9823 30436
rect 9789 30334 9823 30368
rect 9789 30266 9823 30300
rect 9789 30198 9823 30232
rect 9789 30148 9823 30164
rect 10040 30806 10074 30812
rect 10040 30738 10074 30772
rect 10040 30670 10074 30704
rect 10040 30602 10074 30636
rect 10040 30534 10074 30568
rect 10040 30466 10074 30500
rect 10040 30398 10074 30432
rect 10040 30330 10074 30364
rect 10040 30262 10074 30296
rect 10040 30194 10074 30228
rect 10040 30148 10074 30160
rect 14153 30788 14199 30815
rect 14153 30747 14159 30788
rect 14193 30747 14199 30788
rect 14153 30716 14199 30747
rect 14153 30679 14159 30716
rect 14193 30679 14199 30716
rect 14153 30645 14199 30679
rect 14153 30610 14159 30645
rect 14193 30610 14199 30645
rect 14153 30577 14199 30610
rect 14153 30538 14159 30577
rect 14193 30538 14199 30577
rect 14153 30509 14199 30538
rect 14153 30466 14159 30509
rect 14193 30466 14199 30509
rect 14153 30441 14199 30466
rect 14153 30394 14159 30441
rect 14193 30394 14199 30441
rect 14153 30373 14199 30394
rect 14153 30322 14159 30373
rect 14193 30322 14199 30373
rect 14153 30305 14199 30322
rect 14153 30250 14159 30305
rect 14193 30250 14199 30305
rect 14153 30237 14199 30250
rect 14153 30178 14159 30237
rect 14193 30178 14199 30237
rect 14153 30169 14199 30178
rect 9783 30130 9829 30148
rect 9783 30028 9789 30130
rect 9823 30028 9829 30130
rect 9783 30024 9829 30028
rect 9783 29960 9789 30024
rect 9823 29960 9829 30024
rect 9783 29952 9829 29960
rect 9783 29892 9789 29952
rect 9823 29892 9829 29952
rect 9783 29880 9829 29892
rect 9783 29824 9789 29880
rect 9823 29824 9829 29880
rect 9783 29808 9829 29824
rect 9783 29756 9789 29808
rect 9823 29756 9829 29808
rect 9783 29736 9829 29756
rect 9783 29690 9789 29736
rect 9823 29690 9829 29736
rect 10034 30126 10080 30148
rect 10034 30062 10040 30126
rect 10074 30062 10080 30126
rect 10034 30058 10080 30062
rect 10034 29956 10040 30058
rect 10074 30049 10080 30058
rect 14153 30106 14159 30169
rect 14193 30106 14199 30169
rect 14153 30101 14199 30106
rect 14153 30049 14159 30101
rect 10074 30043 14159 30049
rect 10074 30009 10108 30043
rect 10146 30009 10185 30043
rect 10227 30009 10258 30043
rect 10312 30009 10331 30043
rect 10397 30009 10404 30043
rect 10438 30009 10448 30043
rect 10511 30009 10533 30043
rect 10584 30009 10618 30043
rect 10657 30009 10696 30043
rect 10737 30009 10769 30043
rect 10822 30009 10842 30043
rect 10907 30009 10915 30043
rect 10949 30009 10958 30043
rect 11022 30009 11043 30043
rect 11095 30009 11128 30043
rect 11168 30009 11207 30043
rect 11247 30009 11279 30043
rect 11332 30009 11351 30043
rect 11417 30009 11423 30043
rect 11457 30009 11468 30043
rect 11529 30009 11553 30043
rect 11601 30009 11638 30043
rect 11673 30009 11711 30043
rect 11757 30009 11783 30043
rect 11842 30009 11855 30043
rect 11889 30009 11893 30043
rect 11961 30009 11978 30043
rect 12033 30009 12063 30043
rect 12105 30009 12143 30043
rect 12182 30009 12215 30043
rect 12267 30009 12287 30043
rect 12352 30009 12359 30043
rect 12393 30009 12403 30043
rect 12465 30009 12488 30043
rect 12537 30009 12573 30043
rect 12609 30009 12647 30043
rect 12692 30009 12719 30043
rect 12777 30009 12791 30043
rect 12825 30009 12828 30043
rect 12862 30009 12863 30043
rect 12897 30009 12913 30043
rect 12969 30009 12998 30043
rect 13041 30009 13079 30043
rect 13117 30009 13151 30043
rect 13201 30009 13223 30043
rect 13285 30009 13295 30043
rect 13329 30009 13335 30043
rect 13401 30009 13419 30043
rect 13473 30009 13503 30043
rect 13545 30009 13583 30043
rect 13621 30009 13655 30043
rect 13705 30009 13727 30043
rect 13789 30009 13799 30043
rect 13833 30009 13839 30043
rect 13905 30009 13923 30043
rect 13977 30009 14007 30043
rect 14049 30009 14087 30043
rect 14125 30034 14159 30043
rect 14193 30034 14199 30101
rect 14125 30033 14199 30034
rect 14125 30009 14159 30033
rect 10074 30003 14159 30009
rect 10074 29956 10080 30003
rect 10034 29952 10080 29956
rect 14153 29999 14159 30003
rect 14193 29999 14199 30033
rect 14153 29996 14199 29999
rect 10034 29888 10040 29952
rect 10074 29888 10080 29952
rect 10207 29919 10219 29953
rect 10257 29919 10297 29953
rect 10338 29919 10371 29953
rect 10423 29919 10445 29953
rect 10508 29919 10519 29953
rect 10553 29919 10559 29953
rect 10626 29919 10643 29953
rect 10699 29919 10738 29953
rect 10772 29919 10811 29953
rect 10845 29919 10884 29953
rect 10918 29919 10957 29953
rect 10991 29919 11007 29953
rect 11063 29919 11079 29953
rect 11139 29919 11148 29953
rect 11212 29919 11217 29953
rect 11285 29919 11286 29953
rect 11320 29919 11324 29953
rect 11389 29919 11397 29953
rect 11458 29919 11470 29953
rect 11527 29919 11543 29953
rect 11596 29919 11616 29953
rect 11665 29919 11689 29953
rect 11734 29919 11762 29953
rect 11803 29919 11835 29953
rect 11872 29919 11907 29953
rect 11942 29919 11976 29953
rect 12015 29919 12045 29953
rect 12088 29919 12114 29953
rect 12161 29919 12183 29953
rect 12234 29919 12252 29953
rect 12307 29919 12321 29953
rect 12380 29919 12390 29953
rect 12453 29919 12459 29953
rect 12526 29919 12528 29953
rect 12562 29919 12565 29953
rect 12631 29919 12638 29953
rect 12700 29919 12711 29953
rect 12769 29919 12784 29953
rect 12838 29919 12857 29953
rect 12907 29919 12930 29953
rect 12976 29919 13003 29953
rect 13045 29919 13076 29953
rect 13114 29919 13149 29953
rect 13183 29919 13218 29953
rect 13256 29919 13287 29953
rect 13329 29919 13356 29953
rect 13402 29919 13425 29953
rect 13475 29919 13494 29953
rect 13548 29919 13563 29953
rect 13621 29919 13632 29953
rect 13694 29919 13701 29953
rect 13767 29919 13771 29953
rect 13805 29919 13806 29953
rect 13840 29919 13841 29953
rect 13875 29919 13880 29953
rect 13945 29919 13981 29953
rect 14015 29919 14031 29953
rect 14153 29931 14159 29996
rect 14193 29931 14199 29996
rect 14153 29924 14199 29931
rect 10034 29880 10080 29888
rect 10034 29820 10040 29880
rect 10074 29820 10080 29880
rect 10034 29808 10080 29820
rect 10034 29752 10040 29808
rect 10074 29752 10080 29808
rect 10034 29736 10080 29752
rect 10034 29690 10040 29736
rect 9789 29654 9823 29688
rect 9789 29586 9823 29620
rect 9789 29518 9823 29552
rect 9789 29450 9823 29484
rect 9789 29382 9823 29416
rect 9789 29314 9823 29348
rect 9789 29246 9823 29280
rect 9789 29178 9823 29212
rect 9789 29110 9823 29144
rect 9789 29042 9823 29076
rect 9789 28974 9823 29008
rect 10074 29690 10080 29736
rect 14153 29863 14159 29924
rect 14193 29863 14199 29924
rect 14153 29852 14199 29863
rect 14153 29795 14159 29852
rect 14193 29795 14199 29852
rect 14153 29780 14199 29795
rect 14153 29727 14159 29780
rect 14193 29727 14199 29780
rect 14153 29708 14199 29727
rect 10040 29650 10074 29684
rect 10040 29582 10074 29616
rect 10040 29514 10074 29548
rect 10040 29446 10074 29480
rect 10040 29378 10074 29412
rect 10040 29310 10074 29344
rect 10040 29242 10074 29276
rect 10040 29174 10074 29208
rect 10040 29106 10074 29140
rect 10040 29038 10074 29072
rect 10040 28991 10074 29004
rect 14153 29659 14159 29708
rect 14193 29659 14199 29708
rect 14153 29636 14199 29659
rect 14153 29591 14159 29636
rect 14193 29591 14199 29636
rect 14153 29564 14199 29591
rect 14153 29523 14159 29564
rect 14193 29523 14199 29564
rect 14153 29492 14199 29523
rect 14153 29455 14159 29492
rect 14193 29455 14199 29492
rect 14153 29421 14199 29455
rect 14153 29386 14159 29421
rect 14193 29386 14199 29421
rect 14153 29353 14199 29386
rect 14153 29314 14159 29353
rect 14193 29314 14199 29353
rect 14153 29285 14199 29314
rect 14153 29242 14159 29285
rect 14193 29242 14199 29285
rect 14153 29217 14199 29242
rect 14153 29170 14159 29217
rect 14193 29170 14199 29217
rect 14153 29149 14199 29170
rect 14153 29098 14159 29149
rect 14193 29098 14199 29149
rect 14153 29081 14199 29098
rect 14153 29026 14159 29081
rect 14193 29026 14199 29081
rect 14153 29013 14199 29026
rect 9789 28906 9823 28940
rect 9789 28838 9823 28872
rect 9789 28770 9823 28804
rect 9789 28702 9823 28736
rect 9789 28634 9823 28668
rect 9789 28566 9823 28600
rect 9789 28498 9823 28532
rect 9789 28430 9823 28464
rect 9789 28362 9823 28396
rect 9789 28294 9823 28328
rect 9789 28226 9823 28260
rect 9789 28158 9823 28192
rect 9789 28090 9823 28124
rect 9789 28022 9823 28056
rect 10034 28970 10080 28991
rect 10034 28936 10040 28970
rect 10074 28936 10080 28970
rect 10034 28932 10080 28936
rect 10034 28868 10040 28932
rect 10074 28868 10080 28932
rect 10034 28860 10080 28868
rect 10034 28800 10040 28860
rect 10074 28800 10080 28860
rect 10034 28788 10080 28800
rect 10034 28732 10040 28788
rect 10074 28732 10080 28788
rect 10034 28716 10080 28732
rect 10034 28664 10040 28716
rect 10074 28664 10080 28716
rect 10034 28644 10080 28664
rect 10034 28596 10040 28644
rect 10074 28596 10080 28644
rect 10034 28572 10080 28596
rect 10034 28528 10040 28572
rect 10074 28528 10080 28572
rect 10162 28903 10196 28944
rect 10162 28828 10196 28869
rect 10162 28753 10196 28794
rect 10162 28678 10196 28719
rect 10162 28604 10196 28644
rect 11018 28903 11052 28944
rect 11018 28828 11052 28869
rect 11018 28753 11052 28794
rect 11018 28678 11052 28719
rect 11018 28604 11052 28644
rect 11874 28903 11908 28944
rect 11874 28828 11908 28869
rect 11874 28753 11908 28794
rect 11874 28678 11908 28719
rect 11874 28604 11908 28644
rect 12730 28903 12764 28944
rect 12730 28828 12764 28869
rect 12730 28753 12764 28794
rect 12730 28678 12764 28719
rect 12730 28604 12764 28644
rect 13586 28903 13620 28944
rect 13586 28828 13620 28869
rect 13586 28753 13620 28794
rect 13586 28678 13620 28719
rect 13586 28604 13620 28644
rect 14042 28903 14076 28944
rect 14042 28828 14076 28869
rect 14042 28753 14076 28794
rect 14042 28678 14076 28719
rect 14042 28604 14076 28644
rect 14153 28954 14159 29013
rect 14193 28954 14199 29013
rect 14153 28945 14199 28954
rect 14153 28882 14159 28945
rect 14193 28882 14199 28945
rect 14153 28877 14199 28882
rect 14153 28810 14159 28877
rect 14193 28810 14199 28877
rect 14153 28809 14199 28810
rect 14153 28775 14159 28809
rect 14193 28775 14199 28809
rect 14153 28772 14199 28775
rect 14153 28707 14159 28772
rect 14193 28707 14199 28772
rect 14153 28700 14199 28707
rect 14153 28639 14159 28700
rect 14193 28639 14199 28700
rect 14153 28628 14199 28639
rect 14153 28571 14159 28628
rect 14193 28571 14199 28628
rect 10034 28500 10080 28528
rect 10034 28460 10040 28500
rect 10074 28460 10080 28500
rect 10034 28428 10080 28460
rect 10034 28392 10040 28428
rect 10074 28392 10080 28428
rect 10034 28358 10080 28392
rect 10034 28322 10040 28358
rect 10074 28322 10080 28358
rect 10034 28290 10080 28322
rect 10034 28250 10040 28290
rect 10074 28250 10080 28290
rect 10034 28222 10080 28250
rect 10034 28178 10040 28222
rect 10074 28178 10080 28222
rect 10034 28154 10080 28178
rect 10034 28106 10040 28154
rect 10074 28106 10080 28154
rect 10034 28086 10080 28106
rect 10034 28034 10040 28086
rect 10074 28034 10080 28086
rect 10034 28022 10080 28034
rect 14153 28556 14199 28571
rect 14153 28503 14159 28556
rect 14193 28503 14199 28556
rect 14153 28484 14199 28503
rect 14153 28435 14159 28484
rect 14193 28435 14199 28484
rect 14153 28412 14199 28435
rect 14153 28367 14159 28412
rect 14193 28367 14199 28412
rect 14153 28340 14199 28367
rect 14153 28299 14159 28340
rect 14193 28299 14199 28340
rect 14153 28268 14199 28299
rect 14153 28231 14159 28268
rect 14193 28231 14199 28268
rect 14153 28197 14199 28231
rect 14153 28162 14159 28197
rect 14193 28162 14199 28197
rect 14153 28129 14199 28162
rect 14153 28090 14159 28129
rect 14193 28090 14199 28129
rect 14153 28061 14199 28090
rect 9789 27954 9823 27988
rect 9789 27886 9823 27920
rect 9789 27818 9823 27852
rect 10040 28018 10074 28022
rect 10040 27950 10074 27984
rect 10040 27882 10074 27916
rect 10040 27795 10074 27848
rect 14153 28018 14159 28061
rect 14193 28018 14199 28061
rect 14153 27993 14199 28018
rect 14153 27946 14159 27993
rect 14193 27946 14199 27993
rect 14153 27925 14199 27946
rect 14153 27874 14159 27925
rect 14193 27874 14199 27925
rect 14153 27857 14199 27874
rect 14153 27823 14159 27857
rect 14193 27823 14199 27857
rect 14153 27795 14199 27823
rect 9789 27750 9823 27784
rect 10034 27789 14199 27795
rect 10034 27755 10049 27789
rect 10083 27755 10108 27789
rect 10155 27755 10176 27789
rect 10227 27755 10244 27789
rect 10299 27755 10312 27789
rect 10371 27755 10380 27789
rect 10443 27755 10448 27789
rect 10515 27755 10516 27789
rect 10550 27755 10553 27789
rect 10618 27755 10625 27789
rect 10686 27755 10697 27789
rect 10754 27755 10769 27789
rect 10822 27755 10841 27789
rect 10890 27755 10913 27789
rect 10958 27755 10985 27789
rect 11026 27755 11057 27789
rect 11094 27755 11128 27789
rect 11163 27755 11196 27789
rect 11235 27755 11264 27789
rect 11307 27755 11332 27789
rect 11379 27755 11400 27789
rect 11451 27755 11468 27789
rect 11523 27755 11536 27789
rect 11595 27755 11604 27789
rect 11667 27755 11672 27789
rect 11739 27755 11740 27789
rect 11774 27755 11777 27789
rect 11842 27755 11849 27789
rect 11910 27755 11921 27789
rect 11978 27755 11993 27789
rect 12046 27755 12065 27789
rect 12114 27755 12137 27789
rect 12182 27755 12209 27789
rect 12250 27755 12281 27789
rect 12318 27755 12352 27789
rect 12387 27755 12420 27789
rect 12459 27755 12488 27789
rect 12531 27755 12556 27789
rect 12603 27755 12624 27789
rect 12675 27755 12692 27789
rect 12747 27755 12760 27789
rect 12819 27755 12828 27789
rect 12891 27755 12896 27789
rect 12963 27755 12964 27789
rect 12998 27755 13001 27789
rect 13066 27755 13073 27789
rect 13134 27755 13145 27789
rect 13202 27755 13217 27789
rect 13270 27755 13289 27789
rect 13338 27755 13361 27789
rect 13406 27755 13433 27789
rect 13474 27755 13505 27789
rect 13542 27755 13576 27789
rect 13611 27755 13644 27789
rect 13683 27755 13712 27789
rect 13755 27755 13780 27789
rect 13827 27755 13848 27789
rect 13899 27755 13916 27789
rect 13971 27755 13984 27789
rect 14043 27755 14052 27789
rect 14115 27755 14153 27789
rect 14187 27755 14199 27789
rect 10034 27749 14199 27755
rect 14399 34506 14405 34574
rect 14439 34506 14445 34574
rect 14399 34502 14445 34506
rect 14399 34438 14405 34502
rect 14439 34438 14445 34502
rect 14399 34430 14445 34438
rect 14399 34370 14405 34430
rect 14439 34370 14445 34430
rect 14399 34358 14445 34370
rect 14399 34302 14405 34358
rect 14439 34302 14445 34358
rect 14399 34286 14445 34302
rect 14399 34234 14405 34286
rect 14439 34234 14445 34286
rect 14399 34214 14445 34234
rect 14399 34166 14405 34214
rect 14439 34166 14445 34214
rect 14399 34142 14445 34166
rect 14399 34098 14405 34142
rect 14439 34098 14445 34142
rect 14399 34070 14445 34098
rect 14399 34030 14405 34070
rect 14439 34030 14445 34070
rect 14399 33998 14445 34030
rect 14399 33962 14405 33998
rect 14439 33962 14445 33998
rect 14399 33928 14445 33962
rect 14399 33892 14405 33928
rect 14439 33892 14445 33928
rect 14399 33860 14445 33892
rect 14399 33820 14405 33860
rect 14439 33820 14445 33860
rect 14399 33792 14445 33820
rect 14399 33748 14405 33792
rect 14439 33748 14445 33792
rect 14399 33724 14445 33748
rect 14399 33676 14405 33724
rect 14439 33676 14445 33724
rect 14399 33656 14445 33676
rect 14399 33604 14405 33656
rect 14439 33604 14445 33656
rect 14399 33588 14445 33604
rect 14399 33532 14405 33588
rect 14439 33532 14445 33588
rect 14399 33520 14445 33532
rect 14399 33460 14405 33520
rect 14439 33460 14445 33520
rect 14399 33452 14445 33460
rect 14399 33388 14405 33452
rect 14439 33388 14445 33452
rect 14399 33384 14445 33388
rect 14399 33282 14405 33384
rect 14439 33282 14445 33384
rect 14399 33278 14445 33282
rect 14399 33214 14405 33278
rect 14439 33214 14445 33278
rect 14399 33206 14445 33214
rect 14399 33146 14405 33206
rect 14439 33146 14445 33206
rect 14399 33134 14445 33146
rect 14399 33078 14405 33134
rect 14439 33078 14445 33134
rect 14399 33062 14445 33078
rect 14399 33010 14405 33062
rect 14439 33010 14445 33062
rect 14399 32990 14445 33010
rect 14399 32942 14405 32990
rect 14439 32942 14445 32990
rect 14399 32918 14445 32942
rect 14399 32874 14405 32918
rect 14439 32874 14445 32918
rect 14399 32846 14445 32874
rect 14399 32806 14405 32846
rect 14439 32806 14445 32846
rect 14399 32774 14445 32806
rect 14399 32738 14405 32774
rect 14439 32738 14445 32774
rect 14399 32704 14445 32738
rect 14399 32668 14405 32704
rect 14439 32668 14445 32704
rect 14399 32636 14445 32668
rect 14399 32596 14405 32636
rect 14439 32596 14445 32636
rect 14399 32568 14445 32596
rect 14399 32524 14405 32568
rect 14439 32524 14445 32568
rect 14399 32500 14445 32524
rect 14399 32452 14405 32500
rect 14439 32452 14445 32500
rect 14399 32432 14445 32452
rect 14399 32380 14405 32432
rect 14439 32380 14445 32432
rect 14399 32364 14445 32380
rect 14399 32308 14405 32364
rect 14439 32308 14445 32364
rect 14399 32296 14445 32308
rect 14399 32236 14405 32296
rect 14439 32236 14445 32296
rect 14399 32228 14445 32236
rect 14399 32164 14405 32228
rect 14439 32164 14445 32228
rect 14399 32160 14445 32164
rect 14399 32058 14405 32160
rect 14439 32058 14445 32160
rect 14399 32054 14445 32058
rect 14399 31990 14405 32054
rect 14439 31990 14445 32054
rect 14399 31982 14445 31990
rect 14399 31922 14405 31982
rect 14439 31922 14445 31982
rect 14399 31910 14445 31922
rect 14399 31854 14405 31910
rect 14439 31854 14445 31910
rect 14399 31838 14445 31854
rect 14399 31786 14405 31838
rect 14439 31786 14445 31838
rect 14399 31766 14445 31786
rect 14399 31718 14405 31766
rect 14439 31718 14445 31766
rect 14399 31694 14445 31718
rect 14399 31650 14405 31694
rect 14439 31650 14445 31694
rect 14399 31622 14445 31650
rect 14399 31582 14405 31622
rect 14439 31582 14445 31622
rect 14399 31550 14445 31582
rect 14399 31514 14405 31550
rect 14439 31514 14445 31550
rect 14399 31480 14445 31514
rect 14399 31444 14405 31480
rect 14439 31444 14445 31480
rect 14399 31412 14445 31444
rect 14399 31372 14405 31412
rect 14439 31372 14445 31412
rect 14399 31344 14445 31372
rect 14399 31300 14405 31344
rect 14439 31300 14445 31344
rect 14399 31276 14445 31300
rect 14399 31228 14405 31276
rect 14439 31228 14445 31276
rect 14399 31208 14445 31228
rect 14399 31156 14405 31208
rect 14439 31156 14445 31208
rect 14399 31140 14445 31156
rect 14399 31084 14405 31140
rect 14439 31084 14445 31140
rect 14399 31072 14445 31084
rect 14399 31012 14405 31072
rect 14439 31012 14445 31072
rect 14399 31004 14445 31012
rect 14399 30940 14405 31004
rect 14439 30940 14445 31004
rect 14399 30936 14445 30940
rect 14399 30834 14405 30936
rect 14439 30834 14445 30936
rect 14399 30830 14445 30834
rect 14399 30766 14405 30830
rect 14439 30766 14445 30830
rect 14399 30758 14445 30766
rect 14399 30698 14405 30758
rect 14439 30698 14445 30758
rect 14399 30686 14445 30698
rect 14399 30630 14405 30686
rect 14439 30630 14445 30686
rect 14399 30614 14445 30630
rect 14399 30562 14405 30614
rect 14439 30562 14445 30614
rect 14399 30542 14445 30562
rect 14399 30494 14405 30542
rect 14439 30494 14445 30542
rect 14399 30470 14445 30494
rect 14399 30426 14405 30470
rect 14439 30426 14445 30470
rect 14399 30398 14445 30426
rect 14399 30358 14405 30398
rect 14439 30358 14445 30398
rect 14399 30326 14445 30358
rect 14399 30290 14405 30326
rect 14439 30290 14445 30326
rect 14399 30256 14445 30290
rect 14399 30220 14405 30256
rect 14439 30220 14445 30256
rect 14399 30188 14445 30220
rect 14399 30148 14405 30188
rect 14439 30148 14445 30188
rect 14399 30120 14445 30148
rect 14399 30076 14405 30120
rect 14439 30076 14445 30120
rect 14399 30052 14445 30076
rect 14399 30004 14405 30052
rect 14439 30004 14445 30052
rect 14399 29984 14445 30004
rect 14399 29932 14405 29984
rect 14439 29932 14445 29984
rect 14399 29916 14445 29932
rect 14399 29860 14405 29916
rect 14439 29860 14445 29916
rect 14399 29848 14445 29860
rect 14399 29788 14405 29848
rect 14439 29788 14445 29848
rect 14399 29780 14445 29788
rect 14399 29716 14405 29780
rect 14439 29716 14445 29780
rect 14399 29712 14445 29716
rect 14399 29610 14405 29712
rect 14439 29610 14445 29712
rect 14399 29606 14445 29610
rect 14399 29542 14405 29606
rect 14439 29542 14445 29606
rect 14399 29534 14445 29542
rect 14399 29474 14405 29534
rect 14439 29474 14445 29534
rect 14399 29462 14445 29474
rect 14399 29406 14405 29462
rect 14439 29406 14445 29462
rect 14399 29390 14445 29406
rect 14399 29338 14405 29390
rect 14439 29338 14445 29390
rect 14399 29318 14445 29338
rect 14399 29270 14405 29318
rect 14439 29270 14445 29318
rect 14399 29246 14445 29270
rect 14399 29202 14405 29246
rect 14439 29202 14445 29246
rect 14399 29174 14445 29202
rect 14399 29134 14405 29174
rect 14439 29134 14445 29174
rect 14399 29102 14445 29134
rect 14399 29066 14405 29102
rect 14439 29066 14445 29102
rect 14399 29032 14445 29066
rect 14399 28996 14405 29032
rect 14439 28996 14445 29032
rect 14399 28964 14445 28996
rect 14399 28924 14405 28964
rect 14439 28924 14445 28964
rect 14399 28896 14445 28924
rect 14399 28852 14405 28896
rect 14439 28852 14445 28896
rect 14399 28828 14445 28852
rect 14399 28780 14405 28828
rect 14439 28780 14445 28828
rect 14399 28760 14445 28780
rect 14399 28708 14405 28760
rect 14439 28708 14445 28760
rect 14399 28692 14445 28708
rect 14399 28636 14405 28692
rect 14439 28636 14445 28692
rect 14399 28624 14445 28636
rect 14399 28564 14405 28624
rect 14439 28564 14445 28624
rect 14399 28556 14445 28564
rect 14399 28492 14405 28556
rect 14439 28492 14445 28556
rect 14399 28488 14445 28492
rect 14399 28386 14405 28488
rect 14439 28386 14445 28488
rect 14399 28382 14445 28386
rect 14399 28318 14405 28382
rect 14439 28318 14445 28382
rect 14399 28310 14445 28318
rect 14399 28250 14405 28310
rect 14439 28250 14445 28310
rect 14399 28238 14445 28250
rect 14399 28182 14405 28238
rect 14439 28182 14445 28238
rect 14399 28166 14445 28182
rect 14399 28114 14405 28166
rect 14439 28114 14445 28166
rect 14399 28094 14445 28114
rect 14399 28046 14405 28094
rect 14439 28046 14445 28094
rect 14399 28022 14445 28046
rect 14399 27978 14405 28022
rect 14439 27978 14445 28022
rect 14399 27950 14445 27978
rect 14399 27910 14405 27950
rect 14439 27910 14445 27950
rect 14399 27878 14445 27910
rect 14399 27842 14405 27878
rect 14439 27842 14445 27878
rect 14399 27808 14445 27842
rect 14399 27772 14405 27808
rect 14439 27772 14445 27808
rect 9789 27682 9823 27716
rect 9789 27614 9823 27648
rect 9789 27546 9823 27580
rect 9783 27512 9789 27542
rect 14399 27740 14445 27772
rect 14399 27700 14405 27740
rect 14439 27700 14445 27740
rect 14399 27672 14445 27700
rect 14399 27628 14405 27672
rect 14439 27628 14445 27672
rect 14399 27604 14445 27628
rect 14399 27570 14405 27604
rect 14439 27570 14445 27604
rect 14399 27542 14445 27570
rect 9823 27512 9829 27542
rect 12426 27536 14445 27542
rect 12426 27530 12500 27536
rect 9783 27490 9829 27512
rect 9783 27444 9789 27490
rect 9823 27444 9829 27490
rect 11994 27482 12059 27516
rect 12093 27482 12157 27516
rect 12426 27496 12432 27530
rect 12466 27502 12500 27530
rect 12544 27502 12568 27536
rect 12616 27502 12636 27536
rect 12688 27502 12704 27536
rect 12760 27502 12772 27536
rect 12832 27502 12840 27536
rect 12904 27502 12908 27536
rect 13010 27502 13014 27536
rect 13078 27502 13086 27536
rect 13146 27502 13158 27536
rect 13214 27502 13230 27536
rect 13282 27502 13302 27536
rect 13350 27502 13374 27536
rect 13418 27502 13446 27536
rect 13486 27502 13518 27536
rect 13554 27502 13588 27536
rect 13624 27502 13656 27536
rect 13696 27502 13724 27536
rect 13768 27502 13792 27536
rect 13840 27502 13860 27536
rect 13912 27502 13928 27536
rect 13984 27502 13996 27536
rect 14056 27502 14064 27536
rect 14128 27502 14132 27536
rect 14166 27502 14183 27536
rect 14234 27502 14255 27536
rect 14302 27502 14327 27536
rect 14370 27502 14399 27536
rect 14433 27502 14445 27536
rect 12466 27496 14445 27502
rect 9783 27418 9829 27444
rect 9783 27376 9789 27418
rect 9823 27376 9829 27418
rect 9783 27346 9829 27376
rect 9783 27308 9789 27346
rect 9823 27308 9829 27346
rect 9783 27274 9829 27308
rect 9783 27240 9789 27274
rect 9823 27240 9829 27274
rect 9783 27206 9829 27240
rect 9783 27168 9789 27206
rect 9823 27168 9829 27206
rect 9783 27138 9829 27168
rect 9783 27096 9789 27138
rect 9823 27096 9829 27138
rect 9783 27070 9829 27096
rect 9783 27024 9789 27070
rect 9823 27024 9829 27070
rect 9783 27002 9829 27024
rect 9783 26952 9789 27002
rect 9823 26952 9829 27002
rect 9783 26934 9829 26952
rect 9783 26880 9789 26934
rect 9823 26880 9829 26934
rect 9783 26866 9829 26880
rect 9783 26808 9789 26866
rect 9823 26808 9829 26866
rect 9783 26798 9829 26808
rect 9783 26736 9789 26798
rect 9823 26736 9829 26798
rect 9783 26730 9829 26736
rect 9783 26664 9789 26730
rect 9823 26664 9829 26730
rect 10105 27455 10139 27471
rect 10105 27382 10139 27421
rect 10105 27309 10139 27348
rect 10105 27236 10139 27275
rect 10105 27163 10139 27202
rect 10105 27090 10139 27124
rect 10105 27017 10139 27052
rect 10105 26943 10139 26983
rect 10105 26869 10139 26909
rect 10105 26795 10139 26835
rect 10105 26721 10139 26761
rect 10105 26671 10139 26687
rect 12426 27458 12472 27496
rect 12426 27390 12432 27458
rect 12466 27390 12472 27458
rect 12426 27386 12472 27390
rect 12426 27322 12432 27386
rect 12466 27322 12472 27386
rect 12426 27314 12472 27322
rect 12426 27254 12432 27314
rect 12466 27254 12472 27314
rect 12426 27242 12472 27254
rect 12426 27186 12432 27242
rect 12466 27186 12472 27242
rect 12426 27170 12472 27186
rect 12426 27118 12432 27170
rect 12466 27118 12472 27170
rect 12426 27098 12472 27118
rect 12426 27050 12432 27098
rect 12466 27050 12472 27098
rect 12426 27026 12472 27050
rect 12426 26982 12432 27026
rect 12466 26982 12472 27026
rect 12426 26954 12472 26982
rect 12426 26914 12432 26954
rect 12466 26914 12472 26954
rect 12426 26882 12472 26914
rect 12426 26846 12432 26882
rect 12466 26846 12472 26882
rect 12426 26812 12472 26846
rect 12426 26776 12432 26812
rect 12466 26776 12472 26812
rect 12426 26744 12472 26776
rect 12426 26704 12432 26744
rect 12466 26704 12472 26744
rect 12426 26676 12472 26704
rect 9783 26662 9829 26664
rect 9783 26628 9789 26662
rect 9823 26628 9829 26662
rect 9783 26626 9829 26628
rect 11994 26626 12059 26660
rect 12093 26626 12157 26660
rect 12426 26632 12432 26676
rect 12466 26632 12472 26676
rect 9783 26560 9789 26626
rect 9823 26560 9829 26626
rect 9783 26554 9829 26560
rect 9783 26492 9789 26554
rect 9823 26492 9829 26554
rect 9783 26482 9829 26492
rect 9783 26448 9789 26482
rect 9823 26448 9829 26482
rect 9783 26410 9829 26448
rect 12426 26608 12472 26632
rect 12426 26560 12432 26608
rect 12466 26560 12472 26608
rect 12426 26540 12472 26560
rect 12426 26488 12432 26540
rect 12466 26488 12472 26540
rect 12426 26472 12472 26488
rect 12426 26438 12432 26472
rect 12466 26438 12472 26472
rect 12426 26410 12472 26438
rect 9783 26376 9789 26410
rect 9823 26404 12472 26410
rect 9823 26376 9857 26404
rect 9783 26370 9857 26376
rect 9891 26370 9906 26404
rect 9959 26370 9978 26404
rect 10027 26370 10050 26404
rect 10095 26370 10122 26404
rect 10163 26370 10194 26404
rect 10231 26370 10265 26404
rect 10300 26370 10333 26404
rect 10372 26370 10401 26404
rect 10444 26370 10469 26404
rect 10516 26370 10537 26404
rect 10588 26370 10605 26404
rect 10660 26370 10673 26404
rect 10732 26370 10741 26404
rect 10804 26370 10809 26404
rect 10876 26370 10877 26404
rect 10911 26370 10914 26404
rect 10979 26370 10986 26404
rect 11047 26370 11058 26404
rect 11115 26370 11130 26404
rect 11183 26370 11202 26404
rect 11251 26370 11274 26404
rect 11319 26370 11346 26404
rect 11387 26370 11418 26404
rect 11455 26370 11489 26404
rect 11524 26370 11557 26404
rect 11596 26370 11625 26404
rect 11668 26370 11693 26404
rect 11740 26370 11761 26404
rect 11812 26370 11829 26404
rect 11884 26370 11897 26404
rect 11956 26370 11965 26404
rect 12028 26370 12033 26404
rect 12100 26370 12101 26404
rect 12135 26370 12138 26404
rect 12203 26370 12210 26404
rect 12271 26370 12282 26404
rect 12339 26370 12354 26404
rect 12388 26370 12426 26404
rect 12460 26370 12472 26404
rect 9783 26364 12472 26370
rect 130 17343 2270 17344
rect 130 17309 176 17343
rect 210 17309 244 17343
rect 278 17309 312 17343
rect 346 17309 380 17343
rect 414 17309 448 17343
rect 482 17309 516 17343
rect 550 17309 584 17343
rect 618 17309 652 17343
rect 686 17309 720 17343
rect 754 17309 788 17343
rect 822 17309 856 17343
rect 890 17309 924 17343
rect 958 17309 992 17343
rect 1026 17309 1060 17343
rect 1094 17309 1128 17343
rect 1162 17309 1196 17343
rect 1230 17309 1264 17343
rect 1298 17309 1332 17343
rect 1366 17309 1400 17343
rect 1434 17309 1468 17343
rect 1502 17309 1536 17343
rect 1570 17309 1604 17343
rect 1638 17309 1672 17343
rect 1706 17309 1740 17343
rect 1774 17309 1808 17343
rect 1842 17309 1876 17343
rect 1910 17309 1944 17343
rect 1978 17309 2012 17343
rect 2046 17309 2080 17343
rect 2114 17309 2148 17343
rect 2182 17309 2270 17343
rect 130 17308 2270 17309
rect 130 17189 166 17308
rect 2234 17249 2270 17308
rect 2234 17215 2235 17249
rect 2269 17215 2270 17249
rect 164 17155 166 17189
rect 130 17117 166 17155
rect 164 17083 166 17117
rect 130 17045 166 17083
rect 164 17011 166 17045
rect 130 16973 166 17011
rect 246 17161 284 17195
rect 212 16989 318 17161
rect 522 17161 560 17195
rect 488 16989 594 17161
rect 628 16989 716 17191
rect 870 17161 908 17195
rect 836 16989 942 17161
rect 2234 17181 2270 17215
rect 2234 17147 2235 17181
rect 2269 17147 2270 17181
rect 2234 17113 2270 17147
rect 2234 17079 2235 17113
rect 2269 17079 2270 17113
rect 2234 17045 2270 17079
rect 2234 17011 2235 17045
rect 2269 17011 2270 17045
rect 164 16939 166 16973
rect 130 16909 166 16939
rect 130 16908 370 16909
rect 130 16874 234 16908
rect 295 16874 302 16908
rect 367 16874 370 16908
rect 130 16873 370 16874
rect 404 16906 438 16989
rect 628 16906 662 16989
rect 2234 16977 2270 17011
rect 2234 16943 2235 16977
rect 2269 16943 2270 16977
rect 2234 16909 2270 16943
rect 130 12149 166 16873
rect 404 16872 662 16906
rect 698 16908 4906 16909
rect 698 16874 714 16908
rect 748 16874 836 16908
rect 870 16874 904 16908
rect 938 16874 972 16908
rect 1006 16874 1040 16908
rect 1074 16874 1108 16908
rect 1142 16874 1176 16908
rect 1210 16874 1244 16908
rect 1278 16874 1312 16908
rect 1346 16874 1380 16908
rect 1414 16874 1448 16908
rect 1482 16874 1516 16908
rect 1550 16874 1584 16908
rect 1618 16874 1652 16908
rect 1686 16874 1720 16908
rect 1754 16874 1788 16908
rect 1822 16874 1856 16908
rect 1890 16874 1924 16908
rect 1958 16874 1992 16908
rect 2026 16874 2060 16908
rect 2094 16874 2128 16908
rect 2162 16874 2196 16908
rect 2230 16874 2264 16908
rect 2298 16874 2332 16908
rect 2366 16874 2400 16908
rect 2434 16874 2468 16908
rect 2502 16874 2570 16908
rect 2604 16874 2638 16908
rect 2672 16874 2706 16908
rect 2740 16874 2774 16908
rect 2808 16874 2842 16908
rect 2876 16874 2910 16908
rect 2944 16874 2978 16908
rect 3012 16874 3046 16908
rect 3080 16874 3114 16908
rect 3148 16874 3182 16908
rect 3216 16874 3250 16908
rect 3284 16874 3318 16908
rect 3352 16874 3386 16908
rect 3420 16874 3454 16908
rect 3488 16874 3522 16908
rect 3556 16874 3590 16908
rect 3624 16874 3658 16908
rect 3692 16874 3726 16908
rect 3760 16874 3794 16908
rect 3828 16874 3862 16908
rect 3896 16874 3930 16908
rect 3964 16874 3998 16908
rect 4032 16874 4066 16908
rect 4100 16874 4134 16908
rect 4168 16874 4202 16908
rect 4236 16874 4270 16908
rect 4304 16874 4338 16908
rect 4372 16874 4406 16908
rect 4440 16874 4474 16908
rect 4508 16874 4542 16908
rect 4576 16874 4610 16908
rect 4644 16874 4678 16908
rect 4712 16874 4746 16908
rect 4780 16875 4906 16908
rect 4780 16874 4871 16875
rect 698 16873 4871 16874
rect 404 16835 438 16872
rect 236 16789 252 16823
rect 286 16789 320 16823
rect 354 16789 370 16823
rect 248 16695 282 16789
rect 404 16763 438 16801
rect 480 16789 496 16823
rect 530 16789 564 16823
rect 598 16789 632 16823
rect 666 16789 700 16823
rect 734 16789 768 16823
rect 802 16789 818 16823
rect 480 16778 818 16789
rect 480 16744 560 16778
rect 594 16744 632 16778
rect 666 16744 704 16778
rect 738 16744 776 16778
rect 810 16744 818 16778
rect 936 16789 952 16823
rect 986 16789 1020 16823
rect 1054 16789 1088 16823
rect 1122 16789 1156 16823
rect 1190 16789 1224 16823
rect 1258 16789 1274 16823
rect 936 16778 1274 16789
rect 936 16744 944 16778
rect 978 16744 1016 16778
rect 1050 16744 1088 16778
rect 1122 16744 1160 16778
rect 1194 16744 1274 16778
rect 1392 16789 1408 16823
rect 1442 16789 1476 16823
rect 1510 16789 1544 16823
rect 1578 16789 1612 16823
rect 1646 16789 1680 16823
rect 1714 16789 1730 16823
rect 1392 16778 1730 16789
rect 1392 16744 1472 16778
rect 1506 16744 1544 16778
rect 1578 16744 1616 16778
rect 1650 16744 1688 16778
rect 1722 16744 1730 16778
rect 1848 16789 1864 16823
rect 1898 16789 1932 16823
rect 1966 16789 2000 16823
rect 2034 16789 2068 16823
rect 2102 16789 2136 16823
rect 2170 16789 2186 16823
rect 2273 16789 2289 16823
rect 2323 16789 2357 16823
rect 2391 16789 2418 16823
rect 1848 16778 2186 16789
rect 1848 16744 1856 16778
rect 1890 16744 1928 16778
rect 1962 16744 2000 16778
rect 2034 16744 2072 16778
rect 2106 16744 2186 16778
rect 2384 16695 2418 16789
rect 2465 16805 2571 16873
rect 4870 16841 4871 16873
rect 4905 16841 4906 16875
rect 2465 16771 2501 16805
rect 2535 16771 2571 16805
rect 2465 16737 2571 16771
rect 2465 16703 2501 16737
rect 2535 16703 2571 16737
rect 2465 16669 2571 16703
rect 2618 16789 2645 16823
rect 2679 16789 2713 16823
rect 2747 16789 2763 16823
rect 2850 16789 2866 16823
rect 2900 16789 2934 16823
rect 2968 16789 3002 16823
rect 3036 16789 3070 16823
rect 3104 16789 3138 16823
rect 3172 16789 3188 16823
rect 2618 16695 2652 16789
rect 2850 16778 3188 16789
rect 2850 16744 2930 16778
rect 2964 16744 3002 16778
rect 3036 16744 3074 16778
rect 3108 16744 3146 16778
rect 3180 16744 3188 16778
rect 3306 16789 3322 16823
rect 3356 16789 3390 16823
rect 3424 16789 3458 16823
rect 3492 16789 3526 16823
rect 3560 16789 3594 16823
rect 3628 16789 3644 16823
rect 3306 16778 3644 16789
rect 3306 16744 3314 16778
rect 3348 16744 3386 16778
rect 3420 16744 3458 16778
rect 3492 16744 3530 16778
rect 3564 16744 3644 16778
rect 3762 16789 3778 16823
rect 3812 16789 3846 16823
rect 3880 16789 3914 16823
rect 3948 16789 3982 16823
rect 4016 16789 4050 16823
rect 4084 16789 4100 16823
rect 3762 16778 4100 16789
rect 3762 16744 3842 16778
rect 3876 16744 3914 16778
rect 3948 16744 3986 16778
rect 4020 16744 4058 16778
rect 4092 16744 4100 16778
rect 4218 16789 4234 16823
rect 4268 16789 4302 16823
rect 4336 16789 4370 16823
rect 4404 16789 4438 16823
rect 4472 16789 4506 16823
rect 4540 16789 4556 16823
rect 4643 16789 4659 16823
rect 4693 16789 4727 16823
rect 4761 16789 4788 16823
rect 4218 16778 4556 16789
rect 4218 16744 4226 16778
rect 4260 16744 4298 16778
rect 4332 16744 4370 16778
rect 4404 16744 4442 16778
rect 4476 16744 4556 16778
rect 4754 16695 4788 16789
rect 4870 16807 4906 16841
rect 4870 16773 4871 16807
rect 4905 16773 4906 16807
rect 4870 16739 4906 16773
rect 4870 16705 4871 16739
rect 4905 16705 4906 16739
rect 2465 16635 2501 16669
rect 2535 16635 2571 16669
rect 2465 16601 2571 16635
rect 2465 16567 2501 16601
rect 2535 16567 2571 16601
rect 2465 16533 2571 16567
rect 2465 16523 2501 16533
rect 2500 16499 2501 16523
rect 2535 16523 2571 16533
rect 4870 16671 4906 16705
rect 4870 16637 4871 16671
rect 4905 16637 4906 16671
rect 4870 16603 4906 16637
rect 4870 16569 4871 16603
rect 4905 16569 4906 16603
rect 4870 16535 4906 16569
rect 2535 16499 2536 16523
rect 2500 16465 2536 16499
rect 2500 16431 2501 16465
rect 2535 16431 2536 16465
rect 2500 16397 2536 16431
rect 2500 16363 2501 16397
rect 2535 16363 2536 16397
rect 2500 16329 2536 16363
rect 2500 16295 2501 16329
rect 2535 16295 2536 16329
rect 2500 16261 2536 16295
rect 2500 16227 2501 16261
rect 2535 16227 2536 16261
rect 2500 16193 2536 16227
rect 2500 16159 2501 16193
rect 2535 16159 2536 16193
rect 2500 16125 2536 16159
rect 2500 16091 2501 16125
rect 2535 16091 2536 16125
rect 2500 16057 2536 16091
rect 2500 16023 2501 16057
rect 2535 16023 2536 16057
rect 2500 15989 2536 16023
rect 2500 15955 2501 15989
rect 2535 15955 2536 15989
rect 2500 15921 2536 15955
rect 2500 15887 2501 15921
rect 2535 15887 2536 15921
rect 2500 15853 2536 15887
rect 2500 15819 2501 15853
rect 2535 15819 2536 15853
rect 2500 15785 2536 15819
rect 2500 15751 2501 15785
rect 2535 15751 2536 15785
rect 2500 15717 2536 15751
rect 2500 15683 2501 15717
rect 2535 15683 2536 15717
rect 2500 15649 2536 15683
rect 2500 15615 2501 15649
rect 2535 15615 2536 15649
rect 2500 15581 2536 15615
rect 2500 15547 2501 15581
rect 2535 15547 2536 15581
rect 2500 15513 2536 15547
rect 2500 15479 2501 15513
rect 2535 15479 2536 15513
rect 2500 15445 2536 15479
rect 2500 15411 2501 15445
rect 2535 15411 2536 15445
rect 2500 15377 2536 15411
rect 2500 15343 2501 15377
rect 2535 15343 2536 15377
rect 248 15293 282 15337
rect 2384 15293 2418 15337
rect 248 15259 275 15293
rect 309 15259 343 15293
rect 377 15259 393 15293
rect 2273 15259 2289 15293
rect 2323 15259 2357 15293
rect 2391 15259 2418 15293
rect 248 15209 282 15259
rect 2384 15209 2418 15259
rect 2500 15309 2536 15343
rect 4870 16501 4871 16535
rect 4905 16501 4906 16535
rect 4870 16467 4906 16501
rect 4870 16433 4871 16467
rect 4905 16433 4906 16467
rect 4870 16399 4906 16433
rect 4870 16365 4871 16399
rect 4905 16365 4906 16399
rect 4870 16331 4906 16365
rect 4870 16297 4871 16331
rect 4905 16297 4906 16331
rect 4870 16263 4906 16297
rect 4870 16229 4871 16263
rect 4905 16229 4906 16263
rect 4870 16195 4906 16229
rect 4870 16161 4871 16195
rect 4905 16161 4906 16195
rect 4870 16127 4906 16161
rect 4870 16093 4871 16127
rect 4905 16093 4906 16127
rect 4870 16059 4906 16093
rect 4870 16025 4871 16059
rect 4905 16025 4906 16059
rect 4870 15991 4906 16025
rect 4870 15957 4871 15991
rect 4905 15957 4906 15991
rect 4870 15923 4906 15957
rect 4870 15889 4871 15923
rect 4905 15889 4906 15923
rect 4870 15855 4906 15889
rect 4870 15821 4871 15855
rect 4905 15821 4906 15855
rect 4870 15787 4906 15821
rect 4870 15753 4871 15787
rect 4905 15753 4906 15787
rect 4870 15719 4906 15753
rect 4870 15685 4871 15719
rect 4905 15685 4906 15719
rect 4870 15651 4906 15685
rect 4870 15617 4871 15651
rect 4905 15617 4906 15651
rect 4870 15583 4906 15617
rect 4870 15549 4871 15583
rect 4905 15549 4906 15583
rect 4870 15515 4906 15549
rect 4870 15481 4871 15515
rect 4905 15481 4906 15515
rect 4870 15447 4906 15481
rect 4870 15413 4871 15447
rect 4905 15413 4906 15447
rect 4870 15379 4906 15413
rect 4870 15345 4871 15379
rect 4905 15345 4906 15379
rect 2500 15275 2501 15309
rect 2535 15275 2536 15309
rect 2500 15241 2536 15275
rect 2500 15207 2501 15241
rect 2535 15207 2536 15241
rect 2618 15293 2652 15337
rect 4754 15293 4788 15337
rect 2618 15259 2645 15293
rect 2679 15259 2713 15293
rect 2747 15259 2763 15293
rect 4643 15259 4659 15293
rect 4693 15259 4727 15293
rect 4761 15259 4788 15293
rect 2618 15209 2652 15259
rect 4754 15209 4788 15259
rect 4870 15311 4906 15345
rect 4870 15277 4871 15311
rect 4905 15277 4906 15311
rect 4870 15243 4906 15277
rect 4870 15209 4871 15243
rect 4905 15209 4906 15243
rect 2500 15173 2536 15207
rect 2500 15139 2501 15173
rect 2535 15139 2536 15173
rect 2500 15105 2536 15139
rect 2500 15071 2501 15105
rect 2535 15071 2536 15105
rect 2500 15037 2536 15071
rect 2500 15003 2501 15037
rect 2535 15003 2536 15037
rect 2500 14969 2536 15003
rect 2500 14935 2501 14969
rect 2535 14935 2536 14969
rect 2500 14901 2536 14935
rect 2500 14867 2501 14901
rect 2535 14867 2536 14901
rect 2500 14833 2536 14867
rect 2500 14799 2501 14833
rect 2535 14799 2536 14833
rect 2500 14765 2536 14799
rect 2500 14731 2501 14765
rect 2535 14731 2536 14765
rect 2500 14697 2536 14731
rect 2500 14663 2501 14697
rect 2535 14663 2536 14697
rect 2500 14629 2536 14663
rect 2500 14595 2501 14629
rect 2535 14595 2536 14629
rect 2500 14561 2536 14595
rect 2500 14527 2501 14561
rect 2535 14527 2536 14561
rect 2500 14493 2536 14527
rect 2500 14459 2501 14493
rect 2535 14459 2536 14493
rect 2500 14425 2536 14459
rect 2500 14391 2501 14425
rect 2535 14391 2536 14425
rect 2500 14357 2536 14391
rect 2500 14323 2501 14357
rect 2535 14323 2536 14357
rect 2500 14289 2536 14323
rect 2500 14255 2501 14289
rect 2535 14255 2536 14289
rect 2500 14221 2536 14255
rect 2500 14187 2501 14221
rect 2535 14187 2536 14221
rect 2500 14153 2536 14187
rect 2500 14119 2501 14153
rect 2535 14119 2536 14153
rect 2500 14085 2536 14119
rect 2500 14051 2501 14085
rect 2535 14051 2536 14085
rect 2500 14017 2536 14051
rect 2500 13983 2501 14017
rect 2535 13983 2536 14017
rect 2500 13949 2536 13983
rect 2500 13915 2501 13949
rect 2535 13915 2536 13949
rect 2500 13881 2536 13915
rect 2500 13847 2501 13881
rect 2535 13847 2536 13881
rect 2500 13813 2536 13847
rect 248 13763 282 13807
rect 2384 13763 2418 13807
rect 248 13729 275 13763
rect 309 13729 343 13763
rect 377 13729 393 13763
rect 480 13729 488 13763
rect 530 13729 560 13763
rect 598 13729 632 13763
rect 666 13729 700 13763
rect 738 13729 768 13763
rect 810 13729 818 13763
rect 936 13729 944 13763
rect 986 13729 1016 13763
rect 1054 13729 1088 13763
rect 1122 13729 1156 13763
rect 1194 13729 1224 13763
rect 1266 13729 1274 13763
rect 1392 13729 1400 13763
rect 1442 13729 1472 13763
rect 1510 13729 1544 13763
rect 1578 13729 1612 13763
rect 1650 13729 1680 13763
rect 1722 13729 1730 13763
rect 1848 13729 1856 13763
rect 1898 13729 1928 13763
rect 1966 13729 2000 13763
rect 2034 13729 2068 13763
rect 2106 13729 2136 13763
rect 2178 13729 2186 13763
rect 2273 13729 2289 13763
rect 2323 13729 2357 13763
rect 2391 13729 2418 13763
rect 248 13679 282 13729
rect 2384 13679 2418 13729
rect 2500 13779 2501 13813
rect 2535 13779 2536 13813
rect 4870 15175 4906 15209
rect 4870 15141 4871 15175
rect 4905 15141 4906 15175
rect 4870 15107 4906 15141
rect 4870 15073 4871 15107
rect 4905 15073 4906 15107
rect 4870 15039 4906 15073
rect 4870 15005 4871 15039
rect 4905 15005 4906 15039
rect 4870 14971 4906 15005
rect 4870 14937 4871 14971
rect 4905 14937 4906 14971
rect 4870 14903 4906 14937
rect 4870 14869 4871 14903
rect 4905 14869 4906 14903
rect 4870 14835 4906 14869
rect 4870 14801 4871 14835
rect 4905 14801 4906 14835
rect 4870 14767 4906 14801
rect 4870 14733 4871 14767
rect 4905 14733 4906 14767
rect 4870 14699 4906 14733
rect 4870 14665 4871 14699
rect 4905 14665 4906 14699
rect 4870 14631 4906 14665
rect 4870 14597 4871 14631
rect 4905 14597 4906 14631
rect 4870 14563 4906 14597
rect 4870 14529 4871 14563
rect 4905 14529 4906 14563
rect 4870 14495 4906 14529
rect 4870 14461 4871 14495
rect 4905 14461 4906 14495
rect 4870 14427 4906 14461
rect 4870 14393 4871 14427
rect 4905 14393 4906 14427
rect 4870 14359 4906 14393
rect 4870 14325 4871 14359
rect 4905 14325 4906 14359
rect 4870 14291 4906 14325
rect 4870 14257 4871 14291
rect 4905 14257 4906 14291
rect 4870 14223 4906 14257
rect 4870 14189 4871 14223
rect 4905 14189 4906 14223
rect 4870 14155 4906 14189
rect 4870 14121 4871 14155
rect 4905 14121 4906 14155
rect 4870 14087 4906 14121
rect 4870 14053 4871 14087
rect 4905 14053 4906 14087
rect 4870 14019 4906 14053
rect 4870 13985 4871 14019
rect 4905 13985 4906 14019
rect 4870 13951 4906 13985
rect 4870 13917 4871 13951
rect 4905 13917 4906 13951
rect 4870 13883 4906 13917
rect 4870 13849 4871 13883
rect 4905 13849 4906 13883
rect 4870 13815 4906 13849
rect 2500 13745 2536 13779
rect 2500 13711 2501 13745
rect 2535 13711 2536 13745
rect 2500 13677 2536 13711
rect 2618 13763 2652 13807
rect 4754 13763 4788 13807
rect 2618 13729 2645 13763
rect 2679 13729 2713 13763
rect 2747 13729 2763 13763
rect 2850 13729 2858 13763
rect 2900 13729 2930 13763
rect 2968 13729 3002 13763
rect 3036 13729 3070 13763
rect 3108 13729 3138 13763
rect 3180 13729 3188 13763
rect 3306 13729 3314 13763
rect 3356 13729 3386 13763
rect 3424 13729 3458 13763
rect 3492 13729 3526 13763
rect 3564 13729 3594 13763
rect 3636 13729 3644 13763
rect 3762 13729 3770 13763
rect 3812 13729 3842 13763
rect 3880 13729 3914 13763
rect 3948 13729 3982 13763
rect 4020 13729 4050 13763
rect 4092 13729 4100 13763
rect 4218 13729 4226 13763
rect 4268 13729 4298 13763
rect 4336 13729 4370 13763
rect 4404 13729 4438 13763
rect 4476 13729 4506 13763
rect 4548 13729 4556 13763
rect 4643 13729 4659 13763
rect 4693 13729 4727 13763
rect 4761 13729 4788 13763
rect 2618 13679 2652 13729
rect 4754 13679 4788 13729
rect 4870 13781 4871 13815
rect 4905 13781 4906 13815
rect 4870 13747 4906 13781
rect 4870 13713 4871 13747
rect 4905 13713 4906 13747
rect 4870 13679 4906 13713
rect 2500 13643 2501 13677
rect 2535 13643 2536 13677
rect 2500 13609 2536 13643
rect 2500 13575 2501 13609
rect 2535 13575 2536 13609
rect 2500 13541 2536 13575
rect 2500 13507 2501 13541
rect 2535 13507 2536 13541
rect 2500 13473 2536 13507
rect 2500 13439 2501 13473
rect 2535 13439 2536 13473
rect 2500 13405 2536 13439
rect 2500 13371 2501 13405
rect 2535 13371 2536 13405
rect 2500 13337 2536 13371
rect 2500 13303 2501 13337
rect 2535 13303 2536 13337
rect 2500 13269 2536 13303
rect 2500 13235 2501 13269
rect 2535 13235 2536 13269
rect 2500 13201 2536 13235
rect 2500 13167 2501 13201
rect 2535 13167 2536 13201
rect 2500 13133 2536 13167
rect 2500 13099 2501 13133
rect 2535 13099 2536 13133
rect 2500 13065 2536 13099
rect 2500 13031 2501 13065
rect 2535 13031 2536 13065
rect 2500 12997 2536 13031
rect 2500 12963 2501 12997
rect 2535 12963 2536 12997
rect 2500 12929 2536 12963
rect 2500 12895 2501 12929
rect 2535 12895 2536 12929
rect 2500 12861 2536 12895
rect 2500 12827 2501 12861
rect 2535 12827 2536 12861
rect 2500 12793 2536 12827
rect 2500 12759 2501 12793
rect 2535 12759 2536 12793
rect 2500 12725 2536 12759
rect 2500 12691 2501 12725
rect 2535 12691 2536 12725
rect 2500 12657 2536 12691
rect 2500 12623 2501 12657
rect 2535 12623 2536 12657
rect 2500 12589 2536 12623
rect 2500 12555 2501 12589
rect 2535 12555 2536 12589
rect 2500 12521 2536 12555
rect 2500 12487 2501 12521
rect 2535 12487 2536 12521
rect 2500 12453 2536 12487
rect 2500 12419 2501 12453
rect 2535 12419 2536 12453
rect 2500 12385 2536 12419
rect 2500 12351 2501 12385
rect 2535 12351 2536 12385
rect 2500 12317 2536 12351
rect 3230 13584 3264 13625
rect 3230 13508 3264 13550
rect 3230 13432 3264 13474
rect 3230 13356 3264 13398
rect 3230 13280 3264 13322
rect 3230 13204 3264 13246
rect 3230 13128 3264 13170
rect 3230 13052 3264 13094
rect 3230 12976 3264 13018
rect 3230 12900 3264 12942
rect 3230 12824 3264 12866
rect 3230 12748 3264 12790
rect 3230 12672 3264 12714
rect 3230 12596 3264 12638
rect 3230 12520 3264 12562
rect 3230 12444 3264 12486
rect 3230 12368 3264 12410
rect 4870 13645 4871 13679
rect 4905 13645 4906 13679
rect 4870 13611 4906 13645
rect 4870 13577 4871 13611
rect 4905 13577 4906 13611
rect 4870 13543 4906 13577
rect 4870 13509 4871 13543
rect 4905 13509 4906 13543
rect 4870 13475 4906 13509
rect 4870 13441 4871 13475
rect 4905 13441 4906 13475
rect 4870 13407 4906 13441
rect 4870 13373 4871 13407
rect 4905 13373 4906 13407
rect 4870 13339 4906 13373
rect 4870 13305 4871 13339
rect 4905 13305 4906 13339
rect 4870 13271 4906 13305
rect 4870 13237 4871 13271
rect 4905 13237 4906 13271
rect 4870 13203 4906 13237
rect 4870 13169 4871 13203
rect 4905 13169 4906 13203
rect 4870 13135 4906 13169
rect 4870 13101 4871 13135
rect 4905 13101 4906 13135
rect 4870 13067 4906 13101
rect 4870 13033 4871 13067
rect 4905 13033 4906 13067
rect 4870 12999 4906 13033
rect 4870 12965 4871 12999
rect 4905 12965 4906 12999
rect 4870 12931 4906 12965
rect 4870 12897 4871 12931
rect 4905 12897 4906 12931
rect 4870 12863 4906 12897
rect 4870 12829 4871 12863
rect 4905 12829 4906 12863
rect 4870 12795 4906 12829
rect 4870 12761 4871 12795
rect 4905 12761 4906 12795
rect 4870 12727 4906 12761
rect 4870 12693 4871 12727
rect 4905 12693 4906 12727
rect 4870 12659 4906 12693
rect 4870 12625 4871 12659
rect 4905 12625 4906 12659
rect 4870 12591 4906 12625
rect 4870 12557 4871 12591
rect 4905 12557 4906 12591
rect 4870 12523 4906 12557
rect 4870 12489 4871 12523
rect 4905 12489 4906 12523
rect 4870 12455 4906 12489
rect 4870 12421 4871 12455
rect 4905 12421 4906 12455
rect 4870 12387 4906 12421
rect 4870 12353 4871 12387
rect 4905 12353 4906 12387
rect 2500 12283 2501 12317
rect 2535 12283 2536 12317
rect 248 12233 282 12277
rect 2384 12233 2418 12277
rect 2500 12249 2536 12283
rect 4870 12319 4906 12353
rect 4870 12285 4871 12319
rect 4905 12285 4906 12319
rect 2500 12245 2501 12249
rect 248 12199 275 12233
rect 309 12199 343 12233
rect 377 12199 393 12233
rect 480 12199 488 12233
rect 530 12199 560 12233
rect 598 12199 632 12233
rect 666 12199 700 12233
rect 738 12199 768 12233
rect 810 12199 818 12233
rect 936 12199 944 12233
rect 986 12199 1016 12233
rect 1054 12199 1088 12233
rect 1122 12199 1156 12233
rect 1194 12199 1224 12233
rect 1266 12199 1274 12233
rect 1392 12199 1400 12233
rect 1442 12199 1472 12233
rect 1510 12199 1544 12233
rect 1578 12199 1612 12233
rect 1650 12199 1680 12233
rect 1722 12199 1730 12233
rect 1848 12199 1856 12233
rect 1898 12199 1928 12233
rect 1966 12199 2000 12233
rect 2034 12199 2068 12233
rect 2106 12199 2136 12233
rect 2178 12199 2186 12233
rect 2273 12199 2289 12233
rect 2323 12199 2357 12233
rect 2391 12199 2418 12233
rect 2465 12215 2501 12245
rect 2535 12245 2536 12249
rect 2535 12215 2571 12245
rect 2465 12181 2571 12215
rect 2618 12233 2652 12277
rect 4754 12233 4788 12277
rect 2618 12199 2645 12233
rect 2679 12199 2713 12233
rect 2747 12199 2763 12233
rect 2850 12199 2858 12233
rect 2900 12199 2930 12233
rect 2968 12199 3002 12233
rect 3036 12199 3070 12233
rect 3108 12199 3138 12233
rect 3180 12199 3188 12233
rect 3306 12199 3314 12233
rect 3356 12199 3386 12233
rect 3424 12199 3458 12233
rect 3492 12199 3526 12233
rect 3564 12199 3594 12233
rect 3636 12199 3644 12233
rect 3762 12199 3770 12233
rect 3812 12199 3842 12233
rect 3880 12199 3914 12233
rect 3948 12199 3982 12233
rect 4020 12199 4050 12233
rect 4092 12199 4100 12233
rect 4218 12199 4226 12233
rect 4268 12199 4298 12233
rect 4336 12199 4370 12233
rect 4404 12199 4438 12233
rect 4476 12199 4506 12233
rect 4548 12199 4556 12233
rect 4643 12199 4659 12233
rect 4693 12199 4727 12233
rect 4761 12199 4788 12233
rect 2465 12149 2501 12181
rect 130 12148 2501 12149
rect 2535 12149 2571 12181
rect 4870 12182 4906 12285
rect 4870 12149 4871 12182
rect 2535 12148 4871 12149
rect 4905 12148 4906 12182
rect 130 12114 179 12148
rect 213 12114 251 12148
rect 285 12114 291 12148
rect 357 12114 359 12148
rect 393 12114 395 12148
rect 461 12114 467 12148
rect 529 12114 563 12148
rect 597 12114 631 12148
rect 665 12114 699 12148
rect 733 12114 767 12148
rect 801 12114 835 12148
rect 869 12114 903 12148
rect 937 12114 971 12148
rect 1005 12114 1039 12148
rect 1073 12114 1107 12148
rect 1141 12114 1175 12148
rect 1209 12114 1243 12148
rect 1277 12114 1311 12148
rect 1345 12114 1379 12148
rect 1413 12114 1447 12148
rect 1481 12114 1515 12148
rect 1549 12114 1583 12148
rect 1617 12114 1651 12148
rect 1685 12114 1719 12148
rect 1753 12114 1787 12148
rect 1821 12114 1855 12148
rect 1889 12114 1923 12148
rect 1957 12114 1991 12148
rect 2025 12114 2059 12148
rect 2093 12114 2127 12148
rect 2161 12114 2195 12148
rect 2229 12114 2263 12148
rect 2297 12114 2331 12148
rect 2365 12114 2399 12148
rect 2463 12114 2501 12148
rect 2535 12114 2573 12148
rect 2630 12114 2664 12148
rect 2698 12114 2732 12148
rect 2766 12114 2800 12148
rect 2834 12114 2868 12148
rect 2902 12114 2936 12148
rect 2970 12114 3004 12148
rect 3038 12114 3072 12148
rect 3106 12114 3140 12148
rect 3174 12114 3208 12148
rect 3242 12114 3276 12148
rect 3310 12114 3344 12148
rect 3378 12114 3412 12148
rect 3446 12114 3480 12148
rect 3514 12114 3548 12148
rect 3582 12114 3616 12148
rect 3650 12114 3684 12148
rect 3718 12114 3752 12148
rect 3786 12114 3820 12148
rect 3854 12114 3888 12148
rect 3922 12114 3956 12148
rect 3990 12114 4024 12148
rect 4058 12114 4092 12148
rect 4126 12114 4160 12148
rect 4194 12114 4228 12148
rect 4262 12114 4296 12148
rect 4330 12114 4364 12148
rect 4398 12114 4432 12148
rect 4466 12114 4500 12148
rect 4534 12114 4568 12148
rect 4602 12114 4636 12148
rect 4670 12114 4704 12148
rect 4738 12114 4772 12148
rect 4806 12114 4906 12148
rect 130 12113 4906 12114
rect 5059 15813 5684 15814
rect 5059 15780 5140 15813
rect 5059 15746 5060 15780
rect 5094 15779 5140 15780
rect 5174 15779 5208 15813
rect 5242 15779 5276 15813
rect 5310 15779 5344 15813
rect 5378 15779 5412 15813
rect 5446 15779 5480 15813
rect 5514 15779 5548 15813
rect 5582 15779 5616 15813
rect 5650 15779 5684 15813
rect 5094 15778 5684 15779
rect 5094 15746 5095 15778
rect 5059 15712 5095 15746
rect 5059 15678 5060 15712
rect 5094 15678 5095 15712
rect 5238 15698 5248 15732
rect 5282 15730 5320 15732
rect 5354 15730 5392 15732
rect 5426 15730 5464 15732
rect 5288 15698 5320 15730
rect 5238 15696 5254 15698
rect 5288 15696 5322 15698
rect 5356 15696 5390 15730
rect 5426 15698 5458 15730
rect 5498 15698 5508 15732
rect 5424 15696 5458 15698
rect 5492 15696 5508 15698
rect 5059 15644 5095 15678
rect 5059 15610 5060 15644
rect 5094 15610 5095 15644
rect 5059 15576 5095 15610
rect 5648 15686 5684 15778
rect 5648 15652 5649 15686
rect 5683 15652 5684 15686
rect 5648 15618 5684 15652
rect 5648 15584 5649 15618
rect 5683 15584 5684 15618
rect 5059 15542 5060 15576
rect 5094 15542 5095 15576
rect 5059 15508 5095 15542
rect 5059 15474 5060 15508
rect 5094 15474 5095 15508
rect 5059 15440 5095 15474
rect 5059 15406 5060 15440
rect 5094 15406 5095 15440
rect 5059 15372 5095 15406
rect 5059 15338 5060 15372
rect 5094 15338 5095 15372
rect 5059 15304 5095 15338
rect 5059 15270 5060 15304
rect 5094 15270 5095 15304
rect 5059 15236 5095 15270
rect 5059 15202 5060 15236
rect 5094 15202 5095 15236
rect 5059 15168 5095 15202
rect 5059 15134 5060 15168
rect 5094 15134 5095 15168
rect 5059 15100 5095 15134
rect 5180 15508 5214 15546
rect 5180 15436 5214 15474
rect 5180 15364 5214 15402
rect 5180 15292 5214 15330
rect 5180 15220 5214 15258
rect 5180 15148 5214 15186
rect 5356 15497 5390 15546
rect 5356 15414 5390 15463
rect 5356 15331 5390 15380
rect 5356 15248 5390 15297
rect 5356 15164 5390 15214
rect 5532 15508 5566 15546
rect 5532 15436 5566 15474
rect 5532 15364 5566 15402
rect 5532 15292 5566 15330
rect 5532 15220 5566 15258
rect 5532 15148 5566 15186
rect 5648 15550 5684 15584
rect 5648 15516 5649 15550
rect 5683 15516 5684 15550
rect 5648 15482 5684 15516
rect 5648 15448 5649 15482
rect 5683 15448 5684 15482
rect 5648 15414 5684 15448
rect 5648 15380 5649 15414
rect 5683 15380 5684 15414
rect 5648 15346 5684 15380
rect 5648 15312 5649 15346
rect 5683 15312 5684 15346
rect 5648 15278 5684 15312
rect 5648 15244 5649 15278
rect 5683 15244 5684 15278
rect 5648 15210 5684 15244
rect 5648 15176 5649 15210
rect 5683 15176 5684 15210
rect 5648 15142 5684 15176
rect 5059 15066 5060 15100
rect 5094 15066 5095 15100
rect 5059 14974 5095 15066
rect 5648 15108 5649 15142
rect 5683 15108 5684 15142
rect 5648 15074 5684 15108
rect 5648 15040 5649 15074
rect 5683 15040 5684 15074
rect 5648 15006 5684 15040
rect 5648 14974 5649 15006
rect 5059 14973 5649 14974
rect 5059 14939 5093 14973
rect 5127 14939 5161 14973
rect 5195 14939 5229 14973
rect 5263 14939 5297 14973
rect 5331 14939 5365 14973
rect 5399 14939 5433 14973
rect 5467 14939 5501 14973
rect 5535 14939 5569 14973
rect 5603 14972 5649 14973
rect 5683 14972 5684 15006
rect 5603 14939 5684 14972
rect 5059 14859 5684 14939
rect 5059 14858 6339 14859
rect 5059 14824 5093 14858
rect 5127 14824 5161 14858
rect 5195 14824 5229 14858
rect 5263 14824 5297 14858
rect 5331 14824 5365 14858
rect 5399 14824 5433 14858
rect 5467 14824 5501 14858
rect 5535 14824 5569 14858
rect 5603 14824 5637 14858
rect 5671 14824 5705 14858
rect 5739 14824 5773 14858
rect 5807 14824 5841 14858
rect 5875 14824 5909 14858
rect 5943 14824 5977 14858
rect 6011 14824 6045 14858
rect 6079 14824 6113 14858
rect 6147 14824 6181 14858
rect 6215 14825 6339 14858
rect 6215 14824 6304 14825
rect 5059 14823 6304 14824
rect 5059 14769 5095 14823
rect 5059 14735 5060 14769
rect 5094 14735 5095 14769
rect 6303 14791 6304 14823
rect 6338 14791 6339 14825
rect 6303 14757 6339 14791
rect 5059 14701 5095 14735
rect 5059 14667 5060 14701
rect 5094 14667 5095 14701
rect 5176 14707 5192 14741
rect 5226 14707 5242 14741
rect 5176 14673 5242 14707
rect 5596 14707 5612 14741
rect 5646 14707 5662 14741
rect 5059 14633 5095 14667
rect 5192 14671 5226 14673
rect 5596 14661 5662 14707
rect 5059 14599 5060 14633
rect 5094 14599 5095 14633
rect 5059 14565 5095 14599
rect 5059 14531 5060 14565
rect 5094 14531 5095 14565
rect 5596 14627 5612 14661
rect 5646 14627 5662 14661
rect 5596 14589 5662 14627
rect 5596 14555 5612 14589
rect 5646 14555 5662 14589
rect 5596 14549 5662 14555
rect 5736 14707 5752 14741
rect 5786 14707 5802 14741
rect 5736 14661 5802 14707
rect 5736 14627 5756 14661
rect 5790 14627 5802 14661
rect 5736 14589 5802 14627
rect 5736 14555 5756 14589
rect 5790 14555 5802 14589
rect 5736 14549 5802 14555
rect 5876 14707 5892 14741
rect 5926 14707 5942 14741
rect 5876 14661 5942 14707
rect 6016 14707 6032 14741
rect 6066 14707 6082 14741
rect 6016 14673 6082 14707
rect 5876 14627 5892 14661
rect 5926 14627 5942 14661
rect 5876 14589 5942 14627
rect 5876 14555 5892 14589
rect 5926 14555 5942 14589
rect 5876 14549 5942 14555
rect 6020 14661 6082 14673
rect 6020 14627 6036 14661
rect 6070 14627 6082 14661
rect 6020 14589 6082 14627
rect 6020 14555 6036 14589
rect 6070 14555 6082 14589
rect 6020 14549 6082 14555
rect 6156 14707 6172 14741
rect 6206 14707 6222 14741
rect 6156 14660 6222 14707
rect 6156 14626 6172 14660
rect 6206 14626 6222 14660
rect 6156 14588 6222 14626
rect 6156 14554 6172 14588
rect 6206 14554 6222 14588
rect 6156 14548 6222 14554
rect 6303 14723 6304 14757
rect 6338 14723 6339 14757
rect 6303 14689 6339 14723
rect 6303 14655 6304 14689
rect 6338 14655 6339 14689
rect 6303 14621 6339 14655
rect 6303 14587 6304 14621
rect 6338 14587 6339 14621
rect 6303 14553 6339 14587
rect 5059 14497 5095 14531
rect 5059 14463 5060 14497
rect 5094 14463 5095 14497
rect 5059 14429 5095 14463
rect 5059 14395 5060 14429
rect 5094 14395 5095 14429
rect 5059 14361 5095 14395
rect 5059 14327 5060 14361
rect 5094 14327 5095 14361
rect 5059 14293 5095 14327
rect 5059 14259 5060 14293
rect 5094 14259 5095 14293
rect 5059 14225 5095 14259
rect 5059 14191 5060 14225
rect 5094 14191 5095 14225
rect 5059 14157 5095 14191
rect 5059 14123 5060 14157
rect 5094 14123 5095 14157
rect 5059 14089 5095 14123
rect 5059 14055 5060 14089
rect 5094 14055 5095 14089
rect 5059 14021 5095 14055
rect 5059 13987 5060 14021
rect 5094 13987 5095 14021
rect 5059 13953 5095 13987
rect 5059 13919 5060 13953
rect 5094 13919 5095 13953
rect 5059 13885 5095 13919
rect 5059 13851 5060 13885
rect 5094 13851 5095 13885
rect 6303 14519 6304 14553
rect 6338 14519 6339 14553
rect 6303 14485 6339 14519
rect 6303 14451 6304 14485
rect 6338 14451 6339 14485
rect 6303 14417 6339 14451
rect 6303 14383 6304 14417
rect 6338 14383 6339 14417
rect 6303 14349 6339 14383
rect 6303 14315 6304 14349
rect 6338 14315 6339 14349
rect 6303 14281 6339 14315
rect 6303 14247 6304 14281
rect 6338 14247 6339 14281
rect 6303 14213 6339 14247
rect 6303 14179 6304 14213
rect 6338 14179 6339 14213
rect 6303 14145 6339 14179
rect 6303 14111 6304 14145
rect 6338 14111 6339 14145
rect 6303 14077 6339 14111
rect 6303 14043 6304 14077
rect 6338 14043 6339 14077
rect 6303 14009 6339 14043
rect 6303 13975 6304 14009
rect 6338 13975 6339 14009
rect 6303 13941 6339 13975
rect 6303 13907 6304 13941
rect 6338 13907 6339 13941
rect 5059 13817 5095 13851
rect 5059 13783 5060 13817
rect 5094 13783 5095 13817
rect 5059 13749 5095 13783
rect 5316 13876 5382 13882
rect 5316 13840 5332 13876
rect 5366 13840 5382 13876
rect 5316 13804 5382 13840
rect 5316 13770 5332 13804
rect 5366 13770 5382 13804
rect 5316 13764 5382 13770
rect 5456 13876 5522 13882
rect 5456 13874 5476 13876
rect 5456 13840 5472 13874
rect 5510 13842 5522 13876
rect 5506 13840 5522 13842
rect 5456 13804 5522 13840
rect 5456 13770 5476 13804
rect 5510 13770 5522 13804
rect 5456 13764 5522 13770
rect 6303 13873 6339 13907
rect 6303 13839 6304 13873
rect 6338 13839 6339 13873
rect 6303 13805 6339 13839
rect 6303 13771 6304 13805
rect 6338 13771 6339 13805
rect 5059 13715 5060 13749
rect 5094 13715 5095 13749
rect 5059 13681 5095 13715
rect 5059 13647 5060 13681
rect 5094 13647 5095 13681
rect 5059 13613 5095 13647
rect 5059 13579 5060 13613
rect 5094 13579 5095 13613
rect 5059 13545 5095 13579
rect 5059 13511 5060 13545
rect 5094 13511 5095 13545
rect 5059 13477 5095 13511
rect 5059 13443 5060 13477
rect 5094 13443 5095 13477
rect 5059 13409 5095 13443
rect 5059 13375 5060 13409
rect 5094 13375 5095 13409
rect 5059 13341 5095 13375
rect 5059 13307 5060 13341
rect 5094 13307 5095 13341
rect 5059 13273 5095 13307
rect 5059 13239 5060 13273
rect 5094 13239 5095 13273
rect 5059 13205 5095 13239
rect 5059 13171 5060 13205
rect 5094 13171 5095 13205
rect 5059 13137 5095 13171
rect 5059 13103 5060 13137
rect 5094 13103 5095 13137
rect 5059 13069 5095 13103
rect 5059 13035 5060 13069
rect 5094 13035 5095 13069
rect 5059 13001 5095 13035
rect 5059 12967 5060 13001
rect 5094 12967 5095 13001
rect 5059 12933 5095 12967
rect 5059 12899 5060 12933
rect 5094 12899 5095 12933
rect 5059 12865 5095 12899
rect 5059 12831 5060 12865
rect 5094 12831 5095 12865
rect 5059 12797 5095 12831
rect 5059 12763 5060 12797
rect 5094 12763 5095 12797
rect 5059 12729 5095 12763
rect 5059 12695 5060 12729
rect 5094 12695 5095 12729
rect 5059 12661 5095 12695
rect 5059 12627 5060 12661
rect 5094 12627 5095 12661
rect 5059 12593 5095 12627
rect 5059 12559 5060 12593
rect 5094 12559 5095 12593
rect 5059 12525 5095 12559
rect 5059 12491 5060 12525
rect 5094 12491 5095 12525
rect 5059 12457 5095 12491
rect 5059 12423 5060 12457
rect 5094 12423 5095 12457
rect 5059 12389 5095 12423
rect 5059 12355 5060 12389
rect 5094 12355 5095 12389
rect 5059 12321 5095 12355
rect 5059 12287 5060 12321
rect 5094 12287 5095 12321
rect 5059 12253 5095 12287
rect 5059 12219 5060 12253
rect 5094 12219 5095 12253
rect 5059 12185 5095 12219
rect 5059 12151 5060 12185
rect 5094 12151 5095 12185
rect 5059 12117 5095 12151
rect 350 12079 507 12113
rect 350 12045 351 12079
rect 385 12045 472 12079
rect 506 12045 507 12079
rect 350 12011 507 12045
rect 350 11977 351 12011
rect 385 11977 472 12011
rect 506 11977 507 12011
rect 2500 12078 2536 12113
rect 2500 12044 2501 12078
rect 2535 12044 2536 12078
rect 2500 12010 2536 12044
rect 350 11943 507 11977
rect 847 11971 863 12005
rect 900 11971 931 12005
rect 972 11971 981 12005
rect 1083 11971 1097 12005
rect 1133 11971 1167 12005
rect 1203 11971 1217 12005
rect 1319 11971 1333 12005
rect 1369 11971 1403 12005
rect 1439 11971 1453 12005
rect 1555 11971 1569 12005
rect 1605 11971 1639 12005
rect 1675 11971 1689 12005
rect 1791 11971 1805 12005
rect 1841 11971 1875 12005
rect 1911 11971 1925 12005
rect 2027 11971 2041 12005
rect 2077 11971 2111 12005
rect 2147 11971 2161 12005
rect 2500 11976 2501 12010
rect 2535 11976 2536 12010
rect 4528 12079 4686 12113
rect 4528 12045 4529 12079
rect 4563 12078 4686 12079
rect 4563 12045 4651 12078
rect 4528 12044 4651 12045
rect 4685 12044 4686 12078
rect 4528 12011 4686 12044
rect 350 11909 351 11943
rect 385 11909 472 11943
rect 506 11909 507 11943
rect 350 11875 507 11909
rect 350 11841 351 11875
rect 385 11841 472 11875
rect 506 11841 507 11875
rect 350 11807 507 11841
rect 350 11773 351 11807
rect 385 11773 472 11807
rect 506 11773 507 11807
rect 350 11739 507 11773
rect 350 11705 351 11739
rect 385 11705 472 11739
rect 506 11705 507 11739
rect 350 11671 507 11705
rect 350 11637 351 11671
rect 385 11637 472 11671
rect 506 11637 507 11671
rect 350 11603 507 11637
rect 350 11569 351 11603
rect 385 11569 472 11603
rect 506 11569 507 11603
rect 350 11535 507 11569
rect 350 11501 351 11535
rect 385 11501 472 11535
rect 506 11501 507 11535
rect 350 11467 507 11501
rect 350 11433 351 11467
rect 385 11433 472 11467
rect 506 11433 507 11467
rect 350 11399 507 11433
rect 350 11365 351 11399
rect 385 11365 472 11399
rect 506 11365 507 11399
rect 350 11331 507 11365
rect 350 11297 351 11331
rect 385 11297 472 11331
rect 506 11297 507 11331
rect 350 11263 507 11297
rect 350 11229 351 11263
rect 385 11229 472 11263
rect 506 11229 507 11263
rect 350 11195 507 11229
rect 350 11161 351 11195
rect 385 11161 472 11195
rect 506 11161 507 11195
rect 350 11127 507 11161
rect 350 11093 351 11127
rect 385 11093 472 11127
rect 506 11093 507 11127
rect 350 11059 507 11093
rect 350 11025 351 11059
rect 385 11025 472 11059
rect 506 11025 507 11059
rect 350 10991 507 11025
rect 350 10957 351 10991
rect 385 10957 472 10991
rect 506 10957 507 10991
rect 350 10923 507 10957
rect 350 10889 351 10923
rect 385 10889 472 10923
rect 506 10889 507 10923
rect 350 10855 507 10889
rect 350 10821 351 10855
rect 385 10821 472 10855
rect 506 10821 507 10855
rect 350 10787 507 10821
rect 350 10753 351 10787
rect 385 10753 472 10787
rect 506 10753 507 10787
rect 350 10719 507 10753
rect 350 10685 351 10719
rect 385 10685 472 10719
rect 506 10685 507 10719
rect 350 10651 507 10685
rect 350 10617 351 10651
rect 385 10617 472 10651
rect 506 10617 507 10651
rect 350 10583 507 10617
rect 350 10549 351 10583
rect 385 10549 472 10583
rect 506 10549 507 10583
rect 350 10515 507 10549
rect 350 10481 351 10515
rect 385 10481 472 10515
rect 506 10481 507 10515
rect 350 10447 507 10481
rect 350 10413 351 10447
rect 385 10413 472 10447
rect 506 10413 507 10447
rect 350 10379 507 10413
rect 350 10345 351 10379
rect 385 10345 472 10379
rect 506 10345 507 10379
rect 350 10311 507 10345
rect 350 10277 351 10311
rect 385 10277 472 10311
rect 506 10277 507 10311
rect 350 10243 507 10277
rect 350 10209 351 10243
rect 385 10209 472 10243
rect 506 10209 507 10243
rect 350 10175 507 10209
rect 350 10141 351 10175
rect 385 10141 472 10175
rect 506 10141 507 10175
rect 350 10107 507 10141
rect 350 10073 351 10107
rect 385 10073 472 10107
rect 506 10073 507 10107
rect 350 10039 507 10073
rect 350 10005 351 10039
rect 385 10005 472 10039
rect 506 10005 507 10039
rect 350 9971 507 10005
rect 350 9937 351 9971
rect 385 9937 472 9971
rect 506 9937 507 9971
rect 350 9903 507 9937
rect 350 9869 351 9903
rect 385 9869 472 9903
rect 506 9869 507 9903
rect 661 11926 697 11960
rect 661 11892 662 11926
rect 696 11892 697 11926
rect 661 11858 697 11892
rect 661 11824 662 11858
rect 696 11824 697 11858
rect 661 11790 697 11824
rect 661 11756 662 11790
rect 696 11756 697 11790
rect 661 11722 697 11756
rect 661 11688 662 11722
rect 696 11688 697 11722
rect 661 11654 697 11688
rect 661 11620 662 11654
rect 696 11620 697 11654
rect 661 11586 697 11620
rect 661 11552 662 11586
rect 696 11552 697 11586
rect 661 11518 697 11552
rect 661 11484 662 11518
rect 696 11484 697 11518
rect 661 11450 697 11484
rect 661 11416 662 11450
rect 696 11416 697 11450
rect 661 11382 697 11416
rect 661 11348 662 11382
rect 696 11348 697 11382
rect 661 11314 697 11348
rect 661 11280 662 11314
rect 696 11280 697 11314
rect 661 11246 697 11280
rect 661 11212 662 11246
rect 696 11212 697 11246
rect 661 11178 697 11212
rect 661 11144 662 11178
rect 696 11144 697 11178
rect 661 11110 697 11144
rect 661 11076 662 11110
rect 696 11076 697 11110
rect 661 11042 697 11076
rect 661 11008 662 11042
rect 696 11008 697 11042
rect 661 10974 697 11008
rect 661 10940 662 10974
rect 696 10940 697 10974
rect 661 10906 697 10940
rect 661 10872 662 10906
rect 696 10872 697 10906
rect 661 10838 697 10872
rect 661 10804 662 10838
rect 696 10804 697 10838
rect 661 10770 697 10804
rect 661 10736 662 10770
rect 696 10736 697 10770
rect 661 10702 697 10736
rect 661 10668 662 10702
rect 696 10668 697 10702
rect 661 10634 697 10668
rect 661 10600 662 10634
rect 696 10600 697 10634
rect 661 10566 697 10600
rect 661 10532 662 10566
rect 696 10532 697 10566
rect 661 10498 697 10532
rect 661 10464 662 10498
rect 696 10464 697 10498
rect 661 10430 697 10464
rect 661 10396 662 10430
rect 696 10396 697 10430
rect 661 10362 697 10396
rect 661 10328 662 10362
rect 696 10328 697 10362
rect 661 10294 697 10328
rect 661 10260 662 10294
rect 696 10260 697 10294
rect 661 10226 697 10260
rect 661 10192 662 10226
rect 696 10192 697 10226
rect 661 10158 697 10192
rect 661 10124 662 10158
rect 696 10124 697 10158
rect 661 10090 697 10124
rect 661 10056 662 10090
rect 696 10056 697 10090
rect 661 10022 697 10056
rect 661 9988 662 10022
rect 696 9988 697 10022
rect 661 9887 697 9988
rect 2311 11859 2347 11960
rect 2311 11825 2312 11859
rect 2346 11825 2347 11859
rect 2311 11791 2347 11825
rect 2311 11757 2312 11791
rect 2346 11757 2347 11791
rect 2311 11723 2347 11757
rect 2311 11689 2312 11723
rect 2346 11689 2347 11723
rect 2311 11655 2347 11689
rect 2311 11621 2312 11655
rect 2346 11621 2347 11655
rect 2311 11587 2347 11621
rect 2311 11553 2312 11587
rect 2346 11553 2347 11587
rect 2311 11519 2347 11553
rect 2311 11485 2312 11519
rect 2346 11485 2347 11519
rect 2311 11451 2347 11485
rect 2311 11417 2312 11451
rect 2346 11417 2347 11451
rect 2311 11383 2347 11417
rect 2311 11349 2312 11383
rect 2346 11349 2347 11383
rect 2311 11315 2347 11349
rect 2311 11281 2312 11315
rect 2346 11281 2347 11315
rect 2311 11247 2347 11281
rect 2311 11213 2312 11247
rect 2346 11213 2347 11247
rect 2311 11179 2347 11213
rect 2311 11145 2312 11179
rect 2346 11145 2347 11179
rect 2311 11111 2347 11145
rect 2311 11077 2312 11111
rect 2346 11077 2347 11111
rect 2311 11043 2347 11077
rect 2311 11009 2312 11043
rect 2346 11009 2347 11043
rect 2311 10975 2347 11009
rect 2311 10941 2312 10975
rect 2346 10941 2347 10975
rect 2311 10907 2347 10941
rect 2311 10873 2312 10907
rect 2346 10873 2347 10907
rect 2311 10839 2347 10873
rect 2311 10805 2312 10839
rect 2346 10805 2347 10839
rect 2311 10771 2347 10805
rect 2311 10737 2312 10771
rect 2346 10737 2347 10771
rect 2311 10703 2347 10737
rect 2311 10669 2312 10703
rect 2346 10669 2347 10703
rect 2311 10635 2347 10669
rect 2311 10601 2312 10635
rect 2346 10601 2347 10635
rect 2311 10567 2347 10601
rect 2311 10533 2312 10567
rect 2346 10533 2347 10567
rect 2311 10499 2347 10533
rect 2311 10465 2312 10499
rect 2346 10465 2347 10499
rect 2311 10431 2347 10465
rect 2311 10397 2312 10431
rect 2346 10397 2347 10431
rect 2311 10363 2347 10397
rect 2311 10329 2312 10363
rect 2346 10329 2347 10363
rect 2311 10295 2347 10329
rect 2311 10261 2312 10295
rect 2346 10261 2347 10295
rect 2311 10227 2347 10261
rect 2311 10193 2312 10227
rect 2346 10193 2347 10227
rect 2311 10159 2347 10193
rect 2311 10125 2312 10159
rect 2346 10125 2347 10159
rect 2311 10091 2347 10125
rect 2311 10057 2312 10091
rect 2346 10057 2347 10091
rect 2311 10023 2347 10057
rect 2500 11942 2536 11976
rect 2875 11971 2889 12005
rect 2925 11971 2959 12005
rect 2995 11971 3009 12005
rect 3111 11971 3125 12005
rect 3161 11971 3195 12005
rect 3231 11971 3245 12005
rect 3347 11971 3361 12005
rect 3397 11971 3431 12005
rect 3467 11971 3481 12005
rect 3583 11971 3597 12005
rect 3633 11971 3667 12005
rect 3703 11971 3717 12005
rect 3819 11971 3833 12005
rect 3869 11971 3903 12005
rect 3939 11971 3953 12005
rect 4055 11971 4064 12005
rect 4105 11971 4136 12005
rect 4173 11971 4189 12005
rect 4528 11977 4529 12011
rect 4563 12010 4686 12011
rect 4563 11977 4651 12010
rect 4528 11976 4651 11977
rect 4685 11976 4686 12010
rect 2500 11908 2501 11942
rect 2535 11908 2536 11942
rect 2500 11874 2536 11908
rect 2500 11840 2501 11874
rect 2535 11840 2536 11874
rect 2500 11806 2536 11840
rect 2500 11772 2501 11806
rect 2535 11772 2536 11806
rect 2500 11738 2536 11772
rect 2500 11704 2501 11738
rect 2535 11704 2536 11738
rect 2500 11670 2536 11704
rect 2500 11636 2501 11670
rect 2535 11636 2536 11670
rect 2500 11602 2536 11636
rect 2500 11568 2501 11602
rect 2535 11568 2536 11602
rect 2500 11534 2536 11568
rect 2500 11500 2501 11534
rect 2535 11500 2536 11534
rect 2500 11466 2536 11500
rect 2500 11432 2501 11466
rect 2535 11432 2536 11466
rect 2500 11398 2536 11432
rect 2500 11364 2501 11398
rect 2535 11364 2536 11398
rect 2500 11330 2536 11364
rect 2500 11296 2501 11330
rect 2535 11296 2536 11330
rect 2500 11262 2536 11296
rect 2500 11228 2501 11262
rect 2535 11228 2536 11262
rect 2500 11194 2536 11228
rect 2500 11160 2501 11194
rect 2535 11160 2536 11194
rect 2500 11126 2536 11160
rect 2500 11092 2501 11126
rect 2535 11092 2536 11126
rect 2500 11058 2536 11092
rect 2500 11024 2501 11058
rect 2535 11024 2536 11058
rect 2500 10990 2536 11024
rect 2500 10956 2501 10990
rect 2535 10956 2536 10990
rect 2500 10922 2536 10956
rect 2500 10888 2501 10922
rect 2535 10888 2536 10922
rect 2500 10854 2536 10888
rect 2500 10820 2501 10854
rect 2535 10820 2536 10854
rect 2500 10786 2536 10820
rect 2500 10752 2501 10786
rect 2535 10752 2536 10786
rect 2500 10718 2536 10752
rect 2500 10684 2501 10718
rect 2535 10684 2536 10718
rect 2500 10650 2536 10684
rect 2500 10616 2501 10650
rect 2535 10616 2536 10650
rect 2500 10582 2536 10616
rect 2500 10548 2501 10582
rect 2535 10548 2536 10582
rect 2500 10514 2536 10548
rect 2500 10480 2501 10514
rect 2535 10480 2536 10514
rect 2500 10446 2536 10480
rect 2500 10412 2501 10446
rect 2535 10412 2536 10446
rect 2500 10378 2536 10412
rect 2500 10344 2501 10378
rect 2535 10344 2536 10378
rect 2500 10310 2536 10344
rect 2500 10276 2501 10310
rect 2535 10276 2536 10310
rect 2500 10242 2536 10276
rect 2500 10208 2501 10242
rect 2535 10208 2536 10242
rect 2500 10174 2536 10208
rect 2500 10140 2501 10174
rect 2535 10140 2536 10174
rect 2500 10106 2536 10140
rect 2500 10072 2501 10106
rect 2535 10072 2536 10106
rect 2500 10038 2536 10072
rect 2311 9989 2312 10023
rect 2346 9989 2347 10023
rect 2311 9955 2347 9989
rect 2311 9921 2312 9955
rect 2346 9921 2347 9955
rect 350 9835 507 9869
rect 350 9801 351 9835
rect 385 9801 472 9835
rect 506 9801 507 9835
rect 350 9767 507 9801
rect 350 9733 351 9767
rect 385 9733 472 9767
rect 506 9733 507 9767
rect 350 9699 507 9733
rect 350 9665 351 9699
rect 385 9698 507 9699
rect 542 9879 627 9885
rect 542 9845 569 9879
rect 603 9845 627 9879
rect 1015 9875 1049 9919
rect 1487 9875 1521 9919
rect 1959 9875 1993 9919
rect 2311 9887 2347 9921
rect 2381 10019 2466 10025
rect 2381 9985 2405 10019
rect 2439 9985 2466 10019
rect 2381 9947 2466 9985
rect 2381 9913 2405 9947
rect 2439 9913 2466 9947
rect 542 9807 627 9845
rect 847 9841 863 9875
rect 897 9841 931 9875
rect 965 9841 1099 9875
rect 1133 9841 1167 9875
rect 1201 9841 1335 9875
rect 1369 9841 1403 9875
rect 1437 9841 1571 9875
rect 1605 9841 1639 9875
rect 1673 9841 1807 9875
rect 1841 9841 1875 9875
rect 1909 9841 2043 9875
rect 2077 9841 2111 9875
rect 2145 9841 2161 9875
rect 542 9773 569 9807
rect 603 9773 627 9807
rect 385 9665 386 9698
rect 350 9631 386 9665
rect 350 9597 351 9631
rect 385 9597 386 9631
rect 350 9563 386 9597
rect 542 9653 627 9773
rect 662 9733 2347 9734
rect 662 9699 710 9733
rect 744 9699 778 9733
rect 812 9699 846 9733
rect 880 9699 914 9733
rect 948 9699 982 9733
rect 1016 9699 1050 9733
rect 1084 9699 1118 9733
rect 1152 9699 1186 9733
rect 1220 9699 1254 9733
rect 1288 9699 1322 9733
rect 1356 9699 1390 9733
rect 1424 9699 1458 9733
rect 1492 9699 1526 9733
rect 1560 9699 1594 9733
rect 1628 9699 1662 9733
rect 1696 9699 1730 9733
rect 1764 9699 1798 9733
rect 1832 9699 1866 9733
rect 1900 9699 1934 9733
rect 1968 9699 2002 9733
rect 2036 9699 2070 9733
rect 2104 9699 2138 9733
rect 2172 9699 2206 9733
rect 2240 9699 2274 9733
rect 2308 9699 2347 9733
rect 662 9698 2347 9699
rect 2381 9653 2466 9913
rect 2500 10004 2501 10038
rect 2535 10004 2536 10038
rect 2689 11926 2725 11960
rect 2689 11892 2690 11926
rect 2724 11892 2725 11926
rect 2689 11858 2725 11892
rect 2689 11824 2690 11858
rect 2724 11824 2725 11858
rect 2689 11790 2725 11824
rect 2689 11756 2690 11790
rect 2724 11756 2725 11790
rect 2689 11722 2725 11756
rect 2689 11688 2690 11722
rect 2724 11688 2725 11722
rect 2689 11654 2725 11688
rect 2689 11620 2690 11654
rect 2724 11620 2725 11654
rect 2689 11586 2725 11620
rect 2689 11552 2690 11586
rect 2724 11552 2725 11586
rect 2689 11518 2725 11552
rect 2689 11484 2690 11518
rect 2724 11484 2725 11518
rect 2689 11450 2725 11484
rect 2689 11416 2690 11450
rect 2724 11416 2725 11450
rect 2689 11382 2725 11416
rect 2689 11348 2690 11382
rect 2724 11348 2725 11382
rect 2689 11314 2725 11348
rect 2689 11280 2690 11314
rect 2724 11280 2725 11314
rect 2689 11246 2725 11280
rect 2689 11212 2690 11246
rect 2724 11212 2725 11246
rect 2689 11178 2725 11212
rect 2689 11144 2690 11178
rect 2724 11144 2725 11178
rect 2689 11110 2725 11144
rect 2689 11076 2690 11110
rect 2724 11076 2725 11110
rect 2689 11042 2725 11076
rect 2689 11008 2690 11042
rect 2724 11008 2725 11042
rect 2689 10974 2725 11008
rect 2689 10940 2690 10974
rect 2724 10940 2725 10974
rect 2689 10906 2725 10940
rect 2689 10872 2690 10906
rect 2724 10872 2725 10906
rect 2689 10838 2725 10872
rect 2689 10804 2690 10838
rect 2724 10804 2725 10838
rect 2689 10770 2725 10804
rect 2689 10736 2690 10770
rect 2724 10736 2725 10770
rect 2689 10702 2725 10736
rect 2689 10668 2690 10702
rect 2724 10668 2725 10702
rect 2689 10634 2725 10668
rect 2689 10600 2690 10634
rect 2724 10600 2725 10634
rect 2689 10566 2725 10600
rect 2689 10532 2690 10566
rect 2724 10532 2725 10566
rect 2689 10498 2725 10532
rect 2689 10464 2690 10498
rect 2724 10464 2725 10498
rect 2689 10430 2725 10464
rect 2689 10396 2690 10430
rect 2724 10396 2725 10430
rect 2689 10362 2725 10396
rect 2689 10328 2690 10362
rect 2724 10328 2725 10362
rect 2689 10294 2725 10328
rect 2689 10260 2690 10294
rect 2724 10260 2725 10294
rect 2689 10226 2725 10260
rect 2689 10192 2690 10226
rect 2724 10192 2725 10226
rect 2689 10158 2725 10192
rect 2689 10124 2690 10158
rect 2724 10124 2725 10158
rect 2689 10090 2725 10124
rect 2689 10056 2690 10090
rect 2724 10056 2725 10090
rect 2500 9970 2536 10004
rect 2500 9936 2501 9970
rect 2535 9936 2536 9970
rect 2500 9902 2536 9936
rect 2500 9868 2501 9902
rect 2535 9868 2536 9902
rect 2500 9834 2536 9868
rect 2500 9800 2501 9834
rect 2535 9800 2536 9834
rect 2500 9766 2536 9800
rect 2500 9732 2501 9766
rect 2535 9732 2536 9766
rect 2500 9698 2536 9732
rect 2570 10019 2655 10025
rect 2570 9985 2597 10019
rect 2631 9985 2655 10019
rect 2570 9947 2655 9985
rect 2570 9913 2597 9947
rect 2631 9913 2655 9947
rect 2570 9653 2655 9913
rect 2689 10022 2725 10056
rect 2689 9988 2690 10022
rect 2724 9988 2725 10022
rect 2689 9887 2725 9988
rect 4339 11859 4375 11960
rect 4339 11825 4340 11859
rect 4374 11825 4375 11859
rect 4339 11791 4375 11825
rect 4339 11757 4340 11791
rect 4374 11757 4375 11791
rect 4339 11723 4375 11757
rect 4339 11689 4340 11723
rect 4374 11689 4375 11723
rect 4339 11655 4375 11689
rect 4339 11621 4340 11655
rect 4374 11621 4375 11655
rect 4339 11587 4375 11621
rect 4339 11553 4340 11587
rect 4374 11553 4375 11587
rect 4339 11519 4375 11553
rect 4339 11485 4340 11519
rect 4374 11485 4375 11519
rect 4339 11451 4375 11485
rect 4339 11417 4340 11451
rect 4374 11417 4375 11451
rect 4339 11383 4375 11417
rect 4339 11349 4340 11383
rect 4374 11349 4375 11383
rect 4339 11315 4375 11349
rect 4339 11281 4340 11315
rect 4374 11281 4375 11315
rect 4339 11247 4375 11281
rect 4339 11213 4340 11247
rect 4374 11213 4375 11247
rect 4339 11179 4375 11213
rect 4339 11145 4340 11179
rect 4374 11145 4375 11179
rect 4339 11111 4375 11145
rect 4339 11077 4340 11111
rect 4374 11077 4375 11111
rect 4339 11043 4375 11077
rect 4339 11009 4340 11043
rect 4374 11009 4375 11043
rect 4339 10975 4375 11009
rect 4339 10941 4340 10975
rect 4374 10941 4375 10975
rect 4339 10907 4375 10941
rect 4339 10873 4340 10907
rect 4374 10873 4375 10907
rect 4339 10839 4375 10873
rect 4339 10805 4340 10839
rect 4374 10805 4375 10839
rect 4339 10771 4375 10805
rect 4339 10737 4340 10771
rect 4374 10737 4375 10771
rect 4339 10703 4375 10737
rect 4339 10669 4340 10703
rect 4374 10669 4375 10703
rect 4339 10635 4375 10669
rect 4339 10601 4340 10635
rect 4374 10601 4375 10635
rect 4339 10567 4375 10601
rect 4339 10533 4340 10567
rect 4374 10533 4375 10567
rect 4339 10499 4375 10533
rect 4339 10465 4340 10499
rect 4374 10465 4375 10499
rect 4339 10431 4375 10465
rect 4339 10397 4340 10431
rect 4374 10397 4375 10431
rect 4339 10363 4375 10397
rect 4339 10329 4340 10363
rect 4374 10329 4375 10363
rect 4339 10295 4375 10329
rect 4339 10261 4340 10295
rect 4374 10261 4375 10295
rect 4339 10227 4375 10261
rect 4339 10193 4340 10227
rect 4374 10193 4375 10227
rect 4339 10159 4375 10193
rect 4339 10125 4340 10159
rect 4374 10125 4375 10159
rect 4339 10091 4375 10125
rect 4339 10057 4340 10091
rect 4374 10057 4375 10091
rect 4339 10023 4375 10057
rect 4528 11943 4686 11976
rect 4528 11909 4529 11943
rect 4563 11942 4686 11943
rect 4563 11909 4651 11942
rect 4528 11908 4651 11909
rect 4685 11908 4686 11942
rect 4528 11875 4686 11908
rect 4528 11841 4529 11875
rect 4563 11874 4686 11875
rect 4563 11841 4651 11874
rect 4528 11840 4651 11841
rect 4685 11840 4686 11874
rect 4528 11807 4686 11840
rect 4528 11773 4529 11807
rect 4563 11806 4686 11807
rect 4563 11773 4651 11806
rect 4528 11772 4651 11773
rect 4685 11772 4686 11806
rect 4528 11739 4686 11772
rect 4528 11705 4529 11739
rect 4563 11738 4686 11739
rect 4563 11705 4651 11738
rect 4528 11704 4651 11705
rect 4685 11704 4686 11738
rect 4528 11671 4686 11704
rect 4528 11637 4529 11671
rect 4563 11670 4686 11671
rect 4563 11637 4651 11670
rect 4528 11636 4651 11637
rect 4685 11636 4686 11670
rect 4528 11603 4686 11636
rect 4528 11569 4529 11603
rect 4563 11602 4686 11603
rect 4563 11569 4651 11602
rect 4528 11568 4651 11569
rect 4685 11568 4686 11602
rect 4528 11535 4686 11568
rect 4528 11501 4529 11535
rect 4563 11534 4686 11535
rect 4563 11501 4651 11534
rect 4528 11500 4651 11501
rect 4685 11500 4686 11534
rect 4528 11467 4686 11500
rect 4528 11433 4529 11467
rect 4563 11466 4686 11467
rect 4563 11433 4651 11466
rect 4528 11432 4651 11433
rect 4685 11432 4686 11466
rect 4528 11399 4686 11432
rect 4528 11365 4529 11399
rect 4563 11398 4686 11399
rect 4563 11365 4651 11398
rect 4528 11364 4651 11365
rect 4685 11364 4686 11398
rect 4528 11331 4686 11364
rect 4528 11297 4529 11331
rect 4563 11330 4686 11331
rect 4563 11297 4651 11330
rect 4528 11296 4651 11297
rect 4685 11296 4686 11330
rect 4528 11263 4686 11296
rect 4528 11229 4529 11263
rect 4563 11262 4686 11263
rect 4563 11229 4651 11262
rect 4528 11228 4651 11229
rect 4685 11228 4686 11262
rect 4528 11195 4686 11228
rect 4528 11161 4529 11195
rect 4563 11194 4686 11195
rect 4563 11161 4651 11194
rect 4528 11160 4651 11161
rect 4685 11160 4686 11194
rect 4528 11127 4686 11160
rect 4528 11093 4529 11127
rect 4563 11126 4686 11127
rect 4563 11093 4651 11126
rect 4528 11092 4651 11093
rect 4685 11092 4686 11126
rect 4528 11059 4686 11092
rect 4528 11025 4529 11059
rect 4563 11058 4686 11059
rect 4563 11025 4651 11058
rect 4528 11024 4651 11025
rect 4685 11024 4686 11058
rect 4528 10991 4686 11024
rect 4528 10957 4529 10991
rect 4563 10990 4686 10991
rect 4563 10957 4651 10990
rect 4528 10956 4651 10957
rect 4685 10956 4686 10990
rect 4528 10923 4686 10956
rect 4528 10889 4529 10923
rect 4563 10922 4686 10923
rect 4563 10889 4651 10922
rect 4528 10888 4651 10889
rect 4685 10888 4686 10922
rect 4528 10855 4686 10888
rect 4528 10821 4529 10855
rect 4563 10854 4686 10855
rect 4563 10821 4651 10854
rect 4528 10820 4651 10821
rect 4685 10820 4686 10854
rect 4528 10787 4686 10820
rect 4528 10753 4529 10787
rect 4563 10786 4686 10787
rect 4563 10753 4651 10786
rect 4528 10752 4651 10753
rect 4685 10752 4686 10786
rect 4528 10719 4686 10752
rect 4528 10685 4529 10719
rect 4563 10718 4686 10719
rect 4563 10685 4651 10718
rect 4528 10684 4651 10685
rect 4685 10684 4686 10718
rect 4528 10651 4686 10684
rect 4528 10617 4529 10651
rect 4563 10650 4686 10651
rect 4563 10617 4651 10650
rect 4528 10616 4651 10617
rect 4685 10616 4686 10650
rect 4528 10583 4686 10616
rect 4528 10549 4529 10583
rect 4563 10582 4686 10583
rect 4563 10549 4651 10582
rect 4528 10548 4651 10549
rect 4685 10548 4686 10582
rect 4528 10515 4686 10548
rect 4528 10481 4529 10515
rect 4563 10514 4686 10515
rect 4563 10481 4651 10514
rect 4528 10480 4651 10481
rect 4685 10480 4686 10514
rect 4528 10447 4686 10480
rect 4528 10413 4529 10447
rect 4563 10446 4686 10447
rect 4563 10413 4651 10446
rect 4528 10412 4651 10413
rect 4685 10412 4686 10446
rect 4528 10379 4686 10412
rect 4528 10345 4529 10379
rect 4563 10378 4686 10379
rect 4563 10345 4651 10378
rect 4528 10344 4651 10345
rect 4685 10344 4686 10378
rect 4528 10311 4686 10344
rect 4528 10277 4529 10311
rect 4563 10310 4686 10311
rect 4563 10277 4651 10310
rect 4528 10276 4651 10277
rect 4685 10276 4686 10310
rect 4528 10243 4686 10276
rect 4528 10209 4529 10243
rect 4563 10242 4686 10243
rect 4563 10209 4651 10242
rect 4528 10208 4651 10209
rect 4685 10208 4686 10242
rect 4528 10175 4686 10208
rect 4528 10141 4529 10175
rect 4563 10174 4686 10175
rect 4563 10141 4651 10174
rect 4528 10140 4651 10141
rect 4685 10140 4686 10174
rect 4528 10107 4686 10140
rect 4528 10073 4529 10107
rect 4563 10106 4686 10107
rect 4563 10073 4651 10106
rect 4528 10072 4651 10073
rect 4685 10072 4686 10106
rect 5059 12083 5060 12117
rect 5094 12083 5095 12117
rect 5059 12049 5095 12083
rect 5059 12015 5060 12049
rect 5094 12015 5095 12049
rect 5059 11981 5095 12015
rect 5059 11947 5060 11981
rect 5094 11947 5095 11981
rect 5059 11913 5095 11947
rect 5059 11879 5060 11913
rect 5094 11879 5095 11913
rect 5059 11845 5095 11879
rect 5059 11811 5060 11845
rect 5094 11811 5095 11845
rect 5059 11777 5095 11811
rect 5059 11743 5060 11777
rect 5094 11743 5095 11777
rect 5059 11709 5095 11743
rect 5059 11675 5060 11709
rect 5094 11675 5095 11709
rect 5059 11641 5095 11675
rect 5059 11607 5060 11641
rect 5094 11607 5095 11641
rect 5059 11573 5095 11607
rect 5059 11539 5060 11573
rect 5094 11539 5095 11573
rect 5059 11505 5095 11539
rect 5059 11471 5060 11505
rect 5094 11471 5095 11505
rect 5059 11437 5095 11471
rect 5059 11403 5060 11437
rect 5094 11403 5095 11437
rect 5059 11369 5095 11403
rect 5059 11335 5060 11369
rect 5094 11335 5095 11369
rect 5059 11301 5095 11335
rect 5059 11267 5060 11301
rect 5094 11267 5095 11301
rect 5059 11233 5095 11267
rect 5059 11199 5060 11233
rect 5094 11199 5095 11233
rect 5059 11165 5095 11199
rect 5059 11131 5060 11165
rect 5094 11131 5095 11165
rect 5059 11097 5095 11131
rect 5059 11063 5060 11097
rect 5094 11063 5095 11097
rect 5059 11029 5095 11063
rect 5059 10995 5060 11029
rect 5094 10995 5095 11029
rect 5059 10961 5095 10995
rect 5059 10927 5060 10961
rect 5094 10927 5095 10961
rect 5059 10893 5095 10927
rect 5059 10859 5060 10893
rect 5094 10859 5095 10893
rect 5059 10825 5095 10859
rect 5059 10791 5060 10825
rect 5094 10791 5095 10825
rect 5059 10757 5095 10791
rect 5059 10723 5060 10757
rect 5094 10723 5095 10757
rect 5059 10689 5095 10723
rect 5059 10655 5060 10689
rect 5094 10655 5095 10689
rect 5059 10621 5095 10655
rect 5059 10587 5060 10621
rect 5094 10587 5095 10621
rect 5059 10553 5095 10587
rect 5059 10519 5060 10553
rect 5094 10519 5095 10553
rect 5059 10485 5095 10519
rect 5059 10451 5060 10485
rect 5094 10451 5095 10485
rect 5059 10417 5095 10451
rect 5059 10383 5060 10417
rect 5094 10383 5095 10417
rect 6303 13737 6339 13771
rect 6303 13703 6304 13737
rect 6338 13703 6339 13737
rect 6303 13669 6339 13703
rect 6303 13635 6304 13669
rect 6338 13635 6339 13669
rect 6303 13601 6339 13635
rect 6303 13567 6304 13601
rect 6338 13567 6339 13601
rect 6303 13533 6339 13567
rect 6303 13499 6304 13533
rect 6338 13499 6339 13533
rect 6303 13465 6339 13499
rect 6303 13431 6304 13465
rect 6338 13431 6339 13465
rect 6303 13397 6339 13431
rect 6303 13363 6304 13397
rect 6338 13363 6339 13397
rect 6303 13329 6339 13363
rect 6303 13295 6304 13329
rect 6338 13295 6339 13329
rect 6303 13261 6339 13295
rect 6303 13227 6304 13261
rect 6338 13227 6339 13261
rect 6303 13193 6339 13227
rect 6303 13159 6304 13193
rect 6338 13159 6339 13193
rect 6303 13125 6339 13159
rect 6303 13091 6304 13125
rect 6338 13091 6339 13125
rect 6303 13057 6339 13091
rect 6303 13023 6304 13057
rect 6338 13023 6339 13057
rect 6303 12989 6339 13023
rect 6303 12955 6304 12989
rect 6338 12955 6339 12989
rect 6303 12921 6339 12955
rect 6303 12887 6304 12921
rect 6338 12887 6339 12921
rect 6303 12853 6339 12887
rect 6303 12819 6304 12853
rect 6338 12819 6339 12853
rect 6303 12785 6339 12819
rect 6303 12751 6304 12785
rect 6338 12751 6339 12785
rect 6303 12717 6339 12751
rect 6303 12683 6304 12717
rect 6338 12683 6339 12717
rect 6303 12649 6339 12683
rect 6303 12615 6304 12649
rect 6338 12615 6339 12649
rect 6303 12581 6339 12615
rect 6303 12547 6304 12581
rect 6338 12547 6339 12581
rect 6303 12513 6339 12547
rect 6303 12479 6304 12513
rect 6338 12479 6339 12513
rect 6303 12445 6339 12479
rect 6303 12411 6304 12445
rect 6338 12411 6339 12445
rect 6303 12377 6339 12411
rect 6303 12343 6304 12377
rect 6338 12343 6339 12377
rect 6303 12309 6339 12343
rect 6303 12275 6304 12309
rect 6338 12275 6339 12309
rect 6303 12241 6339 12275
rect 6303 12207 6304 12241
rect 6338 12207 6339 12241
rect 6303 12173 6339 12207
rect 6303 12139 6304 12173
rect 6338 12139 6339 12173
rect 6303 12105 6339 12139
rect 6303 12071 6304 12105
rect 6338 12071 6339 12105
rect 6303 12037 6339 12071
rect 6303 12003 6304 12037
rect 6338 12003 6339 12037
rect 6303 11969 6339 12003
rect 6303 11935 6304 11969
rect 6338 11935 6339 11969
rect 6303 11901 6339 11935
rect 6303 11867 6304 11901
rect 6338 11867 6339 11901
rect 6303 11833 6339 11867
rect 6303 11799 6304 11833
rect 6338 11799 6339 11833
rect 6303 11765 6339 11799
rect 6303 11731 6304 11765
rect 6338 11731 6339 11765
rect 6303 11697 6339 11731
rect 6303 11663 6304 11697
rect 6338 11663 6339 11697
rect 6303 11629 6339 11663
rect 6303 11595 6304 11629
rect 6338 11595 6339 11629
rect 6303 11561 6339 11595
rect 6303 11527 6304 11561
rect 6338 11527 6339 11561
rect 6303 11493 6339 11527
rect 6303 11459 6304 11493
rect 6338 11459 6339 11493
rect 6303 11425 6339 11459
rect 6303 11391 6304 11425
rect 6338 11391 6339 11425
rect 6303 11357 6339 11391
rect 6303 11323 6304 11357
rect 6338 11323 6339 11357
rect 6303 11289 6339 11323
rect 6303 11255 6304 11289
rect 6338 11255 6339 11289
rect 6303 11221 6339 11255
rect 6303 11187 6304 11221
rect 6338 11187 6339 11221
rect 6303 11153 6339 11187
rect 6303 11119 6304 11153
rect 6338 11119 6339 11153
rect 6303 11085 6339 11119
rect 6303 11051 6304 11085
rect 6338 11051 6339 11085
rect 6303 10972 6339 11051
rect 6303 10938 6304 10972
rect 6338 10938 6339 10972
rect 6303 10904 6339 10938
rect 6303 10870 6304 10904
rect 6338 10870 6339 10904
rect 6303 10836 6339 10870
rect 6303 10802 6304 10836
rect 6338 10802 6339 10836
rect 6303 10768 6339 10802
rect 6303 10734 6304 10768
rect 6338 10734 6339 10768
rect 6303 10700 6339 10734
rect 6303 10666 6304 10700
rect 6338 10666 6339 10700
rect 6303 10632 6339 10666
rect 6303 10598 6304 10632
rect 6338 10598 6339 10632
rect 6303 10564 6339 10598
rect 6303 10530 6304 10564
rect 6338 10530 6339 10564
rect 6303 10496 6339 10530
rect 6303 10462 6304 10496
rect 6338 10462 6339 10496
rect 6303 10428 6339 10462
rect 6303 10394 6304 10428
rect 6338 10394 6339 10428
rect 5059 10349 5095 10383
rect 5059 10315 5060 10349
rect 5094 10315 5095 10349
rect 5059 10281 5095 10315
rect 5316 10381 5382 10387
rect 5316 10347 5332 10381
rect 5366 10347 5382 10381
rect 5316 10309 5382 10347
rect 5059 10247 5060 10281
rect 5094 10247 5095 10281
rect 5192 10263 5226 10265
rect 5316 10275 5332 10309
rect 5366 10275 5382 10309
rect 5059 10213 5095 10247
rect 5059 10179 5060 10213
rect 5094 10179 5095 10213
rect 5176 10229 5242 10263
rect 5176 10195 5192 10229
rect 5226 10195 5242 10229
rect 5316 10229 5382 10275
rect 5316 10195 5332 10229
rect 5366 10195 5382 10229
rect 5456 10381 5522 10387
rect 5456 10347 5472 10381
rect 5506 10347 5522 10381
rect 5456 10309 5522 10347
rect 5456 10275 5472 10309
rect 5506 10275 5522 10309
rect 5456 10229 5522 10275
rect 5456 10195 5472 10229
rect 5506 10195 5522 10229
rect 5596 10381 5662 10387
rect 5596 10347 5616 10381
rect 5650 10347 5662 10381
rect 5596 10309 5662 10347
rect 5596 10275 5616 10309
rect 5650 10275 5662 10309
rect 5596 10229 5662 10275
rect 5596 10195 5612 10229
rect 5646 10195 5662 10229
rect 5736 10381 5802 10387
rect 5736 10347 5752 10381
rect 5786 10347 5802 10381
rect 5736 10309 5802 10347
rect 5736 10275 5752 10309
rect 5786 10275 5802 10309
rect 5736 10229 5802 10275
rect 5736 10195 5752 10229
rect 5786 10195 5802 10229
rect 5876 10381 5942 10387
rect 5876 10347 5896 10381
rect 5930 10347 5942 10381
rect 5876 10309 5942 10347
rect 5876 10275 5896 10309
rect 5930 10275 5942 10309
rect 5876 10229 5942 10275
rect 5876 10195 5892 10229
rect 5926 10195 5942 10229
rect 6016 10381 6082 10387
rect 6016 10347 6032 10381
rect 6066 10347 6082 10381
rect 6016 10309 6082 10347
rect 6016 10275 6032 10309
rect 6066 10275 6082 10309
rect 6016 10229 6082 10275
rect 6016 10195 6032 10229
rect 6066 10195 6082 10229
rect 6156 10381 6222 10387
rect 6156 10347 6172 10381
rect 6206 10347 6222 10381
rect 6156 10309 6222 10347
rect 6156 10275 6172 10309
rect 6206 10275 6222 10309
rect 6156 10229 6222 10275
rect 6156 10195 6172 10229
rect 6206 10195 6222 10229
rect 6303 10360 6339 10394
rect 6303 10326 6304 10360
rect 6338 10326 6339 10360
rect 6303 10292 6339 10326
rect 6303 10258 6304 10292
rect 6338 10258 6339 10292
rect 6303 10224 6339 10258
rect 5059 10145 5095 10179
rect 5059 10111 5060 10145
rect 5094 10113 5095 10145
rect 6303 10190 6304 10224
rect 6338 10190 6339 10224
rect 6303 10113 6339 10190
rect 5094 10112 6339 10113
rect 5094 10111 5183 10112
rect 5059 10078 5183 10111
rect 5217 10078 5251 10112
rect 5285 10078 5319 10112
rect 5353 10078 5387 10112
rect 5421 10078 5455 10112
rect 5489 10078 5523 10112
rect 5557 10078 5591 10112
rect 5625 10078 5659 10112
rect 5693 10078 5727 10112
rect 5761 10078 5795 10112
rect 5829 10078 5863 10112
rect 5897 10078 5931 10112
rect 5965 10078 5999 10112
rect 6033 10078 6067 10112
rect 6101 10078 6135 10112
rect 6169 10078 6203 10112
rect 6237 10078 6271 10112
rect 6305 10078 6339 10112
rect 5059 10077 6339 10078
rect 4339 9989 4340 10023
rect 4374 9989 4375 10023
rect 4339 9955 4375 9989
rect 4339 9921 4340 9955
rect 4374 9921 4375 9955
rect 3043 9875 3077 9919
rect 3515 9875 3549 9919
rect 3987 9875 4021 9919
rect 4339 9887 4375 9921
rect 4409 10036 4494 10042
rect 4409 10002 4433 10036
rect 4467 10002 4494 10036
rect 4409 9964 4494 10002
rect 4409 9930 4433 9964
rect 4467 9930 4494 9964
rect 2875 9841 2891 9875
rect 2925 9841 2959 9875
rect 2993 9841 3127 9875
rect 3161 9841 3195 9875
rect 3229 9841 3363 9875
rect 3397 9841 3431 9875
rect 3465 9841 3599 9875
rect 3633 9841 3667 9875
rect 3701 9841 3835 9875
rect 3869 9841 3903 9875
rect 3937 9841 4071 9875
rect 4105 9841 4139 9875
rect 4173 9841 4189 9875
rect 2689 9733 4375 9734
rect 2689 9699 2728 9733
rect 2762 9699 2796 9733
rect 2830 9699 2864 9733
rect 2898 9699 2932 9733
rect 2966 9699 3000 9733
rect 3034 9699 3068 9733
rect 3102 9699 3136 9733
rect 3170 9699 3204 9733
rect 3238 9699 3272 9733
rect 3306 9699 3340 9733
rect 3374 9699 3408 9733
rect 3442 9699 3476 9733
rect 3510 9699 3544 9733
rect 3578 9699 3612 9733
rect 3646 9699 3680 9733
rect 3714 9699 3748 9733
rect 3782 9699 3816 9733
rect 3850 9699 3884 9733
rect 3918 9699 3952 9733
rect 3986 9699 4020 9733
rect 4054 9699 4088 9733
rect 4122 9699 4156 9733
rect 4190 9699 4224 9733
rect 4258 9699 4292 9733
rect 4326 9699 4375 9733
rect 2689 9698 4375 9699
rect 4409 9653 4494 9930
rect 4528 10039 4686 10072
rect 4528 10005 4529 10039
rect 4563 10038 4686 10039
rect 4563 10005 4651 10038
rect 4528 10004 4651 10005
rect 4685 10004 4686 10038
rect 4528 9971 4686 10004
rect 4528 9937 4529 9971
rect 4563 9970 4686 9971
rect 4563 9937 4651 9970
rect 4528 9936 4651 9937
rect 4685 9936 4686 9970
rect 4528 9903 4686 9936
rect 4528 9869 4529 9903
rect 4563 9902 4686 9903
rect 4563 9869 4651 9902
rect 4528 9868 4651 9869
rect 4685 9868 4686 9902
rect 4528 9835 4686 9868
rect 4528 9801 4529 9835
rect 4563 9834 4686 9835
rect 4563 9801 4651 9834
rect 4528 9800 4651 9801
rect 4685 9800 4686 9834
rect 4528 9767 4686 9800
rect 4528 9733 4529 9767
rect 4563 9766 4686 9767
rect 4563 9733 4651 9766
rect 4528 9732 4651 9733
rect 4685 9734 4686 9766
rect 4685 9733 6054 9734
rect 4685 9732 4762 9733
rect 4528 9699 4762 9732
rect 4796 9699 4830 9733
rect 4864 9699 4898 9733
rect 4932 9699 4966 9733
rect 5000 9699 5034 9733
rect 5068 9699 5102 9733
rect 5136 9699 5170 9733
rect 5204 9699 5238 9733
rect 5272 9699 5306 9733
rect 5340 9699 5374 9733
rect 5408 9699 5442 9733
rect 5476 9699 5510 9733
rect 5544 9699 5578 9733
rect 5612 9699 5646 9733
rect 5680 9699 5714 9733
rect 5748 9699 5782 9733
rect 5816 9699 5850 9733
rect 5884 9699 5918 9733
rect 5952 9699 5986 9733
rect 6020 9699 6054 9733
rect 4528 9698 6054 9699
rect 4528 9660 4686 9698
rect 542 9638 660 9653
rect 542 9604 548 9638
rect 582 9604 620 9638
rect 654 9604 660 9638
rect 542 9589 660 9604
rect 2348 9638 2688 9653
rect 2348 9604 2354 9638
rect 2388 9604 2426 9638
rect 2460 9604 2576 9638
rect 2610 9604 2648 9638
rect 2682 9604 2688 9638
rect 2348 9589 2688 9604
rect 4376 9638 4494 9653
rect 4376 9604 4382 9638
rect 4416 9604 4454 9638
rect 4488 9604 4494 9638
rect 4376 9589 4494 9604
rect 6018 9650 6054 9698
rect 6018 9616 6019 9650
rect 6053 9616 6054 9650
rect 350 9529 351 9563
rect 385 9529 386 9563
rect 6018 9582 6054 9616
rect 6018 9548 6019 9582
rect 6053 9548 6054 9582
rect 350 9495 386 9529
rect 350 9461 351 9495
rect 385 9461 386 9495
rect 350 9427 386 9461
rect 350 9393 351 9427
rect 385 9393 386 9427
rect 350 9359 386 9393
rect 350 9325 351 9359
rect 385 9325 386 9359
rect 350 9291 386 9325
rect 350 9257 351 9291
rect 385 9257 386 9291
rect 350 9223 386 9257
rect 350 9189 351 9223
rect 385 9189 386 9223
rect 350 9155 386 9189
rect 350 9121 351 9155
rect 385 9121 386 9155
rect 350 9087 386 9121
rect 350 9053 351 9087
rect 385 9053 386 9087
rect 350 9019 386 9053
rect 350 8985 351 9019
rect 385 8985 386 9019
rect 350 8951 386 8985
rect 350 8917 351 8951
rect 385 8917 386 8951
rect 350 8883 386 8917
rect 350 8849 351 8883
rect 385 8849 386 8883
rect 350 8815 386 8849
rect 350 8781 351 8815
rect 385 8781 386 8815
rect 350 8747 386 8781
rect 350 8713 351 8747
rect 385 8713 386 8747
rect 350 8679 386 8713
rect 350 8645 351 8679
rect 385 8645 386 8679
rect 350 8611 386 8645
rect 350 8577 351 8611
rect 385 8577 386 8611
rect 350 8543 386 8577
rect 350 8509 351 8543
rect 385 8509 386 8543
rect 350 8475 386 8509
rect 350 8441 351 8475
rect 385 8441 386 8475
rect 350 8407 386 8441
rect 350 8373 351 8407
rect 385 8373 386 8407
rect 350 8339 386 8373
rect 350 8305 351 8339
rect 385 8305 386 8339
rect 350 8271 386 8305
rect 350 8237 351 8271
rect 385 8237 386 8271
rect 350 8203 386 8237
rect 350 8169 351 8203
rect 385 8169 386 8203
rect 350 8135 386 8169
rect 350 8101 351 8135
rect 385 8101 386 8135
rect 350 8067 386 8101
rect 350 8033 351 8067
rect 385 8033 386 8067
rect 350 7999 386 8033
rect 350 7965 351 7999
rect 385 7965 386 7999
rect 350 7931 386 7965
rect 350 7897 351 7931
rect 385 7897 386 7931
rect 350 7863 386 7897
rect 350 7829 351 7863
rect 385 7829 386 7863
rect 350 7795 386 7829
rect 350 7761 351 7795
rect 385 7761 386 7795
rect 350 7727 386 7761
rect 350 7693 351 7727
rect 385 7693 386 7727
rect 350 7659 386 7693
rect 350 7625 351 7659
rect 385 7625 386 7659
rect 350 7591 386 7625
rect 350 7557 351 7591
rect 385 7557 386 7591
rect 350 7523 386 7557
rect 350 7489 351 7523
rect 385 7489 386 7523
rect 350 7455 386 7489
rect 350 7421 351 7455
rect 385 7421 386 7455
rect 350 7387 386 7421
rect 350 7353 351 7387
rect 385 7353 386 7387
rect 350 7319 386 7353
rect 350 7285 351 7319
rect 385 7285 386 7319
rect 350 7251 386 7285
rect 350 7217 351 7251
rect 385 7217 386 7251
rect 350 7183 386 7217
rect 350 7149 351 7183
rect 385 7149 386 7183
rect 350 7115 386 7149
rect 350 7081 351 7115
rect 385 7081 386 7115
rect 350 7047 386 7081
rect 350 7013 351 7047
rect 385 7013 386 7047
rect 350 6979 386 7013
rect 350 6945 351 6979
rect 385 6945 386 6979
rect 350 6911 386 6945
rect 350 6877 351 6911
rect 385 6877 386 6911
rect 350 6843 386 6877
rect 350 6809 351 6843
rect 385 6809 386 6843
rect 350 6775 386 6809
rect 350 6741 351 6775
rect 385 6741 386 6775
rect 350 6707 386 6741
rect 350 6673 351 6707
rect 385 6673 386 6707
rect 350 6639 386 6673
rect 350 6605 351 6639
rect 385 6605 386 6639
rect 350 6571 386 6605
rect 350 6537 351 6571
rect 385 6537 386 6571
rect 350 6503 386 6537
rect 350 6469 351 6503
rect 385 6469 386 6503
rect 350 6435 386 6469
rect 350 6401 351 6435
rect 385 6401 386 6435
rect 350 6367 386 6401
rect 350 6333 351 6367
rect 385 6333 386 6367
rect 350 6299 386 6333
rect 350 6265 351 6299
rect 385 6265 386 6299
rect 350 6231 386 6265
rect 350 6197 351 6231
rect 385 6197 386 6231
rect 350 6163 386 6197
rect 350 6129 351 6163
rect 385 6129 386 6163
rect 350 6095 386 6129
rect 350 6061 351 6095
rect 385 6061 386 6095
rect 350 6027 386 6061
rect 350 5993 351 6027
rect 385 5993 386 6027
rect 350 5959 386 5993
rect 350 5925 351 5959
rect 385 5925 386 5959
rect 350 5891 386 5925
rect 350 5857 351 5891
rect 385 5857 386 5891
rect 350 5823 386 5857
rect 350 5789 351 5823
rect 385 5789 386 5823
rect 350 5755 386 5789
rect 350 5721 351 5755
rect 385 5721 386 5755
rect 350 5687 386 5721
rect 350 5653 351 5687
rect 385 5653 386 5687
rect 350 5619 386 5653
rect 350 5585 351 5619
rect 385 5585 386 5619
rect 350 5551 386 5585
rect 350 5517 351 5551
rect 385 5517 386 5551
rect 350 5483 386 5517
rect 350 5449 351 5483
rect 385 5449 386 5483
rect 350 5415 386 5449
rect 350 5381 351 5415
rect 385 5381 386 5415
rect 350 5347 386 5381
rect 350 5313 351 5347
rect 385 5313 386 5347
rect 350 5279 386 5313
rect 350 5245 351 5279
rect 385 5245 386 5279
rect 350 5211 386 5245
rect 350 5177 351 5211
rect 385 5177 386 5211
rect 350 5143 386 5177
rect 350 5109 351 5143
rect 385 5109 386 5143
rect 350 5075 386 5109
rect 350 5041 351 5075
rect 385 5041 386 5075
rect 350 5007 386 5041
rect 350 4973 351 5007
rect 385 4973 386 5007
rect 350 4939 386 4973
rect 350 4905 351 4939
rect 385 4905 386 4939
rect 350 4871 386 4905
rect 350 4837 351 4871
rect 385 4837 386 4871
rect 350 4803 386 4837
rect 350 4769 351 4803
rect 385 4769 386 4803
rect 350 4735 386 4769
rect 350 4701 351 4735
rect 385 4701 386 4735
rect 350 4667 386 4701
rect 350 4633 351 4667
rect 385 4633 386 4667
rect 350 4599 386 4633
rect 350 4565 351 4599
rect 385 4565 386 4599
rect 350 4531 386 4565
rect 350 4497 351 4531
rect 385 4497 386 4531
rect 350 4463 386 4497
rect 350 4429 351 4463
rect 385 4429 386 4463
rect 350 4395 386 4429
rect 350 4361 351 4395
rect 385 4361 386 4395
rect 350 4327 386 4361
rect 350 4293 351 4327
rect 385 4293 386 4327
rect 350 4259 386 4293
rect 350 4225 351 4259
rect 385 4225 386 4259
rect 350 4191 386 4225
rect 350 4157 351 4191
rect 385 4157 386 4191
rect 350 4123 386 4157
rect 350 4089 351 4123
rect 385 4089 386 4123
rect 350 4055 386 4089
rect 350 4021 351 4055
rect 385 4021 386 4055
rect 350 3987 386 4021
rect 350 3953 351 3987
rect 385 3953 386 3987
rect 350 3919 386 3953
rect 350 3885 351 3919
rect 385 3885 386 3919
rect 350 3851 386 3885
rect 350 3817 351 3851
rect 385 3817 386 3851
rect 350 3783 386 3817
rect 350 3749 351 3783
rect 385 3749 386 3783
rect 350 3715 386 3749
rect 350 3681 351 3715
rect 385 3681 386 3715
rect 350 3647 386 3681
rect 350 3613 351 3647
rect 385 3613 386 3647
rect 350 3579 386 3613
rect 350 3545 351 3579
rect 385 3545 386 3579
rect 350 3511 386 3545
rect 350 3477 351 3511
rect 385 3477 386 3511
rect 350 3443 386 3477
rect 350 3409 351 3443
rect 385 3409 386 3443
rect 350 3375 386 3409
rect 350 3341 351 3375
rect 385 3341 386 3375
rect 350 3307 386 3341
rect 350 3273 351 3307
rect 385 3273 386 3307
rect 350 3239 386 3273
rect 350 3205 351 3239
rect 385 3205 386 3239
rect 350 3171 386 3205
rect 350 3137 351 3171
rect 385 3137 386 3171
rect 350 3103 386 3137
rect 350 3069 351 3103
rect 385 3069 386 3103
rect 350 3035 386 3069
rect 350 3001 351 3035
rect 385 3001 386 3035
rect 350 2967 386 3001
rect 350 2933 351 2967
rect 385 2933 386 2967
rect 350 2899 386 2933
rect 350 2865 351 2899
rect 385 2865 386 2899
rect 350 2831 386 2865
rect 350 2797 351 2831
rect 385 2797 386 2831
rect 350 2763 386 2797
rect 350 2729 351 2763
rect 385 2729 386 2763
rect 350 2695 386 2729
rect 350 2661 351 2695
rect 385 2661 386 2695
rect 350 2627 386 2661
rect 350 2593 351 2627
rect 385 2593 386 2627
rect 350 2559 386 2593
rect 350 2525 351 2559
rect 385 2525 386 2559
rect 350 2491 386 2525
rect 350 2457 351 2491
rect 385 2457 386 2491
rect 350 2423 386 2457
rect 350 2389 351 2423
rect 385 2389 386 2423
rect 350 2355 386 2389
rect 350 2321 351 2355
rect 385 2321 386 2355
rect 350 2287 386 2321
rect 350 2253 351 2287
rect 385 2253 386 2287
rect 350 2219 386 2253
rect 350 2185 351 2219
rect 385 2185 386 2219
rect 350 2151 386 2185
rect 350 2117 351 2151
rect 385 2117 386 2151
rect 350 2083 386 2117
rect 350 2049 351 2083
rect 385 2049 386 2083
rect 350 2015 386 2049
rect 350 1981 351 2015
rect 385 1981 386 2015
rect 350 1947 386 1981
rect 350 1913 351 1947
rect 385 1913 386 1947
rect 350 1879 386 1913
rect 350 1845 351 1879
rect 385 1845 386 1879
rect 350 1811 386 1845
rect 350 1777 351 1811
rect 385 1777 386 1811
rect 350 1743 386 1777
rect 350 1709 351 1743
rect 385 1709 386 1743
rect 350 1675 386 1709
rect 350 1641 351 1675
rect 385 1641 386 1675
rect 350 1607 386 1641
rect 350 1573 351 1607
rect 385 1573 386 1607
rect 350 1539 386 1573
rect 350 1505 351 1539
rect 385 1505 386 1539
rect 350 1471 386 1505
rect 350 1437 351 1471
rect 385 1437 386 1471
rect 350 1403 386 1437
rect 350 1369 351 1403
rect 385 1369 386 1403
rect 350 1335 386 1369
rect 350 1301 351 1335
rect 385 1301 386 1335
rect 350 1267 386 1301
rect 350 1233 351 1267
rect 385 1233 386 1267
rect 350 1199 386 1233
rect 350 1165 351 1199
rect 385 1165 386 1199
rect 350 1131 386 1165
rect 350 1097 351 1131
rect 385 1097 386 1131
rect 350 1063 386 1097
rect 350 1029 351 1063
rect 385 1029 386 1063
rect 350 995 386 1029
rect 350 961 351 995
rect 385 961 386 995
rect 350 927 386 961
rect 350 893 351 927
rect 385 893 386 927
rect 350 859 386 893
rect 350 825 351 859
rect 385 825 386 859
rect 350 791 386 825
rect 350 757 351 791
rect 385 757 386 791
rect 350 723 386 757
rect 350 689 351 723
rect 385 689 386 723
rect 350 655 386 689
rect 350 621 351 655
rect 385 621 386 655
rect 350 587 386 621
rect 350 553 351 587
rect 385 553 386 587
rect 539 9544 5865 9545
rect 539 9511 546 9544
rect 539 9477 540 9511
rect 580 9510 618 9544
rect 666 9510 690 9544
rect 734 9510 762 9544
rect 802 9510 834 9544
rect 870 9510 904 9544
rect 940 9510 972 9544
rect 1012 9510 1040 9544
rect 1074 9510 1108 9544
rect 1142 9510 1176 9544
rect 1210 9510 1244 9544
rect 1278 9510 1312 9544
rect 1346 9510 1380 9544
rect 1414 9510 1448 9544
rect 1482 9510 1516 9544
rect 1550 9510 1584 9544
rect 1618 9510 1652 9544
rect 1686 9510 1720 9544
rect 1754 9510 1788 9544
rect 1822 9510 1856 9544
rect 1890 9510 1924 9544
rect 1958 9510 1992 9544
rect 2026 9510 2060 9544
rect 2094 9510 2128 9544
rect 2162 9510 2196 9544
rect 2230 9510 2264 9544
rect 2298 9510 2332 9544
rect 2366 9510 2400 9544
rect 2434 9510 2468 9544
rect 2502 9510 2576 9544
rect 2610 9510 2644 9544
rect 2678 9510 2712 9544
rect 2746 9510 2780 9544
rect 2814 9510 2848 9544
rect 2882 9510 2916 9544
rect 2950 9510 2984 9544
rect 3018 9510 3052 9544
rect 3086 9510 3120 9544
rect 3154 9510 3188 9544
rect 3222 9510 3256 9544
rect 3290 9510 3324 9544
rect 3358 9510 3426 9544
rect 3460 9510 3494 9544
rect 3528 9510 3562 9544
rect 3596 9510 3630 9544
rect 3664 9510 3698 9544
rect 3732 9510 3766 9544
rect 3800 9510 3834 9544
rect 3868 9510 3902 9544
rect 3936 9510 3970 9544
rect 4004 9510 4036 9544
rect 4072 9510 4106 9544
rect 4142 9510 4174 9544
rect 4214 9510 4242 9544
rect 4286 9510 4310 9544
rect 4358 9510 4378 9544
rect 4430 9510 4446 9544
rect 4502 9510 4514 9544
rect 4548 9510 4582 9544
rect 4616 9510 4650 9544
rect 4692 9510 4718 9544
rect 4764 9510 4786 9544
rect 4836 9510 4854 9544
rect 4908 9510 4922 9544
rect 4980 9510 4990 9544
rect 5024 9510 5058 9544
rect 5092 9510 5113 9544
rect 5160 9510 5185 9544
rect 5228 9510 5257 9544
rect 5296 9510 5329 9544
rect 5364 9510 5398 9544
rect 5435 9510 5466 9544
rect 5500 9510 5534 9544
rect 5568 9510 5602 9544
rect 5642 9510 5670 9544
rect 5714 9510 5738 9544
rect 5786 9510 5824 9544
rect 5858 9510 5865 9544
rect 574 9509 5865 9510
rect 574 9477 575 9509
rect 539 9443 575 9477
rect 539 9409 540 9443
rect 574 9409 575 9443
rect 539 9375 575 9409
rect 539 9341 540 9375
rect 574 9341 575 9375
rect 539 9307 575 9341
rect 539 9273 540 9307
rect 574 9273 575 9307
rect 539 9239 575 9273
rect 539 9205 540 9239
rect 574 9205 575 9239
rect 539 9171 575 9205
rect 539 9137 540 9171
rect 574 9137 575 9171
rect 539 9103 575 9137
rect 539 9069 540 9103
rect 574 9069 575 9103
rect 539 9035 575 9069
rect 539 9001 540 9035
rect 574 9001 575 9035
rect 539 8967 575 9001
rect 539 8933 540 8967
rect 574 8933 575 8967
rect 539 8899 575 8933
rect 539 8865 540 8899
rect 574 8865 575 8899
rect 539 8831 575 8865
rect 539 8797 540 8831
rect 574 8797 575 8831
rect 539 8763 575 8797
rect 539 8729 540 8763
rect 574 8729 575 8763
rect 539 8695 575 8729
rect 539 8661 540 8695
rect 574 8661 575 8695
rect 539 8627 575 8661
rect 539 8593 540 8627
rect 574 8593 575 8627
rect 539 8559 575 8593
rect 539 8525 540 8559
rect 574 8525 575 8559
rect 539 8491 575 8525
rect 539 8457 540 8491
rect 574 8457 575 8491
rect 539 8423 575 8457
rect 539 8389 540 8423
rect 574 8389 575 8423
rect 539 8355 575 8389
rect 539 8321 540 8355
rect 574 8321 575 8355
rect 539 8287 575 8321
rect 539 8253 540 8287
rect 574 8253 575 8287
rect 539 8219 575 8253
rect 539 8185 540 8219
rect 574 8185 575 8219
rect 539 8151 575 8185
rect 539 8117 540 8151
rect 574 8117 575 8151
rect 539 8083 575 8117
rect 539 8049 540 8083
rect 574 8049 575 8083
rect 539 8015 575 8049
rect 539 7981 540 8015
rect 574 7981 575 8015
rect 539 7947 575 7981
rect 539 7913 540 7947
rect 574 7913 575 7947
rect 539 7879 575 7913
rect 539 7845 540 7879
rect 574 7845 575 7879
rect 539 7811 575 7845
rect 539 7777 540 7811
rect 574 7777 575 7811
rect 539 7743 575 7777
rect 539 7709 540 7743
rect 574 7709 575 7743
rect 539 7675 575 7709
rect 539 7641 540 7675
rect 574 7641 575 7675
rect 539 7607 575 7641
rect 539 7573 540 7607
rect 574 7573 575 7607
rect 539 7539 575 7573
rect 539 7505 540 7539
rect 574 7505 575 7539
rect 539 7471 575 7505
rect 539 7437 540 7471
rect 574 7437 575 7471
rect 539 7403 575 7437
rect 539 7369 540 7403
rect 574 7369 575 7403
rect 539 7288 575 7369
rect 3356 9396 3392 9509
rect 5829 9475 5865 9509
rect 4421 9425 4437 9459
rect 4471 9425 4501 9459
rect 4539 9425 4573 9459
rect 4607 9425 4641 9459
rect 4679 9425 4709 9459
rect 4743 9425 4759 9459
rect 4877 9425 4893 9459
rect 4927 9425 4957 9459
rect 4995 9425 5029 9459
rect 5063 9425 5097 9459
rect 5135 9425 5165 9459
rect 5199 9425 5215 9459
rect 5333 9425 5349 9459
rect 5383 9425 5413 9459
rect 5451 9425 5485 9459
rect 5519 9425 5553 9459
rect 5591 9425 5621 9459
rect 5655 9425 5671 9459
rect 5829 9441 5830 9475
rect 5864 9441 5865 9475
rect 3356 9362 3357 9396
rect 3391 9362 3392 9396
rect 3356 9328 3392 9362
rect 3356 9294 3357 9328
rect 3391 9294 3392 9328
rect 3356 9260 3392 9294
rect 3356 9226 3357 9260
rect 3391 9226 3392 9260
rect 3356 9192 3392 9226
rect 3356 9158 3357 9192
rect 3391 9158 3392 9192
rect 3356 9124 3392 9158
rect 3356 9090 3357 9124
rect 3391 9090 3392 9124
rect 3356 9056 3392 9090
rect 3356 9022 3357 9056
rect 3391 9022 3392 9056
rect 3356 8988 3392 9022
rect 3356 8954 3357 8988
rect 3391 8954 3392 8988
rect 3356 8920 3392 8954
rect 3356 8886 3357 8920
rect 3391 8886 3392 8920
rect 3356 8852 3392 8886
rect 3356 8818 3357 8852
rect 3391 8818 3392 8852
rect 3356 8784 3392 8818
rect 3356 8750 3357 8784
rect 3391 8750 3392 8784
rect 3356 8716 3392 8750
rect 3356 8682 3357 8716
rect 3391 8682 3392 8716
rect 3356 8648 3392 8682
rect 3356 8614 3357 8648
rect 3391 8614 3392 8648
rect 3356 8580 3392 8614
rect 3356 8546 3357 8580
rect 3391 8546 3392 8580
rect 3356 8512 3392 8546
rect 3356 8478 3357 8512
rect 3391 8478 3392 8512
rect 3356 8444 3392 8478
rect 3356 8410 3357 8444
rect 3391 8410 3392 8444
rect 3356 8376 3392 8410
rect 3356 8342 3357 8376
rect 3391 8342 3392 8376
rect 3356 8308 3392 8342
rect 3356 8274 3357 8308
rect 3391 8274 3392 8308
rect 3356 8240 3392 8274
rect 3356 8206 3357 8240
rect 3391 8206 3392 8240
rect 3356 8172 3392 8206
rect 3356 8138 3357 8172
rect 3391 8138 3392 8172
rect 3356 8104 3392 8138
rect 3356 8070 3357 8104
rect 3391 8070 3392 8104
rect 3356 8036 3392 8070
rect 3356 8002 3357 8036
rect 3391 8002 3392 8036
rect 3356 7968 3392 8002
rect 3356 7934 3357 7968
rect 3391 7934 3392 7968
rect 3356 7900 3392 7934
rect 3356 7866 3357 7900
rect 3391 7866 3392 7900
rect 3356 7832 3392 7866
rect 3356 7798 3357 7832
rect 3391 7798 3392 7832
rect 3356 7764 3392 7798
rect 3356 7730 3357 7764
rect 3391 7730 3392 7764
rect 3356 7696 3392 7730
rect 3356 7662 3357 7696
rect 3391 7662 3392 7696
rect 3356 7628 3392 7662
rect 3356 7594 3357 7628
rect 3391 7594 3392 7628
rect 3356 7560 3392 7594
rect 3356 7526 3357 7560
rect 3391 7526 3392 7560
rect 3356 7492 3392 7526
rect 3356 7458 3357 7492
rect 3391 7458 3392 7492
rect 3356 7424 3392 7458
rect 3356 7390 3357 7424
rect 3391 7390 3392 7424
rect 3356 7356 3392 7390
rect 3356 7322 3357 7356
rect 3391 7322 3392 7356
rect 3356 7288 3392 7322
rect 5829 9407 5865 9441
rect 5829 9373 5830 9407
rect 5864 9373 5865 9407
rect 5829 9339 5865 9373
rect 5829 9305 5830 9339
rect 5864 9305 5865 9339
rect 5829 9271 5865 9305
rect 5829 9237 5830 9271
rect 5864 9237 5865 9271
rect 5829 9203 5865 9237
rect 5829 9169 5830 9203
rect 5864 9169 5865 9203
rect 5829 9135 5865 9169
rect 5829 9101 5830 9135
rect 5864 9101 5865 9135
rect 5829 9067 5865 9101
rect 5829 9033 5830 9067
rect 5864 9033 5865 9067
rect 5829 8999 5865 9033
rect 5829 8965 5830 8999
rect 5864 8965 5865 8999
rect 5829 8931 5865 8965
rect 5829 8897 5830 8931
rect 5864 8897 5865 8931
rect 5829 8863 5865 8897
rect 5829 8829 5830 8863
rect 5864 8829 5865 8863
rect 5829 8795 5865 8829
rect 5829 8761 5830 8795
rect 5864 8761 5865 8795
rect 5829 8727 5865 8761
rect 5829 8693 5830 8727
rect 5864 8693 5865 8727
rect 5829 8659 5865 8693
rect 5829 8625 5830 8659
rect 5864 8625 5865 8659
rect 5829 8591 5865 8625
rect 5829 8557 5830 8591
rect 5864 8557 5865 8591
rect 5829 8523 5865 8557
rect 5829 8489 5830 8523
rect 5864 8489 5865 8523
rect 5829 8455 5865 8489
rect 5829 8421 5830 8455
rect 5864 8421 5865 8455
rect 5829 8387 5865 8421
rect 5829 8353 5830 8387
rect 5864 8353 5865 8387
rect 5829 8319 5865 8353
rect 5829 8285 5830 8319
rect 5864 8285 5865 8319
rect 5829 8251 5865 8285
rect 5829 8217 5830 8251
rect 5864 8217 5865 8251
rect 5829 8183 5865 8217
rect 5829 8149 5830 8183
rect 5864 8149 5865 8183
rect 5829 8115 5865 8149
rect 5829 8081 5830 8115
rect 5864 8081 5865 8115
rect 5829 8047 5865 8081
rect 5829 8013 5830 8047
rect 5864 8013 5865 8047
rect 5829 7979 5865 8013
rect 5829 7945 5830 7979
rect 5864 7945 5865 7979
rect 5829 7911 5865 7945
rect 5829 7877 5830 7911
rect 5864 7877 5865 7911
rect 5829 7843 5865 7877
rect 5829 7809 5830 7843
rect 5864 7809 5865 7843
rect 5829 7775 5865 7809
rect 5829 7741 5830 7775
rect 5864 7741 5865 7775
rect 5829 7707 5865 7741
rect 5829 7673 5830 7707
rect 5864 7673 5865 7707
rect 5829 7639 5865 7673
rect 5829 7605 5830 7639
rect 5864 7605 5865 7639
rect 5829 7571 5865 7605
rect 5829 7537 5830 7571
rect 5864 7537 5865 7571
rect 5829 7503 5865 7537
rect 5829 7469 5830 7503
rect 5864 7469 5865 7503
rect 5829 7435 5865 7469
rect 5829 7401 5830 7435
rect 5864 7401 5865 7435
rect 5829 7367 5865 7401
rect 5829 7333 5830 7367
rect 5864 7333 5865 7367
rect 5829 7299 5865 7333
rect 5829 7288 5830 7299
rect 539 7287 967 7288
rect 539 7253 657 7287
rect 691 7253 729 7287
rect 775 7253 801 7287
rect 859 7253 873 7287
rect 907 7253 909 7287
rect 943 7253 967 7287
rect 1237 7287 1823 7288
rect 539 7252 967 7253
rect 1001 7252 1017 7286
rect 1083 7252 1085 7286
rect 1119 7252 1121 7286
rect 1187 7252 1203 7286
rect 1237 7253 1261 7287
rect 1295 7253 1297 7287
rect 1331 7253 1345 7287
rect 1403 7253 1429 7287
rect 1475 7253 1513 7287
rect 1547 7253 1585 7287
rect 1631 7253 1657 7287
rect 1715 7253 1729 7287
rect 1763 7253 1765 7287
rect 1799 7253 1823 7287
rect 2093 7287 2679 7288
rect 1237 7252 1823 7253
rect 1857 7252 1873 7286
rect 1939 7252 1941 7286
rect 1975 7252 1977 7286
rect 2043 7252 2059 7286
rect 2093 7253 2117 7287
rect 2151 7253 2153 7287
rect 2187 7253 2201 7287
rect 2259 7253 2285 7287
rect 2331 7253 2369 7287
rect 2403 7253 2441 7287
rect 2487 7253 2513 7287
rect 2571 7253 2585 7287
rect 2619 7253 2621 7287
rect 2655 7253 2679 7287
rect 2949 7287 3357 7288
rect 2093 7252 2679 7253
rect 2713 7252 2729 7286
rect 2795 7252 2797 7286
rect 2831 7252 2833 7286
rect 2899 7252 2915 7286
rect 2949 7253 2973 7287
rect 3007 7253 3009 7287
rect 3043 7253 3057 7287
rect 3115 7253 3141 7287
rect 3187 7253 3225 7287
rect 3259 7254 3357 7287
rect 3391 7287 3799 7288
rect 3391 7254 3489 7287
rect 3259 7253 3489 7254
rect 3523 7253 3561 7287
rect 3607 7253 3633 7287
rect 3691 7253 3705 7287
rect 3739 7253 3741 7287
rect 3775 7253 3799 7287
rect 4069 7287 4455 7288
rect 2949 7252 3799 7253
rect 3833 7252 3849 7286
rect 3915 7252 3917 7286
rect 3951 7252 3953 7286
rect 4019 7252 4035 7286
rect 4069 7253 4093 7287
rect 4127 7253 4129 7287
rect 4163 7253 4177 7287
rect 4235 7253 4261 7287
rect 4307 7253 4345 7287
rect 4379 7253 4455 7287
rect 4725 7287 4911 7288
rect 4069 7252 4455 7253
rect 4489 7252 4505 7286
rect 4571 7252 4573 7286
rect 4607 7252 4609 7286
rect 4675 7252 4691 7286
rect 4725 7253 4765 7287
rect 4799 7253 4801 7287
rect 4835 7253 4837 7287
rect 4871 7253 4911 7287
rect 5181 7287 5367 7288
rect 4725 7252 4911 7253
rect 4945 7252 4961 7286
rect 5027 7252 5029 7286
rect 5063 7252 5065 7286
rect 5131 7252 5147 7286
rect 5181 7253 5221 7287
rect 5255 7253 5257 7287
rect 5291 7253 5293 7287
rect 5327 7253 5367 7287
rect 5637 7287 5830 7288
rect 5181 7252 5367 7253
rect 5401 7252 5417 7286
rect 5483 7252 5485 7286
rect 5519 7252 5521 7286
rect 5587 7252 5603 7286
rect 5637 7253 5713 7287
rect 5747 7265 5830 7287
rect 5864 7265 5865 7299
rect 5747 7253 5865 7265
rect 5637 7252 5865 7253
rect 539 7251 575 7252
rect 539 7217 540 7251
rect 574 7217 575 7251
rect 539 7183 575 7217
rect 539 7149 540 7183
rect 574 7149 575 7183
rect 539 7115 575 7149
rect 539 7081 540 7115
rect 574 7081 575 7115
rect 539 7047 575 7081
rect 539 7013 540 7047
rect 574 7013 575 7047
rect 539 6979 575 7013
rect 539 6945 540 6979
rect 574 6945 575 6979
rect 539 6911 575 6945
rect 539 6877 540 6911
rect 574 6877 575 6911
rect 539 6843 575 6877
rect 539 6809 540 6843
rect 574 6809 575 6843
rect 539 6775 575 6809
rect 539 6741 540 6775
rect 574 6741 575 6775
rect 539 6707 575 6741
rect 539 6673 540 6707
rect 574 6673 575 6707
rect 539 6639 575 6673
rect 539 6605 540 6639
rect 574 6605 575 6639
rect 539 6571 575 6605
rect 539 6537 540 6571
rect 574 6537 575 6571
rect 539 6503 575 6537
rect 539 6469 540 6503
rect 574 6469 575 6503
rect 539 6435 575 6469
rect 539 6401 540 6435
rect 574 6401 575 6435
rect 539 6367 575 6401
rect 539 6333 540 6367
rect 574 6333 575 6367
rect 539 6299 575 6333
rect 539 6265 540 6299
rect 574 6265 575 6299
rect 539 6231 575 6265
rect 539 6197 540 6231
rect 574 6197 575 6231
rect 539 6163 575 6197
rect 539 6129 540 6163
rect 574 6129 575 6163
rect 539 6095 575 6129
rect 539 6061 540 6095
rect 574 6061 575 6095
rect 539 6027 575 6061
rect 539 5993 540 6027
rect 574 5993 575 6027
rect 539 5959 575 5993
rect 539 5925 540 5959
rect 574 5925 575 5959
rect 539 5891 575 5925
rect 539 5857 540 5891
rect 574 5857 575 5891
rect 539 5823 575 5857
rect 539 5789 540 5823
rect 574 5789 575 5823
rect 539 5755 575 5789
rect 539 5721 540 5755
rect 574 5721 575 5755
rect 539 5687 575 5721
rect 539 5653 540 5687
rect 574 5653 575 5687
rect 539 5619 575 5653
rect 539 5585 540 5619
rect 574 5585 575 5619
rect 539 5551 575 5585
rect 539 5517 540 5551
rect 574 5517 575 5551
rect 539 5483 575 5517
rect 539 5449 540 5483
rect 574 5449 575 5483
rect 539 5415 575 5449
rect 539 5381 540 5415
rect 574 5381 575 5415
rect 539 5347 575 5381
rect 539 5313 540 5347
rect 574 5313 575 5347
rect 539 5279 575 5313
rect 539 5245 540 5279
rect 574 5245 575 5279
rect 539 5211 575 5245
rect 539 5177 540 5211
rect 574 5177 575 5211
rect 539 5068 575 5177
rect 3356 7220 3392 7252
rect 3356 7186 3357 7220
rect 3391 7186 3392 7220
rect 3356 7152 3392 7186
rect 3356 7118 3357 7152
rect 3391 7118 3392 7152
rect 3356 7084 3392 7118
rect 3356 7050 3357 7084
rect 3391 7050 3392 7084
rect 3356 7016 3392 7050
rect 3356 6982 3357 7016
rect 3391 6982 3392 7016
rect 3356 6948 3392 6982
rect 3356 6914 3357 6948
rect 3391 6914 3392 6948
rect 3356 6880 3392 6914
rect 3356 6846 3357 6880
rect 3391 6846 3392 6880
rect 3356 6812 3392 6846
rect 3356 6778 3357 6812
rect 3391 6778 3392 6812
rect 3356 6744 3392 6778
rect 3356 6710 3357 6744
rect 3391 6710 3392 6744
rect 3356 6676 3392 6710
rect 3356 6642 3357 6676
rect 3391 6642 3392 6676
rect 3356 6608 3392 6642
rect 3356 6574 3357 6608
rect 3391 6574 3392 6608
rect 3356 6540 3392 6574
rect 3356 6506 3357 6540
rect 3391 6506 3392 6540
rect 3356 6472 3392 6506
rect 3356 6438 3357 6472
rect 3391 6438 3392 6472
rect 3356 6404 3392 6438
rect 3356 6370 3357 6404
rect 3391 6370 3392 6404
rect 3356 6336 3392 6370
rect 3356 6302 3357 6336
rect 3391 6302 3392 6336
rect 3356 6268 3392 6302
rect 3356 6234 3357 6268
rect 3391 6234 3392 6268
rect 3356 6200 3392 6234
rect 3356 6166 3357 6200
rect 3391 6166 3392 6200
rect 3356 6132 3392 6166
rect 3356 6098 3357 6132
rect 3391 6098 3392 6132
rect 3356 6064 3392 6098
rect 3356 6030 3357 6064
rect 3391 6030 3392 6064
rect 3356 5996 3392 6030
rect 3356 5962 3357 5996
rect 3391 5962 3392 5996
rect 3356 5928 3392 5962
rect 3356 5894 3357 5928
rect 3391 5894 3392 5928
rect 3356 5860 3392 5894
rect 3356 5826 3357 5860
rect 3391 5826 3392 5860
rect 3356 5792 3392 5826
rect 3356 5758 3357 5792
rect 3391 5758 3392 5792
rect 3356 5724 3392 5758
rect 3356 5690 3357 5724
rect 3391 5690 3392 5724
rect 3356 5656 3392 5690
rect 3356 5622 3357 5656
rect 3391 5622 3392 5656
rect 3356 5588 3392 5622
rect 3356 5554 3357 5588
rect 3391 5554 3392 5588
rect 3356 5520 3392 5554
rect 3356 5486 3357 5520
rect 3391 5486 3392 5520
rect 3356 5452 3392 5486
rect 3356 5418 3357 5452
rect 3391 5418 3392 5452
rect 3356 5384 3392 5418
rect 3356 5350 3357 5384
rect 3391 5350 3392 5384
rect 3356 5316 3392 5350
rect 3356 5282 3357 5316
rect 3391 5282 3392 5316
rect 3356 5248 3392 5282
rect 3356 5214 3357 5248
rect 3391 5214 3392 5248
rect 3356 5180 3392 5214
rect 3356 5146 3357 5180
rect 3391 5146 3392 5180
rect 3356 5112 3392 5146
rect 3356 5078 3357 5112
rect 3391 5078 3392 5112
rect 3356 5068 3392 5078
rect 5829 7231 5865 7252
rect 5829 7197 5830 7231
rect 5864 7197 5865 7231
rect 5829 7163 5865 7197
rect 5829 7129 5830 7163
rect 5864 7129 5865 7163
rect 5829 7095 5865 7129
rect 5829 7061 5830 7095
rect 5864 7061 5865 7095
rect 5829 7027 5865 7061
rect 5829 6993 5830 7027
rect 5864 6993 5865 7027
rect 5829 6959 5865 6993
rect 5829 6925 5830 6959
rect 5864 6925 5865 6959
rect 5829 6891 5865 6925
rect 5829 6857 5830 6891
rect 5864 6857 5865 6891
rect 5829 6823 5865 6857
rect 5829 6789 5830 6823
rect 5864 6789 5865 6823
rect 5829 6755 5865 6789
rect 5829 6721 5830 6755
rect 5864 6721 5865 6755
rect 5829 6687 5865 6721
rect 5829 6653 5830 6687
rect 5864 6653 5865 6687
rect 5829 6619 5865 6653
rect 5829 6585 5830 6619
rect 5864 6585 5865 6619
rect 5829 6551 5865 6585
rect 5829 6517 5830 6551
rect 5864 6517 5865 6551
rect 5829 6483 5865 6517
rect 5829 6449 5830 6483
rect 5864 6449 5865 6483
rect 5829 6415 5865 6449
rect 5829 6381 5830 6415
rect 5864 6381 5865 6415
rect 5829 6347 5865 6381
rect 5829 6313 5830 6347
rect 5864 6313 5865 6347
rect 5829 6279 5865 6313
rect 5829 6245 5830 6279
rect 5864 6245 5865 6279
rect 5829 6211 5865 6245
rect 5829 6177 5830 6211
rect 5864 6177 5865 6211
rect 5829 6143 5865 6177
rect 5829 6109 5830 6143
rect 5864 6109 5865 6143
rect 5829 6075 5865 6109
rect 5829 6041 5830 6075
rect 5864 6041 5865 6075
rect 5829 6007 5865 6041
rect 5829 5973 5830 6007
rect 5864 5973 5865 6007
rect 5829 5939 5865 5973
rect 5829 5905 5830 5939
rect 5864 5905 5865 5939
rect 5829 5871 5865 5905
rect 5829 5837 5830 5871
rect 5864 5837 5865 5871
rect 5829 5803 5865 5837
rect 5829 5769 5830 5803
rect 5864 5769 5865 5803
rect 5829 5735 5865 5769
rect 5829 5701 5830 5735
rect 5864 5701 5865 5735
rect 5829 5667 5865 5701
rect 5829 5633 5830 5667
rect 5864 5633 5865 5667
rect 5829 5599 5865 5633
rect 5829 5565 5830 5599
rect 5864 5565 5865 5599
rect 5829 5531 5865 5565
rect 5829 5497 5830 5531
rect 5864 5497 5865 5531
rect 5829 5463 5865 5497
rect 5829 5429 5830 5463
rect 5864 5429 5865 5463
rect 5829 5395 5865 5429
rect 5829 5361 5830 5395
rect 5864 5361 5865 5395
rect 5829 5327 5865 5361
rect 5829 5293 5830 5327
rect 5864 5293 5865 5327
rect 5829 5259 5865 5293
rect 5829 5225 5830 5259
rect 5864 5225 5865 5259
rect 5829 5191 5865 5225
rect 5829 5157 5830 5191
rect 5864 5157 5865 5191
rect 5829 5123 5865 5157
rect 5829 5089 5830 5123
rect 5864 5089 5865 5123
rect 5829 5068 5865 5089
rect 539 5067 967 5068
rect 539 5048 657 5067
rect 539 5014 540 5048
rect 574 5033 657 5048
rect 691 5033 729 5067
rect 775 5033 801 5067
rect 859 5033 873 5067
rect 907 5033 909 5067
rect 943 5033 967 5067
rect 1237 5067 1823 5068
rect 574 5032 967 5033
rect 1001 5032 1017 5066
rect 1083 5032 1085 5066
rect 1119 5032 1121 5066
rect 1187 5032 1203 5066
rect 1237 5033 1261 5067
rect 1295 5033 1297 5067
rect 1331 5033 1345 5067
rect 1403 5033 1429 5067
rect 1475 5033 1513 5067
rect 1547 5033 1585 5067
rect 1631 5033 1657 5067
rect 1715 5033 1729 5067
rect 1763 5033 1765 5067
rect 1799 5033 1823 5067
rect 2093 5067 2679 5068
rect 1237 5032 1823 5033
rect 1857 5032 1873 5066
rect 1939 5032 1941 5066
rect 1975 5032 1977 5066
rect 2043 5032 2059 5066
rect 2093 5033 2117 5067
rect 2151 5033 2153 5067
rect 2187 5033 2201 5067
rect 2259 5033 2285 5067
rect 2331 5033 2369 5067
rect 2403 5033 2441 5067
rect 2487 5033 2513 5067
rect 2571 5033 2585 5067
rect 2619 5033 2621 5067
rect 2655 5033 2679 5067
rect 2949 5067 3799 5068
rect 2093 5032 2679 5033
rect 2713 5032 2729 5066
rect 2795 5032 2797 5066
rect 2831 5032 2833 5066
rect 2899 5032 2915 5066
rect 2949 5033 2973 5067
rect 3007 5033 3009 5067
rect 3043 5033 3057 5067
rect 3115 5033 3141 5067
rect 3187 5033 3225 5067
rect 3259 5044 3489 5067
rect 3259 5033 3357 5044
rect 2949 5032 3357 5033
rect 574 5014 575 5032
rect 539 4980 575 5014
rect 539 4946 540 4980
rect 574 4946 575 4980
rect 539 4912 575 4946
rect 539 4878 540 4912
rect 574 4878 575 4912
rect 539 4844 575 4878
rect 539 4810 540 4844
rect 574 4810 575 4844
rect 539 4776 575 4810
rect 539 4742 540 4776
rect 574 4742 575 4776
rect 539 4708 575 4742
rect 539 4674 540 4708
rect 574 4674 575 4708
rect 539 4640 575 4674
rect 539 4606 540 4640
rect 574 4606 575 4640
rect 539 4572 575 4606
rect 539 4538 540 4572
rect 574 4538 575 4572
rect 539 4504 575 4538
rect 539 4470 540 4504
rect 574 4470 575 4504
rect 539 4436 575 4470
rect 539 4402 540 4436
rect 574 4402 575 4436
rect 539 4368 575 4402
rect 539 4334 540 4368
rect 574 4334 575 4368
rect 539 4300 575 4334
rect 539 4266 540 4300
rect 574 4266 575 4300
rect 539 4232 575 4266
rect 539 4198 540 4232
rect 574 4198 575 4232
rect 539 4164 575 4198
rect 539 4130 540 4164
rect 574 4130 575 4164
rect 539 4096 575 4130
rect 539 4062 540 4096
rect 574 4062 575 4096
rect 539 4028 575 4062
rect 539 3994 540 4028
rect 574 3994 575 4028
rect 539 3960 575 3994
rect 539 3926 540 3960
rect 574 3926 575 3960
rect 539 3892 575 3926
rect 539 3858 540 3892
rect 574 3858 575 3892
rect 539 3824 575 3858
rect 539 3790 540 3824
rect 574 3790 575 3824
rect 539 3756 575 3790
rect 539 3722 540 3756
rect 574 3722 575 3756
rect 539 3688 575 3722
rect 539 3654 540 3688
rect 574 3654 575 3688
rect 539 3620 575 3654
rect 539 3586 540 3620
rect 574 3586 575 3620
rect 539 3552 575 3586
rect 539 3518 540 3552
rect 574 3518 575 3552
rect 539 3484 575 3518
rect 539 3450 540 3484
rect 574 3450 575 3484
rect 539 3416 575 3450
rect 539 3382 540 3416
rect 574 3382 575 3416
rect 539 3348 575 3382
rect 539 3314 540 3348
rect 574 3314 575 3348
rect 539 3280 575 3314
rect 539 3246 540 3280
rect 574 3246 575 3280
rect 539 3212 575 3246
rect 539 3178 540 3212
rect 574 3178 575 3212
rect 539 3144 575 3178
rect 539 3110 540 3144
rect 574 3110 575 3144
rect 539 3076 575 3110
rect 539 3042 540 3076
rect 574 3042 575 3076
rect 539 3008 575 3042
rect 539 2974 540 3008
rect 574 2974 575 3008
rect 539 2940 575 2974
rect 539 2906 540 2940
rect 574 2906 575 2940
rect 539 2872 575 2906
rect 539 2838 540 2872
rect 574 2849 575 2872
rect 3356 5010 3357 5032
rect 3391 5033 3489 5044
rect 3523 5033 3561 5067
rect 3607 5033 3633 5067
rect 3691 5033 3705 5067
rect 3739 5033 3741 5067
rect 3775 5033 3799 5067
rect 4069 5067 4455 5068
rect 3391 5032 3799 5033
rect 3833 5032 3849 5066
rect 3915 5032 3917 5066
rect 3951 5032 3953 5066
rect 4019 5032 4035 5066
rect 4069 5033 4093 5067
rect 4127 5033 4129 5067
rect 4163 5033 4177 5067
rect 4235 5033 4261 5067
rect 4307 5033 4345 5067
rect 4379 5033 4455 5067
rect 4725 5067 4911 5068
rect 4069 5032 4455 5033
rect 4489 5032 4505 5066
rect 4571 5032 4573 5066
rect 4607 5032 4609 5066
rect 4675 5032 4691 5066
rect 4725 5033 4765 5067
rect 4799 5033 4801 5067
rect 4835 5033 4837 5067
rect 4871 5033 4911 5067
rect 5181 5067 5367 5068
rect 4725 5032 4911 5033
rect 4945 5032 4961 5066
rect 5027 5032 5029 5066
rect 5063 5032 5065 5066
rect 5131 5032 5147 5066
rect 5181 5033 5221 5067
rect 5255 5033 5257 5067
rect 5291 5033 5293 5067
rect 5327 5033 5367 5067
rect 5637 5067 5865 5068
rect 5181 5032 5367 5033
rect 5401 5032 5417 5066
rect 5483 5032 5485 5066
rect 5519 5032 5521 5066
rect 5587 5032 5603 5066
rect 5637 5033 5713 5067
rect 5747 5055 5865 5067
rect 5747 5033 5830 5055
rect 5637 5032 5830 5033
rect 3391 5010 3392 5032
rect 3356 4976 3392 5010
rect 3356 4942 3357 4976
rect 3391 4942 3392 4976
rect 3356 4908 3392 4942
rect 3356 4874 3357 4908
rect 3391 4874 3392 4908
rect 3356 4840 3392 4874
rect 3356 4806 3357 4840
rect 3391 4806 3392 4840
rect 3356 4772 3392 4806
rect 3356 4738 3357 4772
rect 3391 4738 3392 4772
rect 3356 4704 3392 4738
rect 3356 4670 3357 4704
rect 3391 4670 3392 4704
rect 3356 4636 3392 4670
rect 3356 4602 3357 4636
rect 3391 4602 3392 4636
rect 3356 4568 3392 4602
rect 3356 4534 3357 4568
rect 3391 4534 3392 4568
rect 3356 4500 3392 4534
rect 3356 4466 3357 4500
rect 3391 4466 3392 4500
rect 3356 4432 3392 4466
rect 3356 4398 3357 4432
rect 3391 4398 3392 4432
rect 3356 4364 3392 4398
rect 3356 4330 3357 4364
rect 3391 4330 3392 4364
rect 3356 4296 3392 4330
rect 3356 4262 3357 4296
rect 3391 4262 3392 4296
rect 3356 4228 3392 4262
rect 3356 4194 3357 4228
rect 3391 4194 3392 4228
rect 3356 4160 3392 4194
rect 3356 4126 3357 4160
rect 3391 4126 3392 4160
rect 3356 4092 3392 4126
rect 3356 4058 3357 4092
rect 3391 4058 3392 4092
rect 3356 4024 3392 4058
rect 3356 3990 3357 4024
rect 3391 3990 3392 4024
rect 3356 3956 3392 3990
rect 3356 3922 3357 3956
rect 3391 3922 3392 3956
rect 3356 3888 3392 3922
rect 3356 3854 3357 3888
rect 3391 3854 3392 3888
rect 3356 3820 3392 3854
rect 3356 3786 3357 3820
rect 3391 3786 3392 3820
rect 3356 3752 3392 3786
rect 3356 3718 3357 3752
rect 3391 3718 3392 3752
rect 3356 3684 3392 3718
rect 3356 3650 3357 3684
rect 3391 3650 3392 3684
rect 3356 3616 3392 3650
rect 3356 3582 3357 3616
rect 3391 3582 3392 3616
rect 3356 3548 3392 3582
rect 3356 3514 3357 3548
rect 3391 3514 3392 3548
rect 3356 3480 3392 3514
rect 3356 3446 3357 3480
rect 3391 3446 3392 3480
rect 3356 3412 3392 3446
rect 3356 3378 3357 3412
rect 3391 3378 3392 3412
rect 3356 3344 3392 3378
rect 3356 3310 3357 3344
rect 3391 3310 3392 3344
rect 3356 3276 3392 3310
rect 3356 3242 3357 3276
rect 3391 3242 3392 3276
rect 3356 3208 3392 3242
rect 3356 3174 3357 3208
rect 3391 3174 3392 3208
rect 3356 3140 3392 3174
rect 3356 3106 3357 3140
rect 3391 3106 3392 3140
rect 3356 3072 3392 3106
rect 3356 3038 3357 3072
rect 3391 3038 3392 3072
rect 3356 3004 3392 3038
rect 3356 2970 3357 3004
rect 3391 2970 3392 3004
rect 3356 2936 3392 2970
rect 3356 2902 3357 2936
rect 3391 2902 3392 2936
rect 3356 2868 3392 2902
rect 3356 2849 3357 2868
rect 574 2848 967 2849
rect 574 2838 657 2848
rect 539 2814 657 2838
rect 691 2814 729 2848
rect 775 2814 801 2848
rect 859 2814 873 2848
rect 907 2814 909 2848
rect 943 2814 967 2848
rect 1237 2848 1823 2849
rect 539 2813 967 2814
rect 1001 2813 1017 2847
rect 1083 2813 1085 2847
rect 1119 2813 1121 2847
rect 1187 2813 1203 2847
rect 1237 2814 1261 2848
rect 1295 2814 1297 2848
rect 1331 2814 1345 2848
rect 1403 2814 1429 2848
rect 1475 2814 1513 2848
rect 1547 2814 1585 2848
rect 1631 2814 1657 2848
rect 1715 2814 1729 2848
rect 1763 2814 1765 2848
rect 1799 2814 1823 2848
rect 2093 2848 2679 2849
rect 1237 2813 1823 2814
rect 1857 2813 1873 2847
rect 1939 2813 1941 2847
rect 1975 2813 1977 2847
rect 2043 2813 2059 2847
rect 2093 2814 2117 2848
rect 2151 2814 2153 2848
rect 2187 2814 2201 2848
rect 2259 2814 2285 2848
rect 2331 2814 2369 2848
rect 2403 2814 2441 2848
rect 2487 2814 2513 2848
rect 2571 2814 2585 2848
rect 2619 2814 2621 2848
rect 2655 2814 2679 2848
rect 2949 2848 3357 2849
rect 2093 2813 2679 2814
rect 2713 2813 2729 2847
rect 2795 2813 2797 2847
rect 2831 2813 2833 2847
rect 2899 2813 2915 2847
rect 2949 2814 2973 2848
rect 3007 2814 3009 2848
rect 3043 2814 3057 2848
rect 3115 2814 3141 2848
rect 3187 2814 3225 2848
rect 3259 2834 3357 2848
rect 3391 2849 3392 2868
rect 5829 5021 5830 5032
rect 5864 5021 5865 5055
rect 5829 4987 5865 5021
rect 5829 4953 5830 4987
rect 5864 4953 5865 4987
rect 5829 4919 5865 4953
rect 5829 4885 5830 4919
rect 5864 4885 5865 4919
rect 5829 4851 5865 4885
rect 5829 4817 5830 4851
rect 5864 4817 5865 4851
rect 5829 4783 5865 4817
rect 5829 4749 5830 4783
rect 5864 4749 5865 4783
rect 5829 4715 5865 4749
rect 5829 4681 5830 4715
rect 5864 4681 5865 4715
rect 5829 4647 5865 4681
rect 5829 4613 5830 4647
rect 5864 4613 5865 4647
rect 5829 4579 5865 4613
rect 5829 4545 5830 4579
rect 5864 4545 5865 4579
rect 5829 4511 5865 4545
rect 5829 4477 5830 4511
rect 5864 4477 5865 4511
rect 5829 4443 5865 4477
rect 5829 4409 5830 4443
rect 5864 4409 5865 4443
rect 5829 4375 5865 4409
rect 5829 4341 5830 4375
rect 5864 4341 5865 4375
rect 5829 4307 5865 4341
rect 5829 4273 5830 4307
rect 5864 4273 5865 4307
rect 5829 4239 5865 4273
rect 5829 4205 5830 4239
rect 5864 4205 5865 4239
rect 5829 4171 5865 4205
rect 5829 4137 5830 4171
rect 5864 4137 5865 4171
rect 5829 4103 5865 4137
rect 5829 4069 5830 4103
rect 5864 4069 5865 4103
rect 5829 4035 5865 4069
rect 5829 4001 5830 4035
rect 5864 4001 5865 4035
rect 5829 3967 5865 4001
rect 5829 3933 5830 3967
rect 5864 3933 5865 3967
rect 5829 3899 5865 3933
rect 5829 3865 5830 3899
rect 5864 3865 5865 3899
rect 5829 3831 5865 3865
rect 5829 3797 5830 3831
rect 5864 3797 5865 3831
rect 5829 3763 5865 3797
rect 5829 3729 5830 3763
rect 5864 3729 5865 3763
rect 5829 3695 5865 3729
rect 5829 3661 5830 3695
rect 5864 3661 5865 3695
rect 5829 3627 5865 3661
rect 5829 3593 5830 3627
rect 5864 3593 5865 3627
rect 5829 3559 5865 3593
rect 5829 3525 5830 3559
rect 5864 3525 5865 3559
rect 5829 3491 5865 3525
rect 5829 3457 5830 3491
rect 5864 3457 5865 3491
rect 5829 3423 5865 3457
rect 5829 3389 5830 3423
rect 5864 3389 5865 3423
rect 5829 3355 5865 3389
rect 5829 3321 5830 3355
rect 5864 3321 5865 3355
rect 5829 3287 5865 3321
rect 5829 3253 5830 3287
rect 5864 3253 5865 3287
rect 5829 3219 5865 3253
rect 5829 3185 5830 3219
rect 5864 3185 5865 3219
rect 5829 3151 5865 3185
rect 5829 3117 5830 3151
rect 5864 3117 5865 3151
rect 5829 3083 5865 3117
rect 5829 3049 5830 3083
rect 5864 3049 5865 3083
rect 5829 3015 5865 3049
rect 5829 2981 5830 3015
rect 5864 2981 5865 3015
rect 5829 2947 5865 2981
rect 5829 2913 5830 2947
rect 5864 2913 5865 2947
rect 5829 2879 5865 2913
rect 5829 2849 5830 2879
rect 3391 2848 3799 2849
rect 3391 2834 3489 2848
rect 3259 2814 3489 2834
rect 3523 2814 3561 2848
rect 3607 2814 3633 2848
rect 3691 2814 3705 2848
rect 3739 2814 3741 2848
rect 3775 2814 3799 2848
rect 4069 2848 4455 2849
rect 2949 2813 3799 2814
rect 3833 2813 3849 2847
rect 3915 2813 3917 2847
rect 3951 2813 3953 2847
rect 4019 2813 4035 2847
rect 4069 2814 4093 2848
rect 4127 2814 4129 2848
rect 4163 2814 4177 2848
rect 4235 2814 4261 2848
rect 4307 2814 4345 2848
rect 4379 2814 4455 2848
rect 4725 2848 4911 2849
rect 4069 2813 4455 2814
rect 4489 2813 4505 2847
rect 4571 2813 4573 2847
rect 4607 2813 4609 2847
rect 4675 2813 4691 2847
rect 4725 2814 4765 2848
rect 4799 2814 4801 2848
rect 4835 2814 4837 2848
rect 4871 2814 4911 2848
rect 4725 2813 4911 2814
rect 4945 2813 4961 2847
rect 5027 2813 5029 2847
rect 5063 2813 5065 2847
rect 5131 2813 5147 2847
rect 5181 2815 5221 2849
rect 5255 2848 5293 2849
rect 5255 2815 5257 2848
rect 5181 2814 5257 2815
rect 5291 2815 5293 2848
rect 5327 2815 5367 2849
rect 5637 2848 5830 2849
rect 5291 2814 5367 2815
rect 5181 2813 5367 2814
rect 5401 2813 5417 2847
rect 5483 2813 5485 2847
rect 5519 2813 5521 2847
rect 5587 2813 5603 2847
rect 5637 2814 5713 2848
rect 5747 2845 5830 2848
rect 5864 2845 5865 2879
rect 5747 2814 5865 2845
rect 5637 2813 5865 2814
rect 539 2804 575 2813
rect 539 2770 540 2804
rect 574 2770 575 2804
rect 539 2736 575 2770
rect 539 2702 540 2736
rect 574 2702 575 2736
rect 539 2584 575 2702
rect 539 2550 540 2584
rect 574 2550 575 2584
rect 539 2516 575 2550
rect 539 2482 540 2516
rect 574 2482 575 2516
rect 539 2448 575 2482
rect 539 2414 540 2448
rect 574 2414 575 2448
rect 539 2380 575 2414
rect 539 2346 540 2380
rect 574 2346 575 2380
rect 539 2312 575 2346
rect 539 2278 540 2312
rect 574 2278 575 2312
rect 539 2244 575 2278
rect 539 2210 540 2244
rect 574 2210 575 2244
rect 539 2176 575 2210
rect 539 2142 540 2176
rect 574 2142 575 2176
rect 539 2108 575 2142
rect 539 2074 540 2108
rect 574 2074 575 2108
rect 539 2040 575 2074
rect 539 2006 540 2040
rect 574 2006 575 2040
rect 539 1972 575 2006
rect 539 1938 540 1972
rect 574 1938 575 1972
rect 539 1904 575 1938
rect 539 1870 540 1904
rect 574 1870 575 1904
rect 539 1836 575 1870
rect 539 1802 540 1836
rect 574 1802 575 1836
rect 539 1768 575 1802
rect 539 1734 540 1768
rect 574 1734 575 1768
rect 539 1700 575 1734
rect 539 1666 540 1700
rect 574 1666 575 1700
rect 539 1632 575 1666
rect 539 1598 540 1632
rect 574 1598 575 1632
rect 539 1564 575 1598
rect 539 1530 540 1564
rect 574 1530 575 1564
rect 539 1496 575 1530
rect 539 1462 540 1496
rect 574 1462 575 1496
rect 539 1428 575 1462
rect 539 1394 540 1428
rect 574 1394 575 1428
rect 539 1360 575 1394
rect 539 1326 540 1360
rect 574 1326 575 1360
rect 539 1292 575 1326
rect 539 1258 540 1292
rect 574 1258 575 1292
rect 539 1224 575 1258
rect 539 1190 540 1224
rect 574 1190 575 1224
rect 539 1156 575 1190
rect 539 1122 540 1156
rect 574 1122 575 1156
rect 539 1088 575 1122
rect 539 1054 540 1088
rect 574 1054 575 1088
rect 539 1020 575 1054
rect 539 986 540 1020
rect 574 986 575 1020
rect 539 952 575 986
rect 539 918 540 952
rect 574 918 575 952
rect 539 884 575 918
rect 539 850 540 884
rect 574 850 575 884
rect 539 816 575 850
rect 539 782 540 816
rect 574 782 575 816
rect 539 748 575 782
rect 539 714 540 748
rect 574 714 575 748
rect 539 592 575 714
rect 3356 2800 3392 2813
rect 3356 2766 3357 2800
rect 3391 2766 3392 2800
rect 3356 2732 3392 2766
rect 3356 2698 3357 2732
rect 3391 2698 3392 2732
rect 3356 2664 3392 2698
rect 3356 2630 3357 2664
rect 3391 2630 3392 2664
rect 3356 2596 3392 2630
rect 3356 2562 3357 2596
rect 3391 2562 3392 2596
rect 3356 2528 3392 2562
rect 3356 2494 3357 2528
rect 3391 2494 3392 2528
rect 3356 2460 3392 2494
rect 3356 2426 3357 2460
rect 3391 2426 3392 2460
rect 3356 2392 3392 2426
rect 3356 2358 3357 2392
rect 3391 2358 3392 2392
rect 3356 2324 3392 2358
rect 3356 2290 3357 2324
rect 3391 2290 3392 2324
rect 3356 2256 3392 2290
rect 3356 2222 3357 2256
rect 3391 2222 3392 2256
rect 3356 2188 3392 2222
rect 3356 2154 3357 2188
rect 3391 2154 3392 2188
rect 3356 2120 3392 2154
rect 3356 2086 3357 2120
rect 3391 2086 3392 2120
rect 3356 2052 3392 2086
rect 3356 2018 3357 2052
rect 3391 2018 3392 2052
rect 3356 1984 3392 2018
rect 3356 1950 3357 1984
rect 3391 1950 3392 1984
rect 3356 1916 3392 1950
rect 3356 1882 3357 1916
rect 3391 1882 3392 1916
rect 3356 1848 3392 1882
rect 3356 1814 3357 1848
rect 3391 1814 3392 1848
rect 3356 1780 3392 1814
rect 3356 1746 3357 1780
rect 3391 1746 3392 1780
rect 3356 1712 3392 1746
rect 3356 1678 3357 1712
rect 3391 1678 3392 1712
rect 3356 1644 3392 1678
rect 3356 1610 3357 1644
rect 3391 1610 3392 1644
rect 3356 1576 3392 1610
rect 3356 1542 3357 1576
rect 3391 1542 3392 1576
rect 3356 1508 3392 1542
rect 3356 1474 3357 1508
rect 3391 1474 3392 1508
rect 3356 1440 3392 1474
rect 3356 1406 3357 1440
rect 3391 1406 3392 1440
rect 3356 1372 3392 1406
rect 3356 1338 3357 1372
rect 3391 1338 3392 1372
rect 3356 1304 3392 1338
rect 3356 1270 3357 1304
rect 3391 1270 3392 1304
rect 3356 1236 3392 1270
rect 3356 1202 3357 1236
rect 3391 1202 3392 1236
rect 3356 1168 3392 1202
rect 3356 1134 3357 1168
rect 3391 1134 3392 1168
rect 3356 1100 3392 1134
rect 3356 1066 3357 1100
rect 3391 1066 3392 1100
rect 3356 1032 3392 1066
rect 3356 998 3357 1032
rect 3391 998 3392 1032
rect 3356 964 3392 998
rect 3356 930 3357 964
rect 3391 930 3392 964
rect 3356 896 3392 930
rect 3356 862 3357 896
rect 3391 862 3392 896
rect 3356 828 3392 862
rect 3356 794 3357 828
rect 3391 794 3392 828
rect 3356 760 3392 794
rect 3356 726 3357 760
rect 3391 726 3392 760
rect 3356 692 3392 726
rect 3356 658 3357 692
rect 3391 658 3392 692
rect 5829 2811 5865 2813
rect 5829 2777 5830 2811
rect 5864 2777 5865 2811
rect 5829 2743 5865 2777
rect 5829 2709 5830 2743
rect 5864 2709 5865 2743
rect 5829 2675 5865 2709
rect 5829 2641 5830 2675
rect 5864 2641 5865 2675
rect 5829 2607 5865 2641
rect 5829 2573 5830 2607
rect 5864 2573 5865 2607
rect 5829 2539 5865 2573
rect 5829 2505 5830 2539
rect 5864 2505 5865 2539
rect 5829 2471 5865 2505
rect 5829 2437 5830 2471
rect 5864 2437 5865 2471
rect 5829 2403 5865 2437
rect 5829 2369 5830 2403
rect 5864 2369 5865 2403
rect 5829 2335 5865 2369
rect 5829 2301 5830 2335
rect 5864 2301 5865 2335
rect 5829 2267 5865 2301
rect 5829 2233 5830 2267
rect 5864 2233 5865 2267
rect 5829 2199 5865 2233
rect 5829 2165 5830 2199
rect 5864 2165 5865 2199
rect 5829 2131 5865 2165
rect 5829 2097 5830 2131
rect 5864 2097 5865 2131
rect 5829 2063 5865 2097
rect 5829 2029 5830 2063
rect 5864 2029 5865 2063
rect 5829 1995 5865 2029
rect 5829 1961 5830 1995
rect 5864 1961 5865 1995
rect 5829 1927 5865 1961
rect 5829 1893 5830 1927
rect 5864 1893 5865 1927
rect 5829 1859 5865 1893
rect 5829 1825 5830 1859
rect 5864 1825 5865 1859
rect 5829 1791 5865 1825
rect 5829 1757 5830 1791
rect 5864 1757 5865 1791
rect 5829 1723 5865 1757
rect 5829 1689 5830 1723
rect 5864 1689 5865 1723
rect 5829 1655 5865 1689
rect 5829 1621 5830 1655
rect 5864 1621 5865 1655
rect 5829 1587 5865 1621
rect 5829 1553 5830 1587
rect 5864 1553 5865 1587
rect 5829 1519 5865 1553
rect 5829 1485 5830 1519
rect 5864 1485 5865 1519
rect 5829 1451 5865 1485
rect 5829 1417 5830 1451
rect 5864 1417 5865 1451
rect 5829 1383 5865 1417
rect 5829 1349 5830 1383
rect 5864 1349 5865 1383
rect 5829 1315 5865 1349
rect 5829 1281 5830 1315
rect 5864 1281 5865 1315
rect 5829 1247 5865 1281
rect 5829 1213 5830 1247
rect 5864 1213 5865 1247
rect 5829 1179 5865 1213
rect 5829 1145 5830 1179
rect 5864 1145 5865 1179
rect 5829 1111 5865 1145
rect 5829 1077 5830 1111
rect 5864 1077 5865 1111
rect 5829 1043 5865 1077
rect 5829 1009 5830 1043
rect 5864 1009 5865 1043
rect 5829 975 5865 1009
rect 5829 941 5830 975
rect 5864 941 5865 975
rect 5829 907 5865 941
rect 5829 873 5830 907
rect 5864 873 5865 907
rect 5829 839 5865 873
rect 5829 805 5830 839
rect 5864 805 5865 839
rect 5829 771 5865 805
rect 5829 737 5830 771
rect 5864 737 5865 771
rect 5829 703 5865 737
rect 539 591 1021 592
rect 539 557 573 591
rect 607 557 618 591
rect 675 557 690 591
rect 743 557 762 591
rect 811 557 834 591
rect 879 557 906 591
rect 947 557 978 591
rect 1012 557 1021 591
rect 539 556 1021 557
rect 350 403 386 553
rect 1055 501 1161 642
rect 1195 591 1977 592
rect 1195 557 1253 591
rect 1287 557 1321 591
rect 1355 557 1389 591
rect 1423 557 1457 591
rect 1491 557 1525 591
rect 1559 557 1593 591
rect 1627 557 1661 591
rect 1695 557 1729 591
rect 1763 557 1797 591
rect 1831 557 1865 591
rect 1899 557 1977 591
rect 1195 556 1977 557
rect 1089 467 1127 501
rect 2011 501 2117 642
rect 2151 591 2899 592
rect 2151 557 2205 591
rect 2239 557 2273 591
rect 2307 557 2341 591
rect 2375 557 2409 591
rect 2443 557 2559 591
rect 2593 557 2627 591
rect 2661 557 2695 591
rect 2729 557 2763 591
rect 2797 557 2831 591
rect 2865 557 2899 591
rect 2151 556 2899 557
rect 2045 467 2083 501
rect 2933 501 3039 642
rect 3356 624 3392 658
rect 4421 642 4437 676
rect 4471 642 4501 676
rect 4539 642 4573 676
rect 4607 642 4641 676
rect 4679 642 4709 676
rect 4743 642 4759 676
rect 4877 642 4893 676
rect 4927 642 4957 676
rect 4995 642 5029 676
rect 5063 642 5097 676
rect 5135 642 5165 676
rect 5199 642 5215 676
rect 5279 642 5349 676
rect 5383 642 5413 676
rect 5451 642 5485 676
rect 5519 642 5553 676
rect 5591 642 5621 676
rect 5655 642 5671 676
rect 5829 669 5830 703
rect 5864 669 5865 703
rect 3356 592 3357 624
rect 3073 591 3357 592
rect 3073 557 3152 591
rect 3186 557 3220 591
rect 3254 557 3288 591
rect 3322 590 3357 591
rect 3391 592 3392 624
rect 3391 591 3698 592
rect 3391 590 3426 591
rect 3322 557 3426 590
rect 3460 557 3494 591
rect 3528 557 3562 591
rect 3596 557 3630 591
rect 3664 557 3698 591
rect 3073 556 3698 557
rect 2967 467 3005 501
rect 3746 501 3852 642
rect 3907 591 4387 592
rect 3941 557 3979 591
rect 4013 557 4047 591
rect 4085 557 4115 591
rect 4157 557 4183 591
rect 4229 557 4251 591
rect 4301 557 4319 591
rect 4373 557 4387 591
rect 3907 556 4387 557
rect 3780 467 3818 501
rect 4421 501 4527 642
rect 4561 591 4843 592
rect 4561 557 4575 591
rect 4609 557 4639 591
rect 4681 557 4707 591
rect 4753 557 4775 591
rect 4825 557 4843 591
rect 4561 556 4843 557
rect 4455 467 4493 501
rect 4877 501 4983 642
rect 5017 591 5245 592
rect 5017 557 5047 591
rect 5081 557 5109 591
rect 5153 557 5177 591
rect 5225 557 5245 591
rect 5017 556 5245 557
rect 4911 467 4949 501
rect 5279 501 5385 642
rect 5829 592 5865 669
rect 5419 591 5865 592
rect 5419 557 5446 591
rect 5491 557 5518 591
rect 5559 557 5590 591
rect 5627 557 5661 591
rect 5696 557 5729 591
rect 5768 557 5797 591
rect 5831 557 5865 591
rect 5419 556 5865 557
rect 6018 9514 6054 9548
rect 6018 9480 6019 9514
rect 6053 9480 6054 9514
rect 6018 9446 6054 9480
rect 6018 9412 6019 9446
rect 6053 9412 6054 9446
rect 6018 9378 6054 9412
rect 6018 9344 6019 9378
rect 6053 9344 6054 9378
rect 6018 9310 6054 9344
rect 6018 9276 6019 9310
rect 6053 9276 6054 9310
rect 6018 9242 6054 9276
rect 6018 9208 6019 9242
rect 6053 9208 6054 9242
rect 6018 9174 6054 9208
rect 6018 9140 6019 9174
rect 6053 9140 6054 9174
rect 6018 9106 6054 9140
rect 6018 9072 6019 9106
rect 6053 9072 6054 9106
rect 6018 9038 6054 9072
rect 6018 9004 6019 9038
rect 6053 9004 6054 9038
rect 6018 8970 6054 9004
rect 6018 8936 6019 8970
rect 6053 8936 6054 8970
rect 6018 8902 6054 8936
rect 6018 8868 6019 8902
rect 6053 8868 6054 8902
rect 6018 8834 6054 8868
rect 6018 8800 6019 8834
rect 6053 8800 6054 8834
rect 6018 8766 6054 8800
rect 6018 8732 6019 8766
rect 6053 8732 6054 8766
rect 6018 8698 6054 8732
rect 6018 8664 6019 8698
rect 6053 8664 6054 8698
rect 6018 8630 6054 8664
rect 6018 8596 6019 8630
rect 6053 8596 6054 8630
rect 6018 8562 6054 8596
rect 6018 8528 6019 8562
rect 6053 8528 6054 8562
rect 6018 8494 6054 8528
rect 6018 8460 6019 8494
rect 6053 8460 6054 8494
rect 6018 8426 6054 8460
rect 6018 8392 6019 8426
rect 6053 8392 6054 8426
rect 6018 8358 6054 8392
rect 6018 8324 6019 8358
rect 6053 8324 6054 8358
rect 6018 8290 6054 8324
rect 6018 8256 6019 8290
rect 6053 8256 6054 8290
rect 6018 8222 6054 8256
rect 6018 8188 6019 8222
rect 6053 8188 6054 8222
rect 6018 8154 6054 8188
rect 6018 8120 6019 8154
rect 6053 8120 6054 8154
rect 6018 8086 6054 8120
rect 6018 8052 6019 8086
rect 6053 8052 6054 8086
rect 6018 8018 6054 8052
rect 6018 7984 6019 8018
rect 6053 7984 6054 8018
rect 6018 7950 6054 7984
rect 6018 7916 6019 7950
rect 6053 7916 6054 7950
rect 6018 7882 6054 7916
rect 6018 7848 6019 7882
rect 6053 7848 6054 7882
rect 6018 7814 6054 7848
rect 6018 7780 6019 7814
rect 6053 7780 6054 7814
rect 6018 7746 6054 7780
rect 6018 7712 6019 7746
rect 6053 7712 6054 7746
rect 6018 7678 6054 7712
rect 6018 7644 6019 7678
rect 6053 7644 6054 7678
rect 6018 7610 6054 7644
rect 6018 7576 6019 7610
rect 6053 7576 6054 7610
rect 6018 7542 6054 7576
rect 6018 7508 6019 7542
rect 6053 7508 6054 7542
rect 6018 7474 6054 7508
rect 6018 7440 6019 7474
rect 6053 7440 6054 7474
rect 6018 7406 6054 7440
rect 6018 7372 6019 7406
rect 6053 7372 6054 7406
rect 6018 7338 6054 7372
rect 6018 7304 6019 7338
rect 6053 7304 6054 7338
rect 6018 7270 6054 7304
rect 6018 7236 6019 7270
rect 6053 7236 6054 7270
rect 6018 7202 6054 7236
rect 6018 7168 6019 7202
rect 6053 7168 6054 7202
rect 6018 7134 6054 7168
rect 6018 7100 6019 7134
rect 6053 7100 6054 7134
rect 6018 7066 6054 7100
rect 6018 7032 6019 7066
rect 6053 7032 6054 7066
rect 6018 6998 6054 7032
rect 6018 6964 6019 6998
rect 6053 6964 6054 6998
rect 6018 6930 6054 6964
rect 6018 6896 6019 6930
rect 6053 6896 6054 6930
rect 6018 6862 6054 6896
rect 6018 6828 6019 6862
rect 6053 6828 6054 6862
rect 6018 6794 6054 6828
rect 6018 6760 6019 6794
rect 6053 6760 6054 6794
rect 6018 6726 6054 6760
rect 6018 6692 6019 6726
rect 6053 6692 6054 6726
rect 6018 6658 6054 6692
rect 6018 6624 6019 6658
rect 6053 6624 6054 6658
rect 6018 6590 6054 6624
rect 6018 6556 6019 6590
rect 6053 6556 6054 6590
rect 6018 6522 6054 6556
rect 6018 6488 6019 6522
rect 6053 6488 6054 6522
rect 6018 6454 6054 6488
rect 6018 6420 6019 6454
rect 6053 6420 6054 6454
rect 6018 6386 6054 6420
rect 6018 6352 6019 6386
rect 6053 6352 6054 6386
rect 6018 6318 6054 6352
rect 6018 6284 6019 6318
rect 6053 6284 6054 6318
rect 6018 6250 6054 6284
rect 6018 6216 6019 6250
rect 6053 6216 6054 6250
rect 6018 6182 6054 6216
rect 6018 6148 6019 6182
rect 6053 6148 6054 6182
rect 6018 6114 6054 6148
rect 6018 6080 6019 6114
rect 6053 6080 6054 6114
rect 6018 6046 6054 6080
rect 6018 6012 6019 6046
rect 6053 6012 6054 6046
rect 6018 5978 6054 6012
rect 6018 5944 6019 5978
rect 6053 5944 6054 5978
rect 6018 5910 6054 5944
rect 6018 5876 6019 5910
rect 6053 5876 6054 5910
rect 6018 5842 6054 5876
rect 6018 5808 6019 5842
rect 6053 5808 6054 5842
rect 6018 5774 6054 5808
rect 6018 5740 6019 5774
rect 6053 5740 6054 5774
rect 6018 5706 6054 5740
rect 6018 5672 6019 5706
rect 6053 5672 6054 5706
rect 6018 5638 6054 5672
rect 6018 5604 6019 5638
rect 6053 5604 6054 5638
rect 6018 5570 6054 5604
rect 6018 5536 6019 5570
rect 6053 5536 6054 5570
rect 6018 5502 6054 5536
rect 6018 5468 6019 5502
rect 6053 5468 6054 5502
rect 6018 5434 6054 5468
rect 6018 5400 6019 5434
rect 6053 5400 6054 5434
rect 6018 5366 6054 5400
rect 6018 5332 6019 5366
rect 6053 5332 6054 5366
rect 6018 5298 6054 5332
rect 6018 5264 6019 5298
rect 6053 5264 6054 5298
rect 6018 5230 6054 5264
rect 6018 5196 6019 5230
rect 6053 5196 6054 5230
rect 6018 5162 6054 5196
rect 6018 5128 6019 5162
rect 6053 5128 6054 5162
rect 6018 5094 6054 5128
rect 6018 5060 6019 5094
rect 6053 5060 6054 5094
rect 6018 5026 6054 5060
rect 6018 4992 6019 5026
rect 6053 4992 6054 5026
rect 6018 4958 6054 4992
rect 6018 4924 6019 4958
rect 6053 4924 6054 4958
rect 6018 4890 6054 4924
rect 6018 4856 6019 4890
rect 6053 4856 6054 4890
rect 6018 4822 6054 4856
rect 6018 4788 6019 4822
rect 6053 4788 6054 4822
rect 6018 4754 6054 4788
rect 6018 4720 6019 4754
rect 6053 4720 6054 4754
rect 6018 4686 6054 4720
rect 6018 4652 6019 4686
rect 6053 4652 6054 4686
rect 6018 4618 6054 4652
rect 6018 4584 6019 4618
rect 6053 4584 6054 4618
rect 6018 4550 6054 4584
rect 6018 4516 6019 4550
rect 6053 4516 6054 4550
rect 6018 4482 6054 4516
rect 6018 4448 6019 4482
rect 6053 4448 6054 4482
rect 6018 4414 6054 4448
rect 6018 4380 6019 4414
rect 6053 4380 6054 4414
rect 6018 4346 6054 4380
rect 6018 4312 6019 4346
rect 6053 4312 6054 4346
rect 6018 4278 6054 4312
rect 6018 4244 6019 4278
rect 6053 4244 6054 4278
rect 6018 4210 6054 4244
rect 6018 4176 6019 4210
rect 6053 4176 6054 4210
rect 6018 4142 6054 4176
rect 6018 4108 6019 4142
rect 6053 4108 6054 4142
rect 6018 4074 6054 4108
rect 6018 4040 6019 4074
rect 6053 4040 6054 4074
rect 6018 4006 6054 4040
rect 6018 3972 6019 4006
rect 6053 3972 6054 4006
rect 6018 3938 6054 3972
rect 6018 3904 6019 3938
rect 6053 3904 6054 3938
rect 6018 3870 6054 3904
rect 6018 3836 6019 3870
rect 6053 3836 6054 3870
rect 6018 3802 6054 3836
rect 6018 3768 6019 3802
rect 6053 3768 6054 3802
rect 6018 3734 6054 3768
rect 6018 3700 6019 3734
rect 6053 3700 6054 3734
rect 6018 3666 6054 3700
rect 6018 3632 6019 3666
rect 6053 3632 6054 3666
rect 6018 3598 6054 3632
rect 6018 3564 6019 3598
rect 6053 3564 6054 3598
rect 6018 3530 6054 3564
rect 6018 3496 6019 3530
rect 6053 3496 6054 3530
rect 6018 3462 6054 3496
rect 6018 3428 6019 3462
rect 6053 3428 6054 3462
rect 6018 3394 6054 3428
rect 6018 3360 6019 3394
rect 6053 3360 6054 3394
rect 6018 3326 6054 3360
rect 6018 3292 6019 3326
rect 6053 3292 6054 3326
rect 6018 3258 6054 3292
rect 6018 3224 6019 3258
rect 6053 3224 6054 3258
rect 6018 3190 6054 3224
rect 6018 3156 6019 3190
rect 6053 3156 6054 3190
rect 6018 3122 6054 3156
rect 6018 3088 6019 3122
rect 6053 3088 6054 3122
rect 6018 3054 6054 3088
rect 6018 3020 6019 3054
rect 6053 3020 6054 3054
rect 6018 2986 6054 3020
rect 6018 2952 6019 2986
rect 6053 2952 6054 2986
rect 6018 2918 6054 2952
rect 6018 2884 6019 2918
rect 6053 2884 6054 2918
rect 6018 2850 6054 2884
rect 6018 2816 6019 2850
rect 6053 2816 6054 2850
rect 6018 2782 6054 2816
rect 6018 2748 6019 2782
rect 6053 2748 6054 2782
rect 6018 2714 6054 2748
rect 6018 2680 6019 2714
rect 6053 2680 6054 2714
rect 6018 2646 6054 2680
rect 6018 2612 6019 2646
rect 6053 2612 6054 2646
rect 6018 2578 6054 2612
rect 6018 2544 6019 2578
rect 6053 2544 6054 2578
rect 6018 2510 6054 2544
rect 6018 2476 6019 2510
rect 6053 2476 6054 2510
rect 6018 2442 6054 2476
rect 6018 2408 6019 2442
rect 6053 2408 6054 2442
rect 6018 2374 6054 2408
rect 6018 2340 6019 2374
rect 6053 2340 6054 2374
rect 6018 2306 6054 2340
rect 6018 2272 6019 2306
rect 6053 2272 6054 2306
rect 6018 2238 6054 2272
rect 6018 2204 6019 2238
rect 6053 2204 6054 2238
rect 6018 2170 6054 2204
rect 6018 2136 6019 2170
rect 6053 2136 6054 2170
rect 6018 2102 6054 2136
rect 6018 2068 6019 2102
rect 6053 2068 6054 2102
rect 6018 2034 6054 2068
rect 6018 2000 6019 2034
rect 6053 2000 6054 2034
rect 6018 1966 6054 2000
rect 6018 1932 6019 1966
rect 6053 1932 6054 1966
rect 6018 1898 6054 1932
rect 6018 1864 6019 1898
rect 6053 1864 6054 1898
rect 6018 1830 6054 1864
rect 6018 1796 6019 1830
rect 6053 1796 6054 1830
rect 6018 1762 6054 1796
rect 6018 1728 6019 1762
rect 6053 1728 6054 1762
rect 6018 1694 6054 1728
rect 6018 1660 6019 1694
rect 6053 1660 6054 1694
rect 6018 1626 6054 1660
rect 6018 1592 6019 1626
rect 6053 1592 6054 1626
rect 6018 1558 6054 1592
rect 6018 1524 6019 1558
rect 6053 1524 6054 1558
rect 6018 1490 6054 1524
rect 6018 1456 6019 1490
rect 6053 1456 6054 1490
rect 6018 1422 6054 1456
rect 6018 1388 6019 1422
rect 6053 1388 6054 1422
rect 6018 1354 6054 1388
rect 6018 1320 6019 1354
rect 6053 1320 6054 1354
rect 6018 1286 6054 1320
rect 6018 1252 6019 1286
rect 6053 1252 6054 1286
rect 6018 1218 6054 1252
rect 6018 1184 6019 1218
rect 6053 1184 6054 1218
rect 6018 1150 6054 1184
rect 6018 1116 6019 1150
rect 6053 1116 6054 1150
rect 6018 1082 6054 1116
rect 6018 1048 6019 1082
rect 6053 1048 6054 1082
rect 6018 1014 6054 1048
rect 6018 980 6019 1014
rect 6053 980 6054 1014
rect 6018 946 6054 980
rect 6018 912 6019 946
rect 6053 912 6054 946
rect 6018 878 6054 912
rect 6018 844 6019 878
rect 6053 844 6054 878
rect 6018 810 6054 844
rect 6018 776 6019 810
rect 6053 776 6054 810
rect 6018 742 6054 776
rect 6018 708 6019 742
rect 6053 708 6054 742
rect 6018 674 6054 708
rect 6018 640 6019 674
rect 6053 640 6054 674
rect 6018 606 6054 640
rect 6018 572 6019 606
rect 6053 572 6054 606
rect 5313 467 5351 501
rect 6018 538 6054 572
rect 6018 504 6019 538
rect 6053 504 6054 538
rect 6018 435 6054 504
rect 6018 403 6019 435
rect 350 402 6019 403
rect 350 368 384 402
rect 418 368 452 402
rect 486 368 520 402
rect 554 368 588 402
rect 622 368 656 402
rect 690 368 724 402
rect 758 368 792 402
rect 826 368 860 402
rect 894 368 928 402
rect 962 368 996 402
rect 1030 368 1064 402
rect 1098 368 1132 402
rect 1166 368 1200 402
rect 1234 368 1268 402
rect 1302 368 1336 402
rect 1370 368 1404 402
rect 1438 368 1472 402
rect 1506 368 1540 402
rect 1574 368 1608 402
rect 1642 368 1676 402
rect 1710 368 1744 402
rect 1778 368 1812 402
rect 1846 368 1880 402
rect 1914 368 1948 402
rect 1982 368 2016 402
rect 2050 368 2084 402
rect 2118 368 2152 402
rect 2186 368 2220 402
rect 2254 368 2288 402
rect 2322 368 2356 402
rect 2390 368 2424 402
rect 2458 368 2492 402
rect 2526 368 2560 402
rect 2594 368 2628 402
rect 2662 368 2696 402
rect 2730 368 2764 402
rect 2798 368 2832 402
rect 2866 368 2900 402
rect 2934 368 2968 402
rect 3002 368 3036 402
rect 3070 368 3104 402
rect 3138 368 3172 402
rect 3206 368 3240 402
rect 3274 368 3308 402
rect 3342 368 3376 402
rect 3410 368 3444 402
rect 3478 368 3512 402
rect 3546 368 3580 402
rect 3614 368 3648 402
rect 3682 368 3716 402
rect 3750 368 3784 402
rect 3818 368 3852 402
rect 3886 368 3920 402
rect 3954 368 3988 402
rect 4022 368 4056 402
rect 4090 368 4124 402
rect 4158 368 4192 402
rect 4226 368 4260 402
rect 4294 368 4328 402
rect 4362 368 4396 402
rect 4430 368 4464 402
rect 4498 368 4532 402
rect 4566 368 4600 402
rect 4634 368 4668 402
rect 4702 368 4736 402
rect 4770 368 4804 402
rect 4838 368 4872 402
rect 4906 368 4940 402
rect 4974 368 5008 402
rect 5042 368 5076 402
rect 5110 368 5144 402
rect 5178 368 5212 402
rect 5246 368 5280 402
rect 5314 368 5348 402
rect 5382 368 5416 402
rect 5450 368 5484 402
rect 5518 368 5552 402
rect 5586 368 5620 402
rect 5654 368 5688 402
rect 5722 368 5756 402
rect 5790 368 5824 402
rect 5858 368 5892 402
rect 5926 401 6019 402
rect 6053 401 6054 435
rect 5926 368 6054 401
rect 350 367 6054 368
<< viali >>
rect 9795 34762 9829 34796
rect 9867 34762 9901 34796
rect 9939 34762 9951 34796
rect 9951 34762 9973 34796
rect 10011 34762 10019 34796
rect 10019 34762 10045 34796
rect 10083 34762 10087 34796
rect 10087 34762 10117 34796
rect 10155 34762 10189 34796
rect 10227 34762 10257 34796
rect 10257 34762 10261 34796
rect 10299 34762 10325 34796
rect 10325 34762 10333 34796
rect 10371 34762 10393 34796
rect 10393 34762 10405 34796
rect 10443 34762 10461 34796
rect 10461 34762 10477 34796
rect 10515 34762 10529 34796
rect 10529 34762 10549 34796
rect 10587 34762 10597 34796
rect 10597 34762 10621 34796
rect 10659 34762 10665 34796
rect 10665 34762 10693 34796
rect 10731 34762 10733 34796
rect 10733 34762 10765 34796
rect 10803 34762 10835 34796
rect 10835 34762 10837 34796
rect 10875 34762 10903 34796
rect 10903 34762 10909 34796
rect 10947 34762 10971 34796
rect 10971 34762 10981 34796
rect 11019 34762 11039 34796
rect 11039 34762 11053 34796
rect 11091 34762 11107 34796
rect 11107 34762 11125 34796
rect 11163 34762 11175 34796
rect 11175 34762 11197 34796
rect 11235 34762 11243 34796
rect 11243 34762 11269 34796
rect 11307 34762 11311 34796
rect 11311 34762 11341 34796
rect 11379 34762 11413 34796
rect 11451 34762 11481 34796
rect 11481 34762 11485 34796
rect 11523 34762 11549 34796
rect 11549 34762 11557 34796
rect 11595 34762 11617 34796
rect 11617 34762 11629 34796
rect 11667 34762 11685 34796
rect 11685 34762 11701 34796
rect 11739 34762 11753 34796
rect 11753 34762 11773 34796
rect 11811 34762 11821 34796
rect 11821 34762 11845 34796
rect 11883 34762 11889 34796
rect 11889 34762 11917 34796
rect 11955 34762 11957 34796
rect 11957 34762 11989 34796
rect 12027 34762 12059 34796
rect 12059 34762 12061 34796
rect 12099 34762 12127 34796
rect 12127 34762 12133 34796
rect 12171 34762 12195 34796
rect 12195 34762 12205 34796
rect 12243 34762 12263 34796
rect 12263 34762 12277 34796
rect 12315 34762 12331 34796
rect 12331 34762 12349 34796
rect 12387 34762 12399 34796
rect 12399 34762 12421 34796
rect 12459 34762 12467 34796
rect 12467 34762 12493 34796
rect 12531 34762 12535 34796
rect 12535 34762 12565 34796
rect 12603 34762 12637 34796
rect 12675 34762 12705 34796
rect 12705 34762 12709 34796
rect 12747 34762 12773 34796
rect 12773 34762 12781 34796
rect 12819 34762 12841 34796
rect 12841 34762 12853 34796
rect 12891 34762 12909 34796
rect 12909 34762 12925 34796
rect 12963 34762 12977 34796
rect 12977 34762 12997 34796
rect 13035 34762 13045 34796
rect 13045 34762 13069 34796
rect 13107 34762 13113 34796
rect 13113 34762 13141 34796
rect 13179 34762 13181 34796
rect 13181 34762 13213 34796
rect 13251 34762 13283 34796
rect 13283 34762 13285 34796
rect 13323 34762 13351 34796
rect 13351 34762 13357 34796
rect 13395 34762 13419 34796
rect 13419 34762 13429 34796
rect 13467 34762 13487 34796
rect 13487 34762 13501 34796
rect 13539 34762 13555 34796
rect 13555 34762 13573 34796
rect 13611 34762 13623 34796
rect 13623 34762 13645 34796
rect 13683 34762 13691 34796
rect 13691 34762 13717 34796
rect 13755 34762 13759 34796
rect 13759 34762 13789 34796
rect 13827 34762 13861 34796
rect 13899 34762 13929 34796
rect 13929 34762 13933 34796
rect 13971 34762 13997 34796
rect 13997 34762 14005 34796
rect 14043 34762 14065 34796
rect 14065 34762 14077 34796
rect 14115 34762 14133 34796
rect 14133 34762 14149 34796
rect 14187 34762 14201 34796
rect 14201 34762 14221 34796
rect 14259 34762 14269 34796
rect 14269 34762 14293 34796
rect 14331 34762 14337 34796
rect 14337 34762 14365 34796
rect 14405 34756 14439 34790
rect 9789 34694 9823 34708
rect 9789 34674 9823 34694
rect 9789 34626 9823 34636
rect 9789 34602 9823 34626
rect 9789 34558 9823 34564
rect 9789 34530 9823 34558
rect 14405 34704 14439 34718
rect 14405 34684 14439 34704
rect 14405 34612 14439 34646
rect 9789 34490 9823 34492
rect 9789 34458 9823 34490
rect 9789 34388 9823 34420
rect 9789 34386 9823 34388
rect 9789 34320 9823 34348
rect 9789 34314 9823 34320
rect 9789 34252 9823 34276
rect 9789 34242 9823 34252
rect 10046 34512 10080 34546
rect 10118 34512 10147 34546
rect 10147 34512 10152 34546
rect 10190 34512 10215 34546
rect 10215 34512 10224 34546
rect 10262 34512 10283 34546
rect 10283 34512 10296 34546
rect 10334 34512 10351 34546
rect 10351 34512 10368 34546
rect 10406 34512 10419 34546
rect 10419 34512 10440 34546
rect 10478 34512 10487 34546
rect 10487 34512 10512 34546
rect 10550 34512 10555 34546
rect 10555 34512 10584 34546
rect 10622 34512 10623 34546
rect 10623 34512 10656 34546
rect 10694 34512 10725 34546
rect 10725 34512 10728 34546
rect 10766 34512 10793 34546
rect 10793 34512 10800 34546
rect 10838 34512 10861 34546
rect 10861 34512 10872 34546
rect 10910 34512 10929 34546
rect 10929 34512 10944 34546
rect 10982 34512 10997 34546
rect 10997 34512 11016 34546
rect 11054 34512 11065 34546
rect 11065 34512 11088 34546
rect 11126 34512 11133 34546
rect 11133 34512 11160 34546
rect 11198 34512 11201 34546
rect 11201 34512 11232 34546
rect 11270 34512 11303 34546
rect 11303 34512 11304 34546
rect 11342 34512 11371 34546
rect 11371 34512 11376 34546
rect 11414 34512 11439 34546
rect 11439 34512 11448 34546
rect 11486 34512 11507 34546
rect 11507 34512 11520 34546
rect 11558 34512 11575 34546
rect 11575 34512 11592 34546
rect 11630 34512 11643 34546
rect 11643 34512 11664 34546
rect 11702 34512 11711 34546
rect 11711 34512 11736 34546
rect 11774 34512 11779 34546
rect 11779 34512 11808 34546
rect 11846 34512 11847 34546
rect 11847 34512 11880 34546
rect 11918 34512 11949 34546
rect 11949 34512 11952 34546
rect 11990 34512 12017 34546
rect 12017 34512 12024 34546
rect 12062 34512 12085 34546
rect 12085 34512 12096 34546
rect 12134 34512 12153 34546
rect 12153 34512 12168 34546
rect 12206 34512 12221 34546
rect 12221 34512 12240 34546
rect 12278 34512 12289 34546
rect 12289 34512 12312 34546
rect 12350 34512 12357 34546
rect 12357 34512 12384 34546
rect 12422 34512 12425 34546
rect 12425 34512 12456 34546
rect 12494 34512 12527 34546
rect 12527 34512 12528 34546
rect 12566 34512 12595 34546
rect 12595 34512 12600 34546
rect 12638 34512 12663 34546
rect 12663 34512 12672 34546
rect 12710 34512 12731 34546
rect 12731 34512 12744 34546
rect 12782 34512 12799 34546
rect 12799 34512 12816 34546
rect 12854 34512 12867 34546
rect 12867 34512 12888 34546
rect 12926 34512 12935 34546
rect 12935 34512 12960 34546
rect 12998 34512 13003 34546
rect 13003 34512 13032 34546
rect 13070 34512 13071 34546
rect 13071 34512 13104 34546
rect 13142 34512 13173 34546
rect 13173 34512 13176 34546
rect 13214 34512 13241 34546
rect 13241 34512 13248 34546
rect 13286 34512 13309 34546
rect 13309 34512 13320 34546
rect 13358 34512 13377 34546
rect 13377 34512 13392 34546
rect 13430 34512 13445 34546
rect 13445 34512 13464 34546
rect 13502 34512 13513 34546
rect 13513 34512 13536 34546
rect 13574 34512 13581 34546
rect 13581 34512 13608 34546
rect 13646 34512 13649 34546
rect 13649 34512 13680 34546
rect 13718 34512 13751 34546
rect 13751 34512 13752 34546
rect 13790 34512 13819 34546
rect 13819 34512 13824 34546
rect 13862 34512 13887 34546
rect 13887 34512 13896 34546
rect 13934 34512 13955 34546
rect 13955 34512 13968 34546
rect 14006 34512 14023 34546
rect 14023 34512 14040 34546
rect 14078 34512 14091 34546
rect 14091 34512 14112 34546
rect 14159 34506 14193 34540
rect 10219 34420 10223 34454
rect 10223 34420 10253 34454
rect 10292 34420 10297 34454
rect 10297 34420 10326 34454
rect 10365 34420 10371 34454
rect 10371 34420 10399 34454
rect 10438 34420 10445 34454
rect 10445 34420 10472 34454
rect 10510 34420 10519 34454
rect 10519 34420 10544 34454
rect 10582 34420 10592 34454
rect 10592 34420 10616 34454
rect 11105 34420 11113 34454
rect 11113 34420 11139 34454
rect 11178 34420 11182 34454
rect 11182 34420 11212 34454
rect 11251 34420 11285 34454
rect 11324 34420 11355 34454
rect 11355 34420 11358 34454
rect 11397 34420 11424 34454
rect 11424 34420 11431 34454
rect 11470 34420 11493 34454
rect 11493 34420 11504 34454
rect 11543 34420 11562 34454
rect 11562 34420 11577 34454
rect 11616 34420 11631 34454
rect 11631 34420 11650 34454
rect 11689 34420 11700 34454
rect 11700 34420 11723 34454
rect 11762 34420 11769 34454
rect 11769 34420 11796 34454
rect 11835 34420 11838 34454
rect 11838 34420 11869 34454
rect 11908 34420 11941 34454
rect 11941 34420 11942 34454
rect 11981 34420 12010 34454
rect 12010 34420 12015 34454
rect 12054 34420 12079 34454
rect 12079 34420 12088 34454
rect 12127 34420 12148 34454
rect 12148 34420 12161 34454
rect 12200 34420 12217 34454
rect 12217 34420 12234 34454
rect 12273 34420 12286 34454
rect 12286 34420 12307 34454
rect 12346 34420 12355 34454
rect 12355 34420 12380 34454
rect 12419 34420 12424 34454
rect 12424 34420 12453 34454
rect 12492 34420 12493 34454
rect 12493 34420 12526 34454
rect 12565 34420 12597 34454
rect 12597 34420 12599 34454
rect 12638 34420 12666 34454
rect 12666 34420 12672 34454
rect 12711 34420 12735 34454
rect 12735 34420 12745 34454
rect 12784 34420 12804 34454
rect 12804 34420 12818 34454
rect 12857 34420 12873 34454
rect 12873 34420 12891 34454
rect 12930 34420 12942 34454
rect 12942 34420 12964 34454
rect 13003 34420 13011 34454
rect 13011 34420 13037 34454
rect 13076 34420 13080 34454
rect 13080 34420 13110 34454
rect 13149 34420 13183 34454
rect 13222 34420 13252 34454
rect 13252 34420 13256 34454
rect 13295 34420 13321 34454
rect 13321 34420 13329 34454
rect 13368 34420 13390 34454
rect 13390 34420 13402 34454
rect 13441 34420 13459 34454
rect 13459 34420 13475 34454
rect 13514 34420 13528 34454
rect 13528 34420 13548 34454
rect 13587 34420 13597 34454
rect 13597 34420 13621 34454
rect 13660 34420 13666 34454
rect 13666 34420 13694 34454
rect 13733 34420 13735 34454
rect 13735 34420 13767 34454
rect 13806 34420 13840 34454
rect 13880 34420 13911 34454
rect 13911 34420 13914 34454
rect 14159 34434 14193 34468
rect 10040 34410 10074 34420
rect 10040 34386 10074 34410
rect 10040 34342 10074 34348
rect 10040 34314 10074 34342
rect 10040 34274 10074 34276
rect 10040 34242 10074 34274
rect 14159 34385 14193 34396
rect 14159 34362 14193 34385
rect 14159 34317 14193 34324
rect 14159 34290 14193 34317
rect 14159 34249 14193 34252
rect 14159 34218 14193 34249
rect 14159 34147 14193 34180
rect 14159 34146 14193 34147
rect 14159 34079 14193 34108
rect 14159 34074 14193 34079
rect 14159 34011 14193 34036
rect 14159 34002 14193 34011
rect 14159 33943 14193 33964
rect 14159 33930 14193 33943
rect 14159 33875 14193 33892
rect 14159 33858 14193 33875
rect 14159 33807 14193 33820
rect 14159 33786 14193 33807
rect 14159 33739 14193 33748
rect 14159 33714 14193 33739
rect 10040 33594 10074 33596
rect 10040 33562 10074 33594
rect 14159 33671 14193 33676
rect 14159 33642 14193 33671
rect 14159 33603 14193 33604
rect 14159 33570 14193 33603
rect 10040 33492 10074 33524
rect 10040 33490 10074 33492
rect 9842 33453 9876 33487
rect 9842 33380 9876 33414
rect 9842 33307 9876 33341
rect 9842 33233 9876 33267
rect 9842 33159 9876 33193
rect 10040 33424 10074 33452
rect 10040 33418 10074 33424
rect 10040 33356 10074 33380
rect 10040 33346 10074 33356
rect 10040 33288 10074 33308
rect 10040 33274 10074 33288
rect 10040 33220 10074 33236
rect 10040 33202 10074 33220
rect 10040 33152 10074 33164
rect 10040 33130 10074 33152
rect 10162 33533 10196 33567
rect 10162 33458 10196 33492
rect 10162 33383 10196 33417
rect 10162 33308 10196 33342
rect 10162 33233 10196 33267
rect 10162 33159 10196 33193
rect 11018 33533 11052 33567
rect 11018 33458 11052 33492
rect 11018 33383 11052 33417
rect 11018 33308 11052 33342
rect 11018 33233 11052 33267
rect 11018 33159 11052 33193
rect 11874 33533 11908 33567
rect 11874 33458 11908 33492
rect 11874 33383 11908 33417
rect 11874 33308 11908 33342
rect 11874 33233 11908 33267
rect 11874 33159 11908 33193
rect 12730 33533 12764 33567
rect 12730 33458 12764 33492
rect 12730 33383 12764 33417
rect 12730 33308 12764 33342
rect 12730 33233 12764 33267
rect 12730 33159 12764 33193
rect 13586 33533 13620 33567
rect 13586 33458 13620 33492
rect 13586 33383 13620 33417
rect 13586 33308 13620 33342
rect 13586 33233 13620 33267
rect 13586 33159 13620 33193
rect 14042 33533 14076 33567
rect 14042 33458 14076 33492
rect 14042 33383 14076 33417
rect 14042 33308 14076 33342
rect 14042 33233 14076 33267
rect 14042 33159 14076 33193
rect 14159 33501 14193 33532
rect 14159 33498 14193 33501
rect 14159 33433 14193 33452
rect 14159 33418 14193 33433
rect 14159 33365 14193 33380
rect 14159 33346 14193 33365
rect 14159 33297 14193 33308
rect 14159 33274 14193 33297
rect 14159 33229 14193 33236
rect 14159 33202 14193 33229
rect 10040 33084 10074 33092
rect 10040 33058 10074 33084
rect 10040 33016 10074 33020
rect 10040 32986 10074 33016
rect 10040 32914 10074 32948
rect 10040 32846 10074 32876
rect 10040 32842 10074 32846
rect 10040 32778 10074 32804
rect 10040 32770 10074 32778
rect 10040 32710 10074 32732
rect 10040 32698 10074 32710
rect 10040 32642 10074 32660
rect 10040 32626 10074 32642
rect 10040 32574 10074 32588
rect 10040 32554 10074 32574
rect 10040 32506 10074 32516
rect 10040 32482 10074 32506
rect 10040 32438 10074 32444
rect 10040 32410 10074 32438
rect 10040 32370 10074 32372
rect 10040 32338 10074 32370
rect 14159 33161 14193 33164
rect 14159 33130 14193 33161
rect 14159 33059 14193 33092
rect 14159 33058 14193 33059
rect 14159 32991 14193 33020
rect 14159 32986 14193 32991
rect 14159 32923 14193 32948
rect 14159 32914 14193 32923
rect 14159 32855 14193 32876
rect 14159 32842 14193 32855
rect 14159 32787 14193 32804
rect 14159 32770 14193 32787
rect 14159 32719 14193 32732
rect 14159 32698 14193 32719
rect 14159 32651 14193 32660
rect 14159 32626 14193 32651
rect 14159 32583 14193 32588
rect 14159 32554 14193 32583
rect 14159 32515 14193 32516
rect 14159 32482 14193 32515
rect 14159 32413 14193 32444
rect 14159 32410 14193 32413
rect 14159 32345 14193 32372
rect 14159 32338 14193 32345
rect 10040 32268 10074 32300
rect 10040 32266 10074 32268
rect 10112 32260 10142 32294
rect 10142 32260 10146 32294
rect 10185 32260 10193 32294
rect 10193 32260 10219 32294
rect 10258 32260 10278 32294
rect 10278 32260 10292 32294
rect 10331 32260 10363 32294
rect 10363 32260 10365 32294
rect 10404 32260 10438 32294
rect 10477 32260 10482 32294
rect 10482 32260 10511 32294
rect 10550 32260 10567 32294
rect 10567 32260 10584 32294
rect 10623 32260 10652 32294
rect 10652 32260 10657 32294
rect 10696 32260 10703 32294
rect 10703 32260 10730 32294
rect 10769 32260 10788 32294
rect 10788 32260 10803 32294
rect 10842 32260 10873 32294
rect 10873 32260 10876 32294
rect 10915 32260 10949 32294
rect 10988 32260 10992 32294
rect 10992 32260 11022 32294
rect 11061 32260 11077 32294
rect 11077 32260 11095 32294
rect 11134 32260 11162 32294
rect 11162 32260 11168 32294
rect 11207 32260 11213 32294
rect 11213 32260 11241 32294
rect 11279 32260 11298 32294
rect 11298 32260 11313 32294
rect 11351 32260 11383 32294
rect 11383 32260 11385 32294
rect 11423 32260 11457 32294
rect 11495 32260 11502 32294
rect 11502 32260 11529 32294
rect 11567 32260 11587 32294
rect 11587 32260 11601 32294
rect 11639 32260 11672 32294
rect 11672 32260 11673 32294
rect 11711 32260 11723 32294
rect 11723 32260 11745 32294
rect 11783 32260 11808 32294
rect 11808 32260 11817 32294
rect 11855 32260 11889 32294
rect 11927 32260 11961 32294
rect 11999 32260 12012 32294
rect 12012 32260 12033 32294
rect 12071 32260 12097 32294
rect 12097 32260 12105 32294
rect 12143 32260 12148 32294
rect 12148 32260 12177 32294
rect 12215 32260 12233 32294
rect 12233 32260 12249 32294
rect 12287 32260 12318 32294
rect 12318 32260 12321 32294
rect 12359 32260 12393 32294
rect 12431 32260 12437 32294
rect 12437 32260 12465 32294
rect 12503 32260 12522 32294
rect 12522 32260 12537 32294
rect 12575 32260 12607 32294
rect 12607 32260 12609 32294
rect 12647 32260 12658 32294
rect 12658 32260 12681 32294
rect 12719 32260 12743 32294
rect 12743 32260 12753 32294
rect 12791 32260 12825 32294
rect 12863 32260 12897 32294
rect 12935 32260 12947 32294
rect 12947 32260 12969 32294
rect 13007 32260 13032 32294
rect 13032 32260 13041 32294
rect 13079 32260 13083 32294
rect 13083 32260 13113 32294
rect 13151 32260 13167 32294
rect 13167 32260 13185 32294
rect 13223 32260 13251 32294
rect 13251 32260 13257 32294
rect 13295 32260 13329 32294
rect 13367 32260 13369 32294
rect 13369 32260 13401 32294
rect 13439 32260 13453 32294
rect 13453 32260 13473 32294
rect 13511 32260 13537 32294
rect 13537 32260 13545 32294
rect 13583 32260 13587 32294
rect 13587 32260 13617 32294
rect 13655 32260 13671 32294
rect 13671 32260 13689 32294
rect 13727 32260 13755 32294
rect 13755 32260 13761 32294
rect 13799 32260 13833 32294
rect 13871 32260 13873 32294
rect 13873 32260 13905 32294
rect 13943 32260 13957 32294
rect 13957 32260 13977 32294
rect 14015 32260 14041 32294
rect 14041 32260 14049 32294
rect 14087 32260 14091 32294
rect 14091 32260 14121 32294
rect 14159 32277 14193 32300
rect 14159 32266 14193 32277
rect 9534 32168 9568 32202
rect 9611 32168 9645 32202
rect 9688 32168 9722 32202
rect 10219 32168 10223 32202
rect 10223 32168 10253 32202
rect 10304 32168 10331 32202
rect 10331 32168 10338 32202
rect 10389 32168 10405 32202
rect 10405 32168 10423 32202
rect 10474 32168 10479 32202
rect 10479 32168 10508 32202
rect 10559 32168 10592 32202
rect 10592 32168 10593 32202
rect 10643 32168 10665 32202
rect 10665 32168 10677 32202
rect 11105 32168 11113 32202
rect 11113 32168 11139 32202
rect 11178 32168 11182 32202
rect 11182 32168 11212 32202
rect 11251 32168 11285 32202
rect 11324 32168 11355 32202
rect 11355 32168 11358 32202
rect 11397 32168 11424 32202
rect 11424 32168 11431 32202
rect 11470 32168 11493 32202
rect 11493 32168 11504 32202
rect 11543 32168 11562 32202
rect 11562 32168 11577 32202
rect 11616 32168 11631 32202
rect 11631 32168 11650 32202
rect 11689 32168 11700 32202
rect 11700 32168 11723 32202
rect 11762 32168 11769 32202
rect 11769 32168 11796 32202
rect 11835 32168 11838 32202
rect 11838 32168 11869 32202
rect 11908 32168 11941 32202
rect 11941 32168 11942 32202
rect 11981 32168 12010 32202
rect 12010 32168 12015 32202
rect 12054 32168 12079 32202
rect 12079 32168 12088 32202
rect 12127 32168 12148 32202
rect 12148 32168 12161 32202
rect 12200 32168 12217 32202
rect 12217 32168 12234 32202
rect 12273 32168 12286 32202
rect 12286 32168 12307 32202
rect 12346 32168 12355 32202
rect 12355 32168 12380 32202
rect 12419 32168 12424 32202
rect 12424 32168 12453 32202
rect 12492 32168 12493 32202
rect 12493 32168 12526 32202
rect 12565 32168 12597 32202
rect 12597 32168 12599 32202
rect 12638 32168 12666 32202
rect 12666 32168 12672 32202
rect 12711 32168 12735 32202
rect 12735 32168 12745 32202
rect 12784 32168 12804 32202
rect 12804 32168 12818 32202
rect 12857 32168 12873 32202
rect 12873 32168 12891 32202
rect 12930 32168 12942 32202
rect 12942 32168 12964 32202
rect 13003 32168 13011 32202
rect 13011 32168 13037 32202
rect 13076 32168 13080 32202
rect 13080 32168 13110 32202
rect 13149 32168 13183 32202
rect 13222 32168 13252 32202
rect 13252 32168 13256 32202
rect 13295 32168 13321 32202
rect 13321 32168 13329 32202
rect 13368 32168 13390 32202
rect 13390 32168 13402 32202
rect 13441 32168 13459 32202
rect 13459 32168 13475 32202
rect 13514 32168 13528 32202
rect 13528 32168 13548 32202
rect 13587 32168 13597 32202
rect 13597 32168 13621 32202
rect 13660 32168 13666 32202
rect 13666 32168 13694 32202
rect 13733 32168 13735 32202
rect 13735 32168 13767 32202
rect 13806 32168 13840 32202
rect 13880 32168 13911 32202
rect 13911 32168 13914 32202
rect 14159 32209 14193 32228
rect 14159 32194 14193 32209
rect 14159 32141 14193 32156
rect 14159 32122 14193 32141
rect 14159 32073 14193 32084
rect 14159 32050 14193 32073
rect 14159 32005 14193 32012
rect 14159 31978 14193 32005
rect 14159 31937 14193 31940
rect 14159 31906 14193 31937
rect 14159 31835 14193 31868
rect 14159 31834 14193 31835
rect 14159 31767 14193 31796
rect 14159 31762 14193 31767
rect 14159 31699 14193 31724
rect 14159 31690 14193 31699
rect 10040 31554 10074 31578
rect 10040 31544 10074 31554
rect 10040 31486 10074 31506
rect 10040 31472 10074 31486
rect 10040 31418 10074 31434
rect 10040 31400 10074 31418
rect 10040 31350 10074 31362
rect 10040 31328 10074 31350
rect 10040 31282 10074 31290
rect 10040 31256 10074 31282
rect 14159 31631 14193 31652
rect 14159 31618 14193 31631
rect 14159 31563 14193 31580
rect 14159 31546 14193 31563
rect 14159 31495 14193 31508
rect 14159 31474 14193 31495
rect 14159 31427 14193 31436
rect 14159 31402 14193 31427
rect 14159 31359 14193 31364
rect 14159 31330 14193 31359
rect 9789 31116 9823 31146
rect 9789 31112 9823 31116
rect 9789 31048 9823 31074
rect 9789 31040 9823 31048
rect 9789 30980 9823 31002
rect 9789 30968 9823 30980
rect 9789 30912 9823 30930
rect 9789 30896 9823 30912
rect 9789 30844 9823 30858
rect 9789 30824 9823 30844
rect 10040 31214 10074 31218
rect 10040 31184 10074 31214
rect 10040 31112 10074 31146
rect 10040 31044 10074 31074
rect 10040 31040 10074 31044
rect 10040 30976 10074 31002
rect 10040 30968 10074 30976
rect 10040 30908 10074 30930
rect 10040 30896 10074 30908
rect 10162 31248 10196 31282
rect 10162 31173 10196 31207
rect 10162 31098 10196 31132
rect 10162 31023 10196 31057
rect 10162 30948 10196 30982
rect 10162 30874 10196 30908
rect 11018 31248 11052 31282
rect 11018 31173 11052 31207
rect 11018 31098 11052 31132
rect 11018 31023 11052 31057
rect 11018 30948 11052 30982
rect 11018 30874 11052 30908
rect 11874 31248 11908 31282
rect 11874 31173 11908 31207
rect 11874 31098 11908 31132
rect 11874 31023 11908 31057
rect 11874 30948 11908 30982
rect 11874 30874 11908 30908
rect 12730 31248 12764 31282
rect 12730 31173 12764 31207
rect 12730 31098 12764 31132
rect 12730 31023 12764 31057
rect 12730 30948 12764 30982
rect 12730 30874 12764 30908
rect 13586 31248 13620 31282
rect 13586 31173 13620 31207
rect 13586 31098 13620 31132
rect 13586 31023 13620 31057
rect 13586 30948 13620 30982
rect 13586 30874 13620 30908
rect 14042 31248 14076 31282
rect 14042 31173 14076 31207
rect 14042 31098 14076 31132
rect 14042 31023 14076 31057
rect 14042 30948 14076 30982
rect 14042 30874 14076 30908
rect 14159 31291 14193 31292
rect 14159 31258 14193 31291
rect 14159 31189 14193 31220
rect 14159 31186 14193 31189
rect 14159 31121 14193 31148
rect 14159 31114 14193 31121
rect 14159 31053 14193 31076
rect 14159 31042 14193 31053
rect 14159 30985 14193 31004
rect 14159 30970 14193 30985
rect 14159 30917 14193 30932
rect 14159 30898 14193 30917
rect 10040 30840 10074 30858
rect 10040 30824 10074 30840
rect 14159 30849 14193 30860
rect 14159 30826 14193 30849
rect 14159 30781 14193 30788
rect 14159 30754 14193 30781
rect 14159 30713 14193 30716
rect 14159 30682 14193 30713
rect 14159 30611 14193 30644
rect 14159 30610 14193 30611
rect 14159 30543 14193 30572
rect 14159 30538 14193 30543
rect 14159 30475 14193 30500
rect 14159 30466 14193 30475
rect 14159 30407 14193 30428
rect 14159 30394 14193 30407
rect 14159 30339 14193 30356
rect 14159 30322 14193 30339
rect 14159 30271 14193 30284
rect 14159 30250 14193 30271
rect 14159 30203 14193 30212
rect 14159 30178 14193 30203
rect 9789 30062 9823 30096
rect 9789 29994 9823 30024
rect 9789 29990 9823 29994
rect 9789 29926 9823 29952
rect 9789 29918 9823 29926
rect 9789 29858 9823 29880
rect 9789 29846 9823 29858
rect 9789 29790 9823 29808
rect 9789 29774 9823 29790
rect 9789 29722 9823 29736
rect 9789 29702 9823 29722
rect 10040 30092 10074 30096
rect 10040 30062 10074 30092
rect 14159 30135 14193 30140
rect 14159 30106 14193 30135
rect 14159 30067 14193 30068
rect 10040 29990 10074 30024
rect 10112 30009 10142 30043
rect 10142 30009 10146 30043
rect 10185 30009 10193 30043
rect 10193 30009 10219 30043
rect 10258 30009 10278 30043
rect 10278 30009 10292 30043
rect 10331 30009 10363 30043
rect 10363 30009 10365 30043
rect 10404 30009 10438 30043
rect 10477 30009 10482 30043
rect 10482 30009 10511 30043
rect 10550 30009 10567 30043
rect 10567 30009 10584 30043
rect 10623 30009 10652 30043
rect 10652 30009 10657 30043
rect 10696 30009 10703 30043
rect 10703 30009 10730 30043
rect 10769 30009 10788 30043
rect 10788 30009 10803 30043
rect 10842 30009 10873 30043
rect 10873 30009 10876 30043
rect 10915 30009 10949 30043
rect 10988 30009 10992 30043
rect 10992 30009 11022 30043
rect 11061 30009 11077 30043
rect 11077 30009 11095 30043
rect 11134 30009 11162 30043
rect 11162 30009 11168 30043
rect 11207 30009 11213 30043
rect 11213 30009 11241 30043
rect 11279 30009 11298 30043
rect 11298 30009 11313 30043
rect 11351 30009 11383 30043
rect 11383 30009 11385 30043
rect 11423 30009 11457 30043
rect 11495 30009 11502 30043
rect 11502 30009 11529 30043
rect 11567 30009 11587 30043
rect 11587 30009 11601 30043
rect 11639 30009 11672 30043
rect 11672 30009 11673 30043
rect 11711 30009 11723 30043
rect 11723 30009 11745 30043
rect 11783 30009 11808 30043
rect 11808 30009 11817 30043
rect 11855 30009 11889 30043
rect 11927 30009 11961 30043
rect 11999 30009 12012 30043
rect 12012 30009 12033 30043
rect 12071 30009 12097 30043
rect 12097 30009 12105 30043
rect 12143 30009 12148 30043
rect 12148 30009 12177 30043
rect 12215 30009 12233 30043
rect 12233 30009 12249 30043
rect 12287 30009 12318 30043
rect 12318 30009 12321 30043
rect 12359 30009 12393 30043
rect 12431 30009 12437 30043
rect 12437 30009 12465 30043
rect 12503 30009 12522 30043
rect 12522 30009 12537 30043
rect 12575 30009 12607 30043
rect 12607 30009 12609 30043
rect 12647 30009 12658 30043
rect 12658 30009 12681 30043
rect 12719 30009 12743 30043
rect 12743 30009 12753 30043
rect 12791 30009 12825 30043
rect 12863 30009 12897 30043
rect 12935 30009 12947 30043
rect 12947 30009 12969 30043
rect 13007 30009 13032 30043
rect 13032 30009 13041 30043
rect 13079 30009 13083 30043
rect 13083 30009 13113 30043
rect 13151 30009 13167 30043
rect 13167 30009 13185 30043
rect 13223 30009 13251 30043
rect 13251 30009 13257 30043
rect 13295 30009 13329 30043
rect 13367 30009 13369 30043
rect 13369 30009 13401 30043
rect 13439 30009 13453 30043
rect 13453 30009 13473 30043
rect 13511 30009 13537 30043
rect 13537 30009 13545 30043
rect 13583 30009 13587 30043
rect 13587 30009 13617 30043
rect 13655 30009 13671 30043
rect 13671 30009 13689 30043
rect 13727 30009 13755 30043
rect 13755 30009 13761 30043
rect 13799 30009 13833 30043
rect 13871 30009 13873 30043
rect 13873 30009 13905 30043
rect 13943 30009 13957 30043
rect 13957 30009 13977 30043
rect 14015 30009 14041 30043
rect 14041 30009 14049 30043
rect 14087 30009 14091 30043
rect 14091 30009 14121 30043
rect 14159 30034 14193 30067
rect 10040 29922 10074 29952
rect 10040 29918 10074 29922
rect 10219 29919 10223 29953
rect 10223 29919 10253 29953
rect 10304 29919 10331 29953
rect 10331 29919 10338 29953
rect 10389 29919 10405 29953
rect 10405 29919 10423 29953
rect 10474 29919 10479 29953
rect 10479 29919 10508 29953
rect 10559 29919 10592 29953
rect 10592 29919 10593 29953
rect 10643 29919 10665 29953
rect 10665 29919 10677 29953
rect 11105 29919 11113 29953
rect 11113 29919 11139 29953
rect 11178 29919 11182 29953
rect 11182 29919 11212 29953
rect 11251 29919 11285 29953
rect 11324 29919 11355 29953
rect 11355 29919 11358 29953
rect 11397 29919 11424 29953
rect 11424 29919 11431 29953
rect 11470 29919 11493 29953
rect 11493 29919 11504 29953
rect 11543 29919 11562 29953
rect 11562 29919 11577 29953
rect 11616 29919 11631 29953
rect 11631 29919 11650 29953
rect 11689 29919 11700 29953
rect 11700 29919 11723 29953
rect 11762 29919 11769 29953
rect 11769 29919 11796 29953
rect 11835 29919 11838 29953
rect 11838 29919 11869 29953
rect 11908 29919 11941 29953
rect 11941 29919 11942 29953
rect 11981 29919 12010 29953
rect 12010 29919 12015 29953
rect 12054 29919 12079 29953
rect 12079 29919 12088 29953
rect 12127 29919 12148 29953
rect 12148 29919 12161 29953
rect 12200 29919 12217 29953
rect 12217 29919 12234 29953
rect 12273 29919 12286 29953
rect 12286 29919 12307 29953
rect 12346 29919 12355 29953
rect 12355 29919 12380 29953
rect 12419 29919 12424 29953
rect 12424 29919 12453 29953
rect 12492 29919 12493 29953
rect 12493 29919 12526 29953
rect 12565 29919 12597 29953
rect 12597 29919 12599 29953
rect 12638 29919 12666 29953
rect 12666 29919 12672 29953
rect 12711 29919 12735 29953
rect 12735 29919 12745 29953
rect 12784 29919 12804 29953
rect 12804 29919 12818 29953
rect 12857 29919 12873 29953
rect 12873 29919 12891 29953
rect 12930 29919 12942 29953
rect 12942 29919 12964 29953
rect 13003 29919 13011 29953
rect 13011 29919 13037 29953
rect 13076 29919 13080 29953
rect 13080 29919 13110 29953
rect 13149 29919 13183 29953
rect 13222 29919 13252 29953
rect 13252 29919 13256 29953
rect 13295 29919 13321 29953
rect 13321 29919 13329 29953
rect 13368 29919 13390 29953
rect 13390 29919 13402 29953
rect 13441 29919 13459 29953
rect 13459 29919 13475 29953
rect 13514 29919 13528 29953
rect 13528 29919 13548 29953
rect 13587 29919 13597 29953
rect 13597 29919 13621 29953
rect 13660 29919 13666 29953
rect 13666 29919 13694 29953
rect 13733 29919 13735 29953
rect 13735 29919 13767 29953
rect 13806 29919 13840 29953
rect 13880 29919 13911 29953
rect 13911 29919 13914 29953
rect 14159 29965 14193 29996
rect 14159 29962 14193 29965
rect 10040 29854 10074 29880
rect 10040 29846 10074 29854
rect 10040 29786 10074 29808
rect 10040 29774 10074 29786
rect 10040 29718 10074 29736
rect 10040 29702 10074 29718
rect 14159 29897 14193 29924
rect 14159 29890 14193 29897
rect 14159 29829 14193 29852
rect 14159 29818 14193 29829
rect 14159 29761 14193 29780
rect 14159 29746 14193 29761
rect 14159 29693 14193 29708
rect 14159 29674 14193 29693
rect 14159 29625 14193 29636
rect 14159 29602 14193 29625
rect 14159 29557 14193 29564
rect 14159 29530 14193 29557
rect 14159 29489 14193 29492
rect 14159 29458 14193 29489
rect 14159 29387 14193 29420
rect 14159 29386 14193 29387
rect 14159 29319 14193 29348
rect 14159 29314 14193 29319
rect 14159 29251 14193 29276
rect 14159 29242 14193 29251
rect 14159 29183 14193 29204
rect 14159 29170 14193 29183
rect 14159 29115 14193 29132
rect 14159 29098 14193 29115
rect 14159 29047 14193 29060
rect 14159 29026 14193 29047
rect 10040 28902 10074 28932
rect 10040 28898 10074 28902
rect 10040 28834 10074 28860
rect 10040 28826 10074 28834
rect 10040 28766 10074 28788
rect 10040 28754 10074 28766
rect 10040 28698 10074 28716
rect 10040 28682 10074 28698
rect 10040 28630 10074 28644
rect 10040 28610 10074 28630
rect 10040 28562 10074 28572
rect 10040 28538 10074 28562
rect 10162 28944 10196 28978
rect 10162 28869 10196 28903
rect 10162 28794 10196 28828
rect 10162 28719 10196 28753
rect 10162 28644 10196 28678
rect 10162 28570 10196 28604
rect 11018 28944 11052 28978
rect 11018 28869 11052 28903
rect 11018 28794 11052 28828
rect 11018 28719 11052 28753
rect 11018 28644 11052 28678
rect 11018 28570 11052 28604
rect 11874 28944 11908 28978
rect 11874 28869 11908 28903
rect 11874 28794 11908 28828
rect 11874 28719 11908 28753
rect 11874 28644 11908 28678
rect 11874 28570 11908 28604
rect 12730 28944 12764 28978
rect 12730 28869 12764 28903
rect 12730 28794 12764 28828
rect 12730 28719 12764 28753
rect 12730 28644 12764 28678
rect 12730 28570 12764 28604
rect 13586 28944 13620 28978
rect 13586 28869 13620 28903
rect 13586 28794 13620 28828
rect 13586 28719 13620 28753
rect 13586 28644 13620 28678
rect 13586 28570 13620 28604
rect 14042 28944 14076 28978
rect 14042 28869 14076 28903
rect 14042 28794 14076 28828
rect 14042 28719 14076 28753
rect 14042 28644 14076 28678
rect 14042 28570 14076 28604
rect 14159 28979 14193 28988
rect 14159 28954 14193 28979
rect 14159 28911 14193 28916
rect 14159 28882 14193 28911
rect 14159 28843 14193 28844
rect 14159 28810 14193 28843
rect 14159 28741 14193 28772
rect 14159 28738 14193 28741
rect 14159 28673 14193 28700
rect 14159 28666 14193 28673
rect 14159 28605 14193 28628
rect 14159 28594 14193 28605
rect 10040 28494 10074 28500
rect 10040 28466 10074 28494
rect 10040 28426 10074 28428
rect 10040 28394 10074 28426
rect 10040 28324 10074 28356
rect 10040 28322 10074 28324
rect 10040 28256 10074 28284
rect 10040 28250 10074 28256
rect 10040 28188 10074 28212
rect 10040 28178 10074 28188
rect 10040 28120 10074 28140
rect 10040 28106 10074 28120
rect 10040 28052 10074 28068
rect 10040 28034 10074 28052
rect 14159 28537 14193 28556
rect 14159 28522 14193 28537
rect 14159 28469 14193 28484
rect 14159 28450 14193 28469
rect 14159 28401 14193 28412
rect 14159 28378 14193 28401
rect 14159 28333 14193 28340
rect 14159 28306 14193 28333
rect 14159 28265 14193 28268
rect 14159 28234 14193 28265
rect 14159 28163 14193 28196
rect 14159 28162 14193 28163
rect 14159 28095 14193 28124
rect 14159 28090 14193 28095
rect 14159 28027 14193 28052
rect 14159 28018 14193 28027
rect 14159 27959 14193 27980
rect 14159 27946 14193 27959
rect 14159 27891 14193 27908
rect 14159 27874 14193 27891
rect 10049 27755 10083 27789
rect 10121 27755 10142 27789
rect 10142 27755 10155 27789
rect 10193 27755 10210 27789
rect 10210 27755 10227 27789
rect 10265 27755 10278 27789
rect 10278 27755 10299 27789
rect 10337 27755 10346 27789
rect 10346 27755 10371 27789
rect 10409 27755 10414 27789
rect 10414 27755 10443 27789
rect 10481 27755 10482 27789
rect 10482 27755 10515 27789
rect 10553 27755 10584 27789
rect 10584 27755 10587 27789
rect 10625 27755 10652 27789
rect 10652 27755 10659 27789
rect 10697 27755 10720 27789
rect 10720 27755 10731 27789
rect 10769 27755 10788 27789
rect 10788 27755 10803 27789
rect 10841 27755 10856 27789
rect 10856 27755 10875 27789
rect 10913 27755 10924 27789
rect 10924 27755 10947 27789
rect 10985 27755 10992 27789
rect 10992 27755 11019 27789
rect 11057 27755 11060 27789
rect 11060 27755 11091 27789
rect 11129 27755 11162 27789
rect 11162 27755 11163 27789
rect 11201 27755 11230 27789
rect 11230 27755 11235 27789
rect 11273 27755 11298 27789
rect 11298 27755 11307 27789
rect 11345 27755 11366 27789
rect 11366 27755 11379 27789
rect 11417 27755 11434 27789
rect 11434 27755 11451 27789
rect 11489 27755 11502 27789
rect 11502 27755 11523 27789
rect 11561 27755 11570 27789
rect 11570 27755 11595 27789
rect 11633 27755 11638 27789
rect 11638 27755 11667 27789
rect 11705 27755 11706 27789
rect 11706 27755 11739 27789
rect 11777 27755 11808 27789
rect 11808 27755 11811 27789
rect 11849 27755 11876 27789
rect 11876 27755 11883 27789
rect 11921 27755 11944 27789
rect 11944 27755 11955 27789
rect 11993 27755 12012 27789
rect 12012 27755 12027 27789
rect 12065 27755 12080 27789
rect 12080 27755 12099 27789
rect 12137 27755 12148 27789
rect 12148 27755 12171 27789
rect 12209 27755 12216 27789
rect 12216 27755 12243 27789
rect 12281 27755 12284 27789
rect 12284 27755 12315 27789
rect 12353 27755 12386 27789
rect 12386 27755 12387 27789
rect 12425 27755 12454 27789
rect 12454 27755 12459 27789
rect 12497 27755 12522 27789
rect 12522 27755 12531 27789
rect 12569 27755 12590 27789
rect 12590 27755 12603 27789
rect 12641 27755 12658 27789
rect 12658 27755 12675 27789
rect 12713 27755 12726 27789
rect 12726 27755 12747 27789
rect 12785 27755 12794 27789
rect 12794 27755 12819 27789
rect 12857 27755 12862 27789
rect 12862 27755 12891 27789
rect 12929 27755 12930 27789
rect 12930 27755 12963 27789
rect 13001 27755 13032 27789
rect 13032 27755 13035 27789
rect 13073 27755 13100 27789
rect 13100 27755 13107 27789
rect 13145 27755 13168 27789
rect 13168 27755 13179 27789
rect 13217 27755 13236 27789
rect 13236 27755 13251 27789
rect 13289 27755 13304 27789
rect 13304 27755 13323 27789
rect 13361 27755 13372 27789
rect 13372 27755 13395 27789
rect 13433 27755 13440 27789
rect 13440 27755 13467 27789
rect 13505 27755 13508 27789
rect 13508 27755 13539 27789
rect 13577 27755 13610 27789
rect 13610 27755 13611 27789
rect 13649 27755 13678 27789
rect 13678 27755 13683 27789
rect 13721 27755 13746 27789
rect 13746 27755 13755 27789
rect 13793 27755 13814 27789
rect 13814 27755 13827 27789
rect 13865 27755 13882 27789
rect 13882 27755 13899 27789
rect 13937 27755 13950 27789
rect 13950 27755 13971 27789
rect 14009 27755 14018 27789
rect 14018 27755 14043 27789
rect 14081 27755 14086 27789
rect 14086 27755 14115 27789
rect 14153 27755 14187 27789
rect 14405 34540 14439 34574
rect 14405 34472 14439 34502
rect 14405 34468 14439 34472
rect 14405 34404 14439 34430
rect 14405 34396 14439 34404
rect 14405 34336 14439 34358
rect 14405 34324 14439 34336
rect 14405 34268 14439 34286
rect 14405 34252 14439 34268
rect 14405 34200 14439 34214
rect 14405 34180 14439 34200
rect 14405 34132 14439 34142
rect 14405 34108 14439 34132
rect 14405 34064 14439 34070
rect 14405 34036 14439 34064
rect 14405 33996 14439 33998
rect 14405 33964 14439 33996
rect 14405 33894 14439 33926
rect 14405 33892 14439 33894
rect 14405 33826 14439 33854
rect 14405 33820 14439 33826
rect 14405 33758 14439 33782
rect 14405 33748 14439 33758
rect 14405 33690 14439 33710
rect 14405 33676 14439 33690
rect 14405 33622 14439 33638
rect 14405 33604 14439 33622
rect 14405 33554 14439 33566
rect 14405 33532 14439 33554
rect 14405 33486 14439 33494
rect 14405 33460 14439 33486
rect 14405 33418 14439 33422
rect 14405 33388 14439 33418
rect 14405 33316 14439 33350
rect 14405 33248 14439 33278
rect 14405 33244 14439 33248
rect 14405 33180 14439 33206
rect 14405 33172 14439 33180
rect 14405 33112 14439 33134
rect 14405 33100 14439 33112
rect 14405 33044 14439 33062
rect 14405 33028 14439 33044
rect 14405 32976 14439 32990
rect 14405 32956 14439 32976
rect 14405 32908 14439 32918
rect 14405 32884 14439 32908
rect 14405 32840 14439 32846
rect 14405 32812 14439 32840
rect 14405 32772 14439 32774
rect 14405 32740 14439 32772
rect 14405 32670 14439 32702
rect 14405 32668 14439 32670
rect 14405 32602 14439 32630
rect 14405 32596 14439 32602
rect 14405 32534 14439 32558
rect 14405 32524 14439 32534
rect 14405 32466 14439 32486
rect 14405 32452 14439 32466
rect 14405 32398 14439 32414
rect 14405 32380 14439 32398
rect 14405 32330 14439 32342
rect 14405 32308 14439 32330
rect 14405 32262 14439 32270
rect 14405 32236 14439 32262
rect 14405 32194 14439 32198
rect 14405 32164 14439 32194
rect 14405 32092 14439 32126
rect 14405 32024 14439 32054
rect 14405 32020 14439 32024
rect 14405 31956 14439 31982
rect 14405 31948 14439 31956
rect 14405 31888 14439 31910
rect 14405 31876 14439 31888
rect 14405 31820 14439 31838
rect 14405 31804 14439 31820
rect 14405 31752 14439 31766
rect 14405 31732 14439 31752
rect 14405 31684 14439 31694
rect 14405 31660 14439 31684
rect 14405 31616 14439 31622
rect 14405 31588 14439 31616
rect 14405 31548 14439 31550
rect 14405 31516 14439 31548
rect 14405 31446 14439 31478
rect 14405 31444 14439 31446
rect 14405 31378 14439 31406
rect 14405 31372 14439 31378
rect 14405 31310 14439 31334
rect 14405 31300 14439 31310
rect 14405 31242 14439 31262
rect 14405 31228 14439 31242
rect 14405 31174 14439 31190
rect 14405 31156 14439 31174
rect 14405 31106 14439 31118
rect 14405 31084 14439 31106
rect 14405 31038 14439 31046
rect 14405 31012 14439 31038
rect 14405 30970 14439 30974
rect 14405 30940 14439 30970
rect 14405 30868 14439 30902
rect 14405 30800 14439 30830
rect 14405 30796 14439 30800
rect 14405 30732 14439 30758
rect 14405 30724 14439 30732
rect 14405 30664 14439 30686
rect 14405 30652 14439 30664
rect 14405 30596 14439 30614
rect 14405 30580 14439 30596
rect 14405 30528 14439 30542
rect 14405 30508 14439 30528
rect 14405 30460 14439 30470
rect 14405 30436 14439 30460
rect 14405 30392 14439 30398
rect 14405 30364 14439 30392
rect 14405 30324 14439 30326
rect 14405 30292 14439 30324
rect 14405 30222 14439 30254
rect 14405 30220 14439 30222
rect 14405 30154 14439 30182
rect 14405 30148 14439 30154
rect 14405 30086 14439 30110
rect 14405 30076 14439 30086
rect 14405 30018 14439 30038
rect 14405 30004 14439 30018
rect 14405 29950 14439 29966
rect 14405 29932 14439 29950
rect 14405 29882 14439 29894
rect 14405 29860 14439 29882
rect 14405 29814 14439 29822
rect 14405 29788 14439 29814
rect 14405 29746 14439 29750
rect 14405 29716 14439 29746
rect 14405 29644 14439 29678
rect 14405 29576 14439 29606
rect 14405 29572 14439 29576
rect 14405 29508 14439 29534
rect 14405 29500 14439 29508
rect 14405 29440 14439 29462
rect 14405 29428 14439 29440
rect 14405 29372 14439 29390
rect 14405 29356 14439 29372
rect 14405 29304 14439 29318
rect 14405 29284 14439 29304
rect 14405 29236 14439 29246
rect 14405 29212 14439 29236
rect 14405 29168 14439 29174
rect 14405 29140 14439 29168
rect 14405 29100 14439 29102
rect 14405 29068 14439 29100
rect 14405 28998 14439 29030
rect 14405 28996 14439 28998
rect 14405 28930 14439 28958
rect 14405 28924 14439 28930
rect 14405 28862 14439 28886
rect 14405 28852 14439 28862
rect 14405 28794 14439 28814
rect 14405 28780 14439 28794
rect 14405 28726 14439 28742
rect 14405 28708 14439 28726
rect 14405 28658 14439 28670
rect 14405 28636 14439 28658
rect 14405 28590 14439 28598
rect 14405 28564 14439 28590
rect 14405 28522 14439 28526
rect 14405 28492 14439 28522
rect 14405 28420 14439 28454
rect 14405 28352 14439 28382
rect 14405 28348 14439 28352
rect 14405 28284 14439 28310
rect 14405 28276 14439 28284
rect 14405 28216 14439 28238
rect 14405 28204 14439 28216
rect 14405 28148 14439 28166
rect 14405 28132 14439 28148
rect 14405 28080 14439 28094
rect 14405 28060 14439 28080
rect 14405 28012 14439 28022
rect 14405 27988 14439 28012
rect 14405 27944 14439 27950
rect 14405 27916 14439 27944
rect 14405 27876 14439 27878
rect 14405 27844 14439 27876
rect 14405 27774 14439 27806
rect 14405 27772 14439 27774
rect 14405 27706 14439 27734
rect 14405 27700 14439 27706
rect 14405 27638 14439 27662
rect 14405 27628 14439 27638
rect 9789 27478 9823 27490
rect 9789 27456 9823 27478
rect 11960 27482 11994 27516
rect 12059 27482 12093 27516
rect 12157 27482 12191 27516
rect 12432 27496 12466 27530
rect 12510 27502 12534 27536
rect 12534 27502 12544 27536
rect 12582 27502 12602 27536
rect 12602 27502 12616 27536
rect 12654 27502 12670 27536
rect 12670 27502 12688 27536
rect 12726 27502 12738 27536
rect 12738 27502 12760 27536
rect 12798 27502 12806 27536
rect 12806 27502 12832 27536
rect 12870 27502 12874 27536
rect 12874 27502 12904 27536
rect 12942 27502 12976 27536
rect 13014 27502 13044 27536
rect 13044 27502 13048 27536
rect 13086 27502 13112 27536
rect 13112 27502 13120 27536
rect 13158 27502 13180 27536
rect 13180 27502 13192 27536
rect 13230 27502 13248 27536
rect 13248 27502 13264 27536
rect 13302 27502 13316 27536
rect 13316 27502 13336 27536
rect 13374 27502 13384 27536
rect 13384 27502 13408 27536
rect 13446 27502 13452 27536
rect 13452 27502 13480 27536
rect 13518 27502 13520 27536
rect 13520 27502 13552 27536
rect 13590 27502 13622 27536
rect 13622 27502 13624 27536
rect 13662 27502 13690 27536
rect 13690 27502 13696 27536
rect 13734 27502 13758 27536
rect 13758 27502 13768 27536
rect 13806 27502 13826 27536
rect 13826 27502 13840 27536
rect 13878 27502 13894 27536
rect 13894 27502 13912 27536
rect 13950 27502 13962 27536
rect 13962 27502 13984 27536
rect 14022 27502 14030 27536
rect 14030 27502 14056 27536
rect 14094 27502 14098 27536
rect 14098 27502 14128 27536
rect 14183 27502 14200 27536
rect 14200 27502 14217 27536
rect 14255 27502 14268 27536
rect 14268 27502 14289 27536
rect 14327 27502 14336 27536
rect 14336 27502 14361 27536
rect 14399 27502 14433 27536
rect 9789 27410 9823 27418
rect 9789 27384 9823 27410
rect 9789 27342 9823 27346
rect 9789 27312 9823 27342
rect 9789 27240 9823 27274
rect 9789 27172 9823 27202
rect 9789 27168 9823 27172
rect 9789 27104 9823 27130
rect 9789 27096 9823 27104
rect 9789 27036 9823 27058
rect 9789 27024 9823 27036
rect 9789 26968 9823 26986
rect 9789 26952 9823 26968
rect 9789 26900 9823 26914
rect 9789 26880 9823 26900
rect 9789 26832 9823 26842
rect 9789 26808 9823 26832
rect 9789 26764 9823 26770
rect 9789 26736 9823 26764
rect 9789 26696 9823 26698
rect 9789 26664 9823 26696
rect 10105 27129 10139 27158
rect 10105 27124 10139 27129
rect 10105 27056 10139 27086
rect 10105 27052 10139 27056
rect 12432 27424 12466 27458
rect 12432 27356 12466 27386
rect 12432 27352 12466 27356
rect 12432 27288 12466 27314
rect 12432 27280 12466 27288
rect 12432 27220 12466 27242
rect 12432 27208 12466 27220
rect 12432 27152 12466 27170
rect 12432 27136 12466 27152
rect 12432 27084 12466 27098
rect 12432 27064 12466 27084
rect 12432 27016 12466 27026
rect 12432 26992 12466 27016
rect 12432 26948 12466 26954
rect 12432 26920 12466 26948
rect 12432 26880 12466 26882
rect 12432 26848 12466 26880
rect 12432 26778 12466 26810
rect 12432 26776 12466 26778
rect 12432 26710 12466 26738
rect 12432 26704 12466 26710
rect 11960 26626 11994 26660
rect 12059 26626 12093 26660
rect 12157 26626 12191 26660
rect 12432 26642 12466 26666
rect 12432 26632 12466 26642
rect 9789 26594 9823 26626
rect 9789 26592 9823 26594
rect 9789 26526 9823 26554
rect 9789 26520 9823 26526
rect 9789 26448 9823 26482
rect 12432 26574 12466 26594
rect 12432 26560 12466 26574
rect 12432 26506 12466 26522
rect 12432 26488 12466 26506
rect 9789 26376 9823 26410
rect 9906 26370 9925 26404
rect 9925 26370 9940 26404
rect 9978 26370 9993 26404
rect 9993 26370 10012 26404
rect 10050 26370 10061 26404
rect 10061 26370 10084 26404
rect 10122 26370 10129 26404
rect 10129 26370 10156 26404
rect 10194 26370 10197 26404
rect 10197 26370 10228 26404
rect 10266 26370 10299 26404
rect 10299 26370 10300 26404
rect 10338 26370 10367 26404
rect 10367 26370 10372 26404
rect 10410 26370 10435 26404
rect 10435 26370 10444 26404
rect 10482 26370 10503 26404
rect 10503 26370 10516 26404
rect 10554 26370 10571 26404
rect 10571 26370 10588 26404
rect 10626 26370 10639 26404
rect 10639 26370 10660 26404
rect 10698 26370 10707 26404
rect 10707 26370 10732 26404
rect 10770 26370 10775 26404
rect 10775 26370 10804 26404
rect 10842 26370 10843 26404
rect 10843 26370 10876 26404
rect 10914 26370 10945 26404
rect 10945 26370 10948 26404
rect 10986 26370 11013 26404
rect 11013 26370 11020 26404
rect 11058 26370 11081 26404
rect 11081 26370 11092 26404
rect 11130 26370 11149 26404
rect 11149 26370 11164 26404
rect 11202 26370 11217 26404
rect 11217 26370 11236 26404
rect 11274 26370 11285 26404
rect 11285 26370 11308 26404
rect 11346 26370 11353 26404
rect 11353 26370 11380 26404
rect 11418 26370 11421 26404
rect 11421 26370 11452 26404
rect 11490 26370 11523 26404
rect 11523 26370 11524 26404
rect 11562 26370 11591 26404
rect 11591 26370 11596 26404
rect 11634 26370 11659 26404
rect 11659 26370 11668 26404
rect 11706 26370 11727 26404
rect 11727 26370 11740 26404
rect 11778 26370 11795 26404
rect 11795 26370 11812 26404
rect 11850 26370 11863 26404
rect 11863 26370 11884 26404
rect 11922 26370 11931 26404
rect 11931 26370 11956 26404
rect 11994 26370 11999 26404
rect 11999 26370 12028 26404
rect 12066 26370 12067 26404
rect 12067 26370 12100 26404
rect 12138 26370 12169 26404
rect 12169 26370 12172 26404
rect 12210 26370 12237 26404
rect 12237 26370 12244 26404
rect 12282 26370 12305 26404
rect 12305 26370 12316 26404
rect 12354 26370 12388 26404
rect 12426 26370 12460 26404
rect 130 17155 164 17189
rect 130 17083 164 17117
rect 130 17011 164 17045
rect 212 17161 246 17195
rect 284 17161 318 17195
rect 488 17161 522 17195
rect 560 17161 594 17195
rect 836 17161 870 17195
rect 908 17161 942 17195
rect 130 16939 164 16973
rect 261 16874 268 16908
rect 268 16874 295 16908
rect 333 16874 336 16908
rect 336 16874 367 16908
rect 404 16801 438 16835
rect 404 16729 438 16763
rect 560 16744 594 16778
rect 632 16744 666 16778
rect 704 16744 738 16778
rect 776 16744 810 16778
rect 944 16744 978 16778
rect 1016 16744 1050 16778
rect 1088 16744 1122 16778
rect 1160 16744 1194 16778
rect 1472 16744 1506 16778
rect 1544 16744 1578 16778
rect 1616 16744 1650 16778
rect 1688 16744 1722 16778
rect 1856 16744 1890 16778
rect 1928 16744 1962 16778
rect 2000 16744 2034 16778
rect 2072 16744 2106 16778
rect 2930 16744 2964 16778
rect 3002 16744 3036 16778
rect 3074 16744 3108 16778
rect 3146 16744 3180 16778
rect 3314 16744 3348 16778
rect 3386 16744 3420 16778
rect 3458 16744 3492 16778
rect 3530 16744 3564 16778
rect 3842 16744 3876 16778
rect 3914 16744 3948 16778
rect 3986 16744 4020 16778
rect 4058 16744 4092 16778
rect 4226 16744 4260 16778
rect 4298 16744 4332 16778
rect 4370 16744 4404 16778
rect 4442 16744 4476 16778
rect 488 13729 496 13763
rect 496 13729 522 13763
rect 560 13729 564 13763
rect 564 13729 594 13763
rect 632 13729 666 13763
rect 704 13729 734 13763
rect 734 13729 738 13763
rect 776 13729 802 13763
rect 802 13729 810 13763
rect 944 13729 952 13763
rect 952 13729 978 13763
rect 1016 13729 1020 13763
rect 1020 13729 1050 13763
rect 1088 13729 1122 13763
rect 1160 13729 1190 13763
rect 1190 13729 1194 13763
rect 1232 13729 1258 13763
rect 1258 13729 1266 13763
rect 1400 13729 1408 13763
rect 1408 13729 1434 13763
rect 1472 13729 1476 13763
rect 1476 13729 1506 13763
rect 1544 13729 1578 13763
rect 1616 13729 1646 13763
rect 1646 13729 1650 13763
rect 1688 13729 1714 13763
rect 1714 13729 1722 13763
rect 1856 13729 1864 13763
rect 1864 13729 1890 13763
rect 1928 13729 1932 13763
rect 1932 13729 1962 13763
rect 2000 13729 2034 13763
rect 2072 13729 2102 13763
rect 2102 13729 2106 13763
rect 2144 13729 2170 13763
rect 2170 13729 2178 13763
rect 2858 13729 2866 13763
rect 2866 13729 2892 13763
rect 2930 13729 2934 13763
rect 2934 13729 2964 13763
rect 3002 13729 3036 13763
rect 3074 13729 3104 13763
rect 3104 13729 3108 13763
rect 3146 13729 3172 13763
rect 3172 13729 3180 13763
rect 3314 13729 3322 13763
rect 3322 13729 3348 13763
rect 3386 13729 3390 13763
rect 3390 13729 3420 13763
rect 3458 13729 3492 13763
rect 3530 13729 3560 13763
rect 3560 13729 3564 13763
rect 3602 13729 3628 13763
rect 3628 13729 3636 13763
rect 3770 13729 3778 13763
rect 3778 13729 3804 13763
rect 3842 13729 3846 13763
rect 3846 13729 3876 13763
rect 3914 13729 3948 13763
rect 3986 13729 4016 13763
rect 4016 13729 4020 13763
rect 4058 13729 4084 13763
rect 4084 13729 4092 13763
rect 4226 13729 4234 13763
rect 4234 13729 4260 13763
rect 4298 13729 4302 13763
rect 4302 13729 4332 13763
rect 4370 13729 4404 13763
rect 4442 13729 4472 13763
rect 4472 13729 4476 13763
rect 4514 13729 4540 13763
rect 4540 13729 4548 13763
rect 3230 13625 3264 13659
rect 3230 13550 3264 13584
rect 3230 13474 3264 13508
rect 3230 13398 3264 13432
rect 3230 13322 3264 13356
rect 3230 13246 3264 13280
rect 3230 13170 3264 13204
rect 3230 13094 3264 13128
rect 3230 13018 3264 13052
rect 3230 12942 3264 12976
rect 3230 12866 3264 12900
rect 3230 12790 3264 12824
rect 3230 12714 3264 12748
rect 3230 12638 3264 12672
rect 3230 12562 3264 12596
rect 3230 12486 3264 12520
rect 3230 12410 3264 12444
rect 3230 12334 3264 12368
rect 488 12199 496 12233
rect 496 12199 522 12233
rect 560 12199 564 12233
rect 564 12199 594 12233
rect 632 12199 666 12233
rect 704 12199 734 12233
rect 734 12199 738 12233
rect 776 12199 802 12233
rect 802 12199 810 12233
rect 944 12199 952 12233
rect 952 12199 978 12233
rect 1016 12199 1020 12233
rect 1020 12199 1050 12233
rect 1088 12199 1122 12233
rect 1160 12199 1190 12233
rect 1190 12199 1194 12233
rect 1232 12199 1258 12233
rect 1258 12199 1266 12233
rect 1400 12199 1408 12233
rect 1408 12199 1434 12233
rect 1472 12199 1476 12233
rect 1476 12199 1506 12233
rect 1544 12199 1578 12233
rect 1616 12199 1646 12233
rect 1646 12199 1650 12233
rect 1688 12199 1714 12233
rect 1714 12199 1722 12233
rect 1856 12199 1864 12233
rect 1864 12199 1890 12233
rect 1928 12199 1932 12233
rect 1932 12199 1962 12233
rect 2000 12199 2034 12233
rect 2072 12199 2102 12233
rect 2102 12199 2106 12233
rect 2144 12199 2170 12233
rect 2170 12199 2178 12233
rect 2858 12199 2866 12233
rect 2866 12199 2892 12233
rect 2930 12199 2934 12233
rect 2934 12199 2964 12233
rect 3002 12199 3036 12233
rect 3074 12199 3104 12233
rect 3104 12199 3108 12233
rect 3146 12199 3172 12233
rect 3172 12199 3180 12233
rect 3314 12199 3322 12233
rect 3322 12199 3348 12233
rect 3386 12199 3390 12233
rect 3390 12199 3420 12233
rect 3458 12199 3492 12233
rect 3530 12199 3560 12233
rect 3560 12199 3564 12233
rect 3602 12199 3628 12233
rect 3628 12199 3636 12233
rect 3770 12199 3778 12233
rect 3778 12199 3804 12233
rect 3842 12199 3846 12233
rect 3846 12199 3876 12233
rect 3914 12199 3948 12233
rect 3986 12199 4016 12233
rect 4016 12199 4020 12233
rect 4058 12199 4084 12233
rect 4084 12199 4092 12233
rect 4226 12199 4234 12233
rect 4234 12199 4260 12233
rect 4298 12199 4302 12233
rect 4302 12199 4332 12233
rect 4370 12199 4404 12233
rect 4442 12199 4472 12233
rect 4472 12199 4476 12233
rect 4514 12199 4540 12233
rect 4540 12199 4548 12233
rect 179 12114 213 12148
rect 251 12114 285 12148
rect 323 12114 325 12148
rect 325 12114 357 12148
rect 395 12114 427 12148
rect 427 12114 429 12148
rect 467 12114 495 12148
rect 495 12114 501 12148
rect 2429 12114 2433 12148
rect 2433 12114 2463 12148
rect 2501 12147 2535 12148
rect 2501 12114 2535 12147
rect 2573 12114 2596 12148
rect 2596 12114 2607 12148
rect 5248 15730 5282 15732
rect 5320 15730 5354 15732
rect 5392 15730 5426 15732
rect 5464 15730 5498 15732
rect 5248 15698 5254 15730
rect 5254 15698 5282 15730
rect 5320 15698 5322 15730
rect 5322 15698 5354 15730
rect 5392 15698 5424 15730
rect 5424 15698 5426 15730
rect 5464 15698 5492 15730
rect 5492 15698 5498 15730
rect 5180 15546 5214 15580
rect 5180 15474 5214 15508
rect 5180 15402 5214 15436
rect 5180 15330 5214 15364
rect 5180 15258 5214 15292
rect 5180 15186 5214 15220
rect 5180 15114 5214 15148
rect 5356 15546 5390 15580
rect 5356 15463 5390 15497
rect 5356 15380 5390 15414
rect 5356 15297 5390 15331
rect 5356 15214 5390 15248
rect 5356 15130 5390 15164
rect 5532 15546 5566 15580
rect 5532 15474 5566 15508
rect 5532 15402 5566 15436
rect 5532 15330 5566 15364
rect 5532 15258 5566 15292
rect 5532 15186 5566 15220
rect 5532 15114 5566 15148
rect 5192 14741 5226 14743
rect 5192 14709 5226 14741
rect 5192 14637 5226 14671
rect 5612 14627 5646 14661
rect 5612 14555 5646 14589
rect 5756 14627 5790 14661
rect 5756 14555 5790 14589
rect 5892 14627 5926 14661
rect 5892 14555 5926 14589
rect 6036 14627 6070 14661
rect 6036 14555 6070 14589
rect 6172 14626 6206 14660
rect 6172 14554 6206 14588
rect 5332 13874 5366 13876
rect 5332 13842 5366 13874
rect 5332 13770 5366 13804
rect 5476 13874 5510 13876
rect 5476 13842 5506 13874
rect 5506 13842 5510 13874
rect 5476 13770 5510 13804
rect 866 11971 897 12005
rect 897 11971 900 12005
rect 938 11971 965 12005
rect 965 11971 972 12005
rect 1097 11971 1099 12005
rect 1099 11971 1131 12005
rect 1169 11971 1201 12005
rect 1201 11971 1203 12005
rect 1333 11971 1335 12005
rect 1335 11971 1367 12005
rect 1405 11971 1437 12005
rect 1437 11971 1439 12005
rect 1569 11971 1571 12005
rect 1571 11971 1603 12005
rect 1641 11971 1673 12005
rect 1673 11971 1675 12005
rect 1805 11971 1807 12005
rect 1807 11971 1839 12005
rect 1877 11971 1909 12005
rect 1909 11971 1911 12005
rect 2041 11971 2043 12005
rect 2043 11971 2075 12005
rect 2113 11971 2145 12005
rect 2145 11971 2147 12005
rect 2889 11971 2891 12005
rect 2891 11971 2923 12005
rect 2961 11971 2993 12005
rect 2993 11971 2995 12005
rect 3125 11971 3127 12005
rect 3127 11971 3159 12005
rect 3197 11971 3229 12005
rect 3229 11971 3231 12005
rect 3361 11971 3363 12005
rect 3363 11971 3395 12005
rect 3433 11971 3465 12005
rect 3465 11971 3467 12005
rect 3597 11971 3599 12005
rect 3599 11971 3631 12005
rect 3669 11971 3701 12005
rect 3701 11971 3703 12005
rect 3833 11971 3835 12005
rect 3835 11971 3867 12005
rect 3905 11971 3937 12005
rect 3937 11971 3939 12005
rect 4064 11971 4071 12005
rect 4071 11971 4098 12005
rect 4136 11971 4139 12005
rect 4139 11971 4170 12005
rect 569 9845 603 9879
rect 2405 9985 2439 10019
rect 2405 9913 2439 9947
rect 569 9773 603 9807
rect 2597 9985 2631 10019
rect 2597 9913 2631 9947
rect 5332 10347 5366 10381
rect 5192 10265 5226 10299
rect 5332 10275 5366 10309
rect 5192 10195 5226 10227
rect 5472 10347 5506 10381
rect 5472 10275 5506 10309
rect 5616 10347 5650 10381
rect 5616 10275 5650 10309
rect 5752 10347 5786 10381
rect 5752 10275 5786 10309
rect 5896 10347 5930 10381
rect 5896 10275 5930 10309
rect 6032 10347 6066 10381
rect 6032 10275 6066 10309
rect 6172 10347 6206 10381
rect 6172 10275 6206 10309
rect 5192 10193 5226 10195
rect 4433 10002 4467 10036
rect 4433 9930 4467 9964
rect 548 9604 582 9638
rect 620 9604 654 9638
rect 2354 9604 2388 9638
rect 2426 9604 2460 9638
rect 2576 9604 2610 9638
rect 2648 9604 2682 9638
rect 4382 9604 4416 9638
rect 4454 9604 4488 9638
rect 546 9511 580 9544
rect 546 9510 574 9511
rect 574 9510 580 9511
rect 618 9510 632 9544
rect 632 9510 652 9544
rect 690 9510 700 9544
rect 700 9510 724 9544
rect 762 9510 768 9544
rect 768 9510 796 9544
rect 834 9510 836 9544
rect 836 9510 868 9544
rect 906 9510 938 9544
rect 938 9510 940 9544
rect 978 9510 1006 9544
rect 1006 9510 1012 9544
rect 4036 9510 4038 9544
rect 4038 9510 4070 9544
rect 4108 9510 4140 9544
rect 4140 9510 4142 9544
rect 4180 9510 4208 9544
rect 4208 9510 4214 9544
rect 4252 9510 4276 9544
rect 4276 9510 4286 9544
rect 4324 9510 4344 9544
rect 4344 9510 4358 9544
rect 4396 9510 4412 9544
rect 4412 9510 4430 9544
rect 4468 9510 4480 9544
rect 4480 9510 4502 9544
rect 4658 9510 4684 9544
rect 4684 9510 4692 9544
rect 4730 9510 4752 9544
rect 4752 9510 4764 9544
rect 4802 9510 4820 9544
rect 4820 9510 4836 9544
rect 4874 9510 4888 9544
rect 4888 9510 4908 9544
rect 4946 9510 4956 9544
rect 4956 9510 4980 9544
rect 5113 9510 5126 9544
rect 5126 9510 5147 9544
rect 5185 9510 5194 9544
rect 5194 9510 5219 9544
rect 5257 9510 5262 9544
rect 5262 9510 5291 9544
rect 5329 9510 5330 9544
rect 5330 9510 5363 9544
rect 5401 9510 5432 9544
rect 5432 9510 5435 9544
rect 5608 9510 5636 9544
rect 5636 9510 5642 9544
rect 5680 9510 5704 9544
rect 5704 9510 5714 9544
rect 5752 9510 5772 9544
rect 5772 9510 5786 9544
rect 5824 9510 5858 9544
rect 4501 9425 4505 9459
rect 4505 9425 4535 9459
rect 4573 9425 4607 9459
rect 4645 9425 4675 9459
rect 4675 9425 4679 9459
rect 4957 9425 4961 9459
rect 4961 9425 4991 9459
rect 5029 9425 5063 9459
rect 5101 9425 5131 9459
rect 5131 9425 5135 9459
rect 5413 9425 5417 9459
rect 5417 9425 5447 9459
rect 5485 9425 5519 9459
rect 5557 9425 5587 9459
rect 5587 9425 5591 9459
rect 657 7253 691 7287
rect 729 7253 741 7287
rect 741 7253 763 7287
rect 801 7253 825 7287
rect 825 7253 835 7287
rect 873 7253 907 7287
rect 1049 7252 1051 7286
rect 1051 7252 1083 7286
rect 1121 7252 1153 7286
rect 1153 7252 1155 7286
rect 1297 7253 1331 7287
rect 1369 7253 1379 7287
rect 1379 7253 1403 7287
rect 1441 7253 1463 7287
rect 1463 7253 1475 7287
rect 1513 7253 1547 7287
rect 1585 7253 1597 7287
rect 1597 7253 1619 7287
rect 1657 7253 1681 7287
rect 1681 7253 1691 7287
rect 1729 7253 1763 7287
rect 1905 7252 1907 7286
rect 1907 7252 1939 7286
rect 1977 7252 2009 7286
rect 2009 7252 2011 7286
rect 2153 7253 2187 7287
rect 2225 7253 2235 7287
rect 2235 7253 2259 7287
rect 2297 7253 2319 7287
rect 2319 7253 2331 7287
rect 2369 7253 2403 7287
rect 2441 7253 2453 7287
rect 2453 7253 2475 7287
rect 2513 7253 2537 7287
rect 2537 7253 2547 7287
rect 2585 7253 2619 7287
rect 2761 7252 2763 7286
rect 2763 7252 2795 7286
rect 2833 7252 2865 7286
rect 2865 7252 2867 7286
rect 3009 7253 3043 7287
rect 3081 7253 3091 7287
rect 3091 7253 3115 7287
rect 3153 7253 3175 7287
rect 3175 7253 3187 7287
rect 3225 7253 3259 7287
rect 3489 7253 3523 7287
rect 3561 7253 3573 7287
rect 3573 7253 3595 7287
rect 3633 7253 3657 7287
rect 3657 7253 3667 7287
rect 3705 7253 3739 7287
rect 3881 7252 3883 7286
rect 3883 7252 3915 7286
rect 3953 7252 3985 7286
rect 3985 7252 3987 7286
rect 4129 7253 4163 7287
rect 4201 7253 4211 7287
rect 4211 7253 4235 7287
rect 4273 7253 4295 7287
rect 4295 7253 4307 7287
rect 4345 7253 4379 7287
rect 4537 7252 4539 7286
rect 4539 7252 4571 7286
rect 4609 7252 4641 7286
rect 4641 7252 4643 7286
rect 4765 7253 4799 7287
rect 4837 7253 4871 7287
rect 4993 7252 4995 7286
rect 4995 7252 5027 7286
rect 5065 7252 5097 7286
rect 5097 7252 5099 7286
rect 5221 7253 5255 7287
rect 5293 7253 5327 7287
rect 5449 7252 5451 7286
rect 5451 7252 5483 7286
rect 5521 7252 5553 7286
rect 5553 7252 5555 7286
rect 5713 7253 5747 7287
rect 657 5033 691 5067
rect 729 5033 741 5067
rect 741 5033 763 5067
rect 801 5033 825 5067
rect 825 5033 835 5067
rect 873 5033 907 5067
rect 1049 5032 1051 5066
rect 1051 5032 1083 5066
rect 1121 5032 1153 5066
rect 1153 5032 1155 5066
rect 1297 5033 1331 5067
rect 1369 5033 1379 5067
rect 1379 5033 1403 5067
rect 1441 5033 1463 5067
rect 1463 5033 1475 5067
rect 1513 5033 1547 5067
rect 1585 5033 1597 5067
rect 1597 5033 1619 5067
rect 1657 5033 1681 5067
rect 1681 5033 1691 5067
rect 1729 5033 1763 5067
rect 1905 5032 1907 5066
rect 1907 5032 1939 5066
rect 1977 5032 2009 5066
rect 2009 5032 2011 5066
rect 2153 5033 2187 5067
rect 2225 5033 2235 5067
rect 2235 5033 2259 5067
rect 2297 5033 2319 5067
rect 2319 5033 2331 5067
rect 2369 5033 2403 5067
rect 2441 5033 2453 5067
rect 2453 5033 2475 5067
rect 2513 5033 2537 5067
rect 2537 5033 2547 5067
rect 2585 5033 2619 5067
rect 2761 5032 2763 5066
rect 2763 5032 2795 5066
rect 2833 5032 2865 5066
rect 2865 5032 2867 5066
rect 3009 5033 3043 5067
rect 3081 5033 3091 5067
rect 3091 5033 3115 5067
rect 3153 5033 3175 5067
rect 3175 5033 3187 5067
rect 3225 5033 3259 5067
rect 3489 5033 3523 5067
rect 3561 5033 3573 5067
rect 3573 5033 3595 5067
rect 3633 5033 3657 5067
rect 3657 5033 3667 5067
rect 3705 5033 3739 5067
rect 3881 5032 3883 5066
rect 3883 5032 3915 5066
rect 3953 5032 3985 5066
rect 3985 5032 3987 5066
rect 4129 5033 4163 5067
rect 4201 5033 4211 5067
rect 4211 5033 4235 5067
rect 4273 5033 4295 5067
rect 4295 5033 4307 5067
rect 4345 5033 4379 5067
rect 4537 5032 4539 5066
rect 4539 5032 4571 5066
rect 4609 5032 4641 5066
rect 4641 5032 4643 5066
rect 4765 5033 4799 5067
rect 4837 5033 4871 5067
rect 4993 5032 4995 5066
rect 4995 5032 5027 5066
rect 5065 5032 5097 5066
rect 5097 5032 5099 5066
rect 5221 5033 5255 5067
rect 5293 5033 5327 5067
rect 5449 5032 5451 5066
rect 5451 5032 5483 5066
rect 5521 5032 5553 5066
rect 5553 5032 5555 5066
rect 5713 5033 5747 5067
rect 657 2814 691 2848
rect 729 2814 741 2848
rect 741 2814 763 2848
rect 801 2814 825 2848
rect 825 2814 835 2848
rect 873 2814 907 2848
rect 1049 2813 1051 2847
rect 1051 2813 1083 2847
rect 1121 2813 1153 2847
rect 1153 2813 1155 2847
rect 1297 2814 1331 2848
rect 1369 2814 1379 2848
rect 1379 2814 1403 2848
rect 1441 2814 1463 2848
rect 1463 2814 1475 2848
rect 1513 2814 1547 2848
rect 1585 2814 1597 2848
rect 1597 2814 1619 2848
rect 1657 2814 1681 2848
rect 1681 2814 1691 2848
rect 1729 2814 1763 2848
rect 1905 2813 1907 2847
rect 1907 2813 1939 2847
rect 1977 2813 2009 2847
rect 2009 2813 2011 2847
rect 2153 2814 2187 2848
rect 2225 2814 2235 2848
rect 2235 2814 2259 2848
rect 2297 2814 2319 2848
rect 2319 2814 2331 2848
rect 2369 2814 2403 2848
rect 2441 2814 2453 2848
rect 2453 2814 2475 2848
rect 2513 2814 2537 2848
rect 2537 2814 2547 2848
rect 2585 2814 2619 2848
rect 2761 2813 2763 2847
rect 2763 2813 2795 2847
rect 2833 2813 2865 2847
rect 2865 2813 2867 2847
rect 3009 2814 3043 2848
rect 3081 2814 3091 2848
rect 3091 2814 3115 2848
rect 3153 2814 3175 2848
rect 3175 2814 3187 2848
rect 3225 2814 3259 2848
rect 3489 2814 3523 2848
rect 3561 2814 3573 2848
rect 3573 2814 3595 2848
rect 3633 2814 3657 2848
rect 3657 2814 3667 2848
rect 3705 2814 3739 2848
rect 3881 2813 3883 2847
rect 3883 2813 3915 2847
rect 3953 2813 3985 2847
rect 3985 2813 3987 2847
rect 4129 2814 4163 2848
rect 4201 2814 4211 2848
rect 4211 2814 4235 2848
rect 4273 2814 4295 2848
rect 4295 2814 4307 2848
rect 4345 2814 4379 2848
rect 4537 2813 4539 2847
rect 4539 2813 4571 2847
rect 4609 2813 4641 2847
rect 4641 2813 4643 2847
rect 4765 2814 4799 2848
rect 4837 2814 4871 2848
rect 4993 2813 4995 2847
rect 4995 2813 5027 2847
rect 5065 2813 5097 2847
rect 5097 2813 5099 2847
rect 5221 2815 5255 2849
rect 5293 2815 5327 2849
rect 5449 2813 5451 2847
rect 5451 2813 5483 2847
rect 5521 2813 5553 2847
rect 5553 2813 5555 2847
rect 5713 2814 5747 2848
rect 618 557 641 591
rect 641 557 652 591
rect 690 557 709 591
rect 709 557 724 591
rect 762 557 777 591
rect 777 557 796 591
rect 834 557 845 591
rect 845 557 868 591
rect 906 557 913 591
rect 913 557 940 591
rect 978 557 1012 591
rect 1055 467 1089 501
rect 1127 467 1161 501
rect 2011 467 2045 501
rect 2083 467 2117 501
rect 4501 642 4505 676
rect 4505 642 4535 676
rect 4573 642 4607 676
rect 4645 642 4675 676
rect 4675 642 4679 676
rect 4957 642 4961 676
rect 4961 642 4991 676
rect 5029 642 5063 676
rect 5101 642 5131 676
rect 5131 642 5135 676
rect 5413 642 5417 676
rect 5417 642 5447 676
rect 5485 642 5519 676
rect 5557 642 5587 676
rect 5587 642 5591 676
rect 2933 467 2967 501
rect 3005 467 3039 501
rect 3907 557 3941 591
rect 3979 557 4013 591
rect 4051 557 4081 591
rect 4081 557 4085 591
rect 4123 557 4149 591
rect 4149 557 4157 591
rect 4195 557 4217 591
rect 4217 557 4229 591
rect 4267 557 4285 591
rect 4285 557 4301 591
rect 4339 557 4353 591
rect 4353 557 4373 591
rect 3746 467 3780 501
rect 3818 467 3852 501
rect 4575 557 4609 591
rect 4647 557 4673 591
rect 4673 557 4681 591
rect 4719 557 4741 591
rect 4741 557 4753 591
rect 4791 557 4809 591
rect 4809 557 4825 591
rect 4421 467 4455 501
rect 4493 467 4527 501
rect 5047 557 5081 591
rect 5119 557 5143 591
rect 5143 557 5153 591
rect 5191 557 5211 591
rect 5211 557 5225 591
rect 4877 467 4911 501
rect 4949 467 4983 501
rect 5446 557 5457 591
rect 5457 557 5480 591
rect 5518 557 5525 591
rect 5525 557 5552 591
rect 5590 557 5593 591
rect 5593 557 5624 591
rect 5662 557 5695 591
rect 5695 557 5696 591
rect 5734 557 5763 591
rect 5763 557 5768 591
rect 5279 467 5313 501
rect 5351 467 5385 501
<< metal1 >>
rect 9783 34796 14445 34802
rect 9783 34762 9795 34796
rect 9829 34762 9867 34796
rect 9901 34762 9939 34796
rect 9973 34762 10011 34796
rect 10045 34762 10083 34796
rect 10117 34762 10155 34796
rect 10189 34762 10227 34796
rect 10261 34762 10299 34796
rect 10333 34762 10371 34796
rect 10405 34762 10443 34796
rect 10477 34762 10515 34796
rect 10549 34762 10587 34796
rect 10621 34762 10659 34796
rect 10693 34762 10731 34796
rect 10765 34762 10803 34796
rect 10837 34762 10875 34796
rect 10909 34762 10947 34796
rect 10981 34762 11019 34796
rect 11053 34762 11091 34796
rect 11125 34762 11163 34796
rect 11197 34762 11235 34796
rect 11269 34762 11307 34796
rect 11341 34762 11379 34796
rect 11413 34762 11451 34796
rect 11485 34762 11523 34796
rect 11557 34762 11595 34796
rect 11629 34762 11667 34796
rect 11701 34762 11739 34796
rect 11773 34762 11811 34796
rect 11845 34762 11883 34796
rect 11917 34762 11955 34796
rect 11989 34762 12027 34796
rect 12061 34762 12099 34796
rect 12133 34762 12171 34796
rect 12205 34762 12243 34796
rect 12277 34762 12315 34796
rect 12349 34762 12387 34796
rect 12421 34762 12459 34796
rect 12493 34762 12531 34796
rect 12565 34762 12603 34796
rect 12637 34762 12675 34796
rect 12709 34762 12747 34796
rect 12781 34762 12819 34796
rect 12853 34762 12891 34796
rect 12925 34762 12963 34796
rect 12997 34762 13035 34796
rect 13069 34762 13107 34796
rect 13141 34762 13179 34796
rect 13213 34762 13251 34796
rect 13285 34762 13323 34796
rect 13357 34762 13395 34796
rect 13429 34762 13467 34796
rect 13501 34762 13539 34796
rect 13573 34762 13611 34796
rect 13645 34762 13683 34796
rect 13717 34762 13755 34796
rect 13789 34762 13827 34796
rect 13861 34762 13899 34796
rect 13933 34762 13971 34796
rect 14005 34762 14043 34796
rect 14077 34762 14115 34796
rect 14149 34762 14187 34796
rect 14221 34762 14259 34796
rect 14293 34762 14331 34796
rect 14365 34790 14445 34796
rect 14365 34762 14405 34790
rect 9783 34756 14405 34762
rect 14439 34756 14445 34790
rect 9783 34708 9829 34756
rect 9783 34674 9789 34708
rect 9823 34674 9829 34708
rect 9783 34636 9829 34674
rect 9783 34602 9789 34636
rect 9823 34602 9829 34636
rect 9783 34564 9829 34602
rect 9783 34530 9789 34564
rect 9823 34530 9829 34564
rect 14399 34718 14445 34756
rect 14399 34684 14405 34718
rect 14439 34684 14445 34718
rect 14399 34646 14445 34684
rect 14399 34612 14405 34646
rect 14439 34612 14445 34646
rect 14399 34574 14445 34612
rect 12372 34552 12378 34555
rect 9783 34492 9829 34530
rect 9783 34458 9789 34492
rect 9823 34458 9829 34492
rect 9783 34420 9829 34458
rect 9783 34386 9789 34420
rect 9823 34386 9829 34420
rect 9783 34348 9829 34386
rect 9783 34314 9789 34348
rect 9823 34314 9829 34348
rect 9783 34276 9829 34314
rect 9783 34242 9789 34276
rect 9823 34242 9829 34276
rect 9783 34230 9829 34242
rect 10034 34546 12378 34552
rect 12430 34546 12459 34555
rect 12511 34546 12540 34555
rect 12592 34546 12620 34555
rect 12672 34552 12678 34555
rect 12672 34546 14199 34552
rect 10034 34512 10046 34546
rect 10080 34512 10118 34546
rect 10152 34512 10190 34546
rect 10224 34512 10262 34546
rect 10296 34512 10334 34546
rect 10368 34512 10406 34546
rect 10440 34512 10478 34546
rect 10512 34512 10550 34546
rect 10584 34512 10622 34546
rect 10656 34512 10694 34546
rect 10728 34512 10766 34546
rect 10800 34512 10838 34546
rect 10872 34512 10910 34546
rect 10944 34512 10982 34546
rect 11016 34512 11054 34546
rect 11088 34512 11126 34546
rect 11160 34512 11198 34546
rect 11232 34512 11270 34546
rect 11304 34512 11342 34546
rect 11376 34512 11414 34546
rect 11448 34512 11486 34546
rect 11520 34512 11558 34546
rect 11592 34512 11630 34546
rect 11664 34512 11702 34546
rect 11736 34512 11774 34546
rect 11808 34512 11846 34546
rect 11880 34512 11918 34546
rect 11952 34512 11990 34546
rect 12024 34512 12062 34546
rect 12096 34512 12134 34546
rect 12168 34512 12206 34546
rect 12240 34512 12278 34546
rect 12312 34512 12350 34546
rect 12456 34512 12459 34546
rect 12528 34512 12540 34546
rect 12600 34512 12620 34546
rect 12672 34512 12710 34546
rect 12744 34512 12782 34546
rect 12816 34512 12854 34546
rect 12888 34512 12926 34546
rect 12960 34512 12998 34546
rect 13032 34512 13070 34546
rect 13104 34512 13142 34546
rect 13176 34512 13214 34546
rect 13248 34512 13286 34546
rect 13320 34512 13358 34546
rect 13392 34512 13430 34546
rect 13464 34512 13502 34546
rect 13536 34512 13574 34546
rect 13608 34512 13646 34546
rect 13680 34512 13718 34546
rect 13752 34512 13790 34546
rect 13824 34512 13862 34546
rect 13896 34512 13934 34546
rect 13968 34512 14006 34546
rect 14040 34512 14078 34546
rect 14112 34540 14199 34546
rect 14112 34512 14159 34540
rect 10034 34506 12378 34512
rect 10034 34420 10080 34506
rect 12372 34503 12378 34506
rect 12430 34503 12459 34512
rect 12511 34503 12540 34512
rect 12592 34503 12620 34512
rect 12672 34506 14159 34512
rect 14193 34506 14199 34540
rect 12672 34503 12678 34506
rect 14153 34468 14199 34506
rect 10500 34460 10506 34466
rect 10034 34386 10040 34420
rect 10074 34386 10080 34420
rect 10207 34454 10506 34460
rect 10207 34420 10219 34454
rect 10253 34420 10292 34454
rect 10326 34420 10365 34454
rect 10399 34420 10438 34454
rect 10472 34420 10506 34454
rect 10207 34414 10506 34420
rect 10558 34414 10570 34466
rect 10622 34414 10680 34466
rect 10681 34415 10682 34465
rect 10718 34415 10719 34465
rect 10720 34414 10778 34466
rect 10830 34414 10842 34466
rect 10894 34414 10952 34466
rect 10953 34415 10954 34465
rect 10990 34415 10991 34465
rect 10992 34460 11044 34466
rect 13926 34460 13978 34466
rect 13980 34465 14016 34466
rect 10992 34454 13978 34460
rect 10992 34420 11105 34454
rect 11139 34420 11178 34454
rect 11212 34420 11251 34454
rect 11285 34420 11324 34454
rect 11358 34420 11397 34454
rect 11431 34420 11470 34454
rect 11504 34420 11543 34454
rect 11577 34420 11616 34454
rect 11650 34420 11689 34454
rect 11723 34420 11762 34454
rect 11796 34420 11835 34454
rect 11869 34420 11908 34454
rect 11942 34420 11981 34454
rect 12015 34420 12054 34454
rect 12088 34420 12127 34454
rect 12161 34420 12200 34454
rect 12234 34420 12273 34454
rect 12307 34420 12346 34454
rect 12380 34420 12419 34454
rect 12453 34420 12492 34454
rect 12526 34420 12565 34454
rect 12599 34420 12638 34454
rect 12672 34420 12711 34454
rect 12745 34420 12784 34454
rect 12818 34420 12857 34454
rect 12891 34420 12930 34454
rect 12964 34420 13003 34454
rect 13037 34420 13076 34454
rect 13110 34420 13149 34454
rect 13183 34420 13222 34454
rect 13256 34420 13295 34454
rect 13329 34420 13368 34454
rect 13402 34420 13441 34454
rect 13475 34420 13514 34454
rect 13548 34420 13587 34454
rect 13621 34420 13660 34454
rect 13694 34420 13733 34454
rect 13767 34420 13806 34454
rect 13840 34420 13880 34454
rect 13914 34420 13978 34454
rect 10992 34414 13978 34420
rect 13979 34415 14017 34465
rect 14018 34460 14122 34466
rect 13980 34414 14016 34415
rect 14018 34414 14070 34460
rect 10034 34348 10080 34386
rect 10034 34314 10040 34348
rect 10074 34314 10080 34348
rect 14070 34396 14122 34408
rect 14070 34338 14122 34344
rect 14153 34434 14159 34468
rect 14193 34434 14199 34468
rect 14153 34396 14199 34434
rect 14153 34362 14159 34396
rect 14193 34362 14199 34396
rect 10034 34276 10080 34314
rect 10034 34242 10040 34276
rect 10074 34242 10080 34276
rect 10034 34230 10080 34242
rect 14153 34324 14199 34362
rect 14153 34290 14159 34324
rect 14193 34290 14199 34324
rect 14153 34252 14199 34290
rect 14153 34218 14159 34252
rect 14193 34218 14199 34252
rect 14153 34180 14199 34218
rect 14153 34146 14159 34180
rect 14193 34146 14199 34180
rect 14153 34108 14199 34146
rect 14153 34074 14159 34108
rect 14193 34074 14199 34108
rect 14153 34036 14199 34074
rect 14153 34002 14159 34036
rect 14193 34002 14199 34036
rect 14153 33964 14199 34002
rect 14153 33930 14159 33964
rect 14193 33930 14199 33964
rect 14153 33892 14199 33930
rect 14153 33858 14159 33892
rect 14193 33858 14199 33892
rect 14153 33820 14199 33858
rect 14070 33796 14122 33802
rect 14070 33732 14122 33744
rect 10500 33674 10506 33726
rect 10558 33674 10570 33726
rect 10622 33674 13978 33726
rect 13980 33725 14016 33726
rect 13979 33675 14017 33725
rect 14018 33680 14070 33726
rect 13980 33674 14016 33675
rect 14018 33674 14122 33680
rect 14153 33786 14159 33820
rect 14193 33786 14199 33820
rect 14153 33748 14199 33786
rect 14153 33714 14159 33748
rect 14193 33714 14199 33748
rect 14153 33676 14199 33714
rect 10034 33596 10080 33656
rect 10034 33579 10040 33596
rect 9836 33562 10040 33579
rect 10074 33579 10080 33596
rect 14153 33642 14159 33676
rect 14193 33642 14199 33676
rect 14153 33604 14199 33642
rect 14153 33579 14159 33604
rect 10074 33567 12378 33579
rect 10074 33562 10162 33567
rect 9836 33533 10162 33562
rect 10196 33533 11018 33567
rect 11052 33533 11874 33567
rect 11908 33533 12378 33567
rect 9836 33527 12378 33533
rect 12430 33527 12459 33579
rect 12511 33527 12540 33579
rect 12592 33527 12620 33579
rect 12672 33570 14159 33579
rect 14193 33570 14199 33604
rect 12672 33567 14199 33570
rect 12672 33533 12730 33567
rect 12764 33533 13586 33567
rect 13620 33533 14042 33567
rect 14076 33533 14199 33567
rect 12672 33532 14199 33533
rect 12672 33527 14159 33532
rect 9836 33524 14159 33527
rect 9836 33490 10040 33524
rect 10074 33503 14159 33524
rect 10074 33492 12378 33503
rect 10074 33490 10162 33492
rect 9836 33487 10162 33490
rect 9836 33453 9842 33487
rect 9876 33458 10162 33487
rect 10196 33458 11018 33492
rect 11052 33458 11874 33492
rect 11908 33458 12378 33492
rect 9876 33453 12378 33458
rect 9836 33452 12378 33453
rect 9836 33418 10040 33452
rect 10074 33451 12378 33452
rect 12430 33451 12459 33503
rect 12511 33451 12540 33503
rect 12592 33451 12620 33503
rect 12672 33498 14159 33503
rect 14193 33498 14199 33532
rect 12672 33492 14199 33498
rect 12672 33458 12730 33492
rect 12764 33458 13586 33492
rect 13620 33458 14042 33492
rect 14076 33458 14199 33492
rect 12672 33452 14199 33458
rect 12672 33451 14159 33452
rect 10074 33427 14159 33451
rect 10074 33418 12378 33427
rect 9836 33417 12378 33418
rect 9836 33414 10162 33417
rect 9836 33380 9842 33414
rect 9876 33383 10162 33414
rect 10196 33383 11018 33417
rect 11052 33383 11874 33417
rect 11908 33383 12378 33417
rect 9876 33380 12378 33383
rect 9836 33346 10040 33380
rect 10074 33375 12378 33380
rect 12430 33375 12459 33427
rect 12511 33375 12540 33427
rect 12592 33375 12620 33427
rect 12672 33418 14159 33427
rect 14193 33418 14199 33452
rect 12672 33417 14199 33418
rect 12672 33383 12730 33417
rect 12764 33383 13586 33417
rect 13620 33383 14042 33417
rect 14076 33383 14199 33417
rect 12672 33380 14199 33383
rect 12672 33375 14159 33380
rect 10074 33351 14159 33375
rect 10074 33346 12378 33351
rect 9836 33342 12378 33346
rect 9836 33341 10162 33342
rect 9836 33307 9842 33341
rect 9876 33308 10162 33341
rect 10196 33308 11018 33342
rect 11052 33308 11874 33342
rect 11908 33308 12378 33342
rect 9876 33307 10040 33308
rect 9836 33274 10040 33307
rect 10074 33299 12378 33308
rect 12430 33299 12459 33351
rect 12511 33299 12540 33351
rect 12592 33299 12620 33351
rect 12672 33346 14159 33351
rect 14193 33346 14199 33380
rect 12672 33342 14199 33346
rect 12672 33308 12730 33342
rect 12764 33308 13586 33342
rect 13620 33308 14042 33342
rect 14076 33308 14199 33342
rect 12672 33299 14159 33308
rect 10074 33275 14159 33299
rect 10074 33274 12378 33275
rect 9836 33267 12378 33274
rect 9836 33233 9842 33267
rect 9876 33236 10162 33267
rect 9876 33233 10040 33236
rect 9836 33202 10040 33233
rect 10074 33233 10162 33236
rect 10196 33233 11018 33267
rect 11052 33233 11874 33267
rect 11908 33233 12378 33267
rect 10074 33223 12378 33233
rect 12430 33223 12459 33275
rect 12511 33223 12540 33275
rect 12592 33223 12620 33275
rect 12672 33274 14159 33275
rect 14193 33274 14199 33308
rect 12672 33267 14199 33274
rect 12672 33233 12730 33267
rect 12764 33233 13586 33267
rect 13620 33233 14042 33267
rect 14076 33236 14199 33267
rect 14076 33233 14159 33236
rect 12672 33223 14159 33233
rect 10074 33202 14159 33223
rect 14193 33202 14199 33236
rect 9836 33199 14199 33202
rect 9836 33193 12378 33199
rect 9836 33159 9842 33193
rect 9876 33164 10162 33193
rect 9876 33159 10040 33164
rect 9836 33147 10040 33159
rect 10034 33130 10040 33147
rect 10074 33159 10162 33164
rect 10196 33159 11018 33193
rect 11052 33159 11874 33193
rect 11908 33159 12378 33193
rect 10074 33147 12378 33159
rect 12430 33147 12459 33199
rect 12511 33147 12540 33199
rect 12592 33147 12620 33199
rect 12672 33193 14199 33199
rect 12672 33159 12730 33193
rect 12764 33159 13586 33193
rect 13620 33159 14042 33193
rect 14076 33164 14199 33193
rect 14076 33159 14159 33164
rect 12672 33147 14159 33159
rect 10074 33130 10080 33147
rect 10034 33092 10080 33130
rect 10034 33058 10040 33092
rect 10074 33058 10080 33092
rect 10034 33020 10080 33058
rect 10034 32986 10040 33020
rect 10074 32986 10080 33020
rect 10034 32948 10080 32986
rect 10034 32914 10040 32948
rect 10074 32914 10080 32948
rect 10034 32876 10080 32914
rect 10034 32842 10040 32876
rect 10074 32842 10080 32876
rect 10034 32804 10080 32842
rect 10034 32770 10040 32804
rect 10074 32770 10080 32804
rect 10034 32732 10080 32770
rect 10034 32698 10040 32732
rect 10074 32698 10080 32732
rect 10034 32660 10080 32698
rect 10034 32626 10040 32660
rect 10074 32626 10080 32660
rect 10034 32588 10080 32626
rect 10034 32554 10040 32588
rect 10074 32554 10080 32588
rect 10034 32516 10080 32554
rect 10034 32482 10040 32516
rect 10074 32482 10080 32516
rect 10034 32444 10080 32482
rect 10034 32410 10040 32444
rect 10074 32410 10080 32444
rect 10034 32372 10080 32410
rect 10034 32338 10040 32372
rect 10074 32338 10080 32372
rect 10034 32300 10080 32338
rect 14153 33130 14159 33147
rect 14193 33130 14199 33164
rect 14153 33092 14199 33130
rect 14153 33058 14159 33092
rect 14193 33058 14199 33092
rect 14153 33020 14199 33058
rect 14153 32986 14159 33020
rect 14193 32986 14199 33020
rect 14153 32948 14199 32986
rect 14153 32914 14159 32948
rect 14193 32914 14199 32948
rect 14153 32876 14199 32914
rect 14153 32842 14159 32876
rect 14193 32842 14199 32876
rect 14153 32804 14199 32842
rect 14153 32770 14159 32804
rect 14193 32770 14199 32804
rect 14153 32732 14199 32770
rect 14153 32698 14159 32732
rect 14193 32698 14199 32732
rect 14153 32660 14199 32698
rect 14153 32626 14159 32660
rect 14193 32626 14199 32660
rect 14153 32588 14199 32626
rect 14153 32554 14159 32588
rect 14193 32554 14199 32588
rect 14153 32516 14199 32554
rect 14153 32482 14159 32516
rect 14193 32482 14199 32516
rect 14153 32444 14199 32482
rect 14153 32410 14159 32444
rect 14193 32410 14199 32444
rect 14153 32372 14199 32410
rect 14153 32338 14159 32372
rect 14193 32338 14199 32372
rect 12372 32300 12378 32303
rect 10034 32266 10040 32300
rect 10074 32294 12378 32300
rect 12430 32294 12459 32303
rect 12511 32294 12540 32303
rect 12592 32294 12620 32303
rect 12672 32300 12678 32303
rect 14153 32300 14199 32338
rect 12672 32294 14159 32300
rect 10074 32266 10112 32294
rect 10034 32260 10112 32266
rect 10146 32260 10185 32294
rect 10219 32260 10258 32294
rect 10292 32260 10331 32294
rect 10365 32260 10404 32294
rect 10438 32260 10477 32294
rect 10511 32260 10550 32294
rect 10584 32260 10623 32294
rect 10657 32260 10696 32294
rect 10730 32260 10769 32294
rect 10803 32260 10842 32294
rect 10876 32260 10915 32294
rect 10949 32260 10988 32294
rect 11022 32260 11061 32294
rect 11095 32260 11134 32294
rect 11168 32260 11207 32294
rect 11241 32260 11279 32294
rect 11313 32260 11351 32294
rect 11385 32260 11423 32294
rect 11457 32260 11495 32294
rect 11529 32260 11567 32294
rect 11601 32260 11639 32294
rect 11673 32260 11711 32294
rect 11745 32260 11783 32294
rect 11817 32260 11855 32294
rect 11889 32260 11927 32294
rect 11961 32260 11999 32294
rect 12033 32260 12071 32294
rect 12105 32260 12143 32294
rect 12177 32260 12215 32294
rect 12249 32260 12287 32294
rect 12321 32260 12359 32294
rect 12430 32260 12431 32294
rect 12537 32260 12540 32294
rect 12609 32260 12620 32294
rect 12681 32260 12719 32294
rect 12753 32260 12791 32294
rect 12825 32260 12863 32294
rect 12897 32260 12935 32294
rect 12969 32260 13007 32294
rect 13041 32260 13079 32294
rect 13113 32260 13151 32294
rect 13185 32260 13223 32294
rect 13257 32260 13295 32294
rect 13329 32260 13367 32294
rect 13401 32260 13439 32294
rect 13473 32260 13511 32294
rect 13545 32260 13583 32294
rect 13617 32260 13655 32294
rect 13689 32260 13727 32294
rect 13761 32260 13799 32294
rect 13833 32260 13871 32294
rect 13905 32260 13943 32294
rect 13977 32260 14015 32294
rect 14049 32260 14087 32294
rect 14121 32266 14159 32294
rect 14193 32266 14199 32300
rect 14121 32260 14199 32266
rect 10034 32254 12378 32260
rect 12372 32251 12378 32254
rect 12430 32251 12459 32260
rect 12511 32251 12540 32260
rect 12592 32251 12620 32260
rect 12672 32254 14199 32260
rect 12672 32251 12678 32254
rect 14153 32228 14199 32254
rect 10500 32208 10506 32214
rect 9522 32202 10506 32208
rect 10558 32202 10570 32214
rect 10622 32208 10628 32214
rect 10622 32202 10689 32208
rect 9522 32168 9534 32202
rect 9568 32168 9611 32202
rect 9645 32168 9688 32202
rect 9722 32168 10219 32202
rect 10253 32168 10304 32202
rect 10338 32168 10389 32202
rect 10423 32168 10474 32202
rect 10558 32168 10559 32202
rect 10622 32168 10643 32202
rect 10677 32168 10689 32202
rect 9522 32162 10506 32168
rect 10558 32162 10570 32168
rect 10622 32162 10689 32168
rect 10772 32162 10778 32214
rect 10830 32162 10842 32214
rect 10894 32162 10952 32214
rect 10953 32163 10954 32213
rect 10990 32163 10991 32213
rect 10992 32208 11044 32214
rect 13926 32208 13978 32214
rect 13980 32213 14016 32214
rect 10992 32202 13978 32208
rect 10992 32168 11105 32202
rect 11139 32168 11178 32202
rect 11212 32168 11251 32202
rect 11285 32168 11324 32202
rect 11358 32168 11397 32202
rect 11431 32168 11470 32202
rect 11504 32168 11543 32202
rect 11577 32168 11616 32202
rect 11650 32168 11689 32202
rect 11723 32168 11762 32202
rect 11796 32168 11835 32202
rect 11869 32168 11908 32202
rect 11942 32168 11981 32202
rect 12015 32168 12054 32202
rect 12088 32168 12127 32202
rect 12161 32168 12200 32202
rect 12234 32168 12273 32202
rect 12307 32168 12346 32202
rect 12380 32168 12419 32202
rect 12453 32168 12492 32202
rect 12526 32168 12565 32202
rect 12599 32168 12638 32202
rect 12672 32168 12711 32202
rect 12745 32168 12784 32202
rect 12818 32168 12857 32202
rect 12891 32168 12930 32202
rect 12964 32168 13003 32202
rect 13037 32168 13076 32202
rect 13110 32168 13149 32202
rect 13183 32168 13222 32202
rect 13256 32168 13295 32202
rect 13329 32168 13368 32202
rect 13402 32168 13441 32202
rect 13475 32168 13514 32202
rect 13548 32168 13587 32202
rect 13621 32168 13660 32202
rect 13694 32168 13733 32202
rect 13767 32168 13806 32202
rect 13840 32168 13880 32202
rect 13914 32168 13978 32202
rect 10992 32162 13978 32168
rect 13979 32163 14017 32213
rect 14018 32208 14122 32214
rect 13980 32162 14016 32163
rect 14018 32162 14070 32208
rect 14070 32144 14122 32156
rect 14070 32086 14122 32092
rect 14153 32194 14159 32228
rect 14193 32194 14199 32228
rect 14153 32156 14199 32194
rect 14153 32122 14159 32156
rect 14193 32122 14199 32156
rect 14153 32084 14199 32122
rect 14153 32050 14159 32084
rect 14193 32050 14199 32084
rect 14153 32012 14199 32050
rect 14153 31978 14159 32012
rect 14193 31978 14199 32012
rect 14153 31940 14199 31978
rect 14153 31906 14159 31940
rect 14193 31906 14199 31940
rect 14153 31868 14199 31906
rect 14153 31834 14159 31868
rect 14193 31834 14199 31868
rect 14153 31796 14199 31834
rect 14153 31762 14159 31796
rect 14193 31762 14199 31796
rect 14153 31724 14199 31762
rect 14153 31690 14159 31724
rect 14193 31690 14199 31724
rect 14153 31652 14199 31690
rect 10034 31578 10080 31621
rect 10034 31544 10040 31578
rect 10074 31544 10080 31578
rect 10034 31506 10080 31544
rect 10034 31472 10040 31506
rect 10074 31472 10080 31506
rect 10034 31434 10080 31472
rect 10034 31400 10040 31434
rect 10074 31400 10080 31434
rect 10034 31362 10080 31400
rect 10034 31328 10040 31362
rect 10074 31328 10080 31362
rect 10034 31294 10080 31328
rect 14153 31618 14159 31652
rect 14193 31618 14199 31652
rect 14153 31580 14199 31618
rect 14153 31546 14159 31580
rect 14193 31546 14199 31580
rect 14153 31508 14199 31546
rect 14153 31474 14159 31508
rect 14193 31474 14199 31508
rect 14153 31436 14199 31474
rect 14153 31402 14159 31436
rect 14193 31402 14199 31436
rect 14153 31364 14199 31402
rect 14153 31330 14159 31364
rect 14193 31330 14199 31364
rect 14153 31294 14199 31330
rect 10034 31290 11788 31294
rect 10034 31256 10040 31290
rect 10074 31282 11788 31290
rect 10074 31256 10162 31282
rect 10034 31248 10162 31256
rect 10196 31248 11018 31282
rect 11052 31248 11788 31282
rect 10034 31242 11788 31248
rect 11840 31282 11892 31294
rect 11840 31248 11874 31282
rect 11840 31242 11892 31248
rect 11944 31242 12378 31294
rect 12430 31242 12459 31294
rect 12511 31242 12540 31294
rect 12592 31242 12620 31294
rect 12672 31292 14199 31294
rect 12672 31282 14159 31292
rect 12672 31248 12730 31282
rect 12764 31248 13586 31282
rect 13620 31248 14042 31282
rect 14076 31258 14159 31282
rect 14193 31258 14199 31292
rect 14076 31248 14199 31258
rect 12672 31242 14199 31248
rect 10034 31220 14199 31242
rect 10034 31218 14159 31220
rect 10034 31184 10040 31218
rect 10074 31207 11788 31218
rect 10074 31184 10162 31207
rect 9783 31146 9829 31184
rect 9783 31112 9789 31146
rect 9823 31112 9829 31146
rect 9783 31074 9829 31112
rect 9783 31040 9789 31074
rect 9823 31040 9829 31074
rect 9783 31002 9829 31040
rect 9783 30968 9789 31002
rect 9823 30968 9829 31002
rect 9783 30930 9829 30968
rect 9783 30896 9789 30930
rect 9823 30896 9829 30930
rect 9783 30858 9829 30896
rect 9783 30824 9789 30858
rect 9823 30824 9829 30858
rect 9783 30812 9829 30824
rect 10034 31173 10162 31184
rect 10196 31173 11018 31207
rect 11052 31173 11788 31207
rect 10034 31166 11788 31173
rect 11840 31207 11892 31218
rect 11840 31173 11874 31207
rect 11840 31166 11892 31173
rect 11944 31166 12378 31218
rect 12430 31166 12459 31218
rect 12511 31166 12540 31218
rect 12592 31166 12620 31218
rect 12672 31207 14159 31218
rect 12672 31173 12730 31207
rect 12764 31173 13586 31207
rect 13620 31173 14042 31207
rect 14076 31186 14159 31207
rect 14193 31186 14199 31220
rect 14076 31173 14199 31186
rect 12672 31166 14199 31173
rect 10034 31148 14199 31166
rect 10034 31146 14159 31148
rect 10034 31112 10040 31146
rect 10074 31142 14159 31146
rect 10074 31132 11788 31142
rect 10074 31112 10162 31132
rect 10034 31098 10162 31112
rect 10196 31098 11018 31132
rect 11052 31098 11788 31132
rect 10034 31090 11788 31098
rect 11840 31132 11892 31142
rect 11840 31098 11874 31132
rect 11840 31090 11892 31098
rect 11944 31090 12378 31142
rect 12430 31090 12459 31142
rect 12511 31090 12540 31142
rect 12592 31090 12620 31142
rect 12672 31132 14159 31142
rect 12672 31098 12730 31132
rect 12764 31098 13586 31132
rect 13620 31098 14042 31132
rect 14076 31114 14159 31132
rect 14193 31114 14199 31148
rect 14076 31098 14199 31114
rect 12672 31090 14199 31098
rect 10034 31076 14199 31090
rect 10034 31074 14159 31076
rect 10034 31040 10040 31074
rect 10074 31066 14159 31074
rect 10074 31057 11788 31066
rect 10074 31040 10162 31057
rect 10034 31023 10162 31040
rect 10196 31023 11018 31057
rect 11052 31023 11788 31057
rect 10034 31014 11788 31023
rect 11840 31057 11892 31066
rect 11840 31023 11874 31057
rect 11840 31014 11892 31023
rect 11944 31014 12378 31066
rect 12430 31014 12459 31066
rect 12511 31014 12540 31066
rect 12592 31014 12620 31066
rect 12672 31057 14159 31066
rect 12672 31023 12730 31057
rect 12764 31023 13586 31057
rect 13620 31023 14042 31057
rect 14076 31042 14159 31057
rect 14193 31042 14199 31076
rect 14076 31023 14199 31042
rect 12672 31014 14199 31023
rect 10034 31004 14199 31014
rect 10034 31002 14159 31004
rect 10034 30968 10040 31002
rect 10074 30990 14159 31002
rect 10074 30982 11788 30990
rect 10074 30968 10162 30982
rect 10034 30948 10162 30968
rect 10196 30948 11018 30982
rect 11052 30948 11788 30982
rect 10034 30938 11788 30948
rect 11840 30982 11892 30990
rect 11840 30948 11874 30982
rect 11840 30938 11892 30948
rect 11944 30938 12378 30990
rect 12430 30938 12459 30990
rect 12511 30938 12540 30990
rect 12592 30938 12620 30990
rect 12672 30982 14159 30990
rect 12672 30948 12730 30982
rect 12764 30948 13586 30982
rect 13620 30948 14042 30982
rect 14076 30970 14159 30982
rect 14193 30970 14199 31004
rect 14076 30948 14199 30970
rect 12672 30938 14199 30948
rect 10034 30932 14199 30938
rect 10034 30930 14159 30932
rect 10034 30896 10040 30930
rect 10074 30914 14159 30930
rect 10074 30908 11788 30914
rect 10074 30896 10162 30908
rect 10034 30874 10162 30896
rect 10196 30874 11018 30908
rect 11052 30874 11788 30908
rect 10034 30862 11788 30874
rect 11840 30908 11892 30914
rect 11840 30874 11874 30908
rect 11840 30862 11892 30874
rect 11944 30862 12378 30914
rect 12430 30862 12459 30914
rect 12511 30862 12540 30914
rect 12592 30862 12620 30914
rect 12672 30908 14159 30914
rect 12672 30874 12730 30908
rect 12764 30874 13586 30908
rect 13620 30874 14042 30908
rect 14076 30898 14159 30908
rect 14193 30898 14199 30932
rect 14076 30874 14199 30898
rect 12672 30862 14199 30874
rect 10034 30858 10080 30862
rect 10034 30824 10040 30858
rect 10074 30824 10080 30858
rect 10034 30812 10080 30824
rect 14153 30860 14199 30862
rect 14153 30826 14159 30860
rect 14193 30826 14199 30860
rect 14153 30788 14199 30826
rect 14153 30754 14159 30788
rect 14193 30754 14199 30788
rect 14153 30716 14199 30754
rect 14153 30682 14159 30716
rect 14193 30682 14199 30716
rect 14153 30644 14199 30682
rect 14153 30610 14159 30644
rect 14193 30610 14199 30644
rect 14153 30572 14199 30610
rect 14153 30538 14159 30572
rect 14193 30538 14199 30572
rect 14153 30500 14199 30538
rect 14153 30466 14159 30500
rect 14193 30466 14199 30500
rect 14153 30428 14199 30466
rect 14153 30394 14159 30428
rect 14193 30394 14199 30428
rect 14153 30356 14199 30394
rect 14153 30322 14159 30356
rect 14193 30322 14199 30356
rect 14153 30284 14199 30322
rect 14153 30250 14159 30284
rect 14193 30250 14199 30284
rect 14153 30212 14199 30250
rect 14153 30178 14159 30212
rect 14193 30178 14199 30212
rect 9783 30096 9829 30148
rect 9783 30062 9789 30096
rect 9823 30062 9829 30096
rect 9783 30024 9829 30062
rect 9783 29990 9789 30024
rect 9823 29990 9829 30024
rect 9783 29952 9829 29990
rect 9783 29918 9789 29952
rect 9823 29918 9829 29952
rect 9783 29880 9829 29918
rect 9783 29846 9789 29880
rect 9823 29846 9829 29880
rect 9783 29808 9829 29846
rect 9783 29774 9789 29808
rect 9823 29774 9829 29808
rect 9783 29736 9829 29774
rect 9783 29702 9789 29736
rect 9823 29702 9829 29736
rect 9783 29690 9829 29702
rect 10034 30096 10080 30148
rect 10034 30062 10040 30096
rect 10074 30062 10080 30096
rect 10034 30049 10080 30062
rect 14153 30140 14199 30178
rect 14153 30106 14159 30140
rect 14193 30106 14199 30140
rect 14153 30068 14199 30106
rect 11782 30049 11788 30052
rect 10034 30043 11788 30049
rect 11840 30043 11892 30052
rect 11944 30049 11950 30052
rect 14153 30049 14159 30068
rect 11944 30043 14159 30049
rect 10034 30024 10112 30043
rect 10034 29990 10040 30024
rect 10074 30009 10112 30024
rect 10146 30009 10185 30043
rect 10219 30009 10258 30043
rect 10292 30009 10331 30043
rect 10365 30009 10404 30043
rect 10438 30009 10477 30043
rect 10511 30009 10550 30043
rect 10584 30009 10623 30043
rect 10657 30009 10696 30043
rect 10730 30009 10769 30043
rect 10803 30009 10842 30043
rect 10876 30009 10915 30043
rect 10949 30009 10988 30043
rect 11022 30009 11061 30043
rect 11095 30009 11134 30043
rect 11168 30009 11207 30043
rect 11241 30009 11279 30043
rect 11313 30009 11351 30043
rect 11385 30009 11423 30043
rect 11457 30009 11495 30043
rect 11529 30009 11567 30043
rect 11601 30009 11639 30043
rect 11673 30009 11711 30043
rect 11745 30009 11783 30043
rect 11840 30009 11855 30043
rect 11889 30009 11892 30043
rect 11961 30009 11999 30043
rect 12033 30009 12071 30043
rect 12105 30009 12143 30043
rect 12177 30009 12215 30043
rect 12249 30009 12287 30043
rect 12321 30009 12359 30043
rect 12393 30009 12431 30043
rect 12465 30009 12503 30043
rect 12537 30009 12575 30043
rect 12609 30009 12647 30043
rect 12681 30009 12719 30043
rect 12753 30009 12791 30043
rect 12825 30009 12863 30043
rect 12897 30009 12935 30043
rect 12969 30009 13007 30043
rect 13041 30009 13079 30043
rect 13113 30009 13151 30043
rect 13185 30009 13223 30043
rect 13257 30009 13295 30043
rect 13329 30009 13367 30043
rect 13401 30009 13439 30043
rect 13473 30009 13511 30043
rect 13545 30009 13583 30043
rect 13617 30009 13655 30043
rect 13689 30009 13727 30043
rect 13761 30009 13799 30043
rect 13833 30009 13871 30043
rect 13905 30009 13943 30043
rect 13977 30009 14015 30043
rect 14049 30009 14087 30043
rect 14121 30034 14159 30043
rect 14193 30034 14199 30068
rect 14121 30009 14199 30034
rect 10074 30003 11788 30009
rect 10074 29990 10080 30003
rect 11782 30000 11788 30003
rect 11840 30000 11892 30009
rect 11944 30003 14199 30009
rect 11944 30000 11950 30003
rect 10034 29952 10080 29990
rect 14153 29996 14199 30003
rect 10500 29959 10506 29965
rect 10034 29918 10040 29952
rect 10074 29918 10080 29952
rect 10034 29880 10080 29918
rect 10207 29953 10506 29959
rect 10558 29953 10570 29965
rect 10622 29959 10628 29965
rect 10622 29953 10689 29959
rect 10207 29919 10219 29953
rect 10253 29919 10304 29953
rect 10338 29919 10389 29953
rect 10423 29919 10474 29953
rect 10558 29919 10559 29953
rect 10622 29919 10643 29953
rect 10677 29919 10689 29953
rect 10207 29913 10506 29919
rect 10558 29913 10570 29919
rect 10622 29913 10689 29919
rect 10772 29913 10778 29965
rect 10830 29913 10842 29965
rect 10894 29913 10952 29965
rect 10953 29914 10954 29964
rect 10990 29914 10991 29964
rect 10992 29959 11044 29965
rect 13926 29959 13978 29965
rect 13980 29964 14016 29965
rect 10992 29953 13978 29959
rect 10992 29919 11105 29953
rect 11139 29919 11178 29953
rect 11212 29919 11251 29953
rect 11285 29919 11324 29953
rect 11358 29919 11397 29953
rect 11431 29919 11470 29953
rect 11504 29919 11543 29953
rect 11577 29919 11616 29953
rect 11650 29919 11689 29953
rect 11723 29919 11762 29953
rect 11796 29919 11835 29953
rect 11869 29919 11908 29953
rect 11942 29919 11981 29953
rect 12015 29919 12054 29953
rect 12088 29919 12127 29953
rect 12161 29919 12200 29953
rect 12234 29919 12273 29953
rect 12307 29919 12346 29953
rect 12380 29919 12419 29953
rect 12453 29919 12492 29953
rect 12526 29919 12565 29953
rect 12599 29919 12638 29953
rect 12672 29919 12711 29953
rect 12745 29919 12784 29953
rect 12818 29919 12857 29953
rect 12891 29919 12930 29953
rect 12964 29919 13003 29953
rect 13037 29919 13076 29953
rect 13110 29919 13149 29953
rect 13183 29919 13222 29953
rect 13256 29919 13295 29953
rect 13329 29919 13368 29953
rect 13402 29919 13441 29953
rect 13475 29919 13514 29953
rect 13548 29919 13587 29953
rect 13621 29919 13660 29953
rect 13694 29919 13733 29953
rect 13767 29919 13806 29953
rect 13840 29919 13880 29953
rect 13914 29919 13978 29953
rect 10992 29913 13978 29919
rect 13979 29914 14017 29964
rect 14018 29959 14122 29965
rect 13980 29913 14016 29914
rect 14018 29913 14070 29959
rect 10034 29846 10040 29880
rect 10074 29846 10080 29880
rect 10034 29808 10080 29846
rect 14070 29895 14122 29907
rect 14070 29837 14122 29843
rect 14153 29962 14159 29996
rect 14193 29962 14199 29996
rect 14153 29924 14199 29962
rect 14153 29890 14159 29924
rect 14193 29890 14199 29924
rect 14153 29852 14199 29890
rect 10034 29774 10040 29808
rect 10074 29774 10080 29808
rect 10034 29736 10080 29774
rect 10034 29702 10040 29736
rect 10074 29702 10080 29736
rect 10034 29690 10080 29702
rect 14153 29818 14159 29852
rect 14193 29818 14199 29852
rect 14153 29780 14199 29818
rect 14153 29746 14159 29780
rect 14193 29746 14199 29780
rect 14153 29708 14199 29746
rect 14153 29674 14159 29708
rect 14193 29674 14199 29708
rect 14153 29636 14199 29674
rect 14153 29602 14159 29636
rect 14193 29602 14199 29636
rect 14153 29564 14199 29602
rect 14153 29530 14159 29564
rect 14193 29530 14199 29564
rect 14153 29492 14199 29530
rect 14153 29458 14159 29492
rect 14193 29458 14199 29492
rect 14070 29447 14122 29453
rect 14070 29386 14122 29395
tri 8749 29356 8779 29386 se
rect 8779 29383 14122 29386
rect 8779 29356 14070 29383
tri 8741 29348 8749 29356 se
rect 8749 29348 14070 29356
tri 8727 29334 8741 29348 se
rect 8741 29334 14070 29348
tri 8708 29315 8727 29334 se
rect 8727 29325 8792 29334
tri 8792 29325 8801 29334 nw
rect 14070 29325 14122 29331
rect 14153 29420 14199 29458
rect 14153 29386 14159 29420
rect 14193 29386 14199 29420
rect 14153 29348 14199 29386
rect 8727 29315 8782 29325
tri 8782 29315 8792 29325 nw
tri 8707 29314 8708 29315 se
rect 8708 29314 8781 29315
tri 8781 29314 8782 29315 nw
rect 14153 29314 14159 29348
rect 14193 29314 14199 29348
tri 8677 29284 8707 29314 se
rect 8707 29284 8751 29314
tri 8751 29284 8781 29314 nw
tri 8669 29276 8677 29284 se
rect 8677 29276 8743 29284
tri 8743 29276 8751 29284 nw
rect 14153 29276 14199 29314
tri 8635 29242 8669 29276 se
rect 8669 29246 8713 29276
tri 8713 29246 8743 29276 nw
rect 8669 29242 8709 29246
tri 8709 29242 8713 29246 nw
tri 8634 29241 8635 29242 se
rect 8635 29241 8708 29242
tri 8708 29241 8709 29242 nw
tri 8605 29212 8634 29241 se
rect 8634 29212 8679 29241
tri 8679 29212 8708 29241 nw
rect 9721 29240 10900 29246
tri 8597 29204 8605 29212 se
rect 8605 29204 8671 29212
tri 8671 29204 8679 29212 nw
tri 8563 29170 8597 29204 se
rect 8597 29170 8637 29204
tri 8637 29170 8671 29204 nw
rect 9773 29188 9811 29240
rect 9863 29188 10772 29240
rect 10824 29188 10848 29240
tri 8560 29167 8563 29170 se
rect 8563 29167 8634 29170
tri 8634 29167 8637 29170 nw
tri 8533 29140 8560 29167 se
rect 8560 29140 8607 29167
tri 8607 29140 8634 29167 nw
rect 9721 29162 10900 29188
tri 8525 29132 8533 29140 se
rect 8533 29132 8599 29140
tri 8599 29132 8607 29140 nw
tri 8491 29098 8525 29132 se
rect 8525 29104 8571 29132
tri 8571 29104 8599 29132 nw
rect 9773 29110 9811 29162
rect 9863 29110 10772 29162
rect 10824 29110 10848 29162
rect 9721 29104 10900 29110
rect 14153 29242 14159 29276
rect 14193 29242 14199 29276
rect 14153 29204 14199 29242
rect 14153 29170 14159 29204
rect 14193 29170 14199 29204
rect 14153 29132 14199 29170
rect 8525 29098 8565 29104
tri 8565 29098 8571 29104 nw
rect 14153 29098 14159 29132
rect 14193 29098 14199 29132
tri 8486 29093 8491 29098 se
rect 8491 29093 8560 29098
tri 8560 29093 8565 29098 nw
tri 8464 29071 8486 29093 se
rect 8486 29071 8535 29093
rect 4295 29019 4301 29071
rect 4353 29019 4365 29071
rect 4417 29068 8535 29071
tri 8535 29068 8560 29093 nw
rect 4417 29060 8527 29068
tri 8527 29060 8535 29068 nw
rect 14153 29060 14199 29098
rect 4417 29026 8493 29060
tri 8493 29026 8527 29060 nw
rect 14153 29026 14159 29060
rect 14193 29026 14199 29060
rect 4417 29019 8486 29026
tri 8486 29019 8493 29026 nw
rect 10034 28990 10080 28991
rect 14153 28990 14199 29026
rect 10008 28978 11788 28990
rect 10008 28969 10162 28978
rect 5622 28959 10162 28969
rect 5622 28907 5624 28959
rect 5676 28907 5730 28959
rect 5782 28907 5836 28959
rect 5888 28944 10162 28959
rect 10196 28944 11018 28978
rect 11052 28944 11788 28978
rect 5888 28938 11788 28944
rect 11840 28978 11892 28990
rect 11944 28988 14199 28990
rect 11944 28978 14159 28988
rect 11840 28944 11874 28978
rect 11944 28944 12730 28978
rect 12764 28944 13586 28978
rect 13620 28944 14042 28978
rect 14076 28954 14159 28978
rect 14193 28954 14199 28988
rect 14076 28944 14199 28954
rect 11840 28938 11892 28944
rect 11944 28938 14199 28944
rect 5888 28932 14199 28938
rect 5888 28907 10040 28932
rect 5622 28898 10040 28907
rect 10074 28916 14199 28932
rect 10074 28914 14159 28916
rect 10074 28903 11788 28914
rect 10074 28898 10162 28903
rect 5622 28874 10162 28898
rect 5622 28822 5624 28874
rect 5676 28822 5730 28874
rect 5782 28822 5836 28874
rect 5888 28869 10162 28874
rect 10196 28869 11018 28903
rect 11052 28869 11788 28903
rect 5888 28862 11788 28869
rect 11840 28903 11892 28914
rect 11944 28903 14159 28914
rect 11840 28869 11874 28903
rect 11944 28869 12730 28903
rect 12764 28869 13586 28903
rect 13620 28869 14042 28903
rect 14076 28882 14159 28903
rect 14193 28882 14199 28916
rect 14076 28869 14199 28882
rect 11840 28862 11892 28869
rect 11944 28862 14199 28869
rect 5888 28860 14199 28862
rect 5888 28826 10040 28860
rect 10074 28844 14199 28860
rect 10074 28838 14159 28844
rect 10074 28828 11788 28838
rect 10074 28826 10162 28828
rect 5888 28822 10162 28826
rect 5622 28794 10162 28822
rect 10196 28794 11018 28828
rect 11052 28794 11788 28828
rect 5622 28788 11788 28794
rect 5622 28736 5624 28788
rect 5676 28736 5730 28788
rect 5782 28736 5836 28788
rect 5888 28754 10040 28788
rect 10074 28786 11788 28788
rect 11840 28828 11892 28838
rect 11944 28828 14159 28838
rect 11840 28794 11874 28828
rect 11944 28794 12730 28828
rect 12764 28794 13586 28828
rect 13620 28794 14042 28828
rect 14076 28810 14159 28828
rect 14193 28810 14199 28844
rect 14076 28794 14199 28810
rect 11840 28786 11892 28794
rect 11944 28786 14199 28794
rect 10074 28772 14199 28786
rect 10074 28762 14159 28772
rect 10074 28754 11788 28762
rect 5888 28753 11788 28754
rect 5888 28736 10162 28753
rect 5622 28719 10162 28736
rect 10196 28719 11018 28753
rect 11052 28719 11788 28753
rect 5622 28716 11788 28719
rect 5622 28702 10040 28716
rect 5622 28650 5624 28702
rect 5676 28650 5730 28702
rect 5782 28650 5836 28702
rect 5888 28682 10040 28702
rect 10074 28710 11788 28716
rect 11840 28753 11892 28762
rect 11944 28753 14159 28762
rect 11840 28719 11874 28753
rect 11944 28719 12730 28753
rect 12764 28719 13586 28753
rect 13620 28719 14042 28753
rect 14076 28738 14159 28753
rect 14193 28738 14199 28772
rect 14076 28719 14199 28738
rect 11840 28710 11892 28719
rect 11944 28710 14199 28719
rect 10074 28700 14199 28710
rect 10074 28686 14159 28700
rect 10074 28682 11788 28686
rect 5888 28678 11788 28682
rect 5888 28650 10162 28678
rect 5622 28644 10162 28650
rect 10196 28644 11018 28678
rect 11052 28644 11788 28678
rect 5622 28616 10040 28644
rect 5622 28564 5624 28616
rect 5676 28564 5730 28616
rect 5782 28564 5836 28616
rect 5888 28610 10040 28616
rect 10074 28634 11788 28644
rect 11840 28678 11892 28686
rect 11944 28678 14159 28686
rect 11840 28644 11874 28678
rect 11944 28644 12730 28678
rect 12764 28644 13586 28678
rect 13620 28644 14042 28678
rect 14076 28666 14159 28678
rect 14193 28666 14199 28700
rect 14076 28644 14199 28666
rect 11840 28634 11892 28644
rect 11944 28634 14199 28644
rect 10074 28628 14199 28634
rect 10074 28610 14159 28628
rect 5888 28604 11788 28610
rect 5888 28572 10162 28604
rect 5888 28564 10040 28572
rect 5622 28558 10040 28564
rect 10034 28538 10040 28558
rect 10074 28570 10162 28572
rect 10196 28570 11018 28604
rect 11052 28570 11788 28604
rect 10074 28558 11788 28570
rect 11840 28604 11892 28610
rect 11944 28604 14159 28610
rect 11840 28570 11874 28604
rect 11944 28570 12730 28604
rect 12764 28570 13586 28604
rect 13620 28570 14042 28604
rect 14076 28594 14159 28604
rect 14193 28594 14199 28628
rect 14076 28570 14199 28594
rect 11840 28558 11892 28570
rect 11944 28558 14199 28570
rect 10074 28538 10080 28558
tri 11781 28556 11783 28558 ne
rect 11783 28556 12368 28558
tri 12368 28556 12370 28558 nw
rect 14153 28556 14199 28558
rect 10034 28500 10080 28538
tri 11783 28522 11817 28556 ne
rect 11817 28522 12334 28556
tri 12334 28522 12368 28556 nw
rect 14153 28522 14159 28556
rect 14193 28522 14199 28556
rect 10034 28466 10040 28500
rect 10074 28466 10080 28500
tri 11817 28492 11847 28522 ne
rect 11847 28492 12304 28522
tri 12304 28492 12334 28522 nw
tri 11847 28484 11855 28492 ne
rect 11855 28484 12296 28492
tri 12296 28484 12304 28492 nw
rect 14153 28484 14199 28522
rect 10034 28428 10080 28466
tri 11855 28450 11889 28484 ne
rect 11889 28450 12262 28484
tri 12262 28450 12296 28484 nw
rect 14153 28450 14159 28484
rect 14193 28450 14199 28484
rect 10034 28394 10040 28428
rect 10074 28394 10080 28428
tri 11889 28420 11919 28450 ne
rect 11919 28420 12232 28450
tri 12232 28420 12262 28450 nw
tri 11919 28412 11927 28420 ne
rect 11927 28412 12224 28420
tri 12224 28412 12232 28420 nw
rect 14153 28412 14199 28450
rect 10034 28356 10080 28394
tri 11927 28391 11948 28412 ne
rect 10034 28322 10040 28356
rect 10074 28322 10080 28356
rect 10034 28284 10080 28322
rect 10034 28250 10040 28284
rect 10074 28250 10080 28284
rect 10034 28212 10080 28250
rect 10034 28178 10040 28212
rect 10074 28178 10080 28212
rect 10034 28140 10080 28178
rect 10034 28106 10040 28140
rect 10074 28106 10080 28140
rect 10034 28068 10080 28106
rect 10034 28034 10040 28068
rect 10074 28034 10080 28068
rect 10034 28022 10080 28034
rect 11948 27795 12203 28412
tri 12203 28391 12224 28412 nw
rect 14153 28378 14159 28412
rect 14193 28378 14199 28412
rect 14153 28340 14199 28378
rect 14153 28306 14159 28340
rect 14193 28306 14199 28340
rect 14153 28268 14199 28306
rect 14153 28234 14159 28268
rect 14193 28234 14199 28268
rect 14153 28196 14199 28234
rect 14153 28162 14159 28196
rect 14193 28162 14199 28196
rect 14153 28124 14199 28162
rect 14153 28090 14159 28124
rect 14193 28090 14199 28124
rect 14153 28052 14199 28090
rect 14153 28018 14159 28052
rect 14193 28018 14199 28052
rect 14153 27980 14199 28018
rect 14153 27946 14159 27980
rect 14193 27946 14199 27980
rect 14153 27908 14199 27946
rect 14153 27874 14159 27908
rect 14193 27874 14199 27908
rect 14153 27795 14199 27874
rect 10034 27789 14199 27795
rect 10034 27755 10049 27789
rect 10083 27755 10121 27789
rect 10155 27755 10193 27789
rect 10227 27755 10265 27789
rect 10299 27755 10337 27789
rect 10371 27755 10409 27789
rect 10443 27755 10481 27789
rect 10515 27755 10553 27789
rect 10587 27755 10625 27789
rect 10659 27755 10697 27789
rect 10731 27755 10769 27789
rect 10803 27755 10841 27789
rect 10875 27755 10913 27789
rect 10947 27755 10985 27789
rect 11019 27755 11057 27789
rect 11091 27755 11129 27789
rect 11163 27755 11201 27789
rect 11235 27755 11273 27789
rect 11307 27755 11345 27789
rect 11379 27755 11417 27789
rect 11451 27755 11489 27789
rect 11523 27755 11561 27789
rect 11595 27755 11633 27789
rect 11667 27755 11705 27789
rect 11739 27755 11777 27789
rect 11811 27755 11849 27789
rect 11883 27755 11921 27789
rect 11955 27755 11993 27789
rect 12027 27755 12065 27789
rect 12099 27755 12137 27789
rect 12171 27755 12209 27789
rect 12243 27755 12281 27789
rect 12315 27755 12353 27789
rect 12387 27755 12425 27789
rect 12459 27755 12497 27789
rect 12531 27755 12569 27789
rect 12603 27755 12641 27789
rect 12675 27755 12713 27789
rect 12747 27755 12785 27789
rect 12819 27755 12857 27789
rect 12891 27755 12929 27789
rect 12963 27755 13001 27789
rect 13035 27755 13073 27789
rect 13107 27755 13145 27789
rect 13179 27755 13217 27789
rect 13251 27755 13289 27789
rect 13323 27755 13361 27789
rect 13395 27755 13433 27789
rect 13467 27755 13505 27789
rect 13539 27755 13577 27789
rect 13611 27755 13649 27789
rect 13683 27755 13721 27789
rect 13755 27755 13793 27789
rect 13827 27755 13865 27789
rect 13899 27755 13937 27789
rect 13971 27755 14009 27789
rect 14043 27755 14081 27789
rect 14115 27755 14153 27789
rect 14187 27755 14199 27789
rect 10034 27749 14199 27755
rect 14399 34540 14405 34574
rect 14439 34540 14445 34574
rect 14399 34502 14445 34540
rect 14399 34468 14405 34502
rect 14439 34468 14445 34502
rect 14399 34430 14445 34468
rect 14399 34396 14405 34430
rect 14439 34396 14445 34430
rect 14399 34358 14445 34396
rect 14399 34324 14405 34358
rect 14439 34324 14445 34358
rect 14399 34286 14445 34324
rect 14399 34252 14405 34286
rect 14439 34252 14445 34286
rect 14399 34214 14445 34252
rect 14399 34180 14405 34214
rect 14439 34180 14445 34214
rect 14399 34142 14445 34180
rect 14399 34108 14405 34142
rect 14439 34108 14445 34142
rect 14399 34070 14445 34108
rect 14399 34036 14405 34070
rect 14439 34036 14445 34070
rect 14399 33998 14445 34036
rect 14399 33964 14405 33998
rect 14439 33964 14445 33998
rect 14399 33926 14445 33964
rect 14399 33892 14405 33926
rect 14439 33892 14445 33926
rect 14399 33854 14445 33892
rect 14399 33820 14405 33854
rect 14439 33820 14445 33854
rect 14399 33782 14445 33820
rect 14399 33748 14405 33782
rect 14439 33748 14445 33782
rect 14399 33710 14445 33748
rect 14399 33676 14405 33710
rect 14439 33676 14445 33710
rect 14399 33638 14445 33676
rect 14399 33604 14405 33638
rect 14439 33604 14445 33638
rect 14399 33566 14445 33604
rect 14399 33532 14405 33566
rect 14439 33532 14445 33566
rect 14399 33494 14445 33532
rect 14399 33460 14405 33494
rect 14439 33460 14445 33494
rect 14399 33422 14445 33460
rect 14399 33388 14405 33422
rect 14439 33388 14445 33422
rect 14399 33350 14445 33388
rect 14399 33316 14405 33350
rect 14439 33316 14445 33350
rect 14399 33278 14445 33316
rect 14399 33244 14405 33278
rect 14439 33244 14445 33278
rect 14399 33206 14445 33244
rect 14399 33172 14405 33206
rect 14439 33172 14445 33206
rect 14399 33134 14445 33172
rect 14399 33100 14405 33134
rect 14439 33100 14445 33134
rect 14399 33062 14445 33100
rect 14399 33028 14405 33062
rect 14439 33028 14445 33062
rect 14399 32990 14445 33028
rect 14399 32956 14405 32990
rect 14439 32956 14445 32990
rect 14399 32918 14445 32956
rect 14399 32884 14405 32918
rect 14439 32884 14445 32918
rect 14399 32846 14445 32884
rect 14399 32812 14405 32846
rect 14439 32812 14445 32846
rect 14399 32774 14445 32812
rect 14399 32740 14405 32774
rect 14439 32740 14445 32774
rect 14399 32702 14445 32740
rect 14399 32668 14405 32702
rect 14439 32668 14445 32702
rect 14399 32630 14445 32668
rect 14399 32596 14405 32630
rect 14439 32596 14445 32630
rect 14399 32558 14445 32596
rect 14399 32524 14405 32558
rect 14439 32524 14445 32558
rect 14399 32486 14445 32524
rect 14399 32452 14405 32486
rect 14439 32452 14445 32486
rect 14399 32414 14445 32452
rect 14399 32380 14405 32414
rect 14439 32380 14445 32414
rect 14399 32342 14445 32380
rect 14399 32308 14405 32342
rect 14439 32308 14445 32342
rect 14399 32270 14445 32308
rect 14399 32236 14405 32270
rect 14439 32236 14445 32270
rect 14399 32198 14445 32236
rect 14399 32164 14405 32198
rect 14439 32164 14445 32198
rect 14399 32126 14445 32164
rect 14399 32092 14405 32126
rect 14439 32092 14445 32126
rect 14399 32054 14445 32092
rect 14399 32020 14405 32054
rect 14439 32020 14445 32054
rect 14399 31982 14445 32020
rect 14399 31948 14405 31982
rect 14439 31948 14445 31982
rect 14399 31910 14445 31948
rect 14399 31876 14405 31910
rect 14439 31876 14445 31910
rect 14399 31838 14445 31876
rect 14399 31804 14405 31838
rect 14439 31804 14445 31838
rect 14399 31766 14445 31804
rect 14399 31732 14405 31766
rect 14439 31732 14445 31766
rect 14399 31694 14445 31732
rect 14399 31660 14405 31694
rect 14439 31660 14445 31694
rect 14399 31622 14445 31660
rect 14399 31588 14405 31622
rect 14439 31588 14445 31622
rect 14399 31550 14445 31588
rect 14399 31516 14405 31550
rect 14439 31516 14445 31550
rect 14399 31478 14445 31516
rect 14399 31444 14405 31478
rect 14439 31444 14445 31478
rect 14399 31406 14445 31444
rect 14399 31372 14405 31406
rect 14439 31372 14445 31406
rect 14399 31334 14445 31372
rect 14399 31300 14405 31334
rect 14439 31300 14445 31334
rect 14399 31262 14445 31300
rect 14399 31228 14405 31262
rect 14439 31228 14445 31262
rect 14399 31190 14445 31228
rect 14399 31156 14405 31190
rect 14439 31156 14445 31190
rect 14399 31118 14445 31156
rect 14399 31084 14405 31118
rect 14439 31084 14445 31118
rect 14399 31046 14445 31084
rect 14399 31012 14405 31046
rect 14439 31012 14445 31046
rect 14399 30974 14445 31012
rect 14399 30940 14405 30974
rect 14439 30940 14445 30974
rect 14399 30902 14445 30940
rect 14399 30868 14405 30902
rect 14439 30868 14445 30902
rect 14399 30830 14445 30868
rect 14399 30796 14405 30830
rect 14439 30796 14445 30830
rect 14399 30758 14445 30796
rect 14399 30724 14405 30758
rect 14439 30724 14445 30758
rect 14399 30686 14445 30724
rect 14399 30652 14405 30686
rect 14439 30652 14445 30686
rect 14399 30614 14445 30652
rect 14399 30580 14405 30614
rect 14439 30580 14445 30614
rect 14399 30542 14445 30580
rect 14399 30508 14405 30542
rect 14439 30508 14445 30542
rect 14399 30470 14445 30508
rect 14399 30436 14405 30470
rect 14439 30436 14445 30470
rect 14399 30398 14445 30436
rect 14399 30364 14405 30398
rect 14439 30364 14445 30398
rect 14399 30326 14445 30364
rect 14399 30292 14405 30326
rect 14439 30292 14445 30326
rect 14399 30254 14445 30292
rect 14399 30220 14405 30254
rect 14439 30220 14445 30254
rect 14399 30182 14445 30220
rect 14399 30148 14405 30182
rect 14439 30148 14445 30182
rect 14399 30110 14445 30148
rect 14399 30076 14405 30110
rect 14439 30076 14445 30110
rect 14399 30038 14445 30076
rect 14399 30004 14405 30038
rect 14439 30004 14445 30038
rect 14399 29966 14445 30004
rect 14399 29932 14405 29966
rect 14439 29932 14445 29966
rect 14399 29894 14445 29932
rect 14399 29860 14405 29894
rect 14439 29860 14445 29894
rect 14399 29822 14445 29860
rect 14399 29788 14405 29822
rect 14439 29788 14445 29822
rect 14399 29750 14445 29788
rect 14399 29716 14405 29750
rect 14439 29716 14445 29750
rect 14399 29678 14445 29716
rect 14399 29644 14405 29678
rect 14439 29644 14445 29678
rect 14399 29606 14445 29644
rect 14399 29572 14405 29606
rect 14439 29572 14445 29606
rect 14399 29534 14445 29572
rect 14399 29500 14405 29534
rect 14439 29500 14445 29534
rect 14399 29462 14445 29500
rect 14399 29428 14405 29462
rect 14439 29428 14445 29462
rect 14399 29390 14445 29428
rect 14399 29356 14405 29390
rect 14439 29356 14445 29390
rect 14399 29318 14445 29356
rect 14399 29284 14405 29318
rect 14439 29284 14445 29318
rect 14399 29246 14445 29284
rect 14399 29212 14405 29246
rect 14439 29212 14445 29246
rect 14399 29174 14445 29212
rect 14399 29140 14405 29174
rect 14439 29140 14445 29174
rect 14399 29102 14445 29140
rect 14399 29068 14405 29102
rect 14439 29068 14445 29102
rect 14399 29030 14445 29068
rect 14399 28996 14405 29030
rect 14439 28996 14445 29030
rect 14399 28958 14445 28996
rect 14399 28924 14405 28958
rect 14439 28924 14445 28958
rect 14399 28886 14445 28924
rect 14399 28852 14405 28886
rect 14439 28852 14445 28886
rect 14399 28814 14445 28852
rect 14399 28780 14405 28814
rect 14439 28780 14445 28814
rect 14399 28742 14445 28780
rect 14399 28708 14405 28742
rect 14439 28708 14445 28742
rect 14399 28670 14445 28708
rect 14399 28636 14405 28670
rect 14439 28636 14445 28670
rect 14399 28598 14445 28636
rect 14399 28564 14405 28598
rect 14439 28564 14445 28598
rect 14399 28526 14445 28564
rect 14399 28492 14405 28526
rect 14439 28492 14445 28526
rect 14399 28454 14445 28492
rect 14399 28420 14405 28454
rect 14439 28420 14445 28454
rect 14399 28382 14445 28420
rect 14399 28348 14405 28382
rect 14439 28348 14445 28382
rect 14399 28310 14445 28348
rect 14399 28276 14405 28310
rect 14439 28276 14445 28310
rect 14399 28238 14445 28276
rect 14399 28204 14405 28238
rect 14439 28204 14445 28238
rect 14399 28166 14445 28204
rect 14399 28132 14405 28166
rect 14439 28132 14445 28166
rect 14399 28094 14445 28132
rect 14399 28060 14405 28094
rect 14439 28060 14445 28094
rect 14399 28022 14445 28060
rect 14399 27988 14405 28022
rect 14439 27988 14445 28022
rect 14399 27950 14445 27988
rect 14399 27916 14405 27950
rect 14439 27916 14445 27950
rect 14399 27878 14445 27916
rect 14399 27844 14405 27878
rect 14439 27844 14445 27878
rect 14399 27806 14445 27844
rect 14399 27772 14405 27806
rect 14439 27772 14445 27806
rect 9783 27490 9829 27542
rect 9783 27456 9789 27490
rect 9823 27456 9829 27490
rect 9783 27418 9829 27456
rect 9783 27384 9789 27418
rect 9823 27384 9829 27418
rect 9783 27346 9829 27384
rect 9783 27312 9789 27346
rect 9823 27312 9829 27346
rect 9783 27274 9829 27312
rect 9783 27240 9789 27274
rect 9823 27240 9829 27274
rect 9783 27202 9829 27240
rect 9783 27168 9789 27202
rect 9823 27168 9829 27202
rect 11948 27516 12203 27749
rect 14399 27734 14445 27772
rect 14399 27700 14405 27734
rect 14439 27700 14445 27734
rect 14399 27662 14445 27700
rect 14399 27628 14405 27662
rect 14439 27628 14445 27662
rect 14399 27542 14445 27628
rect 11948 27482 11960 27516
rect 11994 27482 12059 27516
rect 12093 27482 12157 27516
rect 12191 27482 12203 27516
rect 9783 27130 9829 27168
rect 9783 27096 9789 27130
rect 9823 27096 9829 27130
rect 9783 27058 9829 27096
rect 9783 27024 9789 27058
rect 9823 27024 9829 27058
rect 10099 27158 10145 27170
rect 10099 27124 10105 27158
rect 10139 27128 10145 27158
rect 10139 27124 10506 27128
rect 10099 27086 10506 27124
rect 10099 27052 10105 27086
rect 10139 27076 10506 27086
rect 10558 27076 10570 27128
rect 10622 27076 10628 27128
rect 10139 27052 10145 27076
rect 10099 27040 10145 27052
rect 9783 26986 9829 27024
rect 9783 26952 9789 26986
rect 9823 26952 9829 26986
rect 9783 26914 9829 26952
rect 9783 26880 9789 26914
rect 9823 26880 9829 26914
rect 9783 26842 9829 26880
rect 9783 26808 9789 26842
rect 9823 26808 9829 26842
rect 9783 26770 9829 26808
rect 9783 26736 9789 26770
rect 9823 26736 9829 26770
rect 9783 26698 9829 26736
rect 9783 26664 9789 26698
rect 9823 26664 9829 26698
rect 9783 26626 9829 26664
rect 9783 26592 9789 26626
rect 9823 26592 9829 26626
rect 11948 26660 12203 27482
rect 11948 26626 11960 26660
rect 11994 26626 12059 26660
rect 12093 26626 12157 26660
rect 12191 26626 12203 26660
rect 11948 26620 12203 26626
rect 12426 27536 14445 27542
rect 12426 27530 12510 27536
rect 12426 27496 12432 27530
rect 12466 27502 12510 27530
rect 12544 27502 12582 27536
rect 12616 27502 12654 27536
rect 12688 27502 12726 27536
rect 12760 27502 12798 27536
rect 12832 27502 12870 27536
rect 12904 27502 12942 27536
rect 12976 27502 13014 27536
rect 13048 27502 13086 27536
rect 13120 27502 13158 27536
rect 13192 27502 13230 27536
rect 13264 27502 13302 27536
rect 13336 27502 13374 27536
rect 13408 27502 13446 27536
rect 13480 27502 13518 27536
rect 13552 27502 13590 27536
rect 13624 27502 13662 27536
rect 13696 27502 13734 27536
rect 13768 27502 13806 27536
rect 13840 27502 13878 27536
rect 13912 27502 13950 27536
rect 13984 27502 14022 27536
rect 14056 27502 14094 27536
rect 14128 27502 14183 27536
rect 14217 27502 14255 27536
rect 14289 27502 14327 27536
rect 14361 27502 14399 27536
rect 14433 27502 14445 27536
rect 12466 27496 14445 27502
rect 12426 27458 12472 27496
rect 12426 27424 12432 27458
rect 12466 27424 12472 27458
rect 12426 27386 12472 27424
rect 12426 27352 12432 27386
rect 12466 27352 12472 27386
rect 12426 27314 12472 27352
rect 12426 27280 12432 27314
rect 12466 27280 12472 27314
rect 12426 27242 12472 27280
rect 12426 27208 12432 27242
rect 12466 27208 12472 27242
rect 12426 27170 12472 27208
rect 12426 27136 12432 27170
rect 12466 27136 12472 27170
rect 12426 27098 12472 27136
rect 12426 27064 12432 27098
rect 12466 27064 12472 27098
rect 12426 27026 12472 27064
rect 12426 26992 12432 27026
rect 12466 26992 12472 27026
rect 12426 26954 12472 26992
rect 12426 26920 12432 26954
rect 12466 26920 12472 26954
rect 12426 26882 12472 26920
rect 12426 26848 12432 26882
rect 12466 26848 12472 26882
rect 12426 26810 12472 26848
rect 12426 26776 12432 26810
rect 12466 26776 12472 26810
rect 12426 26738 12472 26776
rect 12426 26704 12432 26738
rect 12466 26704 12472 26738
rect 12426 26666 12472 26704
rect 12426 26632 12432 26666
rect 12466 26632 12472 26666
rect 9783 26554 9829 26592
rect 9783 26520 9789 26554
rect 9823 26520 9829 26554
rect 9783 26482 9829 26520
rect 9783 26448 9789 26482
rect 9823 26448 9829 26482
rect 9783 26410 9829 26448
rect 12426 26594 12472 26632
rect 12426 26560 12432 26594
rect 12466 26560 12472 26594
rect 12426 26522 12472 26560
rect 12426 26488 12432 26522
rect 12466 26488 12472 26522
rect 12426 26410 12472 26488
rect 9783 26376 9789 26410
rect 9823 26404 12472 26410
rect 9823 26376 9906 26404
rect 9783 26370 9906 26376
rect 9940 26370 9978 26404
rect 10012 26370 10050 26404
rect 10084 26370 10122 26404
rect 10156 26370 10194 26404
rect 10228 26370 10266 26404
rect 10300 26370 10338 26404
rect 10372 26370 10410 26404
rect 10444 26370 10482 26404
rect 10516 26370 10554 26404
rect 10588 26370 10626 26404
rect 10660 26370 10698 26404
rect 10732 26370 10770 26404
rect 10804 26370 10842 26404
rect 10876 26370 10914 26404
rect 10948 26370 10986 26404
rect 11020 26370 11058 26404
rect 11092 26370 11130 26404
rect 11164 26370 11202 26404
rect 11236 26370 11274 26404
rect 11308 26370 11346 26404
rect 11380 26370 11418 26404
rect 11452 26370 11490 26404
rect 11524 26370 11562 26404
rect 11596 26370 11634 26404
rect 11668 26370 11706 26404
rect 11740 26370 11778 26404
rect 11812 26370 11850 26404
rect 11884 26370 11922 26404
rect 11956 26370 11994 26404
rect 12028 26370 12066 26404
rect 12100 26370 12138 26404
rect 12172 26370 12210 26404
rect 12244 26370 12282 26404
rect 12316 26370 12354 26404
rect 12388 26370 12426 26404
rect 12460 26370 12472 26404
rect 9783 26364 12472 26370
rect -242 17223 -236 17275
rect -184 17223 -172 17275
rect -120 17229 189 17275
tri 1076 17229 1122 17275 se
rect 1122 17229 2223 17275
rect -120 17223 -114 17229
tri -114 17223 -108 17229 nw
tri 1070 17223 1076 17229 se
rect 1076 17223 2223 17229
tri 1048 17201 1070 17223 se
rect 1070 17201 2223 17223
rect -29 17195 955 17201
rect 151 17189 212 17195
rect 164 17161 212 17189
rect 246 17161 284 17195
rect 318 17161 488 17195
rect 522 17161 560 17195
rect 594 17161 836 17195
rect 870 17161 908 17195
rect 942 17161 955 17195
rect 164 17155 955 17161
rect 151 17120 920 17155
tri 920 17120 955 17155 nw
tri 967 17120 1048 17201 se
rect 1048 17120 2223 17201
rect 151 17117 901 17120
rect 164 17101 901 17117
tri 901 17101 920 17120 nw
tri 948 17101 967 17120 se
rect 967 17101 2223 17120
rect 164 17083 170 17101
rect 151 17079 170 17083
rect -29 17073 170 17079
tri 170 17076 195 17101 nw
tri 923 17076 948 17101 se
rect 948 17076 2223 17101
tri 920 17073 923 17076 se
rect 923 17073 2223 17076
tri -29 17045 -1 17073 ne
rect -1 17045 170 17073
tri -1 17011 33 17045 ne
rect 33 17011 130 17045
rect 164 17011 170 17045
tri 33 16973 71 17011 ne
rect 71 16973 170 17011
tri 71 16939 105 16973 ne
rect 105 16939 130 16973
rect 164 16939 170 16973
rect 207 17067 2223 17073
rect 387 16951 2223 17067
rect 207 16942 2223 16951
tri 2809 16945 2852 16988 se
rect 2852 16945 2982 16988
tri 2806 16942 2809 16945 se
rect 2809 16942 2982 16945
tri 2803 16939 2806 16942 se
rect 2806 16939 2982 16942
tri 105 16927 117 16939 ne
rect 117 16927 170 16939
tri 170 16927 182 16939 sw
tri 2793 16929 2803 16939 se
rect 2803 16938 2982 16939
rect 2803 16929 2973 16938
tri 2973 16929 2982 16938 nw
rect 4920 16942 4991 16988
tri 4920 16929 4933 16942 ne
rect 4933 16929 4991 16942
tri 117 16922 122 16927 ne
rect 122 16922 182 16927
tri 182 16922 187 16927 sw
rect 2793 16923 2961 16929
rect 122 16914 187 16922
tri 187 16914 195 16922 sw
rect 122 16908 787 16914
rect 122 16874 261 16908
rect 295 16874 333 16908
rect 367 16875 787 16908
rect 367 16874 379 16875
rect 122 16873 379 16874
rect 174 16868 379 16873
tri 379 16868 386 16875 nw
tri 459 16868 466 16875 ne
rect 466 16868 787 16875
rect 174 16847 178 16868
tri 178 16847 199 16868 nw
tri 1285 16847 1306 16868 ne
rect 1306 16862 1375 16868
tri 1375 16862 1381 16868 nw
tri 2298 16862 2304 16868 ne
rect 2304 16862 2310 16914
rect 2362 16862 2374 16914
rect 2426 16862 2438 16914
rect 2490 16862 2502 16914
rect 2554 16874 2560 16914
rect 2554 16865 2563 16874
tri 2563 16865 2572 16874 nw
rect 2845 16871 2857 16923
rect 2909 16917 2961 16923
tri 2961 16917 2973 16929 nw
tri 4933 16917 4945 16929 ne
rect 2793 16865 2909 16871
tri 2909 16865 2961 16917 nw
rect 4828 16893 4896 16914
tri 4896 16893 4917 16914 sw
rect 4828 16868 4917 16893
tri 3655 16865 3658 16868 ne
rect 3658 16865 3726 16868
rect 2554 16862 2560 16865
tri 2560 16862 2563 16865 nw
tri 3658 16862 3661 16865 ne
rect 3661 16862 3726 16865
rect 1306 16847 1360 16862
tri 1360 16847 1375 16862 nw
tri 3661 16847 3676 16862 ne
rect 3676 16847 3726 16862
tri 174 16843 178 16847 nw
rect 398 16835 444 16847
tri 1306 16843 1310 16847 ne
rect 398 16801 404 16835
rect 438 16801 444 16835
rect 398 16784 444 16801
tri 444 16784 469 16809 sw
tri 1285 16784 1310 16809 se
rect 1310 16784 1356 16847
tri 1356 16843 1360 16847 nw
tri 3676 16843 3680 16847 ne
tri 1356 16784 1381 16809 sw
tri 3655 16784 3680 16809 se
rect 3680 16784 3726 16847
tri 3726 16843 3751 16868 nw
tri 4837 16843 4862 16868 ne
tri 3726 16784 3751 16809 sw
rect 398 16763 469 16784
rect 398 16729 404 16763
rect 438 16738 469 16763
rect 470 16739 471 16783
rect 507 16739 508 16783
rect 509 16778 1244 16784
rect 1246 16783 1282 16784
rect 509 16744 560 16778
rect 594 16744 632 16778
rect 666 16744 704 16778
rect 738 16744 776 16778
rect 810 16744 944 16778
rect 978 16744 1016 16778
rect 1050 16744 1088 16778
rect 1122 16744 1160 16778
rect 1194 16744 1244 16778
rect 509 16738 1244 16744
rect 1245 16739 1283 16783
rect 1246 16738 1282 16739
rect 1284 16738 1382 16784
rect 1384 16783 1420 16784
rect 1383 16739 1421 16783
rect 1422 16778 2157 16784
rect 1422 16744 1472 16778
rect 1506 16744 1544 16778
rect 1578 16744 1616 16778
rect 1650 16744 1688 16778
rect 1722 16744 1856 16778
rect 1890 16744 1928 16778
rect 1962 16744 2000 16778
rect 2034 16744 2072 16778
rect 2106 16744 2157 16778
rect 1384 16738 1420 16739
rect 1422 16738 2157 16744
rect 2158 16739 2159 16783
rect 2195 16739 2196 16783
rect 2197 16738 2268 16784
rect 438 16729 444 16738
rect 398 16654 444 16729
tri 444 16713 469 16738 nw
tri 2197 16713 2222 16738 ne
tri 444 16654 469 16679 sw
tri 2197 16654 2222 16679 se
rect 2222 16654 2268 16738
rect 2768 16738 2839 16784
rect 2840 16739 2841 16783
rect 2877 16739 2878 16783
rect 2879 16778 3614 16784
rect 3616 16783 3652 16784
rect 2879 16744 2930 16778
rect 2964 16744 3002 16778
rect 3036 16744 3074 16778
rect 3108 16744 3146 16778
rect 3180 16744 3314 16778
rect 3348 16744 3386 16778
rect 3420 16744 3458 16778
rect 3492 16744 3530 16778
rect 3564 16744 3614 16778
rect 2879 16738 3614 16744
rect 3615 16739 3653 16783
rect 3616 16738 3652 16739
rect 3654 16738 3752 16784
rect 3754 16783 3790 16784
rect 3753 16739 3791 16783
rect 3792 16778 4527 16784
rect 3792 16744 3842 16778
rect 3876 16744 3914 16778
rect 3948 16744 3986 16778
rect 4020 16744 4058 16778
rect 4092 16744 4226 16778
rect 4260 16744 4298 16778
rect 4332 16744 4370 16778
rect 4404 16744 4442 16778
rect 4476 16744 4527 16778
rect 3754 16738 3790 16739
rect 3792 16738 4527 16744
rect 4528 16739 4529 16783
rect 4565 16739 4566 16783
rect 4567 16738 4638 16784
tri 2268 16654 2293 16679 sw
tri 2743 16654 2768 16679 se
rect 2768 16654 2814 16738
tri 2814 16713 2839 16738 nw
tri 4567 16713 4592 16738 ne
tri 2814 16654 2839 16679 sw
tri 4567 16654 4592 16679 se
rect 4592 16654 4638 16738
rect 398 16648 4638 16654
rect 398 16608 4295 16648
tri 601 16583 626 16608 ne
rect 242 16535 444 16553
rect 288 15325 398 16535
rect 242 15221 444 15325
rect 288 13795 398 15221
tri 621 13795 626 13800 se
rect 626 13795 672 16608
tri 672 16583 697 16608 nw
tri 1057 16583 1082 16608 ne
rect 854 15293 900 15345
rect 855 15291 899 15292
rect 855 15254 899 15255
rect 854 15201 900 15253
tri 672 13795 677 13800 sw
rect 242 13691 444 13795
tri 601 13775 621 13795 se
rect 621 13775 677 13795
tri 677 13775 697 13795 sw
rect 482 13763 816 13775
rect 482 13729 488 13763
rect 522 13729 560 13763
rect 594 13729 632 13763
rect 666 13729 704 13763
rect 738 13729 776 13763
rect 810 13729 816 13763
rect 482 13717 816 13729
rect 854 13763 900 13815
tri 1057 13775 1082 13800 se
rect 1082 13795 1128 16608
tri 1128 16583 1153 16608 nw
tri 1513 16583 1538 16608 ne
rect 1356 16521 1449 16535
rect 1310 15183 1449 15369
rect 1356 13804 1365 13839
tri 1365 13804 1400 13839 nw
rect 1356 13800 1361 13804
tri 1361 13800 1365 13804 nw
tri 1128 13795 1133 13800 sw
tri 1356 13795 1361 13800 nw
tri 1533 13795 1538 13800 se
rect 1538 13795 1584 16608
tri 1584 16583 1609 16608 nw
tri 1969 16583 1994 16608 ne
rect 1766 15293 1812 15345
rect 1767 15291 1811 15292
rect 1767 15254 1811 15255
rect 1766 15201 1812 15253
tri 1584 13795 1589 13800 sw
rect 1082 13775 1133 13795
tri 1133 13775 1153 13795 sw
rect 855 13761 899 13762
rect 854 13725 900 13761
rect 855 13724 899 13725
tri 601 13692 626 13717 ne
rect 288 12265 398 13691
tri 621 12265 626 12270 se
rect 626 12265 672 13717
tri 672 13692 697 13717 nw
rect 854 13671 900 13723
rect 938 13763 1272 13775
rect 938 13729 944 13763
rect 978 13729 1016 13763
rect 1050 13729 1088 13763
rect 1122 13729 1160 13763
rect 1194 13729 1232 13763
rect 1266 13729 1272 13763
rect 938 13717 1272 13729
tri 1057 13692 1082 13717 ne
tri 672 12265 677 12270 sw
tri 601 12245 621 12265 se
rect 621 12245 677 12265
tri 677 12245 697 12265 sw
rect 482 12233 816 12245
rect 482 12199 488 12233
rect 522 12199 560 12233
rect 594 12199 632 12233
rect 666 12199 704 12233
rect 738 12199 776 12233
rect 810 12199 816 12233
rect 482 12187 816 12199
rect 854 12233 900 12285
tri 1057 12245 1082 12270 se
rect 1082 12265 1128 13717
tri 1128 13692 1153 13717 nw
rect 1310 13691 1356 13795
tri 1513 13775 1533 13795 se
rect 1533 13775 1589 13795
tri 1589 13775 1609 13795 sw
rect 1394 13763 1728 13775
rect 1394 13729 1400 13763
rect 1434 13729 1472 13763
rect 1506 13729 1544 13763
rect 1578 13729 1616 13763
rect 1650 13729 1688 13763
rect 1722 13729 1728 13763
rect 1394 13717 1728 13729
rect 1766 13763 1812 13815
tri 1969 13775 1994 13800 se
rect 1994 13795 2040 16608
tri 2040 16583 2065 16608 nw
tri 2971 16583 2996 16608 ne
rect 2222 16535 2424 16553
rect 2459 16535 2460 16553
rect 2576 16535 2577 16553
rect 2612 16535 2649 16553
rect 2658 16535 2814 16553
rect 2268 15325 2378 16535
rect 2658 15325 2768 16535
rect 2222 15221 2424 15325
rect 2612 15221 2814 15325
tri 2040 13795 2045 13800 sw
rect 2268 13795 2378 15221
rect 2658 13795 2768 15221
tri 2991 13795 2996 13800 se
rect 2996 13795 3042 16608
tri 3042 16583 3067 16608 nw
tri 3427 16583 3452 16608 ne
rect 3224 15293 3270 15345
rect 3225 15291 3269 15292
rect 3225 15254 3269 15255
rect 3224 15201 3270 15253
tri 3042 13795 3047 13800 sw
rect 1994 13775 2045 13795
tri 2045 13775 2065 13795 sw
rect 1767 13761 1811 13762
rect 1766 13725 1812 13761
rect 1767 13724 1811 13725
tri 1513 13692 1538 13717 ne
tri 1356 13671 1376 13691 sw
rect 1356 13659 1376 13671
tri 1376 13659 1388 13671 sw
rect 1356 13653 1388 13659
tri 1388 13653 1394 13659 sw
rect 1356 12285 1376 12309
tri 1376 12285 1400 12309 nw
rect 1356 12270 1361 12285
tri 1361 12270 1376 12285 nw
tri 1128 12265 1133 12270 sw
tri 1356 12265 1361 12270 nw
tri 1533 12265 1538 12270 se
rect 1538 12265 1584 13717
tri 1584 13692 1609 13717 nw
rect 1766 13671 1812 13723
rect 1850 13763 2184 13775
rect 1850 13729 1856 13763
rect 1890 13729 1928 13763
rect 1962 13729 2000 13763
rect 2034 13729 2072 13763
rect 2106 13729 2144 13763
rect 2178 13729 2184 13763
rect 1850 13717 2184 13729
tri 1969 13692 1994 13717 ne
tri 1584 12265 1589 12270 sw
rect 1082 12245 1133 12265
tri 1133 12245 1153 12265 sw
tri 1513 12245 1533 12265 se
rect 1533 12245 1589 12265
tri 1589 12245 1609 12265 sw
rect 855 12231 899 12232
rect 854 12195 900 12231
rect 855 12194 899 12195
tri 532 12179 540 12187 ne
rect 540 12179 615 12187
tri 174 12162 191 12179 sw
tri 540 12162 557 12179 ne
rect 174 12154 191 12162
tri 191 12154 199 12162 sw
rect 167 12148 513 12154
rect 167 12137 179 12148
rect 122 12114 179 12137
rect 213 12114 251 12148
rect 285 12114 323 12148
rect 357 12114 395 12148
rect 429 12114 467 12148
rect 501 12114 513 12148
rect 122 9739 513 12114
rect 557 9879 615 12179
tri 615 12162 640 12187 nw
rect 854 12153 900 12193
rect 938 12233 1272 12245
rect 938 12199 944 12233
rect 978 12199 1016 12233
rect 1050 12199 1088 12233
rect 1122 12199 1160 12233
rect 1194 12199 1232 12233
rect 1266 12199 1272 12233
rect 938 12187 1272 12199
rect 1394 12233 1728 12245
rect 1394 12199 1400 12233
rect 1434 12199 1472 12233
rect 1506 12199 1544 12233
rect 1578 12199 1616 12233
rect 1650 12199 1688 12233
rect 1722 12199 1728 12233
rect 1394 12187 1728 12199
rect 1766 12233 1812 12285
tri 1969 12245 1994 12270 se
rect 1994 12245 2040 13717
tri 2040 13692 2065 13717 nw
rect 2222 13691 2424 13795
rect 2612 13691 2814 13795
tri 2971 13775 2991 13795 se
rect 2991 13775 3047 13795
tri 3047 13775 3067 13795 sw
rect 2852 13763 3186 13775
rect 2852 13729 2858 13763
rect 2892 13729 2930 13763
rect 2964 13729 3002 13763
rect 3036 13729 3074 13763
rect 3108 13729 3146 13763
rect 3180 13729 3186 13763
rect 2852 13717 3186 13729
rect 3224 13763 3270 13815
tri 3427 13775 3452 13800 se
rect 3452 13795 3498 16608
tri 3498 16583 3523 16608 nw
tri 3883 16583 3908 16608 ne
tri 3645 16524 3656 16535 se
rect 3656 16524 3680 16535
rect 3645 16521 3680 16524
rect 3726 16524 3750 16535
tri 3750 16524 3761 16535 sw
rect 3726 16521 3761 16524
rect 3645 15183 3761 15369
rect 3645 13830 3680 13839
tri 3645 13815 3660 13830 ne
rect 3660 13815 3680 13830
tri 3660 13804 3671 13815 ne
rect 3671 13804 3680 13815
tri 3671 13800 3675 13804 ne
rect 3675 13800 3680 13804
tri 3498 13795 3503 13800 sw
tri 3675 13795 3680 13800 ne
rect 3726 13830 3761 13839
rect 3726 13815 3746 13830
tri 3746 13815 3761 13830 nw
rect 3726 13804 3735 13815
tri 3735 13804 3746 13815 nw
tri 3726 13795 3735 13804 nw
tri 3903 13795 3908 13800 se
rect 3908 13795 3954 16608
tri 3954 16583 3979 16608 nw
tri 4213 16583 4238 16608 ne
rect 4238 16596 4295 16608
rect 4347 16608 4638 16648
rect 4347 16596 4410 16608
rect 4238 16584 4410 16596
rect 4238 16583 4295 16584
tri 4238 16553 4268 16583 ne
rect 4268 16553 4295 16583
tri 4268 16535 4286 16553 ne
rect 4286 16535 4295 16553
tri 4286 16526 4295 16535 ne
rect 4347 16532 4410 16584
tri 4410 16583 4435 16608 nw
rect 4295 16526 4410 16532
tri 4295 16521 4300 16526 ne
rect 4300 16521 4410 16526
tri 4300 16457 4364 16521 ne
rect 4136 15293 4182 15345
rect 4137 15291 4181 15292
rect 4137 15254 4181 15255
rect 4136 15201 4182 15253
tri 3954 13795 3959 13800 sw
rect 3452 13775 3503 13795
tri 3503 13775 3523 13795 sw
rect 3225 13761 3269 13762
rect 3224 13725 3270 13761
rect 3225 13724 3269 13725
tri 2971 13692 2996 13717 ne
tri 2040 12245 2065 12270 sw
rect 2268 12265 2378 13691
rect 2658 12265 2768 13691
tri 2991 12265 2996 12270 se
rect 2996 12265 3042 13717
tri 3042 13692 3067 13717 nw
rect 3224 13659 3270 13723
rect 3308 13763 3642 13775
rect 3308 13729 3314 13763
rect 3348 13729 3386 13763
rect 3420 13729 3458 13763
rect 3492 13729 3530 13763
rect 3564 13729 3602 13763
rect 3636 13729 3642 13763
rect 3308 13717 3642 13729
tri 3427 13692 3452 13717 ne
rect 3224 13625 3230 13659
rect 3264 13625 3270 13659
rect 3224 13584 3270 13625
rect 3224 13550 3230 13584
rect 3264 13550 3270 13584
rect 3224 13508 3270 13550
rect 3224 13474 3230 13508
rect 3264 13474 3270 13508
rect 3224 13432 3270 13474
rect 3224 13398 3230 13432
rect 3264 13398 3270 13432
rect 3224 13356 3270 13398
rect 3224 13322 3230 13356
rect 3264 13322 3270 13356
rect 3224 13280 3270 13322
rect 3224 13246 3230 13280
rect 3264 13246 3270 13280
rect 3224 13204 3270 13246
rect 3224 13170 3230 13204
rect 3264 13170 3270 13204
rect 3224 13128 3270 13170
rect 3224 13094 3230 13128
rect 3264 13094 3270 13128
rect 3224 13052 3270 13094
rect 3224 13018 3230 13052
rect 3264 13018 3270 13052
rect 3224 12976 3270 13018
rect 3224 12942 3230 12976
rect 3264 12942 3270 12976
rect 3224 12900 3270 12942
rect 3224 12866 3230 12900
rect 3264 12866 3270 12900
rect 3224 12824 3270 12866
rect 3224 12790 3230 12824
rect 3264 12790 3270 12824
rect 3224 12748 3270 12790
rect 3224 12714 3230 12748
rect 3264 12714 3270 12748
rect 3224 12672 3270 12714
rect 3224 12638 3230 12672
rect 3264 12638 3270 12672
rect 3224 12596 3270 12638
rect 3224 12562 3230 12596
rect 3264 12562 3270 12596
rect 3224 12520 3270 12562
rect 3224 12486 3230 12520
rect 3264 12486 3270 12520
rect 3224 12444 3270 12486
rect 3224 12410 3230 12444
rect 3264 12410 3270 12444
rect 3224 12368 3270 12410
rect 3224 12334 3230 12368
rect 3264 12334 3270 12368
rect 3224 12270 3270 12334
tri 2971 12245 2991 12265 se
rect 2991 12245 3042 12265
tri 3042 12245 3067 12270 sw
tri 3451 12269 3452 12270 se
rect 3452 12269 3498 13717
tri 3498 13692 3523 13717 nw
rect 3680 13691 3726 13795
tri 3883 13775 3903 13795 se
rect 3903 13775 3959 13795
tri 3959 13775 3979 13795 sw
rect 3764 13763 4098 13775
rect 3764 13729 3770 13763
rect 3804 13729 3842 13763
rect 3876 13729 3914 13763
rect 3948 13729 3986 13763
rect 4020 13729 4058 13763
rect 4092 13729 4098 13763
rect 3764 13717 4098 13729
rect 4136 13763 4182 13815
tri 4339 13775 4364 13800 se
rect 4364 13795 4410 16521
rect 4638 16535 4794 16553
rect 4638 15325 4748 16535
rect 4592 15221 4794 15325
tri 4410 13795 4415 13800 sw
rect 4638 13795 4748 15221
rect 4364 13775 4415 13795
tri 4415 13775 4435 13795 sw
rect 4137 13761 4181 13762
rect 4136 13725 4182 13761
rect 4137 13724 4181 13725
tri 3883 13692 3908 13717 ne
tri 3645 13656 3680 13691 se
rect 3645 13653 3680 13656
tri 3726 13671 3746 13691 sw
rect 3726 13656 3746 13671
tri 3746 13656 3761 13671 sw
rect 3726 13653 3761 13656
rect 3645 12300 3680 12309
tri 3645 12270 3675 12300 ne
rect 3675 12270 3680 12300
rect 3225 12268 3269 12269
tri 3450 12268 3451 12269 se
rect 3451 12268 3498 12269
rect 1767 12231 1811 12232
rect 1766 12195 1812 12231
rect 1767 12194 1811 12195
tri 900 12153 925 12178 sw
tri 1741 12153 1766 12178 se
rect 1766 12153 1812 12193
rect 1850 12233 2184 12245
rect 2852 12233 3186 12245
rect 1850 12199 1856 12233
rect 1890 12199 1928 12233
rect 1962 12199 2000 12233
rect 2034 12199 2072 12233
rect 2106 12199 2144 12233
rect 2178 12199 2184 12233
tri 2184 12199 2203 12218 sw
rect 1850 12187 2203 12199
tri 2203 12187 2215 12199 sw
tri 2140 12176 2151 12187 ne
rect 2151 12178 2215 12187
tri 2215 12178 2224 12187 sw
tri 2458 12178 2459 12179 se
rect 2459 12178 2577 12233
tri 2833 12199 2852 12218 se
rect 2852 12199 2858 12233
rect 2892 12199 2930 12233
rect 2964 12199 3002 12233
rect 3036 12199 3074 12233
rect 3108 12199 3146 12233
rect 3180 12199 3186 12233
tri 2821 12187 2833 12199 se
rect 2833 12187 3186 12199
rect 3224 12232 3270 12268
tri 3427 12245 3450 12268 se
rect 3450 12265 3498 12268
tri 3498 12265 3503 12270 sw
tri 3675 12265 3680 12270 ne
rect 3726 12300 3761 12309
rect 3726 12285 3746 12300
tri 3746 12285 3761 12300 nw
tri 3726 12265 3746 12285 nw
tri 3903 12265 3908 12270 se
rect 3908 12265 3954 13717
tri 3954 13692 3979 13717 nw
rect 4136 13671 4182 13723
rect 4220 13763 4554 13775
rect 4220 13729 4226 13763
rect 4260 13729 4298 13763
rect 4332 13729 4370 13763
rect 4404 13729 4442 13763
rect 4476 13729 4514 13763
rect 4548 13729 4554 13763
rect 4220 13717 4554 13729
tri 4339 13692 4364 13717 ne
tri 4361 12315 4364 12318 se
rect 4364 12315 4410 13717
tri 4410 13692 4435 13717 nw
rect 4592 13691 4794 13795
tri 4410 12315 4413 12318 sw
rect 4361 12309 4413 12315
tri 3954 12265 3959 12270 sw
rect 3450 12245 3503 12265
tri 3503 12245 3523 12265 sw
tri 3883 12245 3903 12265 se
rect 3903 12245 3959 12265
tri 3959 12245 3979 12265 sw
rect 3225 12231 3269 12232
tri 2813 12179 2821 12187 se
rect 2821 12179 2887 12187
tri 2577 12178 2578 12179 sw
tri 2812 12178 2813 12179 se
rect 2813 12178 2887 12179
tri 2887 12178 2896 12187 nw
rect 2151 12176 2224 12178
tri 2224 12176 2226 12178 sw
tri 2456 12176 2458 12178 se
rect 2458 12176 2578 12178
tri 2578 12176 2580 12178 sw
tri 2810 12176 2812 12178 se
rect 2812 12176 2852 12178
rect 854 12141 1812 12153
tri 2151 12148 2179 12176 ne
rect 2179 12154 2226 12176
tri 2226 12154 2248 12176 sw
tri 2434 12154 2456 12176 se
rect 2456 12154 2580 12176
tri 2580 12154 2602 12176 sw
tri 2788 12154 2810 12176 se
rect 2810 12154 2852 12176
rect 2179 12148 2248 12154
tri 2248 12148 2254 12154 sw
rect 2417 12148 2619 12154
tri 2179 12143 2184 12148 ne
rect 2184 12143 2254 12148
tri 2184 12141 2186 12143 ne
rect 2186 12141 2254 12143
tri 2254 12141 2261 12148 sw
rect 854 12114 1780 12141
tri 1780 12114 1807 12141 nw
tri 2186 12114 2213 12141 ne
rect 2213 12114 2261 12141
tri 2261 12114 2288 12141 sw
rect 2417 12114 2429 12148
rect 2463 12114 2501 12148
rect 2535 12114 2573 12148
rect 2607 12114 2619 12148
tri 2777 12143 2788 12154 se
rect 2788 12143 2852 12154
tri 2852 12143 2887 12178 nw
rect 3224 12153 3270 12230
rect 3308 12233 3642 12245
rect 3308 12199 3314 12233
rect 3348 12199 3386 12233
rect 3420 12199 3458 12233
rect 3492 12199 3530 12233
rect 3564 12199 3602 12233
rect 3636 12199 3642 12233
rect 3308 12187 3642 12199
rect 3764 12233 4098 12245
rect 3764 12199 3770 12233
rect 3804 12199 3842 12233
rect 3876 12199 3914 12233
rect 3948 12199 3986 12233
rect 4020 12199 4058 12233
rect 4092 12199 4098 12233
rect 3764 12187 4098 12199
rect 4136 12233 4182 12285
tri 4336 12245 4361 12270 se
rect 4361 12245 4413 12257
tri 4413 12245 4439 12271 sw
rect 4638 12265 4748 13691
rect 4137 12231 4181 12232
rect 4136 12195 4182 12231
rect 4137 12194 4181 12195
tri 3270 12153 3295 12178 sw
tri 4111 12153 4136 12178 se
rect 4136 12153 4182 12193
rect 4220 12233 4361 12245
rect 4413 12233 4554 12245
rect 4220 12199 4226 12233
rect 4260 12199 4298 12233
rect 4332 12199 4361 12233
rect 4413 12199 4442 12233
rect 4476 12199 4514 12233
rect 4548 12199 4554 12233
rect 4220 12193 4361 12199
rect 4413 12193 4554 12199
rect 4862 12194 4917 16868
rect 4945 15738 4991 16929
tri 4991 15738 5016 15763 sw
rect 4945 15732 5797 15738
rect 4945 15698 5248 15732
rect 5282 15698 5320 15732
rect 5354 15698 5392 15732
rect 5426 15698 5464 15732
rect 5498 15698 5797 15732
rect 4945 15692 5797 15698
tri 5720 15667 5745 15692 ne
rect 4974 15030 5054 15664
rect 5100 15620 5643 15664
tri 5100 15595 5125 15620 nw
tri 5618 15595 5643 15620 ne
rect 5174 15580 5220 15592
rect 5174 15546 5180 15580
rect 5214 15546 5220 15580
rect 5174 15508 5220 15546
rect 5174 15474 5180 15508
rect 5214 15474 5220 15508
rect 5174 15436 5220 15474
rect 5174 15402 5180 15436
rect 5214 15402 5220 15436
rect 5174 15364 5220 15402
rect 5174 15330 5180 15364
rect 5214 15330 5220 15364
rect 5174 15292 5220 15330
rect 5174 15258 5180 15292
rect 5214 15258 5220 15292
tri 5154 15220 5174 15240 se
rect 5174 15220 5220 15258
tri 5152 15218 5154 15220 se
rect 5154 15218 5180 15220
rect 5152 15166 5158 15218
rect 5214 15186 5220 15220
rect 5210 15166 5220 15186
rect 5152 15154 5220 15166
rect 5152 15102 5158 15154
rect 5210 15148 5220 15154
rect 5214 15114 5220 15148
rect 5210 15102 5220 15114
rect 5350 15580 5396 15592
rect 5350 15546 5356 15580
rect 5390 15546 5396 15580
rect 5350 15497 5396 15546
rect 5350 15463 5356 15497
rect 5390 15463 5396 15497
rect 5350 15414 5396 15463
rect 5350 15380 5356 15414
rect 5390 15380 5396 15414
rect 5350 15331 5396 15380
rect 5350 15297 5356 15331
rect 5390 15297 5396 15331
rect 5350 15248 5396 15297
rect 5350 15214 5356 15248
rect 5390 15214 5396 15248
rect 5526 15580 5572 15592
rect 5526 15546 5532 15580
rect 5566 15546 5572 15580
rect 5526 15508 5572 15546
rect 5526 15474 5532 15508
rect 5566 15474 5572 15508
rect 5526 15436 5572 15474
rect 5526 15402 5532 15436
rect 5566 15402 5572 15436
rect 5526 15364 5572 15402
rect 5526 15330 5532 15364
rect 5566 15330 5572 15364
rect 5526 15292 5572 15330
rect 5526 15258 5532 15292
rect 5566 15258 5572 15292
tri 5503 15220 5526 15243 se
rect 5526 15220 5572 15258
rect 5350 15164 5396 15214
rect 5350 15130 5356 15164
rect 5390 15130 5396 15164
rect 5350 15066 5396 15130
tri 5501 15218 5503 15220 se
rect 5503 15218 5532 15220
rect 5501 15166 5507 15218
rect 5566 15186 5572 15220
rect 5559 15166 5572 15186
rect 5501 15154 5572 15166
rect 5501 15102 5507 15154
rect 5559 15148 5572 15154
rect 5566 15114 5572 15148
rect 5559 15102 5572 15114
rect 5351 15064 5395 15065
rect 4974 14911 5100 15030
rect 5745 15028 5797 15692
rect 5837 15273 6414 15286
rect 5837 15093 5961 15273
rect 6077 15093 6283 15273
rect 6399 15093 6414 15273
rect 5837 15080 6414 15093
tri 5797 15028 5820 15051 sw
rect 5351 15027 5395 15028
tri 5100 14911 5193 15004 sw
rect 5350 14946 5396 15026
rect 5745 15026 5820 15028
tri 5820 15026 5822 15028 sw
rect 5745 14974 6414 15026
tri 5396 14946 5424 14974 sw
rect 5350 14940 6213 14946
rect 5350 14911 6161 14940
rect 4974 14864 5193 14911
tri 5193 14864 5240 14911 sw
tri 6111 14864 6158 14911 ne
rect 6158 14888 6161 14911
rect 6158 14876 6213 14888
rect 6158 14864 6161 14876
tri 4974 14861 4977 14864 ne
rect 4977 14861 5687 14864
tri 6158 14861 6161 14864 ne
tri 4977 14821 5017 14861 ne
rect 5017 14821 5687 14861
tri 6786 14855 6825 14894 nw
tri 8024 14858 8060 14894 ne
tri 8106 14858 8142 14894 nw
tri 9341 14858 9377 14894 ne
rect 9377 14858 9380 14894
tri 9377 14855 9380 14858 ne
tri 5017 14818 5020 14821 ne
rect 5020 14818 5687 14821
tri 6158 14818 6161 14821 se
rect 6161 14818 6213 14824
tri 5020 14790 5048 14818 ne
rect 5048 14790 5103 14818
tri 5103 14793 5128 14818 nw
tri 6133 14793 6158 14818 se
rect 6158 14793 6213 14818
tri 6130 14790 6133 14793 se
rect 6133 14790 6213 14793
tri 5048 14749 5089 14790 ne
rect 5089 14749 5103 14790
tri 5089 14743 5095 14749 ne
rect 5095 14743 5103 14749
tri 5095 14735 5103 14743 ne
rect 5180 14743 6213 14790
rect 5180 14709 5192 14743
rect 5226 14732 6213 14743
rect 5226 14709 5238 14732
rect 5180 14671 5238 14709
tri 5238 14707 5263 14732 nw
tri 5295 14707 5320 14732 ne
rect 5320 14707 5378 14732
tri 5378 14707 5403 14732 nw
tri 5575 14707 5600 14732 ne
rect 5600 14707 5658 14732
tri 5658 14707 5683 14732 nw
tri 5855 14707 5880 14732 ne
rect 5880 14707 5938 14732
tri 5938 14707 5963 14732 nw
rect 5321 14705 5377 14706
rect 5601 14705 5657 14706
rect 5180 14637 5192 14671
rect 5226 14637 5238 14671
rect 5600 14669 5658 14705
rect 4220 12187 4554 12193
tri 4182 12153 4207 12178 sw
tri 5155 12153 5180 12178 se
rect 5180 12153 5238 14637
rect 5321 14668 5377 14669
rect 5601 14668 5657 14669
rect 5881 14705 5937 14706
rect 5880 14669 5938 14705
rect 5881 14668 5937 14669
rect 5320 14661 5378 14667
tri 5378 14661 5384 14667 sw
tri 5458 14661 5464 14667 se
rect 5464 14661 5522 14667
rect 5320 14642 5384 14661
tri 5384 14642 5403 14661 sw
tri 5439 14642 5458 14661 se
rect 5458 14642 5522 14661
rect 5320 14574 5522 14642
rect 5320 14555 5384 14574
tri 5384 14555 5403 14574 nw
tri 5439 14555 5458 14574 ne
rect 5458 14555 5522 14574
rect 5320 14554 5383 14555
tri 5383 14554 5384 14555 nw
tri 5458 14554 5459 14555 ne
rect 5459 14554 5522 14555
rect 5320 13876 5378 14554
tri 5378 14549 5383 14554 nw
tri 5459 14549 5464 14554 ne
rect 5320 13842 5332 13876
rect 5366 13842 5378 13876
rect 5320 13804 5378 13842
rect 5320 13770 5332 13804
rect 5366 13770 5378 13804
rect 5320 13764 5378 13770
rect 5464 13876 5522 14554
rect 5600 14661 5658 14667
tri 5658 14661 5664 14667 sw
tri 5738 14661 5744 14667 se
rect 5744 14661 5802 14667
rect 5600 14627 5612 14661
rect 5646 14642 5664 14661
tri 5664 14642 5683 14661 sw
tri 5719 14642 5738 14661 se
rect 5738 14642 5756 14661
rect 5646 14627 5756 14642
rect 5790 14627 5802 14661
rect 5600 14589 5802 14627
rect 5600 14555 5612 14589
rect 5646 14574 5756 14589
rect 5646 14555 5664 14574
tri 5664 14555 5683 14574 nw
tri 5719 14555 5738 14574 ne
rect 5738 14555 5756 14574
rect 5790 14555 5802 14589
rect 5600 14554 5663 14555
tri 5663 14554 5664 14555 nw
tri 5738 14554 5739 14555 ne
rect 5739 14554 5802 14555
rect 5600 14549 5658 14554
tri 5658 14549 5663 14554 nw
tri 5739 14549 5744 14554 ne
rect 5744 14549 5802 14554
rect 5880 14661 5938 14667
tri 5938 14661 5944 14667 sw
tri 6018 14661 6024 14667 se
rect 6024 14661 6082 14667
rect 5880 14627 5892 14661
rect 5926 14642 5944 14661
tri 5944 14642 5963 14661 sw
tri 5999 14642 6018 14661 se
rect 6018 14642 6036 14661
rect 5926 14627 6036 14642
rect 6070 14627 6082 14661
rect 5880 14589 6082 14627
rect 5880 14555 5892 14589
rect 5926 14574 6036 14589
rect 5926 14555 5944 14574
tri 5944 14555 5963 14574 nw
tri 5999 14555 6018 14574 ne
rect 6018 14555 6036 14574
rect 6070 14555 6082 14589
rect 5880 14554 5943 14555
tri 5943 14554 5944 14555 nw
tri 6018 14554 6019 14555 ne
rect 6019 14554 6082 14555
rect 5880 14549 5938 14554
tri 5938 14549 5943 14554 nw
tri 6019 14549 6024 14554 ne
rect 6024 14549 6082 14554
rect 6149 14614 6155 14666
rect 6207 14614 6218 14666
rect 6149 14602 6218 14614
rect 6149 14550 6155 14602
rect 6207 14550 6218 14602
rect 6149 14548 6218 14550
rect 5464 13842 5476 13876
rect 5510 13842 5522 13876
rect 5464 13804 5522 13842
rect 5464 13770 5476 13804
rect 5510 13770 5522 13804
rect 5464 13764 5522 13770
rect 3224 12146 5238 12153
tri 3224 12143 3227 12146 ne
rect 3227 12143 5238 12146
tri 2775 12141 2777 12143 se
rect 2777 12141 2850 12143
tri 2850 12141 2852 12143 nw
tri 3227 12141 3229 12143 ne
rect 3229 12141 5238 12143
rect 854 12108 1774 12114
tri 1774 12108 1780 12114 nw
tri 2213 12108 2219 12114 ne
rect 2219 12108 2288 12114
tri 2288 12108 2294 12114 sw
rect 2417 12108 2619 12114
tri 2742 12108 2775 12141 se
rect 2775 12108 2804 12141
rect 854 12095 1761 12108
tri 1761 12095 1774 12108 nw
tri 2219 12101 2226 12108 ne
rect 2226 12101 2294 12108
tri 2294 12101 2301 12108 sw
tri 2434 12101 2441 12108 ne
rect 2441 12101 2589 12108
tri 2226 12095 2232 12101 ne
rect 2232 12095 2301 12101
tri 2301 12095 2307 12101 sw
tri 2441 12095 2447 12101 ne
rect 2447 12095 2589 12101
tri 2589 12095 2602 12108 nw
tri 2729 12095 2742 12108 se
rect 2742 12095 2804 12108
tri 2804 12095 2850 12141 nw
tri 3229 12095 3275 12141 ne
rect 3275 12095 5238 12141
rect 854 12011 900 12095
tri 900 12070 925 12095 nw
tri 2232 12070 2257 12095 ne
rect 2257 12070 2307 12095
tri 2307 12070 2332 12095 sw
tri 2447 12070 2472 12095 ne
rect 2472 12070 2564 12095
tri 2564 12070 2589 12095 nw
tri 2704 12070 2729 12095 se
rect 2729 12070 2779 12095
tri 2779 12070 2804 12095 nw
tri 4111 12070 4136 12095 ne
tri 2257 12036 2291 12070 ne
rect 2291 12068 2332 12070
tri 2332 12068 2334 12070 sw
tri 2472 12068 2474 12070 ne
rect 2474 12068 2562 12070
tri 2562 12068 2564 12070 nw
tri 2702 12068 2704 12070 se
rect 2704 12068 2777 12070
tri 2777 12068 2779 12070 nw
rect 2291 12036 2334 12068
tri 2334 12036 2366 12068 sw
tri 2474 12047 2495 12068 ne
rect 2495 12047 2541 12068
tri 2541 12047 2562 12068 nw
tri 2681 12047 2702 12068 se
rect 2702 12047 2720 12068
tri 2670 12036 2681 12047 se
rect 2681 12036 2720 12047
tri 900 12011 925 12036 sw
tri 2291 12026 2301 12036 ne
rect 2301 12026 2366 12036
tri 2366 12026 2376 12036 sw
tri 2660 12026 2670 12036 se
rect 2670 12026 2720 12036
tri 2301 12011 2316 12026 ne
rect 2316 12011 2376 12026
tri 2376 12011 2391 12026 sw
tri 2645 12011 2660 12026 se
rect 2660 12011 2720 12026
tri 2720 12011 2777 12068 nw
tri 4111 12011 4136 12036 se
rect 4136 12011 4182 12095
tri 4182 12070 4207 12095 nw
tri 5155 12070 5180 12095 ne
rect 854 12005 2159 12011
tri 2316 12005 2322 12011 ne
rect 2322 12005 2391 12011
tri 2391 12005 2397 12011 sw
tri 2639 12005 2645 12011 se
rect 2645 12005 2714 12011
tri 2714 12005 2720 12011 nw
rect 2877 12005 4182 12011
rect 854 11971 866 12005
rect 900 11971 938 12005
rect 972 11971 1097 12005
rect 1131 11971 1169 12005
rect 1203 11971 1333 12005
rect 1367 11971 1405 12005
rect 1439 11971 1569 12005
rect 1603 11971 1641 12005
rect 1675 11971 1805 12005
rect 1839 11971 1877 12005
rect 1911 11971 2041 12005
rect 2075 11971 2113 12005
rect 2147 11971 2159 12005
tri 2322 11971 2356 12005 ne
rect 2356 11993 2397 12005
tri 2397 11993 2409 12005 sw
tri 2627 11993 2639 12005 se
rect 2639 11993 2702 12005
tri 2702 11993 2714 12005 nw
rect 2356 11971 2409 11993
tri 2409 11971 2431 11993 sw
tri 2605 11971 2627 11993 se
rect 2627 11971 2680 11993
tri 2680 11971 2702 11993 nw
rect 2877 11971 2889 12005
rect 2923 11971 2961 12005
rect 2995 11971 3125 12005
rect 3159 11971 3197 12005
rect 3231 11971 3361 12005
rect 3395 11971 3433 12005
rect 3467 11971 3597 12005
rect 3631 11971 3669 12005
rect 3703 11971 3833 12005
rect 3867 11971 3905 12005
rect 3939 11971 4064 12005
rect 4098 11971 4136 12005
rect 4170 11971 4182 12005
rect 854 11965 2159 11971
tri 2356 11965 2362 11971 ne
rect 2362 11965 2431 11971
tri 2431 11965 2437 11971 sw
tri 2599 11965 2605 11971 se
rect 2605 11965 2674 11971
tri 2674 11965 2680 11971 nw
rect 2877 11965 4182 11971
tri 984 11951 998 11965 ne
rect 998 11951 1066 11965
tri 1066 11951 1080 11965 nw
tri 1456 11951 1470 11965 ne
rect 1470 11951 1538 11965
tri 1538 11951 1552 11965 nw
tri 1928 11951 1942 11965 ne
rect 1942 11951 2010 11965
tri 2010 11951 2024 11965 nw
tri 2362 11951 2376 11965 ne
rect 2376 11952 2437 11965
tri 2437 11952 2450 11965 sw
tri 2586 11952 2599 11965 se
rect 2599 11952 2661 11965
tri 2661 11952 2674 11965 nw
tri 3012 11952 3025 11965 ne
rect 3025 11952 3095 11965
tri 3095 11952 3108 11965 nw
tri 3484 11952 3497 11965 ne
rect 3497 11952 3567 11965
tri 3567 11952 3580 11965 nw
tri 3956 11952 3969 11965 ne
rect 3969 11952 4039 11965
tri 4039 11952 4052 11965 nw
rect 2376 11951 2450 11952
tri 2450 11951 2451 11952 sw
tri 998 11940 1009 11951 ne
rect 1009 11909 1055 11951
tri 1055 11940 1066 11951 nw
tri 1470 11940 1481 11951 ne
rect 1481 11909 1527 11951
tri 1527 11940 1538 11951 nw
tri 1942 11940 1953 11951 ne
rect 1953 11909 1999 11951
tri 1999 11940 2010 11951 nw
tri 2376 11940 2387 11951 ne
rect 2387 11940 2451 11951
tri 2387 11934 2393 11940 ne
rect 557 9845 569 9879
rect 603 9845 615 9879
rect 557 9807 615 9845
rect 557 9773 569 9807
rect 603 9773 615 9807
rect 557 9767 615 9773
rect 656 9885 819 11909
tri 1242 9904 1245 9907 se
rect 1245 9904 1291 9907
tri 819 9885 838 9904 sw
tri 1223 9885 1242 9904 se
rect 1242 9885 1291 9904
tri 1291 9885 1313 9907 sw
tri 1695 9885 1717 9907 se
rect 1717 9885 1763 9907
rect 656 9879 838 9885
tri 838 9879 844 9885 sw
tri 1217 9879 1223 9885 se
rect 1223 9879 1313 9885
tri 1313 9879 1319 9885 sw
tri 1689 9879 1695 9885 se
rect 1695 9879 1763 9885
tri 1763 9879 1791 9907 sw
tri 2186 9904 2189 9907 se
rect 2189 9904 2352 11909
rect 2393 10019 2451 11940
rect 2393 9985 2405 10019
rect 2439 9985 2451 10019
rect 2393 9947 2451 9985
rect 2393 9913 2405 9947
rect 2439 9913 2451 9947
tri 2585 11951 2586 11952 se
rect 2586 11951 2660 11952
tri 2660 11951 2661 11952 nw
tri 3025 11951 3026 11952 ne
rect 3026 11951 3083 11952
rect 2585 10019 2643 11951
tri 2643 11934 2660 11951 nw
tri 3026 11940 3037 11951 ne
rect 3037 11909 3083 11951
tri 3083 11940 3095 11952 nw
tri 3497 11940 3509 11952 ne
rect 3509 11909 3555 11952
tri 3555 11940 3567 11952 nw
tri 3969 11940 3981 11952 ne
rect 3981 11909 4027 11952
tri 4027 11940 4039 11952 nw
rect 4421 11946 4479 11952
rect 2585 9985 2597 10019
rect 2631 9985 2643 10019
rect 2585 9947 2643 9985
rect 2393 9907 2451 9913
rect 2492 9908 2544 9940
rect 2585 9913 2597 9947
rect 2631 9913 2643 9947
rect 2585 9907 2643 9913
tri 2161 9879 2186 9904 se
rect 2186 9879 2352 9904
tri 2352 9879 2377 9904 sw
rect 2684 9885 2847 11909
tri 4199 9907 4217 9925 se
rect 4217 9924 4380 11909
rect 4473 11894 4479 11946
rect 4421 11882 4479 11894
rect 4473 11830 4479 11882
rect 4421 10036 4479 11830
rect 4421 10002 4433 10036
rect 4467 10002 4479 10036
rect 4421 9964 4479 10002
rect 4421 9930 4433 9964
rect 4467 9930 4479 9964
tri 4380 9924 4381 9925 sw
rect 4421 9924 4479 9930
rect 4217 9907 4381 9924
tri 4381 9907 4398 9924 sw
rect 4569 9907 4816 11981
rect 5180 10299 5238 12095
rect 5297 10516 5303 10568
rect 5355 10516 5361 10568
rect 5297 10510 5361 10516
tri 5361 10510 5419 10568 sw
rect 5297 10504 5627 10510
rect 5297 10452 5303 10504
rect 5355 10458 5627 10504
rect 5679 10458 5695 10510
rect 5747 10458 5763 10510
rect 5815 10458 5831 10510
rect 5883 10458 6078 10510
rect 5355 10452 6078 10458
rect 5297 10450 5378 10452
tri 5297 10427 5320 10450 ne
rect 5320 10427 5378 10450
tri 5378 10427 5403 10452 nw
tri 5435 10427 5460 10452 ne
rect 5460 10427 5518 10452
tri 5518 10427 5543 10452 nw
tri 5715 10427 5740 10452 ne
rect 5740 10427 5798 10452
tri 5798 10427 5823 10452 nw
tri 5995 10427 6020 10452 ne
rect 6020 10427 6078 10452
rect 5180 10265 5192 10299
rect 5226 10265 5238 10299
rect 5321 10425 5377 10426
rect 5461 10425 5517 10426
rect 5741 10425 5797 10426
rect 6021 10425 6077 10426
rect 5320 10389 5378 10425
rect 5321 10388 5377 10389
rect 5320 10381 5378 10387
rect 5320 10347 5332 10381
rect 5366 10347 5378 10381
rect 5320 10309 5378 10347
rect 5320 10275 5332 10309
rect 5366 10275 5378 10309
rect 5320 10269 5378 10275
rect 5321 10267 5377 10268
rect 5461 10388 5517 10389
rect 5741 10388 5797 10389
rect 6021 10388 6077 10389
rect 5460 10381 5518 10387
tri 5518 10381 5524 10387 sw
tri 5598 10381 5604 10387 se
rect 5604 10381 5662 10387
rect 5460 10347 5472 10381
rect 5506 10362 5524 10381
tri 5524 10362 5543 10381 sw
tri 5579 10362 5598 10381 se
rect 5598 10362 5616 10381
rect 5506 10347 5616 10362
rect 5650 10347 5662 10381
rect 5460 10309 5662 10347
rect 5460 10275 5472 10309
rect 5506 10294 5616 10309
rect 5506 10275 5524 10294
tri 5524 10275 5543 10294 nw
tri 5579 10275 5598 10294 ne
rect 5598 10275 5616 10294
rect 5650 10275 5662 10309
rect 5460 10269 5518 10275
tri 5518 10269 5524 10275 nw
tri 5598 10269 5604 10275 ne
rect 5604 10269 5662 10275
rect 5740 10381 5798 10387
tri 5798 10381 5804 10387 sw
tri 5878 10381 5884 10387 se
rect 5884 10381 5942 10387
rect 5740 10347 5752 10381
rect 5786 10362 5804 10381
tri 5804 10362 5823 10381 sw
tri 5859 10362 5878 10381 se
rect 5878 10362 5896 10381
rect 5786 10347 5896 10362
rect 5930 10347 5942 10381
rect 5740 10309 5942 10347
rect 5740 10275 5752 10309
rect 5786 10294 5896 10309
rect 5786 10275 5804 10294
tri 5804 10275 5823 10294 nw
tri 5859 10275 5878 10294 ne
rect 5878 10275 5896 10294
rect 5930 10275 5942 10309
rect 5740 10269 5798 10275
tri 5798 10269 5804 10275 nw
tri 5878 10269 5884 10275 ne
rect 5884 10269 5942 10275
rect 6020 10381 6078 10387
rect 6020 10347 6032 10381
rect 6066 10347 6078 10381
rect 6020 10309 6078 10347
rect 6020 10275 6032 10309
rect 6066 10275 6078 10309
rect 6020 10269 6078 10275
rect 6149 10335 6155 10387
rect 6207 10335 6218 10387
rect 6149 10323 6218 10335
rect 6149 10271 6155 10323
rect 6207 10271 6218 10323
rect 6149 10269 6218 10271
rect 5461 10267 5517 10268
rect 5180 10227 5238 10265
rect 5460 10231 5518 10267
rect 5321 10230 5377 10231
rect 5461 10230 5517 10231
rect 5741 10267 5797 10268
rect 5740 10231 5798 10267
rect 5741 10230 5797 10231
rect 6021 10267 6077 10268
rect 6020 10231 6078 10267
rect 6021 10230 6077 10231
rect 5180 10193 5192 10227
rect 5226 10204 5238 10227
tri 5238 10204 5263 10229 sw
tri 5295 10204 5320 10229 se
rect 5320 10204 5378 10229
tri 5378 10204 5403 10229 sw
tri 5435 10204 5460 10229 se
rect 5460 10204 5518 10229
tri 5518 10204 5543 10229 sw
tri 5715 10204 5740 10229 se
rect 5740 10204 5798 10229
tri 5798 10204 5823 10229 sw
tri 5995 10204 6020 10229 se
rect 6020 10204 6078 10229
tri 6078 10204 6103 10229 sw
rect 5226 10193 6109 10204
rect 5180 10146 6109 10193
tri 6295 10146 6298 10149 se
tri 6292 10143 6295 10146 se
rect 6295 10143 6298 10146
tri 5103 10118 5128 10143 sw
tri 6267 10118 6292 10143 se
rect 6292 10118 6298 10143
rect 5103 10117 6298 10118
rect 5051 10091 6298 10117
rect 5051 10072 6344 10091
tri 3270 9904 3273 9907 se
rect 3273 9904 3319 9907
tri 2847 9885 2866 9904 sw
tri 3251 9885 3270 9904 se
rect 3270 9885 3319 9904
rect 2684 9879 2866 9885
tri 2866 9879 2872 9885 sw
tri 3245 9879 3251 9885 se
rect 3251 9879 3319 9885
tri 3319 9879 3347 9907 sw
tri 3717 9879 3745 9907 se
rect 3745 9879 3791 9907
tri 3791 9879 3819 9907 sw
tri 4171 9879 4199 9907 se
rect 4199 9879 4398 9907
tri 4398 9879 4426 9907 sw
rect 656 9837 2377 9879
tri 2377 9837 2419 9879 sw
rect 2684 9837 6115 9879
tri 6115 9837 6157 9879 sw
rect 656 9835 2419 9837
tri 2419 9835 2421 9837 sw
tri 6099 9835 6101 9837 ne
rect 6101 9835 6157 9837
rect 656 9809 2421 9835
tri 2421 9809 2447 9835 sw
tri 6101 9809 6127 9835 ne
rect 6127 9809 6157 9835
rect 656 9797 6087 9809
tri 6087 9797 6099 9809 sw
tri 6127 9797 6139 9809 ne
rect 6139 9797 6157 9809
rect 656 9779 6099 9797
tri 6099 9779 6117 9797 sw
tri 6139 9779 6157 9797 ne
tri 6157 9779 6215 9837 sw
rect 656 9767 6117 9779
tri 6117 9767 6129 9779 sw
tri 6157 9767 6169 9779 ne
rect 6169 9767 6215 9779
tri 6071 9764 6074 9767 ne
rect 6074 9764 6129 9767
tri 6129 9764 6132 9767 sw
tri 6169 9764 6172 9767 ne
rect 6172 9764 6215 9767
tri 513 9739 538 9764 sw
tri 6074 9754 6084 9764 ne
rect 6084 9754 6132 9764
tri 6132 9754 6142 9764 sw
tri 6172 9754 6182 9764 ne
rect 6182 9754 6215 9764
tri 6084 9751 6087 9754 ne
rect 6087 9751 6142 9754
tri 6087 9739 6099 9751 ne
rect 6099 9739 6142 9751
tri 6142 9739 6157 9754 sw
tri 6182 9739 6197 9754 ne
rect 6197 9739 6215 9754
rect 122 9693 683 9739
rect 122 447 360 9693
rect 392 9687 536 9693
tri 536 9687 542 9693 nw
tri 2285 9687 2291 9693 ne
rect 2291 9687 2297 9739
rect 2349 9687 2361 9739
rect 2413 9687 2425 9739
rect 2477 9687 2489 9739
rect 2541 9687 2553 9739
rect 2605 9687 2617 9739
rect 2669 9687 2681 9739
rect 2733 9687 2739 9739
rect 4353 9693 4781 9739
tri 2739 9687 2745 9693 nw
tri 4769 9687 4775 9693 ne
rect 4775 9687 4781 9693
rect 4833 9687 4845 9739
rect 4897 9687 4903 9739
rect 6013 9693 6059 9739
tri 6099 9696 6142 9739 ne
rect 6142 9721 6157 9739
tri 6157 9721 6175 9739 sw
tri 6197 9721 6215 9739 ne
tri 6215 9721 6273 9779 sw
rect 6142 9696 6175 9721
tri 6175 9696 6200 9721 sw
tri 6215 9696 6240 9721 ne
rect 6240 9696 6273 9721
tri 4903 9687 4909 9693 nw
tri 5988 9687 5994 9693 ne
rect 5994 9687 6059 9693
rect 392 9668 517 9687
tri 517 9668 536 9687 nw
tri 5994 9668 6013 9687 ne
rect 392 9661 510 9668
tri 510 9661 517 9668 nw
rect 6013 9661 6059 9687
tri 6142 9661 6177 9696 ne
rect 6177 9681 6200 9696
tri 6200 9681 6215 9696 sw
tri 6240 9681 6255 9696 ne
rect 6255 9684 6273 9696
tri 6273 9684 6310 9721 sw
rect 6255 9681 6365 9684
rect 6177 9663 6215 9681
tri 6215 9663 6233 9681 sw
tri 6255 9663 6273 9681 ne
rect 6273 9663 6365 9681
rect 6177 9661 6233 9663
tri 6233 9661 6235 9663 sw
tri 6273 9661 6275 9663 ne
rect 6275 9661 6365 9663
rect 392 9653 502 9661
tri 502 9653 510 9661 nw
tri 6177 9653 6185 9661 ne
rect 6185 9653 6235 9661
tri 6235 9653 6243 9661 sw
tri 6275 9653 6283 9661 ne
rect 6283 9653 6365 9661
rect 392 9638 487 9653
tri 487 9638 502 9653 nw
rect 542 9638 5525 9653
tri 6185 9638 6200 9653 ne
rect 6200 9638 6243 9653
tri 6243 9638 6258 9653 sw
tri 6283 9638 6298 9653 ne
rect 6298 9638 6365 9653
rect 392 9604 453 9638
tri 453 9604 487 9638 nw
rect 542 9604 548 9638
rect 582 9604 620 9638
rect 654 9604 2354 9638
rect 2388 9604 2426 9638
rect 2460 9604 2576 9638
rect 2610 9604 2648 9638
rect 2682 9604 4382 9638
rect 4416 9604 4454 9638
rect 4488 9604 5525 9638
rect 392 9589 438 9604
tri 438 9589 453 9604 nw
rect 542 9589 5525 9604
rect 392 9564 413 9589
tri 413 9564 438 9589 nw
tri 1054 9564 1079 9589 ne
rect 392 9550 399 9564
tri 399 9550 413 9564 nw
rect 392 9544 393 9550
tri 393 9544 399 9550 nw
rect 534 9544 1024 9550
tri 392 9543 393 9544 nw
rect 534 9510 546 9544
rect 580 9510 618 9544
rect 652 9510 690 9544
rect 724 9510 762 9544
rect 796 9510 834 9544
rect 868 9510 906 9544
rect 940 9510 978 9544
rect 1012 9510 1024 9544
rect 534 9504 1024 9510
rect 1079 9547 1125 9589
tri 1125 9564 1150 9589 nw
tri 1910 9564 1935 9589 ne
rect 1080 9545 1124 9546
rect 1079 9509 1125 9545
rect 1080 9508 1124 9509
rect 534 9363 700 9504
tri 700 9479 725 9504 nw
tri 1068 9479 1079 9490 se
rect 1079 9479 1125 9507
rect 1935 9547 1981 9589
tri 1981 9564 2006 9589 nw
tri 2766 9564 2791 9589 ne
rect 1936 9545 1980 9546
rect 1935 9509 1981 9545
rect 1936 9508 1980 9509
tri 1422 9490 1436 9504 ne
rect 1436 9490 1613 9504
tri 1125 9479 1136 9490 sw
tri 1436 9479 1447 9490 ne
tri 1054 9465 1068 9479 se
rect 1068 9465 1136 9479
tri 1136 9465 1150 9479 sw
rect 1079 9455 1125 9465
tri 1054 9394 1079 9419 ne
rect 534 7293 697 9363
tri 697 9360 700 9363 nw
tri 1063 7318 1079 7334 se
rect 1079 7328 1125 9419
tri 1125 9394 1150 9419 nw
tri 1125 7328 1131 7334 sw
rect 1079 7318 1131 7328
tri 1131 7318 1141 7328 sw
tri 697 7293 722 7318 sw
tri 1038 7293 1063 7318 se
rect 1063 7293 1141 7318
tri 1141 7293 1166 7318 sw
tri 1422 7293 1447 7318 se
rect 1447 7293 1613 9490
tri 1613 9479 1638 9504 nw
tri 1924 9479 1935 9490 se
rect 1935 9479 1981 9507
rect 2791 9547 2837 9589
tri 2837 9564 2862 9589 nw
tri 3886 9564 3911 9589 ne
rect 2792 9545 2836 9546
rect 2791 9509 2837 9545
rect 2792 9508 2836 9509
tri 2278 9490 2292 9504 ne
rect 2292 9490 2469 9504
tri 1981 9479 1992 9490 sw
tri 2292 9479 2303 9490 ne
tri 1910 9465 1924 9479 se
rect 1924 9465 1992 9479
tri 1992 9465 2006 9479 sw
rect 1935 9455 1981 9465
tri 1910 9394 1935 9419 ne
tri 1929 7328 1935 7334 se
rect 1935 7328 1981 9419
tri 1981 9394 2006 9419 nw
tri 1981 7328 1987 7334 sw
tri 1919 7318 1929 7328 se
rect 1929 7318 1987 7328
tri 1987 7318 1997 7328 sw
tri 1613 7293 1638 7318 sw
tri 1894 7293 1919 7318 se
rect 1919 7293 1997 7318
tri 1997 7293 2022 7318 sw
tri 2278 7293 2303 7318 se
rect 2303 7293 2469 9490
tri 2469 9479 2494 9504 nw
tri 2780 9479 2791 9490 se
rect 2791 9479 2837 9507
rect 3268 9504 3480 9550
tri 3268 9490 3282 9504 ne
rect 3282 9490 3455 9504
tri 2837 9479 2848 9490 sw
tri 3282 9479 3293 9490 ne
tri 2766 9465 2780 9479 se
rect 2780 9465 2848 9479
tri 2848 9465 2862 9479 sw
rect 2791 9455 2837 9465
tri 2766 9394 2791 9419 ne
tri 2785 7328 2791 7334 se
rect 2791 7328 2837 9419
tri 2837 9394 2862 9419 nw
tri 3268 9363 3293 9388 se
rect 3293 9363 3455 9490
tri 3455 9479 3480 9504 nw
rect 3911 9547 3957 9589
tri 3957 9564 3982 9589 nw
tri 4542 9564 4567 9589 ne
rect 3912 9545 3956 9546
rect 3911 9509 3957 9545
rect 3912 9508 3956 9509
tri 3900 9479 3911 9490 se
rect 3911 9479 3957 9507
rect 4024 9544 4514 9550
rect 4024 9510 4036 9544
rect 4070 9510 4108 9544
rect 4142 9510 4180 9544
rect 4214 9510 4252 9544
rect 4286 9510 4324 9544
rect 4358 9510 4396 9544
rect 4430 9510 4468 9544
rect 4502 9510 4514 9544
rect 4024 9504 4514 9510
rect 4567 9547 4613 9589
tri 4613 9564 4638 9589 nw
tri 4998 9564 5023 9589 ne
rect 4568 9545 4612 9546
rect 4567 9509 4613 9545
rect 4568 9508 4612 9509
tri 4254 9490 4268 9504 ne
rect 4268 9490 4456 9504
tri 4456 9490 4470 9504 nw
tri 3886 9465 3900 9479 se
rect 3900 9465 3957 9479
tri 3957 9465 3982 9490 sw
tri 4268 9479 4279 9490 ne
rect 3911 9455 3957 9465
tri 3886 9394 3911 9419 ne
tri 3455 9363 3480 9388 sw
tri 2837 7328 2843 7334 sw
tri 2775 7318 2785 7328 se
rect 2785 7318 2843 7328
tri 2843 7318 2853 7328 sw
tri 2469 7293 2494 7318 sw
tri 2750 7293 2775 7318 se
rect 2775 7293 2853 7318
tri 2853 7293 2878 7318 sw
tri 3194 7293 3219 7318 se
rect 3219 7293 3529 9363
tri 3905 7328 3911 7334 se
rect 3911 7328 3957 9419
tri 3957 9394 3982 9419 nw
tri 3957 7328 3963 7334 sw
tri 3895 7318 3905 7328 se
rect 3905 7318 3963 7328
tri 3963 7318 3973 7328 sw
tri 3529 7293 3554 7318 sw
tri 3870 7293 3895 7318 se
rect 3895 7293 3973 7318
tri 3973 7293 3998 7318 sw
tri 4254 7293 4279 7318 se
rect 4279 7293 4445 9490
tri 4445 9479 4456 9490 nw
tri 4556 9479 4567 9490 se
rect 4567 9479 4613 9507
rect 4646 9544 4992 9550
rect 4646 9510 4658 9544
rect 4692 9510 4730 9544
rect 4764 9510 4802 9544
rect 4836 9510 4874 9544
rect 4908 9510 4946 9544
rect 4980 9510 4992 9544
rect 4646 9504 4992 9510
rect 5023 9547 5069 9589
tri 5069 9564 5094 9589 nw
tri 5454 9564 5479 9589 ne
rect 5024 9545 5068 9546
rect 5023 9509 5069 9545
rect 5024 9508 5068 9509
tri 4710 9490 4724 9504 ne
rect 4724 9490 4912 9504
tri 4912 9490 4926 9504 nw
tri 4542 9465 4556 9479 se
rect 4556 9465 4613 9479
tri 4613 9465 4638 9490 sw
tri 4724 9479 4735 9490 ne
rect 4489 9459 4691 9465
rect 4489 9425 4501 9459
rect 4535 9425 4573 9459
rect 4607 9425 4645 9459
rect 4679 9425 4691 9459
rect 4489 9419 4691 9425
tri 4542 9394 4567 9419 ne
tri 4561 7328 4567 7334 se
rect 4567 7328 4613 9419
tri 4613 9394 4638 9419 nw
tri 4613 7328 4619 7334 sw
tri 4551 7318 4561 7328 se
rect 4561 7318 4619 7328
tri 4550 7317 4551 7318 se
rect 4551 7317 4619 7318
tri 4619 7317 4630 7328 sw
tri 4526 7293 4550 7317 se
rect 4550 7293 4630 7317
tri 4630 7293 4654 7317 sw
rect 534 7287 919 7293
rect 534 7253 657 7287
rect 691 7253 729 7287
rect 763 7253 801 7287
rect 835 7253 873 7287
rect 907 7253 919 7287
rect 534 7247 919 7253
tri 1037 7292 1038 7293 se
rect 1038 7292 1166 7293
tri 1166 7292 1167 7293 sw
rect 1037 7286 1167 7292
rect 1037 7252 1049 7286
rect 1083 7252 1121 7286
rect 1155 7252 1167 7286
rect 534 5073 697 7247
tri 697 7222 722 7247 nw
rect 1037 7246 1167 7252
rect 1285 7287 1775 7293
rect 1285 7253 1297 7287
rect 1331 7253 1369 7287
rect 1403 7253 1441 7287
rect 1475 7253 1513 7287
rect 1547 7253 1585 7287
rect 1619 7253 1657 7287
rect 1691 7253 1729 7287
rect 1763 7253 1775 7287
rect 1285 7247 1775 7253
tri 1893 7292 1894 7293 se
rect 1894 7292 2022 7293
tri 2022 7292 2023 7293 sw
rect 1893 7286 2023 7292
rect 1893 7252 1905 7286
rect 1939 7252 1977 7286
rect 2011 7252 2023 7286
tri 1037 7222 1061 7246 ne
rect 1061 7222 1125 7246
tri 1061 7204 1079 7222 ne
tri 1063 5098 1079 5114 se
rect 1079 5098 1125 7222
tri 1125 7204 1167 7246 nw
tri 1422 7222 1447 7247 ne
tri 697 5073 722 5098 sw
tri 1038 5073 1063 5098 se
rect 1063 5073 1125 5098
tri 1125 5073 1166 5114 sw
tri 1422 5073 1447 5098 se
rect 1447 5073 1613 7247
tri 1613 7222 1638 7247 nw
rect 1893 7246 2023 7252
rect 2141 7287 2631 7293
rect 2141 7253 2153 7287
rect 2187 7253 2225 7287
rect 2259 7253 2297 7287
rect 2331 7253 2369 7287
rect 2403 7253 2441 7287
rect 2475 7253 2513 7287
rect 2547 7253 2585 7287
rect 2619 7253 2631 7287
rect 2141 7247 2631 7253
tri 2749 7292 2750 7293 se
rect 2750 7292 2878 7293
tri 2878 7292 2879 7293 sw
rect 2749 7286 2879 7292
rect 2749 7252 2761 7286
rect 2795 7252 2833 7286
rect 2867 7252 2879 7286
tri 2278 7246 2279 7247 ne
rect 2279 7246 2469 7247
tri 1893 7222 1917 7246 ne
rect 1917 7222 1999 7246
tri 1999 7222 2023 7246 nw
tri 2279 7222 2303 7246 ne
tri 1917 7204 1935 7222 ne
tri 1919 5098 1935 5114 se
rect 1935 5098 1981 7222
tri 1981 7204 1999 7222 nw
tri 1613 5073 1638 5098 sw
tri 1894 5073 1919 5098 se
rect 1919 5073 1981 5098
tri 1981 5073 2022 5114 sw
tri 2278 5073 2303 5098 se
rect 2303 5073 2469 7246
tri 2469 7222 2494 7247 nw
rect 2749 7246 2879 7252
rect 2997 7287 3751 7293
rect 2997 7253 3009 7287
rect 3043 7253 3081 7287
rect 3115 7253 3153 7287
rect 3187 7253 3225 7287
rect 3259 7253 3489 7287
rect 3523 7253 3561 7287
rect 3595 7253 3633 7287
rect 3667 7253 3705 7287
rect 3739 7253 3751 7287
rect 2997 7247 3751 7253
tri 3869 7292 3870 7293 se
rect 3870 7292 3998 7293
tri 3998 7292 3999 7293 sw
rect 3869 7286 3999 7292
rect 3869 7252 3881 7286
rect 3915 7252 3953 7286
rect 3987 7252 3999 7286
tri 2749 7222 2773 7246 ne
rect 2773 7222 2837 7246
tri 2773 7204 2791 7222 ne
tri 2775 5098 2791 5114 se
rect 2791 5098 2837 7222
tri 2837 7204 2879 7246 nw
tri 3194 7222 3219 7247 ne
tri 2469 5073 2494 5098 sw
tri 2750 5073 2775 5098 se
rect 2775 5073 2837 5098
tri 2837 5073 2878 5114 sw
tri 3194 5073 3219 5098 se
rect 3219 5073 3529 7247
tri 3529 7222 3554 7247 nw
rect 3869 7246 3999 7252
rect 4117 7287 4445 7293
rect 4117 7253 4129 7287
rect 4163 7253 4201 7287
rect 4235 7253 4273 7287
rect 4307 7253 4345 7287
rect 4379 7253 4445 7287
rect 4117 7247 4445 7253
tri 4254 7246 4255 7247 ne
rect 4255 7246 4445 7247
tri 3869 7222 3893 7246 ne
rect 3893 7222 3975 7246
tri 3975 7222 3999 7246 nw
tri 4255 7222 4279 7246 ne
tri 3893 7204 3911 7222 ne
tri 3895 5098 3911 5114 se
rect 3911 5098 3957 7222
tri 3957 7204 3975 7222 nw
tri 3957 5098 3973 5114 sw
tri 3529 5073 3554 5098 sw
tri 3870 5073 3895 5098 se
rect 3895 5073 3973 5098
tri 3973 5073 3998 5098 sw
tri 4254 5073 4279 5098 se
rect 4279 5073 4445 7246
tri 4525 7292 4526 7293 se
rect 4526 7292 4654 7293
tri 4654 7292 4655 7293 sw
rect 4525 7286 4655 7292
rect 4525 7252 4537 7286
rect 4571 7252 4609 7286
rect 4643 7252 4655 7286
rect 4525 7246 4655 7252
tri 4525 7222 4549 7246 ne
rect 4549 7222 4631 7246
tri 4631 7222 4655 7246 nw
rect 4735 7287 4901 9490
tri 4901 9479 4912 9490 nw
tri 5012 9479 5023 9490 se
rect 5023 9479 5069 9507
rect 5101 9544 5303 9550
rect 5355 9544 5447 9550
rect 5101 9510 5113 9544
rect 5147 9510 5185 9544
rect 5219 9510 5257 9544
rect 5291 9510 5303 9544
rect 5363 9510 5401 9544
rect 5435 9510 5447 9544
rect 5101 9504 5303 9510
tri 5166 9490 5180 9504 ne
rect 5180 9498 5303 9504
rect 5355 9504 5447 9510
rect 5479 9547 5525 9589
tri 6200 9580 6258 9638 ne
tri 6258 9623 6273 9638 sw
tri 6298 9623 6313 9638 ne
rect 6313 9623 6365 9638
rect 6258 9620 6273 9623
tri 6273 9620 6276 9623 sw
tri 6313 9620 6316 9623 ne
rect 6316 9620 6365 9623
rect 6258 9580 6276 9620
tri 6276 9580 6316 9620 sw
tri 6258 9550 6288 9580 ne
rect 6288 9550 6365 9580
rect 5480 9545 5524 9546
rect 5479 9509 5525 9545
rect 5480 9508 5524 9509
rect 5355 9498 5361 9504
rect 5180 9490 5361 9498
tri 5069 9479 5080 9490 sw
tri 5180 9479 5191 9490 ne
rect 5191 9486 5361 9490
tri 4998 9465 5012 9479 se
rect 5012 9465 5080 9479
tri 5080 9465 5094 9479 sw
rect 4945 9459 5147 9465
rect 4945 9425 4957 9459
rect 4991 9425 5029 9459
rect 5063 9425 5101 9459
rect 5135 9425 5147 9459
rect 4945 9419 5147 9425
rect 5191 9434 5303 9486
rect 5355 9434 5361 9486
tri 5361 9477 5388 9504 nw
tri 5466 9477 5479 9490 se
rect 5479 9477 5525 9507
rect 5596 9544 5870 9550
rect 5596 9510 5608 9544
rect 5642 9510 5680 9544
rect 5714 9510 5752 9544
rect 5786 9510 5824 9544
rect 5858 9510 5870 9544
tri 6288 9516 6322 9550 ne
rect 6322 9516 6365 9550
rect 5596 9504 5870 9510
tri 5622 9490 5636 9504 ne
rect 5636 9490 5870 9504
tri 5454 9465 5466 9477 se
rect 5466 9465 5525 9477
tri 5525 9465 5550 9490 sw
tri 5636 9479 5647 9490 ne
tri 4998 9394 5023 9419 ne
tri 5017 7328 5023 7334 se
rect 5023 7328 5069 9419
tri 5069 9394 5094 9419 nw
tri 5007 7318 5017 7328 se
rect 5017 7318 5069 7328
tri 5006 7317 5007 7318 se
rect 5007 7317 5069 7318
tri 5069 7317 5086 7334 sw
tri 4982 7293 5006 7317 se
rect 5006 7293 5086 7317
tri 5086 7293 5110 7317 sw
rect 4735 7253 4765 7287
rect 4799 7253 4837 7287
rect 4871 7253 4901 7287
tri 4549 7204 4567 7222 ne
rect 534 5067 919 5073
rect 534 5033 657 5067
rect 691 5033 729 5067
rect 763 5033 801 5067
rect 835 5033 873 5067
rect 907 5033 919 5067
rect 534 5027 919 5033
tri 1037 5072 1038 5073 se
rect 1038 5072 1166 5073
tri 1166 5072 1167 5073 sw
rect 1037 5066 1167 5072
rect 1037 5032 1049 5066
rect 1083 5032 1121 5066
rect 1155 5032 1167 5066
rect 534 2854 697 5027
tri 697 5002 722 5027 nw
rect 1037 5026 1167 5032
rect 1285 5067 1775 5073
rect 1285 5033 1297 5067
rect 1331 5033 1369 5067
rect 1403 5033 1441 5067
rect 1475 5033 1513 5067
rect 1547 5033 1585 5067
rect 1619 5033 1657 5067
rect 1691 5033 1729 5067
rect 1763 5033 1775 5067
rect 1285 5027 1775 5033
tri 1893 5072 1894 5073 se
rect 1894 5072 2022 5073
tri 2022 5072 2023 5073 sw
rect 1893 5066 2023 5072
rect 1893 5032 1905 5066
rect 1939 5032 1977 5066
rect 2011 5032 2023 5066
tri 1037 5002 1061 5026 ne
rect 1061 5002 1125 5026
tri 1061 4984 1079 5002 ne
tri 1063 2879 1079 2895 se
rect 1079 2879 1125 5002
tri 1125 4984 1167 5026 nw
tri 1422 5002 1447 5027 ne
tri 697 2854 722 2879 sw
tri 1038 2854 1063 2879 se
rect 1063 2854 1125 2879
tri 1125 2854 1166 2895 sw
tri 1422 2854 1447 2879 se
rect 1447 2854 1613 5027
tri 1613 5002 1638 5027 nw
rect 1893 5026 2023 5032
rect 2141 5067 2631 5073
rect 2141 5033 2153 5067
rect 2187 5033 2225 5067
rect 2259 5033 2297 5067
rect 2331 5033 2369 5067
rect 2403 5033 2441 5067
rect 2475 5033 2513 5067
rect 2547 5033 2585 5067
rect 2619 5033 2631 5067
rect 2141 5027 2631 5033
tri 2749 5072 2750 5073 se
rect 2750 5072 2878 5073
tri 2878 5072 2879 5073 sw
rect 2749 5066 2879 5072
rect 2749 5032 2761 5066
rect 2795 5032 2833 5066
rect 2867 5032 2879 5066
tri 1893 5002 1917 5026 ne
rect 1917 5002 1981 5026
tri 1917 4984 1935 5002 ne
tri 1919 2879 1935 2895 se
rect 1935 2879 1981 5002
tri 1981 4984 2023 5026 nw
tri 2278 5002 2303 5027 ne
tri 1613 2854 1638 2879 sw
tri 1894 2854 1919 2879 se
rect 1919 2854 1981 2879
tri 1981 2854 2022 2895 sw
tri 2278 2854 2303 2879 se
rect 2303 2854 2469 5027
tri 2469 5002 2494 5027 nw
rect 2749 5026 2879 5032
rect 2997 5067 3751 5073
rect 2997 5033 3009 5067
rect 3043 5033 3081 5067
rect 3115 5033 3153 5067
rect 3187 5033 3225 5067
rect 3259 5033 3489 5067
rect 3523 5033 3561 5067
rect 3595 5033 3633 5067
rect 3667 5033 3705 5067
rect 3739 5033 3751 5067
rect 2997 5027 3751 5033
tri 3869 5072 3870 5073 se
rect 3870 5072 3998 5073
tri 3998 5072 3999 5073 sw
rect 3869 5066 3999 5072
rect 3869 5032 3881 5066
rect 3915 5032 3953 5066
rect 3987 5032 3999 5066
tri 2749 5002 2773 5026 ne
rect 2773 5002 2837 5026
tri 2773 4984 2791 5002 ne
tri 2775 2879 2791 2895 se
rect 2791 2879 2837 5002
tri 2837 4984 2879 5026 nw
tri 3194 5002 3219 5027 ne
rect 3219 5026 3553 5027
tri 3553 5026 3554 5027 nw
rect 3869 5026 3999 5032
rect 4117 5067 4445 5073
rect 4117 5033 4129 5067
rect 4163 5033 4201 5067
rect 4235 5033 4273 5067
rect 4307 5033 4345 5067
rect 4379 5033 4445 5067
rect 4117 5027 4445 5033
tri 4254 5026 4255 5027 ne
rect 4255 5026 4445 5027
tri 2469 2854 2494 2879 sw
tri 2750 2854 2775 2879 se
rect 2775 2854 2837 2879
tri 2837 2854 2878 2895 sw
tri 3194 2854 3219 2879 se
rect 3219 2855 3529 5026
tri 3529 5002 3553 5026 nw
tri 3869 5002 3893 5026 ne
rect 3893 5002 3975 5026
tri 3975 5002 3999 5026 nw
tri 4255 5002 4279 5026 ne
tri 3893 4984 3911 5002 ne
tri 3895 2879 3911 2895 se
rect 3911 2879 3957 5002
tri 3957 4984 3975 5002 nw
tri 3957 2879 3973 2895 sw
tri 3529 2855 3553 2879 sw
tri 3871 2855 3895 2879 se
rect 3895 2855 3973 2879
tri 3973 2855 3997 2879 sw
tri 4255 2855 4279 2879 se
rect 4279 2855 4445 5026
tri 4525 5072 4567 5114 se
rect 4567 5072 4613 7222
tri 4613 7204 4631 7222 nw
tri 4613 5072 4655 5114 sw
rect 4525 5066 4655 5072
rect 4525 5032 4537 5066
rect 4571 5032 4609 5066
rect 4643 5032 4655 5066
rect 4525 5026 4655 5032
tri 4525 4984 4567 5026 ne
rect 3219 2854 3553 2855
tri 3553 2854 3554 2855 sw
tri 3870 2854 3871 2855 se
rect 3871 2854 3997 2855
tri 3997 2854 3998 2855 sw
tri 4254 2854 4255 2855 se
rect 4255 2854 4445 2855
rect 534 2848 919 2854
rect 534 2814 657 2848
rect 691 2814 729 2848
rect 763 2814 801 2848
rect 835 2814 873 2848
rect 907 2814 919 2848
rect 534 2808 919 2814
tri 1037 2853 1038 2854 se
rect 1038 2853 1166 2854
tri 1166 2853 1167 2854 sw
rect 1037 2847 1167 2853
rect 1037 2813 1049 2847
rect 1083 2813 1121 2847
rect 1155 2813 1167 2847
rect 534 597 697 2808
tri 697 2783 722 2808 nw
rect 1037 2807 1167 2813
rect 1285 2848 1775 2854
rect 1285 2814 1297 2848
rect 1331 2814 1369 2848
rect 1403 2814 1441 2848
rect 1475 2814 1513 2848
rect 1547 2814 1585 2848
rect 1619 2814 1657 2848
rect 1691 2814 1729 2848
rect 1763 2814 1775 2848
rect 1285 2808 1775 2814
tri 1893 2853 1894 2854 se
rect 1894 2853 2022 2854
tri 2022 2853 2023 2854 sw
rect 1893 2847 2023 2853
rect 1893 2813 1905 2847
rect 1939 2813 1977 2847
rect 2011 2813 2023 2847
tri 1037 2783 1061 2807 ne
rect 1061 2783 1125 2807
tri 1061 2765 1079 2783 ne
tri 1054 682 1079 707 se
rect 1079 682 1125 2783
tri 1125 2765 1167 2807 nw
tri 1422 2783 1447 2808 ne
tri 1125 682 1150 707 sw
tri 697 597 722 622 sw
tri 1422 597 1447 622 se
rect 1447 597 1613 2808
tri 1613 2783 1638 2808 nw
rect 1893 2807 2023 2813
rect 2141 2848 2631 2854
rect 2141 2814 2153 2848
rect 2187 2814 2225 2848
rect 2259 2814 2297 2848
rect 2331 2814 2369 2848
rect 2403 2814 2441 2848
rect 2475 2814 2513 2848
rect 2547 2814 2585 2848
rect 2619 2814 2631 2848
rect 2141 2808 2631 2814
tri 2749 2853 2750 2854 se
rect 2750 2853 2878 2854
tri 2878 2853 2879 2854 sw
rect 2749 2847 2879 2853
rect 2749 2813 2761 2847
rect 2795 2813 2833 2847
rect 2867 2813 2879 2847
tri 1893 2783 1917 2807 ne
rect 1917 2783 1981 2807
tri 1917 2765 1935 2783 ne
tri 1910 682 1935 707 se
rect 1935 682 1981 2783
tri 1981 2765 2023 2807 nw
tri 2278 2783 2303 2808 ne
tri 1981 682 2006 707 sw
tri 1613 597 1638 622 sw
tri 2278 597 2303 622 se
rect 2303 597 2469 2808
tri 2469 2783 2494 2808 nw
rect 2749 2807 2879 2813
rect 2997 2848 3751 2854
rect 2997 2814 3009 2848
rect 3043 2814 3081 2848
rect 3115 2814 3153 2848
rect 3187 2814 3225 2848
rect 3259 2814 3489 2848
rect 3523 2814 3561 2848
rect 3595 2814 3633 2848
rect 3667 2814 3705 2848
rect 3739 2814 3751 2848
rect 2997 2808 3751 2814
tri 3869 2853 3870 2854 se
rect 3870 2853 3998 2854
tri 3998 2853 3999 2854 sw
rect 3869 2847 3999 2853
rect 3869 2813 3881 2847
rect 3915 2813 3953 2847
rect 3987 2813 3999 2847
tri 2749 2783 2773 2807 ne
rect 2773 2783 2837 2807
tri 2773 2765 2791 2783 ne
tri 2766 682 2791 707 se
rect 2791 682 2837 2783
tri 2837 2765 2879 2807 nw
tri 3194 2783 3219 2808 ne
rect 3219 2807 3553 2808
tri 3553 2807 3554 2808 nw
rect 3869 2807 3999 2813
rect 4117 2848 4445 2854
rect 4117 2814 4129 2848
rect 4163 2814 4201 2848
rect 4235 2814 4273 2848
rect 4307 2814 4345 2848
rect 4379 2814 4445 2848
rect 4117 2808 4445 2814
tri 4254 2807 4255 2808 ne
rect 4255 2807 4445 2808
tri 2837 682 2862 707 sw
tri 2469 597 2494 622 sw
tri 3194 597 3219 622 se
rect 3219 597 3529 2807
tri 3529 2783 3553 2807 nw
tri 3869 2783 3893 2807 ne
rect 3893 2783 3975 2807
tri 3975 2783 3999 2807 nw
tri 4255 2783 4279 2807 ne
tri 3893 2765 3911 2783 ne
tri 3886 682 3911 707 se
rect 3911 682 3957 2783
tri 3957 2765 3975 2783 nw
tri 3957 682 3982 707 sw
tri 3529 597 3554 622 sw
tri 4254 597 4279 622 se
rect 4279 597 4445 2807
tri 4525 2853 4567 2895 se
rect 4567 2853 4613 5026
tri 4613 4984 4655 5026 nw
rect 4735 5067 4901 7253
tri 4981 7292 4982 7293 se
rect 4982 7292 5110 7293
tri 5110 7292 5111 7293 sw
rect 4981 7286 5111 7292
rect 4981 7252 4993 7286
rect 5027 7252 5065 7286
rect 5099 7252 5111 7286
rect 4981 7246 5111 7252
tri 4981 7222 5005 7246 ne
rect 5005 7222 5069 7246
tri 5005 7204 5023 7222 ne
rect 4735 5033 4765 5067
rect 4799 5033 4837 5067
rect 4871 5033 4901 5067
tri 4613 2853 4655 2895 sw
rect 4525 2847 4655 2853
rect 4525 2813 4537 2847
rect 4571 2813 4609 2847
rect 4643 2813 4655 2847
rect 4525 2807 4655 2813
tri 4525 2765 4567 2807 ne
tri 4542 682 4567 707 se
rect 4567 682 4613 2807
tri 4613 2765 4655 2807 nw
rect 4735 2848 4901 5033
tri 4981 5072 5023 5114 se
rect 5023 5072 5069 7222
tri 5069 7204 5111 7246 nw
rect 5191 7287 5357 9434
tri 5357 9430 5361 9434 nw
rect 5401 9459 5603 9465
rect 5401 9425 5413 9459
rect 5447 9425 5485 9459
rect 5519 9425 5557 9459
rect 5591 9425 5603 9459
rect 5401 9419 5603 9425
tri 5454 9394 5479 9419 ne
tri 5457 7312 5479 7334 se
rect 5479 7312 5525 9419
tri 5525 9394 5550 9419 nw
tri 5525 7312 5547 7334 sw
rect 5191 7253 5221 7287
rect 5255 7253 5293 7287
rect 5327 7253 5357 7287
tri 5069 5072 5111 5114 sw
rect 4981 5066 5111 5072
rect 4981 5032 4993 5066
rect 5027 5032 5065 5066
rect 5099 5032 5111 5066
rect 4981 5026 5111 5032
tri 4981 4984 5023 5026 ne
rect 4735 2814 4765 2848
rect 4799 2814 4837 2848
rect 4871 2814 4901 2848
tri 4613 682 4638 707 sw
rect 4489 676 4691 682
rect 4489 642 4501 676
rect 4535 642 4573 676
rect 4607 642 4645 676
rect 4679 642 4691 676
rect 4489 636 4691 642
tri 4445 597 4470 622 sw
tri 4710 597 4735 622 se
rect 4735 597 4901 2814
tri 4981 2853 5023 2895 se
rect 5023 2853 5069 5026
tri 5069 4984 5111 5026 nw
rect 5191 5067 5357 7253
tri 5437 7292 5457 7312 se
rect 5457 7293 5547 7312
tri 5547 7293 5566 7312 sw
rect 5457 7292 5566 7293
tri 5566 7292 5567 7293 sw
rect 5437 7286 5567 7292
rect 5437 7252 5449 7286
rect 5483 7252 5521 7286
rect 5555 7252 5567 7286
rect 5437 7246 5567 7252
tri 5437 7204 5479 7246 ne
rect 5191 5033 5221 5067
rect 5255 5033 5293 5067
rect 5327 5033 5357 5067
tri 5069 2853 5111 2895 sw
rect 4981 2847 5111 2853
rect 4981 2813 4993 2847
rect 5027 2813 5065 2847
rect 5099 2813 5111 2847
rect 4981 2807 5111 2813
tri 4981 2765 5023 2807 ne
tri 4998 682 5023 707 se
rect 5023 682 5069 2807
tri 5069 2765 5111 2807 nw
rect 5191 2849 5357 5033
tri 5437 5072 5479 5114 se
rect 5479 5072 5525 7246
tri 5525 7204 5567 7246 nw
rect 5647 7287 5870 9490
rect 5647 7253 5713 7287
rect 5747 7253 5870 7287
tri 5525 5072 5567 5114 sw
rect 5437 5066 5567 5072
rect 5437 5032 5449 5066
rect 5483 5032 5521 5066
rect 5555 5032 5567 5066
rect 5437 5026 5567 5032
tri 5437 4984 5479 5026 ne
rect 5191 2815 5221 2849
rect 5255 2815 5293 2849
rect 5327 2815 5357 2849
tri 5069 682 5094 707 sw
rect 4945 676 5147 682
rect 4945 642 4957 676
rect 4991 642 5029 676
rect 5063 642 5101 676
rect 5135 642 5147 676
rect 4945 636 5147 642
tri 4901 597 4926 622 sw
tri 5166 597 5191 622 se
rect 5191 597 5357 2815
tri 5437 2853 5479 2895 se
rect 5479 2853 5525 5026
tri 5525 4984 5567 5026 nw
rect 5647 5067 5870 7253
tri 7831 6185 7858 6212 nw
tri 8308 6185 8335 6212 ne
rect 5647 5033 5713 5067
rect 5747 5033 5870 5067
tri 5525 2853 5567 2895 sw
rect 5437 2847 5567 2853
rect 5437 2813 5449 2847
rect 5483 2813 5521 2847
rect 5555 2813 5567 2847
rect 5437 2807 5567 2813
tri 5437 2765 5479 2807 ne
tri 5454 682 5479 707 se
rect 5479 682 5525 2807
tri 5525 2765 5567 2807 nw
rect 5647 2848 5870 5033
rect 5647 2814 5713 2848
rect 5747 2814 5870 2848
tri 5525 682 5550 707 sw
rect 5401 676 5603 682
rect 5401 642 5413 676
rect 5447 642 5485 676
rect 5519 642 5557 676
rect 5591 642 5603 676
rect 5401 636 5603 642
tri 5637 622 5647 632 se
rect 5647 622 5870 2814
tri 7776 2091 7785 2100 se
tri 7754 2069 7776 2091 se
rect 7776 2069 7785 2091
tri 7831 2091 7840 2100 sw
tri 8326 2091 8335 2100 se
rect 7831 2082 7840 2091
tri 7840 2082 7849 2091 sw
tri 8317 2082 8326 2091 se
rect 8326 2082 8335 2091
rect 7831 2078 7849 2082
tri 7849 2078 7853 2082 sw
tri 8313 2078 8317 2082 se
rect 8317 2078 8335 2082
rect 7831 2069 7853 2078
tri 7853 2069 7862 2078 sw
tri 8304 2069 8313 2078 se
rect 8313 2069 8335 2078
tri 8381 2091 8390 2100 sw
rect 8381 2082 8390 2091
tri 8390 2082 8399 2091 sw
rect 8381 2078 8399 2082
tri 8399 2078 8403 2082 sw
rect 8381 2069 8403 2078
tri 8403 2069 8412 2078 sw
tri 5357 597 5382 622 sw
tri 5612 597 5637 622 se
rect 5637 597 5870 622
tri 534 591 540 597 ne
rect 540 591 5870 597
tri 540 557 574 591 ne
rect 574 557 618 591
rect 652 557 690 591
rect 724 557 762 591
rect 796 557 834 591
rect 868 557 906 591
rect 940 557 978 591
rect 1012 557 3907 591
rect 3941 557 3979 591
rect 4013 557 4051 591
rect 4085 557 4123 591
rect 4157 557 4195 591
rect 4229 557 4267 591
rect 4301 557 4339 591
rect 4373 557 4575 591
rect 4609 557 4647 591
rect 4681 557 4719 591
rect 4753 557 4791 591
rect 4825 557 5047 591
rect 5081 557 5119 591
rect 5153 557 5191 591
rect 5225 557 5446 591
rect 5480 557 5518 591
rect 5552 557 5590 591
rect 5624 557 5662 591
rect 5696 557 5734 591
rect 5768 557 5870 591
tri 574 551 580 557 ne
rect 580 551 5870 557
rect 811 458 817 510
rect 869 458 881 510
rect 933 458 945 510
rect 997 458 1003 510
rect 1004 459 1005 509
rect 1041 459 1042 509
rect 1043 501 1173 510
rect 1043 467 1055 501
rect 1089 467 1127 501
rect 1161 467 1173 501
rect 1043 458 1173 467
rect 1767 458 1773 510
rect 1825 458 1837 510
rect 1889 458 1901 510
rect 1953 458 1959 510
rect 1960 459 1961 509
rect 1997 459 1998 509
rect 1999 501 2129 510
rect 1999 467 2011 501
rect 2045 467 2083 501
rect 2117 467 2129 501
rect 1999 458 2129 467
rect 2921 501 3051 510
rect 2921 467 2933 501
rect 2967 467 3005 501
rect 3039 467 3051 501
rect 2921 458 3051 467
rect 3052 459 3053 509
rect 3089 459 3090 509
rect 3091 458 3097 510
rect 3149 458 3161 510
rect 3213 458 3225 510
rect 3277 458 3283 510
rect 3502 458 3508 510
rect 3560 458 3572 510
rect 3624 458 3636 510
rect 3688 458 3694 510
rect 3695 459 3696 509
rect 3732 459 3733 509
rect 3734 501 3864 510
rect 3734 467 3746 501
rect 3780 467 3818 501
rect 3852 467 3864 501
rect 3734 458 3864 467
rect 4409 501 4539 510
rect 4409 467 4421 501
rect 4455 467 4493 501
rect 4527 467 4539 501
rect 4409 458 4539 467
rect 4540 459 4541 509
rect 4577 459 4578 509
rect 4579 458 4585 510
rect 4637 458 4649 510
rect 4701 458 4825 510
rect 4826 459 4827 509
rect 4863 459 4864 509
rect 4865 501 4995 510
rect 4865 467 4877 501
rect 4911 467 4949 501
rect 4983 467 4995 501
rect 4865 458 4995 467
rect 5267 501 5397 510
rect 5267 467 5279 501
rect 5313 467 5351 501
rect 5385 467 5397 501
rect 5267 458 5397 467
rect 5398 459 5399 509
rect 5435 459 5436 509
rect 5437 458 5443 510
rect 5495 458 5507 510
rect 5559 458 5565 510
tri 6027 447 6028 448 se
rect 6028 447 6059 448
rect 122 408 392 447
tri 392 408 431 447 sw
tri 5988 408 6027 447 se
rect 6027 408 6059 447
rect 122 362 437 408
rect 5967 362 6059 408
<< rmetal1 >>
rect 10680 34465 10682 34466
rect 10680 34415 10681 34465
rect 10680 34414 10682 34415
rect 10718 34465 10720 34466
rect 10719 34415 10720 34465
rect 10718 34414 10720 34415
rect 10952 34465 10954 34466
rect 10952 34415 10953 34465
rect 10952 34414 10954 34415
rect 10990 34465 10992 34466
rect 10991 34415 10992 34465
rect 13978 34465 13980 34466
rect 14016 34465 14018 34466
rect 10990 34414 10992 34415
rect 13978 34415 13979 34465
rect 14017 34415 14018 34465
rect 13978 34414 13980 34415
rect 14016 34414 14018 34415
rect 13978 33725 13980 33726
rect 14016 33725 14018 33726
rect 13978 33675 13979 33725
rect 14017 33675 14018 33725
rect 13978 33674 13980 33675
rect 14016 33674 14018 33675
rect 10952 32213 10954 32214
rect 10952 32163 10953 32213
rect 10952 32162 10954 32163
rect 10990 32213 10992 32214
rect 10991 32163 10992 32213
rect 13978 32213 13980 32214
rect 14016 32213 14018 32214
rect 10990 32162 10992 32163
rect 13978 32163 13979 32213
rect 14017 32163 14018 32213
rect 13978 32162 13980 32163
rect 14016 32162 14018 32163
rect 10952 29964 10954 29965
rect 10952 29914 10953 29964
rect 10952 29913 10954 29914
rect 10990 29964 10992 29965
rect 10991 29914 10992 29964
rect 13978 29964 13980 29965
rect 14016 29964 14018 29965
rect 10990 29913 10992 29914
rect 13978 29914 13979 29964
rect 14017 29914 14018 29964
rect 13978 29913 13980 29914
rect 14016 29913 14018 29914
rect 469 16783 471 16784
rect 469 16739 470 16783
rect 469 16738 471 16739
rect 507 16783 509 16784
rect 508 16739 509 16783
rect 1244 16783 1246 16784
rect 1282 16783 1284 16784
rect 507 16738 509 16739
rect 1244 16739 1245 16783
rect 1283 16739 1284 16783
rect 1244 16738 1246 16739
rect 1282 16738 1284 16739
rect 1382 16783 1384 16784
rect 1420 16783 1422 16784
rect 1382 16739 1383 16783
rect 1421 16739 1422 16783
rect 2157 16783 2159 16784
rect 1382 16738 1384 16739
rect 1420 16738 1422 16739
rect 2157 16739 2158 16783
rect 2157 16738 2159 16739
rect 2195 16783 2197 16784
rect 2196 16739 2197 16783
rect 2195 16738 2197 16739
rect 2839 16783 2841 16784
rect 2839 16739 2840 16783
rect 2839 16738 2841 16739
rect 2877 16783 2879 16784
rect 2878 16739 2879 16783
rect 3614 16783 3616 16784
rect 3652 16783 3654 16784
rect 2877 16738 2879 16739
rect 3614 16739 3615 16783
rect 3653 16739 3654 16783
rect 3614 16738 3616 16739
rect 3652 16738 3654 16739
rect 3752 16783 3754 16784
rect 3790 16783 3792 16784
rect 3752 16739 3753 16783
rect 3791 16739 3792 16783
rect 4527 16783 4529 16784
rect 3752 16738 3754 16739
rect 3790 16738 3792 16739
rect 4527 16739 4528 16783
rect 4527 16738 4529 16739
rect 4565 16783 4567 16784
rect 4566 16739 4567 16783
rect 4565 16738 4567 16739
rect 854 15292 900 15293
rect 854 15291 855 15292
rect 899 15291 900 15292
rect 854 15254 855 15255
rect 899 15254 900 15255
rect 854 15253 900 15254
rect 1766 15292 1812 15293
rect 1766 15291 1767 15292
rect 1811 15291 1812 15292
rect 1766 15254 1767 15255
rect 1811 15254 1812 15255
rect 1766 15253 1812 15254
rect 854 13762 900 13763
rect 854 13761 855 13762
rect 899 13761 900 13762
rect 854 13724 855 13725
rect 899 13724 900 13725
rect 854 13723 900 13724
rect 3224 15292 3270 15293
rect 3224 15291 3225 15292
rect 3269 15291 3270 15292
rect 3224 15254 3225 15255
rect 3269 15254 3270 15255
rect 3224 15253 3270 15254
rect 1766 13762 1812 13763
rect 1766 13761 1767 13762
rect 1811 13761 1812 13762
rect 1766 13724 1767 13725
rect 1811 13724 1812 13725
rect 1766 13723 1812 13724
rect 854 12232 900 12233
rect 854 12231 855 12232
rect 899 12231 900 12232
rect 854 12194 855 12195
rect 899 12194 900 12195
rect 854 12193 900 12194
rect 4136 15292 4182 15293
rect 4136 15291 4137 15292
rect 4181 15291 4182 15292
rect 4136 15254 4137 15255
rect 4181 15254 4182 15255
rect 4136 15253 4182 15254
rect 3224 13762 3270 13763
rect 3224 13761 3225 13762
rect 3269 13761 3270 13762
rect 3224 13724 3225 13725
rect 3269 13724 3270 13725
rect 3224 13723 3270 13724
rect 3224 12269 3270 12270
rect 4136 13762 4182 13763
rect 4136 13761 4137 13762
rect 4181 13761 4182 13762
rect 4136 13724 4137 13725
rect 4181 13724 4182 13725
rect 4136 13723 4182 13724
rect 3224 12268 3225 12269
rect 3269 12268 3270 12269
rect 1766 12232 1812 12233
rect 1766 12231 1767 12232
rect 1811 12231 1812 12232
rect 1766 12194 1767 12195
rect 1811 12194 1812 12195
rect 1766 12193 1812 12194
rect 3224 12231 3225 12232
rect 3269 12231 3270 12232
rect 3224 12230 3270 12231
rect 4136 12232 4182 12233
rect 4136 12231 4137 12232
rect 4181 12231 4182 12232
rect 4136 12194 4137 12195
rect 4181 12194 4182 12195
rect 4136 12193 4182 12194
rect 5350 15065 5396 15066
rect 5350 15064 5351 15065
rect 5395 15064 5396 15065
rect 5350 15027 5351 15028
rect 5395 15027 5396 15028
rect 5350 15026 5396 15027
rect 5320 14706 5378 14707
rect 5320 14705 5321 14706
rect 5377 14705 5378 14706
rect 5600 14706 5658 14707
rect 5600 14705 5601 14706
rect 5657 14705 5658 14706
rect 5320 14668 5321 14669
rect 5377 14668 5378 14669
rect 5320 14667 5378 14668
rect 5600 14668 5601 14669
rect 5657 14668 5658 14669
rect 5600 14667 5658 14668
rect 5880 14706 5938 14707
rect 5880 14705 5881 14706
rect 5937 14705 5938 14706
rect 5880 14668 5881 14669
rect 5937 14668 5938 14669
rect 5880 14667 5938 14668
rect 5320 10426 5378 10427
rect 5320 10425 5321 10426
rect 5377 10425 5378 10426
rect 5460 10426 5518 10427
rect 5460 10425 5461 10426
rect 5517 10425 5518 10426
rect 5740 10426 5798 10427
rect 5740 10425 5741 10426
rect 5797 10425 5798 10426
rect 6020 10426 6078 10427
rect 6020 10425 6021 10426
rect 6077 10425 6078 10426
rect 5320 10388 5321 10389
rect 5377 10388 5378 10389
rect 5320 10387 5378 10388
rect 5320 10268 5378 10269
rect 5320 10267 5321 10268
rect 5377 10267 5378 10268
rect 5460 10388 5461 10389
rect 5517 10388 5518 10389
rect 5460 10387 5518 10388
rect 5740 10388 5741 10389
rect 5797 10388 5798 10389
rect 5740 10387 5798 10388
rect 6020 10388 6021 10389
rect 6077 10388 6078 10389
rect 6020 10387 6078 10388
rect 5460 10268 5518 10269
rect 5460 10267 5461 10268
rect 5517 10267 5518 10268
rect 5320 10230 5321 10231
rect 5377 10230 5378 10231
rect 5320 10229 5378 10230
rect 5460 10230 5461 10231
rect 5517 10230 5518 10231
rect 5460 10229 5518 10230
rect 5740 10268 5798 10269
rect 5740 10267 5741 10268
rect 5797 10267 5798 10268
rect 5740 10230 5741 10231
rect 5797 10230 5798 10231
rect 5740 10229 5798 10230
rect 6020 10268 6078 10269
rect 6020 10267 6021 10268
rect 6077 10267 6078 10268
rect 6020 10230 6021 10231
rect 6077 10230 6078 10231
rect 6020 10229 6078 10230
rect 1079 9546 1125 9547
rect 1079 9545 1080 9546
rect 1124 9545 1125 9546
rect 1079 9508 1080 9509
rect 1124 9508 1125 9509
rect 1079 9507 1125 9508
rect 1935 9546 1981 9547
rect 1935 9545 1936 9546
rect 1980 9545 1981 9546
rect 1935 9508 1936 9509
rect 1980 9508 1981 9509
rect 1935 9507 1981 9508
rect 2791 9546 2837 9547
rect 2791 9545 2792 9546
rect 2836 9545 2837 9546
rect 2791 9508 2792 9509
rect 2836 9508 2837 9509
rect 2791 9507 2837 9508
rect 3911 9546 3957 9547
rect 3911 9545 3912 9546
rect 3956 9545 3957 9546
rect 3911 9508 3912 9509
rect 3956 9508 3957 9509
rect 3911 9507 3957 9508
rect 4567 9546 4613 9547
rect 4567 9545 4568 9546
rect 4612 9545 4613 9546
rect 4567 9508 4568 9509
rect 4612 9508 4613 9509
rect 4567 9507 4613 9508
rect 5023 9546 5069 9547
rect 5023 9545 5024 9546
rect 5068 9545 5069 9546
rect 5023 9508 5024 9509
rect 5068 9508 5069 9509
rect 5023 9507 5069 9508
rect 5479 9546 5525 9547
rect 5479 9545 5480 9546
rect 5524 9545 5525 9546
rect 5479 9508 5480 9509
rect 5524 9508 5525 9509
rect 5479 9507 5525 9508
rect 1003 509 1005 510
rect 1003 459 1004 509
rect 1003 458 1005 459
rect 1041 509 1043 510
rect 1042 459 1043 509
rect 1041 458 1043 459
rect 1959 509 1961 510
rect 1959 459 1960 509
rect 1959 458 1961 459
rect 1997 509 1999 510
rect 1998 459 1999 509
rect 1997 458 1999 459
rect 3051 509 3053 510
rect 3051 459 3052 509
rect 3051 458 3053 459
rect 3089 509 3091 510
rect 3090 459 3091 509
rect 3089 458 3091 459
rect 3694 509 3696 510
rect 3694 459 3695 509
rect 3694 458 3696 459
rect 3732 509 3734 510
rect 3733 459 3734 509
rect 3732 458 3734 459
rect 4539 509 4541 510
rect 4539 459 4540 509
rect 4539 458 4541 459
rect 4577 509 4579 510
rect 4578 459 4579 509
rect 4577 458 4579 459
rect 4825 509 4827 510
rect 4825 459 4826 509
rect 4825 458 4827 459
rect 4863 509 4865 510
rect 4864 459 4865 509
rect 4863 458 4865 459
rect 5397 509 5399 510
rect 5397 459 5398 509
rect 5397 458 5399 459
rect 5435 509 5437 510
rect 5436 459 5437 509
rect 5435 458 5437 459
<< via1 >>
rect 12378 34546 12430 34555
rect 12459 34546 12511 34555
rect 12540 34546 12592 34555
rect 12620 34546 12672 34555
rect 12378 34512 12384 34546
rect 12384 34512 12422 34546
rect 12422 34512 12430 34546
rect 12459 34512 12494 34546
rect 12494 34512 12511 34546
rect 12540 34512 12566 34546
rect 12566 34512 12592 34546
rect 12620 34512 12638 34546
rect 12638 34512 12672 34546
rect 12378 34503 12430 34512
rect 12459 34503 12511 34512
rect 12540 34503 12592 34512
rect 12620 34503 12672 34512
rect 10506 34454 10558 34466
rect 10506 34420 10510 34454
rect 10510 34420 10544 34454
rect 10544 34420 10558 34454
rect 10506 34414 10558 34420
rect 10570 34454 10622 34466
rect 10570 34420 10582 34454
rect 10582 34420 10616 34454
rect 10616 34420 10622 34454
rect 10570 34414 10622 34420
rect 10778 34414 10830 34466
rect 10842 34414 10894 34466
rect 14070 34408 14122 34460
rect 14070 34344 14122 34396
rect 14070 33744 14122 33796
rect 10506 33674 10558 33726
rect 10570 33674 10622 33726
rect 14070 33680 14122 33732
rect 12378 33527 12430 33579
rect 12459 33527 12511 33579
rect 12540 33527 12592 33579
rect 12620 33527 12672 33579
rect 12378 33451 12430 33503
rect 12459 33451 12511 33503
rect 12540 33451 12592 33503
rect 12620 33451 12672 33503
rect 12378 33375 12430 33427
rect 12459 33375 12511 33427
rect 12540 33375 12592 33427
rect 12620 33375 12672 33427
rect 12378 33299 12430 33351
rect 12459 33299 12511 33351
rect 12540 33299 12592 33351
rect 12620 33299 12672 33351
rect 12378 33223 12430 33275
rect 12459 33223 12511 33275
rect 12540 33223 12592 33275
rect 12620 33223 12672 33275
rect 12378 33147 12430 33199
rect 12459 33147 12511 33199
rect 12540 33147 12592 33199
rect 12620 33147 12672 33199
rect 12378 32294 12430 32303
rect 12459 32294 12511 32303
rect 12540 32294 12592 32303
rect 12620 32294 12672 32303
rect 12378 32260 12393 32294
rect 12393 32260 12430 32294
rect 12459 32260 12465 32294
rect 12465 32260 12503 32294
rect 12503 32260 12511 32294
rect 12540 32260 12575 32294
rect 12575 32260 12592 32294
rect 12620 32260 12647 32294
rect 12647 32260 12672 32294
rect 12378 32251 12430 32260
rect 12459 32251 12511 32260
rect 12540 32251 12592 32260
rect 12620 32251 12672 32260
rect 10506 32202 10558 32214
rect 10570 32202 10622 32214
rect 10506 32168 10508 32202
rect 10508 32168 10558 32202
rect 10570 32168 10593 32202
rect 10593 32168 10622 32202
rect 10506 32162 10558 32168
rect 10570 32162 10622 32168
rect 10778 32162 10830 32214
rect 10842 32162 10894 32214
rect 14070 32156 14122 32208
rect 14070 32092 14122 32144
rect 11788 31242 11840 31294
rect 11892 31282 11944 31294
rect 11892 31248 11908 31282
rect 11908 31248 11944 31282
rect 11892 31242 11944 31248
rect 12378 31242 12430 31294
rect 12459 31242 12511 31294
rect 12540 31242 12592 31294
rect 12620 31242 12672 31294
rect 11788 31166 11840 31218
rect 11892 31207 11944 31218
rect 11892 31173 11908 31207
rect 11908 31173 11944 31207
rect 11892 31166 11944 31173
rect 12378 31166 12430 31218
rect 12459 31166 12511 31218
rect 12540 31166 12592 31218
rect 12620 31166 12672 31218
rect 11788 31090 11840 31142
rect 11892 31132 11944 31142
rect 11892 31098 11908 31132
rect 11908 31098 11944 31132
rect 11892 31090 11944 31098
rect 12378 31090 12430 31142
rect 12459 31090 12511 31142
rect 12540 31090 12592 31142
rect 12620 31090 12672 31142
rect 11788 31014 11840 31066
rect 11892 31057 11944 31066
rect 11892 31023 11908 31057
rect 11908 31023 11944 31057
rect 11892 31014 11944 31023
rect 12378 31014 12430 31066
rect 12459 31014 12511 31066
rect 12540 31014 12592 31066
rect 12620 31014 12672 31066
rect 11788 30938 11840 30990
rect 11892 30982 11944 30990
rect 11892 30948 11908 30982
rect 11908 30948 11944 30982
rect 11892 30938 11944 30948
rect 12378 30938 12430 30990
rect 12459 30938 12511 30990
rect 12540 30938 12592 30990
rect 12620 30938 12672 30990
rect 11788 30862 11840 30914
rect 11892 30908 11944 30914
rect 11892 30874 11908 30908
rect 11908 30874 11944 30908
rect 11892 30862 11944 30874
rect 12378 30862 12430 30914
rect 12459 30862 12511 30914
rect 12540 30862 12592 30914
rect 12620 30862 12672 30914
rect 11788 30043 11840 30052
rect 11892 30043 11944 30052
rect 11788 30009 11817 30043
rect 11817 30009 11840 30043
rect 11892 30009 11927 30043
rect 11927 30009 11944 30043
rect 11788 30000 11840 30009
rect 11892 30000 11944 30009
rect 10506 29953 10558 29965
rect 10570 29953 10622 29965
rect 10506 29919 10508 29953
rect 10508 29919 10558 29953
rect 10570 29919 10593 29953
rect 10593 29919 10622 29953
rect 10506 29913 10558 29919
rect 10570 29913 10622 29919
rect 10778 29913 10830 29965
rect 10842 29913 10894 29965
rect 14070 29907 14122 29959
rect 14070 29843 14122 29895
rect 14070 29395 14122 29447
rect 14070 29331 14122 29383
rect 9721 29188 9773 29240
rect 9811 29188 9863 29240
rect 10772 29188 10824 29240
rect 10848 29188 10900 29240
rect 9721 29110 9773 29162
rect 9811 29110 9863 29162
rect 10772 29110 10824 29162
rect 10848 29110 10900 29162
rect 4301 29019 4353 29071
rect 4365 29019 4417 29071
rect 5624 28907 5676 28959
rect 5730 28907 5782 28959
rect 5836 28907 5888 28959
rect 11788 28938 11840 28990
rect 11892 28978 11944 28990
rect 11892 28944 11908 28978
rect 11908 28944 11944 28978
rect 11892 28938 11944 28944
rect 5624 28822 5676 28874
rect 5730 28822 5782 28874
rect 5836 28822 5888 28874
rect 11788 28862 11840 28914
rect 11892 28903 11944 28914
rect 11892 28869 11908 28903
rect 11908 28869 11944 28903
rect 11892 28862 11944 28869
rect 5624 28736 5676 28788
rect 5730 28736 5782 28788
rect 5836 28736 5888 28788
rect 11788 28786 11840 28838
rect 11892 28828 11944 28838
rect 11892 28794 11908 28828
rect 11908 28794 11944 28828
rect 11892 28786 11944 28794
rect 5624 28650 5676 28702
rect 5730 28650 5782 28702
rect 5836 28650 5888 28702
rect 11788 28710 11840 28762
rect 11892 28753 11944 28762
rect 11892 28719 11908 28753
rect 11908 28719 11944 28753
rect 11892 28710 11944 28719
rect 5624 28564 5676 28616
rect 5730 28564 5782 28616
rect 5836 28564 5888 28616
rect 11788 28634 11840 28686
rect 11892 28678 11944 28686
rect 11892 28644 11908 28678
rect 11908 28644 11944 28678
rect 11892 28634 11944 28644
rect 11788 28558 11840 28610
rect 11892 28604 11944 28610
rect 11892 28570 11908 28604
rect 11908 28570 11944 28604
rect 11892 28558 11944 28570
rect 10506 27076 10558 27128
rect 10570 27076 10622 27128
rect -236 17223 -184 17275
rect -172 17223 -120 17275
rect -29 17189 151 17195
rect -29 17155 130 17189
rect 130 17155 151 17189
rect -29 17117 151 17155
rect -29 17083 130 17117
rect 130 17083 151 17117
rect -29 17079 151 17083
rect 207 16951 387 17067
rect 2310 16862 2362 16914
rect 2374 16862 2426 16914
rect 2438 16862 2490 16914
rect 2502 16862 2554 16914
rect 2793 16871 2845 16923
rect 2857 16871 2909 16923
rect 4295 16596 4347 16648
rect 4295 16532 4347 16584
rect 4361 12257 4413 12309
rect 4361 12233 4413 12245
rect 4361 12199 4370 12233
rect 4370 12199 4404 12233
rect 4404 12199 4413 12233
rect 4361 12193 4413 12199
rect 5158 15186 5180 15218
rect 5180 15186 5210 15218
rect 5158 15166 5210 15186
rect 5158 15148 5210 15154
rect 5158 15114 5180 15148
rect 5180 15114 5210 15148
rect 5158 15102 5210 15114
rect 5507 15186 5532 15218
rect 5532 15186 5559 15218
rect 5507 15166 5559 15186
rect 5507 15148 5559 15154
rect 5507 15114 5532 15148
rect 5532 15114 5559 15148
rect 5507 15102 5559 15114
rect 5961 15093 6077 15273
rect 6283 15093 6399 15273
rect 6161 14888 6213 14940
rect 6161 14824 6213 14876
rect 6155 14660 6207 14666
rect 6155 14626 6172 14660
rect 6172 14626 6206 14660
rect 6206 14626 6207 14660
rect 6155 14614 6207 14626
rect 6155 14588 6207 14602
rect 6155 14554 6172 14588
rect 6172 14554 6206 14588
rect 6206 14554 6207 14588
rect 6155 14550 6207 14554
rect 4421 11894 4473 11946
rect 4421 11830 4473 11882
rect 5303 10516 5355 10568
rect 5303 10452 5355 10504
rect 5627 10458 5679 10510
rect 5695 10458 5747 10510
rect 5763 10458 5815 10510
rect 5831 10458 5883 10510
rect 6155 10381 6207 10387
rect 6155 10347 6172 10381
rect 6172 10347 6206 10381
rect 6206 10347 6207 10381
rect 6155 10335 6207 10347
rect 6155 10309 6207 10323
rect 6155 10275 6172 10309
rect 6172 10275 6206 10309
rect 6206 10275 6207 10309
rect 6155 10271 6207 10275
rect 2297 9687 2349 9739
rect 2361 9687 2413 9739
rect 2425 9687 2477 9739
rect 2489 9687 2541 9739
rect 2553 9687 2605 9739
rect 2617 9687 2669 9739
rect 2681 9687 2733 9739
rect 4781 9687 4833 9739
rect 4845 9687 4897 9739
rect 5303 9544 5355 9550
rect 5303 9510 5329 9544
rect 5329 9510 5355 9544
rect 5303 9498 5355 9510
rect 5303 9434 5355 9486
rect 817 458 869 510
rect 881 458 933 510
rect 945 458 997 510
rect 1773 458 1825 510
rect 1837 458 1889 510
rect 1901 458 1953 510
rect 3097 458 3149 510
rect 3161 458 3213 510
rect 3225 458 3277 510
rect 3508 458 3560 510
rect 3572 458 3624 510
rect 3636 458 3688 510
rect 4585 458 4637 510
rect 4649 458 4701 510
rect 5443 458 5495 510
rect 5507 458 5559 510
<< metal2 >>
rect 12372 34503 12378 34555
rect 12430 34503 12459 34555
rect 12511 34503 12540 34555
rect 12592 34503 12620 34555
rect 12672 34503 12678 34555
rect 10500 34414 10506 34466
rect 10558 34414 10570 34466
rect 10622 34414 10628 34466
rect 10500 33726 10628 34414
rect 10500 33674 10506 33726
rect 10558 33674 10570 33726
rect 10622 33674 10628 33726
rect 10500 32214 10628 33674
rect 10500 32162 10506 32214
rect 10558 32162 10570 32214
rect 10622 32162 10628 32214
rect 10500 29965 10628 32162
rect 10500 29913 10506 29965
rect 10558 29913 10570 29965
rect 10622 29913 10628 29965
rect 9721 29240 9863 29246
rect 9773 29188 9811 29240
rect 9721 29162 9863 29188
rect 9773 29110 9811 29162
rect 4295 29019 4301 29071
rect 4353 29019 4365 29071
rect 4417 29019 4423 29071
rect 4295 28990 4364 29019
tri 4364 28990 4393 29019 nw
rect 4295 27614 4347 28990
tri 4347 28973 4364 28990 nw
rect 5621 28959 5889 28969
rect 5621 28907 5624 28959
rect 5676 28907 5730 28959
rect 5782 28907 5836 28959
rect 5888 28907 5889 28959
rect 5621 28874 5889 28907
rect 5621 28822 5624 28874
rect 5676 28822 5730 28874
rect 5782 28822 5836 28874
rect 5888 28822 5889 28874
rect 5621 28788 5889 28822
rect 5621 28736 5624 28788
rect 5676 28736 5730 28788
rect 5782 28736 5836 28788
rect 5888 28736 5889 28788
rect 5621 28702 5889 28736
rect 5621 28650 5624 28702
rect 5676 28650 5730 28702
rect 5782 28650 5836 28702
rect 5888 28650 5889 28702
rect 5621 28616 5889 28650
tri 9712 28634 9721 28643 se
rect 9721 28634 9863 29110
rect 5621 28564 5624 28616
rect 5676 28564 5730 28616
rect 5782 28564 5836 28616
rect 5888 28564 5889 28616
tri 9688 28610 9712 28634 se
rect 9712 28610 9863 28634
tri 9644 28566 9688 28610 se
rect 9688 28583 9863 28610
rect 9688 28566 9846 28583
tri 9846 28566 9863 28583 nw
rect 5621 28041 5889 28564
tri 9272 28558 9280 28566 se
rect 9280 28558 9838 28566
tri 9838 28558 9846 28566 nw
tri 9133 28419 9272 28558 se
rect 9272 28424 9704 28558
tri 9704 28424 9838 28558 nw
rect 9272 28419 9335 28424
tri 9335 28419 9340 28424 nw
rect 5621 28034 5882 28041
tri 5882 28034 5889 28041 nw
tri 9056 28034 9133 28111 se
rect 9133 28051 9275 28419
tri 9275 28359 9335 28419 nw
rect 9133 28034 9258 28051
tri 9258 28034 9275 28051 nw
rect 5621 27837 5810 28034
tri 5810 27962 5882 28034 nw
tri 5810 27837 5871 27898 sw
rect 8805 27892 9116 28034
tri 9116 27892 9258 28034 nw
tri 8805 27837 8860 27892 nw
rect 5621 27819 5871 27837
tri 5871 27819 5889 27837 sw
rect 5621 27614 5889 27819
rect 10500 27128 10628 29913
rect 10772 34414 10778 34466
rect 10830 34414 10842 34466
rect 10894 34414 10900 34466
rect 10772 32214 10900 34414
rect 10772 32162 10778 32214
rect 10830 32162 10842 32214
rect 10894 32162 10900 32214
rect 10772 29965 10900 32162
rect 12372 33579 12678 34503
rect 12372 33527 12378 33579
rect 12430 33527 12459 33579
rect 12511 33527 12540 33579
rect 12592 33527 12620 33579
rect 12672 33527 12678 33579
rect 12372 33503 12678 33527
rect 12372 33451 12378 33503
rect 12430 33451 12459 33503
rect 12511 33451 12540 33503
rect 12592 33451 12620 33503
rect 12672 33451 12678 33503
rect 12372 33427 12678 33451
rect 12372 33375 12378 33427
rect 12430 33375 12459 33427
rect 12511 33375 12540 33427
rect 12592 33375 12620 33427
rect 12672 33375 12678 33427
rect 12372 33351 12678 33375
rect 12372 33299 12378 33351
rect 12430 33299 12459 33351
rect 12511 33299 12540 33351
rect 12592 33299 12620 33351
rect 12672 33299 12678 33351
rect 12372 33275 12678 33299
rect 12372 33223 12378 33275
rect 12430 33223 12459 33275
rect 12511 33223 12540 33275
rect 12592 33223 12620 33275
rect 12672 33223 12678 33275
rect 12372 33199 12678 33223
rect 12372 33147 12378 33199
rect 12430 33147 12459 33199
rect 12511 33147 12540 33199
rect 12592 33147 12620 33199
rect 12672 33147 12678 33199
rect 12372 32303 12678 33147
rect 12372 32251 12378 32303
rect 12430 32251 12459 32303
rect 12511 32251 12540 32303
rect 12592 32251 12620 32303
rect 12672 32251 12678 32303
rect 12372 31294 12678 32251
rect 10772 29913 10778 29965
rect 10830 29913 10842 29965
rect 10894 29913 10900 29965
rect 10772 29240 10900 29913
rect 10824 29188 10848 29240
rect 10772 29162 10900 29188
rect 10824 29110 10848 29162
rect 10772 29104 10900 29110
rect 11782 31242 11788 31294
rect 11840 31242 11892 31294
rect 11944 31242 11950 31294
rect 11782 31218 11950 31242
rect 11782 31166 11788 31218
rect 11840 31166 11892 31218
rect 11944 31166 11950 31218
rect 11782 31142 11950 31166
rect 11782 31090 11788 31142
rect 11840 31090 11892 31142
rect 11944 31090 11950 31142
rect 11782 31066 11950 31090
rect 11782 31014 11788 31066
rect 11840 31014 11892 31066
rect 11944 31014 11950 31066
rect 11782 30990 11950 31014
rect 11782 30938 11788 30990
rect 11840 30938 11892 30990
rect 11944 30938 11950 30990
rect 11782 30914 11950 30938
rect 11782 30862 11788 30914
rect 11840 30862 11892 30914
rect 11944 30862 11950 30914
rect 12372 31242 12378 31294
rect 12430 31242 12459 31294
rect 12511 31242 12540 31294
rect 12592 31242 12620 31294
rect 12672 31242 12678 31294
rect 12372 31218 12678 31242
rect 12372 31166 12378 31218
rect 12430 31166 12459 31218
rect 12511 31166 12540 31218
rect 12592 31166 12620 31218
rect 12672 31166 12678 31218
rect 12372 31142 12678 31166
rect 12372 31090 12378 31142
rect 12430 31090 12459 31142
rect 12511 31090 12540 31142
rect 12592 31090 12620 31142
rect 12672 31090 12678 31142
rect 12372 31066 12678 31090
rect 12372 31014 12378 31066
rect 12430 31014 12459 31066
rect 12511 31014 12540 31066
rect 12592 31014 12620 31066
rect 12672 31014 12678 31066
rect 12372 30990 12678 31014
rect 12372 30938 12378 30990
rect 12430 30938 12459 30990
rect 12511 30938 12540 30990
rect 12592 30938 12620 30990
rect 12672 30938 12678 30990
rect 12372 30914 12678 30938
rect 12372 30862 12378 30914
rect 12430 30862 12459 30914
rect 12511 30862 12540 30914
rect 12592 30862 12620 30914
rect 12672 30862 12678 30914
rect 14070 34460 14198 34466
rect 14122 34408 14198 34460
rect 14070 34396 14198 34408
rect 14122 34344 14198 34396
rect 14070 33796 14198 34344
rect 14122 33744 14198 33796
rect 14070 33732 14198 33744
rect 14122 33680 14198 33732
rect 14070 32208 14198 33680
rect 14122 32156 14198 32208
rect 14070 32144 14198 32156
rect 14122 32092 14198 32144
rect 11782 30052 11950 30862
rect 11782 30000 11788 30052
rect 11840 30000 11892 30052
rect 11944 30000 11950 30052
rect 11782 28990 11950 30000
rect 14070 29959 14198 32092
rect 14122 29907 14198 29959
rect 14070 29895 14198 29907
rect 14122 29843 14198 29895
rect 14070 29447 14198 29843
rect 14122 29395 14198 29447
rect 14070 29383 14198 29395
rect 14122 29331 14198 29383
rect 14070 29325 14198 29331
rect 11782 28938 11788 28990
rect 11840 28938 11892 28990
rect 11944 28938 11950 28990
rect 11782 28914 11950 28938
rect 11782 28862 11788 28914
rect 11840 28862 11892 28914
rect 11944 28862 11950 28914
rect 11782 28838 11950 28862
rect 11782 28786 11788 28838
rect 11840 28786 11892 28838
rect 11944 28786 11950 28838
rect 11782 28762 11950 28786
rect 11782 28710 11788 28762
rect 11840 28710 11892 28762
rect 11944 28710 11950 28762
rect 11782 28686 11950 28710
rect 11782 28634 11788 28686
rect 11840 28634 11892 28686
rect 11944 28634 11950 28686
rect 11782 28610 11950 28634
rect 11782 28558 11788 28610
rect 11840 28558 11892 28610
rect 11944 28558 11950 28610
rect 10500 27076 10506 27128
rect 10558 27076 10570 27128
rect 10622 27076 10628 27128
rect -242 17223 -236 17275
rect -184 17223 -172 17275
rect -120 17267 -114 17275
tri -114 17267 -106 17275 sw
rect -120 17223 -106 17267
tri -242 17201 -220 17223 ne
rect -220 17201 -106 17223
tri -220 17195 -214 17201 ne
rect -214 17195 -106 17201
tri -214 17139 -158 17195 ne
rect -158 341 -106 17195
rect -78 17195 151 17282
rect 265 17254 647 17282
tri 265 17201 318 17254 ne
rect 318 17201 647 17254
rect -78 17079 -29 17195
tri 318 17090 429 17201 ne
rect -78 16923 151 17079
rect 207 17067 388 17073
rect 387 17060 388 17067
tri 388 17060 401 17073 sw
rect 387 16951 401 17060
tri 151 16923 176 16948 sw
rect 207 16942 401 16951
tri 207 16923 226 16942 ne
rect 226 16923 401 16942
rect -78 16920 176 16923
tri 176 16920 179 16923 sw
tri 226 16920 229 16923 ne
rect 229 16920 401 16923
rect -78 16914 179 16920
tri 179 16914 185 16920 sw
tri 229 16914 235 16920 ne
rect 235 16914 401 16920
rect -78 16870 185 16914
tri 185 16870 229 16914 sw
tri 235 16870 279 16914 ne
rect 279 16870 401 16914
rect -78 341 229 16870
tri 279 16864 285 16870 ne
rect 285 12265 401 16870
tri 410 12193 429 12212 se
rect 429 12193 647 17201
tri 285 12068 410 12193 se
rect 410 12068 647 12193
rect 285 341 647 12068
rect 703 341 755 17282
rect 811 510 1057 17282
rect 811 458 817 510
rect 869 458 881 510
rect 933 458 945 510
rect 997 458 1057 510
rect 811 341 1057 458
rect 1113 341 1165 17282
rect 1221 17238 1603 17282
rect 1221 12257 1273 17238
tri 1273 17210 1301 17238 nw
tri 1481 17210 1509 17238 ne
tri 1301 16923 1320 16942 ne
rect 1320 16923 1462 16942
tri 1462 16923 1481 16942 nw
tri 1320 16914 1329 16923 ne
rect 1329 12309 1453 16923
tri 1453 16914 1462 16923 nw
tri 1273 12257 1294 12278 sw
tri 1488 12257 1509 12278 se
rect 1509 12257 1603 17238
rect 1221 12253 1294 12257
tri 1294 12253 1298 12257 sw
tri 1484 12253 1488 12257 se
rect 1488 12253 1603 12257
rect 1221 341 1603 12253
rect 1659 16862 1993 17282
rect 2185 17254 2455 17282
tri 2185 17201 2238 17254 ne
rect 2238 16993 2455 17254
tri 2455 16993 2497 17035 sw
rect 2238 16945 2497 16993
tri 2497 16945 2545 16993 sw
tri 2817 16953 2857 16993 se
rect 2857 16953 2909 16993
rect 2021 16939 2201 16942
tri 2021 16925 2035 16939 ne
rect 2035 16925 2201 16939
rect 2238 16928 2545 16945
tri 2238 16925 2241 16928 ne
rect 2241 16925 2545 16928
tri 2035 16923 2037 16925 ne
rect 2037 16923 2201 16925
tri 2201 16923 2203 16925 sw
tri 2241 16923 2243 16925 ne
rect 2243 16923 2545 16925
tri 2545 16923 2567 16945 sw
tri 2037 16914 2046 16923 ne
rect 2046 16914 2203 16923
tri 2203 16914 2212 16923 sw
tri 2243 16914 2252 16923 ne
rect 2252 16914 2567 16923
tri 2567 16914 2576 16923 sw
tri 2046 16911 2049 16914 ne
rect 2049 16911 2212 16914
tri 2212 16911 2215 16914 sw
tri 2252 16911 2255 16914 ne
rect 2255 16911 2310 16914
tri 2049 16887 2073 16911 ne
rect 2073 16887 2215 16911
tri 1993 16862 2018 16887 sw
tri 2073 16862 2098 16887 ne
rect 2098 16871 2215 16887
tri 2215 16871 2255 16911 sw
tri 2255 16871 2295 16911 ne
rect 2295 16871 2310 16911
rect 2098 16862 2255 16871
tri 2255 16862 2264 16871 sw
tri 2295 16862 2304 16871 ne
rect 2304 16862 2310 16871
rect 2362 16862 2374 16914
rect 2426 16862 2438 16914
rect 2490 16862 2502 16914
rect 2554 16891 2576 16914
tri 2576 16891 2599 16914 sw
rect 2554 16862 2599 16891
rect 1659 16807 2018 16862
tri 2018 16807 2073 16862 sw
tri 2098 16807 2153 16862 ne
rect 2153 16853 2264 16862
tri 2264 16853 2273 16862 sw
tri 2304 16853 2313 16862 ne
rect 2313 16853 2599 16862
rect 2153 16817 2273 16853
tri 2273 16817 2309 16853 sw
tri 2313 16817 2349 16853 ne
rect 2349 16817 2599 16853
rect 2153 16807 2309 16817
rect 1659 16759 2073 16807
tri 2073 16759 2121 16807 sw
tri 2153 16759 2201 16807 ne
rect 2201 16785 2309 16807
tri 2309 16785 2341 16817 sw
tri 2349 16785 2381 16817 ne
rect 2381 16785 2599 16817
rect 2201 16759 2341 16785
rect 1659 16751 2121 16759
tri 2121 16751 2129 16759 sw
tri 2201 16751 2209 16759 ne
rect 2209 16751 2341 16759
rect 1659 16745 2129 16751
tri 2129 16745 2135 16751 sw
tri 2209 16745 2215 16751 ne
rect 2215 16745 2341 16751
tri 2341 16745 2381 16785 sw
tri 2381 16745 2421 16785 ne
rect 2421 16745 2599 16785
rect 1659 16729 2135 16745
tri 2135 16729 2151 16745 sw
tri 2215 16729 2231 16745 ne
rect 2231 16729 2381 16745
tri 2421 16729 2437 16745 ne
rect 1659 16695 2151 16729
tri 2151 16695 2185 16729 sw
tri 2231 16695 2265 16729 ne
rect 1659 16671 2185 16695
tri 2185 16671 2209 16695 sw
rect 1659 510 2209 16671
rect 2265 12265 2381 16729
tri 2431 12235 2437 12241 se
rect 2437 12235 2599 16745
rect 2649 12265 2765 16953
tri 2809 16945 2817 16953 se
rect 2817 16945 2909 16953
tri 2793 16929 2809 16945 se
rect 2809 16929 2909 16945
rect 2793 16923 2909 16929
rect 2845 16871 2857 16923
rect 2793 16865 2909 16871
rect 2793 16853 2897 16865
tri 2897 16853 2909 16865 nw
rect 2793 16825 2869 16853
tri 2869 16825 2897 16853 nw
tri 2909 16825 2937 16853 se
rect 2937 16825 3283 16953
tri 2389 12193 2431 12235 se
rect 2431 12193 2599 12235
tri 2599 12193 2641 12235 sw
rect 1659 458 1773 510
rect 1825 458 1837 510
rect 1889 458 1901 510
rect 1953 458 2209 510
rect 1659 341 2209 458
tri 2265 12069 2389 12193 se
rect 2389 12069 2641 12193
tri 2641 12069 2765 12193 sw
rect 2265 9739 2765 12069
rect 2265 9687 2297 9739
rect 2349 9687 2361 9739
rect 2413 9687 2425 9739
rect 2477 9687 2489 9739
rect 2541 9687 2553 9739
rect 2605 9687 2617 9739
rect 2669 9687 2681 9739
rect 2733 9687 2765 9739
rect 2265 341 2765 9687
rect 2793 341 2845 16825
tri 2845 16801 2869 16825 nw
tri 2901 16817 2909 16825 se
rect 2909 16817 3283 16825
rect 2901 510 3283 16817
rect 2901 458 3097 510
rect 3149 458 3161 510
rect 3213 458 3225 510
rect 3277 458 3283 510
rect 2901 341 3283 458
rect 3339 341 3391 16845
rect 3419 16748 3484 16953
rect 3512 16821 3628 16953
rect 3656 16861 3721 16953
rect 3749 16900 3801 16953
tri 3749 16888 3761 16900 ne
rect 3761 16888 3801 16900
tri 3801 16888 3835 16922 sw
rect 3857 16907 4239 16953
tri 3857 16888 3876 16907 ne
rect 3876 16888 4239 16907
tri 3656 16849 3668 16861 ne
rect 3668 16860 3721 16861
tri 3721 16860 3749 16888 sw
tri 3761 16881 3768 16888 ne
rect 3768 16881 3835 16888
tri 3835 16881 3842 16888 sw
tri 3876 16881 3883 16888 ne
rect 3883 16881 4239 16888
tri 3768 16860 3789 16881 ne
rect 3789 16866 3842 16881
tri 3842 16866 3857 16881 sw
tri 3883 16866 3898 16881 ne
rect 3898 16866 4239 16881
rect 3789 16860 3857 16866
rect 3668 16849 3749 16860
tri 3749 16849 3760 16860 sw
tri 3789 16849 3800 16860 ne
rect 3800 16849 3857 16860
tri 3857 16849 3874 16866 sw
tri 3898 16849 3915 16866 ne
rect 3915 16849 4239 16866
tri 3628 16821 3656 16849 sw
tri 3668 16821 3696 16849 ne
rect 3696 16848 3760 16849
tri 3760 16848 3761 16849 sw
tri 3800 16848 3801 16849 ne
rect 3801 16848 3874 16849
rect 3696 16821 3761 16848
rect 3512 16817 3656 16821
tri 3656 16817 3660 16821 sw
tri 3696 16819 3698 16821 ne
rect 3698 16819 3761 16821
tri 3761 16819 3790 16848 sw
tri 3801 16819 3830 16848 ne
rect 3830 16819 3874 16848
tri 3874 16819 3904 16849 sw
tri 3915 16819 3945 16849 ne
rect 3945 16819 4239 16849
tri 3698 16817 3700 16819 ne
rect 3700 16817 3790 16819
tri 3790 16817 3792 16819 sw
tri 3830 16817 3832 16819 ne
rect 3832 16817 3904 16819
tri 3904 16817 3906 16819 sw
tri 3945 16817 3947 16819 ne
rect 3947 16817 4239 16819
rect 3512 16800 3660 16817
tri 3512 16788 3524 16800 ne
rect 3524 16796 3660 16800
tri 3660 16796 3681 16817 sw
tri 3700 16796 3721 16817 ne
rect 3721 16808 3792 16817
tri 3792 16808 3801 16817 sw
tri 3832 16808 3841 16817 ne
rect 3841 16808 3906 16817
rect 3721 16807 3801 16808
tri 3801 16807 3802 16808 sw
tri 3841 16807 3842 16808 ne
rect 3842 16807 3906 16808
tri 3906 16807 3916 16817 sw
tri 3947 16807 3957 16817 ne
rect 3957 16807 4239 16817
rect 3721 16796 3802 16807
rect 3524 16788 3681 16796
tri 3484 16748 3524 16788 sw
tri 3524 16748 3564 16788 ne
rect 3564 16756 3681 16788
tri 3681 16756 3721 16796 sw
tri 3721 16756 3761 16796 ne
rect 3761 16767 3802 16796
tri 3802 16767 3842 16807 sw
tri 3842 16792 3857 16807 ne
rect 3857 16792 3916 16807
tri 3857 16767 3882 16792 ne
rect 3882 16774 3916 16792
tri 3916 16774 3949 16807 sw
tri 3957 16774 3990 16807 ne
rect 3990 16774 4239 16807
rect 3882 16767 3949 16774
rect 3761 16756 3842 16767
rect 3564 16748 3721 16756
rect 3419 16723 3524 16748
tri 3524 16723 3549 16748 sw
tri 3564 16723 3589 16748 ne
rect 3589 16727 3721 16748
tri 3721 16727 3750 16756 sw
tri 3761 16727 3790 16756 ne
rect 3790 16752 3842 16756
tri 3842 16752 3857 16767 sw
tri 3882 16752 3897 16767 ne
rect 3897 16752 3949 16767
rect 3790 16733 3857 16752
tri 3857 16733 3876 16752 sw
tri 3897 16733 3916 16752 ne
rect 3916 16733 3949 16752
tri 3949 16733 3990 16774 sw
rect 3790 16727 3876 16733
tri 3876 16727 3882 16733 sw
rect 3589 16723 3750 16727
rect 3419 16716 3549 16723
tri 3549 16716 3556 16723 sw
tri 3589 16716 3596 16723 ne
rect 3596 16716 3750 16723
tri 3750 16716 3761 16727 sw
rect 3419 16684 3556 16716
tri 3556 16684 3588 16716 sw
tri 3596 16684 3628 16716 ne
rect 3628 16684 3761 16716
tri 3790 16700 3817 16727 ne
rect 3419 16683 3588 16684
tri 3588 16683 3589 16684 sw
rect 3419 12235 3589 16683
tri 3628 16667 3645 16684 ne
rect 3645 12265 3761 16684
tri 3589 12235 3595 12241 sw
tri 3811 12235 3817 12241 se
rect 3817 12235 3882 16727
tri 3916 16718 3931 16733 ne
rect 3931 16718 3990 16733
tri 3990 16718 4046 16774 ne
tri 3931 16711 3938 16718 ne
rect 3419 12216 3595 12235
tri 3595 12216 3614 12235 sw
tri 3792 12216 3811 12235 se
rect 3811 12216 3882 12235
rect 3419 510 3882 12216
rect 3419 458 3508 510
rect 3560 458 3572 510
rect 3624 458 3636 510
rect 3688 458 3882 510
rect 3419 341 3882 458
rect 3938 341 3990 16718
rect 4046 16485 4239 16774
rect 4295 16648 4347 16953
rect 4295 16584 4347 16596
rect 4295 16526 4347 16532
tri 4239 16485 4264 16510 sw
tri 4378 16485 4403 16510 se
rect 4403 16485 4536 16953
rect 4046 12371 4536 16485
rect 4046 11952 4305 12371
tri 4305 12339 4337 12371 nw
tri 4437 12339 4469 12371 ne
rect 4361 12309 4413 12315
rect 4361 12245 4413 12257
rect 4361 11987 4413 12193
rect 4469 12068 4536 12371
rect 4592 12265 4708 16953
tri 4536 12068 4708 12240 sw
rect 4469 12033 4708 12068
tri 4469 12009 4493 12033 ne
rect 4493 12009 4708 12033
tri 4361 11963 4385 11987 ne
rect 4385 11976 4413 11987
tri 4413 11976 4446 12009 sw
tri 4493 11976 4526 12009 ne
rect 4385 11963 4446 11976
tri 4305 11952 4316 11963 sw
tri 4385 11952 4396 11963 ne
rect 4396 11952 4446 11963
tri 4446 11952 4470 11976 sw
rect 4046 11946 4316 11952
tri 4316 11946 4322 11952 sw
tri 4396 11946 4402 11952 ne
rect 4402 11946 4473 11952
rect 4046 11935 4322 11946
tri 4322 11935 4333 11946 sw
tri 4402 11935 4413 11946 ne
rect 4413 11935 4421 11946
rect 4046 11927 4333 11935
tri 4333 11927 4341 11935 sw
tri 4413 11927 4421 11935 ne
rect 4046 11906 4341 11927
tri 4341 11906 4362 11927 sw
rect 4046 11768 4362 11906
rect 4421 11882 4473 11894
rect 4421 11824 4473 11830
tri 4362 11768 4394 11800 sw
tri 4494 11768 4526 11800 se
rect 4526 11768 4708 12009
rect 4046 510 4708 11768
rect 4046 458 4585 510
rect 4637 458 4649 510
rect 4701 458 4708 510
rect 4046 341 4708 458
rect 4764 9739 4914 16953
rect 4764 9687 4781 9739
rect 4833 9687 4845 9739
rect 4897 9687 4914 9739
rect 4764 341 4914 9687
rect 4973 15224 5241 15252
rect 4973 15218 5235 15224
tri 5235 15218 5241 15224 nw
rect 5297 15218 5565 15252
rect 4973 15166 5158 15218
rect 5210 15166 5216 15218
tri 5216 15199 5235 15218 nw
rect 4973 15154 5216 15166
rect 4973 15102 5158 15154
rect 5210 15130 5216 15154
rect 5297 15166 5507 15218
rect 5559 15166 5565 15218
rect 5297 15154 5565 15166
tri 5216 15130 5217 15131 sw
rect 5210 15111 5217 15130
tri 5217 15111 5236 15130 sw
tri 5278 15111 5297 15130 se
rect 5297 15111 5507 15154
rect 5210 15102 5507 15111
rect 5559 15102 5565 15154
rect 4973 10624 5565 15102
rect 4973 9378 5241 10624
tri 5241 10592 5273 10624 nw
tri 5385 10592 5417 10624 ne
rect 5297 10516 5303 10568
rect 5355 10516 5361 10568
rect 5297 10504 5361 10516
rect 5297 10452 5303 10504
rect 5355 10452 5361 10504
rect 5297 9550 5361 10452
rect 5297 9498 5303 9550
rect 5355 9498 5361 9550
rect 5297 9486 5361 9498
rect 5297 9434 5303 9486
rect 5355 9434 5361 9486
tri 5241 9378 5273 9410 sw
tri 5385 9378 5417 9410 se
rect 5417 9378 5565 10624
rect 5621 10510 5889 15279
rect 5621 10458 5627 10510
rect 5679 10458 5695 10510
rect 5747 10458 5763 10510
rect 5815 10458 5831 10510
rect 5883 10458 5889 10510
rect 5945 15273 6099 15279
rect 5945 15093 5961 15273
rect 6077 15093 6099 15273
rect 6269 15273 6414 15279
rect 5945 14824 6099 15093
rect 6161 14940 6213 15252
rect 6161 14876 6213 14888
tri 6099 14824 6113 14838 sw
rect 5945 14818 6113 14824
tri 6113 14818 6119 14824 sw
rect 6161 14818 6213 14824
rect 5945 14724 6119 14818
tri 6119 14724 6213 14818 sw
rect 5945 14666 6213 14724
rect 5945 14614 6155 14666
rect 6207 14614 6213 14666
rect 5945 14602 6213 14614
rect 5945 14550 6155 14602
rect 6207 14550 6213 14602
rect 5945 10387 6213 14550
rect 5945 10335 6155 10387
rect 6207 10335 6213 10387
rect 5945 10323 6213 10335
rect 5945 10271 6155 10323
rect 6207 10271 6213 10323
rect 4973 510 5565 9378
rect 4973 458 5443 510
rect 5495 458 5507 510
rect 5559 458 5565 510
rect 4973 393 5565 458
rect 4973 341 5513 393
tri 5513 341 5565 393 nw
rect 5621 341 5889 10142
rect 5945 341 6213 10271
rect 6269 15093 6283 15273
rect 6399 15093 6414 15273
rect 6269 341 6414 15093
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 2631 0 1 9913
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 603 0 1 9773
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 0 1 2576 1 0 9604
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform 0 1 548 1 0 9604
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform 0 -1 4488 1 0 9604
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 0 -1 2460 1 0 9604
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform 1 0 5332 0 -1 13876
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 6036 0 -1 14661
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 5892 0 -1 14661
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 5756 0 -1 14661
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 5612 0 -1 14661
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform 1 0 6172 0 -1 14660
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1707688321
transform 1 0 5192 0 -1 14743
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1707688321
transform 1 0 5476 0 -1 13876
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1707688321
transform 1 0 5472 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1707688321
transform 1 0 5332 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1707688321
transform 1 0 5192 0 1 10193
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1707688321
transform 1 0 2405 0 1 9913
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1707688321
transform 1 0 4433 0 1 9930
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1707688321
transform 1 0 5616 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_20
timestamp 1707688321
transform 1 0 5752 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_21
timestamp 1707688321
transform 1 0 5896 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_22
timestamp 1707688321
transform 1 0 6032 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_23
timestamp 1707688321
transform 1 0 6172 0 1 10275
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 1155 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 1155 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 2867 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 5099 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 5555 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 4871 0 1 5033
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 5327 0 1 5033
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 1155 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 2867 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 5099 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 5555 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 5327 0 1 2815
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 5555 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 5099 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform -1 0 4871 0 1 7253
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform -1 0 2867 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform -1 0 4983 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform -1 0 3039 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform -1 0 594 0 -1 17195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform -1 0 318 0 -1 17195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform -1 0 942 0 -1 17195
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 0 -1 438 1 0 16729
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 5279 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 4421 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 3746 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 2011 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 1055 0 -1 501
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 1 0 1905 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 1 0 3881 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1707688321
transform 1 0 4537 0 1 5032
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1707688321
transform 1 0 866 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1707688321
transform 1 0 1097 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1707688321
transform 1 0 1333 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1707688321
transform 1 0 1569 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1707688321
transform 1 0 1805 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1707688321
transform 1 0 2041 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1707688321
transform 1 0 4064 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1707688321
transform 1 0 3833 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1707688321
transform 1 0 3597 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1707688321
transform 1 0 3361 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1707688321
transform 1 0 3125 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1707688321
transform 1 0 2889 0 1 11971
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1707688321
transform 1 0 1905 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1707688321
transform 1 0 3881 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1707688321
transform 1 0 4537 0 1 2813
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1707688321
transform 1 0 4765 0 1 2814
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1707688321
transform 1 0 5221 0 1 7253
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_47
timestamp 1707688321
transform 1 0 4537 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_48
timestamp 1707688321
transform 1 0 3881 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_49
timestamp 1707688321
transform 1 0 1905 0 1 7252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_50
timestamp 1707688321
transform 1 0 261 0 1 16874
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 1 0 5047 0 -1 591
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 1 0 5413 0 -1 676
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 1 0 4957 0 -1 676
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 1 0 4501 0 -1 676
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 1 0 2429 0 1 12114
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 1 0 5413 0 1 9425
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 1 0 4957 0 1 9425
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 1 0 4501 0 1 9425
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform -1 0 5768 0 -1 591
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1707688321
transform 1 0 5113 0 -1 9544
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_2
timestamp 1707688321
transform 1 0 4658 0 -1 9544
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_3
timestamp 1707688321
transform 1 0 179 0 1 12114
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform 1 0 1209 0 -1 591
box -12 -6 766 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1707688321
transform -1 0 3083 0 1 9425
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1707688321
transform -1 0 4203 0 1 9425
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_2
timestamp 1707688321
transform -1 0 3083 0 -1 676
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_3
timestamp 1707688321
transform -1 0 4203 0 -1 676
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_4
timestamp 1707688321
transform 0 -1 5683 1 0 15114
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_5
timestamp 1707688321
transform 1 0 1689 0 -1 676
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_6
timestamp 1707688321
transform 1 0 833 0 -1 676
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_7
timestamp 1707688321
transform 1 0 1689 0 1 9425
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_8
timestamp 1707688321
transform 1 0 833 0 1 9425
box -12 -6 550 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform -1 0 3180 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1707688321
transform -1 0 1547 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1707688321
transform -1 0 4092 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_3
timestamp 1707688321
transform -1 0 2403 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_4
timestamp 1707688321
transform -1 0 3259 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_5
timestamp 1707688321
transform -1 0 4379 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_6
timestamp 1707688321
transform -1 0 1547 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_7
timestamp 1707688321
transform -1 0 2403 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_8
timestamp 1707688321
transform -1 0 3259 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_9
timestamp 1707688321
transform -1 0 4379 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_10
timestamp 1707688321
transform -1 0 4379 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_11
timestamp 1707688321
transform -1 0 3259 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_12
timestamp 1707688321
transform -1 0 1547 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_13
timestamp 1707688321
transform -1 0 2403 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_14
timestamp 1707688321
transform -1 0 1722 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_15
timestamp 1707688321
transform -1 0 810 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_16
timestamp 1707688321
transform 0 -1 164 1 0 16939
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_17
timestamp 1707688321
transform 1 0 4575 0 -1 591
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_18
timestamp 1707688321
transform 1 0 5608 0 -1 9544
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_19
timestamp 1707688321
transform 1 0 4226 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_20
timestamp 1707688321
transform 1 0 3314 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_21
timestamp 1707688321
transform 1 0 657 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_22
timestamp 1707688321
transform 1 0 1513 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_23
timestamp 1707688321
transform 1 0 2369 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_24
timestamp 1707688321
transform 1 0 3489 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_25
timestamp 1707688321
transform 1 0 657 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_26
timestamp 1707688321
transform 1 0 1513 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_27
timestamp 1707688321
transform 1 0 2369 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_28
timestamp 1707688321
transform 1 0 3489 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_29
timestamp 1707688321
transform 1 0 3489 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_30
timestamp 1707688321
transform 1 0 2369 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_31
timestamp 1707688321
transform 1 0 1513 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_32
timestamp 1707688321
transform 1 0 657 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_33
timestamp 1707688321
transform 1 0 5248 0 1 15698
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_34
timestamp 1707688321
transform 1 0 944 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_35
timestamp 1707688321
transform 1 0 1856 0 1 16744
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 1 0 618 0 -1 591
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1707688321
transform 0 -1 5094 -1 0 15652
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_1
timestamp 1707688321
transform 1 0 3088 0 -1 591
box -12 -6 622 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1707688321
transform 1 0 1189 0 -1 9544
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_1
timestamp 1707688321
transform 1 0 2184 0 -1 591
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_2
timestamp 1707688321
transform 1 0 2045 0 -1 9544
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_3
timestamp 1707688321
transform 1 0 201 0 1 17235
box -12 -6 694 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform 1 0 5142 0 1 10078
box -12 -6 1126 40
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1707688321
transform 0 -1 5566 1 0 15114
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_1
timestamp 1707688321
transform 0 -1 5214 1 0 15114
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_2
timestamp 1707688321
transform 1 0 3907 0 -1 591
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_3
timestamp 1707688321
transform 1 0 546 0 -1 9544
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_4
timestamp 1707688321
transform 1 0 4036 0 -1 9544
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 5747 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform -1 0 5747 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1707688321
transform -1 0 5747 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1707688321
transform 1 0 4345 0 1 5033
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1707688321
transform 1 0 4345 0 1 2814
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1707688321
transform 1 0 4345 0 1 7253
box 0 0 1 1
use L1M1_CDNS_52468879185941  L1M1_CDNS_52468879185941_0
timestamp 1707688321
transform 0 -1 2724 -1 0 11897
box -12 -6 1990 40
use L1M1_CDNS_52468879185941  L1M1_CDNS_52468879185941_1
timestamp 1707688321
transform 0 -1 4374 -1 0 11897
box -12 -6 1990 40
use L1M1_CDNS_52468879185947  L1M1_CDNS_52468879185947_0
timestamp 1707688321
transform 0 1 5060 -1 0 14807
box -12 -6 2566 40
use L1M1_CDNS_52468879185950  L1M1_CDNS_52468879185950_0
timestamp 1707688321
transform 0 -1 386 -1 0 12062
box -12 -6 11638 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1707688321
transform 1 0 2889 0 -1 9544
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_1
timestamp 1707688321
transform 1 0 5132 0 1 14824
box -12 -6 982 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_0
timestamp 1707688321
transform 0 -1 2418 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_1
timestamp 1707688321
transform 0 -1 2652 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_2
timestamp 1707688321
transform 0 -1 2808 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_3
timestamp 1707688321
transform 0 -1 3264 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_4
timestamp 1707688321
transform 0 -1 3720 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_5
timestamp 1707688321
transform 0 -1 4176 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_6
timestamp 1707688321
transform 0 -1 2262 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_7
timestamp 1707688321
transform 0 -1 1806 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_8
timestamp 1707688321
transform 0 -1 1350 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_9
timestamp 1707688321
transform 0 -1 894 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_10
timestamp 1707688321
transform 0 -1 4632 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_11
timestamp 1707688321
transform 0 -1 4788 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_12
timestamp 1707688321
transform 0 -1 438 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_13
timestamp 1707688321
transform 0 -1 282 1 0 15337
box -12 -6 1198 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_0
timestamp 1707688321
transform 1 0 4540 0 -1 9733
box -12 -6 1486 40
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_0
timestamp 1707688321
transform -1 0 2705 0 1 16874
box -12 -6 1918 40
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_1
timestamp 1707688321
transform 0 1 5060 1 0 10119
box -12 -6 1918 40
use L1M1_CDNS_524688791851039  L1M1_CDNS_524688791851039_0
timestamp 1707688321
transform 0 1 131 -1 0 16839
box -12 -6 4654 40
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_0
timestamp 1707688321
transform 0 1 4226 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_1
timestamp 1707688321
transform 0 1 3770 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_2
timestamp 1707688321
transform 0 1 3314 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_3
timestamp 1707688321
transform 0 1 2858 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_4
timestamp 1707688321
transform 0 1 1856 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_5
timestamp 1707688321
transform 0 1 1400 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_6
timestamp 1707688321
transform 0 1 944 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_7
timestamp 1707688321
transform 0 1 488 -1 0 12233
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_8
timestamp 1707688321
transform 0 1 4226 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_9
timestamp 1707688321
transform 0 1 3770 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_10
timestamp 1707688321
transform 0 1 3314 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_11
timestamp 1707688321
transform 0 1 2858 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_12
timestamp 1707688321
transform 0 1 1856 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_13
timestamp 1707688321
transform 0 1 1400 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_14
timestamp 1707688321
transform 0 1 944 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_15
timestamp 1707688321
transform 0 1 488 1 0 13729
box 0 0 1 1
use L1M1_CDNS_524688791851095  L1M1_CDNS_524688791851095_0
timestamp 1707688321
transform 0 1 3357 1 0 654
box -12 -6 8542 40
use L1M1_CDNS_524688791851096  L1M1_CDNS_524688791851096_0
timestamp 1707688321
transform 0 -1 574 1 0 626
box -12 -6 8470 40
use L1M1_CDNS_524688791851096  L1M1_CDNS_524688791851096_1
timestamp 1707688321
transform 0 -1 5864 1 0 626
box -12 -6 8470 40
use L1M1_CDNS_524688791851097  L1M1_CDNS_524688791851097_0
timestamp 1707688321
transform -1 0 4816 0 1 16874
box -12 -6 1774 40
use L1M1_CDNS_524688791851098  L1M1_CDNS_524688791851098_0
timestamp 1707688321
transform 0 -1 2571 1 0 12241
box -12 -6 4294 112
use L1M1_CDNS_524688791851099  L1M1_CDNS_524688791851099_0
timestamp 1707688321
transform -1 0 2313 0 -1 9733
box -12 -6 1630 40
use L1M1_CDNS_524688791851099  L1M1_CDNS_524688791851099_1
timestamp 1707688321
transform 1 0 2723 0 -1 9733
box -12 -6 1630 40
use L1M1_CDNS_524688791851100  L1M1_CDNS_524688791851100_0
timestamp 1707688321
transform 0 1 6304 1 0 10084
box -12 -6 4726 40
use L1M1_CDNS_524688791851101  L1M1_CDNS_524688791851101_0
timestamp 1707688321
transform 1 0 449 0 -1 402
box -12 -6 5518 40
use L1M1_CDNS_524688791851102  L1M1_CDNS_524688791851102_0
timestamp 1707688321
transform 0 -1 6053 1 0 424
box -12 -6 8974 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_0
timestamp 1707688321
transform 0 -1 2346 -1 0 11897
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_1
timestamp 1707688321
transform 0 -1 696 -1 0 11897
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_2
timestamp 1707688321
transform 0 -1 4563 -1 0 11969
box -12 -6 2062 40
use L1M1_CDNS_524688791851103  L1M1_CDNS_524688791851103_3
timestamp 1707688321
transform 0 -1 4685 -1 0 11969
box -12 -6 2062 40
use L1M1_CDNS_524688791851104  L1M1_CDNS_524688791851104_0
timestamp 1707688321
transform 0 -1 4905 -1 0 16857
box -12 -6 4582 40
use L1M1_CDNS_524688791851105  L1M1_CDNS_524688791851105_0
timestamp 1707688321
transform 0 -1 2535 -1 0 12042
box -12 -6 2134 40
use L1M1_CDNS_524688791851106  L1M1_CDNS_524688791851106_0
timestamp 1707688321
transform 0 -1 507 -1 0 12062
box -12 -6 2350 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 4347 -1 0 16654
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 1 4361 -1 0 12315
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 4903 0 1 9687
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform -1 0 -114 0 -1 17275
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 4421 1 0 11824
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 -1 6213 1 0 14818
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 1 0 5437 0 1 458
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 1 0 4579 0 1 458
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 1 6283 1 0 15087
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1707688321
transform 0 1 5961 1 0 15087
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 0 1 207 1 0 16945
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 0 1 -29 1 0 17073
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform -1 0 3283 0 1 458
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1707688321
transform 1 0 3502 0 1 458
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1707688321
transform 1 0 1767 0 1 458
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1707688321
transform 1 0 811 0 1 458
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform -1 0 2560 0 1 16862
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 2793 -1 0 16929
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform -1 0 5361 0 1 10452
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform -1 0 5361 0 1 9434
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform -1 0 6213 0 1 14550
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1707688321
transform -1 0 6213 0 1 10271
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_5
timestamp 1707688321
transform 1 0 5152 0 1 15102
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_6
timestamp 1707688321
transform 1 0 5501 0 1 15102
box 0 0 1 1
use M1M2_CDNS_52468879185965  M1M2_CDNS_52468879185965_0
timestamp 1707688321
transform 0 -1 2544 -1 0 12116
box 0 0 2176 52
use M1M2_CDNS_524688791851020  M1M2_CDNS_524688791851020_0
timestamp 1707688321
transform 0 -1 4816 -1 0 11981
box 0 0 1984 52
use M1M2_CDNS_524688791851033  M1M2_CDNS_524688791851033_0
timestamp 1707688321
transform 0 1 4862 -1 0 16873
box 0 0 4672 52
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1707688321
transform 0 -1 1481 1 0 16942
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_1
timestamp 1707688321
transform 0 -1 2201 1 0 16942
box 0 0 256 180
use M1M2_CDNS_524688791851107  M1M2_CDNS_524688791851107_0
timestamp 1707688321
transform 0 1 1333 -1 0 15183
box 0 0 1344 116
use M1M2_CDNS_524688791851107  M1M2_CDNS_524688791851107_1
timestamp 1707688321
transform 0 1 1333 -1 0 13653
box 0 0 1344 116
use M1M2_CDNS_524688791851107  M1M2_CDNS_524688791851107_2
timestamp 1707688321
transform 0 1 3645 -1 0 13653
box 0 0 1344 116
use M1M2_CDNS_524688791851107  M1M2_CDNS_524688791851107_3
timestamp 1707688321
transform 0 1 3645 -1 0 15183
box 0 0 1344 116
use M1M2_CDNS_524688791851108  M1M2_CDNS_524688791851108_0
timestamp 1707688321
transform 0 -1 174 -1 0 16873
box 0 0 4736 52
use M1M2_CDNS_524688791851109  M1M2_CDNS_524688791851109_0
timestamp 1707688321
transform 0 1 122 -1 0 12077
box 0 0 11712 52
use M1M2_CDNS_524688791851110  M1M2_CDNS_524688791851110_0
timestamp 1707688321
transform 0 1 4592 1 0 12265
box 0 0 4288 116
use M1M2_CDNS_524688791851110  M1M2_CDNS_524688791851110_1
timestamp 1707688321
transform 0 1 2649 1 0 12265
box 0 0 4288 116
use M1M2_CDNS_524688791851110  M1M2_CDNS_524688791851110_2
timestamp 1707688321
transform 0 1 285 1 0 12265
box 0 0 4288 116
use M1M2_CDNS_524688791851110  M1M2_CDNS_524688791851110_3
timestamp 1707688321
transform 0 1 2265 1 0 12265
box 0 0 4288 116
use M1M2_CDNS_524688791851111  M1M2_CDNS_524688791851111_0
timestamp 1707688321
transform 0 1 3645 1 0 15369
box 0 0 1152 116
use M1M2_CDNS_524688791851111  M1M2_CDNS_524688791851111_1
timestamp 1707688321
transform 0 1 1333 1 0 15369
box 0 0 1152 116
use M1M2_CDNS_524688791851112  M1M2_CDNS_524688791851112_0
timestamp 1707688321
transform 0 1 2460 1 0 12137
box 0 0 4416 116
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_0
timestamp 1707688321
transform 1 0 2291 0 1 9687
box 0 0 1 1
use M1M2_CDNS_524688791851114  M1M2_CDNS_524688791851114_0
timestamp 1707688321
transform 0 -1 5103 1 0 10117
box 0 0 1920 52
use M1M2_CDNS_524688791851115  M1M2_CDNS_524688791851115_0
timestamp 1707688321
transform 0 -1 5103 -1 0 14864
box 0 0 2624 52
use nDFres_CDNS_524688791851138  nDFres_CDNS_524688791851138_0
timestamp 1707688321
transform 0 -1 5389 1 0 10297
box -68 -26 3543 106
use nDFres_CDNS_524688791851138  nDFres_CDNS_524688791851138_1
timestamp 1707688321
transform 0 -1 5529 1 0 10297
box -68 -26 3543 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_0
timestamp 1707688321
transform 0 -1 5249 -1 0 14639
box -68 -26 4410 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_1
timestamp 1707688321
transform 0 -1 5669 -1 0 14639
box -68 -26 4410 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_2
timestamp 1707688321
transform 0 -1 5809 -1 0 14639
box -68 -26 4410 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_3
timestamp 1707688321
transform 0 -1 5949 -1 0 14639
box -68 -26 4410 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_4
timestamp 1707688321
transform 0 -1 6089 -1 0 14639
box -68 -26 4410 106
use nDFres_CDNS_524688791851139  nDFres_CDNS_524688791851139_5
timestamp 1707688321
transform 0 -1 6229 -1 0 14639
box -68 -26 4410 106
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_0
timestamp 1707688321
transform 1 0 2414 0 1 7377
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_1
timestamp 1707688321
transform 1 0 2414 0 1 2938
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_2
timestamp 1707688321
transform 1 0 3534 0 1 5163
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_3
timestamp 1707688321
transform 1 0 2414 0 1 5163
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_4
timestamp 1707688321
transform 1 0 2414 0 1 724
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_5
timestamp 1707688321
transform 1 0 3534 0 1 724
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_6
timestamp 1707688321
transform 1 0 3534 0 1 2938
box -79 -26 879 2026
use nfet_CDNS_524688791851116  nfet_CDNS_524688791851116_7
timestamp 1707688321
transform 1 0 3534 0 1 7377
box -79 -26 879 2026
use nfet_CDNS_524688791851118  nfet_CDNS_524688791851118_0
timestamp 1707688321
transform 1 0 4390 0 1 724
box -79 -26 1391 2026
use nfet_CDNS_524688791851118  nfet_CDNS_524688791851118_1
timestamp 1707688321
transform 1 0 4390 0 1 2938
box -79 -26 1391 2026
use nfet_CDNS_524688791851118  nfet_CDNS_524688791851118_2
timestamp 1707688321
transform 1 0 4390 0 1 7377
box -79 -26 1391 2026
use nfet_CDNS_524688791851118  nfet_CDNS_524688791851118_3
timestamp 1707688321
transform 1 0 4390 0 1 5163
box -79 -26 1391 2026
use nfet_CDNS_524688791851119  nfet_CDNS_524688791851119_0
timestamp 1707688321
transform 1 0 5225 0 -1 15648
box -82 -26 375 626
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_0
timestamp 1707688321
transform -1 0 1712 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_1
timestamp 1707688321
transform -1 0 1948 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_2
timestamp 1707688321
transform -1 0 2184 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_3
timestamp 1707688321
transform -1 0 1004 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_4
timestamp 1707688321
transform -1 0 1240 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_5
timestamp 1707688321
transform -1 0 1476 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_6
timestamp 1707688321
transform -1 0 3504 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_7
timestamp 1707688321
transform -1 0 3268 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_8
timestamp 1707688321
transform -1 0 3032 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_9
timestamp 1707688321
transform -1 0 4212 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_10
timestamp 1707688321
transform -1 0 3976 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851120  nfet_CDNS_524688791851120_11
timestamp 1707688321
transform -1 0 3740 0 1 9923
box -79 -26 259 2026
use nfet_CDNS_524688791851121  nfet_CDNS_524688791851121_0
timestamp 1707688321
transform -1 0 2358 0 1 5163
box -79 -26 1735 2026
use nfet_CDNS_524688791851121  nfet_CDNS_524688791851121_1
timestamp 1707688321
transform -1 0 2358 0 1 7377
box -79 -26 1735 2026
use nfet_CDNS_524688791851121  nfet_CDNS_524688791851121_2
timestamp 1707688321
transform -1 0 2358 0 1 2938
box -79 -26 1735 2026
use nfet_CDNS_524688791851121  nfet_CDNS_524688791851121_3
timestamp 1707688321
transform -1 0 2358 0 1 724
box -79 -26 1735 2026
use nfet_CDNS_524688791851122  nfet_CDNS_524688791851122_0
timestamp 1707688321
transform 0 -1 12187 -1 0 27471
box -79 -32 879 2032
use nfet_CDNS_524688791851123  nfet_CDNS_524688791851123_0
timestamp 1707688321
transform -1 0 14031 0 -1 32120
box -79 -32 479 2032
use nfet_CDNS_524688791851123  nfet_CDNS_524688791851123_1
timestamp 1707688321
transform -1 0 14031 0 -1 29871
box -79 -32 479 2032
use nfet_CDNS_524688791851123  nfet_CDNS_524688791851123_2
timestamp 1707688321
transform -1 0 14031 0 -1 34372
box -79 -32 479 2032
use nfet_CDNS_524688791851123  nfet_CDNS_524688791851123_3
timestamp 1707688321
transform 1 0 9431 0 -1 33483
box -79 -32 479 2032
use nfet_CDNS_524688791851124  nfet_CDNS_524688791851124_0
timestamp 1707688321
transform -1 0 13575 0 -1 32120
box -79 -32 3447 2032
use nfet_CDNS_524688791851124  nfet_CDNS_524688791851124_1
timestamp 1707688321
transform -1 0 13575 0 -1 29871
box -79 -32 3447 2032
use nfet_CDNS_524688791851124  nfet_CDNS_524688791851124_2
timestamp 1707688321
transform -1 0 13575 0 -1 34372
box -79 -32 3447 2032
use pfet_CDNS_524688791851131  pfet_CDNS_524688791851131_0
timestamp 1707688321
transform -1 0 3675 0 1 12281
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_0
timestamp 1707688321
transform -1 0 3675 0 1 13811
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_1
timestamp 1707688321
transform -1 0 4587 0 1 13811
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_2
timestamp 1707688321
transform -1 0 4587 0 1 12281
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_3
timestamp 1707688321
transform -1 0 1305 0 1 13811
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_4
timestamp 1707688321
transform -1 0 2217 0 1 13811
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_5
timestamp 1707688321
transform -1 0 1305 0 1 12281
box -119 -66 975 1466
use pfet_CDNS_524688791851133  pfet_CDNS_524688791851133_6
timestamp 1707688321
transform -1 0 2217 0 1 12281
box -119 -66 975 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_0
timestamp 1707688321
transform -1 0 2763 0 1 13811
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_1
timestamp 1707688321
transform -1 0 2763 0 1 12281
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_2
timestamp 1707688321
transform -1 0 393 0 1 12281
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_3
timestamp 1707688321
transform -1 0 393 0 1 13811
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_4
timestamp 1707688321
transform 1 0 4643 0 1 12281
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_5
timestamp 1707688321
transform 1 0 4643 0 1 13811
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_6
timestamp 1707688321
transform 1 0 2273 0 1 13811
box -119 -66 219 1466
use pfet_CDNS_524688791851134  pfet_CDNS_524688791851134_7
timestamp 1707688321
transform 1 0 2273 0 1 12281
box -119 -66 219 1466
use pfet_CDNS_524688791851135  pfet_CDNS_524688791851135_0
timestamp 1707688321
transform -1 0 4587 0 1 15341
box -119 -66 975 1466
use pfet_CDNS_524688791851135  pfet_CDNS_524688791851135_1
timestamp 1707688321
transform -1 0 3675 0 1 15341
box -119 -66 975 1466
use pfet_CDNS_524688791851135  pfet_CDNS_524688791851135_2
timestamp 1707688321
transform -1 0 2217 0 1 15341
box -119 -66 975 1466
use pfet_CDNS_524688791851135  pfet_CDNS_524688791851135_3
timestamp 1707688321
transform -1 0 1305 0 1 15341
box -119 -66 975 1466
use pfet_CDNS_524688791851136  pfet_CDNS_524688791851136_0
timestamp 1707688321
transform -1 0 2763 0 1 15341
box -119 -66 219 1466
use pfet_CDNS_524688791851136  pfet_CDNS_524688791851136_1
timestamp 1707688321
transform -1 0 393 0 1 15341
box -119 -66 219 1466
use pfet_CDNS_524688791851136  pfet_CDNS_524688791851136_2
timestamp 1707688321
transform 1 0 4643 0 1 15341
box -119 -66 219 1466
use pfet_CDNS_524688791851136  pfet_CDNS_524688791851136_3
timestamp 1707688321
transform 1 0 2273 0 1 15341
box -119 -66 219 1466
use pfet_CDNS_524688791851137  pfet_CDNS_524688791851137_0
timestamp 1707688321
transform -1 0 861 0 -1 17187
box -119 -66 687 266
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 4777 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 -1 4777 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 -1 4777 -1 0 15309
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 -1 2407 -1 0 15309
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 -1 2407 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 -1 2407 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 1 2629 -1 0 15309
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 1 2629 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 0 1 2629 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1707688321
transform 0 1 259 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1707688321
transform 0 1 259 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1707688321
transform 0 1 259 -1 0 15309
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_12
timestamp 1707688321
transform 0 1 2027 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_13
timestamp 1707688321
transform 0 1 1791 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_14
timestamp 1707688321
transform 0 1 1555 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_15
timestamp 1707688321
transform 0 1 1319 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_16
timestamp 1707688321
transform 0 1 1083 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_17
timestamp 1707688321
transform 0 1 847 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_18
timestamp 1707688321
transform 0 1 2875 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_19
timestamp 1707688321
transform 0 1 3111 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_20
timestamp 1707688321
transform 0 1 3347 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_21
timestamp 1707688321
transform 0 1 3583 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_22
timestamp 1707688321
transform 0 1 3819 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_23
timestamp 1707688321
transform 0 1 4055 -1 0 9891
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_24
timestamp 1707688321
transform 0 1 2629 1 0 16773
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_25
timestamp 1707688321
transform 0 1 236 1 0 16773
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_26
timestamp 1707688321
transform 0 1 847 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_27
timestamp 1707688321
transform 0 1 1083 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_28
timestamp 1707688321
transform 0 1 1319 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_29
timestamp 1707688321
transform 0 1 1555 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_30
timestamp 1707688321
transform 0 1 1791 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_31
timestamp 1707688321
transform 0 1 2027 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_32
timestamp 1707688321
transform 0 1 4055 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_33
timestamp 1707688321
transform 0 1 3819 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_34
timestamp 1707688321
transform 0 1 3583 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_35
timestamp 1707688321
transform 0 1 3347 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_36
timestamp 1707688321
transform 0 1 3111 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_37
timestamp 1707688321
transform 0 1 2875 1 0 11955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_38
timestamp 1707688321
transform 0 -1 4777 1 0 16773
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_39
timestamp 1707688321
transform 0 -1 2407 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 1857 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1707688321
transform 0 1 3833 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1707688321
transform 0 1 4489 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_3
timestamp 1707688321
transform 0 1 1857 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_4
timestamp 1707688321
transform 0 1 3833 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_5
timestamp 1707688321
transform 0 1 4489 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_6
timestamp 1707688321
transform 0 1 4489 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_7
timestamp 1707688321
transform 0 1 3833 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_8
timestamp 1707688321
transform 0 1 1857 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_9
timestamp 1707688321
transform 0 -1 1203 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_10
timestamp 1707688321
transform 0 -1 2915 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_11
timestamp 1707688321
transform 0 -1 5147 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_12
timestamp 1707688321
transform 0 -1 5603 1 0 5016
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_13
timestamp 1707688321
transform 0 -1 1203 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_14
timestamp 1707688321
transform 0 -1 1203 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_15
timestamp 1707688321
transform 0 -1 2915 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_16
timestamp 1707688321
transform 0 -1 5147 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_17
timestamp 1707688321
transform 0 -1 5603 1 0 2797
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_18
timestamp 1707688321
transform 0 -1 5603 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_19
timestamp 1707688321
transform 0 -1 5147 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_20
timestamp 1707688321
transform 0 -1 2915 1 0 7236
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1707688321
transform 0 1 2850 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_1
timestamp 1707688321
transform 0 1 3306 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_2
timestamp 1707688321
transform 0 1 3762 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_3
timestamp 1707688321
transform 0 1 4218 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_4
timestamp 1707688321
transform 0 1 4218 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_5
timestamp 1707688321
transform 0 1 3762 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_6
timestamp 1707688321
transform 0 1 3306 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_7
timestamp 1707688321
transform 0 1 2850 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_8
timestamp 1707688321
transform 0 1 480 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_9
timestamp 1707688321
transform 0 1 936 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_10
timestamp 1707688321
transform 0 1 1392 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_11
timestamp 1707688321
transform 0 1 1848 -1 0 13779
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_12
timestamp 1707688321
transform 0 1 1848 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_13
timestamp 1707688321
transform 0 1 1392 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_14
timestamp 1707688321
transform 0 1 936 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_15
timestamp 1707688321
transform 0 1 480 -1 0 12249
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_16
timestamp 1707688321
transform 0 1 5333 -1 0 692
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_17
timestamp 1707688321
transform 0 1 4877 -1 0 692
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_18
timestamp 1707688321
transform 0 1 4421 -1 0 692
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_19
timestamp 1707688321
transform 0 1 2850 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_20
timestamp 1707688321
transform 0 1 3306 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_21
timestamp 1707688321
transform 0 1 3762 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_22
timestamp 1707688321
transform 0 1 4218 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_23
timestamp 1707688321
transform 0 1 480 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_24
timestamp 1707688321
transform 0 1 936 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_25
timestamp 1707688321
transform 0 1 1392 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_26
timestamp 1707688321
transform 0 1 1848 1 0 16773
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_27
timestamp 1707688321
transform 0 1 5333 1 0 9409
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_28
timestamp 1707688321
transform 0 1 4877 1 0 9409
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_29
timestamp 1707688321
transform 0 1 4421 1 0 9409
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 1 5238 1 0 15680
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1707688321
transform 0 -1 3187 -1 0 692
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1707688321
transform 0 -1 4307 -1 0 692
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_2
timestamp 1707688321
transform 0 1 1585 -1 0 692
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_3
timestamp 1707688321
transform 0 1 729 -1 0 692
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_4
timestamp 1707688321
transform 0 1 729 1 0 9409
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_5
timestamp 1707688321
transform 0 1 1585 1 0 9409
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_6
timestamp 1707688321
transform 0 -1 4307 1 0 9409
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_7
timestamp 1707688321
transform 0 -1 3187 1 0 9409
box 0 0 66 746
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 1 306 -1 0 17285
box 0 0 66 542
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_0
timestamp 1707688321
transform -1 0 4619 0 -1 16784
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_1
timestamp 1707688321
transform -1 0 2249 0 -1 16784
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_2
timestamp 1707688321
transform 0 1 5350 1 0 14974
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_3
timestamp 1707688321
transform 0 -1 900 1 0 15201
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_4
timestamp 1707688321
transform 0 -1 1812 1 0 15201
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_5
timestamp 1707688321
transform 0 -1 3270 1 0 15201
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_6
timestamp 1707688321
transform 0 -1 4182 1 0 15201
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_7
timestamp 1707688321
transform 1 0 2787 0 -1 16784
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_8
timestamp 1707688321
transform 1 0 417 0 -1 16784
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_0
timestamp 1707688321
transform 0 1 5320 -1 0 10321
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_1
timestamp 1707688321
transform 0 1 5740 1 0 10335
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_2
timestamp 1707688321
transform 0 1 6020 1 0 10335
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_3
timestamp 1707688321
transform 0 1 5460 1 0 10335
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851126  sky130_fd_io__refgen_em1o_CDNS_524688791851126_4
timestamp 1707688321
transform 0 1 5320 1 0 14615
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_0
timestamp 1707688321
transform -1 0 4917 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_1
timestamp 1707688321
transform -1 0 3786 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_2
timestamp 1707688321
transform -1 0 2051 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_3
timestamp 1707688321
transform -1 0 1095 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_4
timestamp 1707688321
transform -1 0 11044 0 -1 29965
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_5
timestamp 1707688321
transform -1 0 11044 0 -1 32214
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_6
timestamp 1707688321
transform -1 0 11044 0 -1 34466
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_7
timestamp 1707688321
transform 1 0 10628 0 -1 34466
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_8
timestamp 1707688321
transform 1 0 5345 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_9
timestamp 1707688321
transform 1 0 4487 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_10
timestamp 1707688321
transform 1 0 2999 0 1 458
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_0
timestamp 1707688321
transform -1 0 14070 0 -1 33726
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_1
timestamp 1707688321
transform -1 0 14070 0 -1 29965
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_2
timestamp 1707688321
transform -1 0 14070 0 -1 32214
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851128  sky130_fd_io__refgen_em1s_CDNS_524688791851128_3
timestamp 1707688321
transform -1 0 14070 0 -1 34466
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_0
timestamp 1707688321
transform -1 0 3844 0 1 16738
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_1
timestamp 1707688321
transform -1 0 1474 0 1 16738
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_2
timestamp 1707688321
transform 0 1 3911 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_3
timestamp 1707688321
transform 0 1 2791 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_4
timestamp 1707688321
transform 0 1 1935 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_5
timestamp 1707688321
transform 0 1 1079 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_6
timestamp 1707688321
transform 0 1 5479 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_7
timestamp 1707688321
transform 0 1 5023 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_8
timestamp 1707688321
transform 0 1 4567 1 0 9455
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_9
timestamp 1707688321
transform 0 -1 3270 1 0 13671
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_10
timestamp 1707688321
transform 0 -1 4182 1 0 13671
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_11
timestamp 1707688321
transform 0 -1 4182 1 0 12141
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_12
timestamp 1707688321
transform 0 -1 3270 1 0 12178
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_13
timestamp 1707688321
transform 0 -1 900 1 0 12141
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_14
timestamp 1707688321
transform 0 -1 1812 1 0 12141
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_15
timestamp 1707688321
transform 0 -1 900 1 0 13671
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_16
timestamp 1707688321
transform 0 -1 1812 1 0 13671
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_17
timestamp 1707688321
transform 1 0 3562 0 1 16738
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_18
timestamp 1707688321
transform 1 0 1192 0 1 16738
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_0
timestamp 1707688321
transform 0 1 5740 -1 0 10321
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_1
timestamp 1707688321
transform 0 1 6020 -1 0 10321
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_2
timestamp 1707688321
transform 0 1 5460 -1 0 10321
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_3
timestamp 1707688321
transform 0 1 5880 1 0 14615
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_4
timestamp 1707688321
transform 0 1 5600 1 0 14615
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851130  sky130_fd_io__refgen_em1s_CDNS_524688791851130_5
timestamp 1707688321
transform 0 1 5320 1 0 10335
box 0 0 1 1
<< labels >>
flabel comment s 13385 27673 13385 27673 0 FreeSans 600 180 0 0 condiode
flabel comment s 12530 33374 12530 33374 0 FreeSans 600 180 0 0 mid
flabel comment s 3963 352 3963 352 3 FreeSans 200 90 0 0 vohref
flabel comment s 3362 352 3362 352 3 FreeSans 200 90 0 0 fb
flabel comment s 1139 352 1139 352 3 FreeSans 200 90 0 0 vohref
flabel comment s 730 352 730 352 3 FreeSans 200 90 0 0 fb_vinref
flabel comment s 972 11953 972 11953 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2994 11953 2994 11953 0 FreeSans 1000 0 0 0 condiode
flabel comment s 3772 16949 3772 16949 3 FreeSans 200 270 0 0 vohref
flabel comment s 3362 16949 3362 16949 3 FreeSans 200 270 0 0 fb
flabel comment s 955 9430 955 9430 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2818 348 2818 348 3 FreeSans 200 90 0 0 vreg_en_h_n
flabel comment s 1139 17272 1139 17272 3 FreeSans 200 270 0 0 vohref
flabel comment s 730 17272 730 17272 3 FreeSans 200 270 0 0 fb_vinref
flabel metal1 s 6371 14974 6414 15026 3 FreeSans 200 180 0 0 en_outop_h_n
port 2 nsew
flabel metal1 s 4920 16942 4949 16988 3 FreeSans 200 0 0 0 en_outop_h_n
port 2 nsew
flabel metal1 s 2201 16942 2223 17275 3 FreeSans 200 180 0 0 vcc_virt_i
port 3 nsew
flabel metal1 s 6339 9516 6365 9580 7 FreeSans 200 0 0 0 res_stack
port 4 nsew
flabel metal1 s 6339 9620 6365 9684 7 FreeSans 200 0 0 0 fb_out
port 5 nsew
flabel metal2 s -158 341 -106 362 3 FreeSans 200 90 0 0 en_outop_h
port 6 nsew
flabel metal2 s 6269 341 6414 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s -78 341 229 362 3 FreeSans 200 90 0 0 vcc_io
port 8 nsew
flabel metal2 s 2265 341 2765 362 3 FreeSans 200 90 0 0 vcc_io
port 8 nsew
flabel metal2 s 4046 341 4708 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 3419 341 3882 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 2937 16935 3283 16953 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 1659 341 2209 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1221 341 1603 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 811 341 1057 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 285 341 647 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 4764 341 4914 362 3 FreeSans 200 90 0 0 vcc_io
port 8 nsew
flabel metal2 s 4973 15224 5241 15252 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 5297 15224 5565 15252 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 5945 341 6213 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 6161 15224 6213 15252 3 FreeSans 200 270 0 0 voutref
port 9 nsew
flabel metal2 s 4403 16935 4536 16953 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 3857 16935 4239 16953 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 5621 341 5889 362 3 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 3656 16935 3721 16953 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 3419 16935 3484 16953 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 2901 341 3283 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1659 17242 1993 17282 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 1221 17243 1603 17282 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 811 17242 1057 17282 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 265 17254 647 17282 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 2649 16935 2765 16953 3 FreeSans 200 270 0 0 vcc_virt_o
port 10 nsew
flabel metal2 s 3512 16935 3628 16953 3 FreeSans 200 270 0 0 vcc_virt_o
port 10 nsew
flabel metal2 s 4592 16935 4708 16953 3 FreeSans 200 270 0 0 vcc_virt_o
port 10 nsew
flabel metal2 s 4764 16935 4914 16953 3 FreeSans 200 270 0 0 vcc_io
port 8 nsew
flabel metal2 s 2185 17254 2455 17282 3 FreeSans 200 180 0 0 vcc_io
port 8 nsew
flabel metal2 s -78 17269 151 17282 3 FreeSans 200 270 0 0 vcc_io
port 8 nsew
flabel metal2 s 4295 16935 4347 16953 3 FreeSans 200 270 0 0 pgate
port 11 nsew
flabel metal2 s 6269 15224 6414 15252 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 5945 15224 6099 15252 3 FreeSans 200 270 0 0 vgnd
port 7 nsew
flabel metal2 s 5317 341 5513 362 3 FreeSans 200 90 0 0 vgnd
port 7 nsew
<< properties >>
string GDS_END 79452966
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79070916
string path 228.400 841.175 228.400 779.600 
<< end >>
