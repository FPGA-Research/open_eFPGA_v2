magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect -197 388 197 397
rect -197 -388 -188 388
rect 188 -388 197 388
rect -197 -397 197 -388
<< via2 >>
rect -188 -388 188 388
<< metal3 >>
rect -193 388 193 393
rect -193 -388 -188 388
rect 188 -388 193 388
rect -193 -393 193 -388
<< properties >>
string GDS_END 34485094
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34481762
<< end >>
