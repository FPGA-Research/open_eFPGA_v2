magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 53 953
<< metal1 >>
rect -6 953 59 956
rect -6 0 0 953
rect 53 0 59 953
rect -6 -3 59 0
<< properties >>
string GDS_END 34509344
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34505756
<< end >>
