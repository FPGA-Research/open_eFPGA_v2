magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 8 157 283 203
rect 637 157 827 203
rect 8 67 827 157
rect 29 -17 63 67
rect 285 21 827 67
<< scnmos >>
rect 86 93 116 177
rect 175 93 205 177
rect 363 47 393 131
rect 450 47 480 131
rect 534 47 564 131
rect 618 47 648 131
rect 716 47 746 177
<< scpmoshvt >>
rect 79 410 109 494
rect 363 413 393 497
rect 176 297 206 381
rect 459 297 489 381
rect 531 297 561 381
rect 618 297 648 381
rect 716 297 746 497
<< ndiff >>
rect 34 149 86 177
rect 34 115 42 149
rect 76 115 86 149
rect 34 93 86 115
rect 116 149 175 177
rect 116 115 131 149
rect 165 115 175 149
rect 116 93 175 115
rect 205 149 257 177
rect 205 115 215 149
rect 249 115 257 149
rect 663 131 716 177
rect 205 93 257 115
rect 311 97 363 131
rect 311 63 319 97
rect 353 63 363 97
rect 311 47 363 63
rect 393 111 450 131
rect 393 77 403 111
rect 437 77 450 111
rect 393 47 450 77
rect 480 97 534 131
rect 480 63 490 97
rect 524 63 534 97
rect 480 47 534 63
rect 564 111 618 131
rect 564 77 574 111
rect 608 77 618 111
rect 564 47 618 77
rect 648 97 716 131
rect 648 63 668 97
rect 702 63 716 97
rect 648 47 716 63
rect 746 135 801 177
rect 746 101 756 135
rect 790 101 801 135
rect 746 47 801 101
<< pdiff >>
rect 27 475 79 494
rect 27 441 35 475
rect 69 441 79 475
rect 27 410 79 441
rect 109 475 161 494
rect 109 441 119 475
rect 153 441 161 475
rect 109 410 161 441
rect 311 475 363 497
rect 311 441 319 475
rect 353 441 363 475
rect 311 413 363 441
rect 393 413 444 497
rect 663 485 716 497
rect 663 451 671 485
rect 705 451 716 485
rect 124 381 161 410
rect 124 297 176 381
rect 206 339 262 381
rect 206 305 216 339
rect 250 305 262 339
rect 206 297 262 305
rect 408 381 444 413
rect 663 417 716 451
rect 663 383 671 417
rect 705 383 716 417
rect 663 381 716 383
rect 408 297 459 381
rect 489 297 531 381
rect 561 297 618 381
rect 648 297 716 381
rect 746 454 801 497
rect 746 420 756 454
rect 790 420 801 454
rect 746 386 801 420
rect 746 352 756 386
rect 790 352 801 386
rect 746 297 801 352
<< ndiffc >>
rect 42 115 76 149
rect 131 115 165 149
rect 215 115 249 149
rect 319 63 353 97
rect 403 77 437 111
rect 490 63 524 97
rect 574 77 608 111
rect 668 63 702 97
rect 756 101 790 135
<< pdiffc >>
rect 35 441 69 475
rect 119 441 153 475
rect 319 441 353 475
rect 671 451 705 485
rect 216 305 250 339
rect 671 383 705 417
rect 756 420 790 454
rect 756 352 790 386
<< poly >>
rect 79 494 109 520
rect 363 497 393 523
rect 716 497 746 523
rect 525 484 591 494
rect 525 450 541 484
rect 575 450 591 484
rect 525 440 591 450
rect 79 265 109 410
rect 176 381 206 407
rect 176 265 206 297
rect 363 265 393 413
rect 459 381 489 407
rect 531 381 561 440
rect 618 381 648 407
rect 459 265 489 297
rect 75 249 129 265
rect 75 215 85 249
rect 119 215 129 249
rect 75 199 129 215
rect 173 249 239 265
rect 173 215 189 249
rect 223 215 239 249
rect 173 199 239 215
rect 302 249 393 265
rect 302 215 312 249
rect 346 215 393 249
rect 302 199 393 215
rect 435 249 489 265
rect 435 215 445 249
rect 479 215 489 249
rect 435 199 489 215
rect 86 177 116 199
rect 175 177 205 199
rect 363 131 393 199
rect 450 131 480 199
rect 531 182 561 297
rect 618 265 648 297
rect 716 265 746 297
rect 603 249 657 265
rect 603 215 613 249
rect 647 215 657 249
rect 603 199 657 215
rect 699 249 753 265
rect 699 215 709 249
rect 743 215 753 249
rect 699 199 753 215
rect 531 152 564 182
rect 534 131 564 152
rect 618 131 648 199
rect 716 177 746 199
rect 86 67 116 93
rect 175 67 205 93
rect 363 21 393 47
rect 450 21 480 47
rect 534 21 564 47
rect 618 21 648 47
rect 716 21 746 47
<< polycont >>
rect 541 450 575 484
rect 85 215 119 249
rect 189 215 223 249
rect 312 215 346 249
rect 445 215 479 249
rect 613 215 647 249
rect 709 215 743 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 475 69 491
rect 17 441 35 475
rect 103 475 169 527
rect 496 484 624 491
rect 103 441 119 475
rect 153 441 169 475
rect 302 441 319 475
rect 353 441 451 475
rect 17 407 69 441
rect 17 373 383 407
rect 17 165 51 373
rect 85 249 155 339
rect 198 305 216 339
rect 250 305 315 339
rect 119 215 155 249
rect 85 199 155 215
rect 189 249 247 265
rect 223 215 247 249
rect 189 199 247 215
rect 281 249 315 305
rect 349 317 383 373
rect 417 391 451 441
rect 496 450 541 484
rect 575 450 624 484
rect 496 425 624 450
rect 658 485 714 527
rect 658 451 671 485
rect 705 451 714 485
rect 658 417 714 451
rect 417 357 624 391
rect 658 383 671 417
rect 705 383 714 417
rect 658 367 714 383
rect 756 454 811 493
rect 790 420 811 454
rect 756 386 811 420
rect 590 333 624 357
rect 790 352 811 386
rect 349 283 479 317
rect 590 299 722 333
rect 756 299 811 352
rect 445 249 479 283
rect 688 265 722 299
rect 281 215 312 249
rect 346 215 366 249
rect 281 165 315 215
rect 445 199 479 215
rect 523 249 654 265
rect 523 215 613 249
rect 647 215 654 249
rect 523 199 654 215
rect 688 249 743 265
rect 688 215 709 249
rect 688 199 743 215
rect 688 165 722 199
rect 17 149 80 165
rect 17 115 42 149
rect 76 115 80 149
rect 17 90 80 115
rect 131 149 165 165
rect 131 17 165 115
rect 215 149 315 165
rect 249 131 315 149
rect 403 131 722 165
rect 777 152 811 299
rect 756 135 811 152
rect 215 90 249 115
rect 403 111 437 131
rect 294 63 319 97
rect 353 63 369 97
rect 294 17 369 63
rect 574 111 608 131
rect 403 61 437 77
rect 474 63 490 97
rect 524 63 540 97
rect 474 17 540 63
rect 790 101 811 135
rect 574 61 608 77
rect 642 63 668 97
rect 702 63 718 97
rect 756 83 811 101
rect 642 17 718 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 581 221 615 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 765 357 799 391 0 FreeSans 400 0 0 0 X
port 9 nsew signal output
flabel locali s 581 425 615 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 D_N
port 4 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or4bb_1
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1097624
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1090576
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
