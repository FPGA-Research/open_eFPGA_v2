##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 18:40:22 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 30.2600 ;
  FOREIGN S_term_RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.57085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.201 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.3682 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.804 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 7.9650 29.9300 8.1350 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.229 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 29.9300 7.2150 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.84245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.697 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8026 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.9355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 6.1250 29.9300 6.2950 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.59425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.405 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.0404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.0875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 29.9300 5.3750 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5072 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 29.9300 16.8750 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 29.9300 15.4950 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1464 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.496 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 14.4050 29.9300 14.5750 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.58865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 29.9300 13.6550 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8516 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.14 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.1050 29.9300 12.2750 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.284 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 29.9300 11.3550 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.426 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.682 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 29.9300 10.4350 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.79945 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.117 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.587 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.8205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 29.9300 9.5150 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.546 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 29.9300 25.1550 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.0650 29.9300 24.2350 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.104 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.6850 29.9300 22.8550 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.5076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.4235 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 29.9300 21.9350 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5669 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.22885 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.752 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 29.9300 21.0150 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.159 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.8584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.656 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 29.9300 19.6350 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.6004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 18.5450 29.9300 18.7150 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 29.9300 17.7950 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.0578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 29.9300 41.7150 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.422 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.226 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 40.6250 29.9300 40.7950 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 29.9300 39.8750 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 29.9300 38.9550 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5165 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 37.4050 29.9300 37.5750 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 29.9300 36.6550 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 29.9300 35.7350 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0728 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.246 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 29.9300 34.3550 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.914 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 29.9300 33.4350 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.428 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 29.9300 32.5150 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9352 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.5615 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.404 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.4250 29.9300 31.5950 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.1548 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.296 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 30.0450 29.9300 30.2150 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.406 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 29.9300 29.2950 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.18105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.213 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4053 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.819 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 29.9300 28.3750 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 29.9300 26.9950 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.594 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 29.9300 26.0750 30.2600 ;
    END
  END N4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7732 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.9733 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.393 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 29.9300 45.8550 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.8638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 79.8711 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 44.7650 29.9300 44.9350 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.8333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 29.9300 44.0150 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.3519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.569 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 29.9300 43.0950 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.7997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.5503 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 29.9300 62.8750 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.3267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.1855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 29.9300 61.9550 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 55.9877 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.937 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 29.9300 60.5750 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9041 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.047 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 29.9300 59.6550 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.856 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8953 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.4528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 29.9300 58.7350 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.2827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.16 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 29.9300 57.8150 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.9616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 126.56 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 29.9300 56.4350 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2804 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.284 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 55.3450 29.9300 55.5150 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1582 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.3428 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 54.4250 29.9300 54.5950 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.154 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.2852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 140.494 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 53.0450 29.9300 53.2150 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4328 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.928 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.2525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.072 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 29.9300 52.2950 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4251 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 18.9079 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 103.855 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 51.2050 29.9300 51.3750 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.19 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.9748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 50.2850 29.9300 50.4550 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.10585 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.301 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.0016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.9305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.6752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 48.9050 29.9300 49.0750 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9226 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4588 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.8459 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 29.9300 48.1550 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.72 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.364 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 38.2852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 186.236 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 29.9300 47.2350 30.2600 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9253 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.4555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 74.2028 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 395.597 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 29.9300 79.4350 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.5776 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.8105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.796 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.1494 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.2987 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 78.3450 29.9300 78.5150 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.952 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8664 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.8836 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 29.9300 77.5950 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.934 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7607 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 118.613 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 29.9300 76.6750 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.577 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.4371 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 29.9300 75.2950 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8044 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.904 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.6978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.4654 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 74.2050 29.9300 74.3750 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.0496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.894 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.3745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 130.94 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 73.2850 29.9300 73.4550 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.561925 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.5316 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.776 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 28.0418 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.091 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 29.9300 72.5350 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.775 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.639 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 31.3808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 152.138 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 29.9300 71.1550 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5086 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.425 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1267 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.6101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.0650 29.9300 70.2350 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.06 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1016 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.0597 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 69.1450 29.9300 69.3150 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.513 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 67.7650 29.9300 67.9350 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.57165 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.849 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.848 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.655 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.928 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 29.9300 67.0150 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 89.7701 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 480.17 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.9250 29.9300 66.0950 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6188 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 65.0050 29.9300 65.1750 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.3796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 147.45 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 63.6250 29.9300 63.7950 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.654 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.8774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.4658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 85.5475 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 447.113 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1998 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.588 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.966 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 3.6739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 13.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3852 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.7393 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.8711 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.7712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.344 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.9255 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.1792 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1312 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.312 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.07013 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.5849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6716 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.122 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.12925 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.456 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.7952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 3.01226 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 11.0377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4428 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.449 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.528 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.9494 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.808 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 60.3399 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 326.088 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.314 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.919 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.6918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.16 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 51.1601 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.157 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.636 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 41.35 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 217.327 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.447 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3226 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.328 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 28.6972 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 153.679 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.632 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.2408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.088 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 28.4053 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.296 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.006 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9155 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.796 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0726 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.1101 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.69065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.989 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.50912 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8126 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.956 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.3812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 41.8285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.5094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.601 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.779 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.28396 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 22.3019 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.45 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.089 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.8468 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.32 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 52.7437 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 278.346 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.969 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.6261 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.4277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4895 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.0783 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 131.006 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.677 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 63.4057 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8505 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.6569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.8396 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.064 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 31.528 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 150.796 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 50.9362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 272.434 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.4395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.584 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6646 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 32.194 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 171.302 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.448 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 36.0311 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 172.06 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.861 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.824 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 43.5349 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 224.843 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3379 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.2948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.376 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 56.0682 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 293.069 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5924 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.854 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.2399 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.814 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7347 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.759 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6302 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 58.272 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.365 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.507 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.5818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 89.4708 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 468.635 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.493 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 28.6600 100.2800 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 26.6200 100.2800 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2401 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.87 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.5538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.424 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 24.9200 100.2800 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 22.8800 100.2800 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5625 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 21.1800 100.2800 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3127 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 19.1400 100.2800 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8505 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 17.4400 100.2800 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 15.7400 100.2800 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 13.7000 100.2800 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.4328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 12.0000 100.2800 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6193 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6738 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.064 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 10.3000 100.2800 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 8.2600 100.2800 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4913 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2305 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 6.5600 100.2800 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8806 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.177 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 4.5200 100.2800 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.986 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.704 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 2.8200 100.2800 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.681 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 1.1200 100.2800 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.165 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 27.6250 100.2800 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.812 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 25.9250 100.2800 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.1145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 24.2250 100.2800 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.355 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.6984 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.136 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 22.5250 100.2800 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.0145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.831 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 20.8250 100.2800 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.826 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8144 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.836 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 19.1250 100.2800 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.521 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 17.4250 100.2800 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2042 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.549 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 15.7250 100.2800 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 14.0250 100.2800 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8874 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.044 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.3944 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.935 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 12.3250 100.2800 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 10.6250 100.2800 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.0084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 8.9250 100.2800 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.7095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.81 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 7.2250 100.2800 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7438 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.228 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.4928 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.427 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 5.5250 100.2800 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4828 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.568 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 3.8250 100.2800 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.4385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 2.1250 100.2800 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.1447 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 0.0000 97.8200 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.2453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.274 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.064 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 22.5299 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 119.069 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 0.0000 95.9800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.264 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1876 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 64.5978 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 346.082 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 72.1447 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 0.0000 94.6000 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8675 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.3035 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.8145 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 0.0000 93.6800 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9814 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.7799 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 0.0000 92.7600 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7715 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.9852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.7987 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 0.0000 91.8400 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2298 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 23.6802 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 127.189 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 0.0000 91.3800 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6395 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.8871 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 99.3082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 0.0000 90.4600 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.7965 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.597 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.0881 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 0.0000 88.6200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.3774 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5455 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.6695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.2201 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 0.0000 87.2400 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.7991 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.2925 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 86.1800 0.0000 86.3200 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.327 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9774 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.2217 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.327 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 85.2600 0.0000 85.4000 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0028 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 54.8868 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 0.0000 84.9400 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0122 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.5024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.424 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 22.8267 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 126.299 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.8800 0.0000 84.0200 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.352 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 26.1925 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.145 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 0.0000 83.1000 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4116 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.9308 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 0.0000 82.6400 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9608 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 29.7750 97.8200 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7934 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.806 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.9488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.864 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 29.7750 96.9000 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4766 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.222 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.417 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.7768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.28 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 29.7750 95.9800 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7782 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.612 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.9216 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.856 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 29.7750 95.0600 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 29.7750 94.6000 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 29.7750 93.6800 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 29.7750 92.7600 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.4255 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 29.7750 91.8400 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.4615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 29.7750 91.3800 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 29.7750 90.4600 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 29.7750 89.5400 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 29.7750 88.6200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 29.7750 88.1600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.5600 29.7750 87.7000 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.192 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.182 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 28.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.2856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.464 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 29.7750 86.7800 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.05 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.024 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 29.7750 85.8600 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9019 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 29.7750 84.9400 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8519 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0335 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.8800 29.7750 84.0200 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5014 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.346 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.573 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.856 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.4478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.192 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 29.7750 83.1000 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7838 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.64 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 29.7750 82.6400 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 94.7200 6.0700 ;
        RECT 5.5600 23.0000 94.7200 25.0000 ;
        RECT 92.7200 15.0600 94.7200 15.5400 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 92.7200 9.6200 94.7200 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 92.7200 20.5000 94.7200 20.9800 ;
      LAYER met4 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 92.7200 4.0700 94.7200 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 97.7200 3.0700 ;
        RECT 2.5600 26.0000 97.7200 28.0000 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 95.7200 12.3400 97.7200 12.8200 ;
        RECT 95.7200 6.9000 97.7200 7.3800 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 95.7200 17.7800 97.7200 18.2600 ;
      LAYER met4 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 95.7200 1.0700 97.7200 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 79.6050 29.7600 100.2800 30.2600 ;
      RECT 78.6850 29.7600 79.0950 30.2600 ;
      RECT 77.7650 29.7600 78.1750 30.2600 ;
      RECT 76.8450 29.7600 77.2550 30.2600 ;
      RECT 75.4650 29.7600 76.3350 30.2600 ;
      RECT 74.5450 29.7600 74.9550 30.2600 ;
      RECT 73.6250 29.7600 74.0350 30.2600 ;
      RECT 72.7050 29.7600 73.1150 30.2600 ;
      RECT 71.3250 29.7600 72.1950 30.2600 ;
      RECT 70.4050 29.7600 70.8150 30.2600 ;
      RECT 69.4850 29.7600 69.8950 30.2600 ;
      RECT 68.1050 29.7600 68.9750 30.2600 ;
      RECT 67.1850 29.7600 67.5950 30.2600 ;
      RECT 66.2650 29.7600 66.6750 30.2600 ;
      RECT 65.3450 29.7600 65.7550 30.2600 ;
      RECT 63.9650 29.7600 64.8350 30.2600 ;
      RECT 63.0450 29.7600 63.4550 30.2600 ;
      RECT 62.1250 29.7600 62.5350 30.2600 ;
      RECT 60.7450 29.7600 61.6150 30.2600 ;
      RECT 59.8250 29.7600 60.2350 30.2600 ;
      RECT 58.9050 29.7600 59.3150 30.2600 ;
      RECT 57.9850 29.7600 58.3950 30.2600 ;
      RECT 56.6050 29.7600 57.4750 30.2600 ;
      RECT 55.6850 29.7600 56.0950 30.2600 ;
      RECT 54.7650 29.7600 55.1750 30.2600 ;
      RECT 53.3850 29.7600 54.2550 30.2600 ;
      RECT 52.4650 29.7600 52.8750 30.2600 ;
      RECT 51.5450 29.7600 51.9550 30.2600 ;
      RECT 50.6250 29.7600 51.0350 30.2600 ;
      RECT 49.2450 29.7600 50.1150 30.2600 ;
      RECT 48.3250 29.7600 48.7350 30.2600 ;
      RECT 47.4050 29.7600 47.8150 30.2600 ;
      RECT 46.0250 29.7600 46.8950 30.2600 ;
      RECT 45.1050 29.7600 45.5150 30.2600 ;
      RECT 44.1850 29.7600 44.5950 30.2600 ;
      RECT 43.2650 29.7600 43.6750 30.2600 ;
      RECT 41.8850 29.7600 42.7550 30.2600 ;
      RECT 40.9650 29.7600 41.3750 30.2600 ;
      RECT 40.0450 29.7600 40.4550 30.2600 ;
      RECT 39.1250 29.7600 39.5350 30.2600 ;
      RECT 37.7450 29.7600 38.6150 30.2600 ;
      RECT 36.8250 29.7600 37.2350 30.2600 ;
      RECT 35.9050 29.7600 36.3150 30.2600 ;
      RECT 34.5250 29.7600 35.3950 30.2600 ;
      RECT 33.6050 29.7600 34.0150 30.2600 ;
      RECT 32.6850 29.7600 33.0950 30.2600 ;
      RECT 31.7650 29.7600 32.1750 30.2600 ;
      RECT 30.3850 29.7600 31.2550 30.2600 ;
      RECT 29.4650 29.7600 29.8750 30.2600 ;
      RECT 28.5450 29.7600 28.9550 30.2600 ;
      RECT 27.1650 29.7600 28.0350 30.2600 ;
      RECT 26.2450 29.7600 26.6550 30.2600 ;
      RECT 25.3250 29.7600 25.7350 30.2600 ;
      RECT 24.4050 29.7600 24.8150 30.2600 ;
      RECT 23.0250 29.7600 23.8950 30.2600 ;
      RECT 22.1050 29.7600 22.5150 30.2600 ;
      RECT 21.1850 29.7600 21.5950 30.2600 ;
      RECT 19.8050 29.7600 20.6750 30.2600 ;
      RECT 18.8850 29.7600 19.2950 30.2600 ;
      RECT 17.9650 29.7600 18.3750 30.2600 ;
      RECT 17.0450 29.7600 17.4550 30.2600 ;
      RECT 15.6650 29.7600 16.5350 30.2600 ;
      RECT 14.7450 29.7600 15.1550 30.2600 ;
      RECT 13.8250 29.7600 14.2350 30.2600 ;
      RECT 12.4450 29.7600 13.3150 30.2600 ;
      RECT 11.5250 29.7600 11.9350 30.2600 ;
      RECT 10.6050 29.7600 11.0150 30.2600 ;
      RECT 9.6850 29.7600 10.0950 30.2600 ;
      RECT 8.3050 29.7600 9.1750 30.2600 ;
      RECT 7.3850 29.7600 7.7950 30.2600 ;
      RECT 6.4650 29.7600 6.8750 30.2600 ;
      RECT 5.5450 29.7600 5.9550 30.2600 ;
      RECT 0.0000 29.7600 5.0350 30.2600 ;
      RECT 0.0000 28.9850 100.2800 29.7600 ;
      RECT 0.5000 28.4750 100.2800 28.9850 ;
      RECT 0.0000 27.9650 100.2800 28.4750 ;
      RECT 0.0000 27.4550 99.7800 27.9650 ;
      RECT 0.0000 26.9450 100.2800 27.4550 ;
      RECT 0.5000 26.4350 100.2800 26.9450 ;
      RECT 0.0000 26.2650 100.2800 26.4350 ;
      RECT 0.0000 25.7550 99.7800 26.2650 ;
      RECT 0.0000 25.2450 100.2800 25.7550 ;
      RECT 0.5000 24.7350 100.2800 25.2450 ;
      RECT 0.0000 24.5650 100.2800 24.7350 ;
      RECT 0.0000 24.0550 99.7800 24.5650 ;
      RECT 0.0000 23.2050 100.2800 24.0550 ;
      RECT 0.5000 22.8650 100.2800 23.2050 ;
      RECT 0.5000 22.6950 99.7800 22.8650 ;
      RECT 0.0000 22.3550 99.7800 22.6950 ;
      RECT 0.0000 21.5050 100.2800 22.3550 ;
      RECT 0.5000 21.1650 100.2800 21.5050 ;
      RECT 0.5000 20.9950 99.7800 21.1650 ;
      RECT 0.0000 20.6550 99.7800 20.9950 ;
      RECT 0.0000 19.4650 100.2800 20.6550 ;
      RECT 0.5000 18.9550 99.7800 19.4650 ;
      RECT 0.0000 17.7650 100.2800 18.9550 ;
      RECT 0.5000 17.2550 99.7800 17.7650 ;
      RECT 0.0000 16.0650 100.2800 17.2550 ;
      RECT 0.5000 15.5550 99.7800 16.0650 ;
      RECT 0.0000 14.3650 100.2800 15.5550 ;
      RECT 0.0000 14.0250 99.7800 14.3650 ;
      RECT 0.5000 13.8550 99.7800 14.0250 ;
      RECT 0.5000 13.5150 100.2800 13.8550 ;
      RECT 0.0000 12.6650 100.2800 13.5150 ;
      RECT 0.0000 12.3250 99.7800 12.6650 ;
      RECT 0.5000 12.1550 99.7800 12.3250 ;
      RECT 0.5000 11.8150 100.2800 12.1550 ;
      RECT 0.0000 10.9650 100.2800 11.8150 ;
      RECT 0.0000 10.6250 99.7800 10.9650 ;
      RECT 0.5000 10.4550 99.7800 10.6250 ;
      RECT 0.5000 10.1150 100.2800 10.4550 ;
      RECT 0.0000 9.2650 100.2800 10.1150 ;
      RECT 0.0000 8.7550 99.7800 9.2650 ;
      RECT 0.0000 8.5850 100.2800 8.7550 ;
      RECT 0.5000 8.0750 100.2800 8.5850 ;
      RECT 0.0000 7.5650 100.2800 8.0750 ;
      RECT 0.0000 7.0550 99.7800 7.5650 ;
      RECT 0.0000 6.8850 100.2800 7.0550 ;
      RECT 0.5000 6.3750 100.2800 6.8850 ;
      RECT 0.0000 5.8650 100.2800 6.3750 ;
      RECT 0.0000 5.3550 99.7800 5.8650 ;
      RECT 0.0000 4.8450 100.2800 5.3550 ;
      RECT 0.5000 4.3350 100.2800 4.8450 ;
      RECT 0.0000 4.1650 100.2800 4.3350 ;
      RECT 0.0000 3.6550 99.7800 4.1650 ;
      RECT 0.0000 3.1450 100.2800 3.6550 ;
      RECT 0.5000 2.6350 100.2800 3.1450 ;
      RECT 0.0000 2.4650 100.2800 2.6350 ;
      RECT 0.0000 1.9550 99.7800 2.4650 ;
      RECT 0.0000 1.4450 100.2800 1.9550 ;
      RECT 0.5000 0.9350 100.2800 1.4450 ;
      RECT 0.0000 0.0000 100.2800 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 100.2800 30.2600 ;
    LAYER met2 ;
      RECT 97.9600 29.6350 100.2800 30.2600 ;
      RECT 97.0400 29.6350 97.5400 30.2600 ;
      RECT 96.1200 29.6350 96.6200 30.2600 ;
      RECT 95.2000 29.6350 95.7000 30.2600 ;
      RECT 94.7400 29.6350 94.7800 30.2600 ;
      RECT 93.8200 29.6350 94.3200 30.2600 ;
      RECT 92.9000 29.6350 93.4000 30.2600 ;
      RECT 91.9800 29.6350 92.4800 30.2600 ;
      RECT 91.5200 29.6350 91.5600 30.2600 ;
      RECT 90.6000 29.6350 91.1000 30.2600 ;
      RECT 89.6800 29.6350 90.1800 30.2600 ;
      RECT 88.7600 29.6350 89.2600 30.2600 ;
      RECT 88.3000 29.6350 88.3400 30.2600 ;
      RECT 87.8400 29.6350 87.8800 30.2600 ;
      RECT 86.9200 29.6350 87.4200 30.2600 ;
      RECT 86.0000 29.6350 86.5000 30.2600 ;
      RECT 85.0800 29.6350 85.5800 30.2600 ;
      RECT 84.1600 29.6350 84.6600 30.2600 ;
      RECT 83.2400 29.6350 83.7400 30.2600 ;
      RECT 82.7800 29.6350 82.8200 30.2600 ;
      RECT 0.0000 29.6350 82.3600 30.2600 ;
      RECT 0.0000 28.9400 100.2800 29.6350 ;
      RECT 0.0000 28.5200 99.6550 28.9400 ;
      RECT 0.0000 27.9200 100.2800 28.5200 ;
      RECT 0.6250 27.5000 100.2800 27.9200 ;
      RECT 0.0000 26.9000 100.2800 27.5000 ;
      RECT 0.0000 26.4800 99.6550 26.9000 ;
      RECT 0.0000 26.2200 100.2800 26.4800 ;
      RECT 0.6250 25.8000 100.2800 26.2200 ;
      RECT 0.0000 25.2000 100.2800 25.8000 ;
      RECT 0.0000 24.7800 99.6550 25.2000 ;
      RECT 0.0000 24.5200 100.2800 24.7800 ;
      RECT 0.6250 24.1000 100.2800 24.5200 ;
      RECT 0.0000 23.1600 100.2800 24.1000 ;
      RECT 0.0000 22.8200 99.6550 23.1600 ;
      RECT 0.6250 22.7400 99.6550 22.8200 ;
      RECT 0.6250 22.4000 100.2800 22.7400 ;
      RECT 0.0000 21.4600 100.2800 22.4000 ;
      RECT 0.0000 21.1200 99.6550 21.4600 ;
      RECT 0.6250 21.0400 99.6550 21.1200 ;
      RECT 0.6250 20.7000 100.2800 21.0400 ;
      RECT 0.0000 19.4200 100.2800 20.7000 ;
      RECT 0.6250 19.0000 99.6550 19.4200 ;
      RECT 0.0000 17.7200 100.2800 19.0000 ;
      RECT 0.6250 17.3000 99.6550 17.7200 ;
      RECT 0.0000 16.0200 100.2800 17.3000 ;
      RECT 0.6250 15.6000 99.6550 16.0200 ;
      RECT 0.0000 14.3200 100.2800 15.6000 ;
      RECT 0.6250 13.9800 100.2800 14.3200 ;
      RECT 0.6250 13.9000 99.6550 13.9800 ;
      RECT 0.0000 13.5600 99.6550 13.9000 ;
      RECT 0.0000 12.6200 100.2800 13.5600 ;
      RECT 0.6250 12.2800 100.2800 12.6200 ;
      RECT 0.6250 12.2000 99.6550 12.2800 ;
      RECT 0.0000 11.8600 99.6550 12.2000 ;
      RECT 0.0000 10.9200 100.2800 11.8600 ;
      RECT 0.6250 10.5800 100.2800 10.9200 ;
      RECT 0.6250 10.5000 99.6550 10.5800 ;
      RECT 0.0000 10.1600 99.6550 10.5000 ;
      RECT 0.0000 9.2200 100.2800 10.1600 ;
      RECT 0.6250 8.8000 100.2800 9.2200 ;
      RECT 0.0000 8.5400 100.2800 8.8000 ;
      RECT 0.0000 8.1200 99.6550 8.5400 ;
      RECT 0.0000 7.5200 100.2800 8.1200 ;
      RECT 0.6250 7.1000 100.2800 7.5200 ;
      RECT 0.0000 6.8400 100.2800 7.1000 ;
      RECT 0.0000 6.4200 99.6550 6.8400 ;
      RECT 0.0000 5.8200 100.2800 6.4200 ;
      RECT 0.6250 5.4000 100.2800 5.8200 ;
      RECT 0.0000 4.8000 100.2800 5.4000 ;
      RECT 0.0000 4.3800 99.6550 4.8000 ;
      RECT 0.0000 4.1200 100.2800 4.3800 ;
      RECT 0.6250 3.7000 100.2800 4.1200 ;
      RECT 0.0000 3.1000 100.2800 3.7000 ;
      RECT 0.0000 2.6800 99.6550 3.1000 ;
      RECT 0.0000 2.4200 100.2800 2.6800 ;
      RECT 0.6250 2.0000 100.2800 2.4200 ;
      RECT 0.0000 1.4000 100.2800 2.0000 ;
      RECT 0.0000 0.9800 99.6550 1.4000 ;
      RECT 0.0000 0.6250 100.2800 0.9800 ;
      RECT 97.9600 0.0000 100.2800 0.6250 ;
      RECT 97.0400 0.0000 97.5400 0.6250 ;
      RECT 96.1200 0.0000 96.6200 0.6250 ;
      RECT 95.2000 0.0000 95.7000 0.6250 ;
      RECT 94.7400 0.0000 94.7800 0.6250 ;
      RECT 93.8200 0.0000 94.3200 0.6250 ;
      RECT 92.9000 0.0000 93.4000 0.6250 ;
      RECT 91.9800 0.0000 92.4800 0.6250 ;
      RECT 91.5200 0.0000 91.5600 0.6250 ;
      RECT 90.6000 0.0000 91.1000 0.6250 ;
      RECT 89.6800 0.0000 90.1800 0.6250 ;
      RECT 88.7600 0.0000 89.2600 0.6250 ;
      RECT 88.3000 0.0000 88.3400 0.6250 ;
      RECT 87.3800 0.0000 87.8800 0.6250 ;
      RECT 86.4600 0.0000 86.9600 0.6250 ;
      RECT 85.5400 0.0000 86.0400 0.6250 ;
      RECT 85.0800 0.0000 85.1200 0.6250 ;
      RECT 84.1600 0.0000 84.6600 0.6250 ;
      RECT 83.2400 0.0000 83.7400 0.6250 ;
      RECT 82.7800 0.0000 82.8200 0.6250 ;
      RECT 0.0000 0.0000 82.3600 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 98.0200 25.7000 100.2800 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 100.2800 25.7000 ;
      RECT 95.0200 22.7000 100.2800 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 100.2800 22.7000 ;
      RECT 95.0200 20.2000 100.2800 21.2800 ;
      RECT 7.8600 20.2000 92.4200 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 98.0200 17.4800 100.2800 18.5600 ;
      RECT 4.8600 17.4800 95.4200 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 95.0200 14.7600 100.2800 15.8400 ;
      RECT 7.8600 14.7600 92.4200 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 98.0200 12.0400 100.2800 13.1200 ;
      RECT 4.8600 12.0400 95.4200 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 95.0200 9.3200 100.2800 10.4000 ;
      RECT 7.8600 9.3200 92.4200 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 100.2800 9.3200 ;
      RECT 98.0200 6.6000 100.2800 7.6800 ;
      RECT 4.8600 6.6000 95.4200 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 100.2800 6.6000 ;
      RECT 95.0200 3.7700 100.2800 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 100.2800 3.7700 ;
      RECT 98.0200 0.7700 100.2800 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 4.8600 25.3000 95.4200 28.3000 ;
      RECT 95.0200 3.7700 95.4200 25.3000 ;
      RECT 7.8600 3.7700 92.4200 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 98.0200 0.7700 100.2800 28.3000 ;
      RECT 4.8600 0.7700 95.4200 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
  END
END S_term_RAM_IO

END LIBRARY
