magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 39714 3456 40000
rect 0 286 286 39714
rect 0 0 3456 286
<< obsli1 >>
rect 120 120 3336 39880
<< obsm1 >>
rect 117 120 3339 39880
<< metal2 >>
rect 695 39341 1295 39782
rect 695 39165 1471 39341
rect 695 38423 1295 39165
rect 2095 39341 2695 39782
rect 1919 39165 2695 39341
rect 2095 38423 2695 39165
rect 695 0 1295 242
rect 1495 0 1895 242
rect 2095 0 2695 242
<< obsm2 >>
rect 115 38367 639 39782
rect 1351 39397 2039 39782
rect 1527 39109 1863 39397
rect 1351 38367 2039 39109
rect 2751 38367 3341 39782
rect 115 298 3341 38367
rect 115 242 639 298
rect 1351 242 1439 298
rect 1951 242 2039 298
rect 2751 242 3341 298
<< metal3 >>
rect 695 0 1295 166
rect 1495 0 1895 166
rect 2095 0 2695 166
<< obsm3 >>
rect 110 286 3346 39714
<< metal4 >>
rect 0 35157 254 39999
rect 3012 35157 3456 40000
rect 0 14007 254 19000
rect 3012 14007 3456 19000
rect 0 12817 254 13707
rect 3202 12817 3456 13707
rect 0 11647 254 12537
rect 3012 11647 3456 12537
rect 0 11281 3456 11347
rect 0 10625 3456 11221
rect 0 10329 254 10565
rect 3012 10329 3456 10565
rect 0 9673 3456 10269
rect 0 9547 3456 9613
rect 0 8317 254 9247
rect 3013 8317 3456 9247
rect 0 7347 254 8037
rect 3012 7347 3456 8037
rect 0 6377 254 7067
rect 3012 6377 3456 7067
rect 0 5167 254 6097
rect 3012 5167 3456 6097
rect 0 3957 254 4887
rect 3012 3957 3456 4887
rect 0 2987 215 3677
rect 3012 2987 3456 3677
rect 0 1777 254 2707
rect 3012 1777 3456 2707
rect 0 407 254 1497
rect 3012 407 3456 1497
<< obsm4 >>
rect 0 39999 3012 40000
rect 334 35077 2932 39999
rect 0 19080 3202 35077
rect 334 13927 2932 19080
rect 0 13787 3202 13927
rect 334 12737 3122 13787
rect 0 12617 3202 12737
rect 334 11567 2932 12617
rect 0 11427 3202 11567
rect 334 10349 2932 10545
rect 0 9327 3202 9467
rect 334 8237 2933 9327
rect 0 8117 3202 8237
rect 334 7267 2932 8117
rect 0 7147 3202 7267
rect 334 6297 2932 7147
rect 0 6177 3202 6297
rect 334 5087 2932 6177
rect 0 4967 3202 5087
rect 334 3877 2932 4967
rect 0 3757 3202 3877
rect 295 2907 2932 3757
rect 0 2787 3202 2907
rect 334 1697 2932 2787
rect 0 1577 3202 1697
rect 334 407 2932 1577
<< metal5 >>
rect 0 35157 254 40000
rect 3012 35157 3456 40000
rect 0 14007 254 18997
rect 3012 14007 3456 18997
rect 0 12837 254 13687
rect 3013 12837 3456 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 3012 11667 3456 12517
rect 3012 9547 3456 11347
rect 0 8337 254 9227
rect 3013 8337 3456 9227
rect 0 7367 254 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 3012 7367 3456 8017
rect 3012 6397 3456 7047
rect 3012 5187 3456 6077
rect 3012 3977 3456 4867
rect 0 3007 215 3657
rect 3012 3007 3456 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 3012 1797 3456 2687
rect 3012 427 3456 1477
<< obsm5 >>
rect 574 34837 2692 40000
rect 215 19317 3013 34837
rect 574 13687 2692 19317
rect 574 12837 2693 13687
rect 574 9227 2692 12837
rect 574 8337 2693 9227
rect 574 3657 2692 8337
rect 535 3007 2692 3657
rect 574 427 2692 3007
<< labels >>
rlabel metal3 s 1495 0 1895 166 6 cpos
port 1 nsew power bidirectional
rlabel metal2 s 1495 0 1895 242 6 cpos
port 1 nsew power bidirectional
rlabel metal3 s 2095 0 2695 166 6 cneg
port 2 nsew ground bidirectional
rlabel metal3 s 695 0 1295 166 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2095 0 2695 242 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 0 1295 242 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1295 39165 1471 39341 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 695 38423 1295 39782 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 1919 39165 2095 39341 6 cneg
port 2 nsew ground bidirectional
rlabel metal2 s 2095 38423 2695 39782 6 cneg
port 2 nsew ground bidirectional
rlabel metal5 s 3012 35157 3456 40000 6 vssio
port 3 nsew ground bidirectional
rlabel metal5 s 3012 5187 3456 6077 6 vssio
port 3 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 vssio
port 3 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 3012 35157 3456 40000 6 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 3012 5167 3456 6097 6 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 vssio
port 3 nsew ground bidirectional
rlabel metal4 s 0 35157 254 39999 6 vssio
port 3 nsew ground bidirectional
rlabel metal5 s 3013 12837 3456 13687 6 vddio_q
port 4 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 vddio_q
port 4 nsew power bidirectional
rlabel metal4 s 3202 12817 3456 13707 6 vddio_q
port 4 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 vddio_q
port 4 nsew power bidirectional
rlabel metal5 s 3012 14007 3456 18997 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 3012 3977 3456 4867 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 3012 14007 3456 19000 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 3012 3957 3456 4887 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 3012 11667 3456 12517 6 vssio_q
port 6 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 vssio_q
port 6 nsew ground bidirectional
rlabel metal4 s 3012 11647 3456 12537 6 vssio_q
port 6 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 vssio_q
port 6 nsew ground bidirectional
rlabel metal5 s 3012 1797 3456 2687 6 vccd
port 7 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 vccd
port 7 nsew power bidirectional
rlabel metal4 s 3012 1777 3456 2707 6 vccd
port 7 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 vccd
port 7 nsew power bidirectional
rlabel metal5 s 3012 7367 3456 8017 6 vssa
port 8 nsew ground bidirectional
rlabel metal5 s 3012 9547 3456 11347 6 vssa
port 8 nsew ground bidirectional
rlabel metal5 s 0 7367 254 8017 6 vssa
port 8 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 3012 7347 3456 8037 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 9547 3456 9613 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 3012 10329 3456 10565 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 11281 3456 11347 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 vssa
port 8 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 vssa
port 8 nsew ground bidirectional
rlabel metal5 s 3012 427 3456 1477 6 vcchib
port 9 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 vcchib
port 9 nsew power bidirectional
rlabel metal4 s 3012 407 3456 1497 6 vcchib
port 9 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 vcchib
port 9 nsew power bidirectional
rlabel metal5 s 3012 6397 3456 7047 6 vswitch
port 10 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 vswitch
port 10 nsew power bidirectional
rlabel metal4 s 3012 6377 3456 7067 6 vswitch
port 10 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 vswitch
port 10 nsew power bidirectional
rlabel metal5 s 3012 3007 3456 3657 6 vdda
port 11 nsew power bidirectional
rlabel metal5 s 0 3007 215 3657 6 vdda
port 11 nsew power bidirectional
rlabel metal4 s 3012 2987 3456 3677 6 vdda
port 11 nsew power bidirectional
rlabel metal4 s 0 2987 215 3677 6 vdda
port 11 nsew power bidirectional
rlabel metal5 s 3013 8337 3456 9227 6 vssd
port 12 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 vssd
port 12 nsew ground bidirectional
rlabel metal4 s 3013 8317 3456 9247 6 vssd
port 12 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 vssd
port 12 nsew ground bidirectional
rlabel metal4 s 0 9673 3456 10269 6 amuxbus_b
port 13 nsew signal bidirectional
rlabel metal4 s 0 10625 3456 11221 6 amuxbus_a
port 14 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 3456 40000
string LEFclass PAD
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 9654072
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8300788
<< end >>
