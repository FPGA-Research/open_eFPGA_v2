magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -68 -26 1749 162
<< ndiff >>
rect -42 119 0 136
rect -42 85 -34 119
rect -42 51 0 85
rect -42 17 -34 51
rect -42 0 0 17
rect 1681 119 1723 136
rect 1715 85 1723 119
rect 1681 51 1723 85
rect 1715 17 1723 51
rect 1681 0 1723 17
<< ndiffc >>
rect -34 85 0 119
rect -34 17 0 51
rect 1681 85 1715 119
rect 1681 17 1715 51
<< ndiffres >>
rect 0 0 1681 136
<< locali >>
rect -34 119 0 135
rect -34 51 0 85
rect -34 1 0 17
rect 1681 119 1715 135
rect 1681 51 1715 85
rect 1681 1 1715 17
use DFL1_CDNS_524688791851252  DFL1_CDNS_524688791851252_0
timestamp 1707688321
transform -1 0 8 0 1 5
box 0 0 1 1
use DFL1_CDNS_524688791851252  DFL1_CDNS_524688791851252_1
timestamp 1707688321
transform 1 0 1673 0 1 5
box 0 0 1 1
<< properties >>
string GDS_END 86902866
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86902360
<< end >>
