magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 2141 53
<< metal1 >>
rect -6 53 2147 56
rect -6 0 0 53
rect 2141 0 2147 53
rect -6 -3 2147 0
<< properties >>
string GDS_END 79043928
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79036116
<< end >>
