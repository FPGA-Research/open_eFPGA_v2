magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 402 217 668 283
rect 58 43 668 217
rect -26 -43 698 43
<< locali >>
rect 121 235 187 345
rect 306 235 372 345
rect 596 99 647 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 166 735 560 751
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 80 415 130 535
rect 166 451 560 701
rect 80 381 555 415
rect 236 199 270 381
rect 489 345 555 381
rect 18 113 200 199
rect 18 79 20 113
rect 54 79 92 113
rect 126 79 164 113
rect 198 79 200 113
rect 236 99 302 199
rect 408 113 526 265
rect 18 73 200 79
rect 408 79 414 113
rect 448 79 486 113
rect 520 79 526 113
rect 408 73 526 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 166 701 200 735
rect 238 701 272 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 20 79 54 113
rect 92 79 126 113
rect 164 79 198 113
rect 414 79 448 113
rect 486 79 520 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 166 735
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 20 113
rect 54 79 92 113
rect 126 79 164 113
rect 198 79 414 113
rect 448 79 486 113
rect 520 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel locali s 306 235 372 345 6 A
port 1 nsew signal input
rlabel locali s 121 235 187 345 6 B
port 2 nsew signal input
rlabel metal1 s 0 51 672 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 672 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 698 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 58 43 668 217 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 402 217 668 283 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 672 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 738 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 672 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 596 99 647 751 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 672 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 376290
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 367608
<< end >>
