magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< obsli1 >>
rect 385 1777 1913 1796
rect 190 1633 256 1699
rect 385 1671 412 1777
rect 1886 1671 1913 1777
rect 385 1659 1913 1671
rect 2042 1633 2108 1699
rect 190 1611 230 1633
rect 2068 1611 2108 1633
rect 41 1563 230 1611
rect 41 1529 60 1563
rect 94 1529 230 1563
rect 41 1491 230 1529
rect 41 1457 60 1491
rect 94 1457 230 1491
rect 41 1419 230 1457
rect 41 1385 60 1419
rect 94 1385 230 1419
rect 41 1347 230 1385
rect 41 1313 60 1347
rect 94 1313 230 1347
rect 41 1275 230 1313
rect 41 1241 60 1275
rect 94 1241 230 1275
rect 41 1203 230 1241
rect 41 1169 60 1203
rect 94 1169 230 1203
rect 41 1131 230 1169
rect 41 1097 60 1131
rect 94 1097 230 1131
rect 41 1059 230 1097
rect 41 1025 60 1059
rect 94 1025 230 1059
rect 41 987 230 1025
rect 41 953 60 987
rect 94 953 230 987
rect 41 915 230 953
rect 41 881 60 915
rect 94 881 230 915
rect 41 843 230 881
rect 41 809 60 843
rect 94 809 230 843
rect 41 771 230 809
rect 41 737 60 771
rect 94 737 230 771
rect 41 699 230 737
rect 41 665 60 699
rect 94 665 230 699
rect 41 627 230 665
rect 41 593 60 627
rect 94 593 230 627
rect 41 555 230 593
rect 41 521 60 555
rect 94 521 230 555
rect 41 483 230 521
rect 41 449 60 483
rect 94 449 230 483
rect 41 411 230 449
rect 41 377 60 411
rect 94 377 230 411
rect 41 339 230 377
rect 41 305 60 339
rect 94 305 230 339
rect 41 267 230 305
rect 41 233 60 267
rect 94 233 230 267
rect 41 185 230 233
rect 352 185 386 1611
rect 508 185 542 1611
rect 664 185 698 1611
rect 820 185 854 1611
rect 976 185 1010 1611
rect 1132 185 1166 1611
rect 1288 185 1322 1611
rect 1444 185 1478 1611
rect 1600 185 1634 1611
rect 1756 185 1790 1611
rect 1912 185 1946 1611
rect 2068 1563 2257 1611
rect 2068 1529 2204 1563
rect 2238 1529 2257 1563
rect 2068 1491 2257 1529
rect 2068 1457 2204 1491
rect 2238 1457 2257 1491
rect 2068 1419 2257 1457
rect 2068 1385 2204 1419
rect 2238 1385 2257 1419
rect 2068 1347 2257 1385
rect 2068 1313 2204 1347
rect 2238 1313 2257 1347
rect 2068 1275 2257 1313
rect 2068 1241 2204 1275
rect 2238 1241 2257 1275
rect 2068 1203 2257 1241
rect 2068 1169 2204 1203
rect 2238 1169 2257 1203
rect 2068 1131 2257 1169
rect 2068 1097 2204 1131
rect 2238 1097 2257 1131
rect 2068 1059 2257 1097
rect 2068 1025 2204 1059
rect 2238 1025 2257 1059
rect 2068 987 2257 1025
rect 2068 953 2204 987
rect 2238 953 2257 987
rect 2068 915 2257 953
rect 2068 881 2204 915
rect 2238 881 2257 915
rect 2068 843 2257 881
rect 2068 809 2204 843
rect 2238 809 2257 843
rect 2068 771 2257 809
rect 2068 737 2204 771
rect 2238 737 2257 771
rect 2068 699 2257 737
rect 2068 665 2204 699
rect 2238 665 2257 699
rect 2068 627 2257 665
rect 2068 593 2204 627
rect 2238 593 2257 627
rect 2068 555 2257 593
rect 2068 521 2204 555
rect 2238 521 2257 555
rect 2068 483 2257 521
rect 2068 449 2204 483
rect 2238 449 2257 483
rect 2068 411 2257 449
rect 2068 377 2204 411
rect 2238 377 2257 411
rect 2068 339 2257 377
rect 2068 305 2204 339
rect 2238 305 2257 339
rect 2068 267 2257 305
rect 2068 233 2204 267
rect 2238 233 2257 267
rect 2068 185 2257 233
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 97 256 163
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 97 2108 163
rect 385 0 1913 19
<< obsli1c >>
rect 412 1671 1886 1777
rect 60 1529 94 1563
rect 60 1457 94 1491
rect 60 1385 94 1419
rect 60 1313 94 1347
rect 60 1241 94 1275
rect 60 1169 94 1203
rect 60 1097 94 1131
rect 60 1025 94 1059
rect 60 953 94 987
rect 60 881 94 915
rect 60 809 94 843
rect 60 737 94 771
rect 60 665 94 699
rect 60 593 94 627
rect 60 521 94 555
rect 60 449 94 483
rect 60 377 94 411
rect 60 305 94 339
rect 60 233 94 267
rect 2204 1529 2238 1563
rect 2204 1457 2238 1491
rect 2204 1385 2238 1419
rect 2204 1313 2238 1347
rect 2204 1241 2238 1275
rect 2204 1169 2238 1203
rect 2204 1097 2238 1131
rect 2204 1025 2238 1059
rect 2204 953 2238 987
rect 2204 881 2238 915
rect 2204 809 2238 843
rect 2204 737 2238 771
rect 2204 665 2238 699
rect 2204 593 2238 627
rect 2204 521 2238 555
rect 2204 449 2238 483
rect 2204 377 2238 411
rect 2204 305 2238 339
rect 2204 233 2238 267
rect 412 19 1886 125
<< metal1 >>
rect 381 1777 1917 1796
rect 381 1671 412 1777
rect 1886 1671 1917 1777
rect 381 1659 1917 1671
rect 41 1563 100 1594
rect 41 1529 60 1563
rect 94 1529 100 1563
rect 41 1491 100 1529
rect 41 1457 60 1491
rect 94 1457 100 1491
rect 41 1419 100 1457
rect 41 1385 60 1419
rect 94 1385 100 1419
rect 41 1347 100 1385
rect 41 1313 60 1347
rect 94 1313 100 1347
rect 41 1275 100 1313
rect 41 1241 60 1275
rect 94 1241 100 1275
rect 41 1203 100 1241
rect 41 1169 60 1203
rect 94 1169 100 1203
rect 41 1131 100 1169
rect 41 1097 60 1131
rect 94 1097 100 1131
rect 41 1059 100 1097
rect 41 1025 60 1059
rect 94 1025 100 1059
rect 41 987 100 1025
rect 41 953 60 987
rect 94 953 100 987
rect 41 915 100 953
rect 41 881 60 915
rect 94 881 100 915
rect 41 843 100 881
rect 41 809 60 843
rect 94 809 100 843
rect 41 771 100 809
rect 41 737 60 771
rect 94 737 100 771
rect 41 699 100 737
rect 41 665 60 699
rect 94 665 100 699
rect 41 627 100 665
rect 41 593 60 627
rect 94 593 100 627
rect 41 555 100 593
rect 41 521 60 555
rect 94 521 100 555
rect 41 483 100 521
rect 41 449 60 483
rect 94 449 100 483
rect 41 411 100 449
rect 41 377 60 411
rect 94 377 100 411
rect 41 339 100 377
rect 41 305 60 339
rect 94 305 100 339
rect 41 267 100 305
rect 41 233 60 267
rect 94 233 100 267
rect 41 202 100 233
rect 2198 1563 2257 1594
rect 2198 1529 2204 1563
rect 2238 1529 2257 1563
rect 2198 1491 2257 1529
rect 2198 1457 2204 1491
rect 2238 1457 2257 1491
rect 2198 1419 2257 1457
rect 2198 1385 2204 1419
rect 2238 1385 2257 1419
rect 2198 1347 2257 1385
rect 2198 1313 2204 1347
rect 2238 1313 2257 1347
rect 2198 1275 2257 1313
rect 2198 1241 2204 1275
rect 2238 1241 2257 1275
rect 2198 1203 2257 1241
rect 2198 1169 2204 1203
rect 2238 1169 2257 1203
rect 2198 1131 2257 1169
rect 2198 1097 2204 1131
rect 2238 1097 2257 1131
rect 2198 1059 2257 1097
rect 2198 1025 2204 1059
rect 2238 1025 2257 1059
rect 2198 987 2257 1025
rect 2198 953 2204 987
rect 2238 953 2257 987
rect 2198 915 2257 953
rect 2198 881 2204 915
rect 2238 881 2257 915
rect 2198 843 2257 881
rect 2198 809 2204 843
rect 2238 809 2257 843
rect 2198 771 2257 809
rect 2198 737 2204 771
rect 2238 737 2257 771
rect 2198 699 2257 737
rect 2198 665 2204 699
rect 2238 665 2257 699
rect 2198 627 2257 665
rect 2198 593 2204 627
rect 2238 593 2257 627
rect 2198 555 2257 593
rect 2198 521 2204 555
rect 2238 521 2257 555
rect 2198 483 2257 521
rect 2198 449 2204 483
rect 2238 449 2257 483
rect 2198 411 2257 449
rect 2198 377 2204 411
rect 2238 377 2257 411
rect 2198 339 2257 377
rect 2198 305 2204 339
rect 2238 305 2257 339
rect 2198 267 2257 305
rect 2198 233 2204 267
rect 2238 233 2257 267
rect 2198 202 2257 233
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< obsm1 >>
rect 343 202 395 1594
rect 499 202 551 1594
rect 655 202 707 1594
rect 811 202 863 1594
rect 967 202 1019 1594
rect 1123 202 1175 1594
rect 1279 202 1331 1594
rect 1435 202 1487 1594
rect 1591 202 1643 1594
rect 1747 202 1799 1594
rect 1903 202 1955 1594
<< metal2 >>
rect 14 1274 2284 1594
rect 14 578 2284 1218
rect 14 202 2284 522
<< labels >>
rlabel metal2 s 14 578 2284 1218 6 DRAIN
port 1 nsew
rlabel metal1 s 381 1659 1917 1796 6 GATE
port 2 nsew
rlabel metal1 s 381 0 1917 137 6 GATE
port 2 nsew
rlabel metal2 s 14 1274 2284 1594 6 SOURCE
port 3 nsew
rlabel metal2 s 14 202 2284 522 6 SOURCE
port 3 nsew
rlabel metal1 s 41 202 100 1594 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 2198 202 2257 1594 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 2284 1796
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8686098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8617662
string device primitive
<< end >>
