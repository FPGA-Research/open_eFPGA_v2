magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 488 226
<< nmos >>
rect 0 0 100 200
rect 156 0 256 200
rect 312 0 412 200
<< ndiff >>
rect -50 0 0 200
rect 412 0 462 200
<< poly >>
rect 0 200 100 226
rect 0 -26 100 0
rect 156 200 256 226
rect 156 -26 256 0
rect 312 200 412 226
rect 312 -26 412 0
<< metal1 >>
rect -51 -16 -5 186
rect 105 -16 151 186
rect 261 -16 307 186
rect 417 -16 463 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1707688321
transform 1 0 256 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_1
timestamp 1707688321
transform 1 0 100 0 1 0
box -26 -26 82 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1707688321
transform 1 0 412 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 128 85 128 85 0 FreeSans 300 0 0 0 D
flabel comment s 284 85 284 85 0 FreeSans 300 0 0 0 S
flabel comment s 440 85 440 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86887254
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86885428
<< end >>
