magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 214 214 1978 1978
<< nwell >>
rect 134 1698 2058 2058
rect 134 494 494 1698
rect 1698 494 2058 1698
rect 134 134 2058 494
<< pwell >>
rect 0 2058 2192 2192
rect 0 134 134 2058
rect 628 628 1564 1564
rect 2058 134 2192 2058
rect 0 0 2192 134
<< ndiff >>
rect 896 1283 1296 1296
rect 896 909 909 1283
rect 1283 909 1296 1283
rect 896 896 1296 909
<< ndiffc >>
rect 909 909 1283 1283
<< psubdiff >>
rect 26 2142 2166 2166
rect 26 2108 50 2142
rect 84 2108 127 2142
rect 161 2108 195 2142
rect 229 2108 263 2142
rect 297 2108 331 2142
rect 365 2108 399 2142
rect 433 2108 467 2142
rect 501 2108 535 2142
rect 569 2108 603 2142
rect 637 2108 671 2142
rect 705 2108 739 2142
rect 773 2108 807 2142
rect 841 2108 875 2142
rect 909 2108 943 2142
rect 977 2108 1011 2142
rect 1045 2108 1079 2142
rect 1113 2108 1147 2142
rect 1181 2108 1215 2142
rect 1249 2108 1283 2142
rect 1317 2108 1351 2142
rect 1385 2108 1419 2142
rect 1453 2108 1487 2142
rect 1521 2108 1555 2142
rect 1589 2108 1623 2142
rect 1657 2108 1691 2142
rect 1725 2108 1759 2142
rect 1793 2108 1827 2142
rect 1861 2108 1895 2142
rect 1929 2108 1963 2142
rect 1997 2108 2031 2142
rect 2065 2108 2108 2142
rect 2142 2108 2166 2142
rect 26 2084 2166 2108
rect 26 2065 108 2084
rect 26 2031 50 2065
rect 84 2031 108 2065
rect 26 1997 108 2031
rect 26 1963 50 1997
rect 84 1963 108 1997
rect 26 1929 108 1963
rect 2084 2065 2166 2084
rect 2084 2031 2108 2065
rect 2142 2031 2166 2065
rect 2084 1997 2166 2031
rect 2084 1963 2108 1997
rect 2142 1963 2166 1997
rect 26 1895 50 1929
rect 84 1895 108 1929
rect 26 1861 108 1895
rect 26 1827 50 1861
rect 84 1827 108 1861
rect 26 1793 108 1827
rect 26 1759 50 1793
rect 84 1759 108 1793
rect 26 1725 108 1759
rect 26 1691 50 1725
rect 84 1691 108 1725
rect 26 1657 108 1691
rect 26 1623 50 1657
rect 84 1623 108 1657
rect 26 1589 108 1623
rect 26 1555 50 1589
rect 84 1555 108 1589
rect 26 1521 108 1555
rect 26 1487 50 1521
rect 84 1487 108 1521
rect 26 1453 108 1487
rect 26 1419 50 1453
rect 84 1419 108 1453
rect 26 1385 108 1419
rect 26 1351 50 1385
rect 84 1351 108 1385
rect 26 1317 108 1351
rect 26 1283 50 1317
rect 84 1283 108 1317
rect 26 1249 108 1283
rect 26 1215 50 1249
rect 84 1215 108 1249
rect 26 1181 108 1215
rect 26 1147 50 1181
rect 84 1147 108 1181
rect 26 1113 108 1147
rect 26 1079 50 1113
rect 84 1079 108 1113
rect 26 1045 108 1079
rect 26 1011 50 1045
rect 84 1011 108 1045
rect 26 977 108 1011
rect 26 943 50 977
rect 84 943 108 977
rect 26 909 108 943
rect 26 875 50 909
rect 84 875 108 909
rect 26 841 108 875
rect 26 807 50 841
rect 84 807 108 841
rect 26 773 108 807
rect 26 739 50 773
rect 84 739 108 773
rect 26 705 108 739
rect 26 671 50 705
rect 84 671 108 705
rect 26 637 108 671
rect 26 603 50 637
rect 84 603 108 637
rect 26 569 108 603
rect 26 535 50 569
rect 84 535 108 569
rect 26 501 108 535
rect 26 467 50 501
rect 84 467 108 501
rect 26 433 108 467
rect 26 399 50 433
rect 84 399 108 433
rect 26 365 108 399
rect 26 331 50 365
rect 84 331 108 365
rect 26 297 108 331
rect 26 263 50 297
rect 84 263 108 297
rect 26 229 108 263
rect 654 1514 1538 1538
rect 654 1480 678 1514
rect 712 1480 773 1514
rect 807 1480 841 1514
rect 875 1480 909 1514
rect 943 1480 977 1514
rect 1011 1480 1045 1514
rect 1079 1480 1113 1514
rect 1147 1480 1181 1514
rect 1215 1480 1249 1514
rect 1283 1480 1317 1514
rect 1351 1480 1385 1514
rect 1419 1480 1480 1514
rect 1514 1480 1538 1514
rect 654 1456 1538 1480
rect 654 1419 736 1456
rect 654 1385 678 1419
rect 712 1385 736 1419
rect 654 1351 736 1385
rect 654 1317 678 1351
rect 712 1317 736 1351
rect 654 1283 736 1317
rect 1456 1419 1538 1456
rect 1456 1385 1480 1419
rect 1514 1385 1538 1419
rect 1456 1351 1538 1385
rect 1456 1317 1480 1351
rect 1514 1317 1538 1351
rect 654 1249 678 1283
rect 712 1249 736 1283
rect 654 1215 736 1249
rect 654 1181 678 1215
rect 712 1181 736 1215
rect 654 1147 736 1181
rect 654 1113 678 1147
rect 712 1113 736 1147
rect 654 1079 736 1113
rect 654 1045 678 1079
rect 712 1045 736 1079
rect 654 1011 736 1045
rect 654 977 678 1011
rect 712 977 736 1011
rect 654 943 736 977
rect 654 909 678 943
rect 712 909 736 943
rect 654 875 736 909
rect 1456 1283 1538 1317
rect 1456 1249 1480 1283
rect 1514 1249 1538 1283
rect 1456 1215 1538 1249
rect 1456 1181 1480 1215
rect 1514 1181 1538 1215
rect 1456 1147 1538 1181
rect 1456 1113 1480 1147
rect 1514 1113 1538 1147
rect 1456 1079 1538 1113
rect 1456 1045 1480 1079
rect 1514 1045 1538 1079
rect 1456 1011 1538 1045
rect 1456 977 1480 1011
rect 1514 977 1538 1011
rect 1456 943 1538 977
rect 1456 909 1480 943
rect 1514 909 1538 943
rect 654 841 678 875
rect 712 841 736 875
rect 654 807 736 841
rect 654 773 678 807
rect 712 773 736 807
rect 654 736 736 773
rect 1456 875 1538 909
rect 1456 841 1480 875
rect 1514 841 1538 875
rect 1456 807 1538 841
rect 1456 773 1480 807
rect 1514 773 1538 807
rect 1456 736 1538 773
rect 654 712 1538 736
rect 654 678 678 712
rect 712 678 773 712
rect 807 678 841 712
rect 875 678 909 712
rect 943 678 977 712
rect 1011 678 1045 712
rect 1079 678 1113 712
rect 1147 678 1181 712
rect 1215 678 1249 712
rect 1283 678 1317 712
rect 1351 678 1385 712
rect 1419 678 1480 712
rect 1514 678 1538 712
rect 654 654 1538 678
rect 2084 1929 2166 1963
rect 2084 1895 2108 1929
rect 2142 1895 2166 1929
rect 2084 1861 2166 1895
rect 2084 1827 2108 1861
rect 2142 1827 2166 1861
rect 2084 1793 2166 1827
rect 2084 1759 2108 1793
rect 2142 1759 2166 1793
rect 2084 1725 2166 1759
rect 2084 1691 2108 1725
rect 2142 1691 2166 1725
rect 2084 1657 2166 1691
rect 2084 1623 2108 1657
rect 2142 1623 2166 1657
rect 2084 1589 2166 1623
rect 2084 1555 2108 1589
rect 2142 1555 2166 1589
rect 2084 1521 2166 1555
rect 2084 1487 2108 1521
rect 2142 1487 2166 1521
rect 2084 1453 2166 1487
rect 2084 1419 2108 1453
rect 2142 1419 2166 1453
rect 2084 1385 2166 1419
rect 2084 1351 2108 1385
rect 2142 1351 2166 1385
rect 2084 1317 2166 1351
rect 2084 1283 2108 1317
rect 2142 1283 2166 1317
rect 2084 1249 2166 1283
rect 2084 1215 2108 1249
rect 2142 1215 2166 1249
rect 2084 1181 2166 1215
rect 2084 1147 2108 1181
rect 2142 1147 2166 1181
rect 2084 1113 2166 1147
rect 2084 1079 2108 1113
rect 2142 1079 2166 1113
rect 2084 1045 2166 1079
rect 2084 1011 2108 1045
rect 2142 1011 2166 1045
rect 2084 977 2166 1011
rect 2084 943 2108 977
rect 2142 943 2166 977
rect 2084 909 2166 943
rect 2084 875 2108 909
rect 2142 875 2166 909
rect 2084 841 2166 875
rect 2084 807 2108 841
rect 2142 807 2166 841
rect 2084 773 2166 807
rect 2084 739 2108 773
rect 2142 739 2166 773
rect 2084 705 2166 739
rect 2084 671 2108 705
rect 2142 671 2166 705
rect 2084 637 2166 671
rect 2084 603 2108 637
rect 2142 603 2166 637
rect 2084 569 2166 603
rect 2084 535 2108 569
rect 2142 535 2166 569
rect 2084 501 2166 535
rect 2084 467 2108 501
rect 2142 467 2166 501
rect 2084 433 2166 467
rect 2084 399 2108 433
rect 2142 399 2166 433
rect 2084 365 2166 399
rect 2084 331 2108 365
rect 2142 331 2166 365
rect 2084 297 2166 331
rect 2084 263 2108 297
rect 2142 263 2166 297
rect 26 195 50 229
rect 84 195 108 229
rect 26 161 108 195
rect 26 127 50 161
rect 84 127 108 161
rect 26 108 108 127
rect 2084 229 2166 263
rect 2084 195 2108 229
rect 2142 195 2166 229
rect 2084 161 2166 195
rect 2084 127 2108 161
rect 2142 127 2166 161
rect 2084 108 2166 127
rect 26 84 2166 108
rect 26 50 50 84
rect 84 50 127 84
rect 161 50 195 84
rect 229 50 263 84
rect 297 50 331 84
rect 365 50 399 84
rect 433 50 467 84
rect 501 50 535 84
rect 569 50 603 84
rect 637 50 671 84
rect 705 50 739 84
rect 773 50 807 84
rect 841 50 875 84
rect 909 50 943 84
rect 977 50 1011 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1181 50 1215 84
rect 1249 50 1283 84
rect 1317 50 1351 84
rect 1385 50 1419 84
rect 1453 50 1487 84
rect 1521 50 1555 84
rect 1589 50 1623 84
rect 1657 50 1691 84
rect 1725 50 1759 84
rect 1793 50 1827 84
rect 1861 50 1895 84
rect 1929 50 1963 84
rect 1997 50 2031 84
rect 2065 50 2108 84
rect 2142 50 2166 84
rect 26 26 2166 50
<< nsubdiff >>
rect 252 1916 1940 1940
rect 252 1882 276 1916
rect 310 1882 365 1916
rect 399 1882 433 1916
rect 467 1882 501 1916
rect 535 1882 569 1916
rect 603 1882 637 1916
rect 671 1882 705 1916
rect 739 1882 773 1916
rect 807 1882 841 1916
rect 875 1882 909 1916
rect 943 1882 977 1916
rect 1011 1882 1045 1916
rect 1079 1882 1113 1916
rect 1147 1882 1181 1916
rect 1215 1882 1249 1916
rect 1283 1882 1317 1916
rect 1351 1882 1385 1916
rect 1419 1882 1453 1916
rect 1487 1882 1521 1916
rect 1555 1882 1589 1916
rect 1623 1882 1657 1916
rect 1691 1882 1725 1916
rect 1759 1882 1793 1916
rect 1827 1882 1882 1916
rect 1916 1882 1940 1916
rect 252 1858 1940 1882
rect 252 1827 334 1858
rect 252 1793 276 1827
rect 310 1793 334 1827
rect 252 1759 334 1793
rect 252 1725 276 1759
rect 310 1725 334 1759
rect 252 1691 334 1725
rect 252 1657 276 1691
rect 310 1657 334 1691
rect 252 1623 334 1657
rect 252 1589 276 1623
rect 310 1589 334 1623
rect 252 1555 334 1589
rect 252 1521 276 1555
rect 310 1521 334 1555
rect 1858 1827 1940 1858
rect 1858 1793 1882 1827
rect 1916 1793 1940 1827
rect 1858 1759 1940 1793
rect 1858 1725 1882 1759
rect 1916 1725 1940 1759
rect 1858 1691 1940 1725
rect 1858 1657 1882 1691
rect 1916 1657 1940 1691
rect 1858 1623 1940 1657
rect 1858 1589 1882 1623
rect 1916 1589 1940 1623
rect 1858 1555 1940 1589
rect 252 1487 334 1521
rect 252 1453 276 1487
rect 310 1453 334 1487
rect 252 1419 334 1453
rect 252 1385 276 1419
rect 310 1385 334 1419
rect 252 1351 334 1385
rect 252 1317 276 1351
rect 310 1317 334 1351
rect 252 1283 334 1317
rect 252 1249 276 1283
rect 310 1249 334 1283
rect 252 1215 334 1249
rect 252 1181 276 1215
rect 310 1181 334 1215
rect 252 1147 334 1181
rect 252 1113 276 1147
rect 310 1113 334 1147
rect 252 1079 334 1113
rect 252 1045 276 1079
rect 310 1045 334 1079
rect 252 1011 334 1045
rect 252 977 276 1011
rect 310 977 334 1011
rect 252 943 334 977
rect 252 909 276 943
rect 310 909 334 943
rect 252 875 334 909
rect 252 841 276 875
rect 310 841 334 875
rect 252 807 334 841
rect 252 773 276 807
rect 310 773 334 807
rect 252 739 334 773
rect 252 705 276 739
rect 310 705 334 739
rect 252 671 334 705
rect 252 637 276 671
rect 310 637 334 671
rect 1858 1521 1882 1555
rect 1916 1521 1940 1555
rect 1858 1487 1940 1521
rect 1858 1453 1882 1487
rect 1916 1453 1940 1487
rect 1858 1419 1940 1453
rect 1858 1385 1882 1419
rect 1916 1385 1940 1419
rect 1858 1351 1940 1385
rect 1858 1317 1882 1351
rect 1916 1317 1940 1351
rect 1858 1283 1940 1317
rect 1858 1249 1882 1283
rect 1916 1249 1940 1283
rect 1858 1215 1940 1249
rect 1858 1181 1882 1215
rect 1916 1181 1940 1215
rect 1858 1147 1940 1181
rect 1858 1113 1882 1147
rect 1916 1113 1940 1147
rect 1858 1079 1940 1113
rect 1858 1045 1882 1079
rect 1916 1045 1940 1079
rect 1858 1011 1940 1045
rect 1858 977 1882 1011
rect 1916 977 1940 1011
rect 1858 943 1940 977
rect 1858 909 1882 943
rect 1916 909 1940 943
rect 1858 875 1940 909
rect 1858 841 1882 875
rect 1916 841 1940 875
rect 1858 807 1940 841
rect 1858 773 1882 807
rect 1916 773 1940 807
rect 1858 739 1940 773
rect 1858 705 1882 739
rect 1916 705 1940 739
rect 1858 671 1940 705
rect 252 603 334 637
rect 252 569 276 603
rect 310 569 334 603
rect 252 535 334 569
rect 252 501 276 535
rect 310 501 334 535
rect 252 467 334 501
rect 252 433 276 467
rect 310 433 334 467
rect 252 399 334 433
rect 252 365 276 399
rect 310 365 334 399
rect 252 334 334 365
rect 1858 637 1882 671
rect 1916 637 1940 671
rect 1858 603 1940 637
rect 1858 569 1882 603
rect 1916 569 1940 603
rect 1858 535 1940 569
rect 1858 501 1882 535
rect 1916 501 1940 535
rect 1858 467 1940 501
rect 1858 433 1882 467
rect 1916 433 1940 467
rect 1858 399 1940 433
rect 1858 365 1882 399
rect 1916 365 1940 399
rect 1858 334 1940 365
rect 252 310 1940 334
rect 252 276 276 310
rect 310 276 365 310
rect 399 276 433 310
rect 467 276 501 310
rect 535 276 569 310
rect 603 276 637 310
rect 671 276 705 310
rect 739 276 773 310
rect 807 276 841 310
rect 875 276 909 310
rect 943 276 977 310
rect 1011 276 1045 310
rect 1079 276 1113 310
rect 1147 276 1181 310
rect 1215 276 1249 310
rect 1283 276 1317 310
rect 1351 276 1385 310
rect 1419 276 1453 310
rect 1487 276 1521 310
rect 1555 276 1589 310
rect 1623 276 1657 310
rect 1691 276 1725 310
rect 1759 276 1793 310
rect 1827 276 1882 310
rect 1916 276 1940 310
rect 252 252 1940 276
<< psubdiffcont >>
rect 50 2108 84 2142
rect 127 2108 161 2142
rect 195 2108 229 2142
rect 263 2108 297 2142
rect 331 2108 365 2142
rect 399 2108 433 2142
rect 467 2108 501 2142
rect 535 2108 569 2142
rect 603 2108 637 2142
rect 671 2108 705 2142
rect 739 2108 773 2142
rect 807 2108 841 2142
rect 875 2108 909 2142
rect 943 2108 977 2142
rect 1011 2108 1045 2142
rect 1079 2108 1113 2142
rect 1147 2108 1181 2142
rect 1215 2108 1249 2142
rect 1283 2108 1317 2142
rect 1351 2108 1385 2142
rect 1419 2108 1453 2142
rect 1487 2108 1521 2142
rect 1555 2108 1589 2142
rect 1623 2108 1657 2142
rect 1691 2108 1725 2142
rect 1759 2108 1793 2142
rect 1827 2108 1861 2142
rect 1895 2108 1929 2142
rect 1963 2108 1997 2142
rect 2031 2108 2065 2142
rect 2108 2108 2142 2142
rect 50 2031 84 2065
rect 50 1963 84 1997
rect 2108 2031 2142 2065
rect 2108 1963 2142 1997
rect 50 1895 84 1929
rect 50 1827 84 1861
rect 50 1759 84 1793
rect 50 1691 84 1725
rect 50 1623 84 1657
rect 50 1555 84 1589
rect 50 1487 84 1521
rect 50 1419 84 1453
rect 50 1351 84 1385
rect 50 1283 84 1317
rect 50 1215 84 1249
rect 50 1147 84 1181
rect 50 1079 84 1113
rect 50 1011 84 1045
rect 50 943 84 977
rect 50 875 84 909
rect 50 807 84 841
rect 50 739 84 773
rect 50 671 84 705
rect 50 603 84 637
rect 50 535 84 569
rect 50 467 84 501
rect 50 399 84 433
rect 50 331 84 365
rect 50 263 84 297
rect 678 1480 712 1514
rect 773 1480 807 1514
rect 841 1480 875 1514
rect 909 1480 943 1514
rect 977 1480 1011 1514
rect 1045 1480 1079 1514
rect 1113 1480 1147 1514
rect 1181 1480 1215 1514
rect 1249 1480 1283 1514
rect 1317 1480 1351 1514
rect 1385 1480 1419 1514
rect 1480 1480 1514 1514
rect 678 1385 712 1419
rect 678 1317 712 1351
rect 1480 1385 1514 1419
rect 1480 1317 1514 1351
rect 678 1249 712 1283
rect 678 1181 712 1215
rect 678 1113 712 1147
rect 678 1045 712 1079
rect 678 977 712 1011
rect 678 909 712 943
rect 1480 1249 1514 1283
rect 1480 1181 1514 1215
rect 1480 1113 1514 1147
rect 1480 1045 1514 1079
rect 1480 977 1514 1011
rect 1480 909 1514 943
rect 678 841 712 875
rect 678 773 712 807
rect 1480 841 1514 875
rect 1480 773 1514 807
rect 678 678 712 712
rect 773 678 807 712
rect 841 678 875 712
rect 909 678 943 712
rect 977 678 1011 712
rect 1045 678 1079 712
rect 1113 678 1147 712
rect 1181 678 1215 712
rect 1249 678 1283 712
rect 1317 678 1351 712
rect 1385 678 1419 712
rect 1480 678 1514 712
rect 2108 1895 2142 1929
rect 2108 1827 2142 1861
rect 2108 1759 2142 1793
rect 2108 1691 2142 1725
rect 2108 1623 2142 1657
rect 2108 1555 2142 1589
rect 2108 1487 2142 1521
rect 2108 1419 2142 1453
rect 2108 1351 2142 1385
rect 2108 1283 2142 1317
rect 2108 1215 2142 1249
rect 2108 1147 2142 1181
rect 2108 1079 2142 1113
rect 2108 1011 2142 1045
rect 2108 943 2142 977
rect 2108 875 2142 909
rect 2108 807 2142 841
rect 2108 739 2142 773
rect 2108 671 2142 705
rect 2108 603 2142 637
rect 2108 535 2142 569
rect 2108 467 2142 501
rect 2108 399 2142 433
rect 2108 331 2142 365
rect 2108 263 2142 297
rect 50 195 84 229
rect 50 127 84 161
rect 2108 195 2142 229
rect 2108 127 2142 161
rect 50 50 84 84
rect 127 50 161 84
rect 195 50 229 84
rect 263 50 297 84
rect 331 50 365 84
rect 399 50 433 84
rect 467 50 501 84
rect 535 50 569 84
rect 603 50 637 84
rect 671 50 705 84
rect 739 50 773 84
rect 807 50 841 84
rect 875 50 909 84
rect 943 50 977 84
rect 1011 50 1045 84
rect 1079 50 1113 84
rect 1147 50 1181 84
rect 1215 50 1249 84
rect 1283 50 1317 84
rect 1351 50 1385 84
rect 1419 50 1453 84
rect 1487 50 1521 84
rect 1555 50 1589 84
rect 1623 50 1657 84
rect 1691 50 1725 84
rect 1759 50 1793 84
rect 1827 50 1861 84
rect 1895 50 1929 84
rect 1963 50 1997 84
rect 2031 50 2065 84
rect 2108 50 2142 84
<< nsubdiffcont >>
rect 276 1882 310 1916
rect 365 1882 399 1916
rect 433 1882 467 1916
rect 501 1882 535 1916
rect 569 1882 603 1916
rect 637 1882 671 1916
rect 705 1882 739 1916
rect 773 1882 807 1916
rect 841 1882 875 1916
rect 909 1882 943 1916
rect 977 1882 1011 1916
rect 1045 1882 1079 1916
rect 1113 1882 1147 1916
rect 1181 1882 1215 1916
rect 1249 1882 1283 1916
rect 1317 1882 1351 1916
rect 1385 1882 1419 1916
rect 1453 1882 1487 1916
rect 1521 1882 1555 1916
rect 1589 1882 1623 1916
rect 1657 1882 1691 1916
rect 1725 1882 1759 1916
rect 1793 1882 1827 1916
rect 1882 1882 1916 1916
rect 276 1793 310 1827
rect 276 1725 310 1759
rect 276 1657 310 1691
rect 276 1589 310 1623
rect 276 1521 310 1555
rect 1882 1793 1916 1827
rect 1882 1725 1916 1759
rect 1882 1657 1916 1691
rect 1882 1589 1916 1623
rect 276 1453 310 1487
rect 276 1385 310 1419
rect 276 1317 310 1351
rect 276 1249 310 1283
rect 276 1181 310 1215
rect 276 1113 310 1147
rect 276 1045 310 1079
rect 276 977 310 1011
rect 276 909 310 943
rect 276 841 310 875
rect 276 773 310 807
rect 276 705 310 739
rect 276 637 310 671
rect 1882 1521 1916 1555
rect 1882 1453 1916 1487
rect 1882 1385 1916 1419
rect 1882 1317 1916 1351
rect 1882 1249 1916 1283
rect 1882 1181 1916 1215
rect 1882 1113 1916 1147
rect 1882 1045 1916 1079
rect 1882 977 1916 1011
rect 1882 909 1916 943
rect 1882 841 1916 875
rect 1882 773 1916 807
rect 1882 705 1916 739
rect 276 569 310 603
rect 276 501 310 535
rect 276 433 310 467
rect 276 365 310 399
rect 1882 637 1916 671
rect 1882 569 1916 603
rect 1882 501 1916 535
rect 1882 433 1916 467
rect 1882 365 1916 399
rect 276 276 310 310
rect 365 276 399 310
rect 433 276 467 310
rect 501 276 535 310
rect 569 276 603 310
rect 637 276 671 310
rect 705 276 739 310
rect 773 276 807 310
rect 841 276 875 310
rect 909 276 943 310
rect 977 276 1011 310
rect 1045 276 1079 310
rect 1113 276 1147 310
rect 1181 276 1215 310
rect 1249 276 1283 310
rect 1317 276 1351 310
rect 1385 276 1419 310
rect 1453 276 1487 310
rect 1521 276 1555 310
rect 1589 276 1623 310
rect 1657 276 1691 310
rect 1725 276 1759 310
rect 1793 276 1827 310
rect 1882 276 1916 310
<< locali >>
rect 34 2142 2158 2158
rect 34 2108 50 2142
rect 84 2108 127 2142
rect 177 2108 195 2142
rect 249 2108 263 2142
rect 321 2108 331 2142
rect 393 2108 399 2142
rect 465 2108 467 2142
rect 501 2108 503 2142
rect 569 2108 575 2142
rect 637 2108 647 2142
rect 705 2108 719 2142
rect 773 2108 791 2142
rect 841 2108 863 2142
rect 909 2108 935 2142
rect 977 2108 1007 2142
rect 1045 2108 1079 2142
rect 1113 2108 1147 2142
rect 1185 2108 1215 2142
rect 1257 2108 1283 2142
rect 1329 2108 1351 2142
rect 1401 2108 1419 2142
rect 1473 2108 1487 2142
rect 1545 2108 1555 2142
rect 1617 2108 1623 2142
rect 1689 2108 1691 2142
rect 1725 2108 1727 2142
rect 1793 2108 1799 2142
rect 1861 2108 1871 2142
rect 1929 2108 1943 2142
rect 1997 2108 2015 2142
rect 2065 2108 2108 2142
rect 2142 2108 2158 2142
rect 34 2092 2158 2108
rect 34 2065 100 2092
rect 34 2015 50 2065
rect 84 2015 100 2065
rect 34 1997 100 2015
rect 34 1943 50 1997
rect 84 1943 100 1997
rect 34 1929 100 1943
rect 2092 2065 2158 2092
rect 2092 2015 2108 2065
rect 2142 2015 2158 2065
rect 2092 1997 2158 2015
rect 2092 1943 2108 1997
rect 2142 1943 2158 1997
rect 34 1871 50 1929
rect 84 1871 100 1929
rect 34 1861 100 1871
rect 34 1799 50 1861
rect 84 1799 100 1861
rect 34 1793 100 1799
rect 34 1727 50 1793
rect 84 1727 100 1793
rect 34 1725 100 1727
rect 34 1691 50 1725
rect 84 1691 100 1725
rect 34 1689 100 1691
rect 34 1623 50 1689
rect 84 1623 100 1689
rect 34 1617 100 1623
rect 34 1555 50 1617
rect 84 1555 100 1617
rect 34 1545 100 1555
rect 34 1487 50 1545
rect 84 1487 100 1545
rect 34 1473 100 1487
rect 34 1419 50 1473
rect 84 1419 100 1473
rect 34 1401 100 1419
rect 34 1351 50 1401
rect 84 1351 100 1401
rect 34 1329 100 1351
rect 34 1283 50 1329
rect 84 1283 100 1329
rect 34 1257 100 1283
rect 34 1215 50 1257
rect 84 1215 100 1257
rect 34 1185 100 1215
rect 34 1147 50 1185
rect 84 1147 100 1185
rect 34 1113 100 1147
rect 34 1079 50 1113
rect 84 1079 100 1113
rect 34 1045 100 1079
rect 34 1007 50 1045
rect 84 1007 100 1045
rect 34 977 100 1007
rect 34 935 50 977
rect 84 935 100 977
rect 34 909 100 935
rect 34 863 50 909
rect 84 863 100 909
rect 34 841 100 863
rect 34 791 50 841
rect 84 791 100 841
rect 34 773 100 791
rect 34 719 50 773
rect 84 719 100 773
rect 34 705 100 719
rect 34 647 50 705
rect 84 647 100 705
rect 34 637 100 647
rect 34 575 50 637
rect 84 575 100 637
rect 34 569 100 575
rect 34 503 50 569
rect 84 503 100 569
rect 34 501 100 503
rect 34 467 50 501
rect 84 467 100 501
rect 34 465 100 467
rect 34 399 50 465
rect 84 399 100 465
rect 34 393 100 399
rect 34 331 50 393
rect 84 331 100 393
rect 34 321 100 331
rect 34 263 50 321
rect 84 263 100 321
rect 34 249 100 263
rect 260 1916 1932 1932
rect 260 1882 276 1916
rect 310 1882 359 1916
rect 399 1882 431 1916
rect 467 1882 501 1916
rect 537 1882 569 1916
rect 609 1882 637 1916
rect 681 1882 705 1916
rect 753 1882 773 1916
rect 825 1882 841 1916
rect 897 1882 909 1916
rect 969 1882 977 1916
rect 1041 1882 1045 1916
rect 1147 1882 1151 1916
rect 1215 1882 1223 1916
rect 1283 1882 1295 1916
rect 1351 1882 1367 1916
rect 1419 1882 1439 1916
rect 1487 1882 1511 1916
rect 1555 1882 1583 1916
rect 1623 1882 1655 1916
rect 1691 1882 1725 1916
rect 1761 1882 1793 1916
rect 1833 1882 1882 1916
rect 1916 1882 1932 1916
rect 260 1866 1932 1882
rect 260 1833 326 1866
rect 260 1793 276 1833
rect 310 1793 326 1833
rect 260 1761 326 1793
rect 260 1725 276 1761
rect 310 1725 326 1761
rect 260 1691 326 1725
rect 260 1655 276 1691
rect 310 1655 326 1691
rect 260 1623 326 1655
rect 260 1583 276 1623
rect 310 1583 326 1623
rect 260 1555 326 1583
rect 260 1511 276 1555
rect 310 1511 326 1555
rect 1866 1833 1932 1866
rect 1866 1793 1882 1833
rect 1916 1793 1932 1833
rect 1866 1761 1932 1793
rect 1866 1725 1882 1761
rect 1916 1725 1932 1761
rect 1866 1691 1932 1725
rect 1866 1655 1882 1691
rect 1916 1655 1932 1691
rect 1866 1623 1932 1655
rect 1866 1583 1882 1623
rect 1916 1583 1932 1623
rect 1866 1555 1932 1583
rect 260 1487 326 1511
rect 260 1439 276 1487
rect 310 1439 326 1487
rect 260 1419 326 1439
rect 260 1367 276 1419
rect 310 1367 326 1419
rect 260 1351 326 1367
rect 260 1295 276 1351
rect 310 1295 326 1351
rect 260 1283 326 1295
rect 260 1223 276 1283
rect 310 1223 326 1283
rect 260 1215 326 1223
rect 260 1151 276 1215
rect 310 1151 326 1215
rect 260 1147 326 1151
rect 260 1045 276 1147
rect 310 1045 326 1147
rect 260 1041 326 1045
rect 260 977 276 1041
rect 310 977 326 1041
rect 260 969 326 977
rect 260 909 276 969
rect 310 909 326 969
rect 260 897 326 909
rect 260 841 276 897
rect 310 841 326 897
rect 260 825 326 841
rect 260 773 276 825
rect 310 773 326 825
rect 260 753 326 773
rect 260 705 276 753
rect 310 705 326 753
rect 260 681 326 705
rect 260 637 276 681
rect 310 637 326 681
rect 662 1514 1530 1530
rect 662 1480 678 1514
rect 712 1480 755 1514
rect 807 1480 827 1514
rect 875 1480 899 1514
rect 943 1480 971 1514
rect 1011 1480 1043 1514
rect 1079 1480 1113 1514
rect 1149 1480 1181 1514
rect 1221 1480 1249 1514
rect 1293 1480 1317 1514
rect 1365 1480 1385 1514
rect 1437 1480 1480 1514
rect 1514 1480 1530 1514
rect 662 1464 1530 1480
rect 662 1437 728 1464
rect 662 1385 678 1437
rect 712 1385 728 1437
rect 662 1365 728 1385
rect 662 1317 678 1365
rect 712 1317 728 1365
rect 662 1293 728 1317
rect 1464 1437 1530 1464
rect 1464 1385 1480 1437
rect 1514 1385 1530 1437
rect 1464 1365 1530 1385
rect 1464 1317 1480 1365
rect 1514 1317 1530 1365
rect 662 1249 678 1293
rect 712 1249 728 1293
rect 662 1221 728 1249
rect 662 1181 678 1221
rect 712 1181 728 1221
rect 662 1149 728 1181
rect 662 1113 678 1149
rect 712 1113 728 1149
rect 662 1079 728 1113
rect 662 1043 678 1079
rect 712 1043 728 1079
rect 662 1011 728 1043
rect 662 971 678 1011
rect 712 971 728 1011
rect 662 943 728 971
rect 662 899 678 943
rect 712 899 728 943
rect 662 875 728 899
rect 893 1283 1299 1299
rect 893 909 909 1283
rect 1283 909 1299 1283
rect 893 893 1299 909
rect 1464 1293 1530 1317
rect 1464 1249 1480 1293
rect 1514 1249 1530 1293
rect 1464 1221 1530 1249
rect 1464 1181 1480 1221
rect 1514 1181 1530 1221
rect 1464 1149 1530 1181
rect 1464 1113 1480 1149
rect 1514 1113 1530 1149
rect 1464 1079 1530 1113
rect 1464 1043 1480 1079
rect 1514 1043 1530 1079
rect 1464 1011 1530 1043
rect 1464 971 1480 1011
rect 1514 971 1530 1011
rect 1464 943 1530 971
rect 1464 899 1480 943
rect 1514 899 1530 943
rect 662 827 678 875
rect 712 827 728 875
rect 662 807 728 827
rect 662 755 678 807
rect 712 755 728 807
rect 662 728 728 755
rect 1464 875 1530 899
rect 1464 827 1480 875
rect 1514 827 1530 875
rect 1464 807 1530 827
rect 1464 755 1480 807
rect 1514 755 1530 807
rect 1464 728 1530 755
rect 662 712 1530 728
rect 662 678 678 712
rect 712 678 755 712
rect 807 678 827 712
rect 875 678 899 712
rect 943 678 971 712
rect 1011 678 1043 712
rect 1079 678 1113 712
rect 1149 678 1181 712
rect 1221 678 1249 712
rect 1293 678 1317 712
rect 1365 678 1385 712
rect 1437 678 1480 712
rect 1514 678 1530 712
rect 662 662 1530 678
rect 1866 1511 1882 1555
rect 1916 1511 1932 1555
rect 1866 1487 1932 1511
rect 1866 1439 1882 1487
rect 1916 1439 1932 1487
rect 1866 1419 1932 1439
rect 1866 1367 1882 1419
rect 1916 1367 1932 1419
rect 1866 1351 1932 1367
rect 1866 1295 1882 1351
rect 1916 1295 1932 1351
rect 1866 1283 1932 1295
rect 1866 1223 1882 1283
rect 1916 1223 1932 1283
rect 1866 1215 1932 1223
rect 1866 1151 1882 1215
rect 1916 1151 1932 1215
rect 1866 1147 1932 1151
rect 1866 1045 1882 1147
rect 1916 1045 1932 1147
rect 1866 1041 1932 1045
rect 1866 977 1882 1041
rect 1916 977 1932 1041
rect 1866 969 1932 977
rect 1866 909 1882 969
rect 1916 909 1932 969
rect 1866 897 1932 909
rect 1866 841 1882 897
rect 1916 841 1932 897
rect 1866 825 1932 841
rect 1866 773 1882 825
rect 1916 773 1932 825
rect 1866 753 1932 773
rect 1866 705 1882 753
rect 1916 705 1932 753
rect 1866 681 1932 705
rect 260 609 326 637
rect 260 569 276 609
rect 310 569 326 609
rect 260 537 326 569
rect 260 501 276 537
rect 310 501 326 537
rect 260 467 326 501
rect 260 431 276 467
rect 310 431 326 467
rect 260 399 326 431
rect 260 359 276 399
rect 310 359 326 399
rect 260 326 326 359
rect 1866 637 1882 681
rect 1916 637 1932 681
rect 1866 609 1932 637
rect 1866 569 1882 609
rect 1916 569 1932 609
rect 1866 537 1932 569
rect 1866 501 1882 537
rect 1916 501 1932 537
rect 1866 467 1932 501
rect 1866 431 1882 467
rect 1916 431 1932 467
rect 1866 399 1932 431
rect 1866 359 1882 399
rect 1916 359 1932 399
rect 1866 326 1932 359
rect 260 310 1932 326
rect 260 276 276 310
rect 310 276 359 310
rect 399 276 431 310
rect 467 276 501 310
rect 537 276 569 310
rect 609 276 637 310
rect 681 276 705 310
rect 753 276 773 310
rect 825 276 841 310
rect 897 276 909 310
rect 969 276 977 310
rect 1041 276 1045 310
rect 1147 276 1151 310
rect 1215 276 1223 310
rect 1283 276 1295 310
rect 1351 276 1367 310
rect 1419 276 1439 310
rect 1487 276 1511 310
rect 1555 276 1583 310
rect 1623 276 1655 310
rect 1691 276 1725 310
rect 1761 276 1793 310
rect 1833 276 1882 310
rect 1916 276 1932 310
rect 260 260 1932 276
rect 2092 1929 2158 1943
rect 2092 1871 2108 1929
rect 2142 1871 2158 1929
rect 2092 1861 2158 1871
rect 2092 1799 2108 1861
rect 2142 1799 2158 1861
rect 2092 1793 2158 1799
rect 2092 1727 2108 1793
rect 2142 1727 2158 1793
rect 2092 1725 2158 1727
rect 2092 1691 2108 1725
rect 2142 1691 2158 1725
rect 2092 1689 2158 1691
rect 2092 1623 2108 1689
rect 2142 1623 2158 1689
rect 2092 1617 2158 1623
rect 2092 1555 2108 1617
rect 2142 1555 2158 1617
rect 2092 1545 2158 1555
rect 2092 1487 2108 1545
rect 2142 1487 2158 1545
rect 2092 1473 2158 1487
rect 2092 1419 2108 1473
rect 2142 1419 2158 1473
rect 2092 1401 2158 1419
rect 2092 1351 2108 1401
rect 2142 1351 2158 1401
rect 2092 1329 2158 1351
rect 2092 1283 2108 1329
rect 2142 1283 2158 1329
rect 2092 1257 2158 1283
rect 2092 1215 2108 1257
rect 2142 1215 2158 1257
rect 2092 1185 2158 1215
rect 2092 1147 2108 1185
rect 2142 1147 2158 1185
rect 2092 1113 2158 1147
rect 2092 1079 2108 1113
rect 2142 1079 2158 1113
rect 2092 1045 2158 1079
rect 2092 1007 2108 1045
rect 2142 1007 2158 1045
rect 2092 977 2158 1007
rect 2092 935 2108 977
rect 2142 935 2158 977
rect 2092 909 2158 935
rect 2092 863 2108 909
rect 2142 863 2158 909
rect 2092 841 2158 863
rect 2092 791 2108 841
rect 2142 791 2158 841
rect 2092 773 2158 791
rect 2092 719 2108 773
rect 2142 719 2158 773
rect 2092 705 2158 719
rect 2092 647 2108 705
rect 2142 647 2158 705
rect 2092 637 2158 647
rect 2092 575 2108 637
rect 2142 575 2158 637
rect 2092 569 2158 575
rect 2092 503 2108 569
rect 2142 503 2158 569
rect 2092 501 2158 503
rect 2092 467 2108 501
rect 2142 467 2158 501
rect 2092 465 2158 467
rect 2092 399 2108 465
rect 2142 399 2158 465
rect 2092 393 2158 399
rect 2092 331 2108 393
rect 2142 331 2158 393
rect 2092 321 2158 331
rect 2092 263 2108 321
rect 2142 263 2158 321
rect 34 195 50 249
rect 84 195 100 249
rect 34 177 100 195
rect 34 127 50 177
rect 84 127 100 177
rect 34 100 100 127
rect 2092 249 2158 263
rect 2092 195 2108 249
rect 2142 195 2158 249
rect 2092 177 2158 195
rect 2092 127 2108 177
rect 2142 127 2158 177
rect 2092 100 2158 127
rect 34 84 2158 100
rect 34 50 50 84
rect 84 50 127 84
rect 177 50 195 84
rect 249 50 263 84
rect 321 50 331 84
rect 393 50 399 84
rect 465 50 467 84
rect 501 50 503 84
rect 569 50 575 84
rect 637 50 647 84
rect 705 50 719 84
rect 773 50 791 84
rect 841 50 863 84
rect 909 50 935 84
rect 977 50 1007 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1185 50 1215 84
rect 1257 50 1283 84
rect 1329 50 1351 84
rect 1401 50 1419 84
rect 1473 50 1487 84
rect 1545 50 1555 84
rect 1617 50 1623 84
rect 1689 50 1691 84
rect 1725 50 1727 84
rect 1793 50 1799 84
rect 1861 50 1871 84
rect 1929 50 1943 84
rect 1997 50 2015 84
rect 2065 50 2108 84
rect 2142 50 2158 84
rect 34 34 2158 50
<< viali >>
rect 50 2108 84 2142
rect 143 2108 161 2142
rect 161 2108 177 2142
rect 215 2108 229 2142
rect 229 2108 249 2142
rect 287 2108 297 2142
rect 297 2108 321 2142
rect 359 2108 365 2142
rect 365 2108 393 2142
rect 431 2108 433 2142
rect 433 2108 465 2142
rect 503 2108 535 2142
rect 535 2108 537 2142
rect 575 2108 603 2142
rect 603 2108 609 2142
rect 647 2108 671 2142
rect 671 2108 681 2142
rect 719 2108 739 2142
rect 739 2108 753 2142
rect 791 2108 807 2142
rect 807 2108 825 2142
rect 863 2108 875 2142
rect 875 2108 897 2142
rect 935 2108 943 2142
rect 943 2108 969 2142
rect 1007 2108 1011 2142
rect 1011 2108 1041 2142
rect 1079 2108 1113 2142
rect 1151 2108 1181 2142
rect 1181 2108 1185 2142
rect 1223 2108 1249 2142
rect 1249 2108 1257 2142
rect 1295 2108 1317 2142
rect 1317 2108 1329 2142
rect 1367 2108 1385 2142
rect 1385 2108 1401 2142
rect 1439 2108 1453 2142
rect 1453 2108 1473 2142
rect 1511 2108 1521 2142
rect 1521 2108 1545 2142
rect 1583 2108 1589 2142
rect 1589 2108 1617 2142
rect 1655 2108 1657 2142
rect 1657 2108 1689 2142
rect 1727 2108 1759 2142
rect 1759 2108 1761 2142
rect 1799 2108 1827 2142
rect 1827 2108 1833 2142
rect 1871 2108 1895 2142
rect 1895 2108 1905 2142
rect 1943 2108 1963 2142
rect 1963 2108 1977 2142
rect 2015 2108 2031 2142
rect 2031 2108 2049 2142
rect 2108 2108 2142 2142
rect 50 2031 84 2049
rect 50 2015 84 2031
rect 50 1963 84 1977
rect 50 1943 84 1963
rect 2108 2031 2142 2049
rect 2108 2015 2142 2031
rect 2108 1963 2142 1977
rect 2108 1943 2142 1963
rect 50 1895 84 1905
rect 50 1871 84 1895
rect 50 1827 84 1833
rect 50 1799 84 1827
rect 50 1759 84 1761
rect 50 1727 84 1759
rect 50 1657 84 1689
rect 50 1655 84 1657
rect 50 1589 84 1617
rect 50 1583 84 1589
rect 50 1521 84 1545
rect 50 1511 84 1521
rect 50 1453 84 1473
rect 50 1439 84 1453
rect 50 1385 84 1401
rect 50 1367 84 1385
rect 50 1317 84 1329
rect 50 1295 84 1317
rect 50 1249 84 1257
rect 50 1223 84 1249
rect 50 1181 84 1185
rect 50 1151 84 1181
rect 50 1079 84 1113
rect 50 1011 84 1041
rect 50 1007 84 1011
rect 50 943 84 969
rect 50 935 84 943
rect 50 875 84 897
rect 50 863 84 875
rect 50 807 84 825
rect 50 791 84 807
rect 50 739 84 753
rect 50 719 84 739
rect 50 671 84 681
rect 50 647 84 671
rect 50 603 84 609
rect 50 575 84 603
rect 50 535 84 537
rect 50 503 84 535
rect 50 433 84 465
rect 50 431 84 433
rect 50 365 84 393
rect 50 359 84 365
rect 50 297 84 321
rect 50 287 84 297
rect 276 1882 310 1916
rect 359 1882 365 1916
rect 365 1882 393 1916
rect 431 1882 433 1916
rect 433 1882 465 1916
rect 503 1882 535 1916
rect 535 1882 537 1916
rect 575 1882 603 1916
rect 603 1882 609 1916
rect 647 1882 671 1916
rect 671 1882 681 1916
rect 719 1882 739 1916
rect 739 1882 753 1916
rect 791 1882 807 1916
rect 807 1882 825 1916
rect 863 1882 875 1916
rect 875 1882 897 1916
rect 935 1882 943 1916
rect 943 1882 969 1916
rect 1007 1882 1011 1916
rect 1011 1882 1041 1916
rect 1079 1882 1113 1916
rect 1151 1882 1181 1916
rect 1181 1882 1185 1916
rect 1223 1882 1249 1916
rect 1249 1882 1257 1916
rect 1295 1882 1317 1916
rect 1317 1882 1329 1916
rect 1367 1882 1385 1916
rect 1385 1882 1401 1916
rect 1439 1882 1453 1916
rect 1453 1882 1473 1916
rect 1511 1882 1521 1916
rect 1521 1882 1545 1916
rect 1583 1882 1589 1916
rect 1589 1882 1617 1916
rect 1655 1882 1657 1916
rect 1657 1882 1689 1916
rect 1727 1882 1759 1916
rect 1759 1882 1761 1916
rect 1799 1882 1827 1916
rect 1827 1882 1833 1916
rect 1882 1882 1916 1916
rect 276 1827 310 1833
rect 276 1799 310 1827
rect 276 1759 310 1761
rect 276 1727 310 1759
rect 276 1657 310 1689
rect 276 1655 310 1657
rect 276 1589 310 1617
rect 276 1583 310 1589
rect 276 1521 310 1545
rect 276 1511 310 1521
rect 1882 1827 1916 1833
rect 1882 1799 1916 1827
rect 1882 1759 1916 1761
rect 1882 1727 1916 1759
rect 1882 1657 1916 1689
rect 1882 1655 1916 1657
rect 1882 1589 1916 1617
rect 1882 1583 1916 1589
rect 276 1453 310 1473
rect 276 1439 310 1453
rect 276 1385 310 1401
rect 276 1367 310 1385
rect 276 1317 310 1329
rect 276 1295 310 1317
rect 276 1249 310 1257
rect 276 1223 310 1249
rect 276 1181 310 1185
rect 276 1151 310 1181
rect 276 1079 310 1113
rect 276 1011 310 1041
rect 276 1007 310 1011
rect 276 943 310 969
rect 276 935 310 943
rect 276 875 310 897
rect 276 863 310 875
rect 276 807 310 825
rect 276 791 310 807
rect 276 739 310 753
rect 276 719 310 739
rect 276 671 310 681
rect 276 647 310 671
rect 678 1480 712 1514
rect 755 1480 773 1514
rect 773 1480 789 1514
rect 827 1480 841 1514
rect 841 1480 861 1514
rect 899 1480 909 1514
rect 909 1480 933 1514
rect 971 1480 977 1514
rect 977 1480 1005 1514
rect 1043 1480 1045 1514
rect 1045 1480 1077 1514
rect 1115 1480 1147 1514
rect 1147 1480 1149 1514
rect 1187 1480 1215 1514
rect 1215 1480 1221 1514
rect 1259 1480 1283 1514
rect 1283 1480 1293 1514
rect 1331 1480 1351 1514
rect 1351 1480 1365 1514
rect 1403 1480 1419 1514
rect 1419 1480 1437 1514
rect 1480 1480 1514 1514
rect 678 1419 712 1437
rect 678 1403 712 1419
rect 678 1351 712 1365
rect 678 1331 712 1351
rect 1480 1419 1514 1437
rect 1480 1403 1514 1419
rect 1480 1351 1514 1365
rect 1480 1331 1514 1351
rect 678 1283 712 1293
rect 678 1259 712 1283
rect 678 1215 712 1221
rect 678 1187 712 1215
rect 678 1147 712 1149
rect 678 1115 712 1147
rect 678 1045 712 1077
rect 678 1043 712 1045
rect 678 977 712 1005
rect 678 971 712 977
rect 678 909 712 933
rect 678 899 712 909
rect 935 935 1257 1257
rect 1480 1283 1514 1293
rect 1480 1259 1514 1283
rect 1480 1215 1514 1221
rect 1480 1187 1514 1215
rect 1480 1147 1514 1149
rect 1480 1115 1514 1147
rect 1480 1045 1514 1077
rect 1480 1043 1514 1045
rect 1480 977 1514 1005
rect 1480 971 1514 977
rect 1480 909 1514 933
rect 1480 899 1514 909
rect 678 841 712 861
rect 678 827 712 841
rect 678 773 712 789
rect 678 755 712 773
rect 1480 841 1514 861
rect 1480 827 1514 841
rect 1480 773 1514 789
rect 1480 755 1514 773
rect 678 678 712 712
rect 755 678 773 712
rect 773 678 789 712
rect 827 678 841 712
rect 841 678 861 712
rect 899 678 909 712
rect 909 678 933 712
rect 971 678 977 712
rect 977 678 1005 712
rect 1043 678 1045 712
rect 1045 678 1077 712
rect 1115 678 1147 712
rect 1147 678 1149 712
rect 1187 678 1215 712
rect 1215 678 1221 712
rect 1259 678 1283 712
rect 1283 678 1293 712
rect 1331 678 1351 712
rect 1351 678 1365 712
rect 1403 678 1419 712
rect 1419 678 1437 712
rect 1480 678 1514 712
rect 1882 1521 1916 1545
rect 1882 1511 1916 1521
rect 1882 1453 1916 1473
rect 1882 1439 1916 1453
rect 1882 1385 1916 1401
rect 1882 1367 1916 1385
rect 1882 1317 1916 1329
rect 1882 1295 1916 1317
rect 1882 1249 1916 1257
rect 1882 1223 1916 1249
rect 1882 1181 1916 1185
rect 1882 1151 1916 1181
rect 1882 1079 1916 1113
rect 1882 1011 1916 1041
rect 1882 1007 1916 1011
rect 1882 943 1916 969
rect 1882 935 1916 943
rect 1882 875 1916 897
rect 1882 863 1916 875
rect 1882 807 1916 825
rect 1882 791 1916 807
rect 1882 739 1916 753
rect 1882 719 1916 739
rect 276 603 310 609
rect 276 575 310 603
rect 276 535 310 537
rect 276 503 310 535
rect 276 433 310 465
rect 276 431 310 433
rect 276 365 310 393
rect 276 359 310 365
rect 1882 671 1916 681
rect 1882 647 1916 671
rect 1882 603 1916 609
rect 1882 575 1916 603
rect 1882 535 1916 537
rect 1882 503 1916 535
rect 1882 433 1916 465
rect 1882 431 1916 433
rect 1882 365 1916 393
rect 1882 359 1916 365
rect 276 276 310 310
rect 359 276 365 310
rect 365 276 393 310
rect 431 276 433 310
rect 433 276 465 310
rect 503 276 535 310
rect 535 276 537 310
rect 575 276 603 310
rect 603 276 609 310
rect 647 276 671 310
rect 671 276 681 310
rect 719 276 739 310
rect 739 276 753 310
rect 791 276 807 310
rect 807 276 825 310
rect 863 276 875 310
rect 875 276 897 310
rect 935 276 943 310
rect 943 276 969 310
rect 1007 276 1011 310
rect 1011 276 1041 310
rect 1079 276 1113 310
rect 1151 276 1181 310
rect 1181 276 1185 310
rect 1223 276 1249 310
rect 1249 276 1257 310
rect 1295 276 1317 310
rect 1317 276 1329 310
rect 1367 276 1385 310
rect 1385 276 1401 310
rect 1439 276 1453 310
rect 1453 276 1473 310
rect 1511 276 1521 310
rect 1521 276 1545 310
rect 1583 276 1589 310
rect 1589 276 1617 310
rect 1655 276 1657 310
rect 1657 276 1689 310
rect 1727 276 1759 310
rect 1759 276 1761 310
rect 1799 276 1827 310
rect 1827 276 1833 310
rect 1882 276 1916 310
rect 2108 1895 2142 1905
rect 2108 1871 2142 1895
rect 2108 1827 2142 1833
rect 2108 1799 2142 1827
rect 2108 1759 2142 1761
rect 2108 1727 2142 1759
rect 2108 1657 2142 1689
rect 2108 1655 2142 1657
rect 2108 1589 2142 1617
rect 2108 1583 2142 1589
rect 2108 1521 2142 1545
rect 2108 1511 2142 1521
rect 2108 1453 2142 1473
rect 2108 1439 2142 1453
rect 2108 1385 2142 1401
rect 2108 1367 2142 1385
rect 2108 1317 2142 1329
rect 2108 1295 2142 1317
rect 2108 1249 2142 1257
rect 2108 1223 2142 1249
rect 2108 1181 2142 1185
rect 2108 1151 2142 1181
rect 2108 1079 2142 1113
rect 2108 1011 2142 1041
rect 2108 1007 2142 1011
rect 2108 943 2142 969
rect 2108 935 2142 943
rect 2108 875 2142 897
rect 2108 863 2142 875
rect 2108 807 2142 825
rect 2108 791 2142 807
rect 2108 739 2142 753
rect 2108 719 2142 739
rect 2108 671 2142 681
rect 2108 647 2142 671
rect 2108 603 2142 609
rect 2108 575 2142 603
rect 2108 535 2142 537
rect 2108 503 2142 535
rect 2108 433 2142 465
rect 2108 431 2142 433
rect 2108 365 2142 393
rect 2108 359 2142 365
rect 2108 297 2142 321
rect 2108 287 2142 297
rect 50 229 84 249
rect 50 215 84 229
rect 50 161 84 177
rect 50 143 84 161
rect 2108 229 2142 249
rect 2108 215 2142 229
rect 2108 161 2142 177
rect 2108 143 2142 161
rect 50 50 84 84
rect 143 50 161 84
rect 161 50 177 84
rect 215 50 229 84
rect 229 50 249 84
rect 287 50 297 84
rect 297 50 321 84
rect 359 50 365 84
rect 365 50 393 84
rect 431 50 433 84
rect 433 50 465 84
rect 503 50 535 84
rect 535 50 537 84
rect 575 50 603 84
rect 603 50 609 84
rect 647 50 671 84
rect 671 50 681 84
rect 719 50 739 84
rect 739 50 753 84
rect 791 50 807 84
rect 807 50 825 84
rect 863 50 875 84
rect 875 50 897 84
rect 935 50 943 84
rect 943 50 969 84
rect 1007 50 1011 84
rect 1011 50 1041 84
rect 1079 50 1113 84
rect 1151 50 1181 84
rect 1181 50 1185 84
rect 1223 50 1249 84
rect 1249 50 1257 84
rect 1295 50 1317 84
rect 1317 50 1329 84
rect 1367 50 1385 84
rect 1385 50 1401 84
rect 1439 50 1453 84
rect 1453 50 1473 84
rect 1511 50 1521 84
rect 1521 50 1545 84
rect 1583 50 1589 84
rect 1589 50 1617 84
rect 1655 50 1657 84
rect 1657 50 1689 84
rect 1727 50 1759 84
rect 1759 50 1761 84
rect 1799 50 1827 84
rect 1827 50 1833 84
rect 1871 50 1895 84
rect 1895 50 1905 84
rect 1943 50 1963 84
rect 1963 50 1977 84
rect 2015 50 2031 84
rect 2031 50 2049 84
rect 2108 50 2142 84
<< metal1 >>
rect 38 2142 2154 2154
rect 38 2108 50 2142
rect 84 2108 143 2142
rect 177 2108 215 2142
rect 249 2108 287 2142
rect 321 2108 359 2142
rect 393 2108 431 2142
rect 465 2108 503 2142
rect 537 2108 575 2142
rect 609 2108 647 2142
rect 681 2108 719 2142
rect 753 2108 791 2142
rect 825 2108 863 2142
rect 897 2108 935 2142
rect 969 2108 1007 2142
rect 1041 2108 1079 2142
rect 1113 2108 1151 2142
rect 1185 2108 1223 2142
rect 1257 2108 1295 2142
rect 1329 2108 1367 2142
rect 1401 2108 1439 2142
rect 1473 2108 1511 2142
rect 1545 2108 1583 2142
rect 1617 2108 1655 2142
rect 1689 2108 1727 2142
rect 1761 2108 1799 2142
rect 1833 2108 1871 2142
rect 1905 2108 1943 2142
rect 1977 2108 2015 2142
rect 2049 2108 2108 2142
rect 2142 2108 2154 2142
rect 38 2096 2154 2108
rect 38 2049 96 2096
rect 38 2015 50 2049
rect 84 2015 96 2049
rect 38 1977 96 2015
rect 38 1943 50 1977
rect 84 1943 96 1977
rect 38 1905 96 1943
rect 2096 2049 2154 2096
rect 2096 2015 2108 2049
rect 2142 2015 2154 2049
rect 2096 1977 2154 2015
rect 2096 1943 2108 1977
rect 2142 1943 2154 1977
rect 38 1871 50 1905
rect 84 1871 96 1905
rect 38 1833 96 1871
rect 38 1799 50 1833
rect 84 1799 96 1833
rect 38 1761 96 1799
rect 38 1727 50 1761
rect 84 1727 96 1761
rect 38 1689 96 1727
rect 38 1655 50 1689
rect 84 1655 96 1689
rect 38 1617 96 1655
rect 38 1583 50 1617
rect 84 1583 96 1617
rect 38 1545 96 1583
rect 38 1511 50 1545
rect 84 1511 96 1545
rect 38 1473 96 1511
rect 38 1439 50 1473
rect 84 1439 96 1473
rect 38 1401 96 1439
rect 38 1367 50 1401
rect 84 1367 96 1401
rect 38 1329 96 1367
rect 38 1295 50 1329
rect 84 1295 96 1329
rect 38 1257 96 1295
rect 38 1223 50 1257
rect 84 1223 96 1257
rect 38 1185 96 1223
rect 38 1151 50 1185
rect 84 1151 96 1185
rect 38 1113 96 1151
rect 38 1079 50 1113
rect 84 1079 96 1113
rect 38 1041 96 1079
rect 38 1007 50 1041
rect 84 1007 96 1041
rect 38 969 96 1007
rect 38 935 50 969
rect 84 935 96 969
rect 38 897 96 935
rect 38 863 50 897
rect 84 863 96 897
rect 38 825 96 863
rect 38 791 50 825
rect 84 791 96 825
rect 38 753 96 791
rect 38 719 50 753
rect 84 719 96 753
rect 38 681 96 719
rect 38 647 50 681
rect 84 647 96 681
rect 38 609 96 647
rect 38 575 50 609
rect 84 575 96 609
rect 38 537 96 575
rect 38 503 50 537
rect 84 503 96 537
rect 38 465 96 503
rect 38 431 50 465
rect 84 431 96 465
rect 38 393 96 431
rect 38 359 50 393
rect 84 359 96 393
rect 38 321 96 359
rect 38 287 50 321
rect 84 287 96 321
rect 38 249 96 287
rect 264 1916 1928 1928
rect 264 1882 276 1916
rect 310 1882 359 1916
rect 393 1882 431 1916
rect 465 1882 503 1916
rect 537 1882 575 1916
rect 609 1882 647 1916
rect 681 1882 719 1916
rect 753 1882 791 1916
rect 825 1882 863 1916
rect 897 1882 935 1916
rect 969 1882 1007 1916
rect 1041 1882 1079 1916
rect 1113 1882 1151 1916
rect 1185 1882 1223 1916
rect 1257 1882 1295 1916
rect 1329 1882 1367 1916
rect 1401 1882 1439 1916
rect 1473 1882 1511 1916
rect 1545 1882 1583 1916
rect 1617 1882 1655 1916
rect 1689 1882 1727 1916
rect 1761 1882 1799 1916
rect 1833 1882 1882 1916
rect 1916 1882 1928 1916
rect 264 1870 1928 1882
rect 264 1833 322 1870
rect 264 1799 276 1833
rect 310 1799 322 1833
rect 264 1761 322 1799
rect 264 1727 276 1761
rect 310 1727 322 1761
rect 264 1689 322 1727
rect 264 1655 276 1689
rect 310 1655 322 1689
rect 264 1617 322 1655
rect 264 1583 276 1617
rect 310 1583 322 1617
rect 264 1545 322 1583
rect 264 1511 276 1545
rect 310 1511 322 1545
rect 1870 1833 1928 1870
rect 1870 1799 1882 1833
rect 1916 1799 1928 1833
rect 1870 1761 1928 1799
rect 1870 1727 1882 1761
rect 1916 1727 1928 1761
rect 1870 1689 1928 1727
rect 1870 1655 1882 1689
rect 1916 1655 1928 1689
rect 1870 1617 1928 1655
rect 1870 1583 1882 1617
rect 1916 1583 1928 1617
rect 1870 1545 1928 1583
rect 264 1473 322 1511
rect 264 1439 276 1473
rect 310 1439 322 1473
rect 264 1401 322 1439
rect 264 1367 276 1401
rect 310 1367 322 1401
rect 264 1329 322 1367
rect 264 1295 276 1329
rect 310 1295 322 1329
rect 264 1257 322 1295
rect 264 1223 276 1257
rect 310 1223 322 1257
rect 264 1185 322 1223
rect 264 1151 276 1185
rect 310 1151 322 1185
rect 264 1113 322 1151
rect 264 1079 276 1113
rect 310 1079 322 1113
rect 264 1041 322 1079
rect 264 1007 276 1041
rect 310 1007 322 1041
rect 264 969 322 1007
rect 264 935 276 969
rect 310 935 322 969
rect 264 897 322 935
rect 264 863 276 897
rect 310 863 322 897
rect 264 825 322 863
rect 264 791 276 825
rect 310 791 322 825
rect 264 753 322 791
rect 264 719 276 753
rect 310 719 322 753
rect 264 681 322 719
rect 264 647 276 681
rect 310 647 322 681
rect 666 1514 1526 1526
rect 666 1480 678 1514
rect 712 1480 755 1514
rect 789 1480 827 1514
rect 861 1480 899 1514
rect 933 1480 971 1514
rect 1005 1480 1043 1514
rect 1077 1480 1115 1514
rect 1149 1480 1187 1514
rect 1221 1480 1259 1514
rect 1293 1480 1331 1514
rect 1365 1480 1403 1514
rect 1437 1480 1480 1514
rect 1514 1480 1526 1514
rect 666 1468 1526 1480
rect 666 1437 724 1468
rect 666 1403 678 1437
rect 712 1403 724 1437
rect 666 1365 724 1403
rect 666 1331 678 1365
rect 712 1331 724 1365
rect 666 1293 724 1331
rect 666 1259 678 1293
rect 712 1259 724 1293
rect 1468 1437 1526 1468
rect 1468 1403 1480 1437
rect 1514 1403 1526 1437
rect 1468 1365 1526 1403
rect 1468 1331 1480 1365
rect 1514 1331 1526 1365
rect 1468 1293 1526 1331
rect 666 1221 724 1259
rect 666 1187 678 1221
rect 712 1187 724 1221
rect 666 1149 724 1187
rect 666 1115 678 1149
rect 712 1115 724 1149
rect 666 1077 724 1115
rect 666 1043 678 1077
rect 712 1043 724 1077
rect 666 1005 724 1043
rect 666 971 678 1005
rect 712 971 724 1005
rect 666 933 724 971
rect 666 899 678 933
rect 712 899 724 933
rect 923 1257 1269 1269
rect 923 935 935 1257
rect 1257 935 1269 1257
rect 923 923 1269 935
rect 1468 1259 1480 1293
rect 1514 1259 1526 1293
rect 1468 1221 1526 1259
rect 1468 1187 1480 1221
rect 1514 1187 1526 1221
rect 1468 1149 1526 1187
rect 1468 1115 1480 1149
rect 1514 1115 1526 1149
rect 1468 1077 1526 1115
rect 1468 1043 1480 1077
rect 1514 1043 1526 1077
rect 1468 1005 1526 1043
rect 1468 971 1480 1005
rect 1514 971 1526 1005
rect 1468 933 1526 971
rect 666 861 724 899
rect 666 827 678 861
rect 712 827 724 861
rect 666 789 724 827
rect 666 755 678 789
rect 712 755 724 789
rect 666 724 724 755
rect 1468 899 1480 933
rect 1514 899 1526 933
rect 1468 861 1526 899
rect 1468 827 1480 861
rect 1514 827 1526 861
rect 1468 789 1526 827
rect 1468 755 1480 789
rect 1514 755 1526 789
rect 1468 724 1526 755
rect 666 712 1526 724
rect 666 678 678 712
rect 712 678 755 712
rect 789 678 827 712
rect 861 678 899 712
rect 933 678 971 712
rect 1005 678 1043 712
rect 1077 678 1115 712
rect 1149 678 1187 712
rect 1221 678 1259 712
rect 1293 678 1331 712
rect 1365 678 1403 712
rect 1437 678 1480 712
rect 1514 678 1526 712
rect 666 666 1526 678
rect 1870 1511 1882 1545
rect 1916 1511 1928 1545
rect 1870 1473 1928 1511
rect 1870 1439 1882 1473
rect 1916 1439 1928 1473
rect 1870 1401 1928 1439
rect 1870 1367 1882 1401
rect 1916 1367 1928 1401
rect 1870 1329 1928 1367
rect 1870 1295 1882 1329
rect 1916 1295 1928 1329
rect 1870 1257 1928 1295
rect 1870 1223 1882 1257
rect 1916 1223 1928 1257
rect 1870 1185 1928 1223
rect 1870 1151 1882 1185
rect 1916 1151 1928 1185
rect 1870 1113 1928 1151
rect 1870 1079 1882 1113
rect 1916 1079 1928 1113
rect 1870 1041 1928 1079
rect 1870 1007 1882 1041
rect 1916 1007 1928 1041
rect 1870 969 1928 1007
rect 1870 935 1882 969
rect 1916 935 1928 969
rect 1870 897 1928 935
rect 1870 863 1882 897
rect 1916 863 1928 897
rect 1870 825 1928 863
rect 1870 791 1882 825
rect 1916 791 1928 825
rect 1870 753 1928 791
rect 1870 719 1882 753
rect 1916 719 1928 753
rect 1870 681 1928 719
rect 264 609 322 647
rect 264 575 276 609
rect 310 575 322 609
rect 264 537 322 575
rect 264 503 276 537
rect 310 503 322 537
rect 264 465 322 503
rect 264 431 276 465
rect 310 431 322 465
rect 264 393 322 431
rect 264 359 276 393
rect 310 359 322 393
rect 264 322 322 359
rect 1870 647 1882 681
rect 1916 647 1928 681
rect 1870 609 1928 647
rect 1870 575 1882 609
rect 1916 575 1928 609
rect 1870 537 1928 575
rect 1870 503 1882 537
rect 1916 503 1928 537
rect 1870 465 1928 503
rect 1870 431 1882 465
rect 1916 431 1928 465
rect 1870 393 1928 431
rect 1870 359 1882 393
rect 1916 359 1928 393
rect 1870 322 1928 359
rect 264 310 1928 322
rect 264 276 276 310
rect 310 276 359 310
rect 393 276 431 310
rect 465 276 503 310
rect 537 276 575 310
rect 609 276 647 310
rect 681 276 719 310
rect 753 276 791 310
rect 825 276 863 310
rect 897 276 935 310
rect 969 276 1007 310
rect 1041 276 1079 310
rect 1113 276 1151 310
rect 1185 276 1223 310
rect 1257 276 1295 310
rect 1329 276 1367 310
rect 1401 276 1439 310
rect 1473 276 1511 310
rect 1545 276 1583 310
rect 1617 276 1655 310
rect 1689 276 1727 310
rect 1761 276 1799 310
rect 1833 276 1882 310
rect 1916 276 1928 310
rect 264 264 1928 276
rect 2096 1905 2154 1943
rect 2096 1871 2108 1905
rect 2142 1871 2154 1905
rect 2096 1833 2154 1871
rect 2096 1799 2108 1833
rect 2142 1799 2154 1833
rect 2096 1761 2154 1799
rect 2096 1727 2108 1761
rect 2142 1727 2154 1761
rect 2096 1689 2154 1727
rect 2096 1655 2108 1689
rect 2142 1655 2154 1689
rect 2096 1617 2154 1655
rect 2096 1583 2108 1617
rect 2142 1583 2154 1617
rect 2096 1545 2154 1583
rect 2096 1511 2108 1545
rect 2142 1511 2154 1545
rect 2096 1473 2154 1511
rect 2096 1439 2108 1473
rect 2142 1439 2154 1473
rect 2096 1401 2154 1439
rect 2096 1367 2108 1401
rect 2142 1367 2154 1401
rect 2096 1329 2154 1367
rect 2096 1295 2108 1329
rect 2142 1295 2154 1329
rect 2096 1257 2154 1295
rect 2096 1223 2108 1257
rect 2142 1223 2154 1257
rect 2096 1185 2154 1223
rect 2096 1151 2108 1185
rect 2142 1151 2154 1185
rect 2096 1113 2154 1151
rect 2096 1079 2108 1113
rect 2142 1079 2154 1113
rect 2096 1041 2154 1079
rect 2096 1007 2108 1041
rect 2142 1007 2154 1041
rect 2096 969 2154 1007
rect 2096 935 2108 969
rect 2142 935 2154 969
rect 2096 897 2154 935
rect 2096 863 2108 897
rect 2142 863 2154 897
rect 2096 825 2154 863
rect 2096 791 2108 825
rect 2142 791 2154 825
rect 2096 753 2154 791
rect 2096 719 2108 753
rect 2142 719 2154 753
rect 2096 681 2154 719
rect 2096 647 2108 681
rect 2142 647 2154 681
rect 2096 609 2154 647
rect 2096 575 2108 609
rect 2142 575 2154 609
rect 2096 537 2154 575
rect 2096 503 2108 537
rect 2142 503 2154 537
rect 2096 465 2154 503
rect 2096 431 2108 465
rect 2142 431 2154 465
rect 2096 393 2154 431
rect 2096 359 2108 393
rect 2142 359 2154 393
rect 2096 321 2154 359
rect 2096 287 2108 321
rect 2142 287 2154 321
rect 38 215 50 249
rect 84 215 96 249
rect 38 177 96 215
rect 38 143 50 177
rect 84 143 96 177
rect 38 96 96 143
rect 2096 249 2154 287
rect 2096 215 2108 249
rect 2142 215 2154 249
rect 2096 177 2154 215
rect 2096 143 2108 177
rect 2142 143 2154 177
rect 2096 96 2154 143
rect 38 84 2154 96
rect 38 50 50 84
rect 84 50 143 84
rect 177 50 215 84
rect 249 50 287 84
rect 321 50 359 84
rect 393 50 431 84
rect 465 50 503 84
rect 537 50 575 84
rect 609 50 647 84
rect 681 50 719 84
rect 753 50 791 84
rect 825 50 863 84
rect 897 50 935 84
rect 969 50 1007 84
rect 1041 50 1079 84
rect 1113 50 1151 84
rect 1185 50 1223 84
rect 1257 50 1295 84
rect 1329 50 1367 84
rect 1401 50 1439 84
rect 1473 50 1511 84
rect 1545 50 1583 84
rect 1617 50 1655 84
rect 1689 50 1727 84
rect 1761 50 1799 84
rect 1833 50 1871 84
rect 1905 50 1943 84
rect 1977 50 2015 84
rect 2049 50 2108 84
rect 2142 50 2154 84
rect 38 38 2154 50
<< properties >>
string GDS_END 8885666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8840726
string path 7.850 12.350 7.850 46.950 46.950 46.950 46.950 7.850 3.350 7.850 
<< end >>
