magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -79 -26 935 110
<< mvnmos >>
rect 0 0 400 84
rect 456 0 856 84
<< mvndiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 400 46 456 84
rect 400 12 411 46
rect 445 12 456 46
rect 400 0 456 12
rect 856 46 909 84
rect 856 12 867 46
rect 901 12 909 46
rect 856 0 909 12
<< mvndiffc >>
rect -45 12 -11 46
rect 411 12 445 46
rect 867 12 901 46
<< poly >>
rect 0 84 400 116
rect 456 84 856 116
rect 0 -32 400 0
rect 456 -32 856 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 411 46 445 62
rect 411 -4 445 12
rect 867 46 901 62
rect 867 -4 901 12
use DFL1sd2_CDNS_52468879185467  DFL1sd2_CDNS_52468879185467_0
timestamp 1707688321
transform 1 0 400 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185271  DFL1sd_CDNS_52468879185271_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185271  DFL1sd_CDNS_52468879185271_1
timestamp 1707688321
transform 1 0 856 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 428 29 428 29 0 FreeSans 300 0 0 0 D
flabel comment s 884 29 884 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 89250856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89249472
<< end >>
