magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -1274 4473 -131 4708
rect -1274 4163 -1106 4473
rect -1869 4116 -1106 4163
rect -299 4116 -131 4473
rect -1869 4007 -131 4116
rect -1869 3995 -1106 4007
rect -1869 3588 -1701 3995
rect -837 3588 -328 3634
rect -1869 3466 -328 3588
rect -1869 3281 -479 3466
rect -647 3274 -479 3281
rect -299 3274 -131 4007
rect -647 3106 -131 3274
rect 853 2048 1769 2216
rect 853 1461 930 2048
rect 1601 1461 1769 2048
rect 853 1395 1769 1461
rect 841 805 1769 871
rect 841 218 1009 805
rect 1601 218 1769 805
rect 841 50 1769 218
<< pwell >>
rect -71 4581 1678 4667
rect -71 2369 15 4581
rect 920 4544 1190 4581
rect 920 2369 1190 2406
rect 1592 2369 1678 4581
rect -71 2362 1678 2369
rect -71 2283 1915 2362
rect -71 -17 15 2283
rect 695 2276 1915 2283
rect 695 1336 781 2276
rect 695 1335 791 1336
rect 1829 1335 1915 2276
rect 695 1250 1915 1335
rect 695 1016 791 1250
rect 1829 1016 1915 1250
rect 695 931 1915 1016
rect 695 930 791 931
rect 695 -10 781 930
rect 1829 -10 1915 931
rect 695 -17 1915 -10
rect -71 -103 1915 -17
<< mvpsubdiff >>
rect -45 4607 88 4641
rect 122 4607 156 4641
rect 190 4607 224 4641
rect 258 4607 292 4641
rect 326 4607 360 4641
rect 394 4607 428 4641
rect 462 4607 496 4641
rect 530 4607 564 4641
rect 598 4607 632 4641
rect 666 4607 700 4641
rect 734 4607 768 4641
rect 802 4607 836 4641
rect 870 4607 904 4641
rect 938 4607 972 4641
rect 1006 4607 1040 4641
rect 1074 4607 1108 4641
rect 1142 4607 1176 4641
rect 1210 4607 1244 4641
rect 1278 4607 1312 4641
rect 1346 4607 1380 4641
rect 1414 4607 1448 4641
rect 1482 4607 1516 4641
rect 1550 4607 1584 4641
rect -45 4539 -11 4573
rect -45 4471 -11 4505
rect 946 4570 1164 4607
rect 1618 4553 1652 4641
rect -45 4403 -11 4437
rect -45 4335 -11 4369
rect -45 4267 -11 4301
rect -45 4199 -11 4233
rect -45 4131 -11 4165
rect -45 4063 -11 4097
rect -45 3995 -11 4029
rect -45 3927 -11 3961
rect -45 3859 -11 3893
rect -45 3791 -11 3825
rect -45 3723 -11 3757
rect -45 3655 -11 3689
rect -45 3587 -11 3621
rect -45 3519 -11 3553
rect -45 3451 -11 3485
rect -45 3383 -11 3417
rect -45 3315 -11 3349
rect -45 3247 -11 3281
rect -45 3179 -11 3213
rect -45 3111 -11 3145
rect -45 3043 -11 3077
rect -45 2975 -11 3009
rect -45 2907 -11 2941
rect -45 2839 -11 2873
rect -45 2771 -11 2805
rect -45 2703 -11 2737
rect -45 2635 -11 2669
rect -45 2567 -11 2601
rect -45 2343 -11 2533
rect 1618 4485 1652 4519
rect 1618 4417 1652 4451
rect 1618 4349 1652 4383
rect 1618 4281 1652 4315
rect 1618 4213 1652 4247
rect 1618 4145 1652 4179
rect 1618 4077 1652 4111
rect 1618 4009 1652 4043
rect 1618 3941 1652 3975
rect 1618 3873 1652 3907
rect 1618 3805 1652 3839
rect 1618 3737 1652 3771
rect 1618 3669 1652 3703
rect 1618 3601 1652 3635
rect 1618 3533 1652 3567
rect 1618 3465 1652 3499
rect 1618 3397 1652 3431
rect 1618 3329 1652 3363
rect 1618 3261 1652 3295
rect 1618 3193 1652 3227
rect 1618 3125 1652 3159
rect 1618 3057 1652 3091
rect 1618 2989 1652 3023
rect 1618 2921 1652 2955
rect 1618 2853 1652 2887
rect 1618 2785 1652 2819
rect 1618 2717 1652 2751
rect 1618 2649 1652 2683
rect 1618 2581 1652 2615
rect 1618 2513 1652 2547
rect 946 2343 1164 2380
rect 1618 2445 1652 2479
rect 1618 2377 1652 2411
rect -45 2309 88 2343
rect 122 2309 156 2343
rect 190 2309 224 2343
rect 258 2309 292 2343
rect 326 2309 360 2343
rect 394 2309 428 2343
rect 462 2309 496 2343
rect 530 2309 564 2343
rect 598 2309 632 2343
rect 666 2309 700 2343
rect 734 2309 768 2343
rect 802 2309 836 2343
rect 870 2309 904 2343
rect 938 2309 972 2343
rect 1006 2309 1040 2343
rect 1074 2309 1108 2343
rect 1142 2309 1176 2343
rect 1210 2309 1244 2343
rect 1278 2309 1312 2343
rect 1346 2309 1380 2343
rect 1414 2309 1448 2343
rect 1482 2309 1516 2343
rect 1550 2336 1652 2343
rect 1550 2309 1686 2336
rect -45 2303 -11 2309
rect -45 2235 -11 2269
rect -45 2167 -11 2201
rect -45 2099 -11 2133
rect -45 2031 -11 2065
rect -45 1963 -11 1997
rect -45 1895 -11 1929
rect -45 1827 -11 1861
rect -45 1759 -11 1793
rect -45 1691 -11 1725
rect -45 1623 -11 1657
rect 721 2302 1686 2309
rect 1720 2302 1754 2336
rect 1788 2302 1889 2336
rect 721 2275 755 2302
rect 721 2207 755 2241
rect 721 2139 755 2173
rect 1855 2240 1889 2302
rect 1855 2169 1889 2206
rect 721 2071 755 2105
rect 721 2003 755 2037
rect 721 1935 755 1969
rect 721 1867 755 1901
rect 721 1799 755 1833
rect 721 1731 755 1765
rect 721 1663 755 1697
rect -45 1555 -11 1589
rect 721 1595 755 1629
rect -45 1487 -11 1521
rect 721 1527 755 1561
rect -45 1419 -11 1453
rect 721 1459 755 1493
rect 1855 2098 1889 2135
rect 1855 2027 1889 2064
rect 1855 1956 1889 1993
rect 1855 1885 1889 1922
rect 1855 1814 1889 1851
rect 1855 1743 1889 1780
rect 1855 1672 1889 1709
rect 1855 1601 1889 1638
rect 1855 1530 1889 1567
rect 1855 1459 1889 1496
rect -45 1351 -11 1385
rect -45 1283 -11 1317
rect -45 1215 -11 1249
rect -45 1147 -11 1181
rect -45 1079 -11 1113
rect -45 1011 -11 1045
rect -45 943 -11 977
rect -45 875 -11 909
rect -45 807 -11 841
rect -45 739 -11 773
rect 721 1391 755 1425
rect 1855 1388 1889 1425
rect 721 1323 755 1357
rect 755 1309 765 1310
rect 1855 1309 1889 1354
rect 755 1289 1889 1309
rect 721 1276 1889 1289
rect 721 1255 765 1276
rect 755 1221 765 1255
rect 721 1187 765 1221
rect 755 1153 765 1187
rect 721 1119 765 1153
rect 755 1085 765 1119
rect 721 1051 765 1085
rect 755 1017 765 1051
rect 721 990 765 1017
rect 1855 990 1889 1276
rect 721 983 1889 990
rect 755 957 1889 983
rect 755 956 765 957
rect 721 915 755 949
rect 1855 948 1889 957
rect 721 847 755 881
rect 1855 875 1889 914
rect 721 779 755 813
rect -45 671 -11 705
rect 721 711 755 745
rect -45 603 -11 637
rect -45 535 -11 569
rect -45 467 -11 501
rect -45 399 -11 433
rect -45 331 -11 365
rect -45 263 -11 297
rect -45 195 -11 229
rect -45 127 -11 161
rect -45 59 -11 93
rect -45 -9 -11 25
rect 721 643 755 677
rect 721 575 755 609
rect 721 507 755 541
rect 721 439 755 473
rect 721 371 755 405
rect 721 303 755 337
rect 721 235 755 269
rect 721 167 755 201
rect 721 99 755 133
rect 1855 802 1889 841
rect 1855 729 1889 768
rect 1855 656 1889 695
rect 1855 583 1889 622
rect 1855 511 1889 549
rect 1855 439 1889 477
rect 1855 367 1889 405
rect 1855 295 1889 333
rect 1855 223 1889 261
rect 1855 151 1889 189
rect 721 -36 755 65
rect 1855 79 1889 117
rect 1855 7 1889 45
rect 1855 -36 1889 -27
rect -45 -77 75 -43
rect 109 -77 143 -43
rect 177 -77 211 -43
rect 245 -77 279 -43
rect 313 -77 347 -43
rect 381 -77 415 -43
rect 449 -77 483 -43
rect 517 -77 551 -43
rect 585 -77 619 -43
rect 653 -77 687 -43
rect 721 -70 789 -36
rect 823 -70 857 -36
rect 891 -70 925 -36
rect 959 -70 993 -36
rect 1027 -70 1061 -36
rect 1095 -70 1129 -36
rect 1163 -70 1197 -36
rect 1231 -70 1265 -36
rect 1299 -70 1333 -36
rect 1367 -70 1401 -36
rect 1435 -70 1469 -36
rect 1503 -70 1537 -36
rect 1571 -70 1605 -36
rect 1639 -70 1673 -36
rect 1707 -70 1741 -36
rect 1775 -70 1889 -36
rect 721 -77 1889 -70
<< mvnsubdiff >>
rect -1207 4607 -1082 4641
rect -1048 4607 -1014 4641
rect -980 4607 -946 4641
rect -912 4607 -878 4641
rect -844 4607 -810 4641
rect -776 4607 -742 4641
rect -708 4607 -674 4641
rect -640 4607 -606 4641
rect -572 4607 -538 4641
rect -504 4607 -470 4641
rect -436 4607 -402 4641
rect -368 4607 -334 4641
rect -300 4607 -266 4641
rect -1207 4539 -1173 4573
rect -1207 4471 -1173 4505
rect -1207 4403 -1173 4437
rect -232 4532 -198 4641
rect -232 4464 -198 4498
rect -1207 4335 -1173 4369
rect -1207 4267 -1173 4301
rect -1207 4199 -1173 4233
rect -1802 4062 -1717 4096
rect -1683 4062 -1649 4096
rect -1615 4062 -1581 4096
rect -1547 4062 -1513 4096
rect -1479 4062 -1445 4096
rect -1411 4062 -1377 4096
rect -1343 4062 -1309 4096
rect -1275 4062 -1241 4096
rect -1207 4062 -1173 4165
rect -232 4396 -198 4430
rect -232 4328 -198 4362
rect -232 4260 -198 4294
rect -232 4192 -198 4226
rect -232 4124 -198 4158
rect -1802 4028 -1768 4062
rect -232 4056 -198 4090
rect -1802 3960 -1768 3994
rect -232 3988 -198 4022
rect -1802 3892 -1768 3926
rect -1802 3824 -1768 3858
rect -1802 3756 -1768 3790
rect -1802 3688 -1768 3722
rect -1802 3620 -1768 3654
rect -232 3920 -198 3954
rect -232 3852 -198 3886
rect -232 3784 -198 3818
rect -232 3716 -198 3750
rect -1802 3552 -1768 3586
rect -1802 3484 -1768 3518
rect -232 3581 -198 3682
rect -232 3513 -198 3547
rect -1802 3416 -1768 3450
rect -232 3445 -198 3479
rect -1802 3348 -1734 3382
rect -1700 3348 -1666 3382
rect -1632 3348 -1598 3382
rect -1564 3348 -1530 3382
rect -1496 3348 -1462 3382
rect -1428 3348 -1394 3382
rect -1360 3348 -1326 3382
rect -1292 3348 -1258 3382
rect -1224 3348 -1190 3382
rect -1156 3348 -1122 3382
rect -1088 3348 -1054 3382
rect -1020 3348 -986 3382
rect -952 3348 -918 3382
rect -884 3348 -850 3382
rect -816 3348 -782 3382
rect -748 3348 -714 3382
rect -680 3348 -546 3382
rect -580 3343 -546 3348
rect -580 3275 -546 3309
rect -580 3173 -546 3241
rect -232 3377 -198 3411
rect -232 3309 -198 3343
rect -232 3241 -198 3275
rect -512 3173 -478 3207
rect -444 3173 -410 3207
rect -376 3173 -342 3207
rect -308 3173 -198 3207
rect 919 2115 953 2149
rect 987 2115 1021 2149
rect 1055 2115 1089 2149
rect 1123 2115 1157 2149
rect 1191 2115 1225 2149
rect 1259 2115 1293 2149
rect 1327 2115 1361 2149
rect 1395 2115 1429 2149
rect 1463 2115 1497 2149
rect 1531 2115 1565 2149
rect 1599 2115 1702 2149
rect 1668 2047 1702 2081
rect 1668 1979 1702 2013
rect 1668 1911 1702 1945
rect 1668 1843 1702 1877
rect 1668 1775 1702 1809
rect 1668 1707 1702 1741
rect 1668 1639 1702 1673
rect 1668 1571 1702 1605
rect 1668 1461 1702 1537
rect 908 771 942 805
rect 908 703 942 737
rect 908 635 942 669
rect 908 567 942 601
rect 908 499 942 533
rect 908 431 942 465
rect 908 363 942 397
rect 908 295 942 329
rect 908 117 942 261
rect 1668 729 1702 805
rect 1668 661 1702 695
rect 1668 593 1702 627
rect 1668 525 1702 559
rect 1668 457 1702 491
rect 1668 389 1702 423
rect 1668 321 1702 355
rect 1668 253 1702 287
rect 1668 185 1702 219
rect 976 117 1010 151
rect 1044 117 1078 151
rect 1112 117 1146 151
rect 1180 117 1214 151
rect 1248 117 1282 151
rect 1316 117 1350 151
rect 1384 117 1418 151
rect 1452 117 1486 151
rect 1520 117 1554 151
rect 1588 117 1702 151
<< mvpsubdiffcont >>
rect 88 4607 122 4641
rect 156 4607 190 4641
rect 224 4607 258 4641
rect 292 4607 326 4641
rect 360 4607 394 4641
rect 428 4607 462 4641
rect 496 4607 530 4641
rect 564 4607 598 4641
rect 632 4607 666 4641
rect 700 4607 734 4641
rect 768 4607 802 4641
rect 836 4607 870 4641
rect 904 4607 938 4641
rect 972 4607 1006 4641
rect 1040 4607 1074 4641
rect 1108 4607 1142 4641
rect 1176 4607 1210 4641
rect 1244 4607 1278 4641
rect 1312 4607 1346 4641
rect 1380 4607 1414 4641
rect 1448 4607 1482 4641
rect 1516 4607 1550 4641
rect 1584 4607 1618 4641
rect -45 4573 -11 4607
rect -45 4505 -11 4539
rect 1618 4519 1652 4553
rect -45 4437 -11 4471
rect -45 4369 -11 4403
rect -45 4301 -11 4335
rect -45 4233 -11 4267
rect -45 4165 -11 4199
rect -45 4097 -11 4131
rect -45 4029 -11 4063
rect -45 3961 -11 3995
rect -45 3893 -11 3927
rect -45 3825 -11 3859
rect -45 3757 -11 3791
rect -45 3689 -11 3723
rect -45 3621 -11 3655
rect -45 3553 -11 3587
rect -45 3485 -11 3519
rect -45 3417 -11 3451
rect -45 3349 -11 3383
rect -45 3281 -11 3315
rect -45 3213 -11 3247
rect -45 3145 -11 3179
rect -45 3077 -11 3111
rect -45 3009 -11 3043
rect -45 2941 -11 2975
rect -45 2873 -11 2907
rect -45 2805 -11 2839
rect -45 2737 -11 2771
rect -45 2669 -11 2703
rect -45 2601 -11 2635
rect -45 2533 -11 2567
rect 1618 4451 1652 4485
rect 1618 4383 1652 4417
rect 1618 4315 1652 4349
rect 1618 4247 1652 4281
rect 1618 4179 1652 4213
rect 1618 4111 1652 4145
rect 1618 4043 1652 4077
rect 1618 3975 1652 4009
rect 1618 3907 1652 3941
rect 1618 3839 1652 3873
rect 1618 3771 1652 3805
rect 1618 3703 1652 3737
rect 1618 3635 1652 3669
rect 1618 3567 1652 3601
rect 1618 3499 1652 3533
rect 1618 3431 1652 3465
rect 1618 3363 1652 3397
rect 1618 3295 1652 3329
rect 1618 3227 1652 3261
rect 1618 3159 1652 3193
rect 1618 3091 1652 3125
rect 1618 3023 1652 3057
rect 1618 2955 1652 2989
rect 1618 2887 1652 2921
rect 1618 2819 1652 2853
rect 1618 2751 1652 2785
rect 1618 2683 1652 2717
rect 1618 2615 1652 2649
rect 1618 2547 1652 2581
rect 1618 2479 1652 2513
rect 1618 2411 1652 2445
rect 1618 2343 1652 2377
rect 88 2309 122 2343
rect 156 2309 190 2343
rect 224 2309 258 2343
rect 292 2309 326 2343
rect 360 2309 394 2343
rect 428 2309 462 2343
rect 496 2309 530 2343
rect 564 2309 598 2343
rect 632 2309 666 2343
rect 700 2309 734 2343
rect 768 2309 802 2343
rect 836 2309 870 2343
rect 904 2309 938 2343
rect 972 2309 1006 2343
rect 1040 2309 1074 2343
rect 1108 2309 1142 2343
rect 1176 2309 1210 2343
rect 1244 2309 1278 2343
rect 1312 2309 1346 2343
rect 1380 2309 1414 2343
rect 1448 2309 1482 2343
rect 1516 2309 1550 2343
rect -45 2269 -11 2303
rect -45 2201 -11 2235
rect -45 2133 -11 2167
rect -45 2065 -11 2099
rect -45 1997 -11 2031
rect -45 1929 -11 1963
rect -45 1861 -11 1895
rect -45 1793 -11 1827
rect -45 1725 -11 1759
rect -45 1657 -11 1691
rect -45 1589 -11 1623
rect 1686 2302 1720 2336
rect 1754 2302 1788 2336
rect 721 2241 755 2275
rect 721 2173 755 2207
rect 1855 2206 1889 2240
rect 721 2105 755 2139
rect 721 2037 755 2071
rect 721 1969 755 2003
rect 721 1901 755 1935
rect 721 1833 755 1867
rect 721 1765 755 1799
rect 721 1697 755 1731
rect 721 1629 755 1663
rect -45 1521 -11 1555
rect 721 1561 755 1595
rect -45 1453 -11 1487
rect 721 1493 755 1527
rect 1855 2135 1889 2169
rect 1855 2064 1889 2098
rect 1855 1993 1889 2027
rect 1855 1922 1889 1956
rect 1855 1851 1889 1885
rect 1855 1780 1889 1814
rect 1855 1709 1889 1743
rect 1855 1638 1889 1672
rect 1855 1567 1889 1601
rect 1855 1496 1889 1530
rect 721 1425 755 1459
rect -45 1385 -11 1419
rect -45 1317 -11 1351
rect -45 1249 -11 1283
rect -45 1181 -11 1215
rect -45 1113 -11 1147
rect -45 1045 -11 1079
rect -45 977 -11 1011
rect -45 909 -11 943
rect -45 841 -11 875
rect -45 773 -11 807
rect -45 705 -11 739
rect 721 1357 755 1391
rect 1855 1425 1889 1459
rect 721 1289 755 1323
rect 1855 1354 1889 1388
rect 721 1221 755 1255
rect 721 1153 755 1187
rect 721 1085 755 1119
rect 721 1017 755 1051
rect 721 949 755 983
rect 721 881 755 915
rect 1855 914 1889 948
rect 721 813 755 847
rect 1855 841 1889 875
rect 721 745 755 779
rect -45 637 -11 671
rect 721 677 755 711
rect -45 569 -11 603
rect -45 501 -11 535
rect -45 433 -11 467
rect -45 365 -11 399
rect -45 297 -11 331
rect -45 229 -11 263
rect -45 161 -11 195
rect -45 93 -11 127
rect -45 25 -11 59
rect -45 -43 -11 -9
rect 721 609 755 643
rect 721 541 755 575
rect 721 473 755 507
rect 721 405 755 439
rect 721 337 755 371
rect 721 269 755 303
rect 721 201 755 235
rect 721 133 755 167
rect 1855 768 1889 802
rect 1855 695 1889 729
rect 1855 622 1889 656
rect 1855 549 1889 583
rect 1855 477 1889 511
rect 1855 405 1889 439
rect 1855 333 1889 367
rect 1855 261 1889 295
rect 1855 189 1889 223
rect 1855 117 1889 151
rect 721 65 755 99
rect 1855 45 1889 79
rect 1855 -27 1889 7
rect 75 -77 109 -43
rect 143 -77 177 -43
rect 211 -77 245 -43
rect 279 -77 313 -43
rect 347 -77 381 -43
rect 415 -77 449 -43
rect 483 -77 517 -43
rect 551 -77 585 -43
rect 619 -77 653 -43
rect 687 -77 721 -43
rect 789 -70 823 -36
rect 857 -70 891 -36
rect 925 -70 959 -36
rect 993 -70 1027 -36
rect 1061 -70 1095 -36
rect 1129 -70 1163 -36
rect 1197 -70 1231 -36
rect 1265 -70 1299 -36
rect 1333 -70 1367 -36
rect 1401 -70 1435 -36
rect 1469 -70 1503 -36
rect 1537 -70 1571 -36
rect 1605 -70 1639 -36
rect 1673 -70 1707 -36
rect 1741 -70 1775 -36
<< mvnsubdiffcont >>
rect -1082 4607 -1048 4641
rect -1014 4607 -980 4641
rect -946 4607 -912 4641
rect -878 4607 -844 4641
rect -810 4607 -776 4641
rect -742 4607 -708 4641
rect -674 4607 -640 4641
rect -606 4607 -572 4641
rect -538 4607 -504 4641
rect -470 4607 -436 4641
rect -402 4607 -368 4641
rect -334 4607 -300 4641
rect -266 4607 -232 4641
rect -1207 4573 -1173 4607
rect -1207 4505 -1173 4539
rect -1207 4437 -1173 4471
rect -232 4498 -198 4532
rect -1207 4369 -1173 4403
rect -1207 4301 -1173 4335
rect -1207 4233 -1173 4267
rect -1207 4165 -1173 4199
rect -1717 4062 -1683 4096
rect -1649 4062 -1615 4096
rect -1581 4062 -1547 4096
rect -1513 4062 -1479 4096
rect -1445 4062 -1411 4096
rect -1377 4062 -1343 4096
rect -1309 4062 -1275 4096
rect -1241 4062 -1207 4096
rect -232 4430 -198 4464
rect -232 4362 -198 4396
rect -232 4294 -198 4328
rect -232 4226 -198 4260
rect -232 4158 -198 4192
rect -232 4090 -198 4124
rect -1802 3994 -1768 4028
rect -232 4022 -198 4056
rect -1802 3926 -1768 3960
rect -1802 3858 -1768 3892
rect -1802 3790 -1768 3824
rect -1802 3722 -1768 3756
rect -1802 3654 -1768 3688
rect -1802 3586 -1768 3620
rect -232 3954 -198 3988
rect -232 3886 -198 3920
rect -232 3818 -198 3852
rect -232 3750 -198 3784
rect -232 3682 -198 3716
rect -1802 3518 -1768 3552
rect -232 3547 -198 3581
rect -1802 3450 -1768 3484
rect -1802 3382 -1768 3416
rect -232 3479 -198 3513
rect -232 3411 -198 3445
rect -1734 3348 -1700 3382
rect -1666 3348 -1632 3382
rect -1598 3348 -1564 3382
rect -1530 3348 -1496 3382
rect -1462 3348 -1428 3382
rect -1394 3348 -1360 3382
rect -1326 3348 -1292 3382
rect -1258 3348 -1224 3382
rect -1190 3348 -1156 3382
rect -1122 3348 -1088 3382
rect -1054 3348 -1020 3382
rect -986 3348 -952 3382
rect -918 3348 -884 3382
rect -850 3348 -816 3382
rect -782 3348 -748 3382
rect -714 3348 -680 3382
rect -580 3309 -546 3343
rect -580 3241 -546 3275
rect -232 3343 -198 3377
rect -232 3275 -198 3309
rect -232 3207 -198 3241
rect -546 3173 -512 3207
rect -478 3173 -444 3207
rect -410 3173 -376 3207
rect -342 3173 -308 3207
rect 953 2115 987 2149
rect 1021 2115 1055 2149
rect 1089 2115 1123 2149
rect 1157 2115 1191 2149
rect 1225 2115 1259 2149
rect 1293 2115 1327 2149
rect 1361 2115 1395 2149
rect 1429 2115 1463 2149
rect 1497 2115 1531 2149
rect 1565 2115 1599 2149
rect 1668 2081 1702 2115
rect 1668 2013 1702 2047
rect 1668 1945 1702 1979
rect 1668 1877 1702 1911
rect 1668 1809 1702 1843
rect 1668 1741 1702 1775
rect 1668 1673 1702 1707
rect 1668 1605 1702 1639
rect 1668 1537 1702 1571
rect 908 737 942 771
rect 908 669 942 703
rect 908 601 942 635
rect 908 533 942 567
rect 908 465 942 499
rect 908 397 942 431
rect 908 329 942 363
rect 908 261 942 295
rect 1668 695 1702 729
rect 1668 627 1702 661
rect 1668 559 1702 593
rect 1668 491 1702 525
rect 1668 423 1702 457
rect 1668 355 1702 389
rect 1668 287 1702 321
rect 1668 219 1702 253
rect 1668 151 1702 185
rect 942 117 976 151
rect 1010 117 1044 151
rect 1078 117 1112 151
rect 1146 117 1180 151
rect 1214 117 1248 151
rect 1282 117 1316 151
rect 1350 117 1384 151
rect 1418 117 1452 151
rect 1486 117 1520 151
rect 1554 117 1588 151
<< poly >>
rect -1063 4557 -963 4573
rect -1063 4523 -1030 4557
rect -996 4523 -963 4557
rect -1063 4489 -963 4523
rect -1063 4455 -1030 4489
rect -996 4455 -963 4489
rect -1063 4433 -963 4455
rect -907 4557 -807 4573
rect -907 4523 -874 4557
rect -840 4523 -807 4557
rect -907 4489 -807 4523
rect -907 4455 -874 4489
rect -840 4455 -807 4489
rect -907 4433 -807 4455
rect -751 4557 -651 4573
rect -751 4523 -718 4557
rect -684 4523 -651 4557
rect -751 4489 -651 4523
rect -751 4455 -718 4489
rect -684 4455 -651 4489
rect -751 4433 -651 4455
rect -595 4557 -495 4573
rect -595 4523 -562 4557
rect -528 4523 -495 4557
rect -595 4489 -495 4523
rect -595 4455 -562 4489
rect -528 4455 -495 4489
rect -595 4433 -495 4455
rect -439 4557 -339 4573
rect -439 4523 -406 4557
rect -372 4523 -339 4557
rect -439 4489 -339 4523
rect -439 4455 -406 4489
rect -372 4455 -339 4489
rect -439 4433 -339 4455
rect -439 4039 -339 4081
rect -864 4023 -495 4039
rect -864 3989 -848 4023
rect -814 3989 -773 4023
rect -739 3989 -697 4023
rect -663 3989 -621 4023
rect -587 3989 -545 4023
rect -511 3989 -495 4023
rect -864 3973 -495 3989
rect -864 3967 -764 3973
rect -595 3967 -495 3973
rect -439 4023 -305 4039
rect -439 3989 -423 4023
rect -389 3989 -355 4023
rect -321 3989 -305 4023
rect -439 3973 -305 3989
rect -439 3967 -339 3973
rect -1632 3573 -1232 3615
rect -1176 3573 -1076 3615
rect -1632 3557 -1076 3573
rect -1632 3523 -1616 3557
rect -1582 3523 -1546 3557
rect -1512 3523 -1476 3557
rect -1442 3523 -1406 3557
rect -1372 3523 -1336 3557
rect -1302 3523 -1266 3557
rect -1232 3523 -1196 3557
rect -1162 3523 -1126 3557
rect -1092 3523 -1076 3557
rect -1632 3507 -1076 3523
rect -1020 3573 -920 3615
rect -439 3607 -339 3615
rect -1020 3557 -886 3573
rect -1020 3523 -1004 3557
rect -970 3523 -936 3557
rect -902 3523 -886 3557
rect -1020 3507 -886 3523
rect 147 4557 327 4573
rect 147 4523 163 4557
rect 197 4523 254 4557
rect 288 4523 327 4557
rect 147 4501 327 4523
rect 383 4557 563 4573
rect 383 4523 399 4557
rect 433 4523 513 4557
rect 547 4523 563 4557
rect 383 4501 563 4523
rect 619 4557 799 4573
rect 619 4523 635 4557
rect 669 4523 749 4557
rect 783 4523 799 4557
rect 619 4501 799 4523
rect 1311 4557 1491 4573
rect 1311 4523 1327 4557
rect 1361 4523 1441 4557
rect 1475 4523 1491 4557
rect 1311 4501 1491 4523
rect 147 2427 327 2449
rect 147 2393 163 2427
rect 197 2393 254 2427
rect 288 2393 327 2427
rect 147 2377 327 2393
rect 383 2427 563 2449
rect 383 2393 399 2427
rect 433 2393 513 2427
rect 547 2393 563 2427
rect 383 2377 563 2393
rect 619 2427 799 2449
rect 619 2393 635 2427
rect 669 2393 749 2427
rect 783 2393 799 2427
rect 619 2377 799 2393
rect 1311 2427 1491 2449
rect 1311 2393 1327 2427
rect 1361 2393 1441 2427
rect 1475 2393 1491 2427
rect 1311 2377 1491 2393
rect 119 1603 239 1609
rect 105 1587 239 1603
rect 105 1553 121 1587
rect 155 1553 189 1587
rect 223 1553 239 1587
rect 105 1537 239 1553
rect 295 1603 415 1609
rect 471 1603 591 1609
rect 295 1587 591 1603
rect 295 1553 311 1587
rect 345 1553 387 1587
rect 421 1553 464 1587
rect 498 1553 541 1587
rect 575 1553 591 1587
rect 295 1537 591 1553
rect 135 1479 335 1495
rect 135 1445 151 1479
rect 185 1445 285 1479
rect 319 1445 335 1479
rect 135 1423 335 1445
rect 391 1479 591 1495
rect 391 1445 407 1479
rect 441 1445 541 1479
rect 575 1445 591 1479
rect 391 1423 591 1445
rect 1049 1429 1149 1435
rect 1205 1429 1305 1435
rect 1049 1413 1305 1429
rect 1049 1379 1092 1413
rect 1126 1379 1160 1413
rect 1194 1379 1228 1413
rect 1262 1379 1305 1413
rect 1049 1363 1305 1379
rect 1361 1413 1561 1435
rect 1361 1379 1410 1413
rect 1444 1379 1478 1413
rect 1512 1379 1561 1413
rect 1361 1363 1561 1379
rect 1049 887 1305 903
rect 1049 853 1092 887
rect 1126 853 1160 887
rect 1194 853 1228 887
rect 1262 853 1305 887
rect 1049 837 1305 853
rect 1049 831 1149 837
rect 1205 831 1305 837
rect 1361 887 1561 903
rect 1361 853 1410 887
rect 1444 853 1478 887
rect 1512 853 1561 887
rect 1361 831 1561 853
rect 105 713 239 729
rect 105 679 121 713
rect 155 679 189 713
rect 223 679 239 713
rect 105 663 239 679
rect 119 657 239 663
rect 295 713 591 729
rect 295 679 311 713
rect 345 679 387 713
rect 421 679 464 713
rect 498 679 541 713
rect 575 679 591 713
rect 295 663 591 679
rect 295 657 415 663
rect 471 657 591 663
<< polycont >>
rect -1030 4523 -996 4557
rect -1030 4455 -996 4489
rect -874 4523 -840 4557
rect -874 4455 -840 4489
rect -718 4523 -684 4557
rect -718 4455 -684 4489
rect -562 4523 -528 4557
rect -562 4455 -528 4489
rect -406 4523 -372 4557
rect -406 4455 -372 4489
rect -848 3989 -814 4023
rect -773 3989 -739 4023
rect -697 3989 -663 4023
rect -621 3989 -587 4023
rect -545 3989 -511 4023
rect -423 3989 -389 4023
rect -355 3989 -321 4023
rect -1616 3523 -1582 3557
rect -1546 3523 -1512 3557
rect -1476 3523 -1442 3557
rect -1406 3523 -1372 3557
rect -1336 3523 -1302 3557
rect -1266 3523 -1232 3557
rect -1196 3523 -1162 3557
rect -1126 3523 -1092 3557
rect -1004 3523 -970 3557
rect -936 3523 -902 3557
rect 163 4523 197 4557
rect 254 4523 288 4557
rect 399 4523 433 4557
rect 513 4523 547 4557
rect 635 4523 669 4557
rect 749 4523 783 4557
rect 1327 4523 1361 4557
rect 1441 4523 1475 4557
rect 163 2393 197 2427
rect 254 2393 288 2427
rect 399 2393 433 2427
rect 513 2393 547 2427
rect 635 2393 669 2427
rect 749 2393 783 2427
rect 1327 2393 1361 2427
rect 1441 2393 1475 2427
rect 121 1553 155 1587
rect 189 1553 223 1587
rect 311 1553 345 1587
rect 387 1553 421 1587
rect 464 1553 498 1587
rect 541 1553 575 1587
rect 151 1445 185 1479
rect 285 1445 319 1479
rect 407 1445 441 1479
rect 541 1445 575 1479
rect 1092 1379 1126 1413
rect 1160 1379 1194 1413
rect 1228 1379 1262 1413
rect 1410 1379 1444 1413
rect 1478 1379 1512 1413
rect 1092 853 1126 887
rect 1160 853 1194 887
rect 1228 853 1262 887
rect 1410 853 1444 887
rect 1478 853 1512 887
rect 121 679 155 713
rect 189 679 223 713
rect 311 679 345 713
rect 387 679 421 713
rect 464 679 498 713
rect 541 679 575 713
<< locali >>
rect -1802 4623 -1796 4657
rect -1762 4623 -1721 4657
rect -1687 4623 -1646 4657
rect -1612 4623 -1571 4657
rect -1537 4623 -1496 4657
rect -1462 4623 -1422 4657
rect -1388 4623 -1348 4657
rect -1314 4623 -1274 4657
rect -1240 4623 -1200 4657
rect -1166 4623 -1126 4657
rect -1092 4641 -1052 4657
rect -1018 4641 -978 4657
rect -944 4641 -904 4657
rect -870 4641 -830 4657
rect -796 4641 -756 4657
rect -722 4641 -682 4657
rect -648 4641 -608 4657
rect -574 4641 -534 4657
rect -500 4641 -460 4657
rect -426 4641 -386 4657
rect -352 4641 -312 4657
rect -278 4641 -238 4657
rect -1092 4623 -1082 4641
rect -1018 4623 -1014 4641
rect -1802 4585 -1768 4623
rect -1802 4510 -1768 4551
rect -1207 4607 -1082 4623
rect -1048 4607 -1014 4623
rect -980 4623 -978 4641
rect -912 4623 -904 4641
rect -844 4623 -830 4641
rect -776 4623 -756 4641
rect -708 4623 -682 4641
rect -640 4623 -608 4641
rect -980 4607 -946 4623
rect -912 4607 -878 4623
rect -844 4607 -810 4623
rect -776 4607 -742 4623
rect -708 4607 -674 4623
rect -640 4607 -606 4623
rect -572 4607 -538 4641
rect -500 4623 -470 4641
rect -426 4623 -402 4641
rect -352 4623 -334 4641
rect -278 4623 -266 4641
rect -204 4623 -198 4641
rect -504 4607 -470 4623
rect -436 4607 -402 4623
rect -368 4607 -334 4623
rect -300 4607 -266 4623
rect -1207 4539 -1173 4573
rect -1207 4495 -1173 4505
rect -1802 4435 -1768 4476
rect -1802 4360 -1768 4401
rect -1802 4285 -1768 4326
rect -1802 4210 -1768 4251
rect -1204 4471 -1173 4495
rect -1046 4523 -1030 4557
rect -996 4523 -980 4557
rect -1046 4489 -980 4523
rect -1046 4468 -1030 4489
rect -1238 4437 -1207 4461
rect -1238 4403 -1173 4437
rect -1068 4434 -1030 4468
rect -996 4434 -980 4489
rect -1046 4427 -980 4434
rect -890 4512 -874 4557
rect -840 4512 -824 4557
rect -890 4489 -824 4512
rect -890 4440 -874 4489
rect -840 4440 -824 4489
rect -734 4523 -718 4557
rect -684 4523 -668 4557
rect -734 4489 -668 4523
rect -734 4468 -718 4489
rect -890 4427 -824 4440
rect -756 4434 -718 4468
rect -684 4434 -668 4489
rect -734 4427 -668 4434
rect -578 4512 -562 4557
rect -528 4512 -512 4557
rect -578 4489 -512 4512
rect -578 4440 -562 4489
rect -528 4440 -512 4489
rect -422 4523 -406 4557
rect -372 4523 -356 4557
rect -422 4489 -356 4523
rect -422 4455 -406 4489
rect -372 4455 -356 4489
rect -232 4535 -198 4623
rect -232 4464 -198 4498
rect -578 4427 -512 4440
rect -1238 4389 -1207 4403
rect -1204 4355 -1173 4369
rect -1238 4335 -1173 4355
rect -1238 4301 -1207 4335
rect -1238 4283 -1173 4301
rect -1204 4267 -1173 4283
rect -1802 4135 -1768 4176
rect -1207 4199 -1173 4233
rect -1207 4152 -1173 4165
rect -1802 4096 -1768 4101
rect -1336 4118 -1288 4152
rect -1254 4118 -1207 4152
rect -1108 4260 -1074 4319
rect -1108 4167 -1074 4226
rect -948 4321 -914 4359
rect -948 4249 -914 4287
rect -796 4260 -762 4319
rect -796 4167 -762 4226
rect -636 4250 -602 4359
rect -484 4260 -450 4319
rect -484 4167 -450 4226
rect -416 4174 -363 4455
rect -232 4396 -198 4430
rect -416 4140 -410 4174
rect -376 4140 -363 4174
rect -1370 4096 -1173 4118
rect -1802 4062 -1730 4096
rect -1683 4062 -1649 4096
rect -1612 4062 -1581 4096
rect -1547 4062 -1513 4096
rect -1479 4062 -1445 4096
rect -1411 4062 -1377 4096
rect -1343 4062 -1309 4096
rect -1275 4062 -1241 4096
rect -1207 4062 -1173 4096
rect -416 4102 -363 4140
rect -328 4260 -294 4319
rect -328 4167 -294 4226
rect -232 4328 -198 4341
rect -232 4260 -198 4268
rect -232 4192 -198 4195
rect -232 4156 -198 4158
rect -416 4068 -410 4102
rect -376 4068 -363 4102
rect -1802 4060 -1768 4062
rect -416 4023 -363 4068
rect -232 4083 -198 4090
rect -1802 3985 -1768 3994
rect -864 4022 -848 4023
rect -814 4022 -773 4023
rect -739 4022 -697 4023
rect -864 3989 -852 4022
rect -814 3989 -775 4022
rect -739 3989 -698 4022
rect -663 3989 -621 4023
rect -818 3988 -775 3989
rect -741 3988 -698 3989
rect -664 3988 -621 3989
rect -587 3988 -545 4023
rect -511 3989 -495 4023
rect -439 3989 -423 4023
rect -389 3989 -355 4023
rect -321 3989 -305 4023
rect -232 4010 -198 4022
rect -232 3937 -198 3954
rect -1802 3910 -1768 3926
rect -1802 3835 -1768 3858
rect -1802 3760 -1768 3790
rect -1802 3688 -1768 3722
rect -1677 3864 -1643 3902
rect -1677 3792 -1643 3830
rect -1677 3719 -1643 3758
rect -1221 3855 -1187 3902
rect -232 3864 -198 3886
rect -1221 3774 -1187 3821
rect -1221 3693 -1187 3740
rect -1065 3765 -1031 3803
rect -1065 3693 -1031 3731
rect -987 3672 -953 3710
rect -1802 3620 -1768 3651
rect -1802 3552 -1768 3576
rect -987 3557 -953 3638
rect -909 3714 -875 3752
rect -909 3642 -875 3680
rect -753 3765 -719 3803
rect -753 3693 -719 3731
rect -640 3765 -606 3803
rect -640 3693 -606 3731
rect -484 3765 -450 3803
rect -484 3693 -450 3731
rect -328 3765 -294 3803
rect -328 3693 -294 3731
rect -232 3791 -198 3818
rect -232 3718 -198 3750
rect -232 3645 -198 3682
rect -232 3581 -198 3611
rect -1632 3523 -1625 3557
rect -1582 3523 -1546 3557
rect -1508 3523 -1476 3557
rect -1424 3523 -1406 3557
rect -1340 3523 -1336 3557
rect -1302 3523 -1290 3557
rect -1232 3523 -1206 3557
rect -1162 3523 -1126 3557
rect -1088 3523 -1076 3557
rect -1020 3523 -1004 3557
rect -970 3523 -936 3557
rect -902 3523 -886 3557
rect -1802 3484 -1768 3502
rect -1802 3416 -1768 3428
rect -232 3513 -198 3539
rect -232 3445 -198 3467
rect -1768 3354 -1734 3382
rect -1802 3348 -1734 3354
rect -1696 3348 -1666 3382
rect -1619 3348 -1598 3382
rect -1542 3348 -1530 3382
rect -1465 3348 -1462 3382
rect -1428 3348 -1422 3382
rect -1360 3348 -1345 3382
rect -1292 3348 -1268 3382
rect -1224 3348 -1191 3382
rect -1156 3348 -1122 3382
rect -1080 3348 -1054 3382
rect -1003 3348 -986 3382
rect -926 3348 -918 3382
rect -884 3348 -883 3382
rect -816 3348 -806 3382
rect -748 3348 -729 3382
rect -680 3348 -652 3382
rect -618 3376 -546 3382
rect -618 3348 -580 3376
rect -580 3279 -546 3309
rect -580 3207 -546 3241
rect -232 3377 -198 3395
rect -232 3309 -198 3323
rect -232 3241 -198 3251
rect -580 3173 -574 3207
rect -512 3173 -484 3207
rect -444 3173 -410 3207
rect -360 3173 -342 3207
rect -308 3173 -304 3207
rect -270 3179 -232 3207
rect -270 3173 -198 3179
rect -45 4607 -14 4641
rect 20 4607 60 4641
rect 122 4607 134 4641
rect 190 4607 208 4641
rect 258 4607 282 4641
rect 326 4607 356 4641
rect 394 4607 428 4641
rect 464 4607 496 4641
rect 538 4607 564 4641
rect 612 4607 632 4641
rect 686 4607 700 4641
rect 760 4607 768 4641
rect 834 4607 836 4641
rect 870 4607 874 4641
rect 938 4607 948 4641
rect 1006 4607 1022 4641
rect 1074 4607 1096 4641
rect 1142 4607 1171 4641
rect 1210 4607 1244 4641
rect 1280 4607 1312 4641
rect 1355 4607 1380 4641
rect 1430 4607 1448 4641
rect 1505 4607 1516 4641
rect 1580 4607 1584 4641
rect 1618 4635 1652 4641
rect -11 4573 14 4607
rect -45 4539 14 4573
rect -11 4535 14 4539
rect 147 4523 163 4557
rect 216 4523 254 4557
rect 292 4523 304 4557
rect 338 4523 399 4557
rect 433 4523 513 4557
rect 547 4523 563 4557
rect 619 4523 635 4557
rect 669 4523 749 4557
rect 783 4523 844 4557
rect 954 4546 1156 4607
rect 1618 4562 1652 4601
rect -45 4501 -20 4505
rect -45 4471 -11 4501
rect 338 4449 372 4523
rect 810 4449 844 4523
rect 1266 4523 1327 4557
rect 1361 4523 1441 4557
rect 1475 4523 1491 4557
rect 1266 4449 1300 4523
rect 1618 4489 1652 4519
rect -45 4403 -11 4437
rect 1618 4417 1652 4451
rect -45 4341 -20 4369
rect -45 4335 14 4341
rect -11 4303 14 4335
rect -45 4269 -20 4301
rect -45 4267 14 4269
rect -11 4233 14 4267
rect -45 4231 14 4233
rect -45 4199 -20 4231
rect -11 4165 14 4197
rect -45 4159 14 4165
rect -45 4131 -20 4159
rect -11 4097 14 4125
rect -45 4087 14 4097
rect -45 4063 -20 4087
rect -11 4029 14 4053
rect -45 4015 14 4029
rect -45 3995 -20 4015
rect -11 3961 14 3981
rect -45 3943 14 3961
rect -45 3927 -20 3943
rect -11 3893 14 3909
rect -45 3871 14 3893
rect -45 3859 -20 3871
rect -11 3825 14 3837
rect -45 3799 14 3825
rect -45 3791 -20 3799
rect -11 3757 14 3765
rect -45 3727 14 3757
rect -45 3723 -20 3727
rect -11 3689 14 3693
rect -45 3655 14 3689
rect -45 3587 14 3621
rect -11 3583 14 3587
rect -45 3549 -20 3553
rect -45 3519 14 3549
rect -11 3511 14 3519
rect -45 3477 -20 3485
rect -45 3451 14 3477
rect -11 3439 14 3451
rect -45 3405 -20 3417
rect -45 3383 14 3405
rect -11 3367 14 3383
rect -45 3333 -20 3349
rect -45 3315 14 3333
rect -11 3295 14 3315
rect -45 3261 -20 3281
rect -45 3247 14 3261
rect -11 3223 14 3247
rect -45 3189 -20 3213
rect -45 3179 14 3189
rect -11 3151 14 3179
rect -45 3117 -20 3145
rect -45 3111 14 3117
rect -11 3079 14 3111
rect -45 3045 -20 3077
rect -45 3043 14 3045
rect -11 3009 14 3043
rect -45 3007 14 3009
rect -45 2975 -20 3007
rect -11 2941 14 2973
rect -45 2935 14 2941
rect -45 2907 -20 2935
rect -11 2873 14 2901
rect -45 2863 14 2873
rect -45 2839 -20 2863
rect -11 2805 14 2829
rect -45 2791 14 2805
rect -45 2771 -20 2791
rect -11 2737 14 2757
rect -45 2719 14 2737
rect -45 2703 -20 2719
rect -11 2669 14 2685
rect -45 2647 14 2669
rect -45 2635 -20 2647
rect -11 2601 14 2613
rect -45 2575 14 2601
rect -45 2567 -20 2575
rect -11 2533 14 2541
rect -45 2503 14 2533
rect -45 2469 -20 2503
rect 1618 4349 1652 4382
rect 1618 4281 1652 4309
rect 1618 4213 1652 4236
rect 1618 4145 1652 4163
rect 1618 4077 1652 4090
rect 1618 4009 1652 4017
rect 1618 3941 1652 3943
rect 1618 3903 1652 3907
rect 1618 3829 1652 3839
rect 1618 3755 1652 3771
rect 1618 3681 1652 3703
rect 1618 3607 1652 3635
rect 1618 3533 1652 3567
rect 1618 3465 1652 3499
rect 1618 3397 1652 3425
rect 1618 3329 1652 3351
rect 1618 3261 1652 3277
rect 1618 3193 1652 3203
rect 1618 3125 1652 3129
rect 1618 3089 1652 3091
rect 1618 3015 1652 3023
rect 1618 2941 1652 2955
rect 1618 2867 1652 2887
rect 1618 2793 1652 2819
rect 1618 2719 1652 2751
rect 1618 2649 1652 2683
rect 1618 2581 1652 2611
rect 1618 2513 1652 2537
rect -45 2431 14 2469
rect -45 2397 -20 2431
rect 216 2453 258 2487
rect 182 2427 292 2453
rect 338 2427 372 2471
rect 810 2427 844 2471
rect -45 2359 14 2397
rect 147 2393 163 2427
rect 197 2393 254 2427
rect 288 2393 304 2427
rect 338 2393 399 2427
rect 433 2393 513 2427
rect 547 2393 563 2427
rect 619 2393 635 2427
rect 669 2393 749 2427
rect 783 2393 844 2427
rect 1266 2427 1300 2501
rect 1618 2445 1652 2463
rect -45 2325 -20 2359
rect 954 2343 1156 2404
rect 1266 2393 1327 2427
rect 1361 2393 1441 2427
rect 1475 2393 1491 2427
rect 1618 2377 1652 2389
rect 14 2325 88 2343
rect -45 2309 88 2325
rect 122 2309 156 2343
rect 190 2309 198 2343
rect 258 2309 272 2343
rect 326 2309 346 2343
rect 394 2309 420 2343
rect 462 2309 494 2343
rect 530 2309 564 2343
rect 602 2309 632 2343
rect 676 2309 700 2343
rect 750 2309 768 2343
rect 824 2309 836 2343
rect 898 2309 904 2343
rect 1006 2309 1012 2343
rect 1074 2309 1087 2343
rect 1142 2309 1176 2343
rect 1210 2309 1244 2343
rect 1278 2309 1312 2343
rect 1346 2309 1380 2343
rect 1414 2309 1448 2343
rect 1482 2309 1516 2343
rect 1550 2315 1618 2343
rect 1743 2336 1889 2343
rect 1652 2315 1686 2336
rect 1550 2309 1686 2315
rect 1743 2309 1754 2336
rect -45 2303 14 2309
rect -11 2287 14 2303
rect -45 2253 -20 2269
rect -45 2235 14 2253
rect 250 2239 284 2309
rect 602 2302 1686 2309
rect 1720 2302 1754 2309
rect 1788 2305 1889 2336
rect 1788 2302 1855 2305
rect 602 2275 755 2302
rect -11 2214 14 2235
rect -45 2180 -20 2201
rect -45 2167 14 2180
rect -11 2141 14 2167
rect -45 2107 -20 2133
rect -45 2099 14 2107
rect -11 2068 14 2099
rect -45 2034 -20 2065
rect -45 2031 14 2034
rect -11 1997 14 2031
rect -45 1995 14 1997
rect -45 1963 -20 1995
rect -11 1929 14 1961
rect -45 1922 14 1929
rect -45 1895 -20 1922
rect -11 1861 14 1888
rect -45 1849 14 1861
rect -45 1827 -20 1849
rect 74 2089 108 2141
rect 74 2003 108 2055
rect 74 1917 108 1969
rect 74 1830 108 1883
rect 251 2138 285 2180
rect 251 2061 285 2104
rect 251 1984 285 2027
rect 251 1907 285 1950
rect 251 1830 285 1873
rect 426 2035 479 2239
rect 426 2001 445 2035
rect 426 1951 479 2001
rect 426 1917 445 1951
rect 426 1867 479 1917
rect 426 1833 445 1867
rect -45 1759 -11 1793
rect -45 1691 -11 1725
rect 426 1783 479 1833
rect 426 1749 445 1783
rect 426 1699 479 1749
rect 426 1665 445 1699
rect 602 2237 721 2275
rect 602 2214 755 2237
rect 636 2207 755 2214
rect 636 2180 721 2207
rect 602 2153 721 2180
rect 602 2141 755 2153
rect 1855 2240 1889 2271
rect 1855 2169 1889 2197
rect 636 2139 755 2141
rect 636 2107 721 2139
rect 602 2105 721 2107
rect 919 2115 953 2149
rect 1014 2115 1021 2149
rect 1055 2115 1057 2149
rect 1123 2115 1134 2149
rect 1191 2115 1211 2149
rect 1259 2115 1288 2149
rect 1327 2115 1361 2149
rect 1399 2115 1429 2149
rect 1476 2115 1497 2149
rect 1553 2115 1565 2149
rect 1630 2143 1702 2149
rect 1630 2115 1668 2143
rect 602 2103 755 2105
rect 602 2067 721 2103
rect 636 2037 721 2067
rect 1668 2062 1702 2081
rect 636 2033 755 2037
rect 602 2020 755 2033
rect 602 1993 721 2020
rect 636 1969 721 1993
rect 636 1959 755 1969
rect 602 1937 755 1959
rect 602 1919 721 1937
rect 636 1901 721 1919
rect 636 1885 755 1901
rect 602 1867 755 1885
rect 602 1845 721 1867
rect 636 1820 721 1845
rect 636 1811 755 1820
rect 602 1799 755 1811
rect 602 1771 721 1799
rect 636 1737 721 1771
rect 602 1731 755 1737
rect 602 1697 721 1731
rect -45 1623 -11 1657
rect -45 1555 -11 1589
rect 721 1663 755 1697
rect 721 1613 755 1629
rect 105 1553 120 1587
rect 155 1553 189 1587
rect 236 1553 239 1587
rect 295 1553 311 1587
rect 345 1553 387 1587
rect 426 1553 464 1587
rect 504 1553 541 1587
rect 582 1553 591 1587
rect -45 1487 -11 1521
rect 721 1535 755 1561
rect 1004 1926 1038 1965
rect 1004 1853 1038 1892
rect 1004 1780 1038 1819
rect 1004 1707 1038 1746
rect 1004 1634 1038 1673
rect 1004 1561 1038 1600
rect 1160 1976 1194 2019
rect 1160 1900 1194 1942
rect 1160 1824 1194 1866
rect 1160 1748 1194 1790
rect 1160 1672 1194 1714
rect 1160 1596 1194 1638
rect 1316 1955 1350 2000
rect 1316 1876 1350 1921
rect 1316 1797 1350 1842
rect 1316 1718 1350 1763
rect 1316 1639 1350 1684
rect 1572 1979 1606 2019
rect 1572 1905 1606 1945
rect 1572 1831 1606 1871
rect 1572 1758 1606 1797
rect 1572 1685 1606 1724
rect 1668 1981 1702 2013
rect 1668 1911 1702 1945
rect 1668 1843 1702 1866
rect 1668 1775 1702 1786
rect 1668 1740 1702 1741
rect 1668 1660 1702 1673
rect 1316 1561 1350 1605
rect 1668 1580 1702 1605
rect -45 1419 -11 1453
rect 135 1445 151 1479
rect 191 1445 285 1479
rect 323 1445 335 1479
rect 391 1445 403 1479
rect 441 1445 487 1479
rect 521 1445 541 1479
rect 575 1445 591 1479
rect 721 1459 755 1493
rect 1668 1461 1702 1537
rect 1855 2098 1889 2123
rect 1855 2027 1889 2049
rect 1855 1956 1889 1975
rect 1855 1885 1889 1901
rect 1855 1814 1889 1827
rect 1855 1743 1889 1753
rect 1855 1672 1889 1679
rect 1855 1601 1889 1605
rect 1855 1565 1889 1567
rect 1855 1530 1889 1531
rect 1855 1491 1889 1496
rect -45 1359 -20 1385
rect -45 1351 14 1359
rect -11 1321 14 1351
rect 721 1391 755 1423
rect 1855 1417 1889 1425
rect 1076 1409 1092 1413
rect 1076 1375 1088 1409
rect 1126 1379 1160 1413
rect 1194 1409 1228 1413
rect 1262 1409 1278 1413
rect 1394 1409 1410 1413
rect 1444 1409 1478 1413
rect 1512 1409 1528 1413
rect 1204 1379 1228 1409
rect 1122 1375 1170 1379
rect 1204 1375 1252 1379
rect 1286 1375 1334 1409
rect 1368 1379 1410 1409
rect 1450 1379 1478 1409
rect 1368 1375 1416 1379
rect 1450 1375 1498 1379
rect 1532 1375 1579 1409
rect 721 1343 755 1346
rect -45 1287 -20 1317
rect -45 1283 14 1287
rect -11 1249 14 1283
rect -45 1215 -20 1249
rect -11 1181 14 1215
rect -45 1177 14 1181
rect -45 1147 -20 1177
rect -11 1113 14 1143
rect -45 1105 14 1113
rect -45 1079 -20 1105
rect -11 1045 14 1071
rect -45 1033 14 1045
rect -45 1011 -20 1033
rect -11 977 14 999
rect -45 961 14 977
rect -45 943 -20 961
rect -11 909 14 927
rect -45 889 14 909
rect -45 875 -20 889
rect -11 841 14 855
rect -45 817 14 841
rect -45 807 -20 817
rect 90 1270 124 1309
rect 90 1197 124 1236
rect 636 1323 755 1343
rect 636 1309 721 1323
rect 602 1271 721 1309
rect 636 1269 721 1271
rect 636 1268 755 1269
rect 1855 1343 1889 1354
rect 1855 1270 1889 1309
rect 636 1255 789 1268
rect 636 1237 721 1255
rect 602 1199 721 1237
rect 636 1192 721 1199
rect 755 1192 789 1255
rect 636 1187 789 1192
rect 636 1165 721 1187
rect 90 1123 124 1163
rect 90 1049 124 1089
rect 90 975 124 1015
rect 90 901 124 941
rect 90 827 124 867
rect 346 1086 380 1131
rect 346 1006 380 1052
rect 346 926 380 972
rect 346 846 380 892
rect 602 1153 721 1165
rect 755 1153 789 1187
rect 602 1149 789 1153
rect 602 1127 721 1149
rect 636 1093 721 1127
rect 602 1085 721 1093
rect 755 1085 789 1149
rect 602 1072 789 1085
rect 602 1055 721 1072
rect 636 1021 721 1055
rect 602 1017 721 1021
rect 755 1017 789 1072
rect 602 998 789 1017
rect 1843 1236 1855 1268
rect 1843 1197 1889 1236
rect 1843 1163 1855 1197
rect 1843 1124 1889 1163
rect 1843 1090 1855 1124
rect 1843 1051 1889 1090
rect 1843 1017 1855 1051
rect 1843 998 1889 1017
rect 602 995 755 998
rect 602 983 721 995
rect 636 949 721 983
rect 602 918 755 949
rect 602 911 721 918
rect 636 881 721 911
rect 1855 978 1889 998
rect 1855 905 1889 914
rect 636 877 755 881
rect 602 847 755 877
rect 1076 857 1088 891
rect 1122 887 1170 891
rect 1204 887 1252 891
rect 1076 853 1092 857
rect 1126 853 1160 887
rect 1204 857 1228 887
rect 1286 857 1334 891
rect 1368 887 1416 891
rect 1450 887 1498 891
rect 1368 857 1410 887
rect 1450 857 1478 887
rect 1532 857 1579 891
rect 1194 853 1228 857
rect 1262 853 1278 857
rect 1394 853 1410 857
rect 1444 853 1478 857
rect 1512 853 1528 857
rect 602 839 721 847
rect 636 807 721 839
rect 636 805 755 807
rect 1855 832 1889 841
rect 602 793 755 805
rect -11 773 14 783
rect -45 745 14 773
rect -45 739 -20 745
rect 721 779 755 793
rect -11 705 14 711
rect -45 673 14 705
rect 105 679 117 713
rect 155 679 189 713
rect 236 679 239 713
rect 295 679 311 713
rect 345 679 387 713
rect 423 679 464 713
rect 501 679 541 713
rect 579 679 591 713
rect 721 711 755 730
rect -45 671 -20 673
rect -11 637 14 639
rect -45 603 14 637
rect -11 601 14 603
rect 721 643 755 653
rect -45 567 -20 569
rect -45 535 14 567
rect -11 529 14 535
rect -45 495 -20 501
rect -45 467 14 495
rect -11 457 14 467
rect -45 423 -20 433
rect -45 399 14 423
rect -11 384 14 399
rect -45 350 -20 365
rect -45 331 14 350
rect -11 311 14 331
rect -45 277 -20 297
rect -45 263 14 277
rect -11 238 14 263
rect -45 204 -20 229
rect -45 195 14 204
rect -11 165 14 195
rect -45 131 -20 161
rect -45 127 14 131
rect -11 93 14 127
rect -45 92 14 93
rect -45 59 -20 92
rect 74 487 108 534
rect 426 567 439 601
rect 721 575 755 609
rect 426 528 473 567
rect 74 406 108 453
rect 74 326 108 372
rect 74 246 108 292
rect 74 166 108 212
rect 250 411 284 467
rect 250 321 284 377
rect 250 231 284 287
rect 426 494 439 528
rect 426 456 473 494
rect 426 422 439 456
rect 426 384 473 422
rect 426 350 439 384
rect 74 86 108 132
rect 426 27 473 350
rect 602 541 721 569
rect 602 529 755 541
rect 636 495 721 529
rect 602 473 721 495
rect 602 453 755 473
rect 636 446 755 453
rect 636 419 721 446
rect 602 405 721 419
rect 602 377 755 405
rect 636 371 755 377
rect 636 343 721 371
rect 602 329 721 343
rect 602 303 755 329
rect 602 302 721 303
rect 636 268 721 302
rect 602 246 721 268
rect 602 235 755 246
rect 602 227 721 235
rect 636 201 721 227
rect 636 197 755 201
rect 636 193 721 197
rect 602 152 721 193
rect 636 133 721 152
rect 636 118 755 133
rect 602 114 755 118
rect 908 771 942 805
rect 908 703 942 705
rect 908 667 942 669
rect 908 595 942 601
rect 908 522 942 533
rect 908 449 942 465
rect 908 376 942 397
rect 908 303 942 329
rect 1004 666 1038 705
rect 1004 593 1038 632
rect 1004 520 1038 559
rect 1004 446 1038 486
rect 1004 372 1038 412
rect 1004 298 1038 338
rect 1160 628 1194 670
rect 1160 552 1194 594
rect 1160 476 1194 518
rect 1160 400 1194 442
rect 1160 324 1194 366
rect 908 230 942 261
rect 1160 247 1194 290
rect 1316 661 1350 705
rect 1316 582 1350 627
rect 1668 729 1702 805
rect 1668 661 1702 686
rect 1316 503 1350 548
rect 1316 424 1350 469
rect 1316 345 1350 390
rect 1316 266 1350 311
rect 1572 542 1606 581
rect 1572 469 1606 508
rect 1572 395 1606 435
rect 1572 321 1606 361
rect 1572 247 1606 287
rect 1668 593 1702 606
rect 1668 525 1702 526
rect 1668 480 1702 491
rect 1668 400 1702 423
rect 1668 321 1702 355
rect 1668 253 1702 285
rect 908 157 942 196
rect 1668 185 1702 204
rect 908 117 942 123
rect 976 117 980 151
rect 1044 117 1057 151
rect 1112 117 1134 151
rect 1180 117 1211 151
rect 1248 117 1282 151
rect 1322 117 1350 151
rect 1399 117 1418 151
rect 1476 117 1486 151
rect 1553 117 1554 151
rect 1588 117 1596 151
rect 1630 123 1668 151
rect 1630 117 1702 123
rect 1855 759 1889 768
rect 1855 686 1889 695
rect 1855 613 1889 622
rect 1855 540 1889 549
rect 1855 467 1889 477
rect 1855 394 1889 405
rect 1855 321 1889 333
rect 1855 248 1889 261
rect 1855 175 1889 189
rect 602 65 721 114
rect 602 31 755 65
rect -45 -9 -11 25
rect 602 -3 721 31
rect 602 -36 755 -3
rect 1855 102 1889 117
rect 1855 29 1889 45
rect 1855 -36 1889 -27
rect 602 -43 789 -36
rect -45 -77 75 -43
rect 109 -77 143 -43
rect 177 -77 211 -43
rect 245 -77 279 -43
rect 313 -77 347 -43
rect 381 -77 415 -43
rect 449 -77 483 -43
rect 517 -77 551 -43
rect 585 -77 619 -43
rect 653 -77 687 -43
rect 721 -70 789 -43
rect 823 -70 857 -36
rect 891 -70 925 -36
rect 959 -70 993 -36
rect 1027 -70 1061 -36
rect 1095 -70 1129 -36
rect 1163 -70 1197 -36
rect 1231 -70 1265 -36
rect 1299 -70 1333 -36
rect 1367 -70 1401 -36
rect 1435 -70 1469 -36
rect 1503 -70 1537 -36
rect 1571 -70 1605 -36
rect 1639 -70 1673 -36
rect 1707 -70 1741 -36
rect 1775 -70 1889 -36
rect 721 -77 1889 -70
<< viali >>
rect -1796 4623 -1762 4657
rect -1721 4623 -1687 4657
rect -1646 4623 -1612 4657
rect -1571 4623 -1537 4657
rect -1496 4623 -1462 4657
rect -1422 4623 -1388 4657
rect -1348 4623 -1314 4657
rect -1274 4623 -1240 4657
rect -1200 4623 -1166 4657
rect -1126 4623 -1092 4657
rect -1052 4641 -1018 4657
rect -978 4641 -944 4657
rect -904 4641 -870 4657
rect -830 4641 -796 4657
rect -756 4641 -722 4657
rect -682 4641 -648 4657
rect -608 4641 -574 4657
rect -534 4641 -500 4657
rect -460 4641 -426 4657
rect -386 4641 -352 4657
rect -312 4641 -278 4657
rect -238 4641 -204 4657
rect -1052 4623 -1048 4641
rect -1048 4623 -1018 4641
rect -1802 4551 -1768 4585
rect -1802 4476 -1768 4510
rect -978 4623 -946 4641
rect -946 4623 -944 4641
rect -904 4623 -878 4641
rect -878 4623 -870 4641
rect -830 4623 -810 4641
rect -810 4623 -796 4641
rect -756 4623 -742 4641
rect -742 4623 -722 4641
rect -682 4623 -674 4641
rect -674 4623 -648 4641
rect -608 4623 -606 4641
rect -606 4623 -574 4641
rect -534 4623 -504 4641
rect -504 4623 -500 4641
rect -460 4623 -436 4641
rect -436 4623 -426 4641
rect -386 4623 -368 4641
rect -368 4623 -352 4641
rect -312 4623 -300 4641
rect -300 4623 -278 4641
rect -238 4623 -232 4641
rect -232 4623 -204 4641
rect -1802 4401 -1768 4435
rect -1802 4326 -1768 4360
rect -1802 4251 -1768 4285
rect -1238 4471 -1204 4495
rect -1238 4461 -1207 4471
rect -1207 4461 -1204 4471
rect -1102 4434 -1068 4468
rect -1030 4455 -996 4468
rect -1030 4434 -996 4455
rect -874 4523 -840 4546
rect -874 4512 -840 4523
rect -874 4455 -840 4474
rect -874 4440 -840 4455
rect -790 4434 -756 4468
rect -718 4455 -684 4468
rect -718 4434 -684 4455
rect -562 4523 -528 4546
rect -562 4512 -528 4523
rect -562 4455 -528 4474
rect -562 4440 -528 4455
rect -232 4532 -198 4535
rect -232 4501 -198 4532
rect -1238 4369 -1207 4389
rect -1207 4369 -1204 4389
rect -1238 4355 -1204 4369
rect -948 4359 -914 4393
rect -1238 4267 -1204 4283
rect -1238 4249 -1207 4267
rect -1207 4249 -1204 4267
rect -1802 4176 -1768 4210
rect -1802 4101 -1768 4135
rect -1370 4118 -1336 4152
rect -1288 4118 -1254 4152
rect -1207 4118 -1173 4152
rect -1108 4319 -1074 4353
rect -1108 4226 -1074 4260
rect -636 4359 -602 4393
rect -948 4287 -914 4321
rect -948 4215 -914 4249
rect -796 4319 -762 4353
rect -796 4226 -762 4260
rect -1108 4133 -1074 4167
rect -636 4216 -602 4250
rect -484 4319 -450 4353
rect -484 4226 -450 4260
rect -796 4133 -762 4167
rect -484 4133 -450 4167
rect -232 4362 -198 4375
rect -410 4140 -376 4174
rect -1730 4062 -1717 4096
rect -1717 4062 -1696 4096
rect -1646 4062 -1615 4096
rect -1615 4062 -1612 4096
rect -328 4319 -294 4353
rect -328 4226 -294 4260
rect -328 4133 -294 4167
rect -232 4341 -198 4362
rect -232 4294 -198 4302
rect -232 4268 -198 4294
rect -232 4226 -198 4229
rect -232 4195 -198 4226
rect -410 4068 -376 4102
rect -1802 4028 -1768 4060
rect -1802 4026 -1768 4028
rect -232 4124 -198 4156
rect -232 4122 -198 4124
rect -232 4056 -198 4083
rect -232 4049 -198 4056
rect -852 3989 -848 4022
rect -848 3989 -818 4022
rect -775 3989 -773 4022
rect -773 3989 -741 4022
rect -698 3989 -697 4022
rect -697 3989 -664 4022
rect -621 3989 -587 4022
rect -852 3988 -818 3989
rect -775 3988 -741 3989
rect -698 3988 -664 3989
rect -621 3988 -587 3989
rect -545 3989 -511 4022
rect -545 3988 -511 3989
rect -232 3988 -198 4010
rect -1802 3960 -1768 3985
rect -1802 3951 -1768 3960
rect -232 3976 -198 3988
rect -1802 3892 -1768 3910
rect -1802 3876 -1768 3892
rect -1802 3824 -1768 3835
rect -1802 3801 -1768 3824
rect -1802 3756 -1768 3760
rect -1802 3726 -1768 3756
rect -1677 3902 -1643 3936
rect -1677 3830 -1643 3864
rect -1677 3758 -1643 3792
rect -1677 3685 -1643 3719
rect -1221 3902 -1187 3936
rect -1221 3821 -1187 3855
rect -232 3920 -198 3937
rect -232 3903 -198 3920
rect -232 3852 -198 3864
rect -1221 3740 -1187 3774
rect -1802 3654 -1768 3685
rect -1221 3659 -1187 3693
rect -1065 3803 -1031 3837
rect -753 3803 -719 3837
rect -1065 3731 -1031 3765
rect -909 3752 -875 3786
rect -1065 3659 -1031 3693
rect -987 3710 -953 3744
rect -1802 3651 -1768 3654
rect -1802 3586 -1768 3610
rect -1802 3576 -1768 3586
rect -987 3638 -953 3672
rect -909 3680 -875 3714
rect -753 3731 -719 3765
rect -753 3659 -719 3693
rect -640 3803 -606 3837
rect -640 3731 -606 3765
rect -640 3659 -606 3693
rect -484 3803 -450 3837
rect -484 3731 -450 3765
rect -484 3659 -450 3693
rect -328 3803 -294 3837
rect -328 3731 -294 3765
rect -328 3659 -294 3693
rect -232 3830 -198 3852
rect -232 3784 -198 3791
rect -232 3757 -198 3784
rect -232 3716 -198 3718
rect -232 3684 -198 3716
rect -909 3608 -875 3642
rect -232 3611 -198 3645
rect -1802 3518 -1768 3536
rect -1625 3523 -1616 3557
rect -1616 3523 -1591 3557
rect -1542 3523 -1512 3557
rect -1512 3523 -1508 3557
rect -1458 3523 -1442 3557
rect -1442 3523 -1424 3557
rect -1374 3523 -1372 3557
rect -1372 3523 -1340 3557
rect -1290 3523 -1266 3557
rect -1266 3523 -1256 3557
rect -1206 3523 -1196 3557
rect -1196 3523 -1172 3557
rect -1122 3523 -1092 3557
rect -1092 3523 -1088 3557
rect -232 3547 -198 3573
rect -232 3539 -198 3547
rect -1802 3502 -1768 3518
rect -1802 3450 -1768 3462
rect -1802 3428 -1768 3450
rect -1802 3382 -1768 3388
rect -232 3479 -198 3501
rect -232 3467 -198 3479
rect -232 3411 -198 3429
rect -232 3395 -198 3411
rect -1802 3354 -1768 3382
rect -1730 3348 -1700 3382
rect -1700 3348 -1696 3382
rect -1653 3348 -1632 3382
rect -1632 3348 -1619 3382
rect -1576 3348 -1564 3382
rect -1564 3348 -1542 3382
rect -1499 3348 -1496 3382
rect -1496 3348 -1465 3382
rect -1422 3348 -1394 3382
rect -1394 3348 -1388 3382
rect -1345 3348 -1326 3382
rect -1326 3348 -1311 3382
rect -1268 3348 -1258 3382
rect -1258 3348 -1234 3382
rect -1191 3348 -1190 3382
rect -1190 3348 -1157 3382
rect -1114 3348 -1088 3382
rect -1088 3348 -1080 3382
rect -1037 3348 -1020 3382
rect -1020 3348 -1003 3382
rect -960 3348 -952 3382
rect -952 3348 -926 3382
rect -883 3348 -850 3382
rect -850 3348 -849 3382
rect -806 3348 -782 3382
rect -782 3348 -772 3382
rect -729 3348 -714 3382
rect -714 3348 -695 3382
rect -652 3348 -618 3382
rect -580 3343 -546 3376
rect -580 3342 -546 3343
rect -580 3275 -546 3279
rect -580 3245 -546 3275
rect -232 3343 -198 3357
rect -232 3323 -198 3343
rect -232 3275 -198 3285
rect -232 3251 -198 3275
rect -232 3207 -198 3213
rect -574 3173 -546 3207
rect -546 3173 -540 3207
rect -484 3173 -478 3207
rect -478 3173 -450 3207
rect -394 3173 -376 3207
rect -376 3173 -360 3207
rect -304 3173 -270 3207
rect -232 3179 -198 3207
rect -14 4607 20 4641
rect 60 4607 88 4641
rect 88 4607 94 4641
rect 134 4607 156 4641
rect 156 4607 168 4641
rect 208 4607 224 4641
rect 224 4607 242 4641
rect 282 4607 292 4641
rect 292 4607 316 4641
rect 356 4607 360 4641
rect 360 4607 390 4641
rect 430 4607 462 4641
rect 462 4607 464 4641
rect 504 4607 530 4641
rect 530 4607 538 4641
rect 578 4607 598 4641
rect 598 4607 612 4641
rect 652 4607 666 4641
rect 666 4607 686 4641
rect 726 4607 734 4641
rect 734 4607 760 4641
rect 800 4607 802 4641
rect 802 4607 834 4641
rect 874 4607 904 4641
rect 904 4607 908 4641
rect 948 4607 972 4641
rect 972 4607 982 4641
rect 1022 4607 1040 4641
rect 1040 4607 1056 4641
rect 1096 4607 1108 4641
rect 1108 4607 1130 4641
rect 1171 4607 1176 4641
rect 1176 4607 1205 4641
rect 1246 4607 1278 4641
rect 1278 4607 1280 4641
rect 1321 4607 1346 4641
rect 1346 4607 1355 4641
rect 1396 4607 1414 4641
rect 1414 4607 1430 4641
rect 1471 4607 1482 4641
rect 1482 4607 1505 4641
rect 1546 4607 1550 4641
rect 1550 4607 1580 4641
rect -20 4505 -11 4535
rect -11 4505 14 4535
rect 182 4523 197 4557
rect 197 4523 216 4557
rect 258 4523 288 4557
rect 288 4523 292 4557
rect 1618 4601 1652 4635
rect -20 4501 14 4505
rect 1618 4553 1652 4562
rect 1618 4528 1652 4553
rect 1618 4485 1652 4489
rect 1618 4455 1652 4485
rect 1618 4383 1652 4416
rect 1618 4382 1652 4383
rect -20 4369 -11 4375
rect -11 4369 14 4375
rect -20 4341 14 4369
rect -20 4301 -11 4303
rect -11 4301 14 4303
rect -20 4269 14 4301
rect -20 4199 14 4231
rect -20 4197 -11 4199
rect -11 4197 14 4199
rect -20 4131 14 4159
rect -20 4125 -11 4131
rect -11 4125 14 4131
rect -20 4063 14 4087
rect -20 4053 -11 4063
rect -11 4053 14 4063
rect -20 3995 14 4015
rect -20 3981 -11 3995
rect -11 3981 14 3995
rect -20 3927 14 3943
rect -20 3909 -11 3927
rect -11 3909 14 3927
rect -20 3859 14 3871
rect -20 3837 -11 3859
rect -11 3837 14 3859
rect -20 3791 14 3799
rect -20 3765 -11 3791
rect -11 3765 14 3791
rect -20 3723 14 3727
rect -20 3693 -11 3723
rect -11 3693 14 3723
rect -20 3621 -11 3655
rect -11 3621 14 3655
rect -20 3553 -11 3583
rect -11 3553 14 3583
rect -20 3549 14 3553
rect -20 3485 -11 3511
rect -11 3485 14 3511
rect -20 3477 14 3485
rect -20 3417 -11 3439
rect -11 3417 14 3439
rect -20 3405 14 3417
rect -20 3349 -11 3367
rect -11 3349 14 3367
rect -20 3333 14 3349
rect -20 3281 -11 3295
rect -11 3281 14 3295
rect -20 3261 14 3281
rect -20 3213 -11 3223
rect -11 3213 14 3223
rect -20 3189 14 3213
rect -20 3145 -11 3151
rect -11 3145 14 3151
rect -20 3117 14 3145
rect -20 3077 -11 3079
rect -11 3077 14 3079
rect -20 3045 14 3077
rect -20 2975 14 3007
rect -20 2973 -11 2975
rect -11 2973 14 2975
rect -20 2907 14 2935
rect -20 2901 -11 2907
rect -11 2901 14 2907
rect -20 2839 14 2863
rect -20 2829 -11 2839
rect -11 2829 14 2839
rect -20 2771 14 2791
rect -20 2757 -11 2771
rect -11 2757 14 2771
rect -20 2703 14 2719
rect -20 2685 -11 2703
rect -11 2685 14 2703
rect -20 2635 14 2647
rect -20 2613 -11 2635
rect -11 2613 14 2635
rect -20 2567 14 2575
rect -20 2541 -11 2567
rect -11 2541 14 2567
rect -20 2469 14 2503
rect 1618 4315 1652 4343
rect 1618 4309 1652 4315
rect 1618 4247 1652 4270
rect 1618 4236 1652 4247
rect 1618 4179 1652 4197
rect 1618 4163 1652 4179
rect 1618 4111 1652 4124
rect 1618 4090 1652 4111
rect 1618 4043 1652 4051
rect 1618 4017 1652 4043
rect 1618 3975 1652 3977
rect 1618 3943 1652 3975
rect 1618 3873 1652 3903
rect 1618 3869 1652 3873
rect 1618 3805 1652 3829
rect 1618 3795 1652 3805
rect 1618 3737 1652 3755
rect 1618 3721 1652 3737
rect 1618 3669 1652 3681
rect 1618 3647 1652 3669
rect 1618 3601 1652 3607
rect 1618 3573 1652 3601
rect 1618 3499 1652 3533
rect 1618 3431 1652 3459
rect 1618 3425 1652 3431
rect 1618 3363 1652 3385
rect 1618 3351 1652 3363
rect 1618 3295 1652 3311
rect 1618 3277 1652 3295
rect 1618 3227 1652 3237
rect 1618 3203 1652 3227
rect 1618 3159 1652 3163
rect 1618 3129 1652 3159
rect 1618 3057 1652 3089
rect 1618 3055 1652 3057
rect 1618 2989 1652 3015
rect 1618 2981 1652 2989
rect 1618 2921 1652 2941
rect 1618 2907 1652 2921
rect 1618 2853 1652 2867
rect 1618 2833 1652 2853
rect 1618 2785 1652 2793
rect 1618 2759 1652 2785
rect 1618 2717 1652 2719
rect 1618 2685 1652 2717
rect 1618 2615 1652 2645
rect 1618 2611 1652 2615
rect 1618 2547 1652 2571
rect 1618 2537 1652 2547
rect -20 2397 14 2431
rect 182 2453 216 2487
rect 258 2453 292 2487
rect 1618 2479 1652 2497
rect 1618 2463 1652 2479
rect -20 2325 14 2359
rect 1618 2411 1652 2423
rect 1618 2389 1652 2411
rect 1618 2343 1652 2349
rect 198 2309 224 2343
rect 224 2309 232 2343
rect 272 2309 292 2343
rect 292 2309 306 2343
rect 346 2309 360 2343
rect 360 2309 380 2343
rect 420 2309 428 2343
rect 428 2309 454 2343
rect 494 2309 496 2343
rect 496 2309 528 2343
rect 568 2309 598 2343
rect 598 2309 602 2343
rect 642 2309 666 2343
rect 666 2309 676 2343
rect 716 2309 734 2343
rect 734 2309 750 2343
rect 790 2309 802 2343
rect 802 2309 824 2343
rect 864 2309 870 2343
rect 870 2309 898 2343
rect 938 2309 972 2343
rect 1012 2309 1040 2343
rect 1040 2309 1046 2343
rect 1087 2309 1108 2343
rect 1108 2309 1121 2343
rect 1618 2315 1652 2343
rect 1709 2336 1743 2343
rect 1709 2309 1720 2336
rect 1720 2309 1743 2336
rect -20 2269 -11 2287
rect -11 2269 14 2287
rect -20 2253 14 2269
rect -20 2201 -11 2214
rect -11 2201 14 2214
rect -20 2180 14 2201
rect 251 2180 285 2214
rect -20 2133 -11 2141
rect -11 2133 14 2141
rect -20 2107 14 2133
rect -20 2065 -11 2068
rect -11 2065 14 2068
rect -20 2034 14 2065
rect -20 1963 14 1995
rect -20 1961 -11 1963
rect -11 1961 14 1963
rect -20 1895 14 1922
rect -20 1888 -11 1895
rect -11 1888 14 1895
rect -20 1827 14 1849
rect -20 1815 -11 1827
rect -11 1815 14 1827
rect 74 2141 108 2175
rect 74 2055 108 2089
rect 74 1969 108 2003
rect 74 1883 108 1917
rect 74 1796 108 1830
rect 251 2104 285 2138
rect 251 2027 285 2061
rect 251 1950 285 1984
rect 251 1873 285 1907
rect 251 1796 285 1830
rect 445 2001 479 2035
rect 445 1917 479 1951
rect 445 1833 479 1867
rect 445 1749 479 1783
rect 445 1665 479 1699
rect 721 2241 755 2271
rect 721 2237 755 2241
rect 602 2180 636 2214
rect 721 2173 755 2187
rect 721 2153 755 2173
rect 1855 2271 1889 2305
rect 1855 2206 1889 2231
rect 1855 2197 1889 2206
rect 602 2107 636 2141
rect 980 2115 987 2149
rect 987 2115 1014 2149
rect 1057 2115 1089 2149
rect 1089 2115 1091 2149
rect 1134 2115 1157 2149
rect 1157 2115 1168 2149
rect 1211 2115 1225 2149
rect 1225 2115 1245 2149
rect 1288 2115 1293 2149
rect 1293 2115 1322 2149
rect 1365 2115 1395 2149
rect 1395 2115 1399 2149
rect 1442 2115 1463 2149
rect 1463 2115 1476 2149
rect 1519 2115 1531 2149
rect 1531 2115 1553 2149
rect 1596 2115 1599 2149
rect 1599 2115 1630 2149
rect 1668 2115 1702 2143
rect 721 2071 755 2103
rect 721 2069 755 2071
rect 602 2033 636 2067
rect 1668 2109 1702 2115
rect 721 2003 755 2020
rect 602 1959 636 1993
rect 721 1986 755 2003
rect 1160 2019 1194 2053
rect 721 1935 755 1937
rect 602 1885 636 1919
rect 721 1903 755 1935
rect 602 1811 636 1845
rect 721 1833 755 1854
rect 721 1820 755 1833
rect 602 1737 636 1771
rect 721 1765 755 1771
rect 721 1737 755 1765
rect 721 1595 755 1613
rect 120 1553 121 1587
rect 121 1553 154 1587
rect 202 1553 223 1587
rect 223 1553 236 1587
rect 392 1553 421 1587
rect 421 1553 426 1587
rect 470 1553 498 1587
rect 498 1553 504 1587
rect 548 1553 575 1587
rect 575 1553 582 1587
rect 721 1579 755 1595
rect 721 1527 755 1535
rect 1004 1965 1038 1999
rect 1004 1892 1038 1926
rect 1004 1819 1038 1853
rect 1004 1746 1038 1780
rect 1004 1673 1038 1707
rect 1004 1600 1038 1634
rect 1160 1942 1194 1976
rect 1160 1866 1194 1900
rect 1160 1790 1194 1824
rect 1160 1714 1194 1748
rect 1160 1638 1194 1672
rect 1160 1562 1194 1596
rect 1316 2000 1350 2034
rect 1316 1921 1350 1955
rect 1316 1842 1350 1876
rect 1316 1763 1350 1797
rect 1316 1684 1350 1718
rect 1572 2019 1606 2053
rect 1572 1945 1606 1979
rect 1572 1871 1606 1905
rect 1572 1797 1606 1831
rect 1572 1724 1606 1758
rect 1572 1651 1606 1685
rect 1668 2047 1702 2062
rect 1668 2028 1702 2047
rect 1668 1979 1702 1981
rect 1668 1947 1702 1979
rect 1668 1877 1702 1900
rect 1668 1866 1702 1877
rect 1668 1809 1702 1820
rect 1668 1786 1702 1809
rect 1668 1707 1702 1740
rect 1668 1706 1702 1707
rect 1316 1605 1350 1639
rect 1004 1527 1038 1561
rect 1316 1527 1350 1561
rect 1668 1639 1702 1660
rect 1668 1626 1702 1639
rect 1668 1571 1702 1580
rect 1668 1546 1702 1571
rect 721 1501 755 1527
rect 157 1445 185 1479
rect 185 1445 191 1479
rect 289 1445 319 1479
rect 319 1445 323 1479
rect 403 1445 407 1479
rect 407 1445 437 1479
rect 487 1445 521 1479
rect 1855 2135 1889 2157
rect 1855 2123 1889 2135
rect 1855 2064 1889 2083
rect 1855 2049 1889 2064
rect 1855 1993 1889 2009
rect 1855 1975 1889 1993
rect 1855 1922 1889 1935
rect 1855 1901 1889 1922
rect 1855 1851 1889 1861
rect 1855 1827 1889 1851
rect 1855 1780 1889 1787
rect 1855 1753 1889 1780
rect 1855 1709 1889 1713
rect 1855 1679 1889 1709
rect 1855 1638 1889 1639
rect 1855 1605 1889 1638
rect 1855 1531 1889 1565
rect 721 1425 755 1457
rect 721 1423 755 1425
rect -20 1385 -11 1393
rect -11 1385 14 1393
rect -20 1359 14 1385
rect 1855 1459 1889 1491
rect 1855 1457 1889 1459
rect 721 1357 755 1380
rect 1088 1379 1092 1409
rect 1092 1379 1122 1409
rect 1170 1379 1194 1409
rect 1194 1379 1204 1409
rect 1252 1379 1262 1409
rect 1262 1379 1286 1409
rect 1088 1375 1122 1379
rect 1170 1375 1204 1379
rect 1252 1375 1286 1379
rect 1334 1375 1368 1409
rect 1416 1379 1444 1409
rect 1444 1379 1450 1409
rect 1498 1379 1512 1409
rect 1512 1379 1532 1409
rect 1416 1375 1450 1379
rect 1498 1375 1532 1379
rect 1579 1375 1613 1409
rect 1855 1388 1889 1417
rect 1855 1383 1889 1388
rect 721 1346 755 1357
rect -20 1317 -11 1321
rect -11 1317 14 1321
rect -20 1287 14 1317
rect -20 1215 14 1249
rect -20 1147 14 1177
rect -20 1143 -11 1147
rect -11 1143 14 1147
rect -20 1079 14 1105
rect -20 1071 -11 1079
rect -11 1071 14 1079
rect -20 1011 14 1033
rect -20 999 -11 1011
rect -11 999 14 1011
rect -20 943 14 961
rect -20 927 -11 943
rect -11 927 14 943
rect -20 875 14 889
rect -20 855 -11 875
rect -11 855 14 875
rect -20 807 14 817
rect -20 783 -11 807
rect -11 783 14 807
rect 90 1309 124 1343
rect 90 1236 124 1270
rect 90 1163 124 1197
rect 602 1309 636 1343
rect 721 1289 755 1303
rect 602 1237 636 1271
rect 721 1269 755 1289
rect 1855 1309 1889 1343
rect 721 1221 755 1226
rect 602 1165 636 1199
rect 721 1192 755 1221
rect 90 1089 124 1123
rect 90 1015 124 1049
rect 90 941 124 975
rect 90 867 124 901
rect 90 793 124 827
rect 346 1131 380 1165
rect 346 1052 380 1086
rect 346 972 380 1006
rect 346 892 380 926
rect 346 812 380 846
rect 602 1093 636 1127
rect 721 1119 755 1149
rect 721 1115 755 1119
rect 602 1021 636 1055
rect 721 1051 755 1072
rect 721 1038 755 1051
rect 1855 1236 1889 1270
rect 1855 1163 1889 1197
rect 1855 1090 1889 1124
rect 1855 1017 1889 1051
rect 721 983 755 995
rect 602 949 636 983
rect 721 961 755 983
rect 721 915 755 918
rect 602 877 636 911
rect 721 884 755 915
rect 1855 948 1889 978
rect 1855 944 1889 948
rect 1088 887 1122 891
rect 1170 887 1204 891
rect 1252 887 1286 891
rect 1088 857 1092 887
rect 1092 857 1122 887
rect 1170 857 1194 887
rect 1194 857 1204 887
rect 1252 857 1262 887
rect 1262 857 1286 887
rect 1334 857 1368 891
rect 1416 887 1450 891
rect 1498 887 1532 891
rect 1416 857 1444 887
rect 1444 857 1450 887
rect 1498 857 1512 887
rect 1512 857 1532 887
rect 1579 857 1613 891
rect 1855 875 1889 905
rect 1855 871 1889 875
rect 602 805 636 839
rect 721 813 755 841
rect 721 807 755 813
rect -20 739 14 745
rect -20 711 -11 739
rect -11 711 14 739
rect 721 745 755 764
rect 721 730 755 745
rect 117 679 121 713
rect 121 679 151 713
rect 202 679 223 713
rect 223 679 236 713
rect 389 679 421 713
rect 421 679 423 713
rect 467 679 498 713
rect 498 679 501 713
rect 545 679 575 713
rect 575 679 579 713
rect -20 671 14 673
rect -20 639 -11 671
rect -11 639 14 671
rect 721 677 755 687
rect 721 653 755 677
rect -20 569 -11 601
rect -11 569 14 601
rect -20 567 14 569
rect -20 501 -11 529
rect -11 501 14 529
rect -20 495 14 501
rect -20 433 -11 457
rect -11 433 14 457
rect -20 423 14 433
rect -20 365 -11 384
rect -11 365 14 384
rect -20 350 14 365
rect -20 297 -11 311
rect -11 297 14 311
rect -20 277 14 297
rect -20 229 -11 238
rect -11 229 14 238
rect -20 204 14 229
rect -20 161 -11 165
rect -11 161 14 165
rect -20 131 14 161
rect -20 59 14 92
rect -20 58 -11 59
rect -11 58 14 59
rect 74 534 108 568
rect 439 567 473 601
rect 74 453 108 487
rect 74 372 108 406
rect 74 292 108 326
rect 74 212 108 246
rect 250 467 284 501
rect 250 377 284 411
rect 250 287 284 321
rect 250 197 284 231
rect 439 494 473 528
rect 439 422 473 456
rect 439 350 473 384
rect 74 132 108 166
rect 74 52 108 86
rect 602 495 636 529
rect 721 507 755 529
rect 721 495 755 507
rect 602 419 636 453
rect 721 439 755 446
rect 721 412 755 439
rect 602 343 636 377
rect 721 337 755 363
rect 721 329 755 337
rect 602 268 636 302
rect 721 269 755 280
rect 721 246 755 269
rect 602 193 636 227
rect 721 167 755 197
rect 721 163 755 167
rect 602 118 636 152
rect 908 737 942 739
rect 908 705 942 737
rect 908 635 942 667
rect 908 633 942 635
rect 908 567 942 595
rect 908 561 942 567
rect 908 499 942 522
rect 908 488 942 499
rect 908 431 942 449
rect 908 415 942 431
rect 908 363 942 376
rect 908 342 942 363
rect 908 295 942 303
rect 908 269 942 295
rect 1004 705 1038 739
rect 1316 705 1350 739
rect 1004 632 1038 666
rect 1004 559 1038 593
rect 1004 486 1038 520
rect 1004 412 1038 446
rect 1004 338 1038 372
rect 1004 264 1038 298
rect 1160 670 1194 704
rect 1160 594 1194 628
rect 1160 518 1194 552
rect 1160 442 1194 476
rect 1160 366 1194 400
rect 1160 290 1194 324
rect 908 196 942 230
rect 1160 213 1194 247
rect 1316 627 1350 661
rect 1668 695 1702 720
rect 1668 686 1702 695
rect 1668 627 1702 640
rect 1316 548 1350 582
rect 1316 469 1350 503
rect 1316 390 1350 424
rect 1316 311 1350 345
rect 1316 232 1350 266
rect 1572 581 1606 615
rect 1572 508 1606 542
rect 1572 435 1606 469
rect 1572 361 1606 395
rect 1572 287 1606 321
rect 1572 213 1606 247
rect 1668 606 1702 627
rect 1668 559 1702 560
rect 1668 526 1702 559
rect 1668 457 1702 480
rect 1668 446 1702 457
rect 1668 389 1702 400
rect 1668 366 1702 389
rect 1668 287 1702 319
rect 1668 285 1702 287
rect 1668 219 1702 238
rect 908 123 942 157
rect 1668 204 1702 219
rect 1668 151 1702 157
rect 980 117 1010 151
rect 1010 117 1014 151
rect 1057 117 1078 151
rect 1078 117 1091 151
rect 1134 117 1146 151
rect 1146 117 1168 151
rect 1211 117 1214 151
rect 1214 117 1245 151
rect 1288 117 1316 151
rect 1316 117 1322 151
rect 1365 117 1384 151
rect 1384 117 1399 151
rect 1442 117 1452 151
rect 1452 117 1476 151
rect 1519 117 1520 151
rect 1520 117 1553 151
rect 1596 117 1630 151
rect 1668 123 1702 151
rect 1855 802 1889 832
rect 1855 798 1889 802
rect 1855 729 1889 759
rect 1855 725 1889 729
rect 1855 656 1889 686
rect 1855 652 1889 656
rect 1855 583 1889 613
rect 1855 579 1889 583
rect 1855 511 1889 540
rect 1855 506 1889 511
rect 1855 439 1889 467
rect 1855 433 1889 439
rect 1855 367 1889 394
rect 1855 360 1889 367
rect 1855 295 1889 321
rect 1855 287 1889 295
rect 1855 223 1889 248
rect 1855 214 1889 223
rect 1855 151 1889 175
rect 1855 141 1889 151
rect 721 99 755 114
rect 721 80 755 99
rect 721 -3 755 31
rect 1855 79 1889 102
rect 1855 68 1889 79
rect 1855 7 1889 29
rect 1855 -5 1889 7
<< metal1 >>
rect -1157 5023 -1151 5075
rect -1099 5023 -1074 5075
rect -1022 5023 -996 5075
rect -944 5023 2001 5075
rect 2053 5023 2072 5075
rect 2124 5023 2144 5075
rect 2196 5023 2216 5075
rect 2268 5023 2288 5075
rect 2340 5023 2346 5075
rect -1157 5011 2346 5023
rect -1157 4959 -1151 5011
rect -1099 4959 -1074 5011
rect -1022 4959 -996 5011
rect -944 4959 2001 5011
rect 2053 4959 2072 5011
rect 2124 4959 2144 5011
rect 2196 4959 2216 5011
rect 2268 4959 2288 5011
rect 2340 4959 2346 5011
rect -748 4893 -696 4899
rect -659 4851 -653 4903
rect -601 4851 -589 4903
rect -537 4851 277 4903
rect 329 4851 341 4903
rect 393 4851 405 4903
rect 457 4851 463 4903
rect -748 4829 -696 4841
rect -882 4813 -830 4819
tri -696 4823 -671 4848 sw
rect -696 4777 832 4823
rect -748 4771 832 4777
rect 884 4771 896 4823
rect 948 4771 954 4823
rect -882 4749 -830 4761
tri -830 4743 -805 4768 sw
rect -830 4697 750 4743
rect -882 4691 750 4697
rect 802 4691 814 4743
rect 866 4691 872 4743
rect -1808 4657 -192 4663
rect -1808 4623 -1796 4657
rect -1762 4623 -1721 4657
rect -1687 4623 -1646 4657
rect -1612 4623 -1571 4657
rect -1537 4623 -1496 4657
rect -1462 4623 -1422 4657
rect -1388 4623 -1348 4657
rect -1314 4623 -1274 4657
rect -1240 4623 -1200 4657
rect -1166 4623 -1126 4657
rect -1092 4623 -1052 4657
rect -1018 4623 -978 4657
rect -944 4623 -904 4657
rect -870 4623 -830 4657
rect -796 4623 -756 4657
rect -722 4623 -682 4657
rect -648 4623 -608 4657
rect -574 4623 -534 4657
rect -500 4623 -460 4657
rect -426 4623 -386 4657
rect -352 4623 -312 4657
rect -278 4623 -238 4657
rect -204 4623 -192 4657
tri 511 4647 517 4653 se
rect 517 4647 523 4653
rect -1808 4617 -192 4623
rect -1808 4607 -1745 4617
tri -1745 4607 -1735 4617 nw
tri -263 4607 -253 4617 ne
rect -253 4607 -192 4617
rect -1808 4601 -1751 4607
tri -1751 4601 -1745 4607 nw
tri -253 4601 -247 4607 ne
rect -247 4601 -192 4607
rect -1808 4592 -1760 4601
tri -1760 4592 -1751 4601 nw
tri -247 4592 -238 4601 ne
rect -1808 4585 -1762 4592
tri -1762 4590 -1760 4592 nw
rect -1808 4551 -1802 4585
rect -1768 4551 -1762 4585
rect -1808 4512 -1762 4551
rect -1568 4588 -522 4589
rect -1568 4536 -1562 4588
rect -1510 4536 -1498 4588
rect -1446 4560 -522 4588
rect -1446 4557 -1124 4560
tri -1124 4557 -1121 4560 nw
tri -1080 4557 -1077 4560 ne
rect -1077 4557 -987 4560
tri -987 4557 -984 4560 nw
tri -905 4557 -902 4560 ne
rect -902 4557 -812 4560
tri -812 4557 -809 4560 nw
tri -768 4557 -765 4560 ne
rect -765 4557 -675 4560
tri -675 4557 -672 4560 nw
tri -593 4557 -590 4560 ne
rect -590 4557 -522 4560
rect -1446 4546 -1135 4557
tri -1135 4546 -1124 4557 nw
tri -1077 4546 -1066 4557 ne
rect -1066 4546 -998 4557
tri -998 4546 -987 4557 nw
tri -902 4546 -891 4557 ne
rect -891 4546 -823 4557
tri -823 4546 -812 4557 nw
tri -765 4546 -754 4557 ne
rect -754 4546 -686 4557
tri -686 4546 -675 4557 nw
tri -590 4546 -579 4557 ne
rect -579 4546 -522 4557
rect -1446 4536 -1145 4546
tri -1145 4536 -1135 4546 nw
tri -1066 4536 -1056 4546 ne
rect -1056 4537 -1007 4546
tri -1007 4537 -998 4546 nw
tri -891 4537 -882 4546 ne
rect -882 4537 -874 4546
rect -1056 4536 -1055 4537
rect -1009 4536 -1008 4537
tri -1008 4536 -1007 4537 nw
tri -882 4536 -881 4537 ne
rect -881 4536 -874 4537
rect -1568 4535 -1146 4536
tri -1146 4535 -1145 4536 nw
tri -1056 4535 -1055 4536 ne
rect -1054 4535 -1010 4536
tri -1009 4535 -1008 4536 nw
tri -881 4535 -880 4536 ne
tri -1762 4512 -1742 4532 sw
rect -880 4512 -874 4536
rect -840 4512 -834 4546
tri -834 4535 -823 4546 nw
tri -754 4535 -743 4546 ne
rect -743 4537 -695 4546
tri -695 4537 -686 4546 nw
tri -579 4537 -570 4546 ne
rect -570 4537 -562 4546
rect -697 4536 -696 4537
tri -696 4536 -695 4537 nw
tri -570 4536 -569 4537 ne
rect -569 4536 -562 4537
rect -742 4535 -698 4536
tri -697 4535 -696 4536 nw
tri -569 4535 -568 4536 ne
rect -1808 4510 -1742 4512
rect -1808 4476 -1802 4510
rect -1768 4507 -1742 4510
tri -1742 4507 -1737 4512 sw
rect -1768 4495 -1198 4507
rect -1768 4476 -1238 4495
rect -1808 4461 -1238 4476
rect -1204 4461 -1198 4495
tri -1065 4489 -1055 4499 se
rect -1054 4498 -1010 4499
tri -1009 4498 -1008 4499 sw
rect -1009 4497 -1008 4498
tri -1008 4497 -1007 4498 sw
rect -1055 4489 -1007 4497
tri -1007 4489 -999 4497 sw
tri -1080 4474 -1065 4489 se
rect -1065 4474 -999 4489
tri -999 4474 -984 4489 sw
rect -1808 4435 -1198 4461
rect -1808 4401 -1802 4435
rect -1768 4401 -1198 4435
rect -1808 4389 -1198 4401
rect -1808 4372 -1238 4389
rect -1808 4360 -1745 4372
rect -1808 4326 -1802 4360
rect -1768 4355 -1745 4360
tri -1745 4355 -1728 4372 nw
tri -1576 4355 -1559 4372 ne
rect -1559 4355 -1238 4372
rect -1204 4359 -1198 4389
rect -1114 4468 -984 4474
rect -1114 4434 -1102 4468
rect -1068 4434 -1030 4468
rect -996 4434 -984 4468
rect -1114 4428 -984 4434
rect -880 4474 -834 4512
rect -568 4512 -562 4536
rect -528 4512 -522 4546
tri -753 4489 -743 4499 se
rect -742 4498 -698 4499
tri -697 4498 -696 4499 sw
rect -697 4497 -696 4498
tri -696 4497 -695 4498 sw
rect -743 4489 -695 4497
tri -695 4489 -687 4497 sw
tri -768 4474 -753 4489 se
rect -753 4474 -687 4489
tri -687 4474 -672 4489 sw
rect -880 4440 -874 4474
rect -840 4440 -834 4474
rect -880 4428 -834 4440
rect -802 4468 -672 4474
rect -802 4434 -790 4468
rect -756 4434 -718 4468
rect -684 4434 -672 4468
rect -802 4428 -672 4434
rect -568 4474 -522 4512
rect -238 4535 -192 4601
rect -238 4501 -232 4535
rect -198 4501 -192 4535
rect -238 4489 -192 4501
rect -26 4641 523 4647
rect 575 4641 590 4653
rect 642 4641 658 4653
rect 710 4647 716 4653
tri 716 4647 722 4653 sw
rect 710 4641 1658 4647
rect -26 4607 -14 4641
rect 20 4607 60 4641
rect 94 4607 134 4641
rect 168 4607 208 4641
rect 242 4607 282 4641
rect 316 4607 356 4641
rect 390 4607 430 4641
rect 464 4607 504 4641
rect 575 4607 578 4641
rect 642 4607 652 4641
rect 710 4607 726 4641
rect 760 4607 800 4641
rect 834 4607 874 4641
rect 908 4607 948 4641
rect 982 4607 1022 4641
rect 1056 4607 1096 4641
rect 1130 4607 1171 4641
rect 1205 4607 1246 4641
rect 1280 4607 1321 4641
rect 1355 4607 1396 4641
rect 1430 4607 1471 4641
rect 1505 4607 1546 4641
rect 1580 4635 1658 4641
rect 1580 4607 1618 4635
rect -26 4601 523 4607
rect 575 4601 590 4607
rect 642 4601 658 4607
rect 710 4601 1618 4607
rect 1652 4601 1658 4635
rect -26 4589 33 4601
tri 33 4589 45 4601 nw
tri 1587 4589 1599 4601 ne
rect 1599 4589 1658 4601
rect -26 4535 20 4589
tri 20 4576 33 4589 nw
tri 1599 4576 1612 4589 ne
rect -26 4501 -20 4535
rect 14 4501 20 4535
rect -26 4489 20 4501
rect 170 4557 277 4573
rect 170 4523 182 4557
rect 216 4523 258 4557
rect 170 4521 277 4523
rect 329 4521 341 4573
rect 393 4521 405 4573
rect 457 4545 1306 4573
rect 457 4535 477 4545
tri 477 4535 487 4545 nw
tri 1204 4535 1214 4545 ne
rect 1214 4535 1306 4545
rect 457 4528 470 4535
tri 470 4528 477 4535 nw
tri 1214 4528 1221 4535 ne
rect 1221 4528 1306 4535
rect 457 4521 463 4528
tri 463 4521 470 4528 nw
tri 1221 4521 1228 4528 ne
rect 1228 4521 1306 4528
rect 170 4517 304 4521
tri 304 4517 308 4521 nw
tri 1228 4517 1232 4521 ne
rect 1232 4517 1306 4521
tri 170 4499 188 4517 ne
rect 188 4499 276 4517
tri 188 4489 198 4499 ne
rect 198 4489 276 4499
tri 276 4489 304 4517 nw
rect 568 4489 922 4517
tri 922 4489 950 4517 sw
tri 1232 4489 1260 4517 ne
rect -568 4440 -562 4474
rect -528 4440 -522 4474
tri 198 4473 214 4489 ne
rect -568 4428 -522 4440
rect -1114 4416 -1055 4428
tri -1055 4416 -1043 4428 nw
rect -802 4416 -743 4428
tri -743 4416 -731 4428 nw
rect -1114 4405 -1066 4416
tri -1066 4405 -1055 4416 nw
rect -802 4405 -754 4416
tri -754 4405 -743 4416 nw
rect -342 4415 96 4461
rect -1068 4404 -1067 4405
tri -1067 4404 -1066 4405 nw
rect -1113 4403 -1069 4404
tri -1068 4403 -1067 4404 nw
rect -1114 4367 -1068 4403
tri -1198 4359 -1190 4367 sw
tri -1122 4359 -1114 4367 se
rect -1113 4366 -1069 4367
rect -1114 4359 -1068 4365
rect -1204 4355 -1190 4359
rect -1768 4353 -1747 4355
tri -1747 4353 -1745 4355 nw
tri -1559 4353 -1557 4355 ne
rect -1557 4353 -1190 4355
tri -1190 4353 -1184 4359 sw
tri -1128 4353 -1122 4359 se
rect -1122 4353 -1068 4359
rect -1768 4326 -1762 4353
tri -1762 4338 -1747 4353 nw
tri -1557 4338 -1542 4353 ne
rect -1542 4342 -1184 4353
tri -1184 4342 -1173 4353 sw
tri -1139 4342 -1128 4353 se
rect -1128 4342 -1108 4353
rect -1542 4338 -1108 4342
rect -1808 4285 -1762 4326
tri -1542 4319 -1523 4338 ne
rect -1523 4319 -1108 4338
rect -1074 4319 -1068 4353
tri -1523 4316 -1520 4319 ne
rect -1520 4316 -1068 4319
rect -1808 4251 -1802 4285
rect -1768 4251 -1762 4285
rect -1652 4310 -1600 4316
rect -1808 4249 -1762 4251
tri -1762 4249 -1743 4268 sw
tri -1671 4249 -1652 4268 se
tri -1520 4287 -1491 4316 ne
rect -1491 4287 -1068 4316
tri -1491 4283 -1487 4287 ne
rect -1487 4283 -1068 4287
tri -1487 4266 -1470 4283 ne
rect -1470 4266 -1238 4283
rect -1652 4249 -1600 4258
tri -1600 4249 -1583 4266 sw
tri -1470 4249 -1453 4266 ne
rect -1453 4249 -1238 4266
rect -1204 4260 -1068 4283
rect -1204 4249 -1108 4260
rect -1808 4243 -1743 4249
tri -1743 4243 -1737 4249 sw
tri -1677 4243 -1671 4249 se
rect -1671 4244 -1583 4249
rect -1671 4243 -1652 4244
rect -1808 4210 -1739 4243
rect -1808 4176 -1802 4210
rect -1768 4186 -1739 4210
rect -1738 4187 -1737 4242
rect -1701 4187 -1700 4242
rect -1699 4192 -1652 4243
rect -1600 4243 -1583 4244
tri -1583 4243 -1577 4249 sw
tri -1453 4243 -1447 4249 ne
rect -1447 4243 -1108 4249
rect -1600 4242 -1577 4243
tri -1577 4242 -1576 4243 sw
tri -1447 4242 -1446 4243 ne
rect -1446 4242 -1108 4243
rect -1600 4237 -1576 4242
tri -1576 4237 -1571 4242 sw
tri -1446 4237 -1441 4242 ne
rect -1441 4237 -1108 4242
rect -1600 4226 -1571 4237
tri -1571 4226 -1560 4237 sw
tri -1441 4226 -1430 4237 ne
rect -1430 4226 -1108 4237
rect -1074 4226 -1068 4260
rect -1600 4215 -1560 4226
tri -1560 4215 -1549 4226 sw
tri -1430 4215 -1419 4226 ne
rect -1419 4215 -1068 4226
rect -1600 4204 -1549 4215
tri -1549 4204 -1538 4215 sw
tri -1419 4204 -1408 4215 ne
rect -1408 4204 -1068 4215
rect -954 4393 -908 4405
tri -908 4393 -896 4405 sw
rect -756 4404 -755 4405
tri -755 4404 -754 4405 nw
tri -643 4404 -642 4405 se
rect -642 4404 -596 4405
rect -801 4403 -757 4404
tri -756 4403 -755 4404 nw
tri -644 4403 -643 4404 se
rect -643 4403 -596 4404
rect -954 4359 -948 4393
rect -914 4387 -896 4393
tri -896 4387 -890 4393 sw
rect -914 4381 -830 4387
rect -914 4359 -882 4381
rect -954 4329 -882 4359
rect -954 4321 -830 4329
rect -954 4287 -948 4321
rect -914 4299 -830 4321
rect -914 4287 -882 4299
rect -954 4249 -882 4287
rect -954 4215 -948 4249
rect -914 4247 -882 4249
rect -914 4241 -830 4247
rect -914 4226 -845 4241
tri -845 4226 -830 4241 nw
rect -802 4367 -756 4403
tri -654 4393 -644 4403 se
rect -644 4393 -596 4403
tri -660 4387 -654 4393 se
rect -654 4387 -636 4393
rect -801 4366 -757 4367
rect -802 4353 -756 4365
rect -802 4319 -796 4353
rect -762 4319 -756 4353
rect -802 4260 -756 4319
rect -802 4226 -796 4260
rect -762 4226 -756 4260
rect -914 4216 -855 4226
tri -855 4216 -845 4226 nw
rect -914 4215 -858 4216
rect -954 4213 -858 4215
tri -858 4213 -855 4216 nw
rect -1600 4195 -1538 4204
tri -1538 4195 -1529 4204 sw
tri -1408 4195 -1399 4204 ne
rect -1399 4195 -1068 4204
tri -1068 4195 -1050 4213 sw
rect -954 4203 -868 4213
tri -868 4203 -858 4213 nw
tri -812 4203 -802 4213 se
rect -802 4203 -756 4226
rect -668 4381 -636 4387
rect -602 4359 -596 4393
rect -616 4329 -596 4359
rect -668 4262 -596 4329
rect -616 4250 -596 4262
rect -602 4216 -596 4250
tri -820 4195 -812 4203 se
rect -812 4200 -756 4203
tri -756 4200 -743 4213 sw
rect -616 4210 -596 4216
rect -668 4204 -596 4210
rect -560 4359 -444 4365
rect -508 4307 -496 4359
rect -560 4269 -444 4307
rect -508 4217 -496 4269
rect -812 4195 -743 4200
tri -743 4195 -738 4200 sw
tri -565 4195 -560 4200 se
rect -560 4195 -444 4217
rect -1600 4192 -1529 4195
rect -1699 4186 -1529 4192
tri -1529 4186 -1520 4195 sw
tri -1399 4186 -1390 4195 ne
rect -1390 4186 -1050 4195
rect -1768 4178 -1745 4186
tri -1745 4178 -1737 4186 nw
tri -1560 4178 -1552 4186 ne
rect -1552 4178 -1520 4186
tri -1520 4178 -1512 4186 sw
tri -1390 4178 -1382 4186 ne
rect -1768 4176 -1749 4178
rect -1808 4174 -1749 4176
tri -1749 4174 -1745 4178 nw
tri -1552 4174 -1548 4178 ne
rect -1548 4174 -1512 4178
tri -1512 4174 -1508 4178 sw
rect -1382 4175 -1050 4186
tri -1050 4175 -1030 4195 sw
tri -840 4175 -820 4195 se
rect -820 4175 -738 4195
tri -738 4175 -718 4195 sw
tri -585 4175 -565 4195 se
rect -565 4179 -444 4195
rect -342 4353 -288 4415
tri -288 4390 -263 4415 nw
tri 71 4390 96 4415 ne
rect -342 4319 -328 4353
rect -294 4319 -288 4353
rect -342 4260 -288 4319
rect -342 4226 -328 4260
rect -294 4226 -288 4260
rect -565 4175 -560 4179
rect -1808 4167 -1756 4174
tri -1756 4167 -1749 4174 nw
tri -1548 4167 -1541 4174 ne
rect -1541 4167 -1508 4174
tri -1508 4167 -1501 4174 sw
rect -1382 4167 -560 4175
rect -1808 4164 -1759 4167
tri -1759 4164 -1756 4167 nw
tri -1541 4164 -1538 4167 ne
rect -1538 4164 -1501 4167
tri -1501 4164 -1498 4167 sw
rect -1808 4135 -1762 4164
tri -1762 4161 -1759 4164 nw
tri -1538 4161 -1535 4164 ne
rect -1535 4161 -1498 4164
tri -1535 4152 -1526 4161 ne
rect -1526 4158 -1498 4161
tri -1498 4158 -1492 4164 sw
rect -1526 4152 -1492 4158
tri -1492 4152 -1486 4158 sw
rect -1382 4152 -1108 4167
rect -1808 4101 -1802 4135
rect -1768 4124 -1762 4135
tri -1526 4127 -1501 4152 ne
rect -1501 4127 -1486 4152
tri -1762 4124 -1759 4127 sw
tri -1501 4124 -1498 4127 ne
rect -1498 4124 -1486 4127
tri -1486 4124 -1458 4152 sw
rect -1768 4118 -1759 4124
tri -1759 4118 -1753 4124 sw
tri -1498 4118 -1492 4124 ne
rect -1492 4118 -1458 4124
tri -1458 4118 -1452 4124 sw
rect -1382 4118 -1370 4152
rect -1336 4118 -1288 4152
rect -1254 4118 -1207 4152
rect -1173 4133 -1108 4152
rect -1074 4133 -796 4167
rect -762 4133 -560 4167
rect -1173 4127 -560 4133
rect -508 4127 -496 4179
rect -1173 4121 -444 4127
rect -1173 4118 -453 4121
rect -1768 4106 -1753 4118
tri -1753 4106 -1741 4118 sw
tri -1492 4106 -1480 4118 ne
rect -1480 4112 -1452 4118
tri -1452 4112 -1446 4118 sw
rect -1382 4112 -453 4118
tri -453 4112 -444 4121 nw
rect -416 4174 -370 4186
rect -416 4140 -410 4174
rect -376 4140 -370 4174
rect -1480 4109 -1446 4112
tri -1446 4109 -1443 4112 sw
rect -1480 4106 -1443 4109
tri -1443 4106 -1440 4109 sw
tri -419 4106 -416 4109 se
rect -416 4106 -370 4140
rect -1768 4102 -1741 4106
tri -1741 4102 -1737 4106 sw
rect -1768 4101 -1600 4102
rect -1808 4096 -1600 4101
rect -1808 4062 -1730 4096
rect -1696 4062 -1646 4096
rect -1612 4062 -1600 4096
rect -1808 4060 -1600 4062
rect -1808 4026 -1802 4060
rect -1768 4056 -1600 4060
rect -1572 4100 -1520 4106
tri -1480 4102 -1476 4106 ne
rect -1476 4102 -1440 4106
tri -1440 4102 -1436 4106 sw
tri -423 4102 -419 4106 se
rect -419 4102 -370 4106
rect -1768 4049 -1744 4056
tri -1744 4049 -1737 4056 nw
rect -1768 4026 -1762 4049
tri -1762 4031 -1744 4049 nw
tri -1476 4084 -1458 4102 ne
rect -1458 4084 -1436 4102
tri -1436 4084 -1418 4102 sw
tri -441 4084 -423 4102 se
rect -423 4084 -410 4102
tri -1458 4068 -1442 4084 ne
rect -1442 4068 -410 4084
rect -376 4068 -370 4102
tri -1442 4056 -1430 4068 ne
rect -1430 4056 -370 4068
rect -342 4167 -288 4226
rect -342 4133 -328 4167
rect -294 4133 -288 4167
tri -1520 4049 -1516 4053 sw
rect -1520 4048 -1516 4049
rect -1572 4034 -1516 4048
rect -1808 3985 -1762 4026
rect -1808 3951 -1802 3985
rect -1768 3951 -1762 3985
rect -1520 4028 -1516 4034
tri -1516 4028 -1495 4049 sw
rect -1520 4022 -499 4028
rect -1520 3988 -852 4022
rect -818 3988 -775 4022
rect -741 3988 -698 4022
rect -664 3988 -621 4022
rect -587 3988 -545 4022
rect -511 3988 -499 4022
rect -1520 3982 -499 3988
rect -1572 3976 -499 3982
rect -1808 3948 -1762 3951
tri -1762 3948 -1737 3973 sw
rect -1808 3936 -444 3948
rect -1808 3910 -1677 3936
rect -1808 3876 -1802 3910
rect -1768 3902 -1677 3910
rect -1643 3902 -1221 3936
rect -1187 3902 -444 3936
rect -1768 3882 -444 3902
rect -1768 3876 -1167 3882
rect -1808 3871 -1167 3876
tri -1167 3871 -1156 3882 nw
tri -1018 3871 -1007 3882 ne
rect -1007 3871 -933 3882
tri -933 3871 -922 3882 nw
tri -888 3871 -877 3882 ne
rect -877 3871 -805 3882
tri -805 3871 -794 3882 nw
tri -586 3871 -575 3882 ne
rect -575 3871 -444 3882
rect -1808 3864 -1174 3871
tri -1174 3864 -1167 3871 nw
tri -1007 3864 -1000 3871 ne
rect -1000 3864 -940 3871
tri -940 3864 -933 3871 nw
tri -877 3864 -870 3871 ne
rect -870 3864 -812 3871
tri -812 3864 -805 3871 nw
tri -575 3864 -568 3871 ne
rect -568 3864 -444 3871
rect -1808 3835 -1677 3864
rect -1808 3801 -1802 3835
rect -1768 3830 -1677 3835
rect -1643 3855 -1181 3864
tri -1181 3857 -1174 3864 nw
tri -1000 3857 -993 3864 ne
rect -1643 3830 -1221 3855
rect -1768 3821 -1221 3830
rect -1187 3821 -1181 3855
rect -1768 3801 -1181 3821
rect -1808 3792 -1181 3801
rect -1808 3760 -1677 3792
rect -1808 3726 -1802 3760
rect -1768 3758 -1677 3760
rect -1643 3774 -1181 3792
rect -1643 3758 -1221 3774
rect -1768 3740 -1221 3758
rect -1187 3740 -1181 3774
rect -1768 3726 -1181 3740
rect -1808 3719 -1181 3726
rect -1808 3685 -1677 3719
rect -1643 3693 -1181 3719
rect -1643 3685 -1221 3693
rect -1808 3651 -1802 3685
rect -1768 3673 -1221 3685
rect -1768 3659 -1725 3673
tri -1725 3659 -1711 3673 nw
tri -1344 3659 -1330 3673 ne
rect -1330 3659 -1221 3673
rect -1187 3659 -1181 3693
rect -1768 3651 -1737 3659
rect -1808 3647 -1737 3651
tri -1737 3647 -1725 3659 nw
tri -1330 3647 -1318 3659 ne
rect -1318 3647 -1181 3659
rect -1121 3837 -1025 3849
rect -1121 3803 -1065 3837
rect -1031 3803 -1025 3837
rect -1121 3765 -1025 3803
rect -1121 3731 -1065 3765
rect -1031 3731 -1025 3765
rect -1121 3693 -1025 3731
rect -1121 3659 -1065 3693
rect -1031 3659 -1025 3693
rect -1121 3647 -1025 3659
rect -993 3796 -947 3864
tri -947 3857 -940 3864 nw
tri -870 3857 -863 3864 ne
tri -883 3803 -863 3823 se
rect -863 3803 -819 3864
tri -819 3857 -812 3864 nw
tri -568 3857 -561 3864 ne
tri -887 3799 -883 3803 se
rect -883 3799 -819 3803
tri -888 3798 -887 3799 se
rect -887 3798 -819 3799
rect -992 3794 -948 3795
rect -993 3758 -947 3794
rect -992 3757 -948 3758
rect -993 3744 -947 3756
rect -993 3710 -987 3744
rect -953 3710 -947 3744
rect -993 3672 -947 3710
rect -1808 3638 -1746 3647
tri -1746 3638 -1737 3647 nw
tri -1499 3638 -1492 3645 se
rect -1492 3639 -1440 3645
rect -1808 3624 -1760 3638
tri -1760 3624 -1746 3638 nw
tri -1513 3624 -1499 3638 se
rect -1499 3624 -1492 3638
rect -1808 3610 -1762 3624
tri -1762 3622 -1760 3624 nw
tri -1515 3622 -1513 3624 se
rect -1513 3622 -1492 3624
rect -1808 3576 -1802 3610
rect -1768 3576 -1762 3610
tri -1529 3608 -1515 3622 se
rect -1515 3608 -1492 3622
tri -1530 3607 -1529 3608 se
rect -1529 3607 -1492 3608
tri -1554 3583 -1530 3607 se
rect -1530 3587 -1492 3607
tri -1440 3638 -1433 3645 sw
rect -1121 3638 -1061 3647
tri -1061 3638 -1052 3647 nw
rect -993 3638 -987 3672
rect -953 3638 -947 3672
rect -1440 3608 -1433 3638
tri -1433 3608 -1403 3638 sw
rect -1121 3624 -1075 3638
tri -1075 3624 -1061 3638 nw
rect -993 3626 -947 3638
rect -992 3624 -948 3625
rect -915 3786 -819 3798
rect -915 3752 -909 3786
rect -875 3752 -819 3786
rect -915 3714 -819 3752
rect -915 3680 -909 3714
rect -875 3680 -819 3714
rect -915 3646 -819 3680
rect -759 3837 -713 3849
rect -759 3803 -753 3837
rect -719 3803 -713 3837
rect -759 3765 -713 3803
rect -759 3731 -753 3765
rect -719 3731 -713 3765
rect -759 3693 -713 3731
tri -760 3659 -759 3660 se
rect -759 3659 -753 3693
rect -719 3659 -713 3693
tri -764 3655 -760 3659 se
rect -760 3655 -713 3659
tri -772 3647 -764 3655 se
rect -764 3647 -713 3655
rect -646 3837 -600 3849
rect -646 3803 -640 3837
rect -606 3803 -600 3837
rect -646 3765 -600 3803
rect -646 3731 -640 3765
rect -606 3731 -600 3765
rect -646 3693 -600 3731
rect -646 3659 -640 3693
rect -606 3659 -600 3693
rect -646 3647 -600 3659
rect -915 3645 -820 3646
tri -820 3645 -819 3646 nw
tri -774 3645 -772 3647 se
rect -772 3645 -723 3647
tri -723 3645 -721 3647 nw
rect -645 3645 -601 3646
rect -915 3642 -854 3645
rect -1440 3607 -1403 3608
tri -1403 3607 -1402 3608 sw
rect -1440 3588 -1402 3607
tri -1402 3588 -1383 3607 sw
rect -1440 3587 -1383 3588
rect -1530 3583 -1383 3587
tri -1383 3583 -1378 3588 sw
tri -1126 3583 -1121 3588 se
rect -1121 3583 -1077 3624
tri -1077 3622 -1075 3624 nw
rect -915 3608 -909 3642
rect -875 3611 -854 3642
tri -854 3611 -820 3645 nw
tri -808 3611 -774 3645 se
rect -774 3611 -757 3645
tri -757 3611 -723 3645 nw
rect -875 3609 -856 3611
tri -856 3609 -854 3611 nw
tri -810 3609 -808 3611 se
rect -808 3609 -759 3611
tri -759 3609 -757 3611 nw
rect -646 3609 -600 3645
rect -875 3608 -858 3609
rect -915 3607 -858 3608
tri -858 3607 -856 3609 nw
tri -812 3607 -810 3609 se
rect -810 3607 -761 3609
tri -761 3607 -759 3609 nw
tri -648 3607 -646 3609 se
rect -645 3608 -601 3609
rect -915 3596 -869 3607
tri -869 3596 -858 3607 nw
tri -823 3596 -812 3607 se
rect -812 3596 -772 3607
tri -772 3596 -761 3607 nw
tri -659 3596 -648 3607 se
rect -648 3596 -600 3607
tri -831 3588 -823 3596 se
rect -823 3588 -780 3596
tri -780 3588 -772 3596 nw
tri -667 3588 -659 3596 se
rect -659 3588 -600 3596
tri -1077 3583 -1072 3588 sw
tri -998 3583 -993 3588 se
rect -992 3587 -948 3588
tri -947 3587 -946 3588 sw
tri -832 3587 -831 3588 se
rect -831 3587 -784 3588
rect -947 3586 -946 3587
tri -946 3586 -945 3587 sw
tri -833 3586 -832 3587 se
rect -832 3586 -784 3587
rect -993 3584 -945 3586
tri -945 3584 -943 3586 sw
tri -835 3584 -833 3586 se
rect -833 3584 -784 3586
tri -784 3584 -780 3588 nw
tri -671 3584 -667 3588 se
rect -667 3584 -600 3588
rect -993 3583 -943 3584
tri -943 3583 -942 3584 sw
tri -836 3583 -835 3584 se
rect -835 3583 -785 3584
tri -785 3583 -784 3584 nw
rect -1808 3536 -1762 3576
tri -1564 3573 -1554 3583 se
rect -1554 3575 -1378 3583
rect -1554 3573 -1492 3575
tri -1574 3563 -1564 3573 se
rect -1564 3563 -1492 3573
rect -1808 3502 -1802 3536
rect -1768 3502 -1762 3536
rect -1637 3557 -1492 3563
rect -1440 3573 -1378 3575
tri -1378 3573 -1368 3583 sw
tri -1136 3573 -1126 3583 se
rect -1126 3573 -1072 3583
tri -1072 3573 -1062 3583 sw
tri -1008 3573 -998 3583 se
rect -998 3573 -942 3583
tri -942 3573 -932 3583 sw
tri -846 3573 -836 3583 se
rect -836 3573 -795 3583
tri -795 3573 -785 3583 nw
rect -1440 3563 -1368 3573
tri -1368 3563 -1358 3573 sw
tri -1146 3563 -1136 3573 se
rect -1136 3563 -1062 3573
tri -1062 3563 -1052 3573 sw
tri -1018 3563 -1008 3573 se
rect -1008 3563 -932 3573
tri -932 3563 -922 3573 sw
tri -856 3563 -846 3573 se
rect -846 3563 -805 3573
tri -805 3563 -795 3573 nw
rect -1440 3557 -829 3563
rect -1637 3523 -1625 3557
rect -1591 3523 -1542 3557
rect -1508 3523 -1492 3557
rect -1424 3523 -1374 3557
rect -1340 3523 -1290 3557
rect -1256 3523 -1206 3557
rect -1172 3523 -1122 3557
rect -1088 3539 -829 3557
tri -829 3539 -805 3563 nw
rect -1088 3534 -834 3539
tri -834 3534 -829 3539 nw
rect -1088 3533 -835 3534
tri -835 3533 -834 3534 nw
rect -1088 3532 -836 3533
tri -836 3532 -835 3533 nw
rect -744 3532 -738 3584
rect -686 3532 -674 3584
rect -622 3532 -600 3584
rect -561 3837 -444 3864
rect -561 3803 -484 3837
rect -450 3803 -444 3837
rect -561 3765 -444 3803
rect -561 3731 -484 3765
rect -450 3731 -444 3765
rect -561 3693 -444 3731
rect -561 3659 -484 3693
rect -450 3659 -444 3693
rect -1088 3523 -851 3532
rect -1637 3517 -851 3523
tri -851 3517 -836 3532 nw
rect -1808 3462 -1762 3502
rect -1808 3428 -1802 3462
rect -1768 3428 -1762 3462
rect -1808 3411 -1762 3428
tri -1762 3411 -1760 3413 sw
tri -563 3411 -561 3413 se
rect -561 3411 -444 3659
rect -1808 3395 -1760 3411
tri -1760 3395 -1744 3411 sw
tri -579 3395 -563 3411 se
rect -563 3405 -444 3411
rect -563 3395 -560 3405
rect -1808 3388 -1744 3395
tri -1744 3388 -1737 3395 sw
tri -586 3388 -579 3395 se
rect -579 3388 -560 3395
rect -1808 3354 -1802 3388
rect -1768 3382 -560 3388
rect -1768 3354 -1730 3382
rect -1808 3348 -1730 3354
rect -1696 3348 -1653 3382
rect -1619 3348 -1576 3382
rect -1542 3348 -1499 3382
rect -1465 3348 -1422 3382
rect -1388 3348 -1345 3382
rect -1311 3348 -1268 3382
rect -1234 3348 -1191 3382
rect -1157 3348 -1114 3382
rect -1080 3348 -1037 3382
rect -1003 3348 -960 3382
rect -926 3348 -883 3382
rect -849 3348 -806 3382
rect -772 3348 -729 3382
rect -695 3348 -652 3382
rect -618 3376 -560 3382
rect -618 3348 -580 3376
rect -508 3353 -496 3405
rect -1808 3342 -580 3348
rect -546 3342 -444 3353
tri -611 3323 -592 3342 ne
rect -592 3323 -444 3342
tri -592 3317 -586 3323 ne
rect -586 3315 -444 3323
rect -586 3279 -560 3315
rect -586 3245 -580 3279
rect -508 3263 -496 3315
rect -342 3837 -288 4133
rect -342 3803 -328 3837
rect -294 3803 -288 3837
rect -342 3765 -288 3803
rect -342 3731 -328 3765
rect -294 3731 -288 3765
rect -342 3693 -288 3731
rect -342 3659 -328 3693
rect -294 3659 -288 3693
rect -342 3265 -288 3659
rect -238 4375 -192 4387
rect -238 4359 -232 4375
rect -198 4365 -192 4375
rect -26 4375 20 4387
tri -192 4365 -186 4371 sw
rect -198 4359 -186 4365
rect -238 4302 -186 4307
rect -238 4269 -232 4302
rect -198 4269 -186 4302
rect -238 4195 -232 4217
rect -198 4195 -186 4217
rect -238 4179 -186 4195
rect -238 4122 -232 4127
rect -198 4122 -186 4127
rect -238 4121 -186 4122
rect -238 4083 -192 4121
tri -192 4115 -186 4121 nw
rect -26 4341 -20 4375
rect 14 4341 20 4375
rect -26 4303 20 4341
rect -26 4269 -20 4303
rect 14 4269 20 4303
rect -26 4231 20 4269
rect -26 4197 -20 4231
rect 14 4197 20 4231
rect -26 4159 20 4197
rect -26 4125 -20 4159
rect 14 4125 20 4159
rect -238 4049 -232 4083
rect -198 4049 -192 4083
rect -238 4010 -192 4049
rect -238 3976 -232 4010
rect -198 3976 -192 4010
rect -238 3937 -192 3976
rect -238 3903 -232 3937
rect -198 3903 -192 3937
rect -238 3864 -192 3903
rect -238 3830 -232 3864
rect -198 3830 -192 3864
rect -238 3791 -192 3830
rect -238 3757 -232 3791
rect -198 3757 -192 3791
rect -238 3718 -192 3757
rect -238 3684 -232 3718
rect -198 3684 -192 3718
rect -238 3645 -192 3684
rect -238 3611 -232 3645
rect -198 3611 -192 3645
rect -238 3573 -192 3611
rect -238 3539 -232 3573
rect -198 3539 -192 3573
rect -238 3501 -192 3539
rect -238 3467 -232 3501
rect -198 3467 -192 3501
rect -238 3429 -192 3467
rect -238 3405 -232 3429
rect -198 3411 -192 3429
rect -26 4087 20 4125
rect -26 4053 -20 4087
rect 14 4053 20 4087
rect -26 4015 20 4053
rect -26 3981 -20 4015
rect 14 3981 20 4015
rect -26 3943 20 3981
rect -26 3909 -20 3943
rect 14 3909 20 3943
rect -26 3871 20 3909
rect -26 3837 -20 3871
rect 14 3837 20 3871
rect -26 3799 20 3837
rect -26 3765 -20 3799
rect 14 3765 20 3799
rect -26 3727 20 3765
rect -26 3693 -20 3727
rect 14 3693 20 3727
rect -26 3655 20 3693
rect -26 3621 -20 3655
rect 14 3621 20 3655
rect -26 3583 20 3621
rect -26 3549 -20 3583
rect 14 3549 20 3583
rect -26 3511 20 3549
rect -26 3477 -20 3511
rect 14 3477 20 3511
rect -26 3439 20 3477
tri -192 3411 -186 3417 sw
rect -198 3405 -186 3411
rect -238 3323 -232 3353
rect -198 3323 -186 3353
rect -238 3315 -186 3323
rect -546 3245 -444 3263
rect -586 3237 -444 3245
rect -238 3251 -232 3263
rect -198 3251 -186 3263
tri -444 3237 -443 3238 sw
tri -239 3237 -238 3238 se
rect -238 3237 -186 3251
rect -586 3225 -443 3237
rect -1492 3217 -1440 3223
rect -586 3207 -560 3225
rect -586 3173 -574 3207
rect -508 3173 -496 3225
rect -444 3223 -443 3225
tri -443 3223 -429 3237 sw
tri -253 3223 -239 3237 se
rect -239 3225 -186 3237
rect -239 3223 -238 3225
rect -444 3213 -429 3223
tri -429 3213 -419 3223 sw
tri -263 3213 -253 3223 se
rect -253 3213 -238 3223
rect -444 3207 -238 3213
rect -444 3173 -394 3207
rect -360 3173 -304 3207
rect -270 3173 -238 3207
rect -586 3167 -186 3173
rect -26 3405 -20 3439
rect 14 3405 20 3439
rect -26 3367 20 3405
rect -26 3333 -20 3367
rect 14 3333 20 3367
rect -26 3295 20 3333
rect -26 3261 -20 3295
rect 14 3261 20 3295
rect -26 3223 20 3261
rect -26 3189 -20 3223
rect 14 3189 20 3223
rect -1492 3163 -1440 3165
tri -1440 3163 -1439 3164 sw
rect -1492 3151 -1439 3163
tri -1439 3151 -1427 3163 sw
rect -26 3151 20 3189
rect -1572 3143 -1520 3149
rect -1440 3139 -1427 3151
tri -1427 3139 -1415 3151 sw
rect -1440 3117 -105 3139
tri -105 3117 -83 3139 sw
rect -26 3117 -20 3151
rect 14 3117 20 3151
rect -1440 3099 -83 3117
rect -1492 3093 -83 3099
rect -1572 3079 -1520 3091
tri -125 3089 -121 3093 ne
rect -121 3089 -83 3093
tri -83 3089 -55 3117 sw
tri -121 3088 -120 3089 ne
rect -120 3088 -55 3089
tri -55 3088 -54 3089 sw
tri -120 3081 -113 3088 ne
rect -113 3081 -54 3088
tri -1520 3079 -1518 3081 sw
tri -113 3079 -111 3081 ne
rect -111 3079 -54 3081
rect -1572 3077 -1518 3079
rect -1520 3056 -1518 3077
tri -1518 3056 -1495 3079 sw
tri -111 3073 -105 3079 ne
rect -105 3073 -54 3079
tri -105 3068 -100 3073 ne
rect -1520 3045 -179 3056
tri -179 3045 -168 3056 sw
rect -1520 3025 -168 3045
rect -1572 3015 -168 3025
tri -168 3015 -138 3045 sw
rect -1572 3010 -138 3015
tri -199 3007 -196 3010 ne
rect -196 3007 -138 3010
tri -138 3007 -130 3015 sw
tri -196 3005 -194 3007 ne
rect -194 3005 -130 3007
tri -130 3005 -128 3007 sw
tri -194 2990 -179 3005 ne
rect -179 2990 -128 3005
tri -179 2985 -174 2990 ne
rect -1652 2930 -1646 2982
rect -1594 2930 -1580 2982
rect -1528 2973 -253 2982
tri -253 2973 -244 2982 sw
rect -1528 2941 -244 2973
tri -244 2941 -212 2973 sw
rect -1528 2936 -212 2941
rect -1528 2935 -1517 2936
tri -1517 2935 -1516 2936 nw
tri -273 2935 -272 2936 ne
rect -272 2935 -212 2936
tri -212 2935 -206 2941 sw
rect -1528 2931 -1521 2935
tri -1521 2931 -1517 2935 nw
tri -272 2931 -268 2935 ne
rect -268 2931 -206 2935
tri -206 2931 -202 2935 sw
rect -1528 2930 -1522 2931
tri -1522 2930 -1521 2931 nw
tri -268 2930 -267 2931 ne
rect -267 2930 -202 2931
tri -267 2916 -253 2930 ne
rect -253 2916 -202 2930
tri -253 2911 -248 2916 ne
rect -248 1613 -202 2916
rect -174 1672 -128 2990
rect -100 1756 -54 3073
rect -26 3079 20 3117
rect -26 3045 -20 3079
rect 14 3045 20 3079
rect -26 3007 20 3045
rect -26 2973 -20 3007
rect 14 2973 20 3007
rect -26 2935 20 2973
rect -26 2901 -20 2935
rect 14 2901 20 2935
rect -26 2863 20 2901
rect -26 2829 -20 2863
rect 14 2829 20 2863
rect -26 2791 20 2829
rect -26 2757 -20 2791
rect 14 2757 20 2791
rect -26 2719 20 2757
rect -26 2685 -20 2719
rect 14 2685 20 2719
rect -26 2647 20 2685
rect -26 2613 -20 2647
rect 14 2613 20 2647
rect -26 2575 20 2613
rect -26 2541 -20 2575
rect 14 2541 20 2575
rect -26 2503 20 2541
rect -26 2469 -20 2503
rect 14 2469 20 2503
tri 174 2497 214 2537 se
rect 214 2497 260 4489
tri 260 4473 276 4489 nw
rect 568 4473 623 4489
tri 623 4473 639 4489 nw
tri 888 4473 904 4489 ne
rect 904 4473 950 4489
tri 950 4473 966 4489 sw
rect 568 4461 614 4473
tri 614 4464 623 4473 nw
tri 904 4464 913 4473 ne
rect 913 4467 966 4473
rect 913 4464 914 4467
tri 913 4463 914 4464 ne
rect 820 4455 872 4461
rect 820 4391 872 4403
rect 820 4327 872 4339
rect 820 4263 872 4275
rect 1260 4461 1306 4517
rect 1612 4562 1658 4589
rect 1612 4528 1618 4562
rect 1652 4528 1658 4562
rect 1612 4489 1658 4528
rect 914 4403 966 4415
rect 914 4339 966 4351
rect 914 4275 966 4287
rect 914 4217 966 4223
rect 1612 4455 1618 4489
rect 1652 4455 1658 4489
rect 1612 4416 1658 4455
rect 1612 4382 1618 4416
rect 1652 4382 1658 4416
rect 1612 4343 1658 4382
rect 1612 4309 1618 4343
rect 1652 4309 1658 4343
rect 1612 4270 1658 4309
rect 1612 4236 1618 4270
rect 1652 4236 1658 4270
rect 820 4199 872 4211
rect 820 4135 872 4147
rect 820 4071 872 4083
rect 820 4007 872 4019
rect 820 3943 872 3955
rect 820 3879 872 3891
rect 820 3815 872 3827
rect 820 3751 872 3763
rect 820 3687 872 3699
rect 820 3622 872 3635
rect 820 3557 872 3570
rect 820 3492 872 3505
rect 820 3427 872 3440
rect 820 3362 872 3375
rect 820 3297 872 3310
rect 820 3232 872 3245
rect 820 3167 872 3180
rect 820 3102 872 3115
rect 820 3037 872 3050
rect 820 2972 872 2985
rect 820 2907 872 2920
rect 820 2842 872 2855
rect 820 2777 872 2790
rect 820 2712 872 2725
rect 820 2647 872 2660
rect 820 2582 872 2595
tri 260 2497 300 2537 sw
rect 820 2517 872 2530
rect -26 2431 20 2469
tri 170 2493 174 2497 se
rect 174 2493 300 2497
tri 300 2493 304 2497 sw
rect 170 2487 304 2493
rect 170 2453 182 2487
rect 216 2453 258 2487
rect 292 2453 304 2487
rect 820 2459 872 2465
rect 1612 4197 1658 4236
rect 1612 4163 1618 4197
rect 1652 4163 1658 4197
rect 1612 4124 1658 4163
rect 1612 4090 1618 4124
rect 1652 4090 1658 4124
rect 1612 4051 1658 4090
rect 1612 4017 1618 4051
rect 1652 4017 1658 4051
rect 1612 3977 1658 4017
rect 1612 3943 1618 3977
rect 1652 3943 1658 3977
rect 1612 3903 1658 3943
rect 1612 3869 1618 3903
rect 1652 3869 1658 3903
rect 1612 3829 1658 3869
rect 1612 3795 1618 3829
rect 1652 3795 1658 3829
rect 1612 3755 1658 3795
rect 1612 3721 1618 3755
rect 1652 3721 1658 3755
rect 1612 3681 1658 3721
rect 1612 3647 1618 3681
rect 1652 3647 1658 3681
rect 1612 3607 1658 3647
rect 1612 3573 1618 3607
rect 1652 3573 1658 3607
rect 1612 3533 1658 3573
rect 1612 3499 1618 3533
rect 1652 3499 1658 3533
rect 1612 3459 1658 3499
rect 1612 3425 1618 3459
rect 1652 3425 1658 3459
rect 1612 3385 1658 3425
rect 1612 3351 1618 3385
rect 1652 3351 1658 3385
rect 1612 3311 1658 3351
rect 1612 3277 1618 3311
rect 1652 3277 1658 3311
rect 1612 3237 1658 3277
rect 1612 3203 1618 3237
rect 1652 3203 1658 3237
rect 1612 3163 1658 3203
rect 1612 3129 1618 3163
rect 1652 3129 1658 3163
rect 1612 3089 1658 3129
rect 1612 3055 1618 3089
rect 1652 3055 1658 3089
rect 1612 3015 1658 3055
rect 1612 2981 1618 3015
rect 1652 2981 1658 3015
rect 1612 2941 1658 2981
rect 1612 2907 1618 2941
rect 1652 2907 1658 2941
rect 1612 2867 1658 2907
rect 1612 2833 1618 2867
rect 1652 2833 1658 2867
rect 1612 2793 1658 2833
rect 1612 2759 1618 2793
rect 1652 2759 1658 2793
rect 1612 2719 1658 2759
rect 1612 2685 1618 2719
rect 1652 2685 1658 2719
rect 1612 2645 1658 2685
rect 1612 2611 1618 2645
rect 1652 2611 1658 2645
rect 1612 2571 1658 2611
rect 1612 2537 1618 2571
rect 1652 2537 1658 2571
rect 1612 2497 1658 2537
rect 1612 2463 1618 2497
rect 1652 2463 1658 2497
rect 170 2447 304 2453
rect -26 2397 -20 2431
rect 14 2397 20 2431
tri 547 2423 568 2444 se
rect 568 2423 614 2459
tri 614 2423 639 2448 sw
tri 543 2419 547 2423 se
rect 547 2419 1229 2423
rect -26 2359 20 2397
rect -26 2325 -20 2359
rect 14 2325 20 2359
rect -26 2287 20 2325
rect 90 2413 435 2419
rect 142 2377 435 2413
rect 436 2378 437 2418
rect 473 2378 474 2418
rect 475 2377 1229 2419
rect 142 2361 143 2377
rect 90 2349 143 2361
tri 143 2349 171 2377 nw
tri 1148 2349 1176 2377 ne
rect 1176 2349 1229 2377
rect 90 2347 142 2349
tri 142 2348 143 2349 nw
rect 90 2289 142 2295
rect 186 2343 1133 2349
tri 1176 2348 1177 2349 ne
rect 186 2309 198 2343
rect 232 2309 272 2343
rect 306 2309 346 2343
rect 380 2309 420 2343
rect 454 2309 494 2343
rect 528 2309 568 2343
rect 602 2309 642 2343
rect 676 2312 716 2343
rect 750 2312 790 2343
rect 676 2309 715 2312
rect 767 2309 790 2312
rect 824 2309 864 2343
rect 898 2309 938 2343
rect 972 2309 1012 2343
rect 1046 2309 1087 2343
rect 1121 2309 1133 2343
rect 186 2303 715 2309
rect -26 2253 -20 2287
rect 14 2278 20 2287
rect 186 2286 252 2303
tri 252 2286 269 2303 nw
tri 690 2286 707 2303 ne
rect 707 2286 715 2303
tri 20 2278 28 2286 sw
tri 178 2278 186 2286 se
rect 186 2278 244 2286
tri 244 2278 252 2286 nw
tri 707 2278 715 2286 ne
rect 14 2271 28 2278
tri 28 2271 35 2278 sw
tri 171 2271 178 2278 se
rect 178 2271 237 2278
tri 237 2271 244 2278 nw
rect 767 2303 1133 2309
tri 767 2278 792 2303 nw
rect 14 2261 35 2271
tri 35 2261 45 2271 sw
tri 161 2261 171 2271 se
rect 171 2261 227 2271
tri 227 2261 237 2271 nw
rect 14 2253 203 2261
rect -26 2237 203 2253
tri 203 2237 227 2261 nw
rect 715 2245 721 2260
rect 755 2245 767 2260
rect -26 2231 197 2237
tri 197 2231 203 2237 nw
rect -26 2226 192 2231
tri 192 2226 197 2231 nw
rect -26 2215 181 2226
tri 181 2215 192 2226 nw
rect 245 2220 642 2226
rect -26 2214 44 2215
tri 44 2214 45 2215 nw
rect 245 2214 513 2220
rect -26 2180 -20 2214
rect 14 2180 20 2214
tri 20 2190 44 2214 nw
rect -26 2141 20 2180
rect -26 2107 -20 2141
rect 14 2107 20 2141
rect -26 2068 20 2107
rect -26 2034 -20 2068
rect 14 2034 20 2068
rect -26 1995 20 2034
rect -26 1961 -20 1995
rect 14 1961 20 1995
rect -26 1922 20 1961
rect -26 1888 -20 1922
rect 14 1888 20 1922
rect -26 1849 20 1888
rect -26 1815 -20 1849
rect 14 1815 20 1849
rect -26 1803 20 1815
rect 68 2181 142 2187
rect 68 2175 90 2181
rect 68 2141 74 2175
rect 68 2129 90 2141
rect 68 2114 142 2129
rect 68 2089 90 2114
rect 68 2055 74 2089
rect 108 2055 142 2062
rect 68 2046 142 2055
rect 68 2003 90 2046
rect 68 1969 74 2003
rect 108 1978 142 1994
rect 68 1926 90 1969
rect 68 1917 142 1926
rect 68 1883 74 1917
rect 108 1910 142 1917
rect 68 1858 90 1883
rect 68 1842 142 1858
rect 68 1830 90 1842
rect 68 1796 74 1830
rect 68 1790 90 1796
rect 68 1784 142 1790
rect 245 2180 251 2214
rect 285 2180 513 2214
rect 245 2168 513 2180
rect 565 2168 590 2220
rect 245 2151 642 2168
rect 245 2138 513 2151
rect 245 2104 251 2138
rect 285 2104 513 2138
rect 245 2099 513 2104
rect 565 2099 590 2151
rect 245 2096 642 2099
rect 245 2061 291 2096
tri 291 2071 316 2096 nw
tri 488 2071 513 2096 ne
rect 513 2082 642 2096
rect 245 2027 251 2061
rect 285 2027 291 2061
rect 245 1984 291 2027
rect 245 1950 251 1984
rect 285 1950 291 1984
rect 245 1907 291 1950
rect 245 1873 251 1907
rect 285 1873 291 1907
rect 245 1830 291 1873
rect 245 1796 251 1830
rect 285 1796 291 1830
rect 245 1784 291 1796
rect 439 2035 485 2047
rect 439 2001 445 2035
rect 479 2001 485 2035
rect 439 1951 485 2001
rect 439 1917 445 1951
rect 479 1917 485 1951
rect 439 1867 485 1917
rect 439 1833 445 1867
rect 479 1833 485 1867
rect 439 1783 485 1833
tri -54 1756 -35 1775 sw
rect -100 1755 -35 1756
tri -100 1750 -95 1755 ne
rect -95 1750 -35 1755
tri -35 1750 -29 1756 sw
tri 275 1750 281 1756 se
rect 281 1750 287 1756
tri -95 1749 -94 1750 ne
rect -94 1749 287 1750
tri -94 1737 -82 1749 ne
rect -82 1737 287 1749
tri -82 1714 -59 1737 ne
rect -59 1714 287 1737
tri -59 1709 -54 1714 ne
rect -54 1709 287 1714
tri -54 1707 -52 1709 ne
rect -52 1707 287 1709
tri -52 1704 -49 1707 ne
rect -49 1704 287 1707
rect 339 1704 353 1756
rect 405 1704 411 1756
rect 439 1749 445 1783
rect 479 1749 485 1783
rect 439 1725 485 1749
rect 565 2030 590 2082
rect 513 2013 642 2030
rect 565 1961 590 2013
rect 513 1959 602 1961
rect 636 1959 642 1961
rect 513 1944 642 1959
rect 565 1892 590 1944
rect 513 1885 602 1892
rect 636 1885 642 1892
rect 513 1875 642 1885
rect 565 1823 590 1875
rect 513 1811 602 1823
rect 636 1811 642 1823
rect 513 1805 642 1811
rect 565 1753 590 1805
rect 513 1747 602 1753
tri 513 1737 523 1747 ne
rect 523 1737 602 1747
rect 636 1737 642 1753
tri 523 1728 532 1737 ne
rect 532 1728 642 1737
tri 485 1725 488 1728 sw
tri 532 1725 535 1728 ne
rect 535 1725 642 1728
rect 715 2187 767 2193
rect 715 2179 721 2187
rect 755 2179 767 2187
rect 715 2113 767 2127
rect 914 2269 966 2275
rect 914 2205 966 2217
tri 966 2157 989 2180 sw
tri 1154 2157 1177 2180 se
rect 1177 2175 1229 2349
rect 1496 2246 1542 2459
rect 1612 2423 1658 2463
rect 1612 2389 1618 2423
rect 1652 2389 1658 2423
rect 1612 2349 1658 2389
tri 1658 2349 1683 2374 sw
rect 1612 2315 1618 2349
rect 1652 2343 1895 2349
rect 1652 2315 1709 2343
rect 1612 2309 1709 2315
rect 1743 2309 1895 2343
rect 1612 2305 1895 2309
rect 1612 2303 1855 2305
tri 1824 2278 1849 2303 ne
rect 1849 2271 1855 2303
rect 1889 2271 1895 2305
tri 1496 2241 1501 2246 ne
rect 1501 2241 1542 2246
tri 1542 2241 1567 2266 sw
tri 1501 2231 1511 2241 ne
rect 1511 2231 1756 2241
tri 1756 2231 1766 2241 sw
rect 1849 2231 1895 2271
tri 1511 2200 1542 2231 ne
rect 1542 2200 1766 2231
tri 1542 2197 1545 2200 ne
rect 1545 2197 1766 2200
tri 1766 2197 1800 2231 sw
rect 1849 2197 1855 2231
rect 1889 2197 1895 2231
tri 1545 2195 1547 2197 ne
rect 1547 2195 1800 2197
tri 1736 2190 1741 2195 ne
rect 1741 2190 1800 2195
tri 1800 2190 1807 2197 sw
tri 1741 2180 1751 2190 ne
rect 1751 2180 1807 2190
tri 1229 2175 1234 2180 sw
tri 1751 2175 1756 2180 ne
rect 1756 2175 1807 2180
rect 1177 2170 1234 2175
tri 1234 2170 1239 2175 sw
tri 1756 2170 1761 2175 ne
rect 1177 2157 1239 2170
tri 1239 2157 1252 2170 sw
rect 966 2155 989 2157
tri 989 2155 991 2157 sw
tri 1152 2155 1154 2157 se
rect 1154 2155 1252 2157
tri 1252 2155 1254 2157 sw
rect 966 2153 1708 2155
rect 914 2149 1708 2153
rect 914 2141 980 2149
rect 966 2115 980 2141
rect 1014 2115 1057 2149
rect 1091 2115 1134 2149
rect 1168 2115 1211 2149
rect 1245 2115 1288 2149
rect 1322 2115 1365 2149
rect 1399 2115 1442 2149
rect 1476 2115 1519 2149
rect 1553 2115 1596 2149
rect 1630 2143 1708 2149
rect 1630 2115 1668 2143
rect 966 2109 1668 2115
rect 1702 2109 1708 2143
rect 966 2103 1063 2109
tri 1063 2103 1069 2109 nw
tri 1285 2103 1291 2109 ne
rect 1291 2103 1358 2109
rect 966 2089 1044 2103
rect 914 2083 1044 2089
tri 1044 2084 1063 2103 nw
tri 1291 2084 1310 2103 ne
rect 1310 2086 1358 2103
tri 1358 2086 1381 2109 nw
tri 1637 2086 1660 2109 ne
rect 1660 2086 1708 2109
rect 1356 2085 1357 2086
tri 1357 2085 1358 2086 nw
tri 1660 2085 1661 2086 ne
rect 1661 2085 1708 2086
rect 1311 2084 1355 2085
tri 1356 2084 1357 2085 nw
tri 1661 2084 1662 2085 ne
tri 966 2062 987 2083 ne
rect 987 2062 1044 2083
rect 715 2047 767 2061
tri 987 2053 996 2062 ne
rect 996 2053 1044 2062
tri 996 2051 998 2053 ne
rect 998 2051 1044 2053
rect 715 1986 721 1995
rect 755 1986 767 1995
rect 715 1981 767 1986
rect 715 1915 721 1929
rect 755 1915 767 1929
rect 715 1854 767 1863
rect 715 1849 721 1854
rect 755 1849 767 1854
rect 715 1783 767 1797
rect 715 1725 767 1731
rect 999 2049 1043 2050
rect 998 2013 1044 2049
rect 999 2012 1043 2013
rect 998 1999 1044 2011
rect 998 1965 1004 1999
rect 1038 1965 1044 1999
rect 998 1926 1044 1965
rect 998 1892 1004 1926
rect 1038 1892 1044 1926
rect 998 1853 1044 1892
rect 998 1819 1004 1853
rect 1038 1819 1044 1853
rect 998 1780 1044 1819
rect 998 1746 1004 1780
rect 1038 1746 1044 1780
rect 439 1716 488 1725
tri 488 1716 497 1725 sw
rect 439 1714 497 1716
tri 497 1714 499 1716 sw
rect 439 1707 499 1714
tri 499 1707 506 1714 sw
rect 998 1707 1044 1746
rect 439 1699 506 1707
tri -174 1667 -169 1672 ne
rect -169 1667 -128 1672
tri -128 1667 -103 1692 sw
tri -169 1665 -167 1667 ne
rect -167 1665 405 1667
tri -167 1638 -140 1665 ne
rect -140 1661 405 1665
rect -140 1638 353 1661
tri -140 1634 -136 1638 ne
rect -136 1634 353 1638
tri -136 1626 -128 1634 ne
rect -128 1626 353 1634
tri -128 1621 -123 1626 ne
rect -123 1621 353 1626
tri 328 1618 331 1621 ne
rect 331 1618 353 1621
tri -202 1613 -197 1618 sw
tri 331 1613 336 1618 ne
rect 336 1613 353 1618
rect -248 1598 -197 1613
tri -248 1593 -243 1598 ne
rect -243 1596 -197 1598
tri -197 1596 -180 1613 sw
tri 336 1596 353 1613 ne
rect 439 1665 445 1699
rect 479 1697 506 1699
tri 506 1697 516 1707 sw
rect 479 1691 826 1697
tri 826 1691 832 1697 sw
rect 479 1673 832 1691
tri 832 1673 850 1691 sw
rect 998 1673 1004 1707
rect 1038 1673 1044 1707
rect 479 1672 850 1673
tri 850 1672 851 1673 sw
rect 479 1665 851 1672
rect 439 1658 851 1665
tri 851 1658 865 1672 sw
rect 439 1653 865 1658
tri 804 1638 819 1653 ne
rect 819 1638 865 1653
tri 819 1637 820 1638 ne
rect 820 1637 865 1638
tri 820 1634 823 1637 ne
rect 823 1634 865 1637
tri 823 1628 829 1634 ne
rect 715 1619 767 1625
tri 405 1613 410 1618 sw
rect 405 1609 410 1613
rect -243 1593 -180 1596
tri -180 1593 -177 1596 sw
rect 353 1595 410 1609
tri -243 1587 -237 1593 ne
rect -237 1587 190 1593
tri -237 1553 -203 1587 ne
rect -203 1553 120 1587
rect 154 1553 190 1587
tri -203 1552 -202 1553 ne
rect -202 1552 190 1553
tri -202 1547 -197 1552 ne
rect -197 1547 190 1552
tri 178 1541 184 1547 ne
rect 184 1541 190 1547
rect 242 1541 256 1593
rect 308 1541 314 1593
rect 405 1593 410 1595
tri 410 1593 430 1613 sw
rect 405 1587 594 1593
rect 426 1553 470 1587
rect 504 1553 548 1587
rect 582 1553 594 1587
rect 405 1547 594 1553
rect 715 1553 767 1567
rect 353 1537 405 1543
tri 405 1537 415 1547 nw
rect 715 1487 767 1501
rect 829 1492 865 1634
rect 998 1634 1044 1673
rect 998 1600 1004 1634
rect 1038 1600 1044 1634
rect 998 1561 1044 1600
rect 998 1527 1004 1561
rect 1038 1527 1044 1561
rect 998 1515 1044 1527
rect 1154 2053 1200 2065
rect 1154 2019 1160 2053
rect 1194 2019 1200 2053
rect 1154 1976 1200 2019
rect 1154 1942 1160 1976
rect 1194 1942 1200 1976
rect 1154 1900 1200 1942
rect 1154 1866 1160 1900
rect 1194 1866 1200 1900
rect 1154 1824 1200 1866
rect 1154 1790 1160 1824
rect 1194 1797 1200 1824
rect 1310 2048 1356 2084
rect 1311 2047 1355 2048
rect 1310 2034 1356 2046
rect 1310 2000 1316 2034
rect 1350 2000 1356 2034
rect 1310 1955 1356 2000
rect 1310 1921 1316 1955
rect 1350 1921 1356 1955
rect 1310 1876 1356 1921
rect 1310 1842 1316 1876
rect 1350 1842 1356 1876
tri 1200 1797 1202 1799 sw
tri 1308 1797 1310 1799 se
rect 1310 1797 1356 1842
rect 1194 1790 1202 1797
rect 1154 1763 1202 1790
tri 1202 1763 1236 1797 sw
tri 1274 1763 1308 1797 se
rect 1308 1763 1316 1797
rect 1350 1763 1356 1797
rect 1154 1762 1236 1763
tri 1236 1762 1237 1763 sw
rect 1154 1748 1235 1762
rect 1154 1714 1160 1748
rect 1194 1716 1235 1748
rect 1236 1717 1237 1761
rect 1194 1714 1218 1716
rect 1154 1697 1218 1714
tri 1218 1697 1237 1716 nw
tri 1273 1762 1274 1763 se
rect 1274 1762 1356 1763
rect 1273 1717 1274 1761
rect 1275 1718 1356 1762
rect 1275 1716 1316 1718
tri 1273 1697 1292 1716 ne
rect 1292 1697 1316 1716
rect 1154 1691 1212 1697
tri 1212 1691 1218 1697 nw
tri 1292 1691 1298 1697 ne
rect 1298 1691 1316 1697
rect 1154 1684 1205 1691
tri 1205 1684 1212 1691 nw
tri 1298 1684 1305 1691 ne
rect 1305 1684 1316 1691
rect 1350 1684 1356 1718
rect 1154 1672 1200 1684
tri 1200 1679 1205 1684 nw
tri 1305 1679 1310 1684 ne
rect 1154 1638 1160 1672
rect 1194 1638 1200 1672
rect 1154 1596 1200 1638
rect 1154 1562 1160 1596
rect 1194 1562 1200 1596
rect 1154 1550 1200 1562
rect 1155 1548 1199 1549
rect 1154 1512 1200 1548
rect 1310 1639 1356 1684
rect 1310 1605 1316 1639
rect 1350 1605 1356 1639
rect 1566 2053 1612 2065
rect 1566 2019 1572 2053
rect 1606 2019 1612 2053
rect 1566 1979 1612 2019
rect 1566 1945 1572 1979
rect 1606 1945 1612 1979
rect 1566 1905 1612 1945
rect 1566 1871 1572 1905
rect 1606 1871 1612 1905
rect 1566 1831 1612 1871
rect 1566 1797 1572 1831
rect 1606 1797 1612 1831
rect 1566 1758 1612 1797
rect 1566 1724 1572 1758
rect 1606 1724 1612 1758
rect 1566 1685 1612 1724
rect 1566 1651 1572 1685
rect 1606 1651 1612 1685
rect 1566 1639 1612 1651
rect 1567 1637 1611 1638
rect 1662 2062 1708 2085
rect 1662 2028 1668 2062
rect 1702 2028 1708 2062
rect 1662 1981 1708 2028
rect 1662 1947 1668 1981
rect 1702 1947 1708 1981
rect 1662 1900 1708 1947
rect 1662 1866 1668 1900
rect 1702 1866 1708 1900
rect 1662 1820 1708 1866
rect 1662 1786 1668 1820
rect 1702 1786 1708 1820
rect 1662 1740 1708 1786
rect 1662 1706 1668 1740
rect 1702 1706 1708 1740
rect 1662 1660 1708 1706
rect 1310 1561 1356 1605
rect 1662 1626 1668 1660
rect 1702 1626 1708 1660
tri 1545 1580 1566 1601 se
rect 1567 1600 1611 1601
rect 1566 1580 1612 1599
rect 1310 1527 1316 1561
rect 1350 1527 1356 1561
tri 1512 1547 1545 1580 se
rect 1545 1547 1612 1580
rect 1662 1580 1708 1626
tri 1511 1546 1512 1547 se
rect 1512 1546 1573 1547
tri 1573 1546 1574 1547 nw
rect 1662 1546 1668 1580
rect 1702 1546 1708 1580
tri 1504 1539 1511 1546 se
rect 1511 1539 1566 1546
tri 1566 1539 1573 1546 nw
tri 1496 1531 1504 1539 se
rect 1504 1531 1558 1539
tri 1558 1531 1566 1539 nw
rect 1662 1534 1708 1546
rect 1310 1515 1356 1527
tri 1480 1515 1496 1531 se
rect 1496 1515 1518 1531
tri 1477 1512 1480 1515 se
rect 1480 1512 1518 1515
tri 829 1491 830 1492 ne
rect 830 1491 865 1492
tri 865 1491 886 1512 sw
tri 1133 1491 1154 1512 se
rect 1155 1511 1199 1512
tri 1200 1511 1201 1512 sw
tri 1476 1511 1477 1512 se
rect 1477 1511 1518 1512
rect 1200 1510 1201 1511
tri 1201 1510 1202 1511 sw
tri 1475 1510 1476 1511 se
rect 1476 1510 1518 1511
rect 1154 1491 1202 1510
tri 1202 1491 1221 1510 sw
tri 1456 1491 1475 1510 se
rect 1475 1491 1518 1510
tri 1518 1491 1558 1531 nw
tri 830 1487 834 1491 ne
rect 834 1487 886 1491
tri 886 1487 890 1491 sw
tri 1129 1487 1133 1491 se
rect 1133 1487 1221 1491
tri 1221 1487 1225 1491 sw
tri 1452 1487 1456 1491 se
rect 1456 1487 1514 1491
tri 1514 1487 1518 1491 nw
rect -115 1439 78 1485
rect 80 1484 116 1485
rect 79 1440 117 1484
rect 118 1479 339 1485
rect 118 1445 157 1479
rect 191 1445 289 1479
rect 323 1445 339 1479
rect 80 1439 116 1440
rect 118 1439 339 1445
rect 340 1440 341 1484
rect 377 1440 378 1484
rect 379 1479 533 1485
rect 535 1484 571 1485
rect 379 1445 403 1479
rect 437 1445 487 1479
rect 521 1445 533 1479
rect 379 1439 533 1445
rect 534 1440 572 1484
rect 535 1439 571 1440
rect 573 1439 667 1485
rect -115 1423 -54 1439
tri -54 1423 -38 1439 nw
tri 596 1423 612 1439 ne
rect 612 1423 667 1439
rect -115 1417 -60 1423
tri -60 1417 -54 1423 nw
tri 612 1417 618 1423 ne
rect 618 1417 667 1423
rect -115 -100 -63 1417
tri -63 1414 -60 1417 nw
tri 618 1414 621 1417 ne
rect -26 1393 20 1405
rect -26 1359 -20 1393
rect 14 1359 20 1393
rect -26 1321 20 1359
tri 596 1355 621 1380 se
rect 621 1355 667 1417
rect -26 1287 -20 1321
rect 14 1287 20 1321
rect -26 1249 20 1287
rect -26 1215 -20 1249
rect 14 1215 20 1249
rect -26 1177 20 1215
rect -26 1143 -20 1177
rect 14 1143 20 1177
rect -26 1105 20 1143
rect -26 1071 -20 1105
rect 14 1071 20 1105
rect -26 1033 20 1071
rect -26 999 -20 1033
rect 14 999 20 1033
rect -26 961 20 999
rect -26 927 -20 961
rect 14 927 20 961
rect -26 889 20 927
rect -26 855 -20 889
rect 14 855 20 889
rect -26 817 20 855
rect -26 783 -20 817
rect 14 783 20 817
rect -26 745 20 783
rect 84 1349 667 1355
rect 84 1343 513 1349
rect 84 1309 90 1343
rect 124 1309 513 1343
rect 84 1297 513 1309
rect 565 1343 667 1349
rect 565 1309 602 1343
rect 636 1309 667 1343
rect 565 1297 667 1309
rect 84 1272 667 1297
rect 84 1270 513 1272
rect 84 1236 90 1270
rect 124 1236 513 1270
rect 84 1225 513 1236
rect 84 1197 130 1225
tri 130 1200 155 1225 nw
tri 488 1200 513 1225 ne
rect 565 1271 667 1272
rect 565 1237 602 1271
rect 636 1237 667 1271
rect 565 1220 667 1237
rect 84 1163 90 1197
rect 124 1163 130 1197
rect 513 1199 667 1220
rect 513 1195 602 1199
rect 84 1123 130 1163
rect 84 1089 90 1123
rect 124 1089 130 1123
rect 84 1049 130 1089
rect 84 1015 90 1049
rect 124 1015 130 1049
rect 84 975 130 1015
rect 84 941 90 975
rect 124 941 130 975
rect 84 901 130 941
rect 84 867 90 901
rect 124 867 130 901
rect 84 827 130 867
rect 84 793 90 827
rect 124 793 130 827
rect 340 1171 485 1177
rect 340 1165 433 1171
rect 340 1131 346 1165
rect 380 1131 433 1165
rect 340 1119 433 1131
rect 340 1107 485 1119
rect 340 1086 433 1107
rect 340 1052 346 1086
rect 380 1055 433 1086
rect 380 1052 485 1055
rect 340 1049 485 1052
rect 565 1165 602 1195
rect 636 1165 667 1199
rect 565 1143 667 1165
rect 513 1127 667 1143
rect 513 1118 602 1127
rect 565 1093 602 1118
rect 636 1093 667 1127
rect 565 1066 667 1093
rect 513 1055 667 1066
rect 340 1036 452 1049
tri 452 1036 465 1049 nw
rect 513 1041 602 1055
rect 340 1021 437 1036
tri 437 1021 452 1036 nw
tri 498 1021 513 1036 se
rect 340 1017 433 1021
tri 433 1017 437 1021 nw
tri 494 1017 498 1021 se
rect 498 1017 513 1021
rect 340 1008 424 1017
tri 424 1008 433 1017 nw
tri 485 1008 494 1017 se
rect 494 1008 513 1017
rect 340 1006 411 1008
rect 340 972 346 1006
rect 380 995 411 1006
tri 411 995 424 1008 nw
tri 472 995 485 1008 se
rect 485 995 513 1008
rect 380 983 399 995
tri 399 983 411 995 nw
tri 460 983 472 995 se
rect 472 989 513 995
rect 565 1021 602 1041
rect 636 1021 667 1055
rect 565 989 667 1021
rect 472 983 667 989
rect 380 972 386 983
rect 340 926 386 972
tri 386 970 399 983 nw
tri 447 970 460 983 se
rect 460 970 602 983
rect 340 892 346 926
rect 380 892 386 926
rect 340 846 386 892
rect 340 812 346 846
rect 380 812 386 846
rect 340 800 386 812
tri 439 962 447 970 se
rect 447 962 602 970
rect 439 956 602 962
rect 491 949 602 956
rect 636 949 667 983
rect 491 911 667 949
rect 491 904 602 911
rect 439 881 602 904
rect 491 877 602 881
rect 636 877 667 911
rect 491 839 667 877
rect 491 829 602 839
rect 439 805 602 829
rect 636 805 667 839
rect 84 781 130 793
rect 491 753 667 805
rect 439 747 667 753
tri 834 1458 863 1487 ne
rect 863 1458 1485 1487
tri 1485 1458 1514 1487 nw
tri 863 1457 864 1458 ne
rect 864 1457 1484 1458
tri 1484 1457 1485 1458 nw
tri 864 1456 865 1457 ne
rect 865 1456 1483 1457
tri 1483 1456 1484 1457 nw
tri 865 1443 878 1456 ne
rect 878 1443 1470 1456
tri 1470 1443 1483 1456 nw
rect 715 1423 721 1435
rect 755 1423 767 1435
rect 715 1421 767 1423
rect 1076 1409 1625 1415
rect 1076 1375 1088 1409
rect 1122 1375 1170 1409
rect 1204 1375 1252 1409
rect 1286 1375 1334 1409
rect 1368 1375 1416 1409
rect 1450 1375 1498 1409
rect 1532 1375 1573 1409
rect 1076 1369 1573 1375
rect 715 1355 721 1369
rect 755 1355 767 1369
tri 1548 1344 1573 1369 ne
rect 1573 1345 1625 1357
rect 715 1289 721 1303
rect 755 1289 767 1303
tri 767 1270 786 1289 sw
rect 1573 1287 1625 1293
rect 767 1237 786 1270
rect 715 1236 786 1237
tri 786 1236 820 1270 sw
rect 715 1228 820 1236
tri 820 1228 828 1236 sw
rect 715 1226 783 1228
rect 715 1223 721 1226
rect 755 1223 783 1226
rect 767 1171 783 1223
rect 715 1157 783 1171
rect 767 1105 783 1157
rect 715 1091 783 1105
rect 767 1039 783 1091
rect 715 1038 721 1039
rect 755 1038 783 1039
rect 715 1025 807 1038
rect 767 1017 807 1025
tri 807 1017 828 1038 nw
rect 767 978 768 1017
tri 768 978 807 1017 nw
tri 767 977 768 978 nw
rect 715 961 721 973
rect 755 961 767 973
rect 715 959 767 961
rect 1573 973 1625 979
rect 715 894 721 907
rect 755 894 767 907
tri 1556 905 1573 922 se
rect 1573 909 1625 921
tri 1548 897 1556 905 se
rect 1556 897 1573 905
rect 1076 891 1573 897
rect 1076 857 1088 891
rect 1122 857 1170 891
rect 1204 857 1252 891
rect 1286 857 1334 891
rect 1368 857 1416 891
rect 1450 857 1498 891
rect 1532 857 1573 891
rect 1076 851 1625 857
rect 715 841 767 842
rect 715 829 721 841
rect 755 829 767 841
tri 863 808 878 823 se
rect 878 808 1470 823
tri 1470 808 1485 823 sw
tri 853 798 863 808 se
rect 863 806 1485 808
tri 1485 806 1487 808 sw
rect 863 798 1487 806
tri 1487 798 1495 806 sw
tri 1753 798 1761 806 se
rect 1761 798 1807 2175
rect 715 764 767 777
rect -26 711 -20 745
rect 14 711 20 745
rect -26 673 20 711
rect 105 713 325 719
rect 105 679 117 713
rect 151 679 202 713
rect 236 679 273 713
rect 105 673 273 679
rect -26 639 -20 673
rect 14 639 20 673
tri 248 653 268 673 ne
rect 268 661 273 673
rect 268 653 325 661
tri 268 648 273 653 ne
rect -26 601 20 639
rect -26 567 -20 601
rect 14 567 20 601
rect 273 647 325 653
rect 273 589 325 595
rect 353 713 591 719
rect 423 679 467 713
rect 501 679 545 713
rect 579 679 591 713
rect 405 673 591 679
rect 715 699 767 712
rect 405 661 410 673
rect 353 653 410 661
tri 410 653 430 673 nw
rect 353 647 405 653
tri 405 648 410 653 nw
rect 715 641 767 647
tri 829 774 853 798 se
rect 853 781 1495 798
tri 1495 781 1512 798 sw
tri 1736 781 1753 798 se
rect 1753 781 1807 798
rect 853 779 1512 781
rect 853 774 885 779
tri 885 774 890 779 nw
tri 1129 774 1134 779 ne
rect 1134 774 1205 779
rect 829 759 870 774
tri 870 759 885 774 nw
tri 1134 759 1149 774 ne
rect 1149 759 1205 774
tri 1205 759 1225 779 nw
tri 1452 759 1472 779 ne
rect 1472 759 1512 779
tri 1512 759 1534 781 sw
tri 1714 759 1736 781 se
rect 1736 759 1807 781
tri 824 633 829 638 se
rect 829 633 865 759
tri 865 754 870 759 nw
tri 1149 754 1154 759 ne
rect 1154 756 1202 759
tri 1202 756 1205 759 nw
tri 1472 756 1475 759 ne
rect 1475 756 1534 759
rect 1200 755 1201 756
tri 1201 755 1202 756 nw
tri 1475 755 1476 756 ne
rect 1476 755 1534 756
rect 1155 754 1199 755
tri 1200 754 1201 755 nw
tri 1476 754 1477 755 ne
rect 1477 754 1534 755
tri 823 632 824 633 se
rect 824 632 865 633
tri 820 629 823 632 se
rect 823 629 865 632
tri 819 628 820 629 se
rect 820 628 865 629
tri 804 613 819 628 se
rect 819 613 865 628
rect 353 589 405 595
rect 354 587 404 588
rect 433 608 865 613
rect 433 601 852 608
rect -26 529 20 567
rect -26 495 -20 529
rect 14 495 20 529
rect -26 457 20 495
rect -26 423 -20 457
rect 14 423 20 457
rect -26 384 20 423
rect -26 350 -20 384
rect 14 350 20 384
rect -26 311 20 350
rect -26 277 -20 311
rect 14 277 20 311
rect -26 238 20 277
rect -26 204 -20 238
rect 14 204 20 238
rect -26 165 20 204
rect -26 131 -20 165
rect 14 131 20 165
rect -26 92 20 131
rect -26 58 -20 92
rect 14 58 20 92
rect -26 46 20 58
rect 68 574 142 580
rect 68 568 90 574
rect 68 534 74 568
rect 433 567 439 601
rect 473 595 852 601
tri 852 595 865 608 nw
rect 902 739 948 751
rect 902 705 908 739
rect 942 705 948 739
rect 902 667 948 705
rect 902 633 908 667
rect 942 633 948 667
rect 902 595 948 633
rect 473 587 844 595
tri 844 587 852 595 nw
rect 473 575 832 587
tri 832 575 844 587 nw
rect 473 569 826 575
tri 826 569 832 575 nw
rect 473 567 496 569
rect 433 561 496 567
tri 496 561 504 569 nw
rect 902 561 908 595
rect 942 561 948 595
rect 433 559 494 561
tri 494 559 496 561 nw
rect 433 552 487 559
tri 487 552 494 559 nw
rect 433 551 486 552
tri 486 551 487 552 nw
rect 68 522 90 534
tri 331 529 353 551 se
rect 354 550 404 551
rect 353 529 405 549
tri 330 528 331 529 se
rect 331 528 405 529
rect 68 504 142 522
tri 315 513 330 528 se
rect 330 513 405 528
rect 68 487 90 504
rect 68 453 74 487
rect 68 452 90 453
rect 68 434 142 452
rect 68 406 90 434
rect 68 372 74 406
rect 108 372 142 382
rect 68 326 142 372
rect 68 292 74 326
rect 108 292 142 326
rect 68 246 142 292
rect 68 212 74 246
rect 108 212 142 246
rect 68 166 142 212
rect 68 132 74 166
rect 108 132 142 166
rect 244 501 405 513
rect 244 467 250 501
rect 284 497 405 501
rect 433 550 485 551
tri 485 550 486 551 nw
rect 433 528 479 550
tri 479 544 485 550 nw
rect 284 494 350 497
tri 350 494 353 497 nw
rect 433 494 439 528
rect 473 494 479 528
rect 284 488 344 494
tri 344 488 350 494 nw
rect 284 486 342 488
tri 342 486 344 488 nw
rect 284 476 332 486
tri 332 476 342 486 nw
rect 284 467 321 476
rect 244 411 321 467
tri 321 465 332 476 nw
rect 244 377 250 411
rect 284 377 321 411
rect 244 329 321 377
rect 433 456 479 494
rect 433 422 439 456
rect 473 422 479 456
rect 433 384 479 422
rect 433 350 439 384
rect 473 350 479 384
rect 433 338 479 350
rect 596 529 642 541
rect 596 495 602 529
rect 636 495 642 529
rect 596 453 642 495
rect 596 419 602 453
rect 636 419 642 453
rect 596 377 642 419
rect 596 343 602 377
rect 636 343 642 377
tri 321 329 322 330 sw
tri 595 329 596 330 se
rect 596 329 642 343
rect 244 324 322 329
tri 322 324 327 329 sw
tri 590 324 595 329 se
rect 595 324 642 329
rect 244 321 327 324
rect 244 287 250 321
rect 284 305 327 321
tri 327 305 346 324 sw
tri 571 305 590 324 se
rect 590 305 642 324
rect 284 302 642 305
rect 284 299 602 302
rect 284 287 449 299
rect 244 247 449 287
rect 501 247 513 299
rect 565 268 602 299
rect 636 268 642 302
rect 565 247 642 268
rect 244 232 642 247
rect 244 231 449 232
rect 244 197 250 231
rect 284 197 449 231
rect 244 180 449 197
rect 501 180 513 232
rect 565 227 642 232
rect 565 193 602 227
rect 636 193 642 227
rect 565 180 642 193
rect 244 164 642 180
rect 244 137 449 164
rect 68 86 142 132
tri 399 118 418 137 ne
rect 418 118 449 137
tri 418 117 419 118 ne
rect 419 117 449 118
tri 419 114 422 117 ne
rect 422 114 449 117
tri 422 106 430 114 ne
rect 430 112 449 114
rect 501 112 513 164
rect 565 152 642 164
rect 565 118 602 152
rect 636 118 642 152
rect 565 112 642 118
rect 430 106 642 112
rect 715 535 767 541
rect 715 465 767 483
rect 715 412 721 413
rect 755 412 767 413
rect 715 395 767 412
rect 715 329 721 343
rect 755 329 767 343
rect 715 325 767 329
rect 715 255 721 273
rect 755 255 767 273
rect 715 197 767 203
rect 715 185 721 197
rect 755 185 767 197
rect 715 114 767 133
rect 68 52 74 86
rect 108 52 142 86
rect 68 40 142 52
rect 273 79 325 85
rect 273 13 325 27
rect 273 -45 325 -39
rect 274 -47 324 -46
rect 273 -83 325 -47
tri 256 -100 273 -83 se
rect 274 -84 324 -83
rect 273 -100 325 -85
tri 248 -108 256 -100 se
rect 256 -108 325 -100
rect 248 -137 325 -108
rect 353 79 405 85
rect 353 13 405 27
rect 902 522 948 561
rect 902 488 908 522
rect 942 488 948 522
rect 902 449 948 488
rect 902 415 908 449
rect 942 415 948 449
rect 902 376 948 415
rect 902 342 908 376
rect 942 342 948 376
rect 902 303 948 342
rect 902 269 908 303
rect 942 269 948 303
rect 902 230 948 269
rect 998 739 1044 751
rect 998 705 1004 739
rect 1038 705 1044 739
rect 998 666 1044 705
rect 998 632 1004 666
rect 1038 632 1044 666
rect 998 593 1044 632
rect 998 559 1004 593
rect 1038 559 1044 593
rect 998 520 1044 559
rect 998 486 1004 520
rect 1038 486 1044 520
rect 998 446 1044 486
rect 998 412 1004 446
rect 1038 412 1044 446
rect 998 372 1044 412
rect 998 338 1004 372
rect 1038 338 1044 372
rect 998 298 1044 338
rect 1154 718 1200 754
tri 1477 751 1480 754 ne
rect 1480 751 1534 754
rect 1155 717 1199 718
rect 1154 704 1200 716
rect 1154 670 1160 704
rect 1194 670 1200 704
rect 1154 628 1200 670
rect 1154 594 1160 628
rect 1194 594 1200 628
rect 1154 582 1200 594
rect 1310 739 1356 751
rect 1310 705 1316 739
rect 1350 705 1356 739
tri 1480 725 1506 751 ne
rect 1506 732 1534 751
tri 1534 732 1561 759 sw
tri 1687 732 1714 759 se
rect 1714 732 1807 759
rect 1506 725 1561 732
tri 1561 725 1568 732 sw
tri 1506 720 1511 725 ne
rect 1511 720 1568 725
tri 1568 720 1573 725 sw
rect 1662 720 1807 732
tri 1511 719 1512 720 ne
rect 1512 719 1573 720
tri 1573 719 1574 720 sw
rect 1310 661 1356 705
tri 1512 686 1545 719 ne
rect 1545 686 1612 719
tri 1545 665 1566 686 ne
rect 1566 667 1612 686
rect 1567 665 1611 666
rect 1662 686 1668 720
rect 1702 686 1807 720
rect 1310 627 1316 661
rect 1350 627 1356 661
rect 1662 640 1807 686
tri 1200 582 1205 587 sw
tri 1305 582 1310 587 se
rect 1310 582 1356 627
rect 1154 575 1205 582
tri 1205 575 1212 582 sw
tri 1298 575 1305 582 se
rect 1305 575 1316 582
rect 1154 569 1212 575
tri 1212 569 1218 575 sw
tri 1292 569 1298 575 se
rect 1298 569 1316 575
rect 1154 552 1218 569
rect 1154 518 1160 552
rect 1194 551 1218 552
tri 1218 551 1236 569 sw
tri 1274 551 1292 569 se
rect 1292 551 1316 569
rect 1194 550 1236 551
tri 1236 550 1237 551 sw
rect 1194 518 1235 550
rect 1154 504 1235 518
rect 1236 505 1237 549
rect 1154 503 1236 504
tri 1236 503 1237 504 nw
tri 1273 550 1274 551 se
rect 1274 550 1316 551
rect 1273 505 1274 549
rect 1275 548 1316 550
rect 1350 548 1356 582
rect 1275 504 1356 548
tri 1273 503 1274 504 ne
rect 1274 503 1356 504
rect 1154 476 1202 503
rect 1154 442 1160 476
rect 1194 469 1202 476
tri 1202 469 1236 503 nw
tri 1274 469 1308 503 ne
rect 1308 469 1316 503
rect 1350 469 1356 503
rect 1194 442 1200 469
tri 1200 467 1202 469 nw
tri 1308 467 1310 469 ne
rect 1154 400 1200 442
rect 1154 366 1160 400
rect 1194 366 1200 400
rect 1154 324 1200 366
rect 998 264 1004 298
rect 1038 290 1044 298
tri 1044 290 1060 306 sw
rect 1154 290 1160 324
rect 1194 290 1200 324
rect 1038 287 1060 290
tri 1060 287 1063 290 sw
rect 1038 285 1063 287
tri 1063 285 1065 287 sw
rect 1038 272 1065 285
tri 1065 272 1078 285 sw
rect 1038 264 1078 272
rect 998 252 1078 264
tri 998 247 1003 252 ne
rect 1003 247 1078 252
rect 902 196 908 230
rect 942 196 948 230
tri 1003 218 1032 247 ne
rect 1032 220 1078 247
rect 1033 218 1077 219
rect 902 175 948 196
rect 1032 182 1078 218
rect 1154 247 1200 290
rect 1154 213 1160 247
rect 1194 213 1200 247
rect 1154 201 1200 213
rect 1310 424 1356 469
rect 1310 390 1316 424
rect 1350 390 1356 424
rect 1310 345 1356 390
rect 1310 311 1316 345
rect 1350 311 1356 345
rect 1310 266 1356 311
rect 1310 232 1316 266
rect 1350 232 1356 266
rect 1310 220 1356 232
rect 1311 218 1355 219
rect 1310 182 1356 218
rect 1567 628 1611 629
rect 1566 615 1612 627
rect 1566 581 1572 615
rect 1606 581 1612 615
rect 1566 542 1612 581
rect 1566 508 1572 542
rect 1606 508 1612 542
rect 1566 469 1612 508
rect 1566 435 1572 469
rect 1606 435 1612 469
rect 1566 395 1612 435
rect 1566 361 1572 395
rect 1606 361 1612 395
rect 1566 321 1612 361
rect 1566 287 1572 321
rect 1606 287 1612 321
rect 1566 247 1612 287
rect 1566 213 1572 247
rect 1606 213 1612 247
rect 1566 201 1612 213
rect 1662 606 1668 640
rect 1702 606 1807 640
rect 1662 560 1807 606
rect 1662 526 1668 560
rect 1702 526 1807 560
rect 1662 480 1807 526
rect 1662 446 1668 480
rect 1702 446 1807 480
rect 1662 400 1807 446
rect 1662 366 1668 400
rect 1702 366 1807 400
rect 1662 319 1807 366
rect 1662 285 1668 319
rect 1702 285 1807 319
rect 1662 238 1807 285
rect 1662 204 1668 238
rect 1702 204 1807 238
tri 948 175 955 182 sw
tri 1025 175 1032 182 se
rect 1033 181 1077 182
tri 1078 181 1079 182 sw
tri 1309 181 1310 182 se
rect 1311 181 1355 182
tri 1356 181 1357 182 sw
tri 1661 181 1662 182 se
rect 1662 181 1807 204
rect 1078 180 1079 181
tri 1079 180 1080 181 sw
tri 1308 180 1309 181 se
rect 1309 180 1310 181
rect 1356 180 1357 181
tri 1357 180 1358 181 sw
tri 1660 180 1661 181 se
rect 1661 180 1807 181
rect 1032 175 1080 180
tri 1080 175 1085 180 sw
tri 1303 175 1308 180 se
rect 1308 175 1358 180
tri 1358 175 1363 180 sw
tri 1655 175 1660 180 se
rect 1660 175 1807 180
rect 902 157 955 175
tri 955 157 973 175 sw
tri 1007 157 1025 175 se
rect 1025 157 1085 175
tri 1085 157 1103 175 sw
tri 1285 157 1303 175 se
rect 1303 157 1363 175
tri 1363 157 1381 175 sw
tri 1637 157 1655 175 se
rect 1655 157 1807 175
rect 902 123 908 157
rect 942 151 1668 157
rect 942 123 980 151
rect 902 117 980 123
rect 1014 117 1057 151
rect 1091 117 1134 151
rect 1168 117 1211 151
rect 1245 117 1288 151
rect 1322 117 1365 151
rect 1399 117 1442 151
rect 1476 117 1519 151
rect 1553 117 1596 151
rect 1630 123 1668 151
rect 1702 123 1807 157
rect 1630 117 1807 123
rect 902 111 1807 117
rect 1849 2157 1895 2197
rect 1849 2123 1855 2157
rect 1889 2123 1895 2157
rect 1849 2083 1895 2123
rect 1849 2049 1855 2083
rect 1889 2049 1895 2083
rect 1849 2009 1895 2049
rect 1849 1975 1855 2009
rect 1889 1975 1895 2009
rect 1849 1935 1895 1975
rect 1849 1901 1855 1935
rect 1889 1901 1895 1935
rect 1849 1861 1895 1901
rect 1849 1827 1855 1861
rect 1889 1827 1895 1861
rect 1849 1787 1895 1827
rect 1849 1753 1855 1787
rect 1889 1753 1895 1787
rect 1849 1713 1895 1753
rect 1849 1679 1855 1713
rect 1889 1679 1895 1713
rect 1849 1639 1895 1679
rect 1849 1605 1855 1639
rect 1889 1605 1895 1639
rect 1849 1565 1895 1605
rect 1849 1531 1855 1565
rect 1889 1531 1895 1565
rect 1849 1491 1895 1531
rect 1849 1457 1855 1491
rect 1889 1457 1895 1491
rect 1849 1417 1895 1457
rect 1849 1383 1855 1417
rect 1889 1383 1895 1417
rect 1849 1343 1895 1383
rect 1849 1309 1855 1343
rect 1889 1309 1895 1343
rect 1849 1270 1895 1309
rect 1849 1236 1855 1270
rect 1889 1236 1895 1270
rect 1849 1197 1895 1236
rect 1849 1163 1855 1197
rect 1889 1163 1895 1197
rect 1849 1124 1895 1163
rect 1849 1090 1855 1124
rect 1889 1090 1895 1124
rect 1849 1051 1895 1090
rect 1849 1017 1855 1051
rect 1889 1017 1895 1051
rect 1849 978 1895 1017
rect 1849 944 1855 978
rect 1889 944 1895 978
rect 1849 905 1895 944
rect 1849 871 1855 905
rect 1889 871 1895 905
rect 1849 832 1895 871
rect 1849 798 1855 832
rect 1889 798 1895 832
rect 1849 759 1895 798
rect 1849 725 1855 759
rect 1889 725 1895 759
rect 1849 686 1895 725
rect 1849 652 1855 686
rect 1889 652 1895 686
rect 1849 613 1895 652
rect 1849 579 1855 613
rect 1889 579 1895 613
rect 1849 540 1895 579
rect 1849 506 1855 540
rect 1889 506 1895 540
rect 1849 467 1895 506
rect 1849 433 1855 467
rect 1889 433 1895 467
rect 1849 394 1895 433
rect 1849 360 1855 394
rect 1889 360 1895 394
rect 1849 321 1895 360
rect 1849 287 1855 321
rect 1889 287 1895 321
rect 1849 248 1895 287
rect 1849 214 1855 248
rect 1889 214 1895 248
rect 1849 175 1895 214
rect 1849 141 1855 175
rect 1889 141 1895 175
rect 715 43 767 62
rect 1849 102 1895 141
rect 1849 68 1855 102
rect 1889 68 1895 102
rect 1849 29 1895 68
rect 715 -15 767 -9
rect 1573 21 1625 27
rect 353 -45 405 -39
tri 1558 -45 1573 -30 se
rect 1849 -5 1855 29
rect 1889 -5 1895 29
rect 1849 -17 1895 -5
rect 1573 -43 1625 -31
tri 1557 -46 1558 -45 se
rect 1558 -46 1573 -45
rect 354 -47 404 -46
tri 1556 -47 1557 -46 se
rect 1557 -47 1573 -46
rect 353 -83 405 -47
tri 1548 -55 1556 -47 se
rect 1556 -55 1573 -47
rect 354 -84 404 -83
tri 405 -84 406 -83 sw
rect 405 -85 406 -84
tri 406 -85 407 -84 sw
rect 353 -101 407 -85
tri 407 -101 423 -85 sw
tri 1625 -55 1650 -30 sw
rect 1573 -101 1625 -95
rect 353 -108 423 -101
tri 423 -108 430 -101 sw
rect 353 -137 430 -108
<< rmetal1 >>
rect -1055 4536 -1009 4537
rect -1055 4535 -1054 4536
rect -1010 4535 -1009 4536
rect -743 4536 -697 4537
rect -743 4535 -742 4536
rect -698 4535 -697 4536
rect -1055 4498 -1054 4499
rect -1010 4498 -1009 4499
rect -1055 4497 -1009 4498
rect -743 4498 -742 4499
rect -698 4498 -697 4499
rect -743 4497 -697 4498
rect -1114 4404 -1068 4405
rect -1114 4403 -1113 4404
rect -1069 4403 -1068 4404
rect -1114 4366 -1113 4367
rect -1069 4366 -1068 4367
rect -1114 4365 -1068 4366
rect -1739 4242 -1737 4243
rect -1739 4187 -1738 4242
rect -1739 4186 -1737 4187
rect -1701 4242 -1699 4243
rect -1700 4187 -1699 4242
rect -802 4404 -756 4405
rect -802 4403 -801 4404
rect -757 4403 -756 4404
rect -802 4366 -801 4367
rect -757 4366 -756 4367
rect -802 4365 -756 4366
rect -1701 4186 -1699 4187
rect -993 3795 -947 3796
rect -993 3794 -992 3795
rect -948 3794 -947 3795
rect -993 3757 -992 3758
rect -948 3757 -947 3758
rect -993 3756 -947 3757
rect -993 3625 -947 3626
rect -993 3624 -992 3625
rect -948 3624 -947 3625
rect -646 3646 -600 3647
rect -646 3645 -645 3646
rect -601 3645 -600 3646
rect -646 3608 -645 3609
rect -601 3608 -600 3609
rect -646 3607 -600 3608
rect -993 3587 -992 3588
rect -948 3587 -947 3588
rect -993 3586 -947 3587
rect 435 2418 437 2419
rect 435 2378 436 2418
rect 435 2377 437 2378
rect 473 2418 475 2419
rect 474 2378 475 2418
rect 473 2377 475 2378
rect 1310 2085 1356 2086
rect 1310 2084 1311 2085
rect 1355 2084 1356 2085
rect 998 2050 1044 2051
rect 998 2049 999 2050
rect 1043 2049 1044 2050
rect 998 2012 999 2013
rect 1043 2012 1044 2013
rect 998 2011 1044 2012
rect 1310 2047 1311 2048
rect 1355 2047 1356 2048
rect 1310 2046 1356 2047
rect 1235 1761 1237 1762
rect 1235 1717 1236 1761
rect 1235 1716 1237 1717
rect 1273 1761 1275 1762
rect 1274 1717 1275 1761
rect 1273 1716 1275 1717
rect 1154 1549 1200 1550
rect 1154 1548 1155 1549
rect 1199 1548 1200 1549
rect 1566 1638 1612 1639
rect 1566 1637 1567 1638
rect 1611 1637 1612 1638
rect 1566 1600 1567 1601
rect 1611 1600 1612 1601
rect 1566 1599 1612 1600
rect 1154 1511 1155 1512
rect 1199 1511 1200 1512
rect 1154 1510 1200 1511
rect 78 1484 80 1485
rect 116 1484 118 1485
rect 78 1440 79 1484
rect 117 1440 118 1484
rect 339 1484 341 1485
rect 78 1439 80 1440
rect 116 1439 118 1440
rect 339 1440 340 1484
rect 339 1439 341 1440
rect 377 1484 379 1485
rect 378 1440 379 1484
rect 533 1484 535 1485
rect 571 1484 573 1485
rect 377 1439 379 1440
rect 533 1440 534 1484
rect 572 1440 573 1484
rect 533 1439 535 1440
rect 571 1439 573 1440
rect 1154 755 1200 756
rect 1154 754 1155 755
rect 1199 754 1200 755
rect 353 588 405 589
rect 353 587 354 588
rect 404 587 405 588
rect 353 550 354 551
rect 404 550 405 551
rect 353 549 405 550
rect 273 -46 325 -45
rect 273 -47 274 -46
rect 324 -47 325 -46
rect 273 -84 274 -83
rect 324 -84 325 -83
rect 273 -85 325 -84
rect 1154 717 1155 718
rect 1199 717 1200 718
rect 1154 716 1200 717
rect 1566 666 1612 667
rect 1566 665 1567 666
rect 1611 665 1612 666
rect 1235 549 1237 550
rect 1235 505 1236 549
rect 1235 504 1237 505
rect 1273 549 1275 550
rect 1274 505 1275 549
rect 1273 504 1275 505
rect 1032 219 1078 220
rect 1032 218 1033 219
rect 1077 218 1078 219
rect 1310 219 1356 220
rect 1310 218 1311 219
rect 1355 218 1356 219
rect 1566 628 1567 629
rect 1611 628 1612 629
rect 1566 627 1612 628
rect 1032 181 1033 182
rect 1077 181 1078 182
rect 1310 181 1311 182
rect 1355 181 1356 182
rect 1032 180 1078 181
rect 1310 180 1356 181
rect 353 -46 405 -45
rect 353 -47 354 -46
rect 404 -47 405 -46
rect 353 -84 354 -83
rect 404 -84 405 -83
rect 353 -85 405 -84
<< via1 >>
rect -1151 5023 -1099 5075
rect -1074 5023 -1022 5075
rect -996 5023 -944 5075
rect 2001 5023 2053 5075
rect 2072 5023 2124 5075
rect 2144 5023 2196 5075
rect 2216 5023 2268 5075
rect 2288 5023 2340 5075
rect -1151 4959 -1099 5011
rect -1074 4959 -1022 5011
rect -996 4959 -944 5011
rect 2001 4959 2053 5011
rect 2072 4959 2124 5011
rect 2144 4959 2196 5011
rect 2216 4959 2268 5011
rect 2288 4959 2340 5011
rect -748 4841 -696 4893
rect -653 4851 -601 4903
rect -589 4851 -537 4903
rect 277 4851 329 4903
rect 341 4851 393 4903
rect 405 4851 457 4903
rect -882 4761 -830 4813
rect -748 4777 -696 4829
rect 832 4771 884 4823
rect 896 4771 948 4823
rect -882 4697 -830 4749
rect 750 4691 802 4743
rect 814 4691 866 4743
rect -1562 4536 -1510 4588
rect -1498 4536 -1446 4588
rect 523 4641 575 4653
rect 590 4641 642 4653
rect 658 4641 710 4653
rect 523 4607 538 4641
rect 538 4607 575 4641
rect 590 4607 612 4641
rect 612 4607 642 4641
rect 658 4607 686 4641
rect 686 4607 710 4641
rect 523 4601 575 4607
rect 590 4601 642 4607
rect 658 4601 710 4607
rect 277 4557 329 4573
rect 277 4523 292 4557
rect 292 4523 329 4557
rect 277 4521 329 4523
rect 341 4521 393 4573
rect 405 4521 457 4573
rect -1652 4258 -1600 4310
rect -1652 4192 -1600 4244
rect -882 4329 -830 4381
rect -882 4247 -830 4299
rect -668 4359 -636 4381
rect -636 4359 -616 4381
rect -668 4329 -616 4359
rect -668 4250 -616 4262
rect -668 4216 -636 4250
rect -636 4216 -616 4250
rect -668 4210 -616 4216
rect -560 4307 -508 4359
rect -496 4353 -444 4359
rect -496 4319 -484 4353
rect -484 4319 -450 4353
rect -450 4319 -444 4353
rect -496 4307 -444 4319
rect -560 4217 -508 4269
rect -496 4260 -444 4269
rect -496 4226 -484 4260
rect -484 4226 -450 4260
rect -450 4226 -444 4260
rect -496 4217 -444 4226
rect -560 4127 -508 4179
rect -496 4167 -444 4179
rect -496 4133 -484 4167
rect -484 4133 -450 4167
rect -450 4133 -444 4167
rect -496 4127 -444 4133
rect -1572 4048 -1520 4100
rect -1572 3982 -1520 4034
rect -1492 3587 -1440 3639
rect -1492 3557 -1440 3575
rect -1492 3523 -1458 3557
rect -1458 3523 -1440 3557
rect -738 3532 -686 3584
rect -674 3532 -622 3584
rect -560 3376 -508 3405
rect -560 3353 -546 3376
rect -546 3353 -508 3376
rect -496 3353 -444 3405
rect -560 3279 -508 3315
rect -560 3263 -546 3279
rect -546 3263 -508 3279
rect -496 3263 -444 3315
rect -238 4341 -232 4359
rect -232 4341 -198 4359
rect -198 4341 -186 4359
rect -238 4307 -186 4341
rect -238 4268 -232 4269
rect -232 4268 -198 4269
rect -198 4268 -186 4269
rect -238 4229 -186 4268
rect -238 4217 -232 4229
rect -232 4217 -198 4229
rect -198 4217 -186 4229
rect -238 4156 -186 4179
rect -238 4127 -232 4156
rect -232 4127 -198 4156
rect -198 4127 -186 4156
rect -238 3395 -232 3405
rect -232 3395 -198 3405
rect -198 3395 -186 3405
rect -238 3357 -186 3395
rect -238 3353 -232 3357
rect -232 3353 -198 3357
rect -198 3353 -186 3357
rect -238 3285 -186 3315
rect -238 3263 -232 3285
rect -232 3263 -198 3285
rect -198 3263 -186 3285
rect -1492 3165 -1440 3217
rect -560 3207 -508 3225
rect -560 3173 -540 3207
rect -540 3173 -508 3207
rect -496 3207 -444 3225
rect -238 3213 -186 3225
rect -496 3173 -484 3207
rect -484 3173 -450 3207
rect -450 3173 -444 3207
rect -238 3179 -232 3213
rect -232 3179 -198 3213
rect -198 3179 -186 3213
rect -238 3173 -186 3179
rect -1572 3091 -1520 3143
rect -1492 3099 -1440 3151
rect -1572 3025 -1520 3077
rect -1646 2930 -1594 2982
rect -1580 2930 -1528 2982
rect 820 4403 872 4455
rect 820 4339 872 4391
rect 820 4275 872 4327
rect 820 4211 872 4263
rect 914 4415 966 4467
rect 914 4351 966 4403
rect 914 4287 966 4339
rect 914 4223 966 4275
rect 820 4147 872 4199
rect 820 4083 872 4135
rect 820 4019 872 4071
rect 820 3955 872 4007
rect 820 3891 872 3943
rect 820 3827 872 3879
rect 820 3763 872 3815
rect 820 3699 872 3751
rect 820 3635 872 3687
rect 820 3570 872 3622
rect 820 3505 872 3557
rect 820 3440 872 3492
rect 820 3375 872 3427
rect 820 3310 872 3362
rect 820 3245 872 3297
rect 820 3180 872 3232
rect 820 3115 872 3167
rect 820 3050 872 3102
rect 820 2985 872 3037
rect 820 2920 872 2972
rect 820 2855 872 2907
rect 820 2790 872 2842
rect 820 2725 872 2777
rect 820 2660 872 2712
rect 820 2595 872 2647
rect 820 2530 872 2582
rect 820 2465 872 2517
rect 90 2361 142 2413
rect 90 2295 142 2347
rect 715 2309 716 2312
rect 716 2309 750 2312
rect 750 2309 767 2312
rect 715 2271 767 2309
rect 715 2260 721 2271
rect 721 2260 755 2271
rect 755 2260 767 2271
rect 715 2237 721 2245
rect 721 2237 755 2245
rect 755 2237 767 2245
rect 90 2175 142 2181
rect 90 2141 108 2175
rect 108 2141 142 2175
rect 90 2129 142 2141
rect 90 2089 142 2114
rect 90 2062 108 2089
rect 108 2062 142 2089
rect 90 2003 142 2046
rect 90 1994 108 2003
rect 108 1994 142 2003
rect 90 1969 108 1978
rect 108 1969 142 1978
rect 90 1926 142 1969
rect 90 1883 108 1910
rect 108 1883 142 1910
rect 90 1858 142 1883
rect 90 1830 142 1842
rect 90 1796 108 1830
rect 108 1796 142 1830
rect 90 1790 142 1796
rect 513 2168 565 2220
rect 590 2214 642 2220
rect 590 2180 602 2214
rect 602 2180 636 2214
rect 636 2180 642 2214
rect 590 2168 642 2180
rect 513 2099 565 2151
rect 590 2141 642 2151
rect 590 2107 602 2141
rect 602 2107 636 2141
rect 636 2107 642 2141
rect 590 2099 642 2107
rect 287 1704 339 1756
rect 353 1704 405 1756
rect 513 2030 565 2082
rect 590 2067 642 2082
rect 590 2033 602 2067
rect 602 2033 636 2067
rect 636 2033 642 2067
rect 590 2030 642 2033
rect 513 1961 565 2013
rect 590 1993 642 2013
rect 590 1961 602 1993
rect 602 1961 636 1993
rect 636 1961 642 1993
rect 513 1892 565 1944
rect 590 1919 642 1944
rect 590 1892 602 1919
rect 602 1892 636 1919
rect 636 1892 642 1919
rect 513 1823 565 1875
rect 590 1845 642 1875
rect 590 1823 602 1845
rect 602 1823 636 1845
rect 636 1823 642 1845
rect 513 1753 565 1805
rect 590 1771 642 1805
rect 590 1753 602 1771
rect 602 1753 636 1771
rect 636 1753 642 1771
rect 715 2193 767 2237
rect 715 2153 721 2179
rect 721 2153 755 2179
rect 755 2153 767 2179
rect 715 2127 767 2153
rect 715 2103 767 2113
rect 715 2069 721 2103
rect 721 2069 755 2103
rect 755 2069 767 2103
rect 914 2217 966 2269
rect 914 2153 966 2205
rect 914 2089 966 2141
rect 715 2061 767 2069
rect 715 2020 767 2047
rect 715 1995 721 2020
rect 721 1995 755 2020
rect 755 1995 767 2020
rect 715 1937 767 1981
rect 715 1929 721 1937
rect 721 1929 755 1937
rect 755 1929 767 1937
rect 715 1903 721 1915
rect 721 1903 755 1915
rect 755 1903 767 1915
rect 715 1863 767 1903
rect 715 1820 721 1849
rect 721 1820 755 1849
rect 755 1820 767 1849
rect 715 1797 767 1820
rect 715 1771 767 1783
rect 715 1737 721 1771
rect 721 1737 755 1771
rect 755 1737 767 1771
rect 715 1731 767 1737
rect 353 1609 405 1661
rect 715 1613 767 1619
rect 190 1587 242 1593
rect 190 1553 202 1587
rect 202 1553 236 1587
rect 236 1553 242 1587
rect 190 1541 242 1553
rect 256 1541 308 1593
rect 353 1587 405 1595
rect 353 1553 392 1587
rect 392 1553 405 1587
rect 353 1543 405 1553
rect 715 1579 721 1613
rect 721 1579 755 1613
rect 755 1579 767 1613
rect 715 1567 767 1579
rect 715 1535 767 1553
rect 715 1501 721 1535
rect 721 1501 755 1535
rect 755 1501 767 1535
rect 513 1297 565 1349
rect 513 1220 565 1272
rect 433 1119 485 1171
rect 433 1055 485 1107
rect 513 1143 565 1195
rect 513 1066 565 1118
rect 513 989 565 1041
rect 439 904 491 956
rect 439 829 491 881
rect 439 753 491 805
rect 715 1457 767 1487
rect 715 1435 721 1457
rect 721 1435 755 1457
rect 755 1435 767 1457
rect 715 1380 767 1421
rect 715 1369 721 1380
rect 721 1369 755 1380
rect 755 1369 767 1380
rect 1573 1375 1579 1409
rect 1579 1375 1613 1409
rect 1613 1375 1625 1409
rect 715 1346 721 1355
rect 721 1346 755 1355
rect 755 1346 767 1355
rect 715 1303 767 1346
rect 1573 1357 1625 1375
rect 1573 1293 1625 1345
rect 715 1269 721 1289
rect 721 1269 755 1289
rect 755 1269 767 1289
rect 715 1237 767 1269
rect 715 1192 721 1223
rect 721 1192 755 1223
rect 755 1192 767 1223
rect 715 1171 767 1192
rect 715 1149 767 1157
rect 715 1115 721 1149
rect 721 1115 755 1149
rect 755 1115 767 1149
rect 715 1105 767 1115
rect 715 1072 767 1091
rect 715 1039 721 1072
rect 721 1039 755 1072
rect 755 1039 767 1072
rect 715 995 767 1025
rect 715 973 721 995
rect 721 973 755 995
rect 755 973 767 995
rect 715 918 767 959
rect 715 907 721 918
rect 721 907 755 918
rect 755 907 767 918
rect 1573 921 1625 973
rect 715 884 721 894
rect 721 884 755 894
rect 755 884 767 894
rect 715 842 767 884
rect 1573 891 1625 909
rect 1573 857 1579 891
rect 1579 857 1613 891
rect 1613 857 1625 891
rect 715 807 721 829
rect 721 807 755 829
rect 755 807 767 829
rect 715 777 767 807
rect 715 730 721 764
rect 721 730 755 764
rect 755 730 767 764
rect 273 661 325 713
rect 273 595 325 647
rect 353 679 389 713
rect 389 679 405 713
rect 353 661 405 679
rect 715 712 767 730
rect 715 687 767 699
rect 715 653 721 687
rect 721 653 755 687
rect 755 653 767 687
rect 353 595 405 647
rect 715 647 767 653
rect 90 568 142 574
rect 90 534 108 568
rect 108 534 142 568
rect 90 522 142 534
rect 90 487 142 504
rect 90 453 108 487
rect 108 453 142 487
rect 90 452 142 453
rect 90 406 142 434
rect 90 382 108 406
rect 108 382 142 406
rect 449 247 501 299
rect 513 247 565 299
rect 449 180 501 232
rect 513 180 565 232
rect 449 112 501 164
rect 513 112 565 164
rect 715 529 767 535
rect 715 495 721 529
rect 721 495 755 529
rect 755 495 767 529
rect 715 483 767 495
rect 715 446 767 465
rect 715 413 721 446
rect 721 413 755 446
rect 755 413 767 446
rect 715 363 767 395
rect 715 343 721 363
rect 721 343 755 363
rect 755 343 767 363
rect 715 280 767 325
rect 715 273 721 280
rect 721 273 755 280
rect 755 273 767 280
rect 715 246 721 255
rect 721 246 755 255
rect 755 246 767 255
rect 715 203 767 246
rect 715 163 721 185
rect 721 163 755 185
rect 755 163 767 185
rect 715 133 767 163
rect 273 27 325 79
rect 273 -39 325 13
rect 353 27 405 79
rect 353 -39 405 13
rect 715 80 721 114
rect 721 80 755 114
rect 755 80 767 114
rect 715 62 767 80
rect 715 31 767 43
rect 715 -3 721 31
rect 721 -3 755 31
rect 755 -3 767 31
rect 715 -9 767 -3
rect 1573 -31 1625 21
rect 1573 -95 1625 -43
<< metal2 >>
rect -2092 4733 -1618 5075
rect -2092 4697 -1654 4733
tri -1654 4697 -1618 4733 nw
rect -1505 4733 -1185 5075
tri -1505 4697 -1469 4733 ne
rect -1469 4697 -1185 4733
rect -2092 4691 -1660 4697
tri -1660 4691 -1654 4697 nw
tri -1469 4691 -1463 4697 ne
rect -1463 4691 -1185 4697
rect -2092 4653 -1698 4691
tri -1698 4653 -1660 4691 nw
tri -1463 4653 -1425 4691 ne
rect -1425 4653 -1185 4691
rect -2092 2855 -1708 4653
tri -1708 4643 -1698 4653 nw
tri -1425 4643 -1415 4653 ne
rect -1415 4643 -1185 4653
tri -1415 4624 -1396 4643 ne
rect -1568 4536 -1562 4588
rect -1510 4536 -1498 4588
rect -1446 4536 -1440 4588
tri -1517 4521 -1502 4536 ne
rect -1502 4521 -1440 4536
tri -1502 4511 -1492 4521 ne
rect -1652 4310 -1600 4316
rect -1652 4244 -1600 4258
rect -1652 2985 -1600 4192
rect -1572 4100 -1520 4106
rect -1572 4034 -1520 4048
rect -1572 3143 -1520 3982
rect -1492 3639 -1440 4521
rect -1492 3575 -1440 3587
rect -1492 3217 -1440 3523
rect -1492 3151 -1440 3165
rect -1492 3093 -1440 3099
rect -1572 3077 -1520 3091
rect -1572 3019 -1520 3025
tri -1600 2985 -1578 3007 sw
rect -1652 2982 -1578 2985
tri -1578 2982 -1575 2985 sw
rect -1652 2930 -1646 2982
rect -1594 2930 -1580 2982
rect -1528 2930 -1522 2982
tri -1400 2972 -1396 2976 se
rect -1396 2972 -1185 4643
tri -1442 2930 -1400 2972 se
rect -1400 2930 -1185 2972
tri -1452 2920 -1442 2930 se
rect -1442 2920 -1185 2930
tri -1465 2907 -1452 2920 se
rect -1452 2907 -1185 2920
tri -1466 2906 -1465 2907 se
rect -1465 2906 -1185 2907
tri -1708 2855 -1657 2906 sw
tri -1505 2867 -1466 2906 se
rect -1466 2867 -1185 2906
rect -2092 2842 -1657 2855
tri -1657 2842 -1644 2855 sw
rect -2092 2816 -1644 2842
tri -1644 2816 -1618 2842 sw
rect -2092 2498 -1618 2816
rect -1505 2498 -1185 2867
rect -1157 5023 -1151 5075
rect -1099 5023 -1074 5075
rect -1022 5023 -996 5075
rect -944 5023 -938 5075
rect -1157 5011 -938 5023
rect -1157 4959 -1151 5011
rect -1099 4959 -1074 5011
rect -1022 4959 -996 5011
rect -944 4959 -938 5011
rect -1157 4127 -938 4959
rect -748 4893 -696 4899
rect -748 4829 -696 4841
rect -882 4813 -830 4819
rect -882 4749 -830 4761
rect -882 4381 -830 4697
rect -882 4299 -830 4329
rect -882 4241 -830 4247
tri -938 4127 -886 4179 sw
rect -1157 4106 -886 4127
tri -886 4106 -865 4127 sw
rect -1157 4083 -865 4106
tri -865 4083 -842 4106 sw
rect -1157 4071 -842 4083
tri -842 4071 -830 4083 sw
rect -1157 4045 -830 4071
tri -830 4045 -804 4071 sw
rect -1157 2498 -804 4045
rect -748 3584 -696 4777
rect -668 4851 -653 4903
rect -601 4851 -589 4903
rect -537 4851 -531 4903
rect -668 4381 -616 4851
tri -616 4826 -591 4851 nw
tri -143 4467 -103 4507 se
rect -103 4467 217 5075
rect 271 4851 277 4903
rect 329 4851 341 4903
rect 393 4851 405 4903
rect 457 4851 463 4903
tri 271 4826 296 4851 ne
tri 286 4588 296 4598 se
rect 296 4588 348 4851
tri 348 4826 373 4851 nw
rect 517 4653 716 5075
rect 1995 5023 2001 5075
rect 2053 5023 2072 5075
rect 2124 5023 2144 5075
rect 2196 5023 2216 5075
rect 2268 5023 2288 5075
rect 2340 5023 2346 5075
rect 1995 5011 2346 5023
rect 1995 4959 2001 5011
rect 2053 4959 2072 5011
rect 2124 4959 2144 5011
rect 2196 4959 2216 5011
rect 2268 4959 2288 5011
rect 2340 4959 2346 5011
rect 826 4771 832 4823
rect 884 4771 896 4823
rect 948 4811 954 4823
tri 954 4811 966 4823 sw
rect 948 4771 966 4811
tri 889 4746 914 4771 ne
rect 744 4691 750 4743
rect 802 4691 814 4743
rect 866 4691 872 4743
tri 795 4666 820 4691 ne
rect 517 4601 523 4653
rect 575 4601 590 4653
rect 642 4601 658 4653
rect 710 4601 716 4653
tri 348 4588 358 4598 sw
tri 271 4573 286 4588 se
rect 286 4573 358 4588
tri 358 4573 373 4588 sw
rect 271 4521 277 4573
rect 329 4521 341 4573
rect 393 4521 405 4573
rect 457 4521 463 4573
tri -155 4455 -143 4467 se
rect -143 4455 217 4467
tri -207 4403 -155 4455 se
rect -155 4403 217 4455
tri -219 4391 -207 4403 se
rect -207 4391 217 4403
tri -223 4387 -219 4391 se
rect -219 4387 217 4391
tri -245 4365 -223 4387 se
rect -223 4365 217 4387
rect -668 4262 -616 4329
rect -668 4204 -616 4210
rect -560 4359 217 4365
rect -508 4307 -496 4359
rect -444 4307 -238 4359
rect -186 4307 217 4359
rect -560 4269 217 4307
rect -508 4217 -496 4269
rect -444 4217 -238 4269
rect -186 4217 217 4269
rect -560 4179 217 4217
rect -508 4127 -496 4179
rect -444 4127 -238 4179
rect -186 4127 217 4179
rect -560 4121 217 4127
tri -245 4083 -207 4121 ne
rect -207 4083 217 4121
tri -207 4071 -195 4083 ne
rect -195 4071 217 4083
tri -195 4019 -143 4071 ne
rect -143 4019 217 4071
tri -143 4007 -131 4019 ne
rect -131 4007 217 4019
tri -131 3979 -103 4007 ne
tri -696 3584 -671 3609 sw
rect -748 3532 -738 3584
rect -686 3532 -674 3584
rect -622 3532 -616 3584
tri -124 3532 -103 3553 se
rect -103 3532 217 4007
tri -139 3517 -124 3532 se
rect -124 3517 217 3532
tri -151 3505 -139 3517 se
rect -139 3505 217 3517
tri -164 3492 -151 3505 se
rect -151 3492 217 3505
tri -216 3440 -164 3492 se
rect -164 3440 217 3492
tri -229 3427 -216 3440 se
rect -216 3427 217 3440
tri -245 3411 -229 3427 se
rect -229 3411 217 3427
rect -560 3405 217 3411
rect -508 3353 -496 3405
rect -444 3353 -238 3405
rect -186 3353 217 3405
rect -560 3315 217 3353
rect -508 3263 -496 3315
rect -444 3263 -238 3315
rect -186 3263 217 3315
rect -560 3225 217 3263
rect -508 3173 -496 3225
rect -444 3173 -238 3225
rect -186 3173 217 3225
rect -560 3167 217 3173
tri -245 3149 -227 3167 ne
rect -227 3149 217 3167
tri -227 3115 -193 3149 ne
rect -193 3115 217 3149
tri -193 3102 -180 3115 ne
rect -180 3102 217 3115
tri -180 3050 -128 3102 ne
rect -128 3050 217 3102
tri -128 3037 -115 3050 ne
rect -115 3037 217 3050
tri -115 3025 -103 3037 ne
rect -103 2462 217 3037
rect -103 2455 80 2462
tri 80 2455 87 2462 nw
tri 145 2455 152 2462 ne
rect 152 2455 217 2462
rect 517 2465 716 4601
rect 820 4455 872 4691
rect 820 4391 872 4403
rect 820 4327 872 4339
rect 820 4263 872 4275
rect 820 4199 872 4211
rect 820 4135 872 4147
rect 820 4071 872 4083
rect 820 4007 872 4019
rect 820 3943 872 3955
rect 820 3879 872 3891
rect 820 3815 872 3827
rect 820 3751 872 3763
rect 820 3687 872 3699
rect 820 3622 872 3635
rect 820 3557 872 3570
rect 820 3492 872 3505
rect 820 3427 872 3440
rect 820 3362 872 3375
rect 820 3297 872 3310
rect 820 3232 872 3245
rect 820 3167 872 3180
rect 820 3102 872 3115
rect 820 3037 872 3050
rect 820 2972 872 2985
rect 820 2907 872 2920
rect 820 2842 872 2855
rect 820 2777 872 2790
rect 820 2712 872 2725
rect 820 2647 872 2660
rect 820 2582 872 2595
rect 820 2517 872 2530
tri 716 2465 768 2517 sw
rect 517 2459 768 2465
tri 768 2459 774 2465 sw
rect 820 2459 872 2465
rect 914 4467 966 4771
rect 914 4403 966 4415
rect 914 4339 966 4351
rect 914 4275 966 4287
rect -103 343 62 2455
tri 62 2437 80 2455 nw
tri 152 2437 170 2455 ne
rect 90 2413 142 2419
rect 90 2347 142 2361
rect 90 2181 142 2295
rect 90 2114 142 2129
rect 90 2046 142 2062
rect 90 1978 142 1994
rect 90 1910 142 1926
rect 90 1842 142 1858
rect 90 574 142 1790
rect 170 1621 217 2455
tri 513 2451 517 2455 se
rect 517 2451 774 2459
rect 513 2347 774 2451
tri 774 2347 886 2459 sw
rect 513 2312 886 2347
rect 513 2260 715 2312
rect 767 2260 886 2312
rect 513 2245 886 2260
rect 513 2220 715 2245
rect 565 2168 590 2220
rect 642 2193 715 2220
rect 767 2193 886 2245
rect 642 2179 886 2193
rect 642 2168 715 2179
rect 513 2151 715 2168
rect 565 2099 590 2151
rect 642 2127 715 2151
rect 767 2127 886 2179
rect 642 2113 886 2127
rect 642 2099 715 2113
rect 513 2082 715 2099
rect 565 2030 590 2082
rect 642 2061 715 2082
rect 767 2061 886 2113
rect 642 2047 886 2061
rect 642 2030 715 2047
rect 513 2013 715 2030
rect 565 1961 590 2013
rect 642 1995 715 2013
rect 767 1995 886 2047
rect 642 1981 886 1995
rect 642 1961 715 1981
rect 513 1944 715 1961
rect 565 1892 590 1944
rect 642 1929 715 1944
rect 767 1929 886 1981
rect 642 1915 886 1929
rect 642 1892 715 1915
rect 513 1875 715 1892
rect 565 1823 590 1875
rect 642 1863 715 1875
rect 767 1863 886 1915
rect 642 1849 886 1863
rect 642 1823 715 1849
rect 513 1805 715 1823
rect 281 1704 287 1756
rect 339 1704 353 1756
rect 405 1704 485 1756
tri 408 1679 433 1704 ne
rect 353 1661 405 1667
rect 353 1595 405 1609
rect 184 1541 190 1593
rect 242 1541 256 1593
rect 308 1541 325 1593
tri 248 1516 273 1541 ne
rect 90 504 142 522
rect 90 434 142 452
rect 90 376 142 382
tri 62 343 77 358 sw
tri 155 343 170 358 se
rect 170 343 210 1513
rect -103 333 77 343
tri 77 333 87 343 sw
tri 145 333 155 343 se
rect 155 333 210 343
rect -103 86 210 333
rect 273 713 325 1541
rect 273 647 325 661
rect 273 79 325 595
rect 273 13 325 27
rect 273 -45 325 -39
rect 353 713 405 1543
rect 433 1171 485 1704
rect 433 1107 485 1119
rect 433 1049 485 1055
rect 565 1753 590 1805
rect 642 1797 715 1805
rect 767 1797 886 1849
rect 642 1783 886 1797
rect 642 1753 715 1783
rect 513 1731 715 1753
rect 767 1731 886 1783
rect 513 1619 886 1731
rect 914 2269 966 4223
rect 914 2205 966 2217
rect 914 2141 966 2153
rect 914 1800 966 2089
tri 966 1800 988 1822 sw
tri 914 1726 988 1800 ne
tri 988 1726 1062 1800 sw
tri 988 1725 989 1726 ne
rect 989 1725 1062 1726
tri 989 1652 1062 1725 ne
tri 1062 1672 1116 1726 sw
rect 1062 1652 1116 1672
tri 1062 1650 1064 1652 ne
rect 513 1567 715 1619
rect 767 1567 886 1619
rect 513 1553 886 1567
rect 513 1501 715 1553
rect 767 1501 886 1553
rect 513 1487 886 1501
rect 513 1435 715 1487
rect 767 1435 886 1487
rect 1064 1527 1116 1652
rect 1064 1475 1967 1527
rect 513 1421 886 1435
rect 513 1369 715 1421
rect 767 1369 886 1421
rect 513 1355 886 1369
rect 513 1349 715 1355
rect 565 1303 715 1349
rect 767 1303 886 1355
rect 565 1297 886 1303
rect 513 1289 886 1297
rect 513 1272 715 1289
rect 565 1237 715 1272
rect 767 1237 886 1289
rect 565 1223 886 1237
rect 565 1220 715 1223
rect 513 1195 715 1220
rect 565 1171 715 1195
rect 767 1171 886 1223
rect 565 1157 886 1171
rect 565 1143 715 1157
rect 513 1118 715 1143
rect 565 1105 715 1118
rect 767 1105 886 1157
rect 565 1091 886 1105
rect 565 1066 715 1091
rect 513 1041 715 1066
tri 466 989 513 1036 se
rect 565 1039 715 1041
rect 767 1039 886 1091
rect 565 1025 886 1039
rect 565 989 715 1025
tri 460 983 466 989 se
rect 466 983 715 989
tri 450 973 460 983 se
rect 460 973 715 983
rect 767 973 886 1025
tri 439 962 450 973 se
rect 450 962 886 973
tri 436 959 439 962 se
rect 439 959 886 962
rect 353 647 405 661
rect 353 79 405 595
rect 353 13 405 27
tri 433 956 436 959 se
rect 436 956 715 959
rect 433 904 439 956
rect 491 907 715 956
rect 767 907 886 959
rect 491 904 886 907
rect 433 894 886 904
rect 433 881 715 894
rect 433 829 439 881
rect 491 842 715 881
rect 767 842 886 894
rect 491 829 886 842
rect 433 805 715 829
rect 433 753 439 805
rect 491 777 715 805
rect 767 777 886 829
rect 491 764 886 777
rect 491 753 715 764
rect 433 712 715 753
rect 767 712 886 764
rect 433 699 886 712
rect 433 647 715 699
rect 767 647 886 699
rect 433 535 886 647
rect 433 483 715 535
rect 767 483 886 535
rect 433 465 886 483
rect 433 413 715 465
rect 767 413 886 465
rect 433 395 886 413
rect 433 343 715 395
rect 767 343 886 395
rect 433 325 886 343
rect 433 299 715 325
rect 433 247 449 299
rect 501 247 513 299
rect 565 273 715 299
rect 767 273 886 325
rect 565 255 886 273
rect 565 247 715 255
rect 433 232 715 247
rect 433 180 449 232
rect 501 180 513 232
rect 565 203 715 232
rect 767 203 886 255
rect 1573 1409 1625 1415
rect 1573 1345 1625 1357
rect 1573 973 1625 1293
rect 1573 909 1625 921
rect 565 185 886 203
rect 565 180 715 185
rect 433 164 715 180
rect 433 112 449 164
rect 501 112 513 164
rect 565 133 715 164
rect 767 133 886 185
rect 565 114 886 133
rect 565 112 715 114
rect 433 62 715 112
rect 767 62 886 114
rect 433 43 886 62
rect 433 -9 715 43
rect 767 21 886 43
tri 886 21 1068 203 sw
rect 1573 21 1625 857
rect 767 -9 1068 21
rect 433 -15 1068 -9
tri 1068 -15 1104 21 sw
rect 433 -17 1104 -15
tri 433 -22 438 -17 ne
rect 438 -21 1104 -17
tri 1104 -21 1110 -15 sw
rect 438 -22 1528 -21
tri 438 -31 447 -22 ne
rect 447 -31 1528 -22
rect 353 -45 405 -39
tri 447 -43 459 -31 ne
rect 459 -43 1528 -31
tri 459 -45 461 -43 ne
rect 461 -45 1528 -43
tri 461 -95 511 -45 ne
rect 511 -95 1528 -45
tri 511 -101 517 -95 ne
rect 517 -101 1528 -95
rect 1573 -43 1625 -31
rect 1573 -101 1625 -95
tri 517 -313 729 -101 ne
rect 729 -313 1528 -101
rect 1246 -378 1528 -313
rect 1915 -326 1967 1475
rect 1995 1505 2346 4959
rect 1995 -193 2268 1505
tri 2268 1427 2346 1505 nw
tri 2268 -193 2348 -113 sw
rect 1995 -293 2348 -193
tri 1995 -305 2007 -293 ne
rect 2007 -305 2348 -293
tri 1967 -326 1988 -305 sw
tri 2007 -326 2028 -305 ne
rect 1915 -327 1988 -326
tri 1915 -338 1926 -327 ne
rect 1926 -338 1988 -327
tri 1988 -338 2000 -326 sw
tri 1926 -360 1948 -338 ne
rect 1948 -378 2000 -338
rect 2028 -378 2348 -305
use L1M1_CDNS_524688791851292  L1M1_CDNS_524688791851292_0
timestamp 1707688321
transform 1 0 795 0 1 1044
box -12 -6 910 184
use nfet_CDNS_524688791851296  nfet_CDNS_524688791851296_0
timestamp 1707688321
transform 1 0 383 0 1 2475
box -79 -26 259 2026
use nfet_CDNS_524688791851296  nfet_CDNS_524688791851296_1
timestamp 1707688321
transform 1 0 1311 0 1 2475
box -79 -26 259 2026
use nfet_CDNS_524688791851296  nfet_CDNS_524688791851296_2
timestamp 1707688321
transform 1 0 147 0 1 2475
box -79 -26 259 2026
use nfet_CDNS_524688791851296  nfet_CDNS_524688791851296_3
timestamp 1707688321
transform 1 0 619 0 1 2475
box -79 -26 259 2026
use nfet_CDNS_524688791851297  nfet_CDNS_524688791851297_0
timestamp 1707688321
transform -1 0 591 0 1 797
box -82 -26 538 626
use nfet_CDNS_524688791851298  nfet_CDNS_524688791851298_0
timestamp 1707688321
transform -1 0 591 0 1 31
box -82 -26 378 626
use nfet_CDNS_524688791851298  nfet_CDNS_524688791851298_1
timestamp 1707688321
transform -1 0 591 0 -1 2235
box -82 -26 378 626
use nfet_CDNS_524688791851299  nfet_CDNS_524688791851299_0
timestamp 1707688321
transform 1 0 119 0 -1 2235
box -82 -26 202 626
use nfet_CDNS_524688791851299  nfet_CDNS_524688791851299_1
timestamp 1707688321
transform 1 0 119 0 1 31
box -82 -26 202 626
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_0
timestamp 1707688321
transform -1 0 1305 0 1 205
box -119 -66 375 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_1
timestamp 1707688321
transform -1 0 1305 0 -1 2061
box -119 -66 375 666
use pfet_CDNS_524688791851300  pfet_CDNS_524688791851300_0
timestamp 1707688321
transform -1 0 1561 0 1 205
box -119 -66 319 666
use pfet_CDNS_524688791851300  pfet_CDNS_524688791851300_1
timestamp 1707688321
transform -1 0 1561 0 -1 2061
box -119 -66 319 666
use pfet_CDNS_524688791851301  pfet_CDNS_524688791851301_0
timestamp 1707688321
transform -1 0 -339 0 1 3281
box -119 -66 219 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_0
timestamp 1707688321
transform -1 0 -764 0 1 3641
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_1
timestamp 1707688321
transform -1 0 -920 0 1 3641
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_2
timestamp 1707688321
transform -1 0 -963 0 1 4107
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_3
timestamp 1707688321
transform -1 0 -1076 0 1 3641
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_4
timestamp 1707688321
transform -1 0 -495 0 1 4107
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_5
timestamp 1707688321
transform -1 0 -807 0 1 4107
box -122 -66 222 366
use pfet_CDNS_524688791851303  pfet_CDNS_524688791851303_6
timestamp 1707688321
transform -1 0 -651 0 1 4107
box -122 -66 222 366
use pfet_CDNS_524688791851304  pfet_CDNS_524688791851304_0
timestamp 1707688321
transform -1 0 -339 0 1 4107
box -119 -66 222 366
use pfet_CDNS_524688791851304  pfet_CDNS_524688791851304_1
timestamp 1707688321
transform -1 0 -339 0 1 3641
box -119 -66 222 366
use pfet_CDNS_524688791851305  pfet_CDNS_524688791851305_0
timestamp 1707688321
transform -1 0 -1232 0 1 3641
box -122 -66 519 366
use pfet_CDNS_524688791851306  pfet_CDNS_524688791851306_0
timestamp 1707688321
transform -1 0 -495 0 1 3641
box -122 -66 219 366
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 1 -890 -1 0 4573
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 0 1 -734 -1 0 4573
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform 0 1 -578 -1 0 4573
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform 0 1 -422 -1 0 4573
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1707688321
transform 0 1 -1046 -1 0 4573
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 1394 -1 0 1429
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 -1020 -1 0 3573
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 1 1394 1 0 837
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 1076 -1 0 1429
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1707688321
transform 0 1 1076 1 0 837
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1707688321
transform 0 -1 405 -1 0 641
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_0
timestamp 1707688321
transform 1 0 383 0 1 2377
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_0
timestamp 1707688321
transform 0 -1 1612 -1 0 719
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_1
timestamp 1707688321
transform 0 1 -993 -1 0 3678
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_2
timestamp 1707688321
transform 0 1 -1055 -1 0 4589
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_3
timestamp 1707688321
transform 0 1 -743 -1 0 4589
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_4
timestamp 1707688321
transform -1 0 1327 0 1 504
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_5
timestamp 1707688321
transform -1 0 1327 0 -1 1762
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_6
timestamp 1707688321
transform -1 0 431 0 -1 1485
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_7
timestamp 1707688321
transform 0 -1 1612 1 0 1547
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851294  sky130_fd_io__sio_tk_em1o_CDNS_524688791851294_0
timestamp 1707688321
transform -1 0 -1647 0 1 4186
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1707688321
transform 0 -1 405 -1 0 7
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1707688321
transform 0 -1 325 -1 0 7
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_0
timestamp 1707688321
transform 0 -1 -756 -1 0 4457
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_1
timestamp 1707688321
transform 0 -1 -947 -1 0 3848
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_2
timestamp 1707688321
transform 0 -1 -1068 -1 0 4457
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_3
timestamp 1707688321
transform 0 -1 1356 -1 0 2138
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_4
timestamp 1707688321
transform 0 -1 1044 -1 0 2103
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_5
timestamp 1707688321
transform 0 -1 1200 -1 0 808
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_6
timestamp 1707688321
transform 0 -1 -600 -1 0 3699
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_7
timestamp 1707688321
transform -1 0 625 0 -1 1485
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_8
timestamp 1707688321
transform -1 0 170 0 -1 1485
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_9
timestamp 1707688321
transform 0 -1 1200 1 0 1458
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_10
timestamp 1707688321
transform 0 -1 1078 1 0 128
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_11
timestamp 1707688321
transform 0 -1 1356 1 0 128
box 0 0 1 1
use TPL1_CDNS_524688791851290  TPL1_CDNS_524688791851290_0
timestamp 1707688321
transform 1 0 765 0 1 990
box -26 -26 1128 312
use TPL1_CDNS_524688791851291  TPL1_CDNS_524688791851291_0
timestamp 1707688321
transform 0 -1 1164 -1 0 4570
box -26 -26 2216 244
<< labels >>
flabel comment s -12 1337 -12 1337 0 FreeSans 100 90 0 0 li_jumper_ok
flabel comment s -1046 4886 -1046 4886 3 FreeSans 400 270 0 0 vpwr_ka
flabel comment s -1899 2542 -1899 2542 3 FreeSans 400 90 0 0 vcc_io
flabel comment s -1899 4886 -1899 4886 3 FreeSans 400 270 0 0 vcc_io
flabel comment s -1338 4888 -1338 4888 3 FreeSans 400 270 0 0 vnb
flabel metal1 s -115 -100 -63 -73 0 FreeSans 200 0 0 0 nbias
port 5 nsew
flabel metal1 s 273 -137 325 -103 0 FreeSans 200 90 0 0 ie_diff_sel_h_n
port 3 nsew
flabel metal1 s 1573 -101 1625 -84 3 FreeSans 200 90 0 0 vinref
port 4 nsew
flabel metal1 s 353 -137 405 -103 0 FreeSans 200 0 0 0 ie_diff_sel_h
port 2 nsew
flabel metal2 s -103 86 210 119 0 FreeSans 200 0 0 0 vcc_ioq
port 6 nsew
flabel metal2 s 1948 -378 2000 -342 0 FreeSans 200 0 0 0 ng_ctl
port 7 nsew
flabel metal2 s 538 -15 858 11 3 FreeSans 200 90 0 0 vgnd
port 8 nsew
<< properties >>
string GDS_END 86494828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86378102
string path -36.650 80.575 -36.650 77.325 
<< end >>
