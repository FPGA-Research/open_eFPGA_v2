magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 98 157 638 203
rect 1 21 638 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 174 47 204 177
rect 258 47 288 177
rect 446 47 476 177
rect 530 47 560 177
<< scpmoshvt >>
rect 79 369 109 497
rect 267 309 297 497
rect 351 309 381 497
rect 446 297 476 497
rect 530 297 560 497
<< ndiff >>
rect 124 131 174 177
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 174 131
rect 109 55 125 89
rect 159 55 174 89
rect 109 47 174 55
rect 204 124 258 177
rect 204 90 214 124
rect 248 90 258 124
rect 204 47 258 90
rect 288 93 340 177
rect 288 59 298 93
rect 332 59 340 93
rect 288 47 340 59
rect 394 124 446 177
rect 394 90 402 124
rect 436 90 446 124
rect 394 47 446 90
rect 476 169 530 177
rect 476 135 486 169
rect 520 135 530 169
rect 476 47 530 135
rect 560 101 612 177
rect 560 67 570 101
rect 604 67 612 101
rect 560 47 612 67
<< pdiff >>
rect 27 450 79 497
rect 27 416 35 450
rect 69 416 79 450
rect 27 369 79 416
rect 109 485 161 497
rect 109 451 119 485
rect 153 451 161 485
rect 109 369 161 451
rect 215 477 267 497
rect 215 443 223 477
rect 257 443 267 477
rect 215 409 267 443
rect 215 375 223 409
rect 257 375 267 409
rect 215 309 267 375
rect 297 489 351 497
rect 297 455 307 489
rect 341 455 351 489
rect 297 421 351 455
rect 297 387 307 421
rect 341 387 351 421
rect 297 309 351 387
rect 381 477 446 497
rect 381 443 397 477
rect 431 443 446 477
rect 381 409 446 443
rect 381 375 397 409
rect 431 375 446 409
rect 381 309 446 375
rect 396 297 446 309
rect 476 407 530 497
rect 476 373 486 407
rect 520 373 530 407
rect 476 339 530 373
rect 476 305 486 339
rect 520 305 530 339
rect 476 297 530 305
rect 560 477 612 497
rect 560 443 570 477
rect 604 443 612 477
rect 560 409 612 443
rect 560 375 570 409
rect 604 375 612 409
rect 560 297 612 375
<< ndiffc >>
rect 35 72 69 106
rect 125 55 159 89
rect 214 90 248 124
rect 298 59 332 93
rect 402 90 436 124
rect 486 135 520 169
rect 570 67 604 101
<< pdiffc >>
rect 35 416 69 450
rect 119 451 153 485
rect 223 443 257 477
rect 223 375 257 409
rect 307 455 341 489
rect 307 387 341 421
rect 397 443 431 477
rect 397 375 431 409
rect 486 373 520 407
rect 486 305 520 339
rect 570 443 604 477
rect 570 375 604 409
<< poly >>
rect 79 497 109 523
rect 267 497 297 523
rect 351 497 381 523
rect 446 497 476 523
rect 530 497 560 523
rect 79 265 109 369
rect 22 249 109 265
rect 267 294 297 309
rect 351 294 381 309
rect 267 265 381 294
rect 446 265 476 297
rect 530 265 560 297
rect 267 264 385 265
rect 22 215 32 249
rect 66 222 109 249
rect 331 249 385 264
rect 66 215 288 222
rect 22 199 288 215
rect 331 215 341 249
rect 375 215 385 249
rect 331 199 385 215
rect 446 249 623 265
rect 446 215 579 249
rect 613 215 623 249
rect 446 199 623 215
rect 79 192 288 199
rect 79 131 109 192
rect 174 177 204 192
rect 258 177 288 192
rect 446 177 476 199
rect 530 177 560 199
rect 79 21 109 47
rect 174 21 204 47
rect 258 21 288 47
rect 446 21 476 47
rect 530 21 560 47
<< polycont >>
rect 32 215 66 249
rect 341 215 375 249
rect 579 215 613 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 450 69 493
rect 17 416 35 450
rect 103 485 175 527
rect 103 451 119 485
rect 153 451 175 485
rect 103 425 175 451
rect 209 477 257 493
rect 209 443 223 477
rect 17 391 69 416
rect 209 409 257 443
rect 17 357 175 391
rect 17 249 66 323
rect 17 215 32 249
rect 17 199 66 215
rect 100 265 175 357
rect 209 375 223 409
rect 291 489 357 527
rect 291 455 307 489
rect 341 455 357 489
rect 291 421 357 455
rect 291 387 307 421
rect 341 387 357 421
rect 291 379 357 387
rect 397 477 627 493
rect 431 459 570 477
rect 397 409 431 443
rect 604 443 627 477
rect 209 345 257 375
rect 397 345 431 375
rect 209 311 431 345
rect 470 407 536 425
rect 470 373 486 407
rect 520 373 536 407
rect 470 339 536 373
rect 570 409 627 443
rect 604 375 627 409
rect 570 357 627 375
rect 470 305 486 339
rect 520 305 536 339
rect 100 249 436 265
rect 100 215 341 249
rect 375 215 436 249
rect 100 199 436 215
rect 100 165 175 199
rect 470 169 536 305
rect 17 131 175 165
rect 209 131 436 165
rect 17 106 69 131
rect 17 72 35 106
rect 209 124 248 131
rect 17 51 69 72
rect 103 89 175 97
rect 103 55 125 89
rect 159 55 175 89
rect 103 17 175 55
rect 209 90 214 124
rect 388 124 436 131
rect 209 51 248 90
rect 282 93 354 97
rect 282 59 298 93
rect 332 59 354 93
rect 282 17 354 59
rect 388 90 402 124
rect 470 135 486 169
rect 520 135 536 169
rect 570 249 627 323
rect 570 215 579 249
rect 613 215 627 249
rect 570 153 627 215
rect 470 119 536 135
rect 388 85 436 90
rect 570 101 627 119
rect 388 67 570 85
rect 604 67 627 101
rect 388 51 627 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 582 153 616 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 582 289 616 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 490 153 524 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 490 289 524 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 490 357 524 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 TE
port 2 nsew signal input
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 einvp_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 2030880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2024692
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
