magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 1072 29 1130 325
rect 2202 29 2224 325
rect 3231 29 3763 667
rect 0 -77 3817 29
<< pwell >>
rect 3234 1165 3730 1251
<< psubdiff >>
rect 3260 1191 3284 1225
rect 3318 1191 3357 1225
rect 3391 1191 3430 1225
rect 3464 1191 3502 1225
rect 3536 1191 3574 1225
rect 3608 1191 3646 1225
rect 3680 1191 3704 1225
<< nsubdiff >>
rect 3298 607 3332 631
rect 3298 539 3332 573
rect 3298 470 3332 505
rect 3298 401 3332 436
rect 3260 367 3298 377
rect 3260 343 3332 367
rect 36 -41 60 -7
rect 94 -41 130 -7
rect 164 -41 200 -7
rect 234 -41 270 -7
rect 304 -41 340 -7
rect 374 -41 410 -7
rect 444 -41 480 -7
rect 514 -41 549 -7
rect 583 -41 618 -7
rect 652 -41 687 -7
rect 721 -41 756 -7
rect 790 -41 825 -7
rect 859 -41 894 -7
rect 928 -41 963 -7
rect 997 -41 1032 -7
rect 1066 -41 1101 -7
rect 1135 -41 1170 -7
rect 1204 -41 1239 -7
rect 1273 -41 1308 -7
rect 1342 -41 1377 -7
rect 1411 -41 1446 -7
rect 1480 -41 1515 -7
rect 1549 -41 1584 -7
rect 1618 -41 1653 -7
rect 1687 -41 1722 -7
rect 1756 -41 1791 -7
rect 1825 -41 1860 -7
rect 1894 -41 1929 -7
rect 1963 -41 1998 -7
rect 2032 -41 2067 -7
rect 2101 -41 2136 -7
rect 2170 -41 2205 -7
rect 2239 -41 2274 -7
rect 2308 -41 2343 -7
rect 2377 -41 2412 -7
rect 2446 -41 2481 -7
rect 2515 -41 2550 -7
rect 2584 -41 2619 -7
rect 2653 -41 2688 -7
rect 2722 -41 2757 -7
rect 2791 -41 2826 -7
rect 2860 -41 2895 -7
rect 2929 -41 2964 -7
rect 2998 -41 3033 -7
rect 3067 -41 3102 -7
rect 3136 -41 3171 -7
rect 3205 -41 3240 -7
rect 3274 -41 3309 -7
rect 3343 -41 3378 -7
rect 3412 -41 3447 -7
rect 3481 -41 3516 -7
rect 3550 -41 3585 -7
rect 3619 -41 3654 -7
rect 3688 -41 3723 -7
rect 3757 -41 3781 -7
<< psubdiffcont >>
rect 3284 1191 3318 1225
rect 3357 1191 3391 1225
rect 3430 1191 3464 1225
rect 3502 1191 3536 1225
rect 3574 1191 3608 1225
rect 3646 1191 3680 1225
<< nsubdiffcont >>
rect 3298 573 3332 607
rect 3298 505 3332 539
rect 3298 436 3332 470
rect 3298 367 3332 401
rect 60 -41 94 -7
rect 130 -41 164 -7
rect 200 -41 234 -7
rect 270 -41 304 -7
rect 340 -41 374 -7
rect 410 -41 444 -7
rect 480 -41 514 -7
rect 549 -41 583 -7
rect 618 -41 652 -7
rect 687 -41 721 -7
rect 756 -41 790 -7
rect 825 -41 859 -7
rect 894 -41 928 -7
rect 963 -41 997 -7
rect 1032 -41 1066 -7
rect 1101 -41 1135 -7
rect 1170 -41 1204 -7
rect 1239 -41 1273 -7
rect 1308 -41 1342 -7
rect 1377 -41 1411 -7
rect 1446 -41 1480 -7
rect 1515 -41 1549 -7
rect 1584 -41 1618 -7
rect 1653 -41 1687 -7
rect 1722 -41 1756 -7
rect 1791 -41 1825 -7
rect 1860 -41 1894 -7
rect 1929 -41 1963 -7
rect 1998 -41 2032 -7
rect 2067 -41 2101 -7
rect 2136 -41 2170 -7
rect 2205 -41 2239 -7
rect 2274 -41 2308 -7
rect 2343 -41 2377 -7
rect 2412 -41 2446 -7
rect 2481 -41 2515 -7
rect 2550 -41 2584 -7
rect 2619 -41 2653 -7
rect 2688 -41 2722 -7
rect 2757 -41 2791 -7
rect 2826 -41 2860 -7
rect 2895 -41 2929 -7
rect 2964 -41 2998 -7
rect 3033 -41 3067 -7
rect 3102 -41 3136 -7
rect 3171 -41 3205 -7
rect 3240 -41 3274 -7
rect 3309 -41 3343 -7
rect 3378 -41 3412 -7
rect 3447 -41 3481 -7
rect 3516 -41 3550 -7
rect 3585 -41 3619 -7
rect 3654 -41 3688 -7
rect 3723 -41 3757 -7
<< poly >>
rect 3247 789 3651 825
rect 3247 751 3457 789
rect 3247 717 3271 751
rect 3305 717 3339 751
rect 3373 717 3407 751
rect 3441 717 3457 751
rect 3247 701 3457 717
rect 1068 236 1134 243
rect 3292 236 3358 239
rect 1062 227 1140 236
rect 1062 200 1084 227
rect 1068 193 1084 200
rect 1118 200 1140 227
rect 3286 223 3358 236
rect 3286 200 3308 223
rect 1118 193 1134 200
rect 1068 159 1134 193
rect 1068 144 1084 159
rect 1061 125 1084 144
rect 1118 144 1134 159
rect 3292 189 3308 200
rect 3342 189 3358 223
rect 3292 155 3358 189
rect 3292 144 3308 155
rect 1118 125 1140 144
rect 1061 108 1140 125
rect 3286 121 3308 144
rect 3342 121 3358 155
rect 3286 108 3358 121
rect 3292 105 3358 108
rect 3574 81 3674 87
rect 3574 65 3708 81
rect 3574 31 3590 65
rect 3624 31 3658 65
rect 3692 31 3708 65
rect 3574 15 3708 31
<< polycont >>
rect 3271 717 3305 751
rect 3339 717 3373 751
rect 3407 717 3441 751
rect 1084 193 1118 227
rect 1084 125 1118 159
rect 3308 189 3342 223
rect 3308 121 3342 155
rect 3590 31 3624 65
rect 3658 31 3692 65
<< locali >>
rect 3252 1191 3284 1225
rect 3318 1191 3357 1225
rect 3391 1191 3430 1225
rect 3464 1191 3502 1225
rect 3536 1191 3574 1225
rect 3608 1191 3646 1225
rect 3680 1191 3696 1225
rect 3202 1085 3236 1123
rect 3202 1013 3236 1051
rect 3386 1085 3420 1123
rect 3386 1013 3420 1051
rect 3570 1085 3604 1123
rect 3570 1013 3604 1051
rect 3294 819 3328 853
rect 3478 819 3512 853
rect 3662 819 3696 853
rect 3294 785 3297 819
rect 3331 785 3369 819
rect 3403 785 3441 819
rect 3475 785 3513 819
rect 3547 785 3585 819
rect 3619 785 3657 819
rect 3691 785 3696 819
rect 3255 717 3271 751
rect 3305 717 3339 751
rect 3373 717 3407 751
rect 3441 717 3563 751
rect 3447 676 3563 717
rect 3298 607 3332 631
rect 3298 539 3332 573
rect 3298 470 3332 505
rect 3298 401 3332 436
rect 3252 367 3298 377
rect 3252 343 3332 367
rect 982 247 1050 281
rect 1016 97 1050 247
rect 1084 237 1118 275
rect 1084 159 1118 193
rect 1084 109 1118 125
rect 1152 247 1220 281
rect 2226 247 2319 281
rect 980 63 1050 97
rect 1152 97 1186 247
rect 2226 189 2260 247
rect 3447 239 3549 676
rect 3685 607 3719 645
rect 3685 535 3719 573
rect 3685 272 3719 310
rect 2170 155 2260 189
rect 2226 97 2260 155
rect 3308 223 3563 239
rect 3342 189 3563 223
rect 3308 155 3563 189
rect 3342 121 3563 155
rect 3308 105 3563 121
rect 1152 63 1222 97
rect 2226 63 2316 97
rect 3574 31 3590 65
rect 3624 31 3658 65
rect 3692 31 3708 65
rect 36 -41 47 -7
rect 94 -41 121 -7
rect 164 -41 195 -7
rect 234 -41 269 -7
rect 304 -41 340 -7
rect 377 -41 410 -7
rect 451 -41 480 -7
rect 525 -41 549 -7
rect 599 -41 618 -7
rect 673 -41 687 -7
rect 747 -41 756 -7
rect 821 -41 825 -7
rect 859 -41 861 -7
rect 928 -41 935 -7
rect 997 -41 1009 -7
rect 1066 -41 1083 -7
rect 1135 -41 1157 -7
rect 1204 -41 1231 -7
rect 1273 -41 1305 -7
rect 1342 -41 1377 -7
rect 1412 -41 1446 -7
rect 1485 -41 1515 -7
rect 1558 -41 1584 -7
rect 1631 -41 1653 -7
rect 1704 -41 1722 -7
rect 1777 -41 1791 -7
rect 1850 -41 1860 -7
rect 1923 -41 1929 -7
rect 1996 -41 1998 -7
rect 2032 -41 2035 -7
rect 2101 -41 2108 -7
rect 2170 -41 2181 -7
rect 2239 -41 2254 -7
rect 2308 -41 2327 -7
rect 2377 -41 2400 -7
rect 2446 -41 2473 -7
rect 2515 -41 2546 -7
rect 2584 -41 2619 -7
rect 2653 -41 2688 -7
rect 2726 -41 2757 -7
rect 2799 -41 2826 -7
rect 2872 -41 2895 -7
rect 2945 -41 2964 -7
rect 3018 -41 3033 -7
rect 3091 -41 3102 -7
rect 3164 -41 3171 -7
rect 3237 -41 3240 -7
rect 3274 -41 3276 -7
rect 3343 -41 3349 -7
rect 3412 -41 3422 -7
rect 3481 -41 3495 -7
rect 3550 -41 3568 -7
rect 3619 -41 3641 -7
rect 3688 -41 3714 -7
rect 3757 -41 3781 -7
<< viali >>
rect 3202 1123 3236 1157
rect 3202 1051 3236 1085
rect 3202 979 3236 1013
rect 3386 1123 3420 1157
rect 3386 1051 3420 1085
rect 3386 979 3420 1013
rect 3570 1123 3604 1157
rect 3570 1051 3604 1085
rect 3570 979 3604 1013
rect 3297 785 3331 819
rect 3369 785 3403 819
rect 3441 785 3475 819
rect 3513 785 3547 819
rect 3585 785 3619 819
rect 3657 785 3691 819
rect 1084 275 1118 309
rect 1084 227 1118 237
rect 1084 203 1118 227
rect 3685 645 3719 679
rect 3685 573 3719 607
rect 3685 501 3719 535
rect 3685 310 3719 344
rect 3685 238 3719 272
rect 47 -41 60 -7
rect 60 -41 81 -7
rect 121 -41 130 -7
rect 130 -41 155 -7
rect 195 -41 200 -7
rect 200 -41 229 -7
rect 269 -41 270 -7
rect 270 -41 303 -7
rect 343 -41 374 -7
rect 374 -41 377 -7
rect 417 -41 444 -7
rect 444 -41 451 -7
rect 491 -41 514 -7
rect 514 -41 525 -7
rect 565 -41 583 -7
rect 583 -41 599 -7
rect 639 -41 652 -7
rect 652 -41 673 -7
rect 713 -41 721 -7
rect 721 -41 747 -7
rect 787 -41 790 -7
rect 790 -41 821 -7
rect 861 -41 894 -7
rect 894 -41 895 -7
rect 935 -41 963 -7
rect 963 -41 969 -7
rect 1009 -41 1032 -7
rect 1032 -41 1043 -7
rect 1083 -41 1101 -7
rect 1101 -41 1117 -7
rect 1157 -41 1170 -7
rect 1170 -41 1191 -7
rect 1231 -41 1239 -7
rect 1239 -41 1265 -7
rect 1305 -41 1308 -7
rect 1308 -41 1339 -7
rect 1378 -41 1411 -7
rect 1411 -41 1412 -7
rect 1451 -41 1480 -7
rect 1480 -41 1485 -7
rect 1524 -41 1549 -7
rect 1549 -41 1558 -7
rect 1597 -41 1618 -7
rect 1618 -41 1631 -7
rect 1670 -41 1687 -7
rect 1687 -41 1704 -7
rect 1743 -41 1756 -7
rect 1756 -41 1777 -7
rect 1816 -41 1825 -7
rect 1825 -41 1850 -7
rect 1889 -41 1894 -7
rect 1894 -41 1923 -7
rect 1962 -41 1963 -7
rect 1963 -41 1996 -7
rect 2035 -41 2067 -7
rect 2067 -41 2069 -7
rect 2108 -41 2136 -7
rect 2136 -41 2142 -7
rect 2181 -41 2205 -7
rect 2205 -41 2215 -7
rect 2254 -41 2274 -7
rect 2274 -41 2288 -7
rect 2327 -41 2343 -7
rect 2343 -41 2361 -7
rect 2400 -41 2412 -7
rect 2412 -41 2434 -7
rect 2473 -41 2481 -7
rect 2481 -41 2507 -7
rect 2546 -41 2550 -7
rect 2550 -41 2580 -7
rect 2619 -41 2653 -7
rect 2692 -41 2722 -7
rect 2722 -41 2726 -7
rect 2765 -41 2791 -7
rect 2791 -41 2799 -7
rect 2838 -41 2860 -7
rect 2860 -41 2872 -7
rect 2911 -41 2929 -7
rect 2929 -41 2945 -7
rect 2984 -41 2998 -7
rect 2998 -41 3018 -7
rect 3057 -41 3067 -7
rect 3067 -41 3091 -7
rect 3130 -41 3136 -7
rect 3136 -41 3164 -7
rect 3203 -41 3205 -7
rect 3205 -41 3237 -7
rect 3276 -41 3309 -7
rect 3309 -41 3310 -7
rect 3349 -41 3378 -7
rect 3378 -41 3383 -7
rect 3422 -41 3447 -7
rect 3447 -41 3456 -7
rect 3495 -41 3516 -7
rect 3516 -41 3529 -7
rect 3568 -41 3585 -7
rect 3585 -41 3602 -7
rect 3641 -41 3654 -7
rect 3654 -41 3675 -7
rect 3714 -41 3723 -7
rect 3723 -41 3748 -7
<< metal1 >>
rect 3196 1157 3817 1169
rect 3196 1123 3202 1157
rect 3236 1123 3386 1157
rect 3420 1123 3570 1157
rect 3604 1123 3817 1157
rect 3196 1085 3817 1123
rect 3196 1051 3202 1085
rect 3236 1051 3386 1085
rect 3420 1051 3570 1085
rect 3604 1051 3817 1085
rect 3196 1013 3817 1051
rect 3196 979 3202 1013
rect 3236 979 3386 1013
rect 3420 979 3570 1013
rect 3604 979 3817 1013
rect 3196 967 3817 979
rect 2783 773 2789 825
rect 2841 773 2853 825
rect 2905 819 3703 825
rect 2905 785 3297 819
rect 3331 785 3369 819
rect 3403 785 3441 819
rect 3475 785 3513 819
rect 3547 785 3585 819
rect 3619 785 3657 819
rect 3691 785 3703 819
rect 2905 773 3703 785
rect 0 679 3745 691
rect 0 645 3685 679
rect 3719 645 3745 679
rect 0 607 3745 645
rect 0 573 3685 607
rect 3719 573 3745 607
rect 0 535 3745 573
rect 0 501 3685 535
rect 3719 501 3745 535
rect 0 489 3745 501
tri 3693 457 3725 489 ne
rect 3679 344 3725 356
rect 1072 309 1130 315
tri 3677 310 3679 312 se
rect 3679 310 3685 344
rect 3719 310 3725 344
rect 83 226 1005 287
rect 1072 275 1084 309
rect 1118 275 1130 309
tri 3654 287 3677 310 se
rect 3677 287 3725 310
rect 1072 237 1130 275
rect 1072 203 1084 237
rect 1118 203 1130 237
rect 1206 272 3725 287
rect 1206 238 3685 272
rect 3719 238 3725 272
rect 1206 226 3725 238
rect 1072 197 1130 203
tri 994 169 1020 195 sw
tri 1182 169 1208 195 se
rect 144 149 2202 169
tri 144 146 147 149 ne
rect 147 146 2202 149
rect 2282 146 2789 198
rect 2841 146 2853 198
rect 2905 146 3364 198
tri 147 131 162 146 ne
rect 162 131 2202 146
rect 83 39 2911 103
rect 35 -7 3774 9
rect 35 -41 47 -7
rect 81 -41 121 -7
rect 155 -41 195 -7
rect 229 -41 269 -7
rect 303 -41 343 -7
rect 377 -41 417 -7
rect 451 -41 491 -7
rect 525 -41 565 -7
rect 599 -41 639 -7
rect 673 -41 713 -7
rect 747 -41 787 -7
rect 821 -41 861 -7
rect 895 -41 935 -7
rect 969 -41 1009 -7
rect 1043 -41 1083 -7
rect 1117 -41 1157 -7
rect 1191 -41 1231 -7
rect 1265 -41 1305 -7
rect 1339 -41 1378 -7
rect 1412 -41 1451 -7
rect 1485 -41 1524 -7
rect 1558 -41 1597 -7
rect 1631 -41 1670 -7
rect 1704 -41 1743 -7
rect 1777 -41 1816 -7
rect 1850 -41 1889 -7
rect 1923 -41 1962 -7
rect 1996 -41 2035 -7
rect 2069 -41 2108 -7
rect 2142 -41 2181 -7
rect 2215 -41 2254 -7
rect 2288 -41 2327 -7
rect 2361 -41 2400 -7
rect 2434 -41 2473 -7
rect 2507 -41 2546 -7
rect 2580 -41 2619 -7
rect 2653 -41 2692 -7
rect 2726 -41 2765 -7
rect 2799 -41 2838 -7
rect 2872 -41 2911 -7
rect 2945 -41 2984 -7
rect 3018 -41 3057 -7
rect 3091 -41 3130 -7
rect 3164 -41 3203 -7
rect 3237 -41 3276 -7
rect 3310 -41 3349 -7
rect 3383 -41 3422 -7
rect 3456 -41 3495 -7
rect 3529 -41 3568 -7
rect 3602 -41 3641 -7
rect 3675 -41 3714 -7
rect 3748 -41 3774 -7
rect 35 -55 3774 -41
<< via1 >>
rect 2789 773 2841 825
rect 2853 773 2905 825
rect 2789 146 2841 198
rect 2853 146 2905 198
<< metal2 >>
rect 2783 773 2789 825
rect 2841 773 2853 825
rect 2905 773 2911 825
rect 2783 198 2911 773
rect 2783 146 2789 198
rect 2841 146 2853 198
rect 2905 146 2911 198
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 1 0 1084 0 1 203
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 3719 1 0 238
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 1 3685 -1 0 679
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 1 3202 -1 0 1157
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 1 3570 -1 0 1157
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 1 3386 -1 0 1157
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1707688321
transform -1 0 982 0 1 155
box -12 -6 838 40
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 1 0 3297 0 -1 819
box 0 0 1 1
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1707688321
transform -1 0 993 0 1 247
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1707688321
transform -1 0 993 0 1 63
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_2
timestamp 1707688321
transform 1 0 1218 0 1 247
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_3
timestamp 1707688321
transform 1 0 1218 0 1 63
box -12 -6 910 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1707688321
transform 1 0 2294 0 -1 189
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_1
timestamp 1707688321
transform 1 0 1220 0 1 155
box -12 -6 982 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 2911 0 1 146
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 1 0 2783 0 -1 825
box 0 0 1 1
use nfet_CDNS_524688791851199  nfet_CDNS_524688791851199_0
timestamp 1707688321
transform 1 0 3247 0 -1 1051
box -79 -26 483 226
use pfet_CDNS_524688791851196  pfet_CDNS_524688791851196_0
timestamp 1707688321
transform 0 1 36 1 0 108
box -89 -36 217 1036
use pfet_CDNS_524688791851197  pfet_CDNS_524688791851197_0
timestamp 1707688321
transform 0 -1 3260 -1 0 236
box -89 -36 217 1036
use pfet_CDNS_524688791851197  pfet_CDNS_524688791851197_1
timestamp 1707688321
transform 0 -1 2166 -1 0 236
box -89 -36 217 1036
use pfet_CDNS_524688791851198  pfet_CDNS_524688791851198_0
timestamp 1707688321
transform 1 0 3574 0 -1 713
box -89 -36 189 636
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 3708 -1 0 81
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform -1 0 3358 0 -1 239
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform -1 0 1134 0 -1 243
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 3255 -1 0 767
box 0 0 1 1
<< labels >>
flabel comment s 3623 90 3623 90 0 FreeSans 200 180 0 0 ctl_in_n
flabel comment s 3343 283 3343 283 0 FreeSans 200 180 0 0 out
flabel metal1 s 1084 243 1118 275 0 FreeSans 200 0 0 0 ctl_in
port 4 nsew
flabel metal1 s 3685 645 3719 678 0 FreeSans 400 0 0 0 vpwr
port 2 nsew
flabel metal1 s 3202 1123 3236 1157 0 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel locali s 2137 173 2137 173 0 FreeSans 400 0 0 0 n<0>
flabel locali s 3658 31 3692 65 0 FreeSans 400 0 0 0 ctl_in_n
port 5 nsew
flabel locali s 3431 152 3465 186 0 FreeSans 600 0 0 0 din
port 6 nsew
flabel metal2 s 2832 785 2862 815 0 FreeSans 400 0 0 0 out
port 7 nsew
<< properties >>
string GDS_END 85810432
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85797340
string path 0.250 -0.600 95.175 -0.600 
<< end >>
