magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 -36 92 2036
<< pdiff >>
rect 0 1950 56 2000
rect 0 1916 11 1950
rect 45 1916 56 1950
rect 0 1882 56 1916
rect 0 1848 11 1882
rect 45 1848 56 1882
rect 0 1814 56 1848
rect 0 1780 11 1814
rect 45 1780 56 1814
rect 0 1746 56 1780
rect 0 1712 11 1746
rect 45 1712 56 1746
rect 0 1678 56 1712
rect 0 1644 11 1678
rect 45 1644 56 1678
rect 0 1610 56 1644
rect 0 1576 11 1610
rect 45 1576 56 1610
rect 0 1542 56 1576
rect 0 1508 11 1542
rect 45 1508 56 1542
rect 0 1474 56 1508
rect 0 1440 11 1474
rect 45 1440 56 1474
rect 0 1406 56 1440
rect 0 1372 11 1406
rect 45 1372 56 1406
rect 0 1338 56 1372
rect 0 1304 11 1338
rect 45 1304 56 1338
rect 0 1270 56 1304
rect 0 1236 11 1270
rect 45 1236 56 1270
rect 0 1202 56 1236
rect 0 1168 11 1202
rect 45 1168 56 1202
rect 0 1134 56 1168
rect 0 1100 11 1134
rect 45 1100 56 1134
rect 0 1066 56 1100
rect 0 1032 11 1066
rect 45 1032 56 1066
rect 0 998 56 1032
rect 0 964 11 998
rect 45 964 56 998
rect 0 930 56 964
rect 0 896 11 930
rect 45 896 56 930
rect 0 862 56 896
rect 0 828 11 862
rect 45 828 56 862
rect 0 794 56 828
rect 0 760 11 794
rect 45 760 56 794
rect 0 726 56 760
rect 0 692 11 726
rect 45 692 56 726
rect 0 658 56 692
rect 0 624 11 658
rect 45 624 56 658
rect 0 590 56 624
rect 0 556 11 590
rect 45 556 56 590
rect 0 522 56 556
rect 0 488 11 522
rect 45 488 56 522
rect 0 454 56 488
rect 0 420 11 454
rect 45 420 56 454
rect 0 386 56 420
rect 0 352 11 386
rect 45 352 56 386
rect 0 318 56 352
rect 0 284 11 318
rect 45 284 56 318
rect 0 250 56 284
rect 0 216 11 250
rect 45 216 56 250
rect 0 182 56 216
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< pdiffc >>
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 1950 45 1966
rect 11 1882 45 1916
rect 11 1814 45 1848
rect 11 1746 45 1780
rect 11 1678 45 1712
rect 11 1610 45 1644
rect 11 1542 45 1576
rect 11 1474 45 1508
rect 11 1406 45 1440
rect 11 1338 45 1372
rect 11 1270 45 1304
rect 11 1202 45 1236
rect 11 1134 45 1168
rect 11 1066 45 1100
rect 11 998 45 1032
rect 11 930 45 964
rect 11 862 45 896
rect 11 794 45 828
rect 11 726 45 760
rect 11 658 45 692
rect 11 590 45 624
rect 11 522 45 556
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 90860522
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90858406
<< end >>
