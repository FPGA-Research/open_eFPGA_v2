magic
tech sky130A
timestamp 1707688321
<< properties >>
string GDS_END 68190
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 67866
<< end >>
