magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 106 512 1440 844
rect 3783 -835 4173 213
<< pwell >>
rect 706 274 840 360
rect 738 116 811 274
rect 446 8 708 94
rect 1056 8 1250 94
rect 4325 -419 4411 -387
rect 4591 -389 4677 -127
rect 4325 -492 4569 -419
rect 4325 -521 4411 -492
<< mvpsubdiff >>
rect 732 300 756 334
rect 790 300 814 334
rect 472 34 496 68
rect 530 34 624 68
rect 658 34 682 68
rect 1082 34 1106 68
rect 1140 34 1224 68
rect 4617 -177 4651 -153
rect 4617 -305 4651 -211
rect 4617 -363 4651 -339
rect 4351 -437 4385 -413
rect 4351 -495 4385 -471
<< mvnsubdiff >>
rect 186 736 210 770
rect 244 736 308 770
rect 342 736 406 770
rect 440 736 464 770
rect 838 736 862 770
rect 896 736 939 770
rect 973 736 1016 770
rect 1050 736 1074 770
rect 3915 109 3949 133
rect 3915 11 3949 75
rect 3915 -87 3949 -23
rect 3915 -145 3949 -121
rect 3915 -543 3949 -519
rect 3915 -620 3949 -577
rect 3915 -697 3949 -654
rect 3915 -755 3949 -731
<< mvpsubdiffcont >>
rect 756 300 790 334
rect 496 34 530 68
rect 624 34 658 68
rect 1106 34 1140 68
rect 4617 -211 4651 -177
rect 4617 -339 4651 -305
rect 4351 -471 4385 -437
<< mvnsubdiffcont >>
rect 210 736 244 770
rect 308 736 342 770
rect 406 736 440 770
rect 862 736 896 770
rect 939 736 973 770
rect 1016 736 1050 770
rect 3915 75 3949 109
rect 3915 -23 3949 11
rect 3915 -121 3949 -87
rect 3915 -577 3949 -543
rect 3915 -654 3949 -620
rect 3915 -731 3949 -697
<< poly >>
rect 225 530 345 552
rect 225 496 274 530
rect 308 496 345 530
rect 591 504 711 552
rect 225 462 345 496
rect 225 428 274 462
rect 308 428 345 462
rect 225 252 345 428
rect 454 488 711 504
rect 835 498 955 552
rect 1201 504 1321 552
rect 454 454 470 488
rect 504 454 711 488
rect 454 420 711 454
rect 821 482 955 498
rect 821 448 837 482
rect 871 448 905 482
rect 939 448 955 482
rect 821 432 955 448
rect 454 386 470 420
rect 504 386 711 420
rect 454 370 711 386
rect 511 226 711 370
rect 835 226 955 432
rect 997 488 1321 504
rect 997 454 1013 488
rect 1047 454 1321 488
rect 997 420 1321 454
rect 997 386 1013 420
rect 1047 386 1321 420
rect 997 370 1321 386
rect 1121 226 1321 370
rect 4133 45 4433 94
rect 4133 11 4155 45
rect 4189 11 4223 45
rect 4257 11 4433 45
rect 4133 -26 4433 11
rect 4181 -151 4315 -135
rect 4181 -185 4197 -151
rect 4231 -185 4265 -151
rect 4299 -185 4315 -151
rect 4181 -192 4315 -185
rect 4181 -272 4459 -192
rect 4133 -392 4459 -272
rect 4187 -516 4253 -502
rect 4133 -518 4459 -516
rect 4133 -552 4203 -518
rect 4237 -552 4459 -518
rect 4133 -586 4459 -552
rect 4133 -620 4203 -586
rect 4237 -620 4459 -586
rect 4133 -636 4459 -620
rect 4181 -694 4315 -678
rect 4181 -728 4197 -694
rect 4231 -728 4265 -694
rect 4299 -728 4315 -694
rect 4181 -744 4315 -728
<< polycont >>
rect 274 496 308 530
rect 274 428 308 462
rect 470 454 504 488
rect 837 448 871 482
rect 905 448 939 482
rect 470 386 504 420
rect 1013 454 1047 488
rect 1013 386 1047 420
rect 4155 11 4189 45
rect 4223 11 4257 45
rect 4197 -185 4231 -151
rect 4265 -185 4299 -151
rect 4203 -552 4237 -518
rect 4203 -620 4237 -586
rect 4197 -728 4231 -694
rect 4265 -728 4299 -694
<< locali >>
rect 180 770 464 782
rect 180 736 210 770
rect 244 736 308 770
rect 342 736 406 770
rect 440 736 464 770
rect 180 711 464 736
rect 180 677 241 711
rect 275 677 313 711
rect 347 706 464 711
rect 756 770 1074 782
rect 756 736 862 770
rect 896 736 939 770
rect 973 736 1016 770
rect 1050 736 1074 770
rect 756 706 1074 736
rect 756 703 932 706
rect 180 600 347 677
rect 774 669 812 703
rect 846 669 884 703
rect 918 669 932 703
rect 398 600 436 666
rect 232 496 274 530
rect 308 496 338 530
rect 232 462 338 496
rect 232 448 274 462
rect 308 448 338 462
rect 266 428 274 448
rect 266 414 304 428
rect 398 504 432 600
rect 398 498 504 504
rect 432 464 470 498
rect 398 454 470 464
rect 398 420 504 454
rect 180 160 214 198
rect 180 88 214 126
rect 267 34 301 414
rect 398 386 470 420
rect 398 370 504 386
rect 546 482 580 592
rect 756 580 932 669
rect 1003 600 1088 666
rect 1003 504 1037 600
rect 1122 580 1162 782
rect 1260 711 1366 782
rect 1294 677 1332 711
rect 1260 582 1366 677
rect 1122 548 1190 580
rect 1122 514 1128 548
rect 1162 514 1200 548
rect 1003 488 1060 504
rect 546 448 837 482
rect 871 448 905 482
rect 939 448 955 482
rect 1003 470 1013 488
rect 1047 454 1060 488
rect 546 414 564 448
rect 598 414 636 448
rect 1037 436 1060 454
rect 1003 420 1060 436
rect 398 224 432 370
rect 546 242 580 414
rect 821 368 859 402
rect 893 368 924 402
rect 390 22 432 224
rect 466 176 580 242
rect 620 318 756 334
rect 654 284 692 318
rect 726 300 756 318
rect 790 300 814 334
rect 726 284 814 300
rect 620 68 682 284
rect 472 34 496 68
rect 530 34 624 68
rect 658 34 682 68
rect 722 198 756 230
rect 790 198 828 230
rect 722 160 828 198
rect 722 126 756 160
rect 790 126 828 160
rect 722 88 828 126
rect 722 54 756 88
rect 790 54 828 88
rect 722 28 828 54
rect 890 34 924 368
rect 1003 398 1013 420
rect 1047 386 1060 420
rect 1037 370 1060 386
rect 1003 230 1037 364
rect 1122 230 1156 514
rect 986 28 1037 230
rect 1110 164 1156 230
rect 1190 396 1224 408
rect 1190 324 1224 362
rect 1190 68 1224 290
rect 1082 34 1106 68
rect 1140 34 1224 68
rect 1332 160 1366 198
rect 1332 88 1366 126
rect 3903 109 4085 139
rect 3903 75 3915 109
rect 3949 78 4085 109
rect 4487 105 4525 139
rect 4559 105 4597 139
rect 3949 75 3974 78
rect 3903 44 3974 75
rect 4008 44 4085 78
rect 3903 11 4085 44
rect 3903 -23 3915 11
rect 3949 6 4085 11
rect 3949 -23 3974 6
rect 3903 -28 3974 -23
rect 4008 -28 4085 6
rect 4155 53 4237 87
rect 4155 52 4271 53
rect 4155 45 4651 52
rect 4189 11 4223 45
rect 4257 18 4651 45
rect 4257 15 4271 18
rect 4155 -19 4237 11
rect 3903 -87 3979 -28
rect 4461 -79 4663 -71
rect 3903 -121 3915 -87
rect 3949 -121 3979 -87
rect 4019 -113 4187 -79
rect 4221 -113 4663 -79
rect 4019 -117 4085 -113
rect 3903 -145 3979 -121
rect 4181 -151 4315 -113
rect 4181 -185 4187 -151
rect 4231 -185 4265 -151
rect 4299 -185 4315 -151
rect 4443 -227 4509 -147
rect 4093 -245 4509 -227
rect 4093 -261 4237 -245
rect 4203 -279 4237 -261
rect 4271 -261 4509 -245
rect 4617 -177 4651 -153
rect 4203 -317 4271 -279
rect 4617 -301 4651 -211
rect 3903 -455 3982 -437
rect 4016 -455 4105 -437
rect 3903 -493 4105 -455
rect 3903 -527 3982 -493
rect 4016 -527 4105 -493
rect 3903 -543 4105 -527
rect 3903 -577 3915 -543
rect 3949 -565 4105 -543
rect 3949 -577 3982 -565
rect 3903 -599 3982 -577
rect 4016 -599 4105 -565
rect 3903 -613 4105 -599
rect 4203 -518 4237 -317
rect 4351 -335 4367 -301
rect 4401 -305 4651 -301
rect 4401 -335 4617 -305
rect 4351 -339 4617 -335
rect 4351 -363 4651 -339
rect 4351 -373 4401 -363
rect 4351 -407 4367 -373
rect 4351 -437 4401 -407
rect 4455 -437 4657 -403
rect 4385 -471 4401 -437
rect 4487 -471 4525 -437
rect 4559 -471 4597 -437
rect 4631 -471 4657 -437
rect 4351 -495 4401 -471
rect 4203 -586 4237 -552
rect 3903 -620 3979 -613
rect 3903 -654 3915 -620
rect 3949 -654 3979 -620
rect 4455 -509 4657 -471
rect 4283 -571 4317 -533
rect 4317 -605 4651 -571
rect 4203 -636 4237 -620
rect 3903 -697 3979 -654
rect 4455 -684 4657 -667
rect 3903 -731 3915 -697
rect 3949 -731 3979 -697
rect 3903 -755 3979 -731
rect 4019 -694 4215 -684
rect 4249 -694 4287 -684
rect 4019 -718 4197 -694
rect 4249 -718 4265 -694
rect 4321 -718 4657 -684
rect 4019 -769 4085 -718
rect 4181 -728 4197 -718
rect 4231 -728 4265 -718
rect 4299 -728 4315 -718
rect 4181 -741 4315 -728
rect 4179 -905 4217 -871
rect 4251 -905 4289 -871
rect 4323 -905 4361 -871
rect 4395 -905 4617 -871
rect 4145 -928 4617 -905
<< viali >>
rect 241 677 275 711
rect 313 677 347 711
rect 740 669 774 703
rect 812 669 846 703
rect 884 669 918 703
rect 232 414 266 448
rect 304 428 308 448
rect 308 428 338 448
rect 304 414 338 428
rect 398 464 432 498
rect 470 488 504 498
rect 470 464 504 488
rect 180 198 214 232
rect 180 126 214 160
rect 180 54 214 88
rect 1260 677 1294 711
rect 1332 677 1366 711
rect 1128 514 1162 548
rect 1200 514 1234 548
rect 1003 454 1013 470
rect 1013 454 1037 470
rect 564 414 598 448
rect 636 414 670 448
rect 1003 436 1037 454
rect 787 368 821 402
rect 859 368 893 402
rect 620 284 654 318
rect 692 284 726 318
rect 756 198 790 232
rect 756 126 790 160
rect 756 54 790 88
rect 1003 386 1013 398
rect 1013 386 1037 398
rect 1003 364 1037 386
rect 1190 362 1224 396
rect 1190 290 1224 324
rect 1332 198 1366 232
rect 1332 126 1366 160
rect 1332 54 1366 88
rect 4453 105 4487 139
rect 4525 105 4559 139
rect 4597 105 4631 139
rect 3974 44 4008 78
rect 3974 -28 4008 6
rect 4237 53 4271 87
rect 4237 11 4257 15
rect 4257 11 4271 15
rect 4237 -19 4271 11
rect 4187 -113 4221 -79
rect 4187 -185 4197 -151
rect 4197 -185 4221 -151
rect 4237 -279 4271 -245
rect 3982 -455 4016 -421
rect 3982 -527 4016 -493
rect 3982 -599 4016 -565
rect 4237 -351 4271 -317
rect 4367 -335 4401 -301
rect 4367 -407 4401 -373
rect 4453 -471 4487 -437
rect 4525 -471 4559 -437
rect 4597 -471 4631 -437
rect 4283 -533 4317 -499
rect 4283 -605 4317 -571
rect 4215 -694 4249 -684
rect 4287 -694 4321 -684
rect 4215 -718 4231 -694
rect 4231 -718 4249 -694
rect 4287 -718 4299 -694
rect 4299 -718 4321 -694
rect 4145 -905 4179 -871
rect 4217 -905 4251 -871
rect 4289 -905 4323 -871
rect 4361 -905 4395 -871
<< metal1 >>
rect 4125 870 4131 922
rect 4183 870 4189 922
rect 4125 858 4189 870
rect 4125 806 4131 858
rect 4183 806 4189 858
rect 4125 778 4161 806
tri 4161 778 4189 806 nw
rect 235 711 1386 776
rect 235 677 241 711
rect 275 677 313 711
rect 347 703 1260 711
rect 347 677 740 703
rect 235 669 740 677
rect 774 669 812 703
rect 846 669 884 703
rect 918 677 1260 703
rect 1294 677 1332 711
rect 1366 677 1386 711
rect 918 669 1386 677
rect 235 588 1386 669
tri 1287 563 1312 588 ne
tri 253 548 265 560 se
rect 265 548 796 560
tri 245 540 253 548 se
rect 253 540 796 548
rect 245 532 796 540
rect 245 514 332 532
tri 332 514 350 532 nw
tri 552 514 570 532 ne
rect 570 514 664 532
tri 664 514 682 532 nw
tri 766 514 784 532 ne
rect 784 514 796 532
rect 245 509 327 514
tri 327 509 332 514 nw
tri 570 509 575 514 ne
rect 575 509 658 514
rect 325 508 326 509
tri 326 508 327 509 nw
tri 575 508 576 509 ne
rect 576 508 577 509
rect 657 508 658 509
tri 658 508 664 514 nw
tri 784 508 790 514 ne
rect 790 508 796 514
rect 848 508 860 560
rect 912 510 1054 560
rect 1056 559 1084 560
rect 1055 511 1085 559
rect 1086 548 1153 560
rect 1205 548 1217 560
rect 1086 514 1128 548
rect 1056 510 1084 511
rect 1086 510 1153 514
rect 912 508 918 510
tri 918 508 920 510 nw
tri 1114 508 1116 510 ne
rect 1116 508 1153 510
rect 1205 508 1217 514
rect 1269 508 1275 560
rect 246 507 324 508
tri 325 507 326 508 nw
tri 576 507 577 508 ne
rect 578 507 656 508
tri 657 507 658 508 nw
tri 1116 507 1117 508 ne
rect 1117 507 1275 508
tri 1117 504 1120 507 ne
rect 1120 504 1275 507
rect 386 498 516 504
tri 1120 502 1122 504 ne
rect 1122 502 1275 504
rect 1312 500 1386 588
tri 230 464 245 479 se
rect 246 478 324 479
tri 325 478 326 479 sw
rect 325 477 326 478
tri 326 477 327 478 sw
rect 245 464 327 477
tri 327 464 340 477 sw
rect 386 464 398 498
rect 432 464 470 498
rect 504 464 516 498
tri 995 480 997 482 se
rect 997 480 1043 482
tri 568 470 577 479 se
rect 578 478 656 479
tri 657 478 658 479 sw
rect 657 477 658 478
tri 658 477 659 478 sw
rect 577 470 659 477
tri 659 470 666 477 sw
tri 220 454 230 464 se
rect 230 454 340 464
tri 340 454 350 464 sw
rect 386 458 516 464
tri 556 458 568 470 se
rect 568 458 666 470
tri 386 454 390 458 ne
rect 390 454 506 458
rect 220 448 350 454
tri 390 448 396 454 ne
rect 396 448 506 454
tri 506 448 516 458 nw
tri 552 454 556 458 se
rect 556 454 666 458
tri 666 454 682 470 sw
rect 552 448 682 454
rect 220 414 232 448
rect 266 414 304 448
rect 338 414 350 448
tri 396 433 411 448 ne
rect 411 435 493 448
tri 493 435 506 448 nw
rect 491 434 492 435
tri 492 434 493 435 nw
rect 412 433 490 434
tri 491 433 492 434 nw
rect 220 408 350 414
rect 552 414 564 448
rect 598 414 636 448
rect 670 414 682 448
rect 552 408 682 414
rect 775 428 783 480
rect 835 428 847 480
rect 899 428 936 480
rect 938 479 966 480
tri 772 405 775 408 se
rect 775 405 936 428
tri 408 402 411 405 se
rect 412 404 490 405
tri 491 404 492 405 sw
tri 771 404 772 405 se
rect 772 404 936 405
rect 491 403 492 404
tri 492 403 493 404 sw
tri 770 403 771 404 se
rect 771 403 936 404
rect 411 402 493 403
tri 493 402 494 403 sw
tri 769 402 770 403 se
rect 770 402 936 403
tri 386 380 408 402 se
rect 408 380 494 402
tri 494 380 516 402 sw
tri 747 380 769 402 se
rect 769 380 787 402
rect 386 368 787 380
rect 821 368 859 402
rect 893 368 936 402
rect 386 352 936 368
rect 937 353 967 479
rect 968 470 1043 480
rect 968 436 1003 470
rect 1037 436 1043 470
rect 968 398 1043 436
rect 968 364 1003 398
rect 1037 364 1043 398
rect 938 352 966 353
rect 968 352 1043 364
rect 1184 396 1230 408
rect 1184 362 1190 396
rect 1224 362 1230 396
tri 1159 324 1184 349 se
rect 1184 324 1230 362
tri 1230 324 1255 349 sw
rect 220 318 1190 324
rect 220 284 620 318
rect 654 284 692 318
rect 726 290 1190 318
rect 1224 290 1386 324
rect 726 284 1386 290
rect 220 278 1386 284
rect 88 232 1386 250
rect 88 198 180 232
rect 214 198 756 232
rect 790 198 1332 232
rect 1366 198 1386 232
rect 88 160 1386 198
rect 88 126 180 160
rect 214 126 756 160
rect 790 126 1332 160
rect 1366 126 1386 160
rect 88 88 1386 126
rect 88 54 180 88
rect 214 54 756 88
rect 790 54 1332 88
rect 1366 54 1386 88
rect 88 48 1386 54
rect 3909 78 4097 84
rect 3909 44 3974 78
rect 4008 44 4097 78
rect 3909 6 4097 44
rect 3909 -28 3974 6
rect 4008 -28 4097 6
rect 3909 -421 4097 -28
rect 4125 -245 4153 778
tri 4153 770 4161 778 nw
rect 4305 726 4311 778
rect 4363 726 4369 778
rect 4305 714 4369 726
rect 4305 662 4311 714
rect 4363 662 4369 714
rect 4305 630 4337 662
tri 4337 630 4369 662 nw
rect 4213 578 4219 630
rect 4271 578 4277 630
rect 4213 566 4277 578
rect 4213 514 4219 566
rect 4271 514 4277 566
rect 4213 87 4277 514
rect 4213 53 4237 87
rect 4271 53 4277 87
rect 4213 15 4277 53
rect 4213 -19 4237 15
rect 4271 -19 4277 15
rect 4213 -31 4277 -19
rect 4181 -79 4227 -67
rect 4181 -113 4187 -79
rect 4221 -92 4227 -79
tri 4227 -92 4252 -67 sw
rect 4221 -113 4250 -92
rect 4181 -151 4250 -113
rect 4181 -185 4187 -151
rect 4221 -172 4250 -151
rect 4251 -171 4252 -93
rect 4221 -185 4227 -172
rect 4181 -197 4227 -185
tri 4227 -197 4252 -172 nw
tri 4280 -92 4305 -67 se
rect 4305 -92 4333 630
tri 4333 626 4337 630 nw
rect 4435 139 4637 231
rect 4435 105 4453 139
rect 4487 105 4525 139
rect 4559 105 4597 139
rect 4631 105 4637 139
rect 4280 -171 4281 -93
rect 4282 -172 4333 -92
tri 4280 -197 4305 -172 ne
tri 4153 -245 4165 -233 sw
tri 4219 -245 4231 -233 se
rect 4231 -245 4277 -233
rect 4125 -258 4165 -245
tri 4165 -258 4178 -245 sw
rect 4125 -338 4176 -258
rect 4177 -337 4178 -259
tri 4206 -258 4219 -245 se
rect 4219 -258 4237 -245
rect 4206 -337 4207 -259
rect 4208 -279 4237 -258
rect 4271 -279 4277 -245
rect 4208 -317 4277 -279
rect 4208 -338 4237 -317
tri 4206 -351 4219 -338 ne
rect 4219 -351 4237 -338
rect 4271 -351 4277 -317
tri 4219 -363 4231 -351 ne
rect 4231 -363 4277 -351
rect 3909 -455 3982 -421
rect 4016 -455 4097 -421
rect 3909 -493 4097 -455
tri 4293 -471 4305 -459 se
rect 4305 -471 4333 -172
tri 4281 -483 4293 -471 se
rect 4293 -483 4333 -471
rect 3909 -527 3982 -493
rect 4016 -527 4097 -493
rect 3909 -565 4097 -527
rect 3909 -599 3982 -565
rect 4016 -599 4097 -565
rect 3909 -936 4097 -599
tri 4277 -487 4281 -483 se
rect 4281 -487 4333 -483
rect 4277 -499 4333 -487
rect 4277 -533 4283 -499
rect 4317 -533 4333 -499
rect 4277 -571 4333 -533
rect 4277 -605 4283 -571
rect 4317 -605 4333 -571
rect 4277 -617 4333 -605
rect 4278 -619 4332 -618
rect 4361 -301 4407 99
rect 4361 -335 4367 -301
rect 4401 -335 4407 -301
rect 4361 -373 4407 -335
rect 4361 -407 4367 -373
rect 4401 -407 4407 -373
rect 4278 -648 4332 -647
tri 4252 -678 4277 -653 se
rect 4277 -678 4333 -649
rect 4203 -684 4333 -678
rect 4203 -718 4215 -684
rect 4249 -718 4287 -684
rect 4321 -718 4333 -684
rect 4203 -724 4333 -718
tri 4336 -865 4361 -840 se
rect 4361 -865 4407 -407
rect 4133 -871 4407 -865
rect 4133 -905 4145 -871
rect 4179 -905 4217 -871
rect 4251 -905 4289 -871
rect 4323 -905 4361 -871
rect 4395 -905 4407 -871
rect 4133 -911 4407 -905
rect 4435 -437 4637 105
rect 4435 -471 4453 -437
rect 4487 -471 4525 -437
rect 4559 -471 4597 -437
rect 4631 -471 4637 -437
rect 4435 -936 4637 -471
<< rmetal1 >>
rect 245 508 325 509
rect 577 508 657 509
rect 1054 559 1056 560
rect 1084 559 1086 560
rect 1054 511 1055 559
rect 1085 511 1086 559
rect 1054 510 1056 511
rect 1084 510 1086 511
rect 245 507 246 508
rect 324 507 325 508
rect 577 507 578 508
rect 656 507 657 508
rect 245 478 246 479
rect 324 478 325 479
rect 245 477 325 478
rect 577 478 578 479
rect 656 478 657 479
rect 577 477 657 478
rect 411 434 491 435
rect 411 433 412 434
rect 490 433 491 434
rect 936 479 938 480
rect 966 479 968 480
rect 411 404 412 405
rect 490 404 491 405
rect 411 403 491 404
rect 936 353 937 479
rect 967 353 968 479
rect 936 352 938 353
rect 966 352 968 353
rect 4250 -93 4252 -92
rect 4250 -171 4251 -93
rect 4250 -172 4252 -171
rect 4280 -93 4282 -92
rect 4281 -171 4282 -93
rect 4280 -172 4282 -171
rect 4176 -259 4178 -258
rect 4176 -337 4177 -259
rect 4176 -338 4178 -337
rect 4206 -259 4208 -258
rect 4207 -337 4208 -259
rect 4206 -338 4208 -337
rect 4277 -618 4333 -617
rect 4277 -619 4278 -618
rect 4332 -619 4333 -618
rect 4277 -648 4278 -647
rect 4332 -648 4333 -647
rect 4277 -649 4333 -648
<< via1 >>
rect 4131 870 4183 922
rect 4131 806 4183 858
rect 796 508 848 560
rect 860 508 912 560
rect 1153 548 1205 560
rect 1217 548 1269 560
rect 1153 514 1162 548
rect 1162 514 1200 548
rect 1200 514 1205 548
rect 1217 514 1234 548
rect 1234 514 1269 548
rect 1153 508 1205 514
rect 1217 508 1269 514
rect 783 428 835 480
rect 847 428 899 480
rect 4311 726 4363 778
rect 4311 662 4363 714
rect 4219 578 4271 630
rect 4219 514 4271 566
<< metal2 >>
tri 1064 870 1116 922 se
rect 1116 870 4131 922
rect 4183 870 4189 922
tri 1052 858 1064 870 se
rect 1064 858 4189 870
tri 1000 806 1052 858 se
rect 1052 806 4131 858
rect 4183 806 4189 858
tri 972 778 1000 806 se
rect 1000 778 1128 806
tri 1128 778 1156 806 nw
tri 960 766 972 778 se
rect 972 766 1116 778
tri 1116 766 1128 778 nw
tri 1216 766 1228 778 se
rect 1228 766 4311 778
tri 920 726 960 766 se
rect 960 762 1112 766
tri 1112 762 1116 766 nw
tri 1212 762 1216 766 se
rect 1216 762 4311 766
rect 960 726 1076 762
tri 1076 726 1112 762 nw
tri 1176 726 1212 762 se
rect 1212 726 4311 762
rect 4363 726 4369 778
tri 908 714 920 726 se
rect 920 714 1064 726
tri 1064 714 1076 726 nw
tri 1164 714 1176 726 se
rect 1176 714 4369 726
tri 856 662 908 714 se
rect 908 662 1012 714
tri 1012 662 1064 714 nw
tri 1112 662 1164 714 se
rect 1164 662 4311 714
rect 4363 662 4369 714
tri 824 630 856 662 se
rect 856 630 980 662
tri 980 630 1012 662 nw
tri 1080 630 1112 662 se
rect 1112 630 1177 662
tri 1177 630 1209 662 nw
tri 804 610 824 630 se
rect 824 610 960 630
tri 960 610 980 630 nw
tri 1060 610 1080 630 se
rect 1080 622 1169 630
tri 1169 622 1177 630 nw
tri 1209 622 1217 630 se
rect 1217 622 4219 630
rect 1080 610 1157 622
tri 1157 610 1169 622 nw
tri 1197 610 1209 622 se
rect 1209 610 4219 622
tri 790 596 804 610 se
rect 804 596 946 610
tri 946 596 960 610 nw
tri 1046 596 1060 610 se
rect 1060 596 1143 610
tri 1143 596 1157 610 nw
tri 1183 596 1197 610 se
rect 1197 596 4219 610
rect 790 578 928 596
tri 928 578 946 596 nw
tri 1028 578 1046 596 se
rect 1046 578 1125 596
tri 1125 578 1143 596 nw
tri 1165 578 1183 596 se
rect 1183 578 4219 596
rect 4271 578 4277 630
rect 790 560 918 578
tri 918 568 928 578 nw
tri 1018 568 1028 578 se
rect 1028 568 1115 578
tri 1115 568 1125 578 nw
tri 1155 568 1165 578 se
rect 1165 568 4277 578
tri 1016 566 1018 568 se
rect 1018 566 1113 568
tri 1113 566 1115 568 nw
tri 1153 566 1155 568 se
rect 1155 566 4277 568
tri 1015 565 1016 566 se
rect 1016 565 1112 566
tri 1112 565 1113 566 nw
tri 1152 565 1153 566 se
rect 1153 565 4219 566
tri 1010 560 1015 565 se
rect 1015 560 1107 565
tri 1107 560 1112 565 nw
tri 1147 560 1152 565 se
rect 1152 560 4219 565
rect 790 508 796 560
rect 848 508 860 560
rect 912 508 918 560
tri 958 508 1010 560 se
rect 1010 508 1055 560
tri 1055 508 1107 560 nw
rect 1147 508 1153 560
rect 1205 508 1217 560
rect 1269 514 4219 560
rect 4271 514 4277 566
rect 1269 508 1275 514
tri 1275 508 1281 514 nw
tri 930 480 958 508 se
rect 958 480 1027 508
tri 1027 480 1055 508 nw
rect 777 428 783 480
rect 835 428 847 480
rect 899 428 975 480
tri 975 428 1027 480 nw
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 4008 0 1 -28
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 0 1 1260 1 0 677
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 0 -1 347 1 0 677
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform 0 -1 1234 1 0 514
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 1037 -1 0 470
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 1224 -1 0 396
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 504 0 1 464
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 338 0 1 414
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 670 0 1 414
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 893 0 1 368
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 726 0 1 284
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 0 -1 4401 1 0 -407
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 0 -1 4317 1 0 -605
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 0 -1 4271 1 0 -351
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 0 -1 4271 1 0 -19
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 0 -1 4221 1 0 -185
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 4215 0 1 -718
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform -1 0 1366 0 1 54
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1707688321
transform -1 0 790 0 1 54
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1707688321
transform -1 0 214 0 1 54
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1707688321
transform -1 0 4016 0 1 -599
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1707688321
transform 0 -1 918 1 0 669
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_5
timestamp 1707688321
transform 0 -1 4631 1 0 105
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_6
timestamp 1707688321
transform 0 -1 4631 1 0 -471
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform -1 0 4395 0 1 -905
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 1 0 1147 0 1 508
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 1 0 790 0 1 508
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 1 0 777 0 1 428
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 4277 0 -1 630
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform -1 0 4369 0 -1 778
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform -1 0 4189 0 -1 922
box 0 0 1 1
use nfet_CDNS_52468879185346  nfet_CDNS_52468879185346_0
timestamp 1707688321
transform 0 -1 4659 -1 0 94
box -79 -26 199 226
use nfet_CDNS_52468879185346  nfet_CDNS_52468879185346_1
timestamp 1707688321
transform 0 1 4459 -1 0 -516
box -79 -26 199 226
use nfet_CDNS_52468879185346  nfet_CDNS_52468879185346_2
timestamp 1707688321
transform 1 0 835 0 -1 226
box -79 -26 199 226
use nfet_CDNS_52468879185346  nfet_CDNS_52468879185346_3
timestamp 1707688321
transform 1 0 225 0 1 26
box -79 -26 199 226
use nfet_CDNS_52468879185525  nfet_CDNS_52468879185525_0
timestamp 1707688321
transform -1 0 711 0 -1 226
box -79 -26 279 110
use nfet_CDNS_52468879185525  nfet_CDNS_52468879185525_1
timestamp 1707688321
transform -1 0 1321 0 -1 226
box -79 -26 279 110
use nfet_CDNS_52468879185525  nfet_CDNS_52468879185525_2
timestamp 1707688321
transform 0 1 4459 1 0 -392
box -79 -26 279 110
use pfet_CDNS_52468879185526  pfet_CDNS_52468879185526_0
timestamp 1707688321
transform 0 1 4023 -1 0 94
box -119 -66 319 150
use pfet_CDNS_52468879185526  pfet_CDNS_52468879185526_1
timestamp 1707688321
transform 1 0 225 0 -1 662
box -119 -66 319 150
use pfet_CDNS_52468879185527  pfet_CDNS_52468879185527_0
timestamp 1707688321
transform -1 0 711 0 -1 778
box -119 -66 239 266
use pfet_CDNS_52468879185527  pfet_CDNS_52468879185527_1
timestamp 1707688321
transform -1 0 1321 0 -1 778
box -119 -66 239 266
use pfet_CDNS_52468879185527  pfet_CDNS_52468879185527_2
timestamp 1707688321
transform 0 1 3907 1 0 -392
box -119 -66 239 266
use pfet_CDNS_52468879185528  pfet_CDNS_52468879185528_0
timestamp 1707688321
transform 0 1 4023 -1 0 -516
box -119 -66 319 150
use pfet_CDNS_52468879185528  pfet_CDNS_52468879185528_1
timestamp 1707688321
transform 1 0 835 0 -1 662
box -119 -66 319 150
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 -1 324 -1 0 546
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 1 0 4139 0 1 -5
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 4315 -1 0 -678
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 -1 4315 -1 0 -135
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform -1 0 4253 0 -1 -502
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 821 1 0 432
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 1 0 454 0 1 370
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 1 0 997 0 1 370
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185523  sky130_fd_io__tk_em1o_b_CDNS_52468879185523_0
timestamp 1707688321
transform 0 1 4277 -1 0 -565
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185524  sky130_fd_io__tk_em1o_b_CDNS_52468879185524_0
timestamp 1707688321
transform -1 0 4260 0 1 -338
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185524  sky130_fd_io__tk_em1o_b_CDNS_52468879185524_1
timestamp 1707688321
transform -1 0 4334 0 1 -172
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185524  sky130_fd_io__tk_em1o_b_CDNS_52468879185524_2
timestamp 1707688321
transform 0 -1 325 1 0 425
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185524  sky130_fd_io__tk_em1o_b_CDNS_52468879185524_3
timestamp 1707688321
transform 0 -1 491 1 0 351
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_52468879185524  sky130_fd_io__tk_em1o_b_CDNS_52468879185524_4
timestamp 1707688321
transform 0 -1 657 1 0 425
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_52468879185521  sky130_fd_io__tk_em1s_b_CDNS_52468879185521_0
timestamp 1707688321
transform -1 0 1138 0 -1 560
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_52468879185522  sky130_fd_io__tk_em1s_b_CDNS_52468879185522_0
timestamp 1707688321
transform 1 0 884 0 -1 480
box 0 0 1 1
<< labels >>
flabel metal1 s 220 278 250 324 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 1360 500 1386 776 0 FreeSans 200 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 235 588 264 776 0 FreeSans 200 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 1366 278 1386 324 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 4435 -900 4637 -880 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 4145 -900 4191 -880 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 3909 -906 4094 -880 0 FreeSans 200 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 1366 48 1386 250 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 517 541 551 555 0 FreeSans 200 0 0 0 out
port 4 nsew
flabel metal1 s 517 361 551 375 0 FreeSans 200 0 0 0 out_n
port 3 nsew
flabel locali s 4220 -416 4220 -416 0 FreeSans 200 270 0 0 a6
flabel locali s 4348 -95 4348 -95 0 FreeSans 200 270 0 0 a5
flabel locali s 4348 -702 4348 -702 0 FreeSans 200 270 0 0 a7
flabel locali s 735 465 735 465 0 FreeSans 200 0 0 0 a2
flabel locali s 414 337 414 337 0 FreeSans 200 0 0 0 a1
flabel locali s 1021 337 1021 337 0 FreeSans 200 0 0 0 a3
flabel locali s 267 34 301 48 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel metal2 s 4304 737 4304 737 0 FreeSans 200 0 0 0 out_n
flabel metal2 s 4250 583 4250 583 0 FreeSans 200 0 0 0 a4
flabel metal2 s 4154 872 4154 872 0 FreeSans 200 0 0 0 out
<< properties >>
string GDS_END 88544154
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88528372
string path 20.300 18.825 27.500 18.825 
<< end >>
