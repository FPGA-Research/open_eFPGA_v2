magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 35 21 735 203
rect 35 17 62 21
rect 28 -17 62 17
<< scnmos >>
rect 113 47 143 177
rect 197 47 227 177
rect 293 47 323 177
rect 401 47 431 177
rect 509 47 539 177
rect 621 47 651 177
<< scpmoshvt >>
rect 113 297 143 497
rect 197 297 227 497
rect 293 297 323 497
rect 401 297 431 497
rect 509 297 539 497
rect 621 297 651 497
<< ndiff >>
rect 61 161 113 177
rect 61 127 69 161
rect 103 127 113 161
rect 61 93 113 127
rect 61 59 69 93
rect 103 59 113 93
rect 61 47 113 59
rect 143 93 197 177
rect 143 59 153 93
rect 187 59 197 93
rect 143 47 197 59
rect 227 161 293 177
rect 227 127 244 161
rect 278 127 293 161
rect 227 93 293 127
rect 227 59 244 93
rect 278 59 293 93
rect 227 47 293 59
rect 323 93 401 177
rect 323 59 345 93
rect 379 59 401 93
rect 323 47 401 59
rect 431 161 509 177
rect 431 127 458 161
rect 492 127 509 161
rect 431 93 509 127
rect 431 59 458 93
rect 492 59 509 93
rect 431 47 509 59
rect 539 161 621 177
rect 539 127 558 161
rect 592 127 621 161
rect 539 47 621 127
rect 651 93 709 177
rect 651 59 661 93
rect 695 59 709 93
rect 651 47 709 59
<< pdiff >>
rect 46 475 113 497
rect 46 441 60 475
rect 94 441 113 475
rect 46 369 113 441
rect 46 335 60 369
rect 94 335 113 369
rect 46 297 113 335
rect 143 485 197 497
rect 143 451 153 485
rect 187 451 197 485
rect 143 417 197 451
rect 143 383 153 417
rect 187 383 197 417
rect 143 297 197 383
rect 227 297 293 497
rect 323 297 401 497
rect 431 485 509 497
rect 431 451 452 485
rect 486 451 509 485
rect 431 417 509 451
rect 431 383 452 417
rect 486 383 509 417
rect 431 297 509 383
rect 539 297 621 497
rect 651 485 709 497
rect 651 451 661 485
rect 695 451 709 485
rect 651 417 709 451
rect 651 383 661 417
rect 695 383 709 417
rect 651 349 709 383
rect 651 315 661 349
rect 695 315 709 349
rect 651 297 709 315
<< ndiffc >>
rect 69 127 103 161
rect 69 59 103 93
rect 153 59 187 93
rect 244 127 278 161
rect 244 59 278 93
rect 345 59 379 93
rect 458 127 492 161
rect 458 59 492 93
rect 558 127 592 161
rect 661 59 695 93
<< pdiffc >>
rect 60 441 94 475
rect 60 335 94 369
rect 153 451 187 485
rect 153 383 187 417
rect 452 451 486 485
rect 452 383 486 417
rect 661 451 695 485
rect 661 383 695 417
rect 661 315 695 349
<< poly >>
rect 113 497 143 523
rect 197 497 227 523
rect 293 497 323 523
rect 401 497 431 523
rect 509 497 539 523
rect 621 497 651 523
rect 113 265 143 297
rect 197 265 227 297
rect 293 265 323 297
rect 401 265 431 297
rect 509 265 539 297
rect 621 265 651 297
rect 77 249 143 265
rect 77 215 93 249
rect 127 215 143 249
rect 77 199 143 215
rect 185 249 251 265
rect 185 215 201 249
rect 235 215 251 249
rect 185 199 251 215
rect 293 249 359 265
rect 293 215 309 249
rect 343 215 359 249
rect 293 199 359 215
rect 401 249 467 265
rect 401 215 417 249
rect 451 215 467 249
rect 401 199 467 215
rect 509 249 575 265
rect 509 215 525 249
rect 559 215 575 249
rect 509 199 575 215
rect 621 249 714 265
rect 621 215 664 249
rect 698 215 714 249
rect 621 199 714 215
rect 113 177 143 199
rect 197 177 227 199
rect 293 177 323 199
rect 401 177 431 199
rect 509 177 539 199
rect 621 177 651 199
rect 113 21 143 47
rect 197 21 227 47
rect 293 21 323 47
rect 401 21 431 47
rect 509 21 539 47
rect 621 21 651 47
<< polycont >>
rect 93 215 127 249
rect 201 215 235 249
rect 309 215 343 249
rect 417 215 451 249
rect 525 215 559 249
rect 664 215 698 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 475 94 491
rect 17 441 60 475
rect 17 369 94 441
rect 17 335 60 369
rect 137 485 195 527
rect 137 451 153 485
rect 187 451 195 485
rect 137 417 195 451
rect 137 383 153 417
rect 187 383 195 417
rect 137 367 195 383
rect 229 485 502 493
rect 229 459 452 485
rect 17 299 94 335
rect 229 333 263 459
rect 436 451 452 459
rect 486 451 502 485
rect 128 299 263 333
rect 17 165 52 299
rect 128 265 162 299
rect 297 265 362 425
rect 436 417 502 451
rect 661 485 719 527
rect 695 451 719 485
rect 661 417 719 451
rect 436 383 452 417
rect 486 383 627 417
rect 436 367 627 383
rect 89 249 162 265
rect 89 215 93 249
rect 127 215 162 249
rect 201 249 251 265
rect 235 215 251 249
rect 293 249 362 265
rect 293 215 309 249
rect 343 215 362 249
rect 89 199 127 215
rect 201 199 235 215
rect 293 199 362 215
rect 396 249 451 332
rect 396 215 417 249
rect 396 199 451 215
rect 488 249 559 332
rect 488 215 525 249
rect 488 199 559 215
rect 593 165 627 367
rect 695 383 719 417
rect 661 349 719 383
rect 695 315 719 349
rect 661 299 719 315
rect 664 249 719 265
rect 698 215 719 249
rect 664 199 719 215
rect 17 161 119 165
rect 17 127 69 161
rect 103 127 119 161
rect 228 161 508 165
rect 17 93 119 127
rect 17 59 69 93
rect 103 59 119 93
rect 17 51 119 59
rect 153 93 187 129
rect 153 17 187 59
rect 228 127 244 161
rect 278 131 458 161
rect 278 127 294 131
rect 228 93 294 127
rect 442 127 458 131
rect 492 127 508 161
rect 542 161 627 165
rect 542 127 558 161
rect 592 127 627 161
rect 228 59 244 93
rect 278 59 294 93
rect 228 51 294 59
rect 329 93 395 97
rect 329 59 345 93
rect 379 59 395 93
rect 329 17 395 59
rect 442 93 508 127
rect 661 93 719 147
rect 442 59 458 93
rect 492 59 661 93
rect 695 59 719 93
rect 442 51 719 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 28 85 62 119 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 28 425 62 459 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 396 289 430 323 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 212 221 246 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 304 221 338 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 396 221 430 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 672 221 706 255 0 FreeSans 250 0 0 0 B1
port 4 nsew signal input
flabel locali s 488 221 522 255 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 304 289 338 323 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 304 357 338 391 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 488 289 522 323 0 FreeSans 250 0 0 0 B2
port 5 nsew signal input
flabel locali s 28 357 62 391 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o32a_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 1455980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1448936
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
