magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 476 226
<< mvnmos >>
rect 0 0 400 200
<< mvndiff >>
rect -50 0 0 200
rect 400 0 450 200
<< poly >>
rect 0 200 400 232
rect 0 -32 400 0
<< metal1 >>
rect -51 -16 -5 186
rect 405 -16 451 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_1
timestamp 1707688321
transform 1 0 400 0 1 0
box -26 -26 82 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 428 85 428 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6689098
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6688204
<< end >>
