magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 319 1066
<< mvpmos >>
rect 0 0 200 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 200 0 250 1000
<< poly >>
rect 0 1000 200 1026
rect 0 -26 200 0
<< locali >>
rect -45 -4 -11 946
rect 211 -4 245 946
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 1036
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_1
timestamp 1707688321
transform 1 0 200 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 228 471 228 471 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 97342688
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97341670
<< end >>
