magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 35330 -1570 35387 -1554
rect 35364 -1604 35387 -1570
rect 35330 -1620 35387 -1604
<< polycont >>
rect -34 16 0 50
rect 35330 -1604 35364 -1570
<< npolyres >>
rect 0 0 35387 66
rect 35321 -96 35387 0
rect -50 -162 35387 -96
rect -50 -258 16 -162
rect -50 -324 35387 -258
rect 35321 -420 35387 -324
rect -50 -486 35387 -420
rect -50 -582 16 -486
rect -50 -648 35387 -582
rect 35321 -744 35387 -648
rect -50 -810 35387 -744
rect -50 -906 16 -810
rect -50 -972 35387 -906
rect 35321 -1068 35387 -972
rect -50 -1134 35387 -1068
rect -50 -1230 16 -1134
rect -50 -1296 35387 -1230
rect 35321 -1392 35387 -1296
rect -50 -1458 35387 -1392
rect -50 -1554 16 -1458
rect -50 -1620 35330 -1554
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 35330 -1570 35371 -1554
rect 35364 -1604 35371 -1570
rect 35330 -1620 35371 -1604
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_0
timestamp 1707688321
transform 1 0 -50 0 1 0
box 0 0 1 1
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_1
timestamp 1707688321
transform 1 0 35314 0 1 -1620
box 0 0 1 1
<< properties >>
string GDS_END 42938942
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42935834
<< end >>
