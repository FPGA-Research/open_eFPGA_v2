magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -128 -43 580 43
<< psubdiff >>
rect -102 -17 -68 17
<< mvpsubdiff >>
rect -34 -17 2 17
rect 36 -17 72 17
rect 106 -17 141 17
rect 175 -17 210 17
rect 244 -17 279 17
rect 313 -17 348 17
rect 382 -17 417 17
rect 451 -17 486 17
rect 520 -17 554 17
<< psubdiffcont >>
rect -68 -17 -66 17
<< mvpsubdiffcont >>
rect -66 -17 -34 17
rect 2 -17 36 17
rect 72 -17 106 17
rect 141 -17 175 17
rect 210 -17 244 17
rect 279 -17 313 17
rect 348 -17 382 17
rect 417 -17 451 17
rect 486 -17 520 17
<< poly >>
rect 53 1291 349 1297
rect 53 1275 386 1291
rect 53 1241 268 1275
rect 302 1241 336 1275
rect 370 1241 386 1275
rect 53 1225 386 1241
rect 515 1225 635 1297
rect 691 1225 811 1297
rect 867 1225 987 1297
rect 1043 1225 1163 1297
rect 1219 1225 1339 1297
rect 1395 1225 1515 1297
rect 53 1117 173 1225
rect 339 1167 635 1183
rect 339 1133 368 1167
rect 402 1133 436 1167
rect 470 1133 504 1167
rect 538 1133 572 1167
rect 606 1133 635 1167
rect 339 1117 635 1133
<< polycont >>
rect 268 1241 302 1275
rect 336 1241 370 1275
rect 368 1133 402 1167
rect 436 1133 470 1167
rect 504 1133 538 1167
rect 572 1133 606 1167
<< locali >>
rect 8 1685 42 1723
rect 360 1685 394 1723
rect 646 1685 680 1723
rect 998 1685 1032 1723
rect 1350 1685 1384 1723
rect 470 1527 504 1565
rect 470 1455 504 1493
rect 822 1527 856 1565
rect 822 1455 856 1493
rect 1174 1527 1208 1565
rect 1174 1455 1208 1493
rect 1526 1527 1560 1565
rect 1526 1455 1560 1493
rect 184 1037 218 1377
rect 252 1241 268 1275
rect 302 1241 336 1275
rect 370 1241 386 1275
rect 998 1241 1032 1275
rect 352 1133 368 1167
rect 402 1133 436 1167
rect 470 1133 504 1167
rect 538 1133 572 1167
rect 606 1133 622 1167
rect 294 1001 328 1039
rect 294 929 328 967
rect 646 1001 680 1039
rect 646 929 680 967
rect 42 807 80 841
rect 432 807 470 841
rect 294 205 328 243
rect 294 133 328 171
rect 646 205 680 243
rect 646 133 680 171
rect -102 -17 -68 17
rect -34 -17 2 17
rect 36 -17 72 17
rect 106 -17 141 17
rect 175 -17 210 17
rect 244 -17 279 17
rect 313 -17 348 17
rect 382 -17 417 17
rect 451 -17 486 17
rect 520 -17 554 17
<< viali >>
rect 8 1723 42 1757
rect 8 1651 42 1685
rect 360 1723 394 1757
rect 360 1651 394 1685
rect 646 1723 680 1757
rect 646 1651 680 1685
rect 998 1723 1032 1757
rect 998 1651 1032 1685
rect 1350 1723 1384 1757
rect 1350 1651 1384 1685
rect 470 1565 504 1599
rect 470 1493 504 1527
rect 470 1421 504 1455
rect 822 1565 856 1599
rect 822 1493 856 1527
rect 822 1421 856 1455
rect 1174 1565 1208 1599
rect 1174 1493 1208 1527
rect 1174 1421 1208 1455
rect 1526 1565 1560 1599
rect 1526 1493 1560 1527
rect 1526 1421 1560 1455
rect 294 1039 328 1073
rect 294 967 328 1001
rect 294 895 328 929
rect 646 1039 680 1073
rect 646 967 680 1001
rect 646 895 680 929
rect 8 807 42 841
rect 80 807 114 841
rect 398 807 432 841
rect 470 807 504 841
rect 294 243 328 277
rect 294 171 328 205
rect 294 99 328 133
rect 646 243 680 277
rect 646 171 680 205
rect 646 99 680 133
<< metal1 >>
rect 2 1757 1390 1769
rect 2 1723 8 1757
rect 42 1723 360 1757
rect 394 1723 646 1757
rect 680 1723 998 1757
rect 1032 1723 1350 1757
rect 1384 1723 1390 1757
rect 2 1685 1390 1723
rect 2 1651 8 1685
rect 42 1651 360 1685
rect 394 1651 646 1685
rect 680 1651 998 1685
rect 1032 1651 1350 1685
rect 1384 1651 1390 1685
rect 2 1639 1390 1651
rect 464 1599 1576 1611
rect 464 1565 470 1599
rect 504 1565 822 1599
rect 856 1565 1174 1599
rect 1208 1565 1526 1599
rect 1560 1565 1576 1599
rect 464 1527 1576 1565
rect 464 1493 470 1527
rect 504 1493 822 1527
rect 856 1493 1174 1527
rect 1208 1493 1526 1527
rect 1560 1493 1576 1527
rect 464 1455 1576 1493
rect 464 1421 470 1455
rect 504 1421 822 1455
rect 856 1421 1174 1455
rect 1208 1421 1526 1455
rect 1560 1421 1576 1455
rect 464 1409 1576 1421
rect 288 1073 686 1085
rect 288 1039 294 1073
rect 328 1039 646 1073
rect 680 1039 686 1073
rect 288 1001 686 1039
rect 288 967 294 1001
rect 328 967 646 1001
rect 680 967 686 1001
rect 288 929 686 967
rect 288 895 294 929
rect 328 895 646 929
rect 680 895 686 929
rect 288 883 686 895
rect -4 841 516 847
rect -4 807 8 841
rect 42 807 80 841
rect 114 807 398 841
rect 432 807 470 841
rect 504 807 516 841
rect -4 801 516 807
rect 288 277 686 289
rect 288 243 294 277
rect 328 243 646 277
rect 680 243 686 277
rect 288 205 686 243
rect 288 171 294 205
rect 328 171 646 205
rect 680 171 686 205
rect 288 133 686 171
rect 288 99 294 133
rect 328 99 646 133
rect 680 99 686 133
rect 288 87 686 99
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 1 1350 1 0 1651
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 1 8 1 0 1651
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 1 360 1 0 1651
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 1 646 1 0 1651
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 1 998 1 0 1651
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 1 0 8 0 -1 841
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 1 0 398 0 -1 841
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 1560 -1 0 1599
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 856 -1 0 1599
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 504 -1 0 1599
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 -1 1208 -1 0 1599
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 -1 328 1 0 99
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 680 1 0 99
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 328 1 0 895
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 680 1 0 895
box 0 0 1 1
use nfet_CDNS_52468879185124  nfet_CDNS_52468879185124_0
timestamp 1707688321
transform 1 0 53 0 1 91
box -79 -26 199 1026
use nfet_CDNS_524688791851201  nfet_CDNS_524688791851201_0
timestamp 1707688321
transform 1 0 339 0 1 91
box -79 -26 375 1026
use pfet_CDNS_52468879185312  pfet_CDNS_52468879185312_0
timestamp 1707688321
transform 1 0 53 0 -1 2323
box -119 -66 415 1066
use pfet_CDNS_524688791851202  pfet_CDNS_524688791851202_0
timestamp 1707688321
transform 1 0 515 0 -1 2323
box -119 -66 1119 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 252 -1 0 1291
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 -1 622 1 0 1117
box 0 0 1 1
use PYL1_CDNS_52468879185407  PYL1_CDNS_52468879185407_0
timestamp 1707688321
transform 0 -1 1490 -1 0 1291
box 0 0 66 950
<< labels >>
flabel comment s 1015 1235 1015 1235 0 FreeSans 400 0 0 0 ie_n
flabel comment s 488 1175 488 1175 0 FreeSans 400 0 0 0 ie
flabel comment s 198 1165 198 1165 0 FreeSans 400 0 0 0 out
flabel comment s 318 1279 318 1279 0 FreeSans 400 0 0 0 in
flabel metal1 s 416 827 416 827 0 FreeSans 400 0 0 0 n<1>
flabel metal1 s 642 87 663 289 7 FreeSans 400 0 0 0 vgnd
port 1 nsew
flabel metal1 s 1542 1409 1566 1611 7 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 642 883 663 1085 7 FreeSans 400 0 0 0 vgnd
port 1 nsew
flabel locali s 184 1241 218 1275 0 FreeSans 600 0 0 0 out
port 4 nsew
flabel locali s 302 1241 336 1275 0 FreeSans 600 0 0 0 in
port 5 nsew
flabel locali s 998 1241 1032 1275 0 FreeSans 600 0 0 0 ie_n
port 6 nsew
flabel locali s 470 1133 504 1167 0 FreeSans 600 0 0 0 ie
port 7 nsew
<< properties >>
string GDS_END 85761990
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85757434
string path -2.550 0.000 13.850 0.000 
<< end >>
