magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 547 874 568 923
<< obsli1 >>
rect 0 1152 1360 1218
rect 0 1046 66 1152
rect 100 1080 1260 1118
rect 0 1012 611 1046
rect 0 906 66 1012
rect 648 978 712 1080
rect 1294 1046 1360 1152
rect 746 1012 1360 1046
rect 100 940 1260 978
rect 0 872 611 906
rect 0 766 66 872
rect 648 838 712 940
rect 1294 906 1360 1012
rect 746 872 1360 906
rect 100 800 1260 838
rect 0 732 611 766
rect 0 626 66 732
rect 648 698 712 800
rect 1294 766 1360 872
rect 746 732 1360 766
rect 100 660 1260 698
rect 0 592 611 626
rect 0 486 66 592
rect 648 558 712 660
rect 1294 626 1360 732
rect 746 592 1360 626
rect 100 520 1260 558
rect 0 452 611 486
rect 0 346 66 452
rect 648 418 712 520
rect 1294 486 1360 592
rect 746 452 1360 486
rect 100 380 1260 418
rect 0 312 611 346
rect 0 206 66 312
rect 648 278 712 380
rect 1294 346 1360 452
rect 746 312 1360 346
rect 100 240 1260 278
rect 0 172 611 206
rect 0 66 66 172
rect 648 138 712 240
rect 1294 206 1360 312
rect 746 172 1360 206
rect 100 100 1260 138
rect 1294 66 1360 172
rect 0 0 1360 66
<< obsm1 >>
rect 0 1152 1360 1218
rect 0 66 66 1152
rect 94 641 122 1124
rect 150 669 178 1152
rect 206 641 234 1124
rect 262 669 290 1152
rect 318 641 346 1124
rect 374 669 402 1152
rect 430 641 458 1124
rect 486 669 514 1152
rect 542 641 570 1124
rect 598 669 626 1152
rect 654 641 706 1124
rect 734 669 762 1152
rect 790 641 818 1124
rect 846 669 874 1152
rect 902 641 930 1124
rect 958 669 986 1152
rect 1014 641 1042 1124
rect 1070 669 1098 1152
rect 1126 641 1154 1124
rect 1182 669 1210 1152
rect 1238 641 1266 1124
rect 94 577 1266 641
rect 94 94 122 577
rect 150 66 178 549
rect 206 94 234 577
rect 262 66 290 549
rect 318 94 346 577
rect 374 66 402 549
rect 430 94 458 577
rect 486 66 514 549
rect 542 94 570 577
rect 598 66 626 549
rect 654 94 706 577
rect 734 66 762 549
rect 790 94 818 577
rect 846 66 874 549
rect 902 94 930 577
rect 958 66 986 549
rect 1014 94 1042 577
rect 1070 66 1098 549
rect 1126 94 1154 577
rect 1182 66 1210 549
rect 1238 94 1266 577
rect 1294 66 1360 1152
rect 0 0 1360 66
<< obsm2 >>
rect 0 1152 619 1218
rect 0 1068 66 1152
rect 647 1124 713 1218
rect 741 1152 1360 1218
rect 94 1096 1266 1124
rect 0 1040 619 1068
rect 0 956 66 1040
rect 647 1012 713 1096
rect 1294 1068 1360 1152
rect 741 1040 1360 1068
rect 94 984 1266 1012
rect 0 928 619 956
rect 0 844 66 928
rect 647 900 713 984
rect 1294 956 1360 1040
rect 741 928 1360 956
rect 94 872 1266 900
rect 0 816 619 844
rect 0 732 66 816
rect 647 788 713 872
rect 1294 844 1360 928
rect 741 816 1360 844
rect 94 760 1266 788
rect 0 665 619 732
rect 647 637 713 760
rect 1294 732 1360 816
rect 741 665 1360 732
rect 0 581 1360 637
rect 0 486 619 553
rect 0 402 66 486
rect 647 458 713 581
rect 741 486 1360 553
rect 94 430 1266 458
rect 0 374 619 402
rect 0 290 66 374
rect 647 346 713 430
rect 1294 402 1360 486
rect 741 374 1360 402
rect 94 318 1266 346
rect 0 262 619 290
rect 0 178 66 262
rect 647 234 713 318
rect 1294 290 1360 374
rect 741 262 1360 290
rect 94 206 1266 234
rect 0 150 619 178
rect 0 66 66 150
rect 647 122 713 206
rect 1294 178 1360 262
rect 741 150 1360 178
rect 94 94 1266 122
rect 0 0 619 66
rect 647 0 713 94
rect 1294 66 1360 150
rect 741 0 1360 66
<< metal3 >>
rect 0 1152 1360 1218
rect 0 66 66 1152
rect 126 642 194 1092
rect 254 702 322 1152
rect 382 642 450 1092
rect 510 702 578 1152
rect 638 642 722 1092
rect 782 702 850 1152
rect 910 642 978 1092
rect 1038 702 1106 1152
rect 1166 642 1234 1092
rect 126 576 1234 642
rect 126 126 194 576
rect 254 66 322 516
rect 382 126 450 576
rect 510 66 578 516
rect 638 126 722 576
rect 782 66 850 516
rect 910 126 978 576
rect 1038 66 1106 516
rect 1166 126 1234 576
rect 1294 66 1360 1152
rect 0 0 1360 66
<< metal4 >>
rect 0 0 1360 1218
<< labels >>
rlabel metal3 s 1294 66 1360 1152 6 C0
port 1 nsew
rlabel metal3 s 1038 702 1106 1152 6 C0
port 1 nsew
rlabel metal3 s 1038 66 1106 516 6 C0
port 1 nsew
rlabel metal3 s 782 702 850 1152 6 C0
port 1 nsew
rlabel metal3 s 782 66 850 516 6 C0
port 1 nsew
rlabel metal3 s 510 702 578 1152 6 C0
port 1 nsew
rlabel metal3 s 510 66 578 516 6 C0
port 1 nsew
rlabel metal3 s 254 702 322 1152 6 C0
port 1 nsew
rlabel metal3 s 254 66 322 516 6 C0
port 1 nsew
rlabel metal3 s 0 1152 1360 1218 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 1152 6 C0
port 1 nsew
rlabel metal3 s 0 0 1360 66 6 C0
port 1 nsew
rlabel metal3 s 1166 642 1234 1092 6 C1
port 2 nsew
rlabel metal3 s 1166 126 1234 576 6 C1
port 2 nsew
rlabel metal3 s 910 642 978 1092 6 C1
port 2 nsew
rlabel metal3 s 910 126 978 576 6 C1
port 2 nsew
rlabel metal3 s 638 642 722 1092 6 C1
port 2 nsew
rlabel metal3 s 638 126 722 576 6 C1
port 2 nsew
rlabel metal3 s 382 642 450 1092 6 C1
port 2 nsew
rlabel metal3 s 382 126 450 576 6 C1
port 2 nsew
rlabel metal3 s 126 642 194 1092 6 C1
port 2 nsew
rlabel metal3 s 126 576 1234 642 6 C1
port 2 nsew
rlabel metal3 s 126 126 194 576 6 C1
port 2 nsew
rlabel metal4 s 0 0 1360 1218 6 MET4
port 4 nsew
rlabel pwell s 547 874 568 923 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1360 1218
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 303366
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 276488
string device primitive
<< end >>