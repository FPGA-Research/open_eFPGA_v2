magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 161 125
<< metal1 >>
rect -6 125 167 128
rect -6 0 0 125
rect 161 0 167 125
rect -6 -3 167 0
<< properties >>
string GDS_END 87633658
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87632246
<< end >>
