magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 46 -77 3217 683
<< mvnmos >>
rect 125 57 225 657
rect 281 57 381 657
rect 574 57 674 657
rect 730 57 830 657
rect 886 57 986 657
rect 1042 57 1142 657
rect 1198 57 1298 657
rect 1354 57 1454 657
rect 1510 57 1610 657
rect 1666 57 1766 657
rect 1822 57 1922 657
rect 1978 57 2078 657
rect 2134 57 2234 657
rect 2290 57 2390 657
rect 2570 57 2670 657
rect 2726 57 2826 657
rect 2882 57 2982 657
rect 3038 57 3138 657
<< mvndiff >>
rect 72 579 125 657
rect 72 545 80 579
rect 114 545 125 579
rect 72 511 125 545
rect 72 477 80 511
rect 114 477 125 511
rect 72 443 125 477
rect 72 409 80 443
rect 114 409 125 443
rect 72 375 125 409
rect 72 341 80 375
rect 114 341 125 375
rect 72 307 125 341
rect 72 273 80 307
rect 114 273 125 307
rect 72 239 125 273
rect 72 205 80 239
rect 114 205 125 239
rect 72 171 125 205
rect 72 137 80 171
rect 114 137 125 171
rect 72 103 125 137
rect 72 69 80 103
rect 114 69 125 103
rect 72 57 125 69
rect 225 579 281 657
rect 225 545 236 579
rect 270 545 281 579
rect 225 511 281 545
rect 225 477 236 511
rect 270 477 281 511
rect 225 443 281 477
rect 225 409 236 443
rect 270 409 281 443
rect 225 375 281 409
rect 225 341 236 375
rect 270 341 281 375
rect 225 307 281 341
rect 225 273 236 307
rect 270 273 281 307
rect 225 239 281 273
rect 225 205 236 239
rect 270 205 281 239
rect 225 171 281 205
rect 225 137 236 171
rect 270 137 281 171
rect 225 103 281 137
rect 225 69 236 103
rect 270 69 281 103
rect 225 57 281 69
rect 381 579 434 657
rect 381 545 392 579
rect 426 545 434 579
rect 381 511 434 545
rect 381 477 392 511
rect 426 477 434 511
rect 381 443 434 477
rect 381 409 392 443
rect 426 409 434 443
rect 381 375 434 409
rect 381 341 392 375
rect 426 341 434 375
rect 381 307 434 341
rect 381 273 392 307
rect 426 273 434 307
rect 381 239 434 273
rect 381 205 392 239
rect 426 205 434 239
rect 381 171 434 205
rect 381 137 392 171
rect 426 137 434 171
rect 381 103 434 137
rect 381 69 392 103
rect 426 69 434 103
rect 381 57 434 69
rect 521 579 574 657
rect 521 545 529 579
rect 563 545 574 579
rect 521 511 574 545
rect 521 477 529 511
rect 563 477 574 511
rect 521 443 574 477
rect 521 409 529 443
rect 563 409 574 443
rect 521 375 574 409
rect 521 341 529 375
rect 563 341 574 375
rect 521 307 574 341
rect 521 273 529 307
rect 563 273 574 307
rect 521 239 574 273
rect 521 205 529 239
rect 563 205 574 239
rect 521 171 574 205
rect 521 137 529 171
rect 563 137 574 171
rect 521 103 574 137
rect 521 69 529 103
rect 563 69 574 103
rect 521 57 574 69
rect 674 579 730 657
rect 674 545 685 579
rect 719 545 730 579
rect 674 511 730 545
rect 674 477 685 511
rect 719 477 730 511
rect 674 443 730 477
rect 674 409 685 443
rect 719 409 730 443
rect 674 375 730 409
rect 674 341 685 375
rect 719 341 730 375
rect 674 307 730 341
rect 674 273 685 307
rect 719 273 730 307
rect 674 239 730 273
rect 674 205 685 239
rect 719 205 730 239
rect 674 171 730 205
rect 674 137 685 171
rect 719 137 730 171
rect 674 103 730 137
rect 674 69 685 103
rect 719 69 730 103
rect 674 57 730 69
rect 830 579 886 657
rect 830 545 841 579
rect 875 545 886 579
rect 830 511 886 545
rect 830 477 841 511
rect 875 477 886 511
rect 830 443 886 477
rect 830 409 841 443
rect 875 409 886 443
rect 830 375 886 409
rect 830 341 841 375
rect 875 341 886 375
rect 830 307 886 341
rect 830 273 841 307
rect 875 273 886 307
rect 830 239 886 273
rect 830 205 841 239
rect 875 205 886 239
rect 830 171 886 205
rect 830 137 841 171
rect 875 137 886 171
rect 830 103 886 137
rect 830 69 841 103
rect 875 69 886 103
rect 830 57 886 69
rect 986 579 1042 657
rect 986 545 997 579
rect 1031 545 1042 579
rect 986 511 1042 545
rect 986 477 997 511
rect 1031 477 1042 511
rect 986 443 1042 477
rect 986 409 997 443
rect 1031 409 1042 443
rect 986 375 1042 409
rect 986 341 997 375
rect 1031 341 1042 375
rect 986 307 1042 341
rect 986 273 997 307
rect 1031 273 1042 307
rect 986 239 1042 273
rect 986 205 997 239
rect 1031 205 1042 239
rect 986 171 1042 205
rect 986 137 997 171
rect 1031 137 1042 171
rect 986 103 1042 137
rect 986 69 997 103
rect 1031 69 1042 103
rect 986 57 1042 69
rect 1142 579 1198 657
rect 1142 545 1153 579
rect 1187 545 1198 579
rect 1142 511 1198 545
rect 1142 477 1153 511
rect 1187 477 1198 511
rect 1142 443 1198 477
rect 1142 409 1153 443
rect 1187 409 1198 443
rect 1142 375 1198 409
rect 1142 341 1153 375
rect 1187 341 1198 375
rect 1142 307 1198 341
rect 1142 273 1153 307
rect 1187 273 1198 307
rect 1142 239 1198 273
rect 1142 205 1153 239
rect 1187 205 1198 239
rect 1142 171 1198 205
rect 1142 137 1153 171
rect 1187 137 1198 171
rect 1142 103 1198 137
rect 1142 69 1153 103
rect 1187 69 1198 103
rect 1142 57 1198 69
rect 1298 579 1354 657
rect 1298 545 1309 579
rect 1343 545 1354 579
rect 1298 511 1354 545
rect 1298 477 1309 511
rect 1343 477 1354 511
rect 1298 443 1354 477
rect 1298 409 1309 443
rect 1343 409 1354 443
rect 1298 375 1354 409
rect 1298 341 1309 375
rect 1343 341 1354 375
rect 1298 307 1354 341
rect 1298 273 1309 307
rect 1343 273 1354 307
rect 1298 239 1354 273
rect 1298 205 1309 239
rect 1343 205 1354 239
rect 1298 171 1354 205
rect 1298 137 1309 171
rect 1343 137 1354 171
rect 1298 103 1354 137
rect 1298 69 1309 103
rect 1343 69 1354 103
rect 1298 57 1354 69
rect 1454 579 1510 657
rect 1454 545 1465 579
rect 1499 545 1510 579
rect 1454 511 1510 545
rect 1454 477 1465 511
rect 1499 477 1510 511
rect 1454 443 1510 477
rect 1454 409 1465 443
rect 1499 409 1510 443
rect 1454 375 1510 409
rect 1454 341 1465 375
rect 1499 341 1510 375
rect 1454 307 1510 341
rect 1454 273 1465 307
rect 1499 273 1510 307
rect 1454 239 1510 273
rect 1454 205 1465 239
rect 1499 205 1510 239
rect 1454 171 1510 205
rect 1454 137 1465 171
rect 1499 137 1510 171
rect 1454 103 1510 137
rect 1454 69 1465 103
rect 1499 69 1510 103
rect 1454 57 1510 69
rect 1610 579 1666 657
rect 1610 545 1621 579
rect 1655 545 1666 579
rect 1610 511 1666 545
rect 1610 477 1621 511
rect 1655 477 1666 511
rect 1610 443 1666 477
rect 1610 409 1621 443
rect 1655 409 1666 443
rect 1610 375 1666 409
rect 1610 341 1621 375
rect 1655 341 1666 375
rect 1610 307 1666 341
rect 1610 273 1621 307
rect 1655 273 1666 307
rect 1610 239 1666 273
rect 1610 205 1621 239
rect 1655 205 1666 239
rect 1610 171 1666 205
rect 1610 137 1621 171
rect 1655 137 1666 171
rect 1610 103 1666 137
rect 1610 69 1621 103
rect 1655 69 1666 103
rect 1610 57 1666 69
rect 1766 579 1822 657
rect 1766 545 1777 579
rect 1811 545 1822 579
rect 1766 511 1822 545
rect 1766 477 1777 511
rect 1811 477 1822 511
rect 1766 443 1822 477
rect 1766 409 1777 443
rect 1811 409 1822 443
rect 1766 375 1822 409
rect 1766 341 1777 375
rect 1811 341 1822 375
rect 1766 307 1822 341
rect 1766 273 1777 307
rect 1811 273 1822 307
rect 1766 239 1822 273
rect 1766 205 1777 239
rect 1811 205 1822 239
rect 1766 171 1822 205
rect 1766 137 1777 171
rect 1811 137 1822 171
rect 1766 103 1822 137
rect 1766 69 1777 103
rect 1811 69 1822 103
rect 1766 57 1822 69
rect 1922 579 1978 657
rect 1922 545 1933 579
rect 1967 545 1978 579
rect 1922 511 1978 545
rect 1922 477 1933 511
rect 1967 477 1978 511
rect 1922 443 1978 477
rect 1922 409 1933 443
rect 1967 409 1978 443
rect 1922 375 1978 409
rect 1922 341 1933 375
rect 1967 341 1978 375
rect 1922 307 1978 341
rect 1922 273 1933 307
rect 1967 273 1978 307
rect 1922 239 1978 273
rect 1922 205 1933 239
rect 1967 205 1978 239
rect 1922 171 1978 205
rect 1922 137 1933 171
rect 1967 137 1978 171
rect 1922 103 1978 137
rect 1922 69 1933 103
rect 1967 69 1978 103
rect 1922 57 1978 69
rect 2078 579 2134 657
rect 2078 545 2089 579
rect 2123 545 2134 579
rect 2078 511 2134 545
rect 2078 477 2089 511
rect 2123 477 2134 511
rect 2078 443 2134 477
rect 2078 409 2089 443
rect 2123 409 2134 443
rect 2078 375 2134 409
rect 2078 341 2089 375
rect 2123 341 2134 375
rect 2078 307 2134 341
rect 2078 273 2089 307
rect 2123 273 2134 307
rect 2078 239 2134 273
rect 2078 205 2089 239
rect 2123 205 2134 239
rect 2078 171 2134 205
rect 2078 137 2089 171
rect 2123 137 2134 171
rect 2078 103 2134 137
rect 2078 69 2089 103
rect 2123 69 2134 103
rect 2078 57 2134 69
rect 2234 579 2290 657
rect 2234 545 2245 579
rect 2279 545 2290 579
rect 2234 511 2290 545
rect 2234 477 2245 511
rect 2279 477 2290 511
rect 2234 443 2290 477
rect 2234 409 2245 443
rect 2279 409 2290 443
rect 2234 375 2290 409
rect 2234 341 2245 375
rect 2279 341 2290 375
rect 2234 307 2290 341
rect 2234 273 2245 307
rect 2279 273 2290 307
rect 2234 239 2290 273
rect 2234 205 2245 239
rect 2279 205 2290 239
rect 2234 171 2290 205
rect 2234 137 2245 171
rect 2279 137 2290 171
rect 2234 103 2290 137
rect 2234 69 2245 103
rect 2279 69 2290 103
rect 2234 57 2290 69
rect 2390 579 2443 657
rect 2390 545 2401 579
rect 2435 545 2443 579
rect 2390 511 2443 545
rect 2390 477 2401 511
rect 2435 477 2443 511
rect 2390 443 2443 477
rect 2390 409 2401 443
rect 2435 409 2443 443
rect 2390 375 2443 409
rect 2390 341 2401 375
rect 2435 341 2443 375
rect 2390 307 2443 341
rect 2390 273 2401 307
rect 2435 273 2443 307
rect 2390 239 2443 273
rect 2390 205 2401 239
rect 2435 205 2443 239
rect 2390 171 2443 205
rect 2390 137 2401 171
rect 2435 137 2443 171
rect 2390 103 2443 137
rect 2390 69 2401 103
rect 2435 69 2443 103
rect 2390 57 2443 69
rect 2517 579 2570 657
rect 2517 545 2525 579
rect 2559 545 2570 579
rect 2517 511 2570 545
rect 2517 477 2525 511
rect 2559 477 2570 511
rect 2517 443 2570 477
rect 2517 409 2525 443
rect 2559 409 2570 443
rect 2517 375 2570 409
rect 2517 341 2525 375
rect 2559 341 2570 375
rect 2517 307 2570 341
rect 2517 273 2525 307
rect 2559 273 2570 307
rect 2517 239 2570 273
rect 2517 205 2525 239
rect 2559 205 2570 239
rect 2517 171 2570 205
rect 2517 137 2525 171
rect 2559 137 2570 171
rect 2517 103 2570 137
rect 2517 69 2525 103
rect 2559 69 2570 103
rect 2517 57 2570 69
rect 2670 579 2726 657
rect 2670 545 2681 579
rect 2715 545 2726 579
rect 2670 511 2726 545
rect 2670 477 2681 511
rect 2715 477 2726 511
rect 2670 443 2726 477
rect 2670 409 2681 443
rect 2715 409 2726 443
rect 2670 375 2726 409
rect 2670 341 2681 375
rect 2715 341 2726 375
rect 2670 307 2726 341
rect 2670 273 2681 307
rect 2715 273 2726 307
rect 2670 239 2726 273
rect 2670 205 2681 239
rect 2715 205 2726 239
rect 2670 171 2726 205
rect 2670 137 2681 171
rect 2715 137 2726 171
rect 2670 103 2726 137
rect 2670 69 2681 103
rect 2715 69 2726 103
rect 2670 57 2726 69
rect 2826 579 2882 657
rect 2826 545 2837 579
rect 2871 545 2882 579
rect 2826 511 2882 545
rect 2826 477 2837 511
rect 2871 477 2882 511
rect 2826 443 2882 477
rect 2826 409 2837 443
rect 2871 409 2882 443
rect 2826 375 2882 409
rect 2826 341 2837 375
rect 2871 341 2882 375
rect 2826 307 2882 341
rect 2826 273 2837 307
rect 2871 273 2882 307
rect 2826 239 2882 273
rect 2826 205 2837 239
rect 2871 205 2882 239
rect 2826 171 2882 205
rect 2826 137 2837 171
rect 2871 137 2882 171
rect 2826 103 2882 137
rect 2826 69 2837 103
rect 2871 69 2882 103
rect 2826 57 2882 69
rect 2982 579 3038 657
rect 2982 545 2993 579
rect 3027 545 3038 579
rect 2982 511 3038 545
rect 2982 477 2993 511
rect 3027 477 3038 511
rect 2982 443 3038 477
rect 2982 409 2993 443
rect 3027 409 3038 443
rect 2982 375 3038 409
rect 2982 341 2993 375
rect 3027 341 3038 375
rect 2982 307 3038 341
rect 2982 273 2993 307
rect 3027 273 3038 307
rect 2982 239 3038 273
rect 2982 205 2993 239
rect 3027 205 3038 239
rect 2982 171 3038 205
rect 2982 137 2993 171
rect 3027 137 3038 171
rect 2982 103 3038 137
rect 2982 69 2993 103
rect 3027 69 3038 103
rect 2982 57 3038 69
rect 3138 579 3191 657
rect 3138 545 3149 579
rect 3183 545 3191 579
rect 3138 511 3191 545
rect 3138 477 3149 511
rect 3183 477 3191 511
rect 3138 443 3191 477
rect 3138 409 3149 443
rect 3183 409 3191 443
rect 3138 375 3191 409
rect 3138 341 3149 375
rect 3183 341 3191 375
rect 3138 307 3191 341
rect 3138 273 3149 307
rect 3183 273 3191 307
rect 3138 239 3191 273
rect 3138 205 3149 239
rect 3183 205 3191 239
rect 3138 171 3191 205
rect 3138 137 3149 171
rect 3183 137 3191 171
rect 3138 103 3191 137
rect 3138 69 3149 103
rect 3183 69 3191 103
rect 3138 57 3191 69
<< mvndiffc >>
rect 80 545 114 579
rect 80 477 114 511
rect 80 409 114 443
rect 80 341 114 375
rect 80 273 114 307
rect 80 205 114 239
rect 80 137 114 171
rect 80 69 114 103
rect 236 545 270 579
rect 236 477 270 511
rect 236 409 270 443
rect 236 341 270 375
rect 236 273 270 307
rect 236 205 270 239
rect 236 137 270 171
rect 236 69 270 103
rect 392 545 426 579
rect 392 477 426 511
rect 392 409 426 443
rect 392 341 426 375
rect 392 273 426 307
rect 392 205 426 239
rect 392 137 426 171
rect 392 69 426 103
rect 529 545 563 579
rect 529 477 563 511
rect 529 409 563 443
rect 529 341 563 375
rect 529 273 563 307
rect 529 205 563 239
rect 529 137 563 171
rect 529 69 563 103
rect 685 545 719 579
rect 685 477 719 511
rect 685 409 719 443
rect 685 341 719 375
rect 685 273 719 307
rect 685 205 719 239
rect 685 137 719 171
rect 685 69 719 103
rect 841 545 875 579
rect 841 477 875 511
rect 841 409 875 443
rect 841 341 875 375
rect 841 273 875 307
rect 841 205 875 239
rect 841 137 875 171
rect 841 69 875 103
rect 997 545 1031 579
rect 997 477 1031 511
rect 997 409 1031 443
rect 997 341 1031 375
rect 997 273 1031 307
rect 997 205 1031 239
rect 997 137 1031 171
rect 997 69 1031 103
rect 1153 545 1187 579
rect 1153 477 1187 511
rect 1153 409 1187 443
rect 1153 341 1187 375
rect 1153 273 1187 307
rect 1153 205 1187 239
rect 1153 137 1187 171
rect 1153 69 1187 103
rect 1309 545 1343 579
rect 1309 477 1343 511
rect 1309 409 1343 443
rect 1309 341 1343 375
rect 1309 273 1343 307
rect 1309 205 1343 239
rect 1309 137 1343 171
rect 1309 69 1343 103
rect 1465 545 1499 579
rect 1465 477 1499 511
rect 1465 409 1499 443
rect 1465 341 1499 375
rect 1465 273 1499 307
rect 1465 205 1499 239
rect 1465 137 1499 171
rect 1465 69 1499 103
rect 1621 545 1655 579
rect 1621 477 1655 511
rect 1621 409 1655 443
rect 1621 341 1655 375
rect 1621 273 1655 307
rect 1621 205 1655 239
rect 1621 137 1655 171
rect 1621 69 1655 103
rect 1777 545 1811 579
rect 1777 477 1811 511
rect 1777 409 1811 443
rect 1777 341 1811 375
rect 1777 273 1811 307
rect 1777 205 1811 239
rect 1777 137 1811 171
rect 1777 69 1811 103
rect 1933 545 1967 579
rect 1933 477 1967 511
rect 1933 409 1967 443
rect 1933 341 1967 375
rect 1933 273 1967 307
rect 1933 205 1967 239
rect 1933 137 1967 171
rect 1933 69 1967 103
rect 2089 545 2123 579
rect 2089 477 2123 511
rect 2089 409 2123 443
rect 2089 341 2123 375
rect 2089 273 2123 307
rect 2089 205 2123 239
rect 2089 137 2123 171
rect 2089 69 2123 103
rect 2245 545 2279 579
rect 2245 477 2279 511
rect 2245 409 2279 443
rect 2245 341 2279 375
rect 2245 273 2279 307
rect 2245 205 2279 239
rect 2245 137 2279 171
rect 2245 69 2279 103
rect 2401 545 2435 579
rect 2401 477 2435 511
rect 2401 409 2435 443
rect 2401 341 2435 375
rect 2401 273 2435 307
rect 2401 205 2435 239
rect 2401 137 2435 171
rect 2401 69 2435 103
rect 2525 545 2559 579
rect 2525 477 2559 511
rect 2525 409 2559 443
rect 2525 341 2559 375
rect 2525 273 2559 307
rect 2525 205 2559 239
rect 2525 137 2559 171
rect 2525 69 2559 103
rect 2681 545 2715 579
rect 2681 477 2715 511
rect 2681 409 2715 443
rect 2681 341 2715 375
rect 2681 273 2715 307
rect 2681 205 2715 239
rect 2681 137 2715 171
rect 2681 69 2715 103
rect 2837 545 2871 579
rect 2837 477 2871 511
rect 2837 409 2871 443
rect 2837 341 2871 375
rect 2837 273 2871 307
rect 2837 205 2871 239
rect 2837 137 2871 171
rect 2837 69 2871 103
rect 2993 545 3027 579
rect 2993 477 3027 511
rect 2993 409 3027 443
rect 2993 341 3027 375
rect 2993 273 3027 307
rect 2993 205 3027 239
rect 2993 137 3027 171
rect 2993 69 3027 103
rect 3149 545 3183 579
rect 3149 477 3183 511
rect 3149 409 3183 443
rect 3149 341 3183 375
rect 3149 273 3183 307
rect 3149 205 3183 239
rect 3149 137 3183 171
rect 3149 69 3183 103
<< mvpsubdiff >>
rect 72 -51 96 -17
rect 130 -51 166 -17
rect 200 -51 235 -17
rect 269 -51 304 -17
rect 338 -51 373 -17
rect 407 -51 442 -17
rect 476 -51 511 -17
rect 545 -51 580 -17
rect 614 -51 649 -17
rect 683 -51 718 -17
rect 752 -51 787 -17
rect 821 -51 856 -17
rect 890 -51 925 -17
rect 959 -51 994 -17
rect 1028 -51 1063 -17
rect 1097 -51 1132 -17
rect 1166 -51 1201 -17
rect 1235 -51 1270 -17
rect 1304 -51 1339 -17
rect 1373 -51 1408 -17
rect 1442 -51 1477 -17
rect 1511 -51 1546 -17
rect 1580 -51 1615 -17
rect 1649 -51 1684 -17
rect 1718 -51 1753 -17
rect 1787 -51 1822 -17
rect 1856 -51 1891 -17
rect 1925 -51 1960 -17
rect 1994 -51 2029 -17
rect 2063 -51 2098 -17
rect 2132 -51 2167 -17
rect 2201 -51 2236 -17
rect 2270 -51 2305 -17
rect 2339 -51 2374 -17
rect 2408 -51 2443 -17
rect 2477 -51 2512 -17
rect 2546 -51 2581 -17
rect 2615 -51 2650 -17
rect 2684 -51 2719 -17
rect 2753 -51 2788 -17
rect 2822 -51 2857 -17
rect 2891 -51 2926 -17
rect 2960 -51 2995 -17
rect 3029 -51 3064 -17
rect 3098 -51 3133 -17
rect 3167 -51 3191 -17
<< mvpsubdiffcont >>
rect 96 -51 130 -17
rect 166 -51 200 -17
rect 235 -51 269 -17
rect 304 -51 338 -17
rect 373 -51 407 -17
rect 442 -51 476 -17
rect 511 -51 545 -17
rect 580 -51 614 -17
rect 649 -51 683 -17
rect 718 -51 752 -17
rect 787 -51 821 -17
rect 856 -51 890 -17
rect 925 -51 959 -17
rect 994 -51 1028 -17
rect 1063 -51 1097 -17
rect 1132 -51 1166 -17
rect 1201 -51 1235 -17
rect 1270 -51 1304 -17
rect 1339 -51 1373 -17
rect 1408 -51 1442 -17
rect 1477 -51 1511 -17
rect 1546 -51 1580 -17
rect 1615 -51 1649 -17
rect 1684 -51 1718 -17
rect 1753 -51 1787 -17
rect 1822 -51 1856 -17
rect 1891 -51 1925 -17
rect 1960 -51 1994 -17
rect 2029 -51 2063 -17
rect 2098 -51 2132 -17
rect 2167 -51 2201 -17
rect 2236 -51 2270 -17
rect 2305 -51 2339 -17
rect 2374 -51 2408 -17
rect 2443 -51 2477 -17
rect 2512 -51 2546 -17
rect 2581 -51 2615 -17
rect 2650 -51 2684 -17
rect 2719 -51 2753 -17
rect 2788 -51 2822 -17
rect 2857 -51 2891 -17
rect 2926 -51 2960 -17
rect 2995 -51 3029 -17
rect 3064 -51 3098 -17
rect 3133 -51 3167 -17
<< poly >>
rect 125 819 225 835
rect 125 785 160 819
rect 194 785 225 819
rect 125 751 225 785
rect 125 717 160 751
rect 194 717 225 751
rect 125 657 225 717
rect 281 819 381 835
rect 281 785 313 819
rect 347 785 381 819
rect 281 751 381 785
rect 281 717 313 751
rect 347 717 381 751
rect 281 657 381 717
rect 574 739 1454 755
rect 574 705 590 739
rect 624 705 664 739
rect 698 705 738 739
rect 772 705 812 739
rect 846 705 886 739
rect 920 705 960 739
rect 994 705 1034 739
rect 1068 705 1108 739
rect 1142 705 1182 739
rect 1216 705 1256 739
rect 1290 705 1330 739
rect 1364 705 1404 739
rect 1438 705 1454 739
rect 574 689 1454 705
rect 574 657 674 689
rect 730 657 830 689
rect 886 657 986 689
rect 1042 657 1142 689
rect 1198 657 1298 689
rect 1354 657 1454 689
rect 1510 739 2826 755
rect 1510 705 1526 739
rect 1560 705 1596 739
rect 1630 705 1666 739
rect 1700 705 1736 739
rect 1770 705 1806 739
rect 1840 705 1876 739
rect 1910 705 1946 739
rect 1980 705 2016 739
rect 2050 705 2086 739
rect 2120 705 2155 739
rect 2189 705 2224 739
rect 2258 705 2293 739
rect 2327 705 2362 739
rect 2396 705 2431 739
rect 2465 705 2500 739
rect 2534 705 2569 739
rect 2603 705 2638 739
rect 2672 705 2707 739
rect 2741 705 2776 739
rect 2810 705 2826 739
rect 1510 689 2826 705
rect 1510 657 1610 689
rect 1666 657 1766 689
rect 1822 657 1922 689
rect 1978 657 2078 689
rect 2134 657 2234 689
rect 2290 657 2390 689
rect 2570 657 2670 689
rect 2726 657 2826 689
rect 2882 739 3138 755
rect 2882 705 2898 739
rect 2932 705 2993 739
rect 3027 705 3088 739
rect 3122 705 3138 739
rect 2882 689 3138 705
rect 2882 657 2982 689
rect 3038 657 3138 689
rect 125 25 225 57
rect 281 25 381 57
rect 574 25 674 57
rect 730 25 830 57
rect 886 25 986 57
rect 1042 25 1142 57
rect 1198 25 1298 57
rect 1354 25 1454 57
rect 1510 25 1610 57
rect 1666 25 1766 57
rect 1822 25 1922 57
rect 1978 25 2078 57
rect 2134 25 2234 57
rect 2290 25 2390 57
rect 2570 25 2670 57
rect 2726 25 2826 57
rect 2882 25 2982 57
rect 3038 25 3138 57
<< polycont >>
rect 160 785 194 819
rect 160 717 194 751
rect 313 785 347 819
rect 313 717 347 751
rect 590 705 624 739
rect 664 705 698 739
rect 738 705 772 739
rect 812 705 846 739
rect 886 705 920 739
rect 960 705 994 739
rect 1034 705 1068 739
rect 1108 705 1142 739
rect 1182 705 1216 739
rect 1256 705 1290 739
rect 1330 705 1364 739
rect 1404 705 1438 739
rect 1526 705 1560 739
rect 1596 705 1630 739
rect 1666 705 1700 739
rect 1736 705 1770 739
rect 1806 705 1840 739
rect 1876 705 1910 739
rect 1946 705 1980 739
rect 2016 705 2050 739
rect 2086 705 2120 739
rect 2155 705 2189 739
rect 2224 705 2258 739
rect 2293 705 2327 739
rect 2362 705 2396 739
rect 2431 705 2465 739
rect 2500 705 2534 739
rect 2569 705 2603 739
rect 2638 705 2672 739
rect 2707 705 2741 739
rect 2776 705 2810 739
rect 2898 705 2932 739
rect 2993 705 3027 739
rect 3088 705 3122 739
<< locali >>
rect 149 819 202 835
rect 149 785 160 819
rect 194 785 202 819
rect 149 751 202 785
rect 313 819 347 835
rect 313 773 347 785
rect 149 717 160 751
rect 194 717 202 751
rect 323 751 361 773
rect 347 739 361 751
rect 597 739 640 773
rect 674 739 717 773
rect 751 739 794 773
rect 828 739 871 773
rect 905 739 948 773
rect 982 739 1025 773
rect 1059 739 1102 773
rect 1136 739 1179 773
rect 1213 739 1255 773
rect 1289 739 1331 773
rect 1365 739 1407 773
rect 149 677 202 717
rect 313 701 347 717
rect 574 705 590 739
rect 624 705 664 739
rect 698 705 738 739
rect 772 705 812 739
rect 846 705 886 739
rect 920 705 960 739
rect 994 705 1034 739
rect 1068 705 1108 739
rect 1142 705 1182 739
rect 1216 705 1256 739
rect 1290 705 1330 739
rect 1364 705 1404 739
rect 1438 705 1454 739
rect 1510 705 1526 739
rect 1590 705 1596 739
rect 1663 705 1666 739
rect 1700 705 1702 739
rect 1770 705 1775 739
rect 1840 705 1848 739
rect 1910 705 1921 739
rect 1980 705 1994 739
rect 2050 705 2067 739
rect 2120 705 2140 739
rect 2189 705 2213 739
rect 2258 705 2286 739
rect 2327 705 2359 739
rect 2396 705 2431 739
rect 2466 705 2500 739
rect 2539 705 2569 739
rect 2612 705 2638 739
rect 2685 705 2707 739
rect 2758 705 2776 739
rect 2810 705 2826 739
rect 2882 705 2898 739
rect 2932 738 2993 739
rect 3027 738 3088 739
rect 3122 738 3138 739
rect 2947 705 2993 738
rect 3036 705 3088 738
rect 3124 705 3138 738
rect 2947 704 3002 705
rect 3036 704 3090 705
rect 149 643 162 677
rect 196 643 202 677
rect 149 605 202 643
rect 80 579 114 595
rect 149 571 162 605
rect 196 571 202 605
rect 236 579 270 595
rect 80 511 114 545
rect 80 443 114 477
rect 80 375 114 409
rect 80 307 114 341
rect 80 239 114 273
rect 80 171 114 205
rect 80 103 114 137
rect 80 53 114 65
rect 236 511 270 545
rect 236 443 270 477
rect 392 579 426 595
rect 529 579 563 595
rect 685 579 719 595
rect 392 511 426 545
rect 563 545 568 572
rect 530 538 568 545
rect 841 579 875 595
rect 997 579 1031 595
rect 392 443 426 477
rect 236 375 270 409
rect 390 409 392 420
rect 529 511 563 538
rect 685 511 719 545
rect 875 545 881 572
rect 843 538 881 545
rect 1153 579 1187 595
rect 841 511 875 538
rect 529 443 563 477
rect 719 477 724 495
rect 686 461 724 477
rect 997 511 1031 545
rect 1150 545 1153 572
rect 1309 579 1343 595
rect 1187 545 1188 572
rect 1150 538 1188 545
rect 1465 579 1499 595
rect 1621 579 1655 595
rect 426 409 428 420
rect 390 386 428 409
rect 236 307 270 341
rect 236 239 270 273
rect 236 171 270 205
rect 236 103 270 137
rect 236 53 270 69
rect 392 375 426 386
rect 392 307 426 341
rect 392 239 426 273
rect 392 171 426 205
rect 392 103 426 137
rect 392 53 426 69
rect 529 375 563 409
rect 529 307 563 341
rect 529 239 563 273
rect 529 171 563 205
rect 529 103 563 137
rect 529 53 563 69
rect 685 443 719 461
rect 685 375 719 409
rect 685 307 719 341
rect 685 239 719 273
rect 685 171 719 205
rect 685 103 719 137
rect 685 53 719 69
rect 841 443 875 477
rect 1153 511 1187 538
rect 1031 477 1035 495
rect 997 461 1035 477
rect 1309 511 1343 545
rect 1499 545 1505 572
rect 1467 538 1505 545
rect 1777 579 1811 595
rect 841 375 875 409
rect 841 307 875 341
rect 841 239 875 273
rect 841 171 875 205
rect 841 103 875 137
rect 841 53 875 69
rect 997 443 1031 461
rect 997 375 1031 409
rect 997 307 1031 341
rect 997 239 1031 273
rect 997 171 1031 205
rect 997 103 1031 137
rect 997 53 1031 69
rect 1153 443 1187 477
rect 1307 477 1309 495
rect 1465 511 1499 538
rect 1343 477 1345 495
rect 1307 461 1345 477
rect 1153 375 1187 409
rect 1153 307 1187 341
rect 1153 239 1187 273
rect 1153 171 1187 205
rect 1153 103 1187 137
rect 1153 53 1187 69
rect 1309 443 1343 461
rect 1309 375 1343 409
rect 1309 307 1343 341
rect 1309 239 1343 273
rect 1309 171 1343 205
rect 1309 103 1343 137
rect 1309 53 1343 69
rect 1465 443 1499 477
rect 1465 375 1499 409
rect 1465 307 1499 341
rect 1465 239 1499 273
rect 1465 171 1499 205
rect 1465 103 1499 137
rect 1465 53 1499 69
rect 1621 511 1655 545
rect 1933 579 1967 595
rect 1811 545 1815 572
rect 1777 538 1815 545
rect 2089 579 2123 595
rect 2245 579 2279 595
rect 1621 443 1655 477
rect 1621 375 1655 409
rect 1621 307 1655 341
rect 1621 239 1655 273
rect 1621 171 1655 205
rect 1621 103 1655 137
rect 1621 53 1655 65
rect 1777 511 1811 538
rect 1777 443 1811 477
rect 1777 375 1811 409
rect 1777 307 1811 341
rect 1777 239 1811 273
rect 1777 171 1811 205
rect 1777 103 1811 137
rect 1777 53 1811 69
rect 1933 511 1967 545
rect 2077 545 2089 572
rect 2077 538 2115 545
rect 2401 579 2435 595
rect 2525 579 2559 595
rect 1933 443 1967 477
rect 1933 375 1967 409
rect 1933 307 1967 341
rect 1933 239 1967 273
rect 1933 171 1967 205
rect 1933 103 1967 137
rect 1933 53 1967 65
rect 2089 511 2123 538
rect 2089 443 2123 477
rect 2089 375 2123 409
rect 2089 307 2123 341
rect 2089 239 2123 273
rect 2089 171 2123 205
rect 2089 103 2123 137
rect 2089 53 2123 69
rect 2245 511 2279 545
rect 2377 545 2401 572
rect 2377 538 2415 545
rect 2245 443 2279 477
rect 2245 375 2279 409
rect 2245 307 2279 341
rect 2245 239 2279 273
rect 2245 171 2279 205
rect 2245 103 2279 137
rect 2245 53 2279 65
rect 2401 511 2435 538
rect 2525 511 2559 545
rect 2681 579 2715 595
rect 2681 511 2715 545
rect 2401 443 2435 477
rect 2559 477 2586 503
rect 2548 469 2586 477
rect 2837 579 2871 595
rect 2837 511 2871 545
rect 2993 579 3027 595
rect 2993 511 3027 545
rect 2401 375 2435 409
rect 2401 307 2435 341
rect 2401 239 2435 273
rect 2401 171 2435 205
rect 2401 103 2435 137
rect 2401 53 2435 69
rect 2525 443 2559 469
rect 2525 375 2559 409
rect 2525 307 2559 341
rect 2525 239 2559 273
rect 2525 171 2559 205
rect 2525 103 2559 137
rect 2525 53 2559 69
rect 2681 443 2715 477
rect 2871 477 2880 503
rect 2842 469 2880 477
rect 3149 579 3183 595
rect 3149 511 3183 545
rect 2681 375 2715 409
rect 2681 307 2715 341
rect 2681 239 2715 273
rect 2681 171 2715 205
rect 2681 103 2715 137
rect 2681 53 2715 65
rect 2837 443 2871 469
rect 2993 443 3027 477
rect 3128 477 3149 503
rect 3128 469 3166 477
rect 3149 443 3183 469
rect 2837 375 2871 409
rect 2985 409 2993 420
rect 2985 386 3023 409
rect 2837 307 2871 341
rect 2837 239 2871 273
rect 2837 171 2871 205
rect 2837 103 2871 137
rect 2837 53 2871 69
rect 2993 375 3027 386
rect 2993 307 3027 341
rect 2993 239 3027 273
rect 2993 171 3027 205
rect 2993 103 3027 137
rect 2993 53 3027 69
rect 3149 375 3183 409
rect 3149 307 3183 341
rect 3149 239 3183 273
rect 3149 171 3183 205
rect 3149 103 3183 137
rect 3149 53 3183 69
rect 72 -51 77 -17
rect 130 -51 150 -17
rect 200 -51 223 -17
rect 269 -51 296 -17
rect 338 -51 369 -17
rect 407 -51 442 -17
rect 476 -51 511 -17
rect 549 -51 580 -17
rect 622 -51 649 -17
rect 695 -51 718 -17
rect 768 -51 787 -17
rect 841 -51 856 -17
rect 914 -51 925 -17
rect 987 -51 994 -17
rect 1060 -51 1063 -17
rect 1097 -51 1099 -17
rect 1166 -51 1172 -17
rect 1235 -51 1245 -17
rect 1304 -51 1318 -17
rect 1373 -51 1391 -17
rect 1442 -51 1464 -17
rect 1511 -51 1537 -17
rect 1580 -51 1610 -17
rect 1649 -51 1683 -17
rect 1718 -51 1753 -17
rect 1790 -51 1822 -17
rect 1863 -51 1891 -17
rect 1936 -51 1960 -17
rect 2009 -51 2029 -17
rect 2082 -51 2098 -17
rect 2155 -51 2167 -17
rect 2228 -51 2236 -17
rect 2301 -51 2305 -17
rect 2339 -51 2340 -17
rect 2408 -51 2413 -17
rect 2477 -51 2486 -17
rect 2546 -51 2559 -17
rect 2615 -51 2631 -17
rect 2684 -51 2703 -17
rect 2753 -51 2775 -17
rect 2822 -51 2847 -17
rect 2891 -51 2919 -17
rect 2960 -51 2991 -17
rect 3029 -51 3063 -17
rect 3098 -51 3133 -17
rect 3169 -51 3191 -17
<< viali >>
rect 289 751 323 773
rect 289 739 313 751
rect 313 739 323 751
rect 361 739 395 773
rect 563 739 597 773
rect 640 739 674 773
rect 717 739 751 773
rect 794 739 828 773
rect 871 739 905 773
rect 948 739 982 773
rect 1025 739 1059 773
rect 1102 739 1136 773
rect 1179 739 1213 773
rect 1255 739 1289 773
rect 1331 739 1365 773
rect 1407 739 1441 773
rect 1556 705 1560 739
rect 1560 705 1590 739
rect 1629 705 1630 739
rect 1630 705 1663 739
rect 1702 705 1736 739
rect 1775 705 1806 739
rect 1806 705 1809 739
rect 1848 705 1876 739
rect 1876 705 1882 739
rect 1921 705 1946 739
rect 1946 705 1955 739
rect 1994 705 2016 739
rect 2016 705 2028 739
rect 2067 705 2086 739
rect 2086 705 2101 739
rect 2140 705 2155 739
rect 2155 705 2174 739
rect 2213 705 2224 739
rect 2224 705 2247 739
rect 2286 705 2293 739
rect 2293 705 2320 739
rect 2359 705 2362 739
rect 2362 705 2393 739
rect 2432 705 2465 739
rect 2465 705 2466 739
rect 2505 705 2534 739
rect 2534 705 2539 739
rect 2578 705 2603 739
rect 2603 705 2612 739
rect 2651 705 2672 739
rect 2672 705 2685 739
rect 2724 705 2741 739
rect 2741 705 2758 739
rect 2913 705 2932 738
rect 2932 705 2947 738
rect 3002 705 3027 738
rect 3027 705 3036 738
rect 3090 705 3122 738
rect 3122 705 3124 738
rect 2913 704 2947 705
rect 3002 704 3036 705
rect 3090 704 3124 705
rect 162 643 196 677
rect 162 571 196 605
rect 80 137 114 171
rect 80 69 114 99
rect 80 65 114 69
rect 496 545 529 572
rect 529 545 530 572
rect 496 538 530 545
rect 568 538 602 572
rect 356 386 390 420
rect 809 545 841 572
rect 841 545 843 572
rect 809 538 843 545
rect 881 538 915 572
rect 652 477 685 495
rect 685 477 686 495
rect 652 461 686 477
rect 724 461 758 495
rect 1116 538 1150 572
rect 1188 538 1222 572
rect 428 386 462 420
rect 963 461 997 495
rect 1035 461 1069 495
rect 1433 545 1465 572
rect 1465 545 1467 572
rect 1433 538 1467 545
rect 1505 538 1539 572
rect 1273 461 1307 495
rect 1345 461 1379 495
rect 1743 538 1777 572
rect 1815 538 1849 572
rect 1621 137 1655 171
rect 1621 69 1655 99
rect 1621 65 1655 69
rect 2043 538 2077 572
rect 2115 545 2123 572
rect 2123 545 2149 572
rect 2115 538 2149 545
rect 1933 137 1967 171
rect 1933 69 1967 99
rect 1933 65 1967 69
rect 2343 538 2377 572
rect 2415 545 2435 572
rect 2435 545 2449 572
rect 2415 538 2449 545
rect 2245 137 2279 171
rect 2245 69 2279 99
rect 2245 65 2279 69
rect 2514 477 2525 503
rect 2525 477 2548 503
rect 2514 469 2548 477
rect 2586 469 2620 503
rect 2808 477 2837 503
rect 2837 477 2842 503
rect 2808 469 2842 477
rect 2880 469 2914 503
rect 2681 137 2715 171
rect 2681 69 2715 99
rect 2681 65 2715 69
rect 3094 469 3128 503
rect 3166 477 3183 503
rect 3183 477 3200 503
rect 3166 469 3200 477
rect 2951 386 2985 420
rect 3023 409 3027 420
rect 3027 409 3057 420
rect 3023 386 3057 409
rect 77 -51 96 -17
rect 96 -51 111 -17
rect 150 -51 166 -17
rect 166 -51 184 -17
rect 223 -51 235 -17
rect 235 -51 257 -17
rect 296 -51 304 -17
rect 304 -51 330 -17
rect 369 -51 373 -17
rect 373 -51 403 -17
rect 442 -51 476 -17
rect 515 -51 545 -17
rect 545 -51 549 -17
rect 588 -51 614 -17
rect 614 -51 622 -17
rect 661 -51 683 -17
rect 683 -51 695 -17
rect 734 -51 752 -17
rect 752 -51 768 -17
rect 807 -51 821 -17
rect 821 -51 841 -17
rect 880 -51 890 -17
rect 890 -51 914 -17
rect 953 -51 959 -17
rect 959 -51 987 -17
rect 1026 -51 1028 -17
rect 1028 -51 1060 -17
rect 1099 -51 1132 -17
rect 1132 -51 1133 -17
rect 1172 -51 1201 -17
rect 1201 -51 1206 -17
rect 1245 -51 1270 -17
rect 1270 -51 1279 -17
rect 1318 -51 1339 -17
rect 1339 -51 1352 -17
rect 1391 -51 1408 -17
rect 1408 -51 1425 -17
rect 1464 -51 1477 -17
rect 1477 -51 1498 -17
rect 1537 -51 1546 -17
rect 1546 -51 1571 -17
rect 1610 -51 1615 -17
rect 1615 -51 1644 -17
rect 1683 -51 1684 -17
rect 1684 -51 1717 -17
rect 1756 -51 1787 -17
rect 1787 -51 1790 -17
rect 1829 -51 1856 -17
rect 1856 -51 1863 -17
rect 1902 -51 1925 -17
rect 1925 -51 1936 -17
rect 1975 -51 1994 -17
rect 1994 -51 2009 -17
rect 2048 -51 2063 -17
rect 2063 -51 2082 -17
rect 2121 -51 2132 -17
rect 2132 -51 2155 -17
rect 2194 -51 2201 -17
rect 2201 -51 2228 -17
rect 2267 -51 2270 -17
rect 2270 -51 2301 -17
rect 2340 -51 2374 -17
rect 2413 -51 2443 -17
rect 2443 -51 2447 -17
rect 2486 -51 2512 -17
rect 2512 -51 2520 -17
rect 2559 -51 2581 -17
rect 2581 -51 2593 -17
rect 2631 -51 2650 -17
rect 2650 -51 2665 -17
rect 2703 -51 2719 -17
rect 2719 -51 2737 -17
rect 2775 -51 2788 -17
rect 2788 -51 2809 -17
rect 2847 -51 2857 -17
rect 2857 -51 2881 -17
rect 2919 -51 2926 -17
rect 2926 -51 2953 -17
rect 2991 -51 2995 -17
rect 2995 -51 3025 -17
rect 3063 -51 3064 -17
rect 3064 -51 3097 -17
rect 3135 -51 3167 -17
rect 3167 -51 3169 -17
<< metal1 >>
tri 1452 810 1464 822 se
rect 1464 810 2807 822
tri 2807 810 2819 822 sw
tri 1422 780 1452 810 se
rect 1452 780 2819 810
rect 1235 779 2819 780
tri 2819 779 2850 810 sw
rect 277 773 459 779
rect 461 778 497 779
rect 277 739 289 773
rect 323 739 361 773
rect 395 739 459 773
rect 277 733 459 739
rect 460 734 498 778
rect 499 776 2850 779
rect 499 773 1453 776
rect 499 739 563 773
rect 597 739 640 773
rect 674 739 717 773
rect 751 739 794 773
rect 828 739 871 773
rect 905 739 948 773
rect 982 739 1025 773
rect 1059 739 1102 773
rect 1136 739 1179 773
rect 1213 739 1255 773
rect 1289 739 1331 773
rect 1365 739 1407 773
rect 1441 739 1453 773
tri 1453 745 1484 776 nw
tri 2787 745 2818 776 ne
rect 2818 745 2850 776
tri 2850 745 2884 779 sw
tri 1538 739 1544 745 se
rect 1544 744 2770 745
tri 2818 744 2819 745 ne
rect 2819 744 2884 745
tri 2884 744 2885 745 sw
rect 1544 739 2773 744
rect 461 733 497 734
rect 499 733 1453 739
tri 1532 733 1538 739 se
rect 1538 733 1556 739
tri 1504 705 1532 733 se
rect 1532 705 1556 733
rect 1590 705 1629 739
rect 1663 705 1702 739
rect 1736 705 1775 739
rect 1809 705 1848 739
rect 1882 705 1921 739
rect 1955 705 1994 739
rect 2028 705 2067 739
rect 2101 705 2140 739
rect 2174 705 2213 739
rect 2247 705 2286 739
rect 2320 705 2359 739
rect 2393 705 2432 739
rect 2466 705 2505 739
rect 2539 705 2578 739
rect 2612 705 2651 739
rect 2685 705 2724 739
rect 2758 738 2773 739
tri 2773 738 2779 744 sw
tri 2819 738 2825 744 ne
rect 2825 738 3296 744
rect 2758 705 2779 738
tri 1503 704 1504 705 se
rect 1504 704 2779 705
tri 2779 704 2813 738 sw
tri 2825 704 2859 738 ne
rect 2859 704 2913 738
rect 2947 704 3002 738
rect 3036 704 3090 738
rect 3124 704 3296 738
tri 1498 699 1503 704 se
rect 1503 699 2813 704
tri 2813 699 2818 704 sw
tri 2859 699 2864 704 ne
rect 2864 699 3296 704
tri 1488 689 1498 699 se
rect 1498 689 1559 699
rect 156 686 202 689
tri 1485 686 1488 689 se
rect 1488 686 1559 689
tri 1559 686 1572 699 nw
rect 2680 698 2818 699
tri 2818 698 2819 699 sw
tri 2864 698 2865 699 ne
rect 2865 698 3296 699
rect 2680 692 2819 698
tri 2751 686 2757 692 ne
rect 2757 686 2819 692
tri 2819 686 2831 698 sw
rect 156 677 228 686
rect 230 685 266 686
rect 156 643 162 677
rect 196 643 228 677
rect 156 634 228 643
rect 229 635 267 685
rect 230 634 266 635
rect 268 634 1507 686
tri 1507 634 1559 686 nw
tri 2757 674 2769 686 ne
rect 2769 674 2831 686
tri 2831 674 2843 686 sw
tri 2769 670 2773 674 ne
rect 2773 670 2843 674
tri 2773 634 2809 670 ne
rect 2809 634 2843 670
tri 2843 634 2883 674 sw
rect 3244 666 3296 698
rect 3245 664 3295 665
rect 156 605 202 634
rect 156 571 162 605
rect 196 571 202 605
tri 2809 600 2843 634 ne
rect 2843 600 2883 634
tri 2883 600 2917 634 sw
rect 3245 627 3295 628
rect 3244 600 3296 626
tri 2843 578 2865 600 ne
rect 2865 578 3165 600
rect 156 559 202 571
rect 484 572 2461 578
tri 2865 574 2869 578 ne
rect 2869 574 3165 578
rect 484 538 496 572
rect 530 538 568 572
rect 602 538 809 572
rect 843 538 881 572
rect 915 538 1116 572
rect 1150 538 1188 572
rect 1222 538 1433 572
rect 1467 538 1505 572
rect 1539 538 1743 572
rect 1777 538 1815 572
rect 1849 538 2043 572
rect 2077 538 2115 572
rect 2149 538 2343 572
rect 2377 538 2415 572
rect 2449 538 2461 572
tri 2869 548 2895 574 ne
rect 2895 548 3165 574
rect 3166 549 3167 599
rect 3203 549 3204 599
rect 3205 548 3296 600
rect 484 532 2461 538
rect 2502 503 3212 509
rect 344 455 555 501
rect 557 500 593 501
rect 556 456 594 500
rect 595 495 1391 501
rect 595 461 652 495
rect 686 461 724 495
rect 758 461 963 495
rect 997 461 1035 495
rect 1069 461 1273 495
rect 1307 461 1345 495
rect 1379 461 1391 495
rect 2502 469 2514 503
rect 2548 469 2586 503
rect 2620 469 2808 503
rect 2842 469 2880 503
rect 2914 469 3094 503
rect 3128 469 3166 503
rect 3200 469 3212 503
rect 2502 463 3212 469
rect 557 455 593 456
rect 595 455 1391 461
rect 344 426 443 455
rect 344 420 2852 426
rect 344 386 356 420
rect 390 386 428 420
rect 462 386 2852 420
rect 344 380 2852 386
rect 2853 381 2854 425
rect 2890 381 2891 425
rect 2892 420 3069 426
rect 2892 386 2951 420
rect 2985 386 3023 420
rect 3057 386 3069 420
rect 2892 380 3069 386
rect 3244 183 3296 548
rect 65 171 3367 183
rect 65 137 80 171
rect 114 137 1621 171
rect 1655 137 1933 171
rect 1967 137 2245 171
rect 2279 137 2681 171
rect 2715 137 3367 171
rect 65 99 3367 137
rect 65 65 80 99
rect 114 65 1621 99
rect 1655 65 1933 99
rect 1967 65 2245 99
rect 2279 65 2681 99
rect 2715 65 3367 99
rect 65 -6 3367 65
rect 65 -17 3202 -6
rect 65 -51 77 -17
rect 111 -51 150 -17
rect 184 -51 223 -17
rect 257 -51 296 -17
rect 330 -51 369 -17
rect 403 -51 442 -17
rect 476 -51 515 -17
rect 549 -51 588 -17
rect 622 -51 661 -17
rect 695 -51 734 -17
rect 768 -51 807 -17
rect 841 -51 880 -17
rect 914 -51 953 -17
rect 987 -51 1026 -17
rect 1060 -51 1099 -17
rect 1133 -51 1172 -17
rect 1206 -51 1245 -17
rect 1279 -51 1318 -17
rect 1352 -51 1391 -17
rect 1425 -51 1464 -17
rect 1498 -51 1537 -17
rect 1571 -51 1610 -17
rect 1644 -51 1683 -17
rect 1717 -51 1756 -17
rect 1790 -51 1829 -17
rect 1863 -51 1902 -17
rect 1936 -51 1975 -17
rect 2009 -51 2048 -17
rect 2082 -51 2121 -17
rect 2155 -51 2194 -17
rect 2228 -51 2267 -17
rect 2301 -51 2340 -17
rect 2374 -51 2413 -17
rect 2447 -51 2486 -17
rect 2520 -51 2559 -17
rect 2593 -51 2631 -17
rect 2665 -51 2703 -17
rect 2737 -51 2775 -17
rect 2809 -51 2847 -17
rect 2881 -51 2919 -17
rect 2953 -51 2991 -17
rect 3025 -51 3063 -17
rect 3097 -51 3135 -17
rect 3169 -51 3202 -17
rect 65 -56 3202 -51
tri 3202 -56 3252 -6 nw
rect 65 -57 3181 -56
<< rmetal1 >>
rect 459 778 461 779
rect 497 778 499 779
rect 459 734 460 778
rect 498 734 499 778
rect 459 733 461 734
rect 497 733 499 734
rect 228 685 230 686
rect 266 685 268 686
rect 228 635 229 685
rect 267 635 268 685
rect 228 634 230 635
rect 266 634 268 635
rect 3244 665 3296 666
rect 3244 664 3245 665
rect 3295 664 3296 665
rect 3244 627 3245 628
rect 3295 627 3296 628
rect 3244 626 3296 627
rect 3165 599 3167 600
rect 3165 549 3166 599
rect 3165 548 3167 549
rect 3203 599 3205 600
rect 3204 549 3205 599
rect 3203 548 3205 549
rect 555 500 557 501
rect 593 500 595 501
rect 555 456 556 500
rect 594 456 595 500
rect 555 455 557 456
rect 593 455 595 456
rect 2852 425 2854 426
rect 2852 381 2853 425
rect 2852 380 2854 381
rect 2890 425 2892 426
rect 2891 381 2892 425
rect 2890 380 2892 381
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_0
timestamp 1707688321
transform -1 0 2944 0 1 380
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1707688321
transform 0 -1 3296 1 0 574
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1707688321
transform -1 0 3257 0 -1 600
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1707688321
transform -1 0 647 0 1 455
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_1
timestamp 1707688321
transform 1 0 407 0 1 733
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1707688321
transform 1 0 176 0 1 634
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_5595914180883  sky130_fd_pr__nfet_01v8__example_5595914180883_0
timestamp 1707688321
transform -1 0 2826 0 1 57
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_5595914180885  sky130_fd_pr__nfet_01v8__example_5595914180885_0
timestamp 1707688321
transform 1 0 1510 0 1 57
box -1 0 881 1
use sky130_fd_pr__nfet_01v8__example_5595914180886  sky130_fd_pr__nfet_01v8__example_5595914180886_0
timestamp 1707688321
transform -1 0 3138 0 1 57
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_5595914180887  sky130_fd_pr__nfet_01v8__example_5595914180887_0
timestamp 1707688321
transform 1 0 574 0 1 57
box -1 0 881 1
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_0
timestamp 1707688321
transform 1 0 281 0 1 57
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_1
timestamp 1707688321
transform 1 0 125 0 1 57
box -1 0 101 1
<< labels >>
flabel metal1 s 371 396 423 448 3 FreeSans 520 0 0 0 OUT
port 1 nsew
flabel metal1 s 309 733 361 779 3 FreeSans 520 0 0 0 IN1
port 2 nsew
flabel metal1 s 160 624 202 676 3 FreeSans 520 0 0 0 IN2
port 3 nsew
flabel metal1 s 149 92 201 144 3 FreeSans 520 0 0 0 VGND
port 4 nsew
<< properties >>
string GDS_END 70963580
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70943192
<< end >>
