magic
tech sky130B
magscale 1 2
timestamp 1707688321
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_5595914180851  sky130_fd_pr__hvdfl1sd__example_5595914180851_1
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 64843172
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64842246
<< end >>
