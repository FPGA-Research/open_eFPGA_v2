magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< locali >>
rect 179 1160 187 1194
rect 221 1160 259 1194
rect 293 1160 331 1194
rect 365 1160 403 1194
rect 437 1160 475 1194
rect 509 1160 517 1194
rect 179 20 187 54
rect 221 20 259 54
rect 293 20 331 54
rect 365 20 403 54
rect 437 20 475 54
rect 509 20 517 54
<< viali >>
rect 187 1160 221 1194
rect 259 1160 293 1194
rect 331 1160 365 1194
rect 403 1160 437 1194
rect 475 1160 509 1194
rect 187 20 221 54
rect 259 20 293 54
rect 331 20 365 54
rect 403 20 437 54
rect 475 20 509 54
<< obsli1 >>
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 159 98 193 1116
rect 245 98 279 1116
rect 331 98 365 1116
rect 417 98 451 1116
rect 503 98 537 1116
rect 614 1020 648 1058
rect 614 948 648 986
rect 614 876 648 914
rect 614 804 648 842
rect 614 732 648 770
rect 614 660 648 698
rect 614 588 648 626
rect 614 516 648 554
rect 614 444 648 482
rect 614 372 648 410
rect 614 300 648 338
rect 614 228 648 266
rect 614 122 648 194
<< obsli1c >>
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 614 1058 648 1092
rect 614 986 648 1020
rect 614 914 648 948
rect 614 842 648 876
rect 614 770 648 804
rect 614 698 648 732
rect 614 626 648 660
rect 614 554 648 588
rect 614 482 648 516
rect 614 410 648 444
rect 614 338 648 372
rect 614 266 648 300
rect 614 194 648 228
<< metal1 >>
rect 175 1194 521 1214
rect 175 1160 187 1194
rect 221 1160 259 1194
rect 293 1160 331 1194
rect 365 1160 403 1194
rect 437 1160 475 1194
rect 509 1160 521 1194
rect 175 1148 521 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 602 1092 660 1104
rect 602 1058 614 1092
rect 648 1058 660 1092
rect 602 1020 660 1058
rect 602 986 614 1020
rect 648 986 660 1020
rect 602 948 660 986
rect 602 914 614 948
rect 648 914 660 948
rect 602 876 660 914
rect 602 842 614 876
rect 648 842 660 876
rect 602 804 660 842
rect 602 770 614 804
rect 648 770 660 804
rect 602 732 660 770
rect 602 698 614 732
rect 648 698 660 732
rect 602 660 660 698
rect 602 626 614 660
rect 648 626 660 660
rect 602 588 660 626
rect 602 554 614 588
rect 648 554 660 588
rect 602 516 660 554
rect 602 482 614 516
rect 648 482 660 516
rect 602 444 660 482
rect 602 410 614 444
rect 648 410 660 444
rect 602 372 660 410
rect 602 338 614 372
rect 648 338 660 372
rect 602 300 660 338
rect 602 266 614 300
rect 648 266 660 300
rect 602 228 660 266
rect 602 194 614 228
rect 648 194 660 228
rect 602 110 660 194
rect 175 54 521 66
rect 175 20 187 54
rect 221 20 259 54
rect 293 20 331 54
rect 365 20 403 54
rect 437 20 475 54
rect 509 20 521 54
rect 175 0 521 20
<< obsm1 >>
rect 150 110 202 1104
rect 236 110 288 1104
rect 322 110 374 1104
rect 408 110 460 1104
rect 494 110 546 1104
<< metal2 >>
rect 10 632 686 1104
rect 10 110 686 582
<< labels >>
rlabel metal1 s 602 110 660 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 686 1104 6 DRAIN
port 2 nsew
rlabel viali s 475 1160 509 1194 6 GATE
port 3 nsew
rlabel viali s 475 20 509 54 6 GATE
port 3 nsew
rlabel viali s 403 1160 437 1194 6 GATE
port 3 nsew
rlabel viali s 403 20 437 54 6 GATE
port 3 nsew
rlabel viali s 331 1160 365 1194 6 GATE
port 3 nsew
rlabel viali s 331 20 365 54 6 GATE
port 3 nsew
rlabel viali s 259 1160 293 1194 6 GATE
port 3 nsew
rlabel viali s 259 20 293 54 6 GATE
port 3 nsew
rlabel viali s 187 1160 221 1194 6 GATE
port 3 nsew
rlabel viali s 187 20 221 54 6 GATE
port 3 nsew
rlabel locali s 179 1160 517 1194 6 GATE
port 3 nsew
rlabel locali s 179 20 517 54 6 GATE
port 3 nsew
rlabel metal1 s 175 1148 521 1214 6 GATE
port 3 nsew
rlabel metal1 s 175 0 521 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 686 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 696 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9432272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9410370
<< end >>
