magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -95 -26 179 110
<< mvnmos >>
rect 0 0 100 84
<< mvndiff >>
rect -69 46 0 84
rect -69 12 -61 46
rect -27 12 0 46
rect -69 0 0 12
rect 100 46 153 84
rect 100 12 111 46
rect 145 12 153 46
rect 100 0 153 12
<< mvndiffc >>
rect -61 12 -27 46
rect 111 12 145 46
<< poly >>
rect 0 84 100 110
rect 0 -26 100 0
<< locali >>
rect -61 46 -27 62
rect -61 -4 -27 12
rect 111 46 145 62
rect 111 -4 145 12
use DFL1sd_CDNS_52468879185271  DFL1sd_CDNS_52468879185271_0
timestamp 1707688321
transform -1 0 -16 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185271  DFL1sd_CDNS_52468879185271_1
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -44 29 -44 29 0 FreeSans 300 0 0 0 S
flabel comment s 128 29 128 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 70896746
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 70895796
<< end >>
