magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 5111 333 5265 587
rect 6757 333 6911 587
rect 5111 227 6911 333
rect 7311 227 7417 589
rect 8099 227 8205 589
<< pwell >>
rect 4897 1469 7222 1555
rect 4897 1085 5547 1469
rect 6450 1085 7222 1469
rect 4897 167 5051 1085
rect 7000 931 7222 1085
rect 7000 677 7407 931
rect 8109 677 8195 931
rect 7000 589 7459 677
rect 8057 589 8195 677
rect 7000 167 7222 589
rect 4897 13 7222 167
<< psubdiff >>
rect 4923 1505 5101 1529
rect 4957 1471 4991 1505
rect 5025 1495 5101 1505
rect 5135 1495 5170 1529
rect 5204 1495 5239 1529
rect 5273 1495 5308 1529
rect 5342 1495 5377 1529
rect 5411 1495 5511 1529
rect 5545 1495 5584 1529
rect 5618 1495 5656 1529
rect 5690 1495 5728 1529
rect 5762 1495 5800 1529
rect 5834 1495 5868 1529
rect 5902 1495 5936 1529
rect 5970 1495 6008 1529
rect 6042 1495 6080 1529
rect 6114 1495 6148 1529
rect 6182 1495 6216 1529
rect 6250 1495 6288 1529
rect 6322 1495 6356 1529
rect 6390 1495 6424 1529
rect 6458 1495 6568 1529
rect 6602 1495 6646 1529
rect 6680 1495 6724 1529
rect 6758 1495 6802 1529
rect 6836 1495 6880 1529
rect 6914 1495 6958 1529
rect 6992 1505 7196 1529
rect 6992 1495 7026 1505
rect 5025 1471 5521 1495
rect 4923 1461 5521 1471
rect 6476 1471 7026 1495
rect 7060 1471 7094 1505
rect 7128 1471 7162 1505
rect 4923 1436 5101 1461
rect 4957 1402 4991 1436
rect 5025 1427 5101 1436
rect 5135 1427 5170 1461
rect 5204 1427 5239 1461
rect 5273 1427 5308 1461
rect 5342 1427 5377 1461
rect 5411 1427 5521 1461
rect 5025 1412 5521 1427
rect 5025 1402 5487 1412
rect 4923 1393 5487 1402
rect 4923 1367 5101 1393
rect 4957 1333 4991 1367
rect 5025 1359 5101 1367
rect 5135 1359 5170 1393
rect 5204 1359 5239 1393
rect 5273 1359 5308 1393
rect 5342 1359 5377 1393
rect 5411 1378 5487 1393
rect 6476 1461 7196 1471
rect 6476 1427 6568 1461
rect 6602 1427 6646 1461
rect 6680 1427 6724 1461
rect 6758 1427 6802 1461
rect 6836 1427 6880 1461
rect 6914 1427 6958 1461
rect 6992 1436 7196 1461
rect 6992 1427 7026 1436
rect 6476 1424 7026 1427
rect 6510 1402 7026 1424
rect 7060 1402 7094 1436
rect 7128 1402 7162 1436
rect 6510 1393 7196 1402
rect 6510 1390 6568 1393
rect 5411 1359 5521 1378
rect 5025 1333 5521 1359
rect 4923 1331 5521 1333
rect 4923 1325 5487 1331
rect 4923 1298 5101 1325
rect 4957 1264 4991 1298
rect 5025 1291 5101 1298
rect 5135 1291 5170 1325
rect 5204 1291 5239 1325
rect 5273 1291 5308 1325
rect 5342 1291 5377 1325
rect 5411 1297 5487 1325
rect 5411 1291 5521 1297
rect 5025 1264 5521 1291
rect 4923 1250 5521 1264
rect 4923 1229 5487 1250
rect 4957 1195 4991 1229
rect 5025 1216 5487 1229
rect 5025 1195 5521 1216
rect 4923 1169 5521 1195
rect 4923 1160 5487 1169
rect 4957 1126 4991 1160
rect 5025 1145 5487 1160
rect 5025 1126 5323 1145
rect 4923 1111 5323 1126
rect 5357 1111 5393 1145
rect 5427 1135 5487 1145
rect 5427 1111 5521 1135
rect 6476 1359 6568 1390
rect 6602 1359 6646 1393
rect 6680 1359 6724 1393
rect 6758 1359 6802 1393
rect 6836 1359 6880 1393
rect 6914 1359 6958 1393
rect 6992 1367 7196 1393
rect 6992 1359 7026 1367
rect 6476 1343 7026 1359
rect 6510 1333 7026 1343
rect 7060 1333 7094 1367
rect 7128 1333 7162 1367
rect 6510 1325 7196 1333
rect 6510 1309 6568 1325
rect 6476 1291 6568 1309
rect 6602 1291 6646 1325
rect 6680 1291 6724 1325
rect 6758 1291 6802 1325
rect 6836 1291 6880 1325
rect 6914 1291 6958 1325
rect 6992 1298 7196 1325
rect 6992 1291 7026 1298
rect 6476 1264 7026 1291
rect 7060 1264 7094 1298
rect 7128 1264 7162 1298
rect 6476 1262 7196 1264
rect 6510 1229 7196 1262
rect 6510 1228 7026 1229
rect 6476 1195 7026 1228
rect 7060 1195 7094 1229
rect 7128 1195 7162 1229
rect 6476 1160 7196 1195
rect 6476 1145 7026 1160
rect 6476 1111 6500 1145
rect 6534 1111 6579 1145
rect 6613 1111 6657 1145
rect 6691 1126 7026 1145
rect 7060 1126 7094 1160
rect 7128 1126 7162 1160
rect 6691 1111 7196 1126
rect 4923 1091 5025 1111
rect 4957 1057 4991 1091
rect 4923 1022 5025 1057
rect 4957 988 4991 1022
rect 4923 953 5025 988
rect 4957 919 4991 953
rect 4923 884 5025 919
rect 4957 850 4991 884
rect 4923 815 5025 850
rect 4957 781 4991 815
rect 4923 746 5025 781
rect 4957 712 4991 746
rect 7026 1091 7196 1111
rect 7060 1057 7094 1091
rect 7128 1057 7162 1091
rect 7026 1022 7196 1057
rect 7060 988 7094 1022
rect 7128 988 7162 1022
rect 7026 953 7196 988
rect 7060 919 7094 953
rect 7128 919 7162 953
rect 7026 884 7196 919
rect 7060 850 7094 884
rect 7128 850 7162 884
rect 7026 815 7196 850
rect 7060 781 7094 815
rect 7128 781 7162 815
rect 7026 746 7196 781
rect 4923 677 5025 712
rect 4957 643 4991 677
rect 4923 608 5025 643
rect 4957 574 4991 608
rect 7060 712 7094 746
rect 7128 712 7162 746
rect 7026 677 7196 712
rect 7060 643 7094 677
rect 7128 643 7162 677
rect 7026 608 7196 643
rect 7347 881 7381 905
rect 7347 812 7381 847
rect 7347 743 7381 778
rect 7347 673 7381 709
rect 8135 881 8169 905
rect 8135 812 8169 847
rect 8135 743 8169 778
rect 8135 673 8169 709
rect 7381 639 7407 651
rect 7347 615 7407 639
rect 8109 639 8135 651
rect 8109 615 8169 639
rect 4923 538 5025 574
rect 4957 504 4991 538
rect 4923 468 5025 504
rect 4957 434 4991 468
rect 4923 398 5025 434
rect 4957 364 4991 398
rect 4923 328 5025 364
rect 4957 294 4991 328
rect 7060 574 7094 608
rect 7128 574 7162 608
rect 7026 538 7196 574
rect 7060 504 7094 538
rect 7128 504 7162 538
rect 7026 468 7196 504
rect 7060 434 7094 468
rect 7128 434 7162 468
rect 7026 398 7196 434
rect 7060 364 7094 398
rect 7128 364 7162 398
rect 7026 328 7196 364
rect 4923 258 5025 294
rect 7060 294 7094 328
rect 7128 294 7162 328
rect 4957 224 4991 258
rect 4923 141 5025 224
rect 7026 258 7196 294
rect 7060 224 7094 258
rect 7128 224 7162 258
rect 7026 141 7196 224
rect 4923 39 4947 141
rect 6137 107 6172 141
rect 6206 107 6241 141
rect 6275 107 6310 141
rect 6344 107 6379 141
rect 6413 107 6448 141
rect 6482 107 6517 141
rect 6551 107 6586 141
rect 6620 107 6655 141
rect 6689 107 6724 141
rect 6758 107 6793 141
rect 6827 107 6862 141
rect 6896 107 6931 141
rect 6965 107 7000 141
rect 7034 107 7069 141
rect 7103 107 7138 141
rect 7172 107 7196 141
rect 6137 73 7196 107
rect 6137 39 6172 73
rect 6206 39 6241 73
rect 6275 39 6310 73
rect 6344 39 6379 73
rect 6413 39 6448 73
rect 6482 39 6517 73
rect 6551 39 6586 73
rect 6620 39 6655 73
rect 6689 39 6724 73
rect 6758 39 6793 73
rect 6827 39 6862 73
rect 6896 39 6931 73
rect 6965 39 7000 73
rect 7034 39 7069 73
rect 7103 39 7138 73
rect 7172 39 7196 73
<< nsubdiff >>
rect 7407 615 7433 651
rect 8083 615 8109 651
rect 5147 263 5171 297
rect 5205 263 5263 297
rect 5297 263 5333 297
rect 5367 263 5403 297
rect 5437 263 5473 297
rect 5507 263 5543 297
rect 5577 263 5613 297
rect 5647 263 5683 297
rect 5717 263 5753 297
rect 5787 263 5823 297
rect 5857 263 5893 297
rect 5927 263 5963 297
rect 5997 263 6033 297
rect 6067 263 6103 297
rect 6137 263 6173 297
rect 6207 263 6242 297
rect 6276 263 6311 297
rect 6345 263 6380 297
rect 6414 263 6449 297
rect 6483 263 6518 297
rect 6552 263 6587 297
rect 6621 263 6656 297
rect 6690 263 6725 297
rect 6759 263 6817 297
rect 6851 263 6875 297
rect 7347 529 7433 553
rect 7381 517 7433 529
rect 8083 529 8169 553
rect 8083 517 8135 529
rect 7347 460 7381 495
rect 7347 391 7381 426
rect 7347 321 7381 357
rect 7347 263 7381 287
rect 8135 460 8169 495
rect 8135 391 8169 426
rect 8135 321 8169 357
rect 8135 263 8169 287
<< psubdiffcont >>
rect 4923 1471 4957 1505
rect 4991 1471 5025 1505
rect 5101 1495 5135 1529
rect 5170 1495 5204 1529
rect 5239 1495 5273 1529
rect 5308 1495 5342 1529
rect 5377 1495 5411 1529
rect 5511 1495 5545 1529
rect 5584 1495 5618 1529
rect 5656 1495 5690 1529
rect 5728 1495 5762 1529
rect 5800 1495 5834 1529
rect 5868 1495 5902 1529
rect 5936 1495 5970 1529
rect 6008 1495 6042 1529
rect 6080 1495 6114 1529
rect 6148 1495 6182 1529
rect 6216 1495 6250 1529
rect 6288 1495 6322 1529
rect 6356 1495 6390 1529
rect 6424 1495 6458 1529
rect 6568 1495 6602 1529
rect 6646 1495 6680 1529
rect 6724 1495 6758 1529
rect 6802 1495 6836 1529
rect 6880 1495 6914 1529
rect 6958 1495 6992 1529
rect 7026 1471 7060 1505
rect 7094 1471 7128 1505
rect 7162 1471 7196 1505
rect 4923 1402 4957 1436
rect 4991 1402 5025 1436
rect 5101 1427 5135 1461
rect 5170 1427 5204 1461
rect 5239 1427 5273 1461
rect 5308 1427 5342 1461
rect 5377 1427 5411 1461
rect 4923 1333 4957 1367
rect 4991 1333 5025 1367
rect 5101 1359 5135 1393
rect 5170 1359 5204 1393
rect 5239 1359 5273 1393
rect 5308 1359 5342 1393
rect 5377 1359 5411 1393
rect 5487 1378 5521 1412
rect 6568 1427 6602 1461
rect 6646 1427 6680 1461
rect 6724 1427 6758 1461
rect 6802 1427 6836 1461
rect 6880 1427 6914 1461
rect 6958 1427 6992 1461
rect 6476 1390 6510 1424
rect 7026 1402 7060 1436
rect 7094 1402 7128 1436
rect 7162 1402 7196 1436
rect 4923 1264 4957 1298
rect 4991 1264 5025 1298
rect 5101 1291 5135 1325
rect 5170 1291 5204 1325
rect 5239 1291 5273 1325
rect 5308 1291 5342 1325
rect 5377 1291 5411 1325
rect 5487 1297 5521 1331
rect 4923 1195 4957 1229
rect 4991 1195 5025 1229
rect 5487 1216 5521 1250
rect 4923 1126 4957 1160
rect 4991 1126 5025 1160
rect 5323 1111 5357 1145
rect 5393 1111 5427 1145
rect 5487 1135 5521 1169
rect 6568 1359 6602 1393
rect 6646 1359 6680 1393
rect 6724 1359 6758 1393
rect 6802 1359 6836 1393
rect 6880 1359 6914 1393
rect 6958 1359 6992 1393
rect 6476 1309 6510 1343
rect 7026 1333 7060 1367
rect 7094 1333 7128 1367
rect 7162 1333 7196 1367
rect 6568 1291 6602 1325
rect 6646 1291 6680 1325
rect 6724 1291 6758 1325
rect 6802 1291 6836 1325
rect 6880 1291 6914 1325
rect 6958 1291 6992 1325
rect 7026 1264 7060 1298
rect 7094 1264 7128 1298
rect 7162 1264 7196 1298
rect 6476 1228 6510 1262
rect 7026 1195 7060 1229
rect 7094 1195 7128 1229
rect 7162 1195 7196 1229
rect 6500 1111 6534 1145
rect 6579 1111 6613 1145
rect 6657 1111 6691 1145
rect 7026 1126 7060 1160
rect 7094 1126 7128 1160
rect 7162 1126 7196 1160
rect 4923 1057 4957 1091
rect 4991 1057 5025 1091
rect 4923 988 4957 1022
rect 4991 988 5025 1022
rect 4923 919 4957 953
rect 4991 919 5025 953
rect 4923 850 4957 884
rect 4991 850 5025 884
rect 4923 781 4957 815
rect 4991 781 5025 815
rect 4923 712 4957 746
rect 4991 712 5025 746
rect 7026 1057 7060 1091
rect 7094 1057 7128 1091
rect 7162 1057 7196 1091
rect 7026 988 7060 1022
rect 7094 988 7128 1022
rect 7162 988 7196 1022
rect 7026 919 7060 953
rect 7094 919 7128 953
rect 7162 919 7196 953
rect 7026 850 7060 884
rect 7094 850 7128 884
rect 7162 850 7196 884
rect 7026 781 7060 815
rect 7094 781 7128 815
rect 7162 781 7196 815
rect 4923 643 4957 677
rect 4991 643 5025 677
rect 4923 574 4957 608
rect 4991 574 5025 608
rect 7026 712 7060 746
rect 7094 712 7128 746
rect 7162 712 7196 746
rect 7026 643 7060 677
rect 7094 643 7128 677
rect 7162 643 7196 677
rect 7347 847 7381 881
rect 7347 778 7381 812
rect 7347 709 7381 743
rect 7347 639 7381 673
rect 8135 847 8169 881
rect 8135 778 8169 812
rect 8135 709 8169 743
rect 8135 639 8169 673
rect 4923 504 4957 538
rect 4991 504 5025 538
rect 4923 434 4957 468
rect 4991 434 5025 468
rect 4923 364 4957 398
rect 4991 364 5025 398
rect 4923 294 4957 328
rect 4991 294 5025 328
rect 7026 574 7060 608
rect 7094 574 7128 608
rect 7162 574 7196 608
rect 7026 504 7060 538
rect 7094 504 7128 538
rect 7162 504 7196 538
rect 7026 434 7060 468
rect 7094 434 7128 468
rect 7162 434 7196 468
rect 7026 364 7060 398
rect 7094 364 7128 398
rect 7162 364 7196 398
rect 7026 294 7060 328
rect 7094 294 7128 328
rect 7162 294 7196 328
rect 4923 224 4957 258
rect 4991 224 5025 258
rect 7026 224 7060 258
rect 7094 224 7128 258
rect 7162 224 7196 258
rect 4947 39 6137 141
rect 6172 107 6206 141
rect 6241 107 6275 141
rect 6310 107 6344 141
rect 6379 107 6413 141
rect 6448 107 6482 141
rect 6517 107 6551 141
rect 6586 107 6620 141
rect 6655 107 6689 141
rect 6724 107 6758 141
rect 6793 107 6827 141
rect 6862 107 6896 141
rect 6931 107 6965 141
rect 7000 107 7034 141
rect 7069 107 7103 141
rect 7138 107 7172 141
rect 6172 39 6206 73
rect 6241 39 6275 73
rect 6310 39 6344 73
rect 6379 39 6413 73
rect 6448 39 6482 73
rect 6517 39 6551 73
rect 6586 39 6620 73
rect 6655 39 6689 73
rect 6724 39 6758 73
rect 6793 39 6827 73
rect 6862 39 6896 73
rect 6931 39 6965 73
rect 7000 39 7034 73
rect 7069 39 7103 73
rect 7138 39 7172 73
<< nsubdiffcont >>
rect 5171 263 5205 297
rect 5263 263 5297 297
rect 5333 263 5367 297
rect 5403 263 5437 297
rect 5473 263 5507 297
rect 5543 263 5577 297
rect 5613 263 5647 297
rect 5683 263 5717 297
rect 5753 263 5787 297
rect 5823 263 5857 297
rect 5893 263 5927 297
rect 5963 263 5997 297
rect 6033 263 6067 297
rect 6103 263 6137 297
rect 6173 263 6207 297
rect 6242 263 6276 297
rect 6311 263 6345 297
rect 6380 263 6414 297
rect 6449 263 6483 297
rect 6518 263 6552 297
rect 6587 263 6621 297
rect 6656 263 6690 297
rect 6725 263 6759 297
rect 6817 263 6851 297
rect 7347 495 7381 529
rect 7347 426 7381 460
rect 7347 357 7381 391
rect 7347 287 7381 321
rect 8135 495 8169 529
rect 8135 426 8169 460
rect 8135 357 8169 391
rect 8135 287 8169 321
<< poly >>
rect -352 1357 -14 1373
rect -352 1323 -336 1357
rect -302 1323 -268 1357
rect -234 1323 -200 1357
rect -166 1323 -132 1357
rect -98 1323 -64 1357
rect -30 1323 -14 1357
rect -352 1307 -14 1323
rect 5766 1446 5900 1462
rect 5766 1412 5782 1446
rect 5816 1412 5850 1446
rect 5884 1412 5900 1446
rect 5766 1389 5900 1412
rect 6118 1445 6252 1461
rect 6118 1411 6134 1445
rect 6168 1411 6202 1445
rect 6236 1411 6252 1445
rect 6118 1388 6252 1411
rect -346 1301 -226 1307
rect -170 1301 -50 1307
rect -346 939 -50 1053
rect -346 905 -299 939
rect -265 905 -123 939
rect -89 934 -50 939
rect -89 905 278 934
rect -346 871 278 905
rect -346 837 -299 871
rect -265 837 -123 871
rect -89 837 278 871
rect -346 749 278 837
rect 5216 695 5416 745
rect 6606 695 6806 745
rect 5216 679 5928 695
rect 5216 645 5511 679
rect 5545 645 5579 679
rect 5613 645 5647 679
rect 5681 645 5715 679
rect 5749 645 5783 679
rect 5817 645 5851 679
rect 5885 645 5928 679
rect 5216 629 5928 645
rect 5216 583 5672 629
rect 5216 576 5416 583
rect 5472 576 5672 583
rect 5728 577 5928 629
rect 6094 679 6806 695
rect 6094 645 6205 679
rect 6239 645 6273 679
rect 6307 645 6341 679
rect 6375 645 6409 679
rect 6443 645 6477 679
rect 6511 645 6806 679
rect 6094 629 6806 645
rect 6094 576 6294 629
rect 6350 577 6806 629
rect 6606 576 6806 577
rect -346 91 -226 97
rect -170 91 -50 97
rect 6 91 126 97
rect 182 91 302 97
<< polycont >>
rect -336 1323 -302 1357
rect -268 1323 -234 1357
rect -200 1323 -166 1357
rect -132 1323 -98 1357
rect -64 1323 -30 1357
rect 5782 1412 5816 1446
rect 5850 1412 5884 1446
rect 6134 1411 6168 1445
rect 6202 1411 6236 1445
rect -299 905 -265 939
rect -123 905 -89 939
rect -299 837 -265 871
rect -123 837 -89 871
rect 5511 645 5545 679
rect 5579 645 5613 679
rect 5647 645 5681 679
rect 5715 645 5749 679
rect 5783 645 5817 679
rect 5851 645 5885 679
rect 6205 645 6239 679
rect 6273 645 6307 679
rect 6341 645 6375 679
rect 6409 645 6443 679
rect 6477 645 6511 679
<< locali >>
rect 4923 1505 5101 1529
rect 4957 1471 4991 1505
rect 5025 1495 5101 1505
rect 5135 1495 5170 1529
rect 5204 1495 5239 1529
rect 5273 1495 5308 1529
rect 5342 1495 5377 1529
rect 5411 1495 5511 1529
rect 5545 1495 5584 1529
rect 5618 1495 5656 1529
rect 5690 1495 5728 1529
rect 5762 1495 5800 1529
rect 5834 1495 5868 1529
rect 5902 1495 5936 1529
rect 5970 1495 6008 1529
rect 6042 1495 6080 1529
rect 6114 1495 6148 1529
rect 6182 1495 6216 1529
rect 6250 1495 6288 1529
rect 6322 1495 6356 1529
rect 6390 1495 6424 1529
rect 6458 1495 6568 1529
rect 6602 1495 6646 1529
rect 6680 1495 6724 1529
rect 6758 1495 6802 1529
rect 6836 1495 6880 1529
rect 6914 1495 6958 1529
rect 6992 1505 7196 1529
rect 6992 1495 7026 1505
rect 5025 1471 5601 1495
rect 4923 1461 5601 1471
rect 4923 1436 5101 1461
rect -2001 1381 -1963 1415
rect 863 1381 901 1415
rect -2035 1361 -1933 1381
rect -1239 1307 -1165 1373
rect -887 1307 -813 1373
rect -336 1357 -30 1373
rect -302 1323 -268 1357
rect -234 1323 -200 1357
rect -166 1323 -132 1357
rect -98 1323 -64 1357
rect -336 1307 -30 1323
rect 723 1307 761 1341
rect 829 1307 935 1381
rect 4957 1402 4991 1436
rect 5025 1427 5101 1436
rect 5135 1427 5170 1461
rect 5204 1427 5239 1461
rect 5273 1427 5308 1461
rect 5342 1427 5377 1461
rect 5411 1427 5601 1461
rect 6421 1471 7026 1495
rect 7060 1471 7094 1505
rect 7128 1471 7162 1505
rect 6421 1461 7196 1471
rect 5025 1412 5601 1427
rect 5766 1412 5782 1446
rect 5816 1412 5850 1446
rect 5884 1412 5900 1446
rect 6118 1415 6134 1445
rect 5025 1402 5487 1412
rect 4923 1393 5487 1402
rect 4923 1367 5101 1393
rect 1039 1307 1077 1341
rect 4957 1333 4991 1367
rect 5025 1359 5101 1367
rect 5135 1359 5170 1393
rect 5204 1359 5239 1393
rect 5273 1359 5308 1393
rect 5342 1359 5377 1393
rect 5411 1378 5487 1393
rect 5521 1378 5601 1412
rect 5411 1359 5601 1378
rect 5025 1333 5601 1359
rect 4923 1331 5601 1333
rect 4923 1325 5487 1331
rect -391 1169 -357 1207
rect -391 1097 -357 1135
rect -323 939 -249 1307
rect -1975 881 -1937 915
rect -323 905 -299 939
rect -265 905 -249 939
rect -1483 868 -1445 902
rect -744 868 -706 902
rect -481 868 -443 902
rect -323 871 -249 905
rect -323 837 -299 871
rect -265 837 -249 871
rect -391 643 -357 681
rect -391 571 -357 609
rect -601 387 -567 425
rect -1660 274 -1622 308
rect -1500 218 -1466 256
rect -1219 218 -1185 256
rect -867 218 -833 256
rect -323 91 -249 837
rect -215 727 -181 1071
rect -147 939 -73 1307
rect 733 1278 795 1307
rect 4923 1298 5101 1325
rect 733 1244 809 1278
rect 4957 1264 4991 1298
rect 5025 1291 5101 1298
rect 5135 1291 5170 1325
rect 5204 1291 5239 1325
rect 5273 1291 5308 1325
rect 5342 1291 5377 1325
rect 5411 1297 5487 1325
rect 5521 1297 5601 1331
rect 5778 1341 5884 1412
rect 6118 1411 6130 1415
rect 6168 1411 6202 1445
rect 6236 1411 6252 1445
rect 6421 1427 6568 1461
rect 6602 1427 6646 1461
rect 6680 1427 6724 1461
rect 6758 1427 6802 1461
rect 6836 1427 6880 1461
rect 6914 1427 6958 1461
rect 6992 1436 7196 1461
rect 6992 1427 7026 1436
rect 6421 1424 7026 1427
rect 6164 1381 6202 1411
rect 6421 1390 6476 1424
rect 6510 1402 7026 1424
rect 7060 1402 7094 1436
rect 7128 1402 7162 1436
rect 6510 1393 7196 1402
rect 6510 1390 6568 1393
rect 5812 1307 5850 1341
rect 6421 1359 6568 1390
rect 6602 1359 6646 1393
rect 6680 1359 6724 1393
rect 6758 1359 6802 1393
rect 6836 1359 6880 1393
rect 6914 1359 6958 1393
rect 6992 1367 7196 1393
rect 6992 1359 7026 1367
rect 6421 1343 7026 1359
rect 6421 1309 6476 1343
rect 6510 1333 7026 1343
rect 7060 1333 7094 1367
rect 7128 1333 7162 1367
rect 6510 1325 7196 1333
rect 6510 1309 6568 1325
rect 5411 1291 5601 1297
rect 5025 1264 5601 1291
rect 4923 1250 5601 1264
rect -39 1169 -5 1207
rect -39 1097 -5 1135
rect -147 905 -123 939
rect -89 905 -73 939
rect -147 871 -73 905
rect -147 837 -123 871
rect -89 837 -73 871
rect -215 387 -181 425
rect -147 91 -73 837
rect -39 643 -5 681
rect -39 571 -5 609
rect 313 643 347 681
rect 313 571 347 609
rect 137 387 171 425
rect 489 155 523 193
rect 733 124 795 1244
rect 4923 1229 5487 1250
rect 4957 1195 4991 1229
rect 5025 1216 5487 1229
rect 5521 1216 5601 1250
rect 6421 1291 6568 1309
rect 6602 1291 6646 1325
rect 6680 1291 6724 1325
rect 6758 1291 6802 1325
rect 6836 1291 6880 1325
rect 6914 1291 6958 1325
rect 6992 1298 7196 1325
rect 6992 1291 7026 1298
rect 6421 1264 7026 1291
rect 7060 1264 7094 1298
rect 7128 1264 7162 1298
rect 6421 1262 7196 1264
rect 5025 1195 5601 1216
rect 4610 1119 4644 1157
rect 4923 1190 5601 1195
rect 4923 1160 4942 1190
rect 4976 1160 5018 1190
rect 4976 1156 4991 1160
rect 5052 1156 5094 1190
rect 5128 1156 5170 1190
rect 5204 1156 5246 1190
rect 5280 1156 5322 1190
rect 5356 1156 5398 1190
rect 5432 1156 5473 1190
rect 5507 1169 5548 1190
rect 5521 1156 5548 1169
rect 5582 1156 5601 1190
rect 4957 1126 4991 1156
rect 5025 1145 5487 1156
rect 5025 1126 5323 1145
rect 4923 1118 5323 1126
rect 4923 1091 4942 1118
rect 4976 1091 5018 1118
rect 4976 1084 4991 1091
rect 5052 1084 5094 1118
rect 5128 1084 5170 1118
rect 5204 1084 5246 1118
rect 5280 1084 5322 1118
rect 5357 1111 5393 1145
rect 5427 1135 5487 1145
rect 5521 1135 5601 1156
rect 5427 1118 5601 1135
rect 5356 1084 5398 1111
rect 5432 1084 5473 1118
rect 5507 1084 5548 1118
rect 5582 1084 5601 1118
rect 1655 1016 1689 1063
rect 4957 1057 4991 1084
rect 5025 1057 5601 1084
rect 5683 1169 5717 1207
rect 5683 1097 5717 1135
rect 6305 1169 6339 1207
rect 6305 1097 6339 1135
rect 6421 1228 6476 1262
rect 6510 1229 7196 1262
rect 6510 1228 7026 1229
rect 6421 1199 7026 1228
rect 6421 1165 6440 1199
rect 6474 1165 6519 1199
rect 6553 1165 6597 1199
rect 6631 1165 6675 1199
rect 6709 1165 6753 1199
rect 6787 1165 6831 1199
rect 6865 1165 6909 1199
rect 6943 1165 6987 1199
rect 7021 1195 7026 1199
rect 7060 1199 7094 1229
rect 7128 1199 7162 1229
rect 7060 1195 7065 1199
rect 7128 1195 7143 1199
rect 7021 1165 7065 1195
rect 7099 1165 7143 1195
rect 7177 1165 7196 1195
rect 6421 1160 7196 1165
rect 6421 1145 7026 1160
rect 6421 1127 6500 1145
rect 6534 1127 6579 1145
rect 6613 1127 6657 1145
rect 6691 1127 7026 1145
rect 6421 1093 6440 1127
rect 6474 1111 6500 1127
rect 6553 1111 6579 1127
rect 6631 1111 6657 1127
rect 6474 1093 6519 1111
rect 6553 1093 6597 1111
rect 6631 1093 6675 1111
rect 6709 1093 6753 1127
rect 6787 1093 6831 1127
rect 6865 1093 6909 1127
rect 6943 1093 6987 1127
rect 7021 1126 7026 1127
rect 7060 1127 7094 1160
rect 7128 1127 7162 1160
rect 7060 1126 7065 1127
rect 7128 1126 7143 1127
rect 7021 1093 7065 1126
rect 7099 1093 7143 1126
rect 7177 1093 7196 1126
rect 6421 1091 7196 1093
rect 4923 1038 5601 1057
rect 4923 1022 4940 1038
rect 4974 1022 5012 1038
rect 4644 983 4682 1017
rect 4974 1004 4991 1022
rect 5046 1004 5084 1038
rect 5118 1004 5156 1038
rect 5190 1023 5601 1038
rect 5190 1017 5345 1023
rect 5190 1004 5239 1017
rect 4957 988 4991 1004
rect 5025 988 5239 1004
rect 4923 983 5239 988
rect 5273 983 5311 1017
rect 5495 1017 5601 1023
rect 5529 983 5567 1017
rect 6421 1057 7026 1091
rect 7060 1057 7094 1091
rect 7128 1057 7162 1091
rect 6421 1033 7196 1057
rect 6421 1017 6527 1033
rect 6455 983 6493 1017
rect 6677 1022 7196 1033
rect 6677 1017 7026 1022
rect 6711 983 6749 1017
rect 6783 1011 7026 1017
rect 6783 983 7022 1011
rect 7060 988 7094 1022
rect 7128 988 7162 1022
rect 4923 953 5205 983
rect 6677 977 7022 983
rect 7056 977 7094 988
rect 7128 977 7166 988
rect 4957 919 4991 953
rect 5025 919 5205 953
rect 4923 906 5205 919
rect 6817 953 7196 977
rect 6817 919 7026 953
rect 7060 919 7094 953
rect 7128 919 7162 953
rect 6817 907 7196 919
rect 4923 884 5171 906
rect 4957 850 4991 884
rect 5025 850 5171 884
rect 6605 863 6643 897
rect 6849 884 7196 907
rect 4923 815 5171 850
rect 4957 781 4991 815
rect 5025 781 5171 815
rect 4923 773 5171 781
rect 6849 850 7026 884
rect 7060 850 7094 884
rect 7128 850 7162 884
rect 6849 815 7196 850
rect 6849 781 7026 815
rect 7060 781 7094 815
rect 7128 781 7162 815
rect 6849 773 7196 781
rect 4923 746 5025 773
rect 4957 712 4991 746
rect 4923 677 5025 712
rect 4957 643 4991 677
rect 4923 608 5025 643
rect 4957 574 4991 608
rect 4923 538 5025 574
rect 4957 504 4991 538
rect 4923 468 5025 504
rect 4957 434 4991 468
rect 4923 398 5025 434
rect 4957 364 4991 398
rect 5171 486 5205 524
rect 5427 504 5461 773
rect 5939 753 5973 759
rect 5943 719 5981 753
rect 5495 645 5511 679
rect 5545 645 5579 679
rect 5613 645 5647 679
rect 5681 645 5715 679
rect 5761 645 5783 679
rect 5833 645 5851 679
rect 5885 645 5901 679
rect 5939 529 5973 719
rect 6049 679 6083 771
rect 6047 645 6085 679
rect 6189 645 6193 679
rect 6239 645 6265 679
rect 6307 645 6341 679
rect 6375 645 6409 679
rect 6443 645 6477 679
rect 6511 645 6527 679
rect 6049 549 6083 645
rect 5171 414 5205 452
rect 5683 486 5717 524
rect 5683 414 5717 452
rect 6561 549 6595 773
rect 7026 746 7196 773
rect 7060 712 7094 746
rect 7128 712 7162 746
rect 7026 677 7196 712
rect 7060 643 7094 677
rect 7128 643 7162 677
rect 7026 608 7196 643
rect 7060 574 7094 608
rect 7128 574 7162 608
rect 7347 903 7381 905
rect 7525 903 7559 941
rect 8135 903 8169 905
rect 7347 881 7491 903
rect 7381 847 7491 881
rect 8025 881 8169 903
rect 7347 812 7491 847
rect 7381 778 7491 812
rect 7347 743 7491 778
rect 7381 709 7491 743
rect 7347 673 7491 709
rect 7381 667 7491 673
rect 8025 847 8135 881
rect 8025 812 8169 847
rect 8025 778 8135 812
rect 8025 743 8169 778
rect 8025 709 8135 743
rect 8025 673 8169 709
rect 8025 667 8135 673
rect 7381 639 7479 667
rect 7347 638 7479 639
rect 7381 604 7479 638
rect 7347 601 7479 604
rect 8053 639 8135 667
rect 8053 638 8169 639
rect 8053 604 8135 638
rect 8053 601 8169 604
rect 6305 486 6339 524
rect 6305 414 6339 452
rect 6817 486 6851 524
rect 6817 414 6851 452
rect 7026 538 7196 574
rect 7060 504 7094 538
rect 7128 504 7162 538
rect 7026 468 7196 504
rect 7060 434 7094 468
rect 7128 434 7162 468
rect 7026 398 7196 434
rect 4923 328 5025 364
rect 4957 294 4991 328
rect 7060 364 7094 398
rect 7128 364 7162 398
rect 7026 328 7196 364
rect 4923 258 5025 294
rect 5155 263 5171 297
rect 5205 263 5263 297
rect 5297 263 5333 297
rect 5367 263 5403 297
rect 5437 263 5473 297
rect 5507 263 5543 297
rect 5577 263 5613 297
rect 5647 263 5683 297
rect 5717 263 5753 297
rect 5787 263 5823 297
rect 5857 263 5893 297
rect 5927 263 5963 297
rect 5997 263 6033 297
rect 6067 263 6103 297
rect 6137 263 6173 297
rect 6207 263 6242 297
rect 6276 263 6311 297
rect 6345 263 6380 297
rect 6414 263 6449 297
rect 6483 263 6518 297
rect 6552 263 6587 297
rect 6621 263 6656 297
rect 6690 263 6725 297
rect 6759 263 6817 297
rect 6851 263 6867 297
rect 7060 294 7094 328
rect 7128 294 7162 328
rect 7347 564 7463 567
rect 8048 564 8169 567
rect 7347 530 7385 564
rect 7419 530 7457 564
rect 8059 530 8097 564
rect 8131 530 8169 564
rect 7347 529 7463 530
rect 7381 501 7463 529
rect 8048 529 8169 530
rect 8048 501 8135 529
rect 7347 460 7381 495
rect 7347 391 7381 426
rect 7347 321 7381 357
rect 8135 476 8169 495
rect 8135 404 8169 426
rect 8135 321 8169 357
rect 843 155 877 193
rect 1479 155 1513 193
rect 1723 155 1757 193
rect 3131 155 3165 193
rect 4957 224 4991 258
rect 4923 141 5025 224
rect 7026 258 7196 294
rect 7309 263 7347 297
rect 8127 287 8135 297
rect 8127 263 8165 287
rect 7060 224 7094 258
rect 7128 224 7162 258
rect 7026 217 7196 224
rect -2178 43 -2140 77
rect -1239 25 -1165 86
rect -887 25 -813 86
rect 81 35 196 73
rect 293 25 367 91
rect 575 25 609 75
rect 4923 39 4947 141
rect 6137 107 6172 141
rect 6206 107 6241 141
rect 6275 107 6310 141
rect 6344 107 6379 141
rect 6413 107 6448 141
rect 6482 107 6517 141
rect 6551 107 6586 141
rect 6620 107 6655 141
rect 6689 107 6724 141
rect 6758 107 6793 141
rect 6827 107 6862 141
rect 6896 107 6931 141
rect 6965 107 7000 141
rect 7034 107 7069 111
rect 7103 107 7138 111
rect 7172 107 7200 111
rect 6137 73 7200 107
rect 6137 39 6172 73
rect 6206 39 6241 73
rect 6275 39 6310 73
rect 6344 39 6379 73
rect 6413 39 6448 73
rect 6482 39 6517 73
rect 6551 39 6586 73
rect 6620 39 6655 73
rect 6689 39 6724 73
rect 6758 39 6793 73
rect 6827 39 6862 73
rect 6896 39 6931 73
rect 6965 39 7000 73
rect 7034 39 7069 73
rect 7103 39 7138 73
rect 7172 39 7200 73
rect -4754 -171 -4716 -137
rect -4331 -171 -4012 -137
rect -4046 -453 -4012 -171
rect -4046 -525 -4012 -487
rect -4046 -572 -4012 -559
rect -5843 -1630 -5809 -1550
rect -4143 -1574 -4109 -1351
rect -4143 -1596 -4102 -1574
rect -4143 -1730 -4136 -1596
<< viali >>
rect -2035 1381 -2001 1415
rect -1963 1381 -1929 1415
rect 829 1381 863 1415
rect 901 1381 935 1415
rect 689 1307 723 1341
rect 761 1307 795 1341
rect 1005 1307 1039 1341
rect 1077 1307 1111 1341
rect -391 1207 -357 1241
rect -391 1135 -357 1169
rect -391 1063 -357 1097
rect -2009 881 -1975 915
rect -1937 881 -1903 915
rect -1517 868 -1483 902
rect -1445 868 -1411 902
rect -778 868 -744 902
rect -706 868 -672 902
rect -515 868 -481 902
rect -443 868 -409 902
rect -391 681 -357 715
rect -391 609 -357 643
rect -391 537 -357 571
rect -601 425 -567 459
rect -601 353 -567 387
rect -1694 274 -1660 308
rect -1622 274 -1588 308
rect -1500 256 -1466 290
rect -1500 184 -1466 218
rect -1219 256 -1185 290
rect -1219 184 -1185 218
rect -867 256 -833 290
rect -867 184 -833 218
rect 6130 1411 6134 1415
rect 6134 1411 6164 1415
rect 6202 1411 6236 1415
rect 6130 1381 6164 1411
rect 6202 1381 6236 1411
rect 5778 1307 5812 1341
rect 5850 1307 5884 1341
rect -39 1207 -5 1241
rect -39 1135 -5 1169
rect -39 1063 -5 1097
rect -215 425 -181 459
rect -215 353 -181 387
rect -39 681 -5 715
rect -39 609 -5 643
rect -39 537 -5 571
rect 313 681 347 715
rect 313 609 347 643
rect 313 537 347 571
rect 137 425 171 459
rect 137 353 171 387
rect 489 193 523 227
rect 489 121 523 155
rect 4610 1157 4644 1191
rect 4610 1085 4644 1119
rect 4942 1160 4976 1190
rect 5018 1160 5052 1190
rect 4942 1156 4957 1160
rect 4957 1156 4976 1160
rect 5018 1156 5025 1160
rect 5025 1156 5052 1160
rect 5094 1156 5128 1190
rect 5170 1156 5204 1190
rect 5246 1156 5280 1190
rect 5322 1156 5356 1190
rect 5398 1156 5432 1190
rect 5473 1169 5507 1190
rect 5473 1156 5487 1169
rect 5487 1156 5507 1169
rect 5548 1156 5582 1190
rect 4942 1091 4976 1118
rect 5018 1091 5052 1118
rect 4942 1084 4957 1091
rect 4957 1084 4976 1091
rect 5018 1084 5025 1091
rect 5025 1084 5052 1091
rect 5094 1084 5128 1118
rect 5170 1084 5204 1118
rect 5246 1084 5280 1118
rect 5322 1111 5323 1118
rect 5323 1111 5356 1118
rect 5398 1111 5427 1118
rect 5427 1111 5432 1118
rect 5322 1084 5356 1111
rect 5398 1084 5432 1111
rect 5473 1084 5507 1118
rect 5548 1084 5582 1118
rect 5683 1207 5717 1241
rect 5683 1135 5717 1169
rect 5683 1063 5717 1097
rect 6305 1207 6339 1241
rect 6305 1135 6339 1169
rect 6305 1063 6339 1097
rect 6440 1165 6474 1199
rect 6519 1165 6553 1199
rect 6597 1165 6631 1199
rect 6675 1165 6709 1199
rect 6753 1165 6787 1199
rect 6831 1165 6865 1199
rect 6909 1165 6943 1199
rect 6987 1165 7021 1199
rect 7065 1195 7094 1199
rect 7094 1195 7099 1199
rect 7143 1195 7162 1199
rect 7162 1195 7177 1199
rect 7065 1165 7099 1195
rect 7143 1165 7177 1195
rect 6440 1093 6474 1127
rect 6519 1111 6534 1127
rect 6534 1111 6553 1127
rect 6597 1111 6613 1127
rect 6613 1111 6631 1127
rect 6675 1111 6691 1127
rect 6691 1111 6709 1127
rect 6519 1093 6553 1111
rect 6597 1093 6631 1111
rect 6675 1093 6709 1111
rect 6753 1093 6787 1127
rect 6831 1093 6865 1127
rect 6909 1093 6943 1127
rect 6987 1093 7021 1127
rect 7065 1126 7094 1127
rect 7094 1126 7099 1127
rect 7143 1126 7162 1127
rect 7162 1126 7177 1127
rect 7065 1093 7099 1126
rect 7143 1093 7177 1126
rect 4940 1022 4974 1038
rect 5012 1022 5046 1038
rect 4610 983 4644 1017
rect 4682 983 4716 1017
rect 4940 1004 4957 1022
rect 4957 1004 4974 1022
rect 5012 1004 5025 1022
rect 5025 1004 5046 1022
rect 5084 1004 5118 1038
rect 5156 1004 5190 1038
rect 5239 983 5273 1017
rect 5311 983 5345 1017
rect 5495 983 5529 1017
rect 5567 983 5601 1017
rect 6421 983 6455 1017
rect 6493 983 6527 1017
rect 6677 983 6711 1017
rect 6749 983 6783 1017
rect 7022 988 7026 1011
rect 7026 988 7056 1011
rect 7094 988 7128 1011
rect 7166 988 7196 1011
rect 7196 988 7200 1011
rect 7022 977 7056 988
rect 7094 977 7128 988
rect 7166 977 7200 988
rect 6571 863 6605 897
rect 6643 863 6677 897
rect 7525 941 7559 975
rect 5171 524 5205 558
rect 5909 719 5943 753
rect 5981 719 6015 753
rect 5727 645 5749 679
rect 5749 645 5761 679
rect 5799 645 5817 679
rect 5817 645 5833 679
rect 5683 524 5717 558
rect 6013 645 6047 679
rect 6085 645 6119 679
rect 6193 645 6205 679
rect 6205 645 6227 679
rect 6265 645 6273 679
rect 6273 645 6299 679
rect 5171 452 5205 486
rect 5171 380 5205 414
rect 5683 452 5717 486
rect 5683 380 5717 414
rect 6305 524 6339 558
rect 7525 869 7559 903
rect 7347 604 7381 638
rect 8135 604 8169 638
rect 6305 452 6339 486
rect 6305 380 6339 414
rect 6817 524 6851 558
rect 6817 452 6851 486
rect 6817 380 6851 414
rect 7385 530 7419 564
rect 7457 530 7491 564
rect 8025 530 8059 564
rect 8097 530 8131 564
rect 8135 460 8169 476
rect 8135 442 8169 460
rect 8135 391 8169 404
rect 8135 370 8169 391
rect 843 193 877 227
rect 843 121 877 155
rect 1479 193 1513 227
rect 1479 121 1513 155
rect 1723 193 1757 227
rect 1723 121 1757 155
rect 3131 193 3165 227
rect 3131 121 3165 155
rect 7275 263 7309 297
rect 7347 287 7381 297
rect 7347 263 7381 287
rect 8093 263 8127 297
rect 8165 287 8169 297
rect 8169 287 8199 297
rect 8165 263 8199 287
rect 7022 141 7200 217
rect -2212 43 -2178 77
rect -2140 43 -2106 77
rect 7022 111 7034 141
rect 7034 111 7069 141
rect 7069 111 7103 141
rect 7103 111 7138 141
rect 7138 111 7172 141
rect 7172 111 7200 141
rect -4788 -171 -4754 -137
rect -4716 -171 -4682 -137
rect -4046 -487 -4012 -453
rect -4046 -559 -4012 -525
<< metal1 >>
rect 5473 1526 7088 1532
rect 5473 1486 5986 1526
rect 5524 1480 5986 1486
tri 5974 1468 5986 1480 ne
rect 6038 1474 6050 1526
rect 6102 1480 7088 1526
rect 7140 1480 7152 1532
rect 7204 1480 7210 1532
rect 5986 1468 6102 1474
tri 6102 1468 6114 1480 nw
rect -2047 1415 487 1421
tri 487 1415 493 1421 sw
rect 817 1415 6248 1421
rect -2047 1381 -2035 1415
rect -2001 1381 -1963 1415
rect -1929 1413 493 1415
tri 493 1413 495 1415 sw
rect -1929 1381 495 1413
tri 495 1381 527 1413 sw
rect 817 1381 829 1415
rect 863 1381 901 1415
rect 935 1381 6130 1415
rect 6164 1381 6202 1415
rect 6236 1381 6248 1415
rect -2047 1375 527 1381
tri 527 1375 533 1381 sw
rect 817 1375 6248 1381
tri 467 1347 495 1375 ne
rect 495 1347 533 1375
tri 533 1347 561 1375 sw
tri 495 1341 501 1347 ne
rect 501 1341 5896 1347
tri 501 1307 535 1341 ne
rect 535 1307 689 1341
rect 723 1307 761 1341
rect 795 1307 1005 1341
rect 1039 1307 1077 1341
rect 1111 1307 5778 1341
rect 5812 1307 5850 1341
rect 5884 1307 5896 1341
tri 535 1301 541 1307 ne
rect 541 1301 5896 1307
rect -1853 1051 -1781 1253
rect -498 1241 307 1253
rect -498 1207 -391 1241
rect -357 1207 -39 1241
rect -5 1207 307 1241
rect -498 1169 307 1207
rect -498 1135 -391 1169
rect -357 1135 -39 1169
rect -5 1135 307 1169
rect -498 1097 307 1135
rect -498 1063 -391 1097
rect -357 1063 -39 1097
rect -5 1063 307 1097
rect -498 1051 307 1063
rect 327 1051 344 1253
rect 682 1051 792 1253
rect 4656 1244 7977 1253
rect 4656 1241 7861 1244
rect 4656 1207 5683 1241
rect 5717 1207 6305 1241
rect 6339 1207 7861 1241
rect 4604 1191 4650 1203
rect 4604 1157 4610 1191
rect 4644 1157 4650 1191
rect 4604 1119 4650 1157
rect 4604 1085 4610 1119
rect 4644 1085 4650 1119
rect 4604 1073 4650 1085
rect 4656 1199 7861 1207
rect 4656 1190 6440 1199
rect 4656 1156 4942 1190
rect 4976 1156 5018 1190
rect 5052 1156 5094 1190
rect 5128 1156 5170 1190
rect 5204 1156 5246 1190
rect 5280 1156 5322 1190
rect 5356 1156 5398 1190
rect 5432 1156 5473 1190
rect 5507 1156 5548 1190
rect 5582 1169 6440 1190
rect 5582 1156 5683 1169
rect 4656 1135 5683 1156
rect 5717 1135 6305 1169
rect 6339 1165 6440 1169
rect 6474 1165 6519 1199
rect 6553 1165 6597 1199
rect 6631 1165 6675 1199
rect 6709 1165 6753 1199
rect 6787 1165 6831 1199
rect 6865 1165 6909 1199
rect 6943 1165 6987 1199
rect 7021 1165 7065 1199
rect 7099 1165 7143 1199
rect 7177 1165 7861 1199
rect 6339 1135 7861 1165
rect 4656 1127 7861 1135
rect 4656 1118 6440 1127
rect 4656 1084 4942 1118
rect 4976 1084 5018 1118
rect 5052 1084 5094 1118
rect 5128 1084 5170 1118
rect 5204 1084 5246 1118
rect 5280 1084 5322 1118
rect 5356 1084 5398 1118
rect 5432 1084 5473 1118
rect 5507 1084 5548 1118
rect 5582 1097 6440 1118
rect 5582 1084 5683 1097
rect 4656 1063 5683 1084
rect 5717 1063 6305 1097
rect 6339 1093 6440 1097
rect 6474 1093 6519 1127
rect 6553 1093 6597 1127
rect 6631 1093 6675 1127
rect 6709 1093 6753 1127
rect 6787 1093 6831 1127
rect 6865 1093 6909 1127
rect 6943 1093 6987 1127
rect 7021 1093 7065 1127
rect 7099 1093 7143 1127
rect 7177 1093 7861 1127
rect 6339 1064 7861 1093
rect 6339 1063 7977 1064
rect 4656 1051 7977 1063
rect -2291 1038 7210 1051
rect -2291 1023 4940 1038
rect -1853 977 -1787 1023
rect -498 977 301 1023
rect 682 977 792 1023
rect 4598 1017 4940 1023
rect 4598 983 4610 1017
rect 4644 983 4682 1017
rect 4716 1004 4940 1017
rect 4974 1004 5012 1038
rect 5046 1004 5084 1038
rect 5118 1004 5156 1038
rect 5190 1023 7210 1038
rect 5190 1017 7088 1023
rect 5190 1004 5239 1017
rect 4716 983 5239 1004
rect 5273 983 5311 1017
rect 5345 983 5495 1017
rect 5529 983 5567 1017
rect 5601 983 5986 1017
rect 4598 977 5986 983
tri 5961 975 5963 977 ne
rect 5963 975 5986 977
tri 5963 952 5986 975 ne
tri -1318 941 -1310 949 se
rect -1310 941 -1231 949
tri -1338 921 -1318 941 se
rect -1318 921 -1231 941
tri -2532 915 -2526 921 se
rect -2526 915 -1891 921
tri -2566 881 -2532 915 se
rect -2532 881 -2009 915
rect -1975 881 -1937 915
rect -1903 881 -1891 915
tri -1351 908 -1338 921 se
rect -1338 908 -1231 921
rect -1192 911 -1033 940
tri -2572 875 -2566 881 se
rect -2566 875 -1891 881
rect -1529 903 -1231 908
rect -1529 902 -1291 903
tri -1291 902 -1290 903 nw
rect -790 902 -397 908
rect 2933 903 3285 949
rect 4295 909 4329 943
tri -2579 868 -2572 875 se
rect -2572 868 -2513 875
tri -2513 868 -2506 875 nw
rect -1529 868 -1517 902
rect -1483 868 -1445 902
rect -1411 868 -1325 902
tri -1325 868 -1291 902 nw
rect -790 868 -778 902
rect -744 868 -706 902
rect -672 868 -515 902
rect -481 868 -443 902
rect -409 868 -397 902
rect 6102 983 6421 1017
rect 6455 983 6493 1017
rect 6527 983 6677 1017
rect 6711 983 6749 1017
rect 6783 1011 7088 1017
rect 6783 983 7022 1011
rect 6102 977 7022 983
rect 7056 977 7088 1011
rect 6102 975 6125 977
tri 6125 975 6127 977 nw
tri 7004 975 7006 977 ne
rect 7006 975 7088 977
rect 6102 965 6115 975
tri 6115 965 6125 975 nw
tri 7006 965 7016 975 ne
rect 7016 971 7088 975
rect 7140 971 7152 1023
rect 7204 971 7210 1023
rect 7016 965 7210 971
rect 7519 975 7565 987
tri 6102 952 6115 965 nw
rect 7519 941 7525 975
rect 7559 941 7565 975
tri 7494 903 7519 928 se
rect 7519 903 7565 941
rect 7883 925 7917 959
rect 5986 895 6102 901
rect 6559 897 7525 903
tri -2584 863 -2579 868 se
rect -2579 863 -2518 868
tri -2518 863 -2513 868 nw
rect -1529 863 -1330 868
tri -1330 863 -1325 868 nw
tri -2585 862 -2584 863 se
rect -2584 862 -2519 863
tri -2519 862 -2518 863 nw
rect -1529 862 -1331 863
tri -1331 862 -1330 863 nw
rect -790 862 -397 868
rect 6559 863 6571 897
rect 6605 863 6643 897
rect 6677 869 7525 897
rect 7559 869 7565 903
rect 6677 863 7565 869
tri -2590 857 -2585 862 se
rect -2585 857 -2524 862
tri -2524 857 -2519 862 nw
rect 6559 857 7565 863
tri -2592 855 -2590 857 se
rect -2590 855 -2526 857
tri -2526 855 -2524 857 nw
tri -2596 851 -2592 855 se
rect -2592 851 -2530 855
tri -2530 851 -2526 855 nw
tri -2619 425 -2596 448 se
rect -2596 428 -2550 851
tri -2550 831 -2530 851 nw
rect 7861 804 7977 810
rect -2291 715 4656 801
rect 7068 778 7210 800
rect -2291 681 -391 715
rect -357 681 -39 715
rect -5 681 313 715
rect 347 681 4656 715
rect 5897 753 6174 759
rect 5897 719 5909 753
rect 5943 719 5981 753
rect 6015 719 6174 753
rect 5897 713 6174 719
tri 6174 713 6220 759 sw
tri 6153 685 6181 713 ne
rect 6181 685 6220 713
tri 6220 685 6248 713 sw
rect -2291 643 4656 681
rect -2291 609 -391 643
rect -357 609 -39 643
rect -5 609 313 643
rect 347 609 4656 643
rect 5715 679 6131 685
rect 5715 645 5727 679
rect 5761 645 5799 679
rect 5833 645 6013 679
rect 6047 645 6085 679
rect 6119 645 6131 679
rect 5715 639 6131 645
rect 6181 679 6311 685
rect 6181 645 6193 679
rect 6227 645 6265 679
rect 6299 645 6311 679
rect 6181 639 6311 645
rect -2291 571 4656 609
rect 7068 598 7088 778
rect 7204 650 7210 778
tri 7443 682 7445 684 se
rect 7861 682 7977 688
tri 8071 682 8073 684 sw
tri 7436 675 7443 682 se
rect 7443 678 7445 682
rect 8071 678 8073 682
rect 7443 675 8073 678
tri 7210 650 7235 675 sw
tri 7411 650 7436 675 se
rect 7436 650 8073 675
tri 8073 650 8105 682 sw
rect 7204 638 8181 650
rect 7204 604 7347 638
rect 7381 604 8135 638
rect 8169 604 8181 638
rect 7204 598 8181 604
rect -2291 537 -391 571
rect -357 537 -39 571
rect -5 537 313 571
rect 347 537 4656 571
rect -2291 525 4656 537
rect 5127 564 8211 570
rect 5127 558 7385 564
rect 5127 524 5171 558
rect 5205 524 5683 558
rect 5717 524 6305 558
rect 6339 524 6817 558
rect 6851 530 7385 558
rect 7419 530 7457 564
rect 7491 530 7676 564
rect 6851 524 7676 530
rect 5127 512 7676 524
rect 7728 512 7752 564
rect 7804 530 8025 564
rect 8059 530 8097 564
rect 8131 530 8211 564
rect 7804 512 8211 530
rect 5127 489 8211 512
rect 5127 486 7676 489
rect -607 459 177 471
rect -2596 425 -2553 428
tri -2553 425 -2550 428 nw
tri -2630 414 -2619 425 se
rect -2619 414 -2564 425
tri -2564 414 -2553 425 nw
tri -2657 387 -2630 414 se
rect -2630 387 -2591 414
tri -2591 387 -2564 414 nw
rect -1714 406 -1595 456
rect -607 425 -601 459
rect -567 425 -215 459
rect -181 425 137 459
rect 171 425 177 459
rect -607 387 177 425
tri -2662 382 -2657 387 se
rect -2657 382 -2596 387
tri -2596 382 -2591 387 nw
tri -2676 368 -2662 382 se
rect -2662 368 -2616 382
rect -4746 316 -4740 368
rect -4688 316 -4676 368
rect -4624 362 -4618 368
tri -2682 362 -2676 368 se
rect -2676 362 -2616 368
tri -2616 362 -2596 382 nw
tri -2049 380 -2047 382 sw
rect -2049 367 -2047 380
tri -2100 362 -2095 367 ne
rect -2095 362 -2047 367
tri -2047 362 -2029 380 sw
rect -4624 353 -2625 362
tri -2625 353 -2616 362 nw
tri -2095 353 -2086 362 ne
rect -2086 353 -2029 362
tri -2029 353 -2020 362 sw
rect -607 353 -601 387
rect -567 353 -215 387
rect -181 353 137 387
rect 171 353 177 387
rect -4624 341 -2637 353
tri -2637 341 -2625 353 nw
tri -2086 341 -2074 353 ne
rect -2074 341 -2020 353
tri -2020 341 -2008 353 sw
rect -607 341 177 353
rect 5127 452 5171 486
rect 5205 452 5683 486
rect 5717 452 6305 486
rect 6339 452 6817 486
rect 6851 452 7676 486
rect 5127 437 7676 452
rect 7728 437 7752 489
rect 7804 476 8211 489
rect 7804 442 8135 476
rect 8169 442 8211 476
rect 7804 437 8211 442
rect 5127 414 8211 437
rect 5127 380 5171 414
rect 5205 380 5683 414
rect 5717 380 6305 414
rect 6339 380 6817 414
rect 6851 413 8211 414
rect 6851 380 7676 413
rect 5127 361 7676 380
rect 7728 361 7752 413
rect 7804 404 8211 413
rect 7804 370 8135 404
rect 8169 370 8211 404
rect 7804 361 8211 370
rect -4624 316 -2662 341
tri -2662 316 -2637 341 nw
tri -2074 316 -2049 341 ne
rect -2049 316 -2008 341
tri -2008 316 -1983 341 sw
tri -2049 314 -2047 316 ne
rect -2047 314 -1983 316
tri -1983 314 -1981 316 sw
tri -2047 308 -2041 314 ne
rect -2041 308 -1576 314
tri -2041 274 -2007 308 ne
rect -2007 274 -1694 308
rect -1660 274 -1622 308
rect -1588 274 -1576 308
rect 5127 309 8211 361
tri -2007 268 -2001 274 ne
rect -2001 268 -1576 274
rect -1506 290 -827 302
rect -1506 256 -1500 290
rect -1466 256 -1219 290
rect -1185 256 -867 290
rect -833 256 -827 290
rect 5127 297 7682 309
rect 5127 263 7275 297
rect 7309 263 7347 297
rect 7381 263 7682 297
rect 5127 257 7682 263
rect 7734 257 7746 309
rect 7798 297 8211 309
rect 7798 263 8093 297
rect 8127 263 8165 297
rect 8199 263 8211 297
rect 7798 257 8211 263
rect -1506 218 -827 256
rect -1506 184 -1500 218
rect -1466 184 -1219 218
rect -1185 184 -867 218
rect -833 184 -827 218
rect -1506 172 -827 184
rect 483 227 883 239
rect 483 193 489 227
rect 523 193 843 227
rect 877 193 883 227
rect 483 155 883 193
rect 483 121 489 155
rect 523 121 843 155
rect 877 121 883 155
rect 483 109 883 121
rect 1473 227 3171 239
rect 1473 193 1479 227
rect 1513 193 1723 227
rect 1757 193 3131 227
rect 3165 193 3171 227
rect 1473 155 3171 193
rect 1473 121 1479 155
rect 1513 121 1723 155
rect 1757 121 3131 155
rect 3165 121 3171 155
rect 1473 109 3171 121
rect 7016 217 7088 229
rect 7016 111 7022 217
rect 7204 113 7210 229
rect 7200 111 7210 113
rect 7016 99 7210 111
tri -4786 77 -4774 89 se
rect -4774 77 -2094 89
tri -4820 43 -4786 77 se
rect -4786 43 -2212 77
rect -2178 43 -2140 77
rect -2106 43 -2094 77
tri -4826 37 -4820 43 se
rect -4820 37 -2094 43
tri -4870 -7 -4826 37 se
rect -4826 -7 -4796 37
tri -4796 -7 -4752 37 nw
tri -4892 -29 -4870 -7 se
rect -4870 -27 -4816 -7
tri -4816 -27 -4796 -7 nw
rect -4870 -29 -4818 -27
tri -4818 -29 -4816 -27 nw
rect -4550 -29 -4524 -27
tri -4524 -29 -4522 -27 nw
tri -5454 -55 -5428 -29 se
rect -5428 -49 -4838 -29
tri -4838 -49 -4818 -29 nw
rect -4550 -49 -4544 -29
tri -4544 -49 -4524 -29 nw
rect -5428 -55 -4844 -49
tri -4844 -55 -4838 -49 nw
rect -4746 -55 -4694 -49
tri -4550 -55 -4544 -49 nw
rect -5454 -61 -4866 -55
rect -5402 -77 -4866 -61
tri -4866 -77 -4844 -55 nw
rect -5402 -81 -4870 -77
tri -4870 -81 -4866 -77 nw
tri -4750 -81 -4746 -77 se
rect -5454 -125 -5402 -113
tri -5402 -124 -5359 -81 nw
tri -4793 -124 -4750 -81 se
rect -4750 -107 -4746 -81
rect -4750 -119 -4694 -107
rect -4750 -124 -4746 -119
tri -4800 -131 -4793 -124 se
rect -4793 -131 -4746 -124
rect -4800 -137 -4746 -131
tri -4694 -131 -4670 -107 sw
rect -4694 -137 -4670 -131
rect -4800 -171 -4788 -137
rect -4754 -171 -4746 -137
rect -4682 -171 -4670 -137
rect -4800 -177 -4670 -171
rect -5454 -183 -5402 -177
rect -6060 -413 -6026 -211
rect -3992 -413 -3958 -211
rect -6060 -571 -6026 -441
rect -4052 -453 -4006 -441
rect -4052 -487 -4046 -453
rect -4012 -487 -4006 -453
rect -4052 -525 -4006 -487
rect -4052 -559 -4046 -525
rect -4012 -559 -4006 -525
rect -4052 -571 -4006 -559
tri -2850 -782 -2816 -748 ne
tri -2764 -782 -2730 -748 nw
rect -4110 -1208 -4041 -1173
rect -6668 -1562 -6394 -1319
rect -6180 -1332 -6060 -1280
rect -6060 -1562 -6026 -1360
rect -3992 -1562 -3958 -1360
tri -6050 -1635 -5977 -1562 ne
rect -5977 -1635 -4038 -1562
tri -4038 -1635 -3965 -1562 nw
tri -5977 -1636 -5976 -1635 ne
rect -5976 -1636 -4039 -1635
tri -4039 -1636 -4038 -1635 nw
tri -4220 -1708 -4148 -1636 ne
tri -4090 -1687 -4039 -1636 nw
rect -6060 -2207 -6026 -2005
rect -4177 -2207 -4143 -2005
rect -6099 -2235 -3929 -2207
<< via1 >>
rect 5986 1474 6038 1526
rect 6050 1474 6102 1526
rect 7088 1480 7140 1532
rect 7152 1480 7204 1532
rect 7861 1064 7977 1244
rect 5986 901 6102 1017
rect 7088 1011 7140 1023
rect 7088 977 7094 1011
rect 7094 977 7128 1011
rect 7128 977 7140 1011
rect 7088 971 7140 977
rect 7152 1011 7204 1023
rect 7152 977 7166 1011
rect 7166 977 7200 1011
rect 7200 977 7204 1011
rect 7152 971 7204 977
rect 7088 598 7204 778
rect 7861 688 7977 804
rect 7676 512 7728 564
rect 7752 512 7804 564
rect -4740 316 -4688 368
rect -4676 316 -4624 368
rect 7676 437 7728 489
rect 7752 437 7804 489
rect 7676 361 7728 413
rect 7752 361 7804 413
rect 7682 257 7734 309
rect 7746 257 7798 309
rect 7088 217 7204 229
rect 7088 113 7200 217
rect 7200 113 7204 217
rect -5454 -113 -5402 -61
rect -4746 -107 -4694 -55
rect -5454 -177 -5402 -125
rect -4746 -137 -4694 -119
rect -4746 -171 -4716 -137
rect -4716 -171 -4694 -137
<< metal2 >>
rect 5986 1526 6102 1532
rect 6038 1474 6050 1526
rect 5986 1017 6102 1474
rect 5986 895 6102 901
rect 7082 1480 7088 1532
rect 7140 1480 7152 1532
rect 7204 1480 7210 1532
rect 7082 1023 7210 1480
rect 7082 971 7088 1023
rect 7140 971 7152 1023
rect 7204 971 7210 1023
rect 7082 778 7210 971
rect 7082 598 7088 778
rect 7204 598 7210 778
rect 7861 1244 7977 1250
rect 7861 804 7977 1064
rect 7861 682 7977 688
rect -4746 316 -4740 368
rect -4688 316 -4676 368
rect -4624 316 -4618 368
rect -4746 309 -4634 316
tri -4634 309 -4627 316 nw
rect -4746 257 -4686 309
tri -4686 257 -4634 309 nw
rect -4746 -55 -4694 257
tri -4694 249 -4686 257 nw
rect 7082 229 7210 598
rect 7676 564 7804 570
rect 7728 512 7752 564
rect 7676 489 7804 512
rect 7728 437 7752 489
rect 7676 413 7804 437
rect 7728 361 7752 413
rect 7676 309 7804 361
rect 7676 257 7682 309
rect 7734 257 7746 309
rect 7798 257 7804 309
rect 7082 113 7088 229
rect 7204 113 7210 229
rect -5454 -61 -5402 -55
rect -5454 -125 -5402 -113
rect -4746 -119 -4694 -107
rect -4746 -177 -4694 -171
tri -5482 -792 -5454 -764 se
rect -5454 -836 -5402 -177
use hvnTran_CDNS_52468879185633  hvnTran_CDNS_52468879185633_0
timestamp 1707688321
transform 1 0 -346 0 1 1075
box -79 -26 375 226
use hvpTran_CDNS_52468879185530  hvpTran_CDNS_52468879185530_0
timestamp 1707688321
transform -1 0 302 0 -1 723
box -119 -66 767 666
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 -567 -1 0 459
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 8169 -1 0 476
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 -181 -1 0 459
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 -1 171 -1 0 459
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 -1 4644 -1 0 1191
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 0 1 843 -1 0 227
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 1 489 -1 0 227
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 0 1 7525 -1 0 975
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 4716 0 1 983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 6119 0 1 645
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 7381 0 1 263
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 8199 0 1 263
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 7491 0 1 530
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 8131 0 1 530
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform -1 0 5345 0 1 983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform -1 0 5601 0 1 983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform -1 0 795 0 -1 1341
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform -1 0 1111 0 -1 1341
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform -1 0 935 0 -1 1415
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform -1 0 6015 0 -1 753
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform -1 0 6236 0 -1 1415
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform -1 0 5884 0 -1 1341
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform -1 0 6677 0 -1 897
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 0 1 -1500 1 0 184
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 0 1 -1219 1 0 184
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 0 1 -867 1 0 184
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 0 -1 1757 1 0 121
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 0 -1 1513 1 0 121
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 0 -1 3165 1 0 121
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1707688321
transform 1 0 -515 0 -1 902
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1707688321
transform 1 0 -1694 0 -1 308
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1707688321
transform 1 0 -1517 0 -1 902
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1707688321
transform 1 0 -778 0 -1 902
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1707688321
transform 1 0 5727 0 1 645
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1707688321
transform 1 0 6193 0 1 645
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1707688321
transform 1 0 6677 0 1 983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1707688321
transform 1 0 6421 0 1 983
box 0 0 1 1
use L1M1_CDNS_5246887918558  L1M1_CDNS_5246887918558_0
timestamp 1707688321
transform 0 1 7022 -1 0 217
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 -357 -1 0 715
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 -5 -1 0 715
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 347 -1 0 715
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 1 5171 1 0 380
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 1 6817 1 0 380
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 5717 1 0 1063
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 6339 1 0 380
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 6339 1 0 1063
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1707688321
transform 0 -1 5717 1 0 380
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1707688321
transform 0 -1 -5 1 0 1063
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1707688321
transform 0 -1 -357 1 0 1063
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform 0 1 7022 -1 0 1011
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1707688321
transform 1 0 4923 0 1 1492
box -12 -6 550 40
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_0
timestamp 1707688321
transform -1 0 6870 0 1 263
box -12 -6 1414 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1707688321
transform 1 0 6586 0 1 1492
box -12 -6 622 40
use L1M1_CDNS_52468879185333  L1M1_CDNS_52468879185333_0
timestamp 1707688321
transform 0 1 7022 1 0 610
box -12 -6 190 184
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform 1 0 8135 0 1 604
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 1 0 7347 0 1 604
box 0 0 1 1
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1707688321
transform -1 0 6506 0 1 1492
box -12 -6 982 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 7210 0 1 971
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 7210 0 1 1480
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 1 0 7676 0 1 257
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 1 7861 -1 0 1250
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 7861 -1 0 810
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform 0 1 5986 1 0 895
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 1 0 7082 0 1 113
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform -1 0 7210 0 1 598
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 5986 1 0 1468
box 0 0 1 1
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_0
timestamp 1707688321
transform -1 0 6806 0 -1 971
box -79 -26 279 226
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_1
timestamp 1707688321
transform 1 0 5216 0 -1 971
box -79 -26 279 226
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_0
timestamp 1707688321
transform -1 0 6294 0 1 763
box -79 -26 279 626
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_1
timestamp 1707688321
transform 1 0 5728 0 1 763
box -79 -26 279 626
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_0
timestamp 1707688321
transform -1 0 6294 0 1 351
box -89 -36 289 236
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_1
timestamp 1707688321
transform 1 0 5728 0 1 351
box -89 -36 289 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_0
timestamp 1707688321
transform 1 0 6350 0 1 351
box -89 -36 545 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_1
timestamp 1707688321
transform 1 0 5216 0 1 351
box -89 -36 545 236
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 -1 -73 -1 0 955
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 0 -1 -249 -1 0 955
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 6252 1 0 1395
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 -1 5900 1 0 1396
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1707688321
transform 0 -1 6527 -1 0 695
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1707688321
transform 0 -1 5901 -1 0 695
box 0 0 1 1
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_0
timestamp 1707688321
transform 1 0 -352 0 -1 1373
box 0 0 1 1
use PYL1_CDNS_524688791851190  PYL1_CDNS_524688791851190_0
timestamp 1707688321
transform 1 0 -369 0 -1 91
box 0 0 678 66
use sky130_fd_io__com_ctl_ls_1  sky130_fd_io__com_ctl_ls_1_0
timestamp 1707688321
transform 1 0 -6060 0 -1 -121
box -91 0 2150 2319
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_0
timestamp 1707688321
transform -1 0 792 0 -1 1394
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_endcap  sky130_fd_io__sio_hvsbt_endcap_0
timestamp 1707688321
transform -1 0 4627 0 -1 1394
box -84 93 164 1337
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1707688321
transform -1 0 968 0 -1 1394
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1707688321
transform 1 0 -674 0 -1 1394
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x4  sky130_fd_io__sio_hvsbt_inv_x4_0
timestamp 1707688321
transform -1 0 -674 0 -1 1394
box -107 21 811 1369
use sky130_fd_io__sio_hvsbt_inv_x4  sky130_fd_io__sio_hvsbt_inv_x4_1
timestamp 1707688321
transform 1 0 968 0 -1 1394
box -107 21 811 1369
use sky130_fd_io__sio_hvsbt_inv_x8  sky130_fd_io__sio_hvsbt_inv_x8_0
timestamp 1707688321
transform 1 0 3080 0 -1 1394
box -108 21 1517 1369
use sky130_fd_io__sio_hvsbt_inv_x8  sky130_fd_io__sio_hvsbt_inv_x8_1
timestamp 1707688321
transform 1 0 1672 0 -1 1394
box -108 21 1517 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_0
timestamp 1707688321
transform 1 0 330 0 -1 1394
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1707688321
transform -1 0 -1882 0 -1 1394
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_1
timestamp 1707688321
transform -1 0 -1378 0 -1 1394
box -107 21 487 1369
use sky130_fd_io__sio_lvlp_inv_x4  sky130_fd_io__sio_lvlp_inv_x4_0
timestamp 1707688321
transform 1 0 7474 0 -1 1024
box -77 21 645 859
<< labels >>
flabel comment s 1121 1409 1121 1409 0 FreeSans 200 180 0 0 hld_i_h_ls
flabel comment s 5845 1451 5845 1451 0 FreeSans 200 180 0 0 in_c
flabel comment s 6171 1451 6171 1451 0 FreeSans 200 180 0 0 in_t
flabel comment s 6542 737 6542 737 0 FreeSans 200 180 0 0 out_c
flabel comment s 5469 731 5469 731 0 FreeSans 200 180 0 0 out_t
flabel comment s 3413 930 3413 930 0 FreeSans 200 180 0 0 hld_i_h_n
flabel comment s 3406 12 3406 12 0 FreeSans 200 180 0 0 hld_i_h
flabel comment s 1813 12 1813 12 0 FreeSans 200 180 0 0 hld_i_h
flabel comment s 1625 186 1625 186 0 FreeSans 200 180 0 0 hld_i_h
flabel comment s 764 214 764 214 0 FreeSans 200 180 0 0 hld_i_h_ls
flabel comment s 1119 16 1119 16 0 FreeSans 200 180 0 0 hld_i_h_n_ls
flabel comment s 4718 64 4718 64 0 FreeSans 200 180 0 0 hld_i_h_ls
flabel comment s 4849 1337 4849 1337 0 FreeSans 200 180 0 0 hld_i_h_n_ls
flabel comment s 1119 1364 1119 1364 0 FreeSans 200 180 0 0 hld_i_h_n_ls
flabel comment s 888 16 888 16 0 FreeSans 200 180 0 0 hld_i_h_ls
flabel comment s 406 14 406 14 0 FreeSans 200 180 0 0 od_h_n
flabel comment s 591 16 591 16 0 FreeSans 200 180 0 0 hld_h_n
flabel metal1 s -6060 -413 -6026 -211 3 FreeSans 400 0 0 0 vcc_io
port 1 nsew
flabel metal1 s -4110 -1208 -4041 -1173 3 FreeSans 520 0 0 0 hld_ovr
port 4 nsew
flabel metal1 s -4177 -2207 -4143 -2005 3 FreeSans 400 180 0 0 vpwr
port 2 nsew
flabel metal1 s -6043 -312 -6043 -312 3 FreeSans 400 0 0 0 vcc_io
flabel metal1 s -3992 -1562 -3958 -1360 7 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s -6060 -571 -6026 -441 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s -3992 -413 -3958 -211 7 FreeSans 400 0 0 0 vcc_io
port 1 nsew
flabel metal1 s -3975 -312 -3975 -312 7 FreeSans 400 0 0 0 vcc_io
flabel metal1 s -1714 406 -1595 456 3 FreeSans 520 0 0 0 hld_i_ovr_h
port 5 nsew
flabel metal1 s -4160 -2106 -4160 -2106 3 FreeSans 400 180 0 0 vpwr
flabel metal1 s -6060 -2207 -6026 -2005 3 FreeSans 400 0 0 0 vpwr
port 2 nsew
flabel metal1 s -6060 -1562 -6026 -1360 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel metal1 s -6043 -2106 -6043 -2106 3 FreeSans 400 0 0 0 vpwr
flabel metal1 s -6043 -1461 -6043 -1461 3 FreeSans 400 0 0 0 vgnd
flabel metal1 s -3975 -1461 -3975 -1461 7 FreeSans 400 0 0 0 vgnd
flabel metal1 s -17 1051 6 1253 7 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s -374 1051 -351 1253 3 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s -1192 911 -1033 940 3 FreeSans 520 0 0 0 od_i_h
port 6 nsew
flabel metal1 s -6043 -506 -6043 -506 3 FreeSans 400 0 0 0 vgnd
flabel metal1 s 7101 882 7101 882 0 FreeSans 400 0 0 0 hld_i_vpwr_n
flabel metal1 s 4961 1320 4961 1320 0 FreeSans 400 0 0 0 hld_i_h_n_ls
flabel metal1 s 4663 1407 4663 1407 0 FreeSans 400 0 0 0 hld_i_h_ls
flabel metal1 s 1498 212 1498 212 0 FreeSans 400 0 0 0 hld_i_h
flabel metal1 s 154 525 171 801 3 FreeSans 400 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 8042 355 8071 489 3 FreeSans 400 180 0 0 vpwr
port 2 nsew
flabel metal1 s 7883 925 7917 959 0 FreeSans 400 0 0 0 hld_i_vpwr
port 7 nsew
flabel metal1 s 4295 909 4329 943 0 FreeSans 400 0 0 0 hld_i_h_n
port 8 nsew
flabel metal1 s 327 1051 344 1253 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel locali s 81 35 196 73 3 FreeSans 520 0 0 0 enable_h
port 10 nsew
flabel locali s 575 25 609 75 0 FreeSans 400 0 0 0 hld_h_n
port 11 nsew
<< properties >>
string GDS_END 85409484
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85363086
string path -135.700 -1.375 -135.700 -4.575 
<< end >>
