magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 60 614 4074 1730
<< pwell >>
rect 101 72 189 554
rect 2000 466 2134 554
rect 3945 72 4033 554
rect 101 -14 4033 72
<< mvpsubdiff >>
rect 127 494 163 528
rect 127 460 128 494
rect 162 460 163 494
rect 127 426 163 460
rect 127 392 128 426
rect 162 392 163 426
rect 127 358 163 392
rect 127 324 128 358
rect 162 324 163 358
rect 127 290 163 324
rect 127 256 128 290
rect 162 256 163 290
rect 127 222 163 256
rect 127 188 128 222
rect 162 188 163 222
rect 127 154 163 188
rect 127 120 128 154
rect 162 120 163 154
rect 2026 526 2108 528
rect 2026 492 2050 526
rect 2084 492 2108 526
rect 3971 487 4007 528
rect 3971 453 3972 487
rect 4006 453 4007 487
rect 3971 419 4007 453
rect 3971 385 3972 419
rect 4006 385 4007 419
rect 3971 351 4007 385
rect 3971 317 3972 351
rect 4006 317 4007 351
rect 3971 283 4007 317
rect 3971 249 3972 283
rect 4006 249 4007 283
rect 3971 215 4007 249
rect 3971 181 3972 215
rect 4006 181 4007 215
rect 3971 147 4007 181
rect 127 46 163 120
rect 3971 113 3972 147
rect 4006 113 4007 147
rect 3971 79 4007 113
rect 3971 46 3972 79
rect 127 12 161 46
rect 195 12 229 46
rect 263 12 297 46
rect 331 12 365 46
rect 399 12 433 46
rect 467 12 501 46
rect 535 12 569 46
rect 603 12 637 46
rect 671 12 705 46
rect 739 12 773 46
rect 807 12 841 46
rect 875 12 909 46
rect 943 12 977 46
rect 1011 12 1045 46
rect 1079 12 1113 46
rect 1147 12 1181 46
rect 1215 12 1249 46
rect 1283 12 1317 46
rect 1351 12 1385 46
rect 1419 12 1453 46
rect 1487 12 1521 46
rect 1555 12 1589 46
rect 1623 12 1657 46
rect 1691 12 1725 46
rect 1759 12 1793 46
rect 1827 12 1861 46
rect 1895 12 1929 46
rect 1963 12 1997 46
rect 2031 12 2065 46
rect 2099 12 2133 46
rect 2167 12 2201 46
rect 2235 12 2269 46
rect 2303 12 2337 46
rect 2371 12 2405 46
rect 2439 12 2473 46
rect 2507 12 2541 46
rect 2575 12 2609 46
rect 2643 12 2677 46
rect 2711 12 2745 46
rect 2779 12 2813 46
rect 2847 12 2881 46
rect 2915 12 2949 46
rect 2983 12 3017 46
rect 3051 12 3085 46
rect 3119 12 3153 46
rect 3187 12 3221 46
rect 3255 12 3289 46
rect 3323 12 3357 46
rect 3391 12 3425 46
rect 3459 12 3493 46
rect 3527 12 3561 46
rect 3595 12 3629 46
rect 3663 12 3697 46
rect 3731 12 3765 46
rect 3799 12 3833 46
rect 3867 12 3901 46
rect 3935 45 3972 46
rect 4006 45 4007 79
rect 3935 12 4007 45
<< mvnsubdiff >>
rect 127 1662 4007 1663
rect 127 1628 161 1662
rect 195 1628 229 1662
rect 263 1628 297 1662
rect 331 1628 365 1662
rect 399 1628 433 1662
rect 467 1628 501 1662
rect 535 1628 569 1662
rect 603 1628 637 1662
rect 671 1628 705 1662
rect 739 1628 773 1662
rect 807 1628 841 1662
rect 875 1628 909 1662
rect 943 1628 977 1662
rect 1011 1628 1045 1662
rect 1079 1628 1113 1662
rect 1147 1628 1181 1662
rect 1215 1628 1249 1662
rect 1283 1628 1317 1662
rect 1351 1628 1385 1662
rect 1419 1628 1453 1662
rect 1487 1628 1521 1662
rect 1555 1628 1589 1662
rect 1623 1628 1657 1662
rect 1691 1628 1725 1662
rect 1759 1628 1793 1662
rect 1827 1628 1861 1662
rect 1895 1628 1929 1662
rect 1963 1628 1997 1662
rect 2031 1628 2065 1662
rect 2099 1628 2133 1662
rect 2167 1628 2201 1662
rect 2235 1628 2269 1662
rect 2303 1628 2337 1662
rect 2371 1628 2405 1662
rect 2439 1628 2473 1662
rect 2507 1628 2541 1662
rect 2575 1628 2609 1662
rect 2643 1628 2677 1662
rect 2711 1628 2745 1662
rect 2779 1628 2813 1662
rect 2847 1628 2881 1662
rect 2915 1628 2949 1662
rect 2983 1628 3017 1662
rect 3051 1628 3085 1662
rect 3119 1628 3153 1662
rect 3187 1628 3221 1662
rect 3255 1628 3289 1662
rect 3323 1628 3357 1662
rect 3391 1628 3425 1662
rect 3459 1628 3493 1662
rect 3527 1628 3561 1662
rect 3595 1628 3629 1662
rect 3663 1628 3697 1662
rect 3731 1628 3765 1662
rect 3799 1628 3833 1662
rect 3867 1628 3901 1662
rect 3935 1629 4007 1662
rect 3935 1628 3972 1629
rect 127 1627 3972 1628
rect 127 1564 163 1627
rect 127 1530 128 1564
rect 162 1530 163 1564
rect 127 1496 163 1530
rect 127 1462 128 1496
rect 162 1462 163 1496
rect 3971 1595 3972 1627
rect 4006 1595 4007 1629
rect 3971 1561 4007 1595
rect 3971 1527 3972 1561
rect 4006 1527 4007 1561
rect 3971 1493 4007 1527
rect 127 1428 163 1462
rect 127 1394 128 1428
rect 162 1394 163 1428
rect 3971 1459 3972 1493
rect 4006 1459 4007 1493
rect 3971 1425 4007 1459
rect 127 1360 163 1394
rect 127 1326 128 1360
rect 162 1326 163 1360
rect 127 1292 163 1326
rect 127 1258 128 1292
rect 162 1258 163 1292
rect 127 1224 163 1258
rect 127 1190 128 1224
rect 162 1190 163 1224
rect 127 1156 163 1190
rect 127 1122 128 1156
rect 162 1122 163 1156
rect 127 1088 163 1122
rect 127 1054 128 1088
rect 162 1054 163 1088
rect 127 1020 163 1054
rect 127 986 128 1020
rect 162 986 163 1020
rect 127 952 163 986
rect 127 918 128 952
rect 162 918 163 952
rect 127 884 163 918
rect 127 850 128 884
rect 162 850 163 884
rect 127 816 163 850
rect 127 782 128 816
rect 162 782 163 816
rect 127 748 163 782
rect 127 714 128 748
rect 162 714 163 748
rect 3971 1391 3972 1425
rect 4006 1391 4007 1425
rect 3971 1357 4007 1391
rect 3971 1323 3972 1357
rect 4006 1323 4007 1357
rect 3971 1289 4007 1323
rect 3971 1255 3972 1289
rect 4006 1255 4007 1289
rect 3971 1221 4007 1255
rect 3971 1187 3972 1221
rect 4006 1187 4007 1221
rect 3971 1153 4007 1187
rect 3971 1119 3972 1153
rect 4006 1119 4007 1153
rect 3971 1085 4007 1119
rect 3971 1051 3972 1085
rect 4006 1051 4007 1085
rect 3971 1017 4007 1051
rect 3971 983 3972 1017
rect 4006 983 4007 1017
rect 3971 949 4007 983
rect 3971 915 3972 949
rect 4006 915 4007 949
rect 3971 881 4007 915
rect 3971 847 3972 881
rect 4006 847 4007 881
rect 3971 813 4007 847
rect 3971 779 3972 813
rect 4006 779 4007 813
rect 127 680 163 714
rect 3971 680 4007 779
<< mvpsubdiffcont >>
rect 128 460 162 494
rect 128 392 162 426
rect 128 324 162 358
rect 128 256 162 290
rect 128 188 162 222
rect 128 120 162 154
rect 2050 492 2084 526
rect 3972 453 4006 487
rect 3972 385 4006 419
rect 3972 317 4006 351
rect 3972 249 4006 283
rect 3972 181 4006 215
rect 3972 113 4006 147
rect 161 12 195 46
rect 229 12 263 46
rect 297 12 331 46
rect 365 12 399 46
rect 433 12 467 46
rect 501 12 535 46
rect 569 12 603 46
rect 637 12 671 46
rect 705 12 739 46
rect 773 12 807 46
rect 841 12 875 46
rect 909 12 943 46
rect 977 12 1011 46
rect 1045 12 1079 46
rect 1113 12 1147 46
rect 1181 12 1215 46
rect 1249 12 1283 46
rect 1317 12 1351 46
rect 1385 12 1419 46
rect 1453 12 1487 46
rect 1521 12 1555 46
rect 1589 12 1623 46
rect 1657 12 1691 46
rect 1725 12 1759 46
rect 1793 12 1827 46
rect 1861 12 1895 46
rect 1929 12 1963 46
rect 1997 12 2031 46
rect 2065 12 2099 46
rect 2133 12 2167 46
rect 2201 12 2235 46
rect 2269 12 2303 46
rect 2337 12 2371 46
rect 2405 12 2439 46
rect 2473 12 2507 46
rect 2541 12 2575 46
rect 2609 12 2643 46
rect 2677 12 2711 46
rect 2745 12 2779 46
rect 2813 12 2847 46
rect 2881 12 2915 46
rect 2949 12 2983 46
rect 3017 12 3051 46
rect 3085 12 3119 46
rect 3153 12 3187 46
rect 3221 12 3255 46
rect 3289 12 3323 46
rect 3357 12 3391 46
rect 3425 12 3459 46
rect 3493 12 3527 46
rect 3561 12 3595 46
rect 3629 12 3663 46
rect 3697 12 3731 46
rect 3765 12 3799 46
rect 3833 12 3867 46
rect 3901 12 3935 46
rect 3972 45 4006 79
<< mvnsubdiffcont >>
rect 161 1628 195 1662
rect 229 1628 263 1662
rect 297 1628 331 1662
rect 365 1628 399 1662
rect 433 1628 467 1662
rect 501 1628 535 1662
rect 569 1628 603 1662
rect 637 1628 671 1662
rect 705 1628 739 1662
rect 773 1628 807 1662
rect 841 1628 875 1662
rect 909 1628 943 1662
rect 977 1628 1011 1662
rect 1045 1628 1079 1662
rect 1113 1628 1147 1662
rect 1181 1628 1215 1662
rect 1249 1628 1283 1662
rect 1317 1628 1351 1662
rect 1385 1628 1419 1662
rect 1453 1628 1487 1662
rect 1521 1628 1555 1662
rect 1589 1628 1623 1662
rect 1657 1628 1691 1662
rect 1725 1628 1759 1662
rect 1793 1628 1827 1662
rect 1861 1628 1895 1662
rect 1929 1628 1963 1662
rect 1997 1628 2031 1662
rect 2065 1628 2099 1662
rect 2133 1628 2167 1662
rect 2201 1628 2235 1662
rect 2269 1628 2303 1662
rect 2337 1628 2371 1662
rect 2405 1628 2439 1662
rect 2473 1628 2507 1662
rect 2541 1628 2575 1662
rect 2609 1628 2643 1662
rect 2677 1628 2711 1662
rect 2745 1628 2779 1662
rect 2813 1628 2847 1662
rect 2881 1628 2915 1662
rect 2949 1628 2983 1662
rect 3017 1628 3051 1662
rect 3085 1628 3119 1662
rect 3153 1628 3187 1662
rect 3221 1628 3255 1662
rect 3289 1628 3323 1662
rect 3357 1628 3391 1662
rect 3425 1628 3459 1662
rect 3493 1628 3527 1662
rect 3561 1628 3595 1662
rect 3629 1628 3663 1662
rect 3697 1628 3731 1662
rect 3765 1628 3799 1662
rect 3833 1628 3867 1662
rect 3901 1628 3935 1662
rect 128 1530 162 1564
rect 128 1462 162 1496
rect 3972 1595 4006 1629
rect 3972 1527 4006 1561
rect 128 1394 162 1428
rect 3972 1459 4006 1493
rect 128 1326 162 1360
rect 128 1258 162 1292
rect 128 1190 162 1224
rect 128 1122 162 1156
rect 128 1054 162 1088
rect 128 986 162 1020
rect 128 918 162 952
rect 128 850 162 884
rect 128 782 162 816
rect 128 714 162 748
rect 3972 1391 4006 1425
rect 3972 1323 4006 1357
rect 3972 1255 4006 1289
rect 3972 1187 4006 1221
rect 3972 1119 4006 1153
rect 3972 1051 4006 1085
rect 3972 983 4006 1017
rect 3972 915 4006 949
rect 3972 847 4006 881
rect 3972 779 4006 813
<< poly >>
rect 602 1452 878 1468
rect 602 1418 760 1452
rect 794 1418 828 1452
rect 862 1418 878 1452
rect 602 1402 878 1418
rect 1347 1452 1516 1468
rect 1347 1418 1365 1452
rect 1399 1418 1433 1452
rect 1467 1418 1516 1452
rect 1347 1402 1516 1418
rect 602 1396 702 1402
rect 758 1396 878 1402
rect 1396 1396 1516 1402
rect 2618 1452 2787 1468
rect 2618 1418 2667 1452
rect 2701 1418 2735 1452
rect 2769 1418 2787 1452
rect 2618 1402 2787 1418
rect 3207 1452 3343 1468
rect 3207 1418 3225 1452
rect 3259 1418 3293 1452
rect 3327 1418 3343 1452
rect 3207 1402 3343 1418
rect 2618 1396 2738 1402
rect 290 732 390 744
rect 446 732 546 744
rect 245 716 546 732
rect 245 682 261 716
rect 295 682 546 716
rect 245 672 546 682
rect 245 648 311 672
rect 245 614 261 648
rect 295 614 311 648
rect 245 598 311 614
rect 290 186 470 192
rect 526 186 706 192
rect 1420 186 1500 744
rect 1572 732 1672 744
rect 1728 732 1828 744
rect 1884 732 1984 744
rect 2150 732 2250 744
rect 2306 732 2406 744
rect 2462 732 2562 744
rect 1572 716 2017 732
rect 1572 682 1967 716
rect 2001 682 2017 716
rect 1572 672 2017 682
rect 1951 648 2017 672
rect 1951 614 1967 648
rect 2001 614 2017 648
rect 1951 598 2017 614
rect 2117 716 2562 732
rect 2117 682 2133 716
rect 2167 682 2562 716
rect 2117 672 2562 682
rect 2117 648 2183 672
rect 2117 614 2133 648
rect 2167 614 2183 648
rect 2117 598 2183 614
rect 1568 186 1748 192
rect 1804 186 1984 192
rect 290 170 927 186
rect 290 136 807 170
rect 841 136 875 170
rect 909 136 927 170
rect 290 120 927 136
rect 1347 120 1430 186
rect 1972 120 1984 186
rect 2150 186 2330 192
rect 2386 186 2566 192
rect 2634 186 2714 744
rect 3432 732 3532 744
rect 3588 732 3688 744
rect 3744 732 3844 744
rect 3432 716 3877 732
rect 3432 682 3827 716
rect 3861 682 3877 716
rect 3432 672 3877 682
rect 3811 648 3877 672
rect 3811 614 3827 648
rect 3861 614 3877 648
rect 3811 598 3877 614
rect 3428 186 3608 192
rect 3664 186 3844 192
rect 2150 120 2162 186
rect 2704 120 2787 186
rect 3207 120 3290 186
rect 3832 120 3844 186
<< polycont >>
rect 760 1418 794 1452
rect 828 1418 862 1452
rect 1365 1418 1399 1452
rect 1433 1418 1467 1452
rect 2667 1418 2701 1452
rect 2735 1418 2769 1452
rect 3225 1418 3259 1452
rect 3293 1418 3327 1452
rect 261 682 295 716
rect 261 614 295 648
rect 1967 682 2001 716
rect 1967 614 2001 648
rect 2133 682 2167 716
rect 2133 614 2167 648
rect 807 136 841 170
rect 875 136 909 170
rect 3827 682 3861 716
rect 3827 614 3861 648
<< locali >>
rect 127 1662 4007 1663
rect 127 1628 161 1662
rect 195 1628 229 1662
rect 263 1628 297 1662
rect 331 1628 365 1662
rect 399 1628 433 1662
rect 467 1628 501 1662
rect 535 1628 569 1662
rect 603 1628 637 1662
rect 671 1628 705 1662
rect 739 1628 773 1662
rect 807 1628 841 1662
rect 875 1628 909 1662
rect 943 1628 977 1662
rect 1011 1628 1045 1662
rect 1079 1628 1113 1662
rect 1147 1628 1181 1662
rect 1215 1628 1249 1662
rect 1283 1628 1317 1662
rect 1351 1628 1385 1662
rect 1419 1628 1453 1662
rect 1487 1628 1521 1662
rect 1555 1628 1589 1662
rect 1623 1628 1657 1662
rect 1691 1628 1725 1662
rect 1759 1628 1793 1662
rect 1827 1628 1861 1662
rect 1895 1628 1929 1662
rect 1963 1628 1997 1662
rect 2031 1628 2065 1662
rect 2099 1628 2133 1662
rect 2167 1628 2201 1662
rect 2235 1628 2269 1662
rect 2303 1628 2337 1662
rect 2371 1628 2405 1662
rect 2439 1628 2473 1662
rect 2507 1628 2541 1662
rect 2575 1628 2609 1662
rect 2643 1628 2677 1662
rect 2711 1628 2745 1662
rect 2779 1628 2813 1662
rect 2847 1628 2881 1662
rect 2915 1628 2949 1662
rect 2983 1628 3017 1662
rect 3051 1628 3085 1662
rect 3119 1628 3153 1662
rect 3187 1628 3221 1662
rect 3255 1628 3289 1662
rect 3323 1628 3357 1662
rect 3391 1628 3425 1662
rect 3459 1628 3493 1662
rect 3527 1628 3561 1662
rect 3595 1628 3629 1662
rect 3663 1628 3697 1662
rect 3731 1628 3765 1662
rect 3799 1628 3833 1662
rect 3867 1628 3901 1662
rect 3935 1629 4007 1662
rect 3935 1628 3972 1629
rect 127 1627 3972 1628
rect 127 1564 163 1627
rect 3971 1595 3972 1627
rect 4006 1595 4007 1629
rect 127 1530 128 1564
rect 162 1530 163 1564
rect 127 1496 163 1530
rect 127 1462 128 1496
rect 162 1462 163 1496
rect 127 1428 163 1462
rect 469 1587 679 1593
rect 469 1553 483 1587
rect 517 1553 555 1587
rect 589 1553 627 1587
rect 661 1553 679 1587
rect 127 1394 128 1428
rect 162 1394 163 1428
rect 127 1360 163 1394
rect 127 1326 128 1360
rect 162 1326 163 1360
rect 127 1292 163 1326
rect 127 1258 128 1292
rect 162 1258 163 1292
rect 127 1224 163 1258
rect 127 1190 128 1224
rect 162 1190 163 1224
rect 127 1171 163 1190
rect 127 1122 128 1171
rect 162 1122 163 1171
rect 127 1099 163 1122
rect 127 1054 128 1099
rect 162 1054 163 1099
rect 127 1027 163 1054
rect 127 986 128 1027
rect 162 986 163 1027
rect 127 955 163 986
rect 127 918 128 955
rect 162 918 163 955
rect 127 884 163 918
rect 127 849 128 884
rect 162 849 163 884
rect 127 816 163 849
rect 127 777 128 816
rect 162 777 163 816
rect 127 748 163 777
rect 201 1431 307 1437
rect 235 1397 273 1431
rect 201 1114 307 1397
rect 469 1431 679 1553
rect 1683 1587 1793 1593
rect 1683 1553 1685 1587
rect 1719 1553 1757 1587
rect 1791 1553 1793 1587
rect 1523 1513 1629 1519
rect 1557 1479 1595 1513
rect 1331 1452 1483 1468
rect 469 1397 483 1431
rect 517 1397 555 1431
rect 589 1397 627 1431
rect 661 1397 679 1431
rect 744 1418 760 1452
rect 794 1418 828 1452
rect 862 1418 909 1452
rect 1331 1433 1365 1452
rect 1399 1433 1433 1452
rect 1467 1433 1483 1452
rect 201 1080 245 1114
rect 279 1080 307 1114
rect 201 1042 307 1080
rect 201 1008 245 1042
rect 279 1008 307 1042
rect 201 766 307 1008
rect 127 705 128 748
rect 162 705 163 748
rect 127 680 163 705
rect 261 716 295 732
rect 261 658 295 682
rect 235 648 273 658
rect 235 624 261 648
rect 261 598 295 614
rect 341 584 435 1308
rect 363 550 401 584
rect 341 544 435 550
rect 469 732 523 1397
rect 557 1036 591 1074
rect 625 732 679 1397
rect 875 1308 909 1418
rect 1263 1399 1301 1433
rect 1335 1418 1365 1433
rect 1407 1418 1433 1433
rect 1335 1399 1373 1418
rect 1407 1399 1445 1418
rect 1479 1399 1483 1433
rect 977 1357 1011 1395
rect 747 766 909 1308
rect 469 641 679 732
rect 127 510 163 528
rect 127 460 128 510
rect 162 476 200 510
rect 162 460 163 476
rect 127 426 163 460
rect 127 392 128 426
rect 162 392 163 426
rect 127 358 163 392
rect 127 324 128 358
rect 162 324 163 358
rect 127 290 163 324
rect 127 256 128 290
rect 162 256 163 290
rect 127 222 163 256
rect 127 188 128 222
rect 162 188 163 222
rect 127 154 163 188
rect 245 200 375 416
rect 469 214 591 641
rect 645 584 751 590
rect 679 550 717 584
rect 1065 585 1099 623
rect 1175 585 1209 623
rect 245 166 257 200
rect 291 166 329 200
rect 363 166 375 200
rect 245 160 375 166
rect 645 200 751 550
rect 679 166 717 200
rect 1419 186 1483 1399
rect 1523 214 1629 1479
rect 1683 214 1793 1553
rect 1967 1587 2167 1593
rect 1967 1553 1978 1587
rect 2012 1553 2050 1587
rect 2084 1553 2122 1587
rect 2156 1553 2167 1587
rect 1827 1513 1933 1519
rect 1861 1479 1899 1513
rect 1827 416 1933 1479
rect 1967 766 2167 1553
rect 2341 1587 2451 1593
rect 2341 1553 2343 1587
rect 2377 1553 2415 1587
rect 2449 1553 2451 1587
rect 2201 1510 2307 1519
rect 2235 1476 2273 1510
rect 1967 716 2001 732
rect 1967 657 2001 682
rect 1967 585 2001 614
rect 2133 716 2167 732
rect 2133 657 2167 682
rect 2133 585 2167 614
rect 2050 526 2084 542
rect 2050 467 2084 476
rect 2201 416 2307 1476
rect 1827 214 2029 416
rect 2105 214 2307 416
rect 2341 214 2451 1553
rect 3543 1587 3653 1593
rect 3543 1553 3545 1587
rect 3579 1553 3617 1587
rect 3651 1553 3653 1587
rect 2505 1510 2611 1519
rect 2539 1476 2577 1510
rect 2505 214 2611 1476
rect 2651 1452 2803 1468
rect 2651 1418 2667 1452
rect 2701 1418 2735 1452
rect 2769 1418 2803 1452
rect 3191 1452 3343 1468
rect 3191 1433 3225 1452
rect 3259 1433 3293 1452
rect 2651 1402 2803 1418
rect 2651 1117 2715 1402
rect 3209 1418 3225 1433
rect 3281 1418 3293 1433
rect 3327 1418 3343 1452
rect 3209 1399 3247 1418
rect 3281 1399 3343 1418
rect 2651 1083 2666 1117
rect 2700 1083 2715 1117
rect 2651 1045 2715 1083
rect 2651 1011 2666 1045
rect 2700 1011 2715 1045
rect 2837 1045 2871 1083
rect 3279 1043 3343 1399
rect 645 160 751 166
rect 791 170 943 186
rect 127 120 128 154
rect 162 120 163 154
rect 791 136 807 170
rect 841 136 875 170
rect 909 136 943 170
rect 791 120 943 136
rect 1331 180 1483 186
rect 2651 186 2715 1011
rect 3279 1009 3294 1043
rect 3328 1009 3343 1043
rect 2925 585 2959 623
rect 3035 585 3069 623
rect 3279 186 3343 1009
rect 3383 1194 3489 1308
rect 3417 1160 3455 1194
rect 3383 214 3489 1160
rect 3543 214 3653 1553
rect 3827 1587 3933 1593
rect 3861 1553 3899 1587
rect 3827 1427 3933 1553
rect 3827 1393 3871 1427
rect 3905 1393 3933 1427
rect 3827 1355 3933 1393
rect 3827 1321 3871 1355
rect 3905 1321 3933 1355
rect 3687 1194 3793 1308
rect 3721 1160 3759 1194
rect 3687 416 3793 1160
rect 3827 766 3933 1321
rect 3971 1561 4007 1595
rect 3971 1527 3972 1561
rect 4006 1527 4007 1561
rect 3971 1493 4007 1527
rect 3971 1459 3972 1493
rect 4006 1459 4007 1493
rect 3971 1425 4007 1459
rect 3971 1391 3972 1425
rect 4006 1391 4007 1425
rect 3971 1357 4007 1391
rect 3971 1323 3972 1357
rect 4006 1323 4007 1357
rect 3971 1289 4007 1323
rect 3971 1255 3972 1289
rect 4006 1255 4007 1289
rect 3971 1221 4007 1255
rect 3971 1187 3972 1221
rect 4006 1187 4007 1221
rect 3971 1153 4007 1187
rect 3971 1119 3972 1153
rect 4006 1119 4007 1153
rect 3971 1085 4007 1119
rect 3971 1051 3972 1085
rect 4006 1051 4007 1085
rect 3971 1027 4007 1051
rect 3971 983 3972 1027
rect 4006 983 4007 1027
rect 3971 955 4007 983
rect 3971 915 3972 955
rect 4006 915 4007 955
rect 3971 883 4007 915
rect 3971 847 3972 883
rect 4006 847 4007 883
rect 3971 813 4007 847
rect 3971 777 3972 813
rect 4006 777 4007 813
rect 3971 739 4007 777
rect 3827 716 3861 732
rect 3827 657 3861 682
rect 3971 705 3972 739
rect 4006 705 4007 739
rect 3971 680 4007 705
rect 3827 585 3861 614
rect 3971 510 4007 528
rect 3934 476 3972 510
rect 3971 453 3972 476
rect 4006 453 4007 510
rect 3971 419 4007 453
rect 3687 214 3889 416
rect 3971 385 3972 419
rect 4006 385 4007 419
rect 3971 351 4007 385
rect 3971 317 3972 351
rect 4006 317 4007 351
rect 3971 283 4007 317
rect 3971 249 3972 283
rect 4006 249 4007 283
rect 3971 215 4007 249
rect 2651 180 2803 186
rect 1331 120 1972 180
rect 2162 120 2803 180
rect 3191 180 3343 186
rect 3971 181 3972 215
rect 4006 181 4007 215
rect 3191 120 3832 180
rect 3971 147 4007 181
rect 127 46 163 120
rect 3971 113 3972 147
rect 4006 113 4007 147
rect 3971 79 4007 113
rect 3971 47 3972 79
rect 212 46 3972 47
rect 127 12 161 46
rect 195 12 229 46
rect 263 12 297 46
rect 331 12 365 46
rect 399 12 433 46
rect 467 12 501 46
rect 535 12 569 46
rect 603 12 637 46
rect 671 12 705 46
rect 739 12 773 46
rect 807 12 841 46
rect 875 12 909 46
rect 943 12 977 46
rect 1011 12 1045 46
rect 1079 12 1113 46
rect 1147 12 1181 46
rect 1215 12 1249 46
rect 1283 12 1317 46
rect 1351 12 1385 46
rect 1419 12 1453 46
rect 1487 12 1521 46
rect 1555 12 1589 46
rect 1623 12 1657 46
rect 1691 12 1725 46
rect 1759 12 1793 46
rect 1827 12 1861 46
rect 1895 12 1929 46
rect 1963 12 1997 46
rect 2031 12 2065 46
rect 2099 12 2133 46
rect 2167 12 2201 46
rect 2235 12 2269 46
rect 2303 12 2337 46
rect 2371 12 2405 46
rect 2439 12 2473 46
rect 2507 12 2541 46
rect 2575 12 2609 46
rect 2643 12 2677 46
rect 2711 12 2745 46
rect 2779 12 2813 46
rect 2847 12 2881 46
rect 2915 12 2949 46
rect 2983 12 3017 46
rect 3051 12 3085 46
rect 3119 12 3153 46
rect 3187 12 3221 46
rect 3255 12 3289 46
rect 3323 12 3357 46
rect 3391 12 3425 46
rect 3459 12 3493 46
rect 3527 12 3561 46
rect 3595 12 3629 46
rect 3663 12 3697 46
rect 3731 12 3765 46
rect 3799 12 3833 46
rect 3867 12 3901 46
rect 3935 45 3972 46
rect 4006 45 4007 79
rect 3935 12 4007 45
rect 127 11 4007 12
<< viali >>
rect 483 1553 517 1587
rect 555 1553 589 1587
rect 627 1553 661 1587
rect 128 1156 162 1171
rect 128 1137 162 1156
rect 128 1088 162 1099
rect 128 1065 162 1088
rect 128 1020 162 1027
rect 128 993 162 1020
rect 128 952 162 955
rect 128 921 162 952
rect 128 850 162 883
rect 128 849 162 850
rect 128 782 162 811
rect 128 777 162 782
rect 201 1397 235 1431
rect 273 1397 307 1431
rect 1685 1553 1719 1587
rect 1757 1553 1791 1587
rect 1523 1479 1557 1513
rect 1595 1479 1629 1513
rect 483 1397 517 1431
rect 555 1397 589 1431
rect 627 1397 661 1431
rect 245 1080 279 1114
rect 245 1008 279 1042
rect 128 714 162 739
rect 128 705 162 714
rect 201 624 235 658
rect 273 648 307 658
rect 273 624 295 648
rect 295 624 307 648
rect 329 550 363 584
rect 401 550 435 584
rect 557 1074 591 1108
rect 557 1002 591 1036
rect 977 1395 1011 1429
rect 1229 1399 1263 1433
rect 1301 1399 1335 1433
rect 1373 1418 1399 1433
rect 1399 1418 1407 1433
rect 1445 1418 1467 1433
rect 1467 1418 1479 1433
rect 1373 1399 1407 1418
rect 1445 1399 1479 1418
rect 977 1323 1011 1357
rect 128 494 162 510
rect 128 476 162 494
rect 200 476 234 510
rect 1065 623 1099 657
rect 645 550 679 584
rect 717 550 751 584
rect 1065 551 1099 585
rect 1175 623 1209 657
rect 1175 551 1209 585
rect 257 166 291 200
rect 329 166 363 200
rect 645 166 679 200
rect 717 166 751 200
rect 1978 1553 2012 1587
rect 2050 1553 2084 1587
rect 2122 1553 2156 1587
rect 1827 1479 1861 1513
rect 1899 1479 1933 1513
rect 2343 1553 2377 1587
rect 2415 1553 2449 1587
rect 2201 1476 2235 1510
rect 2273 1476 2307 1510
rect 1967 648 2001 657
rect 1967 623 2001 648
rect 1967 551 2001 585
rect 2133 648 2167 657
rect 2133 623 2167 648
rect 2133 551 2167 585
rect 2050 492 2084 510
rect 2050 476 2084 492
rect 3545 1553 3579 1587
rect 3617 1553 3651 1587
rect 2505 1476 2539 1510
rect 2577 1476 2611 1510
rect 3175 1399 3209 1433
rect 3247 1418 3259 1433
rect 3259 1418 3281 1433
rect 3247 1399 3281 1418
rect 2666 1083 2700 1117
rect 2666 1011 2700 1045
rect 2837 1083 2871 1117
rect 2837 1011 2871 1045
rect 3116 1009 3150 1043
rect 3294 1009 3328 1043
rect 2925 623 2959 657
rect 2925 551 2959 585
rect 3035 623 3069 657
rect 3035 551 3069 585
rect 3383 1160 3417 1194
rect 3455 1160 3489 1194
rect 3827 1553 3861 1587
rect 3899 1553 3933 1587
rect 3871 1393 3905 1427
rect 3871 1321 3905 1355
rect 3687 1160 3721 1194
rect 3759 1160 3793 1194
rect 3972 1017 4006 1027
rect 3972 993 4006 1017
rect 3972 949 4006 955
rect 3972 921 4006 949
rect 3972 881 4006 883
rect 3972 849 4006 881
rect 3972 779 4006 811
rect 3972 777 4006 779
rect 3972 705 4006 739
rect 3827 648 3861 657
rect 3827 623 3861 648
rect 3827 551 3861 585
rect 3900 476 3934 510
rect 3972 487 4006 510
rect 3972 476 4006 487
<< metal1 >>
rect 0 1621 398 1673
rect 450 1621 462 1673
rect 514 1621 520 1673
rect 611 1668 1302 1674
rect 1296 1622 1302 1668
rect 1354 1622 1366 1674
rect 1418 1668 3981 1674
rect 1418 1622 1424 1668
rect 0 1587 2513 1593
rect 2515 1592 2551 1593
rect 0 1553 483 1587
rect 517 1553 555 1587
rect 589 1553 627 1587
rect 661 1553 1685 1587
rect 1719 1553 1757 1587
rect 1791 1553 1978 1587
rect 2012 1553 2050 1587
rect 2084 1553 2122 1587
rect 2156 1553 2343 1587
rect 2377 1553 2415 1587
rect 2449 1553 2513 1587
rect 0 1547 2513 1553
rect 2514 1548 2552 1592
rect 2553 1587 3945 1593
rect 2553 1553 3545 1587
rect 3579 1553 3617 1587
rect 3651 1553 3827 1587
rect 3861 1553 3899 1587
rect 3933 1553 3945 1587
rect 2515 1547 2551 1548
rect 2553 1547 3945 1553
rect 3 1473 55 1519
rect 57 1518 93 1519
rect 56 1474 94 1518
rect 95 1513 1945 1519
rect 95 1479 1523 1513
rect 1557 1479 1595 1513
rect 1629 1479 1827 1513
rect 1861 1479 1899 1513
rect 1933 1479 1945 1513
rect 57 1473 93 1474
rect 95 1473 1945 1479
rect 2189 1510 4033 1519
rect 2189 1476 2201 1510
rect 2235 1476 2273 1510
rect 2307 1476 2505 1510
rect 2539 1476 2577 1510
rect 2611 1476 4033 1510
rect 2189 1467 4033 1476
tri 967 1437 971 1441 se
rect 971 1439 1017 1441
tri 1017 1439 1019 1441 sw
rect 971 1437 1019 1439
rect 189 1431 379 1437
rect 189 1397 201 1431
rect 235 1397 273 1431
rect 307 1397 379 1431
rect 189 1391 379 1397
rect 380 1392 381 1436
rect 417 1392 418 1436
rect 419 1431 673 1437
tri 963 1433 967 1437 se
rect 967 1433 1019 1437
tri 1019 1433 1025 1439 sw
rect 1217 1433 2946 1439
rect 419 1397 483 1431
rect 517 1397 555 1431
rect 589 1397 627 1431
rect 661 1397 673 1431
tri 959 1429 963 1433 se
rect 963 1429 1025 1433
rect 419 1391 673 1397
tri 925 1395 959 1429 se
rect 959 1395 977 1429
rect 1011 1399 1025 1429
tri 1025 1399 1059 1433 sw
rect 1217 1399 1229 1433
rect 1263 1399 1301 1433
rect 1335 1399 1373 1433
rect 1407 1399 1445 1433
rect 1479 1399 2946 1433
rect 1011 1395 1059 1399
tri 923 1393 925 1395 se
rect 925 1393 1059 1395
tri 1059 1393 1065 1399 sw
rect 1217 1393 2946 1399
tri 921 1391 923 1393 se
rect 923 1391 1065 1393
tri 893 1363 921 1391 se
rect 921 1387 1065 1391
tri 1065 1387 1071 1393 sw
tri 2934 1387 2940 1393 ne
rect 2940 1387 2946 1393
rect 2998 1387 3010 1439
rect 3062 1393 3074 1439
rect 3075 1394 3076 1438
rect 3112 1394 3113 1438
rect 3114 1433 3293 1439
rect 3114 1399 3175 1433
rect 3209 1399 3247 1433
rect 3281 1399 3293 1433
rect 3114 1393 3293 1399
rect 3368 1433 3420 1439
rect 3062 1387 3068 1393
tri 3068 1387 3074 1393 nw
tri 3367 1387 3368 1388 se
rect 921 1363 1071 1387
tri 1071 1363 1095 1387 sw
tri 3343 1363 3367 1387 se
rect 3367 1381 3368 1387
rect 3367 1369 3420 1381
rect 3367 1363 3368 1369
rect 0 1359 2924 1363
tri 2924 1359 2928 1363 sw
tri 3080 1359 3084 1363 se
rect 3084 1359 3368 1363
rect 0 1357 3368 1359
rect 0 1323 977 1357
rect 1011 1323 3368 1357
rect 0 1317 3368 1323
tri 41 1311 47 1317 ne
rect 47 1311 3420 1317
rect 3859 1427 3917 1433
rect 3859 1393 3871 1427
rect 3905 1393 3917 1427
rect 3859 1355 3917 1393
rect 3859 1321 3871 1355
rect 3905 1321 3917 1355
rect 3859 1315 3917 1321
rect 3957 1432 4021 1433
rect 3957 1380 3963 1432
rect 4015 1380 4021 1432
rect 3957 1368 4021 1380
rect 3957 1316 3963 1368
rect 4015 1316 4021 1368
rect 3957 1315 4021 1316
rect 0 1283 28 1289
tri 28 1283 34 1289 sw
rect 0 1243 4033 1283
tri 0 1231 12 1243 ne
rect 12 1231 4033 1243
rect 459 1197 563 1203
rect 122 1171 168 1183
rect 122 1137 128 1171
rect 162 1137 168 1171
rect 122 1099 168 1137
rect 511 1151 563 1197
rect 564 1152 565 1202
rect 601 1152 602 1202
rect 603 1194 3805 1203
rect 603 1160 3383 1194
rect 3417 1160 3455 1194
rect 3489 1160 3687 1194
rect 3721 1160 3759 1194
rect 3793 1160 3805 1194
rect 603 1151 3805 1160
rect 459 1133 511 1145
rect 122 1065 128 1099
rect 162 1065 168 1099
rect 122 1027 168 1065
rect 122 993 128 1027
rect 162 996 168 1027
rect 239 1114 285 1126
rect 239 1080 245 1114
rect 279 1080 285 1114
rect 239 1045 285 1080
tri 511 1126 536 1151 nw
rect 2654 1117 4033 1123
rect 459 1075 511 1081
rect 545 1108 630 1114
rect 632 1113 668 1114
rect 545 1074 557 1108
rect 591 1074 630 1108
tri 285 1045 309 1069 sw
tri 521 1045 545 1069 se
rect 545 1068 630 1074
rect 631 1069 669 1113
rect 632 1068 668 1069
rect 670 1068 725 1114
rect 545 1045 607 1068
tri 607 1045 630 1068 nw
tri 670 1045 693 1068 ne
rect 693 1045 725 1068
rect 239 1044 309 1045
tri 309 1044 310 1045 sw
tri 520 1044 521 1045 se
rect 521 1044 603 1045
rect 239 1042 603 1044
rect 239 1008 245 1042
rect 279 1036 603 1042
tri 603 1041 607 1045 nw
tri 693 1041 697 1045 ne
rect 279 1008 557 1036
rect 239 1002 557 1008
rect 591 1002 603 1036
tri 168 996 169 997 sw
rect 239 996 603 1002
rect 162 995 169 996
tri 169 995 170 996 sw
rect 162 993 170 995
tri 170 993 172 995 sw
tri 695 993 697 995 se
rect 697 993 725 1045
rect 2654 1083 2666 1117
rect 2700 1083 2837 1117
rect 2871 1083 4033 1117
rect 2654 1077 4033 1083
rect 2654 1049 2927 1077
tri 2927 1049 2955 1077 nw
rect 2654 1045 2921 1049
rect 2654 1011 2666 1045
rect 2700 1011 2837 1045
rect 2871 1043 2921 1045
tri 2921 1043 2927 1049 nw
rect 3104 1043 3358 1049
rect 3360 1048 3396 1049
rect 2871 1011 2887 1043
rect 2654 1009 2887 1011
tri 2887 1009 2921 1043 nw
rect 3104 1009 3116 1043
rect 3150 1009 3294 1043
rect 3328 1009 3358 1043
rect 2654 1005 2883 1009
tri 2883 1005 2887 1009 nw
rect 3104 1003 3358 1009
rect 3359 1004 3397 1048
rect 3360 1003 3396 1004
rect 3398 1003 3517 1049
tri 3954 1027 3966 1039 se
rect 3966 1027 4012 1039
tri 3930 1003 3954 1027 se
rect 3954 1003 3972 1027
tri 3447 995 3455 1003 ne
rect 3455 995 3517 1003
tri 3922 995 3930 1003 se
rect 3930 995 3972 1003
tri 725 993 727 995 sw
tri 3455 993 3457 995 ne
rect 3457 993 3517 995
tri 3920 993 3922 995 se
rect 3922 993 3972 995
rect 4006 993 4012 1027
rect 122 968 172 993
tri 172 968 197 993 sw
tri 670 968 695 993 se
rect 695 968 727 993
tri 727 968 752 993 sw
tri 3457 978 3472 993 ne
rect 122 955 3364 968
tri 3364 955 3377 968 sw
rect 122 921 128 955
rect 162 944 3377 955
tri 3377 944 3388 955 sw
rect 162 921 3388 944
tri 3388 921 3411 944 sw
tri 3449 921 3472 944 se
rect 3472 921 3517 993
tri 3895 968 3920 993 se
rect 3920 968 4012 993
tri 3612 955 3625 968 se
rect 3625 955 4012 968
tri 3601 944 3612 955 se
rect 3612 944 3972 955
tri 3517 921 3540 944 sw
tri 3578 921 3601 944 se
rect 3601 921 3972 944
rect 4006 921 4012 955
rect 122 919 3411 921
tri 3411 919 3413 921 sw
tri 3447 919 3449 921 se
rect 3449 919 3540 921
tri 3540 919 3542 921 sw
tri 3576 919 3578 921 se
rect 3578 919 4012 921
rect 122 883 4012 919
rect 122 849 128 883
rect 162 849 3972 883
rect 4006 849 4012 883
rect 122 811 4012 849
rect 122 777 128 811
rect 162 777 3972 811
rect 4006 777 4012 811
rect 122 739 4012 777
rect 122 705 128 739
rect 162 705 3972 739
rect 4006 705 4012 739
rect 122 692 4012 705
rect 122 590 150 692
tri 150 665 177 692 nw
rect 189 658 1111 664
rect 189 624 201 658
rect 235 624 273 658
rect 307 657 1111 658
rect 307 624 1065 657
rect 189 623 1065 624
rect 1099 623 1111 657
rect 189 618 1111 623
tri 1028 617 1029 618 ne
rect 1029 617 1111 618
tri 150 590 177 617 sw
tri 1029 593 1053 617 ne
rect 122 544 202 590
rect 204 589 240 590
rect 203 545 241 589
rect 242 584 541 590
rect 242 550 329 584
rect 363 550 401 584
rect 435 550 541 584
rect 204 544 240 545
rect 242 544 541 550
rect 542 545 543 589
rect 579 545 580 589
rect 581 584 763 590
rect 581 550 645 584
rect 679 550 717 584
rect 751 550 763 584
rect 581 544 763 550
rect 1053 585 1111 617
rect 1053 551 1065 585
rect 1099 551 1111 585
rect 1053 545 1111 551
rect 1163 657 2013 664
rect 1163 623 1175 657
rect 1209 623 1967 657
rect 2001 623 2013 657
rect 1163 618 2013 623
rect 1163 585 1221 618
tri 1221 593 1246 618 nw
tri 1930 593 1955 618 ne
rect 1163 551 1175 585
rect 1209 551 1221 585
rect 1163 545 1221 551
rect 1955 585 2013 618
rect 1955 551 1967 585
rect 2001 551 2013 585
rect 1955 545 2013 551
rect 2121 657 2971 664
rect 2121 623 2133 657
rect 2167 623 2925 657
rect 2959 623 2971 657
rect 2121 618 2971 623
rect 2121 585 2179 618
tri 2179 593 2204 618 nw
tri 2888 593 2913 618 ne
rect 2121 551 2133 585
rect 2167 551 2179 585
rect 2121 545 2179 551
rect 2913 585 2971 618
rect 2913 551 2925 585
rect 2959 551 2971 585
rect 2913 545 2971 551
rect 3023 657 3081 663
rect 3023 623 3035 657
rect 3069 623 3081 657
rect 3023 591 3081 623
rect 3815 657 3873 663
rect 3815 623 3827 657
rect 3861 623 3873 657
tri 3081 591 3106 616 sw
tri 3790 591 3815 616 se
rect 3815 591 3873 623
rect 3023 585 3873 591
rect 3023 551 3035 585
rect 3069 551 3827 585
rect 3861 551 3873 585
rect 3023 545 3873 551
tri 1489 516 1495 522 se
rect 1495 516 1501 522
rect 0 510 1501 516
rect 0 476 128 510
rect 162 476 200 510
rect 234 476 1501 510
rect 0 470 1501 476
rect 1553 470 1565 522
rect 1617 516 1623 522
tri 1623 516 1629 522 sw
rect 1617 510 4033 516
rect 1617 476 2050 510
rect 2084 476 3900 510
rect 3934 476 3972 510
rect 4006 476 4033 510
rect 1617 470 4033 476
rect 82 454 4033 470
rect 82 402 1501 454
rect 1553 402 1565 454
rect 1617 420 4033 454
rect 1617 402 2270 420
rect 82 376 2270 402
rect 82 324 1501 376
rect 1553 324 1565 376
rect 1617 324 2270 376
rect 82 298 2270 324
rect 82 246 1501 298
rect 1553 246 1565 298
rect 1617 246 2270 298
rect 82 240 2270 246
rect 2386 368 3768 420
rect 3820 368 4033 420
rect 2386 356 4033 368
rect 2386 304 3768 356
rect 3820 304 4033 356
rect 2386 240 4033 304
tri 3953 206 3987 240 ne
rect 3987 206 4033 240
rect 0 200 763 206
rect 0 166 257 200
rect 291 166 329 200
rect 363 166 645 200
rect 679 166 717 200
rect 751 166 763 200
rect 0 160 763 166
tri 3987 160 4033 206 ne
rect 0 80 4033 132
rect 0 6 130 52
rect 1495 6 1501 52
rect 0 0 1501 6
rect 1553 0 1565 52
rect 1617 6 1623 52
rect 1959 6 1965 52
rect 1617 0 1965 6
rect 2017 0 2029 52
rect 2081 0 2093 52
rect 2145 0 2157 52
rect 2209 0 2221 52
rect 2273 6 2331 52
rect 3114 6 3120 52
rect 2273 0 3120 6
rect 3172 0 3184 52
rect 3236 0 3248 52
rect 3300 0 3312 52
rect 3364 0 3376 52
rect 3428 6 3486 52
rect 4000 6 4033 52
rect 3428 0 4033 6
<< rmetal1 >>
rect 2513 1592 2515 1593
rect 2551 1592 2553 1593
rect 2513 1548 2514 1592
rect 2552 1548 2553 1592
rect 2513 1547 2515 1548
rect 2551 1547 2553 1548
rect 55 1518 57 1519
rect 93 1518 95 1519
rect 55 1474 56 1518
rect 94 1474 95 1518
rect 55 1473 57 1474
rect 93 1473 95 1474
rect 379 1436 381 1437
rect 379 1392 380 1436
rect 379 1391 381 1392
rect 417 1436 419 1437
rect 418 1392 419 1436
rect 417 1391 419 1392
rect 3074 1438 3076 1439
rect 3074 1394 3075 1438
rect 3074 1393 3076 1394
rect 3112 1438 3114 1439
rect 3113 1394 3114 1438
rect 3112 1393 3114 1394
rect 563 1202 565 1203
rect 563 1152 564 1202
rect 563 1151 565 1152
rect 601 1202 603 1203
rect 602 1152 603 1202
rect 601 1151 603 1152
rect 630 1113 632 1114
rect 668 1113 670 1114
rect 630 1069 631 1113
rect 669 1069 670 1113
rect 630 1068 632 1069
rect 668 1068 670 1069
rect 3358 1048 3360 1049
rect 3396 1048 3398 1049
rect 3358 1004 3359 1048
rect 3397 1004 3398 1048
rect 3358 1003 3360 1004
rect 3396 1003 3398 1004
rect 202 589 204 590
rect 240 589 242 590
rect 202 545 203 589
rect 241 545 242 589
rect 541 589 543 590
rect 202 544 204 545
rect 240 544 242 545
rect 541 545 542 589
rect 541 544 543 545
rect 579 589 581 590
rect 580 545 581 589
rect 579 544 581 545
<< via1 >>
rect 398 1621 450 1673
rect 462 1621 514 1673
rect 1302 1622 1354 1674
rect 1366 1622 1418 1674
rect 2946 1387 2998 1439
rect 3010 1387 3062 1439
rect 3368 1381 3420 1433
rect 3368 1317 3420 1369
rect 3963 1380 4015 1432
rect 3963 1316 4015 1368
rect 459 1145 511 1197
rect 459 1081 511 1133
rect 1501 470 1553 522
rect 1565 470 1617 522
rect 1501 402 1553 454
rect 1565 402 1617 454
rect 1501 324 1553 376
rect 1565 324 1617 376
rect 1501 246 1553 298
rect 1565 246 1617 298
rect 2270 240 2386 420
rect 3768 368 3820 420
rect 3768 304 3820 356
rect 1501 0 1553 52
rect 1565 0 1617 52
rect 1965 0 2017 52
rect 2029 0 2081 52
rect 2093 0 2145 52
rect 2157 0 2209 52
rect 2221 0 2273 52
rect 3120 0 3172 52
rect 3184 0 3236 52
rect 3248 0 3300 52
rect 3312 0 3364 52
rect 3376 0 3428 52
<< metal2 >>
tri 450 1689 459 1698 se
rect 459 1689 511 1698
rect 82 72 284 1689
rect 312 72 364 1689
tri 441 1680 450 1689 se
rect 450 1680 511 1689
tri 511 1680 520 1689 sw
tri 435 1674 441 1680 se
rect 441 1674 520 1680
tri 434 1673 435 1674 se
rect 435 1673 520 1674
rect 392 1621 398 1673
rect 450 1621 462 1673
rect 514 1621 520 1673
tri 434 1596 459 1621 ne
rect 459 1614 520 1621
rect 459 1197 511 1614
tri 511 1605 520 1614 nw
rect 459 1133 511 1145
rect 459 72 511 1081
rect 571 72 623 1689
rect 729 605 1229 1689
rect 1285 1674 1435 1689
rect 1285 1622 1302 1674
rect 1354 1622 1366 1674
rect 1418 1622 1435 1674
rect 1285 622 1435 1622
rect 729 526 1150 605
tri 1150 526 1229 605 nw
rect 729 522 1146 526
tri 1146 522 1150 526 nw
rect 1494 522 1624 1689
rect 729 470 1094 522
tri 1094 470 1146 522 nw
rect 1494 470 1501 522
rect 1553 470 1565 522
rect 1617 470 1624 522
rect 729 72 1091 470
tri 1091 467 1094 470 nw
rect 1119 72 1435 455
rect 1494 454 1624 470
rect 1494 402 1501 454
rect 1553 402 1565 454
rect 1617 402 1624 454
rect 1494 376 1624 402
rect 1494 324 1501 376
rect 1553 324 1565 376
rect 1617 324 1624 376
rect 1494 298 1624 324
rect 1494 246 1501 298
rect 1553 246 1565 298
rect 1617 246 1624 298
rect 1494 52 1624 246
rect 1680 270 1996 1689
rect 2142 856 2410 1689
tri 2142 795 2203 856 ne
rect 2203 795 2410 856
tri 2203 745 2253 795 ne
tri 1680 240 1710 270 ne
rect 1710 240 1996 270
tri 1710 232 1718 240 ne
rect 1718 232 1996 240
rect 2253 420 2410 795
rect 2253 240 2270 420
rect 2386 240 2410 420
tri 1718 149 1801 232 ne
rect 1801 196 1996 232
tri 1996 196 2032 232 sw
rect 1801 149 2032 196
tri 2032 149 2079 196 sw
tri 2206 149 2253 196 se
rect 2253 149 2410 240
tri 1801 72 1878 149 ne
rect 1878 72 2410 149
rect 2466 1515 2734 1689
tri 2734 1515 2908 1689 sw
rect 2466 1511 2908 1515
tri 2908 1511 2912 1515 sw
rect 2466 72 2912 1511
tri 2940 1439 3016 1515 se
rect 3016 1439 3068 1689
rect 2940 1387 2946 1439
rect 2998 1387 3010 1439
rect 3062 1387 3068 1439
rect 3114 522 3340 1689
rect 3368 1433 3420 1689
rect 3368 1369 3420 1381
rect 3368 1311 3420 1317
tri 3340 522 3344 526 sw
tri 3444 522 3448 526 se
rect 3448 522 3542 1689
tri 3679 1432 3680 1433 se
rect 3680 1432 3732 1689
tri 3627 1380 3679 1432 se
rect 3679 1412 3732 1432
rect 3679 1404 3724 1412
tri 3724 1404 3732 1412 nw
rect 3679 1380 3700 1404
tri 3700 1380 3724 1404 nw
tri 3746 1383 3767 1404 se
rect 3767 1383 3819 1689
tri 3743 1380 3746 1383 se
rect 3746 1380 3816 1383
tri 3816 1380 3819 1383 nw
rect 3847 1432 4030 1689
rect 3847 1380 3963 1432
rect 4015 1380 4030 1432
tri 3615 1368 3627 1380 se
rect 3627 1368 3688 1380
tri 3688 1368 3700 1380 nw
tri 3731 1368 3743 1380 se
rect 3743 1368 3804 1380
tri 3804 1368 3816 1380 nw
rect 3847 1368 4030 1380
tri 3610 1363 3615 1368 se
rect 3615 1363 3683 1368
tri 3683 1363 3688 1368 nw
tri 3726 1363 3731 1368 se
rect 3731 1363 3799 1368
tri 3799 1363 3804 1368 nw
tri 3607 1360 3610 1363 se
rect 3610 1360 3680 1363
tri 3680 1360 3683 1363 nw
tri 3723 1360 3726 1363 se
rect 3726 1360 3796 1363
tri 3796 1360 3799 1363 nw
tri 3597 1350 3607 1360 se
rect 3607 1354 3674 1360
tri 3674 1354 3680 1360 nw
tri 3717 1354 3723 1360 se
rect 3723 1354 3786 1360
rect 3607 1350 3670 1354
tri 3670 1350 3674 1354 nw
tri 3713 1350 3717 1354 se
rect 3717 1350 3786 1354
tri 3786 1350 3796 1360 nw
rect 3114 501 3344 522
tri 3344 501 3365 522 sw
tri 3423 501 3444 522 se
rect 3444 501 3542 522
rect 3114 128 3542 501
rect 3114 72 3486 128
tri 3486 72 3542 128 nw
tri 3587 1340 3597 1350 se
rect 3597 1340 3660 1350
tri 3660 1340 3670 1350 nw
tri 3703 1340 3713 1350 se
rect 3713 1340 3776 1350
tri 3776 1340 3786 1350 nw
tri 3837 1340 3847 1350 se
rect 3847 1340 3963 1368
rect 3587 72 3639 1340
tri 3639 1319 3660 1340 nw
tri 3682 1319 3703 1340 se
rect 3703 1319 3755 1340
tri 3755 1319 3776 1340 nw
tri 3816 1319 3837 1340 se
rect 3837 1319 3963 1340
tri 3679 1316 3682 1319 se
rect 3682 1316 3752 1319
tri 3752 1316 3755 1319 nw
tri 3813 1316 3816 1319 se
rect 3816 1316 3963 1319
rect 4015 1316 4030 1368
tri 3674 1311 3679 1316 se
rect 3679 1311 3738 1316
rect 3674 1302 3738 1311
tri 3738 1302 3752 1316 nw
tri 3799 1302 3813 1316 se
rect 3813 1302 4030 1316
rect 3674 267 3726 1302
tri 3726 1290 3738 1302 nw
tri 3787 1290 3799 1302 se
rect 3799 1290 4030 1302
tri 3762 1265 3787 1290 se
rect 3787 1265 4030 1290
rect 3762 420 4030 1265
rect 3762 368 3768 420
rect 3820 368 4030 420
rect 3762 356 4030 368
rect 3762 304 3768 356
rect 3820 304 4030 356
rect 3762 291 4030 304
tri 3762 270 3783 291 ne
rect 3783 270 4030 291
tri 3726 267 3729 270 sw
tri 3783 267 3786 270 ne
rect 3786 267 4030 270
rect 3674 251 3729 267
tri 3729 251 3745 267 sw
tri 3786 251 3802 267 ne
rect 3802 251 4030 267
rect 3674 249 3745 251
tri 3674 194 3729 249 ne
rect 3729 194 3745 249
tri 3745 194 3802 251 sw
tri 3802 194 3859 251 ne
rect 3859 194 4030 251
tri 3729 121 3802 194 ne
tri 3802 178 3818 194 sw
tri 3859 178 3875 194 ne
rect 3875 178 4030 194
rect 3802 150 3818 178
tri 3818 150 3846 178 sw
tri 3875 150 3903 178 ne
rect 3802 121 3846 150
tri 3846 121 3875 150 sw
tri 3802 100 3823 121 ne
rect 3823 72 3875 121
rect 3903 72 4030 178
rect 1494 0 1501 52
rect 1553 0 1565 52
rect 1617 0 1624 52
rect 1959 0 1965 52
rect 2017 0 2029 52
rect 2081 0 2093 52
rect 2145 0 2157 52
rect 2209 0 2221 52
rect 2273 0 2331 52
rect 3114 0 3120 52
rect 3172 0 3184 52
rect 3236 0 3248 52
rect 3300 0 3312 52
rect 3364 0 3376 52
rect 3428 0 3486 52
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 591 0 1 1002
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 1209 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform -1 0 3861 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 2001 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 2167 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform -1 0 3069 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform -1 0 3905 0 1 1321
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 2666 0 -1 1117
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 2837 0 -1 1117
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 1065 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 2925 0 1 551
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 4006 0 1 476
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 3281 0 -1 1433
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 751 0 -1 200
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 3793 0 -1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 1791 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 1933 0 -1 1513
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 2611 0 -1 1510
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 3651 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 3933 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 0 1 977 1 0 1323
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 0 1 245 1 0 1008
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 201 0 -1 658
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 201 0 -1 1431
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 257 0 -1 200
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 1523 0 -1 1513
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 3383 0 -1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 2201 0 -1 1510
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 2343 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 329 0 -1 584
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 645 0 -1 584
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 128 0 1 476
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 1 0 483 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 1 0 483 0 -1 1431
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 1 0 1978 0 -1 1587
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 0 1 3972 1 0 705
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 1 0 1229 0 -1 1433
box 0 0 1 1
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1707688321
transform 0 1 128 1 0 705
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 2084 0 1 476
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 1 0 3294 0 -1 1043
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1707688321
transform 1 0 3116 0 -1 1043
box 0 0 1 1
use L1M1_CDNS_524688791851066  L1M1_CDNS_524688791851066_0
timestamp 1707688321
transform 1 0 142 0 1 12
box -12 -6 3862 40
use L1M1_CDNS_524688791851146  L1M1_CDNS_524688791851146_0
timestamp 1707688321
transform -1 0 3969 0 -1 1662
box -12 -6 3358 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 511 -1 0 1203
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 1623 0 1 0
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 520 0 1 1621
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform -1 0 1623 0 1 470
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 3368 1 0 1311
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 1 0 1296 0 -1 1674
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 1 0 2940 0 -1 1439
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 1 0 2264 0 1 240
box 0 0 1 1
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1707688321
transform 1 0 1296 0 1 692
box 0 0 128 244
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 1 0 3762 0 -1 420
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 1 0 3957 0 -1 1432
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform -1 0 4024 0 1 240
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 1 0 83 0 1 240
box 0 0 192 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1707688321
transform 1 0 1710 0 1 240
box 0 0 256 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1707688321
transform 1 0 3131 0 1 240
box 0 0 384 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_1
timestamp 1707688321
transform 1 0 2497 0 1 240
box 0 0 384 180
use nfet_CDNS_524688791851149  nfet_CDNS_524688791851149_0
timestamp 1707688321
transform -1 0 1984 0 1 218
box -79 -26 495 226
use nfet_CDNS_524688791851149  nfet_CDNS_524688791851149_1
timestamp 1707688321
transform -1 0 3844 0 1 218
box -79 -26 495 226
use nfet_CDNS_524688791851149  nfet_CDNS_524688791851149_2
timestamp 1707688321
transform 1 0 290 0 1 218
box -79 -26 495 226
use nfet_CDNS_524688791851149  nfet_CDNS_524688791851149_3
timestamp 1707688321
transform 1 0 2150 0 1 218
box -79 -26 495 226
use pfet_CDNS_524688791851147  pfet_CDNS_524688791851147_0
timestamp 1707688321
transform -1 0 878 0 1 770
box -119 -66 239 666
use pfet_CDNS_524688791851147  pfet_CDNS_524688791851147_1
timestamp 1707688321
transform -1 0 2738 0 1 770
box -119 -66 239 666
use pfet_CDNS_524688791851147  pfet_CDNS_524688791851147_2
timestamp 1707688321
transform 1 0 1396 0 1 770
box -119 -66 239 666
use pfet_CDNS_524688791851148  pfet_CDNS_524688791851148_0
timestamp 1707688321
transform -1 0 1984 0 1 770
box -119 -66 531 666
use pfet_CDNS_524688791851148  pfet_CDNS_524688791851148_1
timestamp 1707688321
transform -1 0 3844 0 1 770
box -119 -66 531 666
use pfet_CDNS_524688791851148  pfet_CDNS_524688791851148_2
timestamp 1707688321
transform 1 0 290 0 1 770
box -119 -66 531 666
use pfet_CDNS_524688791851148  pfet_CDNS_524688791851148_3
timestamp 1707688321
transform 1 0 2150 0 1 770
box -119 -66 531 666
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 925 -1 0 186
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 -1 2785 -1 0 1468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 -1 878 -1 0 1468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 3209 -1 0 1468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 1 1349 -1 0 1468
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform -1 0 2017 0 1 598
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform -1 0 3877 0 1 598
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 1 0 245 0 1 598
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 1 0 2117 0 1 598
box 0 0 1 1
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 -1 1972 -1 0 186
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1707688321
transform 0 -1 3832 -1 0 186
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_2
timestamp 1707688321
transform 0 1 2162 -1 0 186
box 0 0 66 542
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_0
timestamp 1707688321
transform -1 0 471 0 -1 1437
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_1
timestamp 1707688321
transform -1 0 633 0 -1 590
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851125  sky130_fd_io__refgen_em1o_CDNS_524688791851125_2
timestamp 1707688321
transform -1 0 3166 0 -1 1439
box 0 0 1 1
use sky130_fd_io__refgen_em1o_CDNS_524688791851127  sky130_fd_io__refgen_em1o_CDNS_524688791851127_0
timestamp 1707688321
transform -1 0 655 0 -1 1203
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_0
timestamp 1707688321
transform -1 0 147 0 -1 1519
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_1
timestamp 1707688321
transform -1 0 2605 0 -1 1593
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_2
timestamp 1707688321
transform 1 0 578 0 -1 1114
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_3
timestamp 1707688321
transform 1 0 150 0 -1 590
box 0 0 1 1
use sky130_fd_io__refgen_em1s_CDNS_524688791851129  sky130_fd_io__refgen_em1s_CDNS_524688791851129_4
timestamp 1707688321
transform 1 0 3306 0 1 1003
box 0 0 1 1
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_0
timestamp 1707688321
transform -1 0 1368 0 1 99
box -107 21 267 1369
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_1
timestamp 1707688321
transform -1 0 3228 0 1 99
box -107 21 267 1369
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_2
timestamp 1707688321
transform 1 0 906 0 1 99
box -107 21 267 1369
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_3
timestamp 1707688321
transform 1 0 2766 0 1 99
box -107 21 267 1369
<< labels >>
flabel comment s 252 1417 252 1417 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 3225 1420 3225 1420 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 341 90 341 90 3 FreeSans 200 90 0 0 ibuf_sel_h_n
flabel comment s 341 1683 341 1683 3 FreeSans 200 270 0 0 ibuf_sel_h_n
flabel comment s 978 114 978 114 3 FreeSans 200 90 0 0 vpwr
flabel comment s 978 1683 978 1683 3 FreeSans 200 270 0 0 vpwr
flabel comment s 4019 1264 4019 1264 3 FreeSans 200 180 0 0 sel_vcc_io_0p4
flabel comment s 12 1264 12 1264 3 FreeSans 200 0 0 0 sel_vcc_io_0p4
flabel comment s 3966 1490 3966 1490 3 FreeSans 200 180 0 0 vohref_op5
flabel comment s 4026 106 4026 106 3 FreeSans 200 180 0 0 vinref
flabel comment s 12 107 12 107 3 FreeSans 200 0 0 0 vinref
flabel comment s 3708 1678 3708 1678 3 FreeSans 200 270 0 0 vref_sel_h
flabel comment s 3612 84 3612 84 3 FreeSans 200 90 0 0 vref_sel_h
flabel comment s 3848 84 3848 84 3 FreeSans 200 90 0 0 vref_sel_h_n
flabel comment s 3791 1685 3791 1685 3 FreeSans 200 270 0 0 vref_sel_h_n
flabel comment s 596 1683 596 1683 3 FreeSans 200 270 0 0 ibuf_sel_h
flabel comment s 597 84 597 84 3 FreeSans 200 90 0 0 ibuf_sel_h
flabel metal1 s 0 470 33 516 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 4000 470 4033 516 3 FreeSans 200 180 0 0 vgnd
port 2 nsew
flabel metal1 s 3 1473 25 1519 3 FreeSans 200 0 0 0 vohref_int
port 3 nsew
flabel metal1 s 4007 1467 4033 1519 3 FreeSans 200 180 0 0 vohref_0p5
port 4 nsew
flabel metal1 s 0 1621 25 1673 3 FreeSans 200 0 0 0 vohref
port 5 nsew
flabel metal1 s 4000 0 4033 52 3 FreeSans 200 180 0 0 vgnd
port 2 nsew
flabel metal1 s 0 0 33 52 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 0 1547 25 1593 3 FreeSans 200 0 0 0 vinref_int
port 6 nsew
flabel metal1 s 0 160 25 206 3 FreeSans 200 0 0 0 vcc_io_ref
port 9 nsew
flabel metal1 s 3971 692 3989 1039 3 FreeSans 200 180 0 0 vcc_io
port 7 nsew
flabel metal1 s 4007 1077 4033 1123 3 FreeSans 200 180 0 0 sel_vohref_0p5
port 8 nsew
flabel metal1 s 0 1317 25 1363 3 FreeSans 200 0 0 0 sel_vcc_io
port 10 nsew
flabel metal2 s 1494 80 1624 113 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 459 72 511 105 3 FreeSans 200 90 0 0 vohref
port 5 nsew
flabel metal2 s 3114 72 3486 105 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 2466 72 2912 105 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 1680 1673 1996 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 2142 1673 2410 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 82 72 284 105 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 459 1673 511 1689 3 FreeSans 200 270 0 0 vohref
port 5 nsew
flabel metal2 s 1579 1672 1579 1672 3 FreeSans 200 270 0 0 vgnd
flabel metal2 s 3016 1673 3068 1689 3 FreeSans 200 270 0 0 sel_vohref
port 11 nsew
flabel metal2 s 3368 1673 3420 1689 3 FreeSans 200 270 0 0 sel_vcc_io
port 10 nsew
flabel metal2 s 1285 1673 1435 1689 3 FreeSans 200 270 0 0 vcc_io
port 7 nsew
flabel metal2 s 3847 1673 4030 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 3448 1673 3542 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 3114 1673 3340 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 2466 1673 2734 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 82 1673 284 1689 3 FreeSans 200 270 0 0 vgnd
port 2 nsew
flabel metal2 s 2142 72 2410 105 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 1878 72 2086 105 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
<< properties >>
string GDS_END 79921328
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79887954
string path 38.975 6.000 38.975 11.500 
<< end >>
