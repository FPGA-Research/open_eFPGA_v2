magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect 119 376 375 392
rect 119 342 135 376
rect 169 342 230 376
rect 264 342 325 376
rect 359 342 375 376
rect 119 326 375 342
rect 431 376 687 392
rect 431 342 447 376
rect 481 342 542 376
rect 576 342 637 376
rect 671 342 687 376
rect 431 326 687 342
rect 119 268 253 284
rect 119 234 135 268
rect 169 234 203 268
rect 237 234 253 268
rect 119 218 253 234
rect 309 268 443 284
rect 309 234 325 268
rect 359 234 393 268
rect 427 234 443 268
rect 309 218 443 234
<< polycont >>
rect 135 342 169 376
rect 230 342 264 376
rect 325 342 359 376
rect 447 342 481 376
rect 542 342 576 376
rect 637 342 671 376
rect 135 234 169 268
rect 203 234 237 268
rect 325 234 359 268
rect 393 234 427 268
<< locali >>
rect 230 556 264 594
rect 74 460 108 498
rect 386 460 420 498
rect 540 490 578 524
rect 698 460 732 498
rect 119 342 131 376
rect 169 342 203 376
rect 264 342 325 376
rect 359 342 375 376
rect 431 342 443 376
rect 481 342 515 376
rect 576 342 637 376
rect 671 342 687 376
rect 165 268 203 278
rect 119 244 131 268
rect 119 234 135 244
rect 169 234 203 268
rect 237 234 253 268
rect 309 234 325 268
rect 380 234 393 268
rect 262 111 300 145
rect 107 24 145 58
rect 417 24 455 58
<< viali >>
rect 230 594 264 628
rect 74 498 108 532
rect 230 522 264 556
rect 74 426 108 460
rect 386 498 420 532
rect 506 490 540 524
rect 578 490 612 524
rect 698 498 732 532
rect 386 426 420 460
rect 698 426 732 460
rect 131 342 135 376
rect 135 342 165 376
rect 203 342 230 376
rect 230 342 237 376
rect 443 342 447 376
rect 447 342 477 376
rect 515 342 542 376
rect 542 342 549 376
rect 131 268 165 278
rect 203 268 237 278
rect 131 244 135 268
rect 135 244 165 268
rect 203 244 237 268
rect 346 234 359 268
rect 359 234 380 268
rect 418 234 427 268
rect 427 234 452 268
rect 228 111 262 145
rect 300 111 334 145
rect 73 24 107 58
rect 145 24 179 58
rect 383 24 417 58
rect 455 24 489 58
<< metal1 >>
rect 66 628 765 690
rect 66 594 230 628
rect 264 594 765 628
rect 66 590 765 594
tri 190 556 224 590 ne
rect 224 556 270 590
tri 270 556 304 590 nw
rect 68 532 114 544
rect 68 498 74 532
rect 108 498 114 532
rect 224 522 230 556
rect 264 522 270 556
rect 224 510 270 522
rect 380 532 426 544
rect 68 460 114 498
rect 380 498 386 532
rect 420 498 426 532
tri 114 460 134 480 sw
tri 360 460 380 480 se
rect 380 460 426 498
rect 494 481 500 533
rect 552 481 566 533
rect 618 481 624 533
rect 692 532 738 544
rect 692 498 698 532
rect 732 498 738 532
tri 426 460 446 480 sw
tri 672 460 692 480 se
rect 692 460 738 498
rect 68 426 74 460
rect 108 446 134 460
tri 134 446 148 460 sw
tri 346 446 360 460 se
rect 360 446 386 460
rect 108 426 386 446
rect 420 446 446 460
tri 446 446 460 460 sw
tri 658 446 672 460 se
rect 672 446 698 460
rect 420 426 698 446
rect 732 426 738 460
rect 68 414 738 426
rect 119 376 249 382
rect 119 342 131 376
rect 165 342 203 376
rect 237 342 249 376
rect 119 278 249 342
rect 431 376 561 382
rect 431 342 443 376
rect 477 342 515 376
rect 549 342 561 376
rect 119 244 131 278
rect 165 244 203 278
rect 237 244 249 278
tri 397 274 431 308 se
rect 431 274 561 342
rect 119 238 249 244
rect 334 268 561 274
rect 334 234 346 268
rect 380 234 418 268
rect 452 234 561 268
rect 334 228 561 234
tri 370 151 419 200 se
rect 419 151 463 200
rect 216 148 463 151
rect 515 148 527 200
rect 579 148 585 200
rect 216 145 390 148
rect 216 111 228 145
rect 262 111 300 145
rect 334 111 390 145
rect 216 105 390 111
tri 390 105 433 148 nw
rect 61 58 501 64
rect 61 24 73 58
rect 107 24 145 58
rect 179 24 383 58
rect 417 24 455 58
rect 489 24 501 58
rect 61 0 501 24
<< via1 >>
rect 500 524 552 533
rect 500 490 506 524
rect 506 490 540 524
rect 540 490 552 524
rect 500 481 552 490
rect 566 524 618 533
rect 566 490 578 524
rect 578 490 612 524
rect 612 490 618 524
rect 566 481 618 490
rect 463 148 515 200
rect 527 148 579 200
<< metal2 >>
rect 494 481 500 533
rect 552 481 566 533
rect 618 481 624 533
rect 533 200 585 481
rect 457 148 463 200
rect 515 148 527 200
rect 579 148 585 200
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_0
timestamp 1707688321
transform 1 0 309 0 1 36
box -82 -32 182 182
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_1
timestamp 1707688321
transform 1 0 153 0 1 36
box -82 -32 182 182
use pfet_CDNS_52468879185703  pfet_CDNS_52468879185703_0
timestamp 1707688321
transform 1 0 119 0 -1 624
box -119 -66 375 266
use pfet_CDNS_52468879185703  pfet_CDNS_52468879185703_1
timestamp 1707688321
transform 1 0 431 0 -1 624
box -119 -66 375 266
<< properties >>
string GDS_END 25724956
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25719460
string path 15.600 12.675 12.350 12.675 
<< end >>
