magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 51673 624 51721
rect 212 51615 268 51624
rect 212 51550 268 51559
rect 0 51453 624 51501
rect 212 51378 268 51387
rect 212 51313 268 51322
rect 0 51199 624 51247
rect 212 51141 268 51150
rect 212 51076 268 51085
rect 0 50979 624 51027
rect 0 50883 624 50931
rect 212 50825 268 50834
rect 212 50760 268 50769
rect 0 50663 624 50711
rect 212 50588 268 50597
rect 212 50523 268 50532
rect 0 50409 624 50457
rect 212 50351 268 50360
rect 212 50286 268 50295
rect 0 50189 624 50237
rect 0 50093 624 50141
rect 212 50035 268 50044
rect 212 49970 268 49979
rect 0 49873 624 49921
rect 212 49798 268 49807
rect 212 49733 268 49742
rect 0 49619 624 49667
rect 212 49561 268 49570
rect 212 49496 268 49505
rect 0 49399 624 49447
rect 0 49303 624 49351
rect 212 49245 268 49254
rect 212 49180 268 49189
rect 0 49083 624 49131
rect 212 49008 268 49017
rect 212 48943 268 48952
rect 0 48829 624 48877
rect 212 48771 268 48780
rect 212 48706 268 48715
rect 0 48609 624 48657
rect 0 48513 624 48561
rect 212 48455 268 48464
rect 212 48390 268 48399
rect 0 48293 624 48341
rect 212 48218 268 48227
rect 212 48153 268 48162
rect 0 48039 624 48087
rect 212 47981 268 47990
rect 212 47916 268 47925
rect 0 47819 624 47867
rect 0 47723 624 47771
rect 212 47665 268 47674
rect 212 47600 268 47609
rect 0 47503 624 47551
rect 212 47428 268 47437
rect 212 47363 268 47372
rect 0 47249 624 47297
rect 212 47191 268 47200
rect 212 47126 268 47135
rect 0 47029 624 47077
rect 0 46933 624 46981
rect 212 46875 268 46884
rect 212 46810 268 46819
rect 0 46713 624 46761
rect 212 46638 268 46647
rect 212 46573 268 46582
rect 0 46459 624 46507
rect 212 46401 268 46410
rect 212 46336 268 46345
rect 0 46239 624 46287
rect 0 46143 624 46191
rect 212 46085 268 46094
rect 212 46020 268 46029
rect 0 45923 624 45971
rect 212 45848 268 45857
rect 212 45783 268 45792
rect 0 45669 624 45717
rect 212 45611 268 45620
rect 212 45546 268 45555
rect 0 45449 624 45497
rect 0 45353 624 45401
rect 212 45295 268 45304
rect 212 45230 268 45239
rect 0 45133 624 45181
rect 212 45058 268 45067
rect 212 44993 268 45002
rect 0 44879 624 44927
rect 212 44821 268 44830
rect 212 44756 268 44765
rect 0 44659 624 44707
rect 0 44563 624 44611
rect 212 44505 268 44514
rect 212 44440 268 44449
rect 0 44343 624 44391
rect 212 44268 268 44277
rect 212 44203 268 44212
rect 0 44089 624 44137
rect 212 44031 268 44040
rect 212 43966 268 43975
rect 0 43869 624 43917
rect 0 43773 624 43821
rect 212 43715 268 43724
rect 212 43650 268 43659
rect 0 43553 624 43601
rect 212 43478 268 43487
rect 212 43413 268 43422
rect 0 43299 624 43347
rect 212 43241 268 43250
rect 212 43176 268 43185
rect 0 43079 624 43127
rect 0 42983 624 43031
rect 212 42925 268 42934
rect 212 42860 268 42869
rect 0 42763 624 42811
rect 212 42688 268 42697
rect 212 42623 268 42632
rect 0 42509 624 42557
rect 212 42451 268 42460
rect 212 42386 268 42395
rect 0 42289 624 42337
rect 0 42193 624 42241
rect 212 42135 268 42144
rect 212 42070 268 42079
rect 0 41973 624 42021
rect 212 41898 268 41907
rect 212 41833 268 41842
rect 0 41719 624 41767
rect 212 41661 268 41670
rect 212 41596 268 41605
rect 0 41499 624 41547
rect 0 41403 624 41451
rect 212 41345 268 41354
rect 212 41280 268 41289
rect 0 41183 624 41231
rect 212 41108 268 41117
rect 212 41043 268 41052
rect 0 40929 624 40977
rect 212 40871 268 40880
rect 212 40806 268 40815
rect 0 40709 624 40757
rect 0 40613 624 40661
rect 212 40555 268 40564
rect 212 40490 268 40499
rect 0 40393 624 40441
rect 212 40318 268 40327
rect 212 40253 268 40262
rect 0 40139 624 40187
rect 212 40081 268 40090
rect 212 40016 268 40025
rect 0 39919 624 39967
rect 0 39823 624 39871
rect 212 39765 268 39774
rect 212 39700 268 39709
rect 0 39603 624 39651
rect 212 39528 268 39537
rect 212 39463 268 39472
rect 0 39349 624 39397
rect 212 39291 268 39300
rect 212 39226 268 39235
rect 0 39129 624 39177
rect 0 39033 624 39081
rect 212 38975 268 38984
rect 212 38910 268 38919
rect 0 38813 624 38861
rect 212 38738 268 38747
rect 212 38673 268 38682
rect 0 38559 624 38607
rect 212 38501 268 38510
rect 212 38436 268 38445
rect 0 38339 624 38387
rect 0 38243 624 38291
rect 212 38185 268 38194
rect 212 38120 268 38129
rect 0 38023 624 38071
rect 212 37948 268 37957
rect 212 37883 268 37892
rect 0 37769 624 37817
rect 212 37711 268 37720
rect 212 37646 268 37655
rect 0 37549 624 37597
rect 0 37453 624 37501
rect 212 37395 268 37404
rect 212 37330 268 37339
rect 0 37233 624 37281
rect 212 37158 268 37167
rect 212 37093 268 37102
rect 0 36979 624 37027
rect 212 36921 268 36930
rect 212 36856 268 36865
rect 0 36759 624 36807
rect 0 36663 624 36711
rect 212 36605 268 36614
rect 212 36540 268 36549
rect 0 36443 624 36491
rect 212 36368 268 36377
rect 212 36303 268 36312
rect 0 36189 624 36237
rect 212 36131 268 36140
rect 212 36066 268 36075
rect 0 35969 624 36017
rect 0 35873 624 35921
rect 212 35815 268 35824
rect 212 35750 268 35759
rect 0 35653 624 35701
rect 212 35578 268 35587
rect 212 35513 268 35522
rect 0 35399 624 35447
rect 212 35341 268 35350
rect 212 35276 268 35285
rect 0 35179 624 35227
rect 0 35083 624 35131
rect 212 35025 268 35034
rect 212 34960 268 34969
rect 0 34863 624 34911
rect 212 34788 268 34797
rect 212 34723 268 34732
rect 0 34609 624 34657
rect 212 34551 268 34560
rect 212 34486 268 34495
rect 0 34389 624 34437
rect 0 34293 624 34341
rect 212 34235 268 34244
rect 212 34170 268 34179
rect 0 34073 624 34121
rect 212 33998 268 34007
rect 212 33933 268 33942
rect 0 33819 624 33867
rect 212 33761 268 33770
rect 212 33696 268 33705
rect 0 33599 624 33647
rect 0 33503 624 33551
rect 212 33445 268 33454
rect 212 33380 268 33389
rect 0 33283 624 33331
rect 212 33208 268 33217
rect 212 33143 268 33152
rect 0 33029 624 33077
rect 212 32971 268 32980
rect 212 32906 268 32915
rect 0 32809 624 32857
rect 0 32713 624 32761
rect 212 32655 268 32664
rect 212 32590 268 32599
rect 0 32493 624 32541
rect 212 32418 268 32427
rect 212 32353 268 32362
rect 0 32239 624 32287
rect 212 32181 268 32190
rect 212 32116 268 32125
rect 0 32019 624 32067
rect 0 31923 624 31971
rect 212 31865 268 31874
rect 212 31800 268 31809
rect 0 31703 624 31751
rect 212 31628 268 31637
rect 212 31563 268 31572
rect 0 31449 624 31497
rect 212 31391 268 31400
rect 212 31326 268 31335
rect 0 31229 624 31277
rect 0 31133 624 31181
rect 212 31075 268 31084
rect 212 31010 268 31019
rect 0 30913 624 30961
rect 212 30838 268 30847
rect 212 30773 268 30782
rect 0 30659 624 30707
rect 212 30601 268 30610
rect 212 30536 268 30545
rect 0 30439 624 30487
rect 0 30343 624 30391
rect 212 30285 268 30294
rect 212 30220 268 30229
rect 0 30123 624 30171
rect 212 30048 268 30057
rect 212 29983 268 29992
rect 0 29869 624 29917
rect 212 29811 268 29820
rect 212 29746 268 29755
rect 0 29649 624 29697
rect 0 29553 624 29601
rect 212 29495 268 29504
rect 212 29430 268 29439
rect 0 29333 624 29381
rect 212 29258 268 29267
rect 212 29193 268 29202
rect 0 29079 624 29127
rect 212 29021 268 29030
rect 212 28956 268 28965
rect 0 28859 624 28907
rect 0 28763 624 28811
rect 212 28705 268 28714
rect 212 28640 268 28649
rect 0 28543 624 28591
rect 212 28468 268 28477
rect 212 28403 268 28412
rect 0 28289 624 28337
rect 212 28231 268 28240
rect 212 28166 268 28175
rect 0 28069 624 28117
rect 0 27973 624 28021
rect 212 27915 268 27924
rect 212 27850 268 27859
rect 0 27753 624 27801
rect 212 27678 268 27687
rect 212 27613 268 27622
rect 0 27499 624 27547
rect 212 27441 268 27450
rect 212 27376 268 27385
rect 0 27279 624 27327
rect 0 27183 624 27231
rect 212 27125 268 27134
rect 212 27060 268 27069
rect 0 26963 624 27011
rect 212 26888 268 26897
rect 212 26823 268 26832
rect 0 26709 624 26757
rect 212 26651 268 26660
rect 212 26586 268 26595
rect 0 26489 624 26537
rect 0 26393 624 26441
rect 212 26335 268 26344
rect 212 26270 268 26279
rect 0 26173 624 26221
rect 212 26098 268 26107
rect 212 26033 268 26042
rect 0 25919 624 25967
rect 212 25861 268 25870
rect 212 25796 268 25805
rect 0 25699 624 25747
rect 0 25603 624 25651
rect 212 25545 268 25554
rect 212 25480 268 25489
rect 0 25383 624 25431
rect 212 25308 268 25317
rect 212 25243 268 25252
rect 0 25129 624 25177
rect 212 25071 268 25080
rect 212 25006 268 25015
rect 0 24909 624 24957
rect 0 24813 624 24861
rect 212 24755 268 24764
rect 212 24690 268 24699
rect 0 24593 624 24641
rect 212 24518 268 24527
rect 212 24453 268 24462
rect 0 24339 624 24387
rect 212 24281 268 24290
rect 212 24216 268 24225
rect 0 24119 624 24167
rect 0 24023 624 24071
rect 212 23965 268 23974
rect 212 23900 268 23909
rect 0 23803 624 23851
rect 212 23728 268 23737
rect 212 23663 268 23672
rect 0 23549 624 23597
rect 212 23491 268 23500
rect 212 23426 268 23435
rect 0 23329 624 23377
rect 0 23233 624 23281
rect 212 23175 268 23184
rect 212 23110 268 23119
rect 0 23013 624 23061
rect 212 22938 268 22947
rect 212 22873 268 22882
rect 0 22759 624 22807
rect 212 22701 268 22710
rect 212 22636 268 22645
rect 0 22539 624 22587
rect 0 22443 624 22491
rect 212 22385 268 22394
rect 212 22320 268 22329
rect 0 22223 624 22271
rect 212 22148 268 22157
rect 212 22083 268 22092
rect 0 21969 624 22017
rect 212 21911 268 21920
rect 212 21846 268 21855
rect 0 21749 624 21797
rect 0 21653 624 21701
rect 212 21595 268 21604
rect 212 21530 268 21539
rect 0 21433 624 21481
rect 212 21358 268 21367
rect 212 21293 268 21302
rect 0 21179 624 21227
rect 212 21121 268 21130
rect 212 21056 268 21065
rect 0 20959 624 21007
rect 0 20863 624 20911
rect 212 20805 268 20814
rect 212 20740 268 20749
rect 0 20643 624 20691
rect 212 20568 268 20577
rect 212 20503 268 20512
rect 0 20389 624 20437
rect 212 20331 268 20340
rect 212 20266 268 20275
rect 0 20169 624 20217
rect 0 20073 624 20121
rect 212 20015 268 20024
rect 212 19950 268 19959
rect 0 19853 624 19901
rect 212 19778 268 19787
rect 212 19713 268 19722
rect 0 19599 624 19647
rect 212 19541 268 19550
rect 212 19476 268 19485
rect 0 19379 624 19427
rect 0 19283 624 19331
rect 212 19225 268 19234
rect 212 19160 268 19169
rect 0 19063 624 19111
rect 212 18988 268 18997
rect 212 18923 268 18932
rect 0 18809 624 18857
rect 212 18751 268 18760
rect 212 18686 268 18695
rect 0 18589 624 18637
rect 0 18493 624 18541
rect 212 18435 268 18444
rect 212 18370 268 18379
rect 0 18273 624 18321
rect 212 18198 268 18207
rect 212 18133 268 18142
rect 0 18019 624 18067
rect 212 17961 268 17970
rect 212 17896 268 17905
rect 0 17799 624 17847
rect 0 17703 624 17751
rect 212 17645 268 17654
rect 212 17580 268 17589
rect 0 17483 624 17531
rect 212 17408 268 17417
rect 212 17343 268 17352
rect 0 17229 624 17277
rect 212 17171 268 17180
rect 212 17106 268 17115
rect 0 17009 624 17057
rect 0 16913 624 16961
rect 212 16855 268 16864
rect 212 16790 268 16799
rect 0 16693 624 16741
rect 212 16618 268 16627
rect 212 16553 268 16562
rect 0 16439 624 16487
rect 212 16381 268 16390
rect 212 16316 268 16325
rect 0 16219 624 16267
rect 0 16123 624 16171
rect 212 16065 268 16074
rect 212 16000 268 16009
rect 0 15903 624 15951
rect 212 15828 268 15837
rect 212 15763 268 15772
rect 0 15649 624 15697
rect 212 15591 268 15600
rect 212 15526 268 15535
rect 0 15429 624 15477
rect 0 15333 624 15381
rect 212 15275 268 15284
rect 212 15210 268 15219
rect 0 15113 624 15161
rect 212 15038 268 15047
rect 212 14973 268 14982
rect 0 14859 624 14907
rect 212 14801 268 14810
rect 212 14736 268 14745
rect 0 14639 624 14687
rect 0 14543 624 14591
rect 212 14485 268 14494
rect 212 14420 268 14429
rect 0 14323 624 14371
rect 212 14248 268 14257
rect 212 14183 268 14192
rect 0 14069 624 14117
rect 212 14011 268 14020
rect 212 13946 268 13955
rect 0 13849 624 13897
rect 0 13753 624 13801
rect 212 13695 268 13704
rect 212 13630 268 13639
rect 0 13533 624 13581
rect 212 13458 268 13467
rect 212 13393 268 13402
rect 0 13279 624 13327
rect 212 13221 268 13230
rect 212 13156 268 13165
rect 0 13059 624 13107
rect 0 12963 624 13011
rect 212 12905 268 12914
rect 212 12840 268 12849
rect 0 12743 624 12791
rect 212 12668 268 12677
rect 212 12603 268 12612
rect 0 12489 624 12537
rect 212 12431 268 12440
rect 212 12366 268 12375
rect 0 12269 624 12317
rect 0 12173 624 12221
rect 212 12115 268 12124
rect 212 12050 268 12059
rect 0 11953 624 12001
rect 212 11878 268 11887
rect 212 11813 268 11822
rect 0 11699 624 11747
rect 212 11641 268 11650
rect 212 11576 268 11585
rect 0 11479 624 11527
rect 0 11383 624 11431
rect 212 11325 268 11334
rect 212 11260 268 11269
rect 0 11163 624 11211
rect 212 11088 268 11097
rect 212 11023 268 11032
rect 0 10909 624 10957
rect 212 10851 268 10860
rect 212 10786 268 10795
rect 0 10689 624 10737
rect 0 10593 624 10641
rect 212 10535 268 10544
rect 212 10470 268 10479
rect 0 10373 624 10421
rect 212 10298 268 10307
rect 212 10233 268 10242
rect 0 10119 624 10167
rect 212 10061 268 10070
rect 212 9996 268 10005
rect 0 9899 624 9947
rect 0 9803 624 9851
rect 212 9745 268 9754
rect 212 9680 268 9689
rect 0 9583 624 9631
rect 212 9508 268 9517
rect 212 9443 268 9452
rect 0 9329 624 9377
rect 212 9271 268 9280
rect 212 9206 268 9215
rect 0 9109 624 9157
rect 0 9013 624 9061
rect 212 8955 268 8964
rect 212 8890 268 8899
rect 0 8793 624 8841
rect 212 8718 268 8727
rect 212 8653 268 8662
rect 0 8539 624 8587
rect 212 8481 268 8490
rect 212 8416 268 8425
rect 0 8319 624 8367
rect 0 8223 624 8271
rect 212 8165 268 8174
rect 212 8100 268 8109
rect 0 8003 624 8051
rect 212 7928 268 7937
rect 212 7863 268 7872
rect 0 7749 624 7797
rect 212 7691 268 7700
rect 212 7626 268 7635
rect 0 7529 624 7577
rect 0 7433 624 7481
rect 212 7375 268 7384
rect 212 7310 268 7319
rect 0 7213 624 7261
rect 212 7138 268 7147
rect 212 7073 268 7082
rect 0 6959 624 7007
rect 212 6901 268 6910
rect 212 6836 268 6845
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 212 6585 268 6594
rect 212 6520 268 6529
rect 0 6423 624 6471
rect 212 6348 268 6357
rect 212 6283 268 6292
rect 0 6169 624 6217
rect 212 6111 268 6120
rect 212 6046 268 6055
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 212 5795 268 5804
rect 212 5730 268 5739
rect 0 5633 624 5681
rect 212 5558 268 5567
rect 212 5493 268 5502
rect 0 5379 624 5427
rect 212 5321 268 5330
rect 212 5256 268 5265
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 212 5005 268 5014
rect 212 4940 268 4949
rect 0 4843 624 4891
rect 212 4768 268 4777
rect 212 4703 268 4712
rect 0 4589 624 4637
rect 212 4531 268 4540
rect 212 4466 268 4475
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 212 4215 268 4224
rect 212 4150 268 4159
rect 0 4053 624 4101
rect 212 3978 268 3987
rect 212 3913 268 3922
rect 0 3799 624 3847
rect 212 3741 268 3750
rect 212 3676 268 3685
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 212 3425 268 3434
rect 212 3360 268 3369
rect 0 3263 624 3311
rect 212 3188 268 3197
rect 212 3123 268 3132
rect 0 3009 624 3057
rect 212 2951 268 2960
rect 212 2886 268 2895
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 212 2635 268 2644
rect 212 2570 268 2579
rect 0 2473 624 2521
rect 212 2398 268 2407
rect 212 2333 268 2342
rect 0 2219 624 2267
rect 212 2161 268 2170
rect 212 2096 268 2105
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 212 1845 268 1854
rect 212 1780 268 1789
rect 0 1683 624 1731
rect 212 1608 268 1617
rect 212 1543 268 1552
rect 0 1429 624 1477
rect 212 1371 268 1380
rect 212 1306 268 1315
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 212 1055 268 1064
rect 212 990 268 999
rect 0 893 624 941
rect 212 818 268 827
rect 212 753 268 762
rect 0 639 624 687
rect 212 581 268 590
rect 212 516 268 525
rect 0 419 624 467
<< via2 >>
rect 212 51559 268 51615
rect 212 51322 268 51378
rect 212 51085 268 51141
rect 212 50769 268 50825
rect 212 50532 268 50588
rect 212 50295 268 50351
rect 212 49979 268 50035
rect 212 49742 268 49798
rect 212 49505 268 49561
rect 212 49189 268 49245
rect 212 48952 268 49008
rect 212 48715 268 48771
rect 212 48399 268 48455
rect 212 48162 268 48218
rect 212 47925 268 47981
rect 212 47609 268 47665
rect 212 47372 268 47428
rect 212 47135 268 47191
rect 212 46819 268 46875
rect 212 46582 268 46638
rect 212 46345 268 46401
rect 212 46029 268 46085
rect 212 45792 268 45848
rect 212 45555 268 45611
rect 212 45239 268 45295
rect 212 45002 268 45058
rect 212 44765 268 44821
rect 212 44449 268 44505
rect 212 44212 268 44268
rect 212 43975 268 44031
rect 212 43659 268 43715
rect 212 43422 268 43478
rect 212 43185 268 43241
rect 212 42869 268 42925
rect 212 42632 268 42688
rect 212 42395 268 42451
rect 212 42079 268 42135
rect 212 41842 268 41898
rect 212 41605 268 41661
rect 212 41289 268 41345
rect 212 41052 268 41108
rect 212 40815 268 40871
rect 212 40499 268 40555
rect 212 40262 268 40318
rect 212 40025 268 40081
rect 212 39709 268 39765
rect 212 39472 268 39528
rect 212 39235 268 39291
rect 212 38919 268 38975
rect 212 38682 268 38738
rect 212 38445 268 38501
rect 212 38129 268 38185
rect 212 37892 268 37948
rect 212 37655 268 37711
rect 212 37339 268 37395
rect 212 37102 268 37158
rect 212 36865 268 36921
rect 212 36549 268 36605
rect 212 36312 268 36368
rect 212 36075 268 36131
rect 212 35759 268 35815
rect 212 35522 268 35578
rect 212 35285 268 35341
rect 212 34969 268 35025
rect 212 34732 268 34788
rect 212 34495 268 34551
rect 212 34179 268 34235
rect 212 33942 268 33998
rect 212 33705 268 33761
rect 212 33389 268 33445
rect 212 33152 268 33208
rect 212 32915 268 32971
rect 212 32599 268 32655
rect 212 32362 268 32418
rect 212 32125 268 32181
rect 212 31809 268 31865
rect 212 31572 268 31628
rect 212 31335 268 31391
rect 212 31019 268 31075
rect 212 30782 268 30838
rect 212 30545 268 30601
rect 212 30229 268 30285
rect 212 29992 268 30048
rect 212 29755 268 29811
rect 212 29439 268 29495
rect 212 29202 268 29258
rect 212 28965 268 29021
rect 212 28649 268 28705
rect 212 28412 268 28468
rect 212 28175 268 28231
rect 212 27859 268 27915
rect 212 27622 268 27678
rect 212 27385 268 27441
rect 212 27069 268 27125
rect 212 26832 268 26888
rect 212 26595 268 26651
rect 212 26279 268 26335
rect 212 26042 268 26098
rect 212 25805 268 25861
rect 212 25489 268 25545
rect 212 25252 268 25308
rect 212 25015 268 25071
rect 212 24699 268 24755
rect 212 24462 268 24518
rect 212 24225 268 24281
rect 212 23909 268 23965
rect 212 23672 268 23728
rect 212 23435 268 23491
rect 212 23119 268 23175
rect 212 22882 268 22938
rect 212 22645 268 22701
rect 212 22329 268 22385
rect 212 22092 268 22148
rect 212 21855 268 21911
rect 212 21539 268 21595
rect 212 21302 268 21358
rect 212 21065 268 21121
rect 212 20749 268 20805
rect 212 20512 268 20568
rect 212 20275 268 20331
rect 212 19959 268 20015
rect 212 19722 268 19778
rect 212 19485 268 19541
rect 212 19169 268 19225
rect 212 18932 268 18988
rect 212 18695 268 18751
rect 212 18379 268 18435
rect 212 18142 268 18198
rect 212 17905 268 17961
rect 212 17589 268 17645
rect 212 17352 268 17408
rect 212 17115 268 17171
rect 212 16799 268 16855
rect 212 16562 268 16618
rect 212 16325 268 16381
rect 212 16009 268 16065
rect 212 15772 268 15828
rect 212 15535 268 15591
rect 212 15219 268 15275
rect 212 14982 268 15038
rect 212 14745 268 14801
rect 212 14429 268 14485
rect 212 14192 268 14248
rect 212 13955 268 14011
rect 212 13639 268 13695
rect 212 13402 268 13458
rect 212 13165 268 13221
rect 212 12849 268 12905
rect 212 12612 268 12668
rect 212 12375 268 12431
rect 212 12059 268 12115
rect 212 11822 268 11878
rect 212 11585 268 11641
rect 212 11269 268 11325
rect 212 11032 268 11088
rect 212 10795 268 10851
rect 212 10479 268 10535
rect 212 10242 268 10298
rect 212 10005 268 10061
rect 212 9689 268 9745
rect 212 9452 268 9508
rect 212 9215 268 9271
rect 212 8899 268 8955
rect 212 8662 268 8718
rect 212 8425 268 8481
rect 212 8109 268 8165
rect 212 7872 268 7928
rect 212 7635 268 7691
rect 212 7319 268 7375
rect 212 7082 268 7138
rect 212 6845 268 6901
rect 212 6529 268 6585
rect 212 6292 268 6348
rect 212 6055 268 6111
rect 212 5739 268 5795
rect 212 5502 268 5558
rect 212 5265 268 5321
rect 212 4949 268 5005
rect 212 4712 268 4768
rect 212 4475 268 4531
rect 212 4159 268 4215
rect 212 3922 268 3978
rect 212 3685 268 3741
rect 212 3369 268 3425
rect 212 3132 268 3188
rect 212 2895 268 2951
rect 212 2579 268 2635
rect 212 2342 268 2398
rect 212 2105 268 2161
rect 212 1789 268 1845
rect 212 1552 268 1608
rect 212 1315 268 1371
rect 212 999 268 1055
rect 212 762 268 818
rect 212 525 268 581
<< metal3 >>
rect 191 51615 289 51636
rect 191 51559 212 51615
rect 268 51559 289 51615
rect 191 51538 289 51559
rect 191 51378 289 51399
rect 191 51322 212 51378
rect 268 51322 289 51378
rect 191 51301 289 51322
rect 191 51141 289 51162
rect 191 51085 212 51141
rect 268 51085 289 51141
rect 191 51064 289 51085
rect 191 50825 289 50846
rect 191 50769 212 50825
rect 268 50769 289 50825
rect 191 50748 289 50769
rect 191 50588 289 50609
rect 191 50532 212 50588
rect 268 50532 289 50588
rect 191 50511 289 50532
rect 191 50351 289 50372
rect 191 50295 212 50351
rect 268 50295 289 50351
rect 191 50274 289 50295
rect 191 50035 289 50056
rect 191 49979 212 50035
rect 268 49979 289 50035
rect 191 49958 289 49979
rect 191 49798 289 49819
rect 191 49742 212 49798
rect 268 49742 289 49798
rect 191 49721 289 49742
rect 191 49561 289 49582
rect 191 49505 212 49561
rect 268 49505 289 49561
rect 191 49484 289 49505
rect 191 49245 289 49266
rect 191 49189 212 49245
rect 268 49189 289 49245
rect 191 49168 289 49189
rect 191 49008 289 49029
rect 191 48952 212 49008
rect 268 48952 289 49008
rect 191 48931 289 48952
rect 191 48771 289 48792
rect 191 48715 212 48771
rect 268 48715 289 48771
rect 191 48694 289 48715
rect 191 48455 289 48476
rect 191 48399 212 48455
rect 268 48399 289 48455
rect 191 48378 289 48399
rect 191 48218 289 48239
rect 191 48162 212 48218
rect 268 48162 289 48218
rect 191 48141 289 48162
rect 191 47981 289 48002
rect 191 47925 212 47981
rect 268 47925 289 47981
rect 191 47904 289 47925
rect 191 47665 289 47686
rect 191 47609 212 47665
rect 268 47609 289 47665
rect 191 47588 289 47609
rect 191 47428 289 47449
rect 191 47372 212 47428
rect 268 47372 289 47428
rect 191 47351 289 47372
rect 191 47191 289 47212
rect 191 47135 212 47191
rect 268 47135 289 47191
rect 191 47114 289 47135
rect 191 46875 289 46896
rect 191 46819 212 46875
rect 268 46819 289 46875
rect 191 46798 289 46819
rect 191 46638 289 46659
rect 191 46582 212 46638
rect 268 46582 289 46638
rect 191 46561 289 46582
rect 191 46401 289 46422
rect 191 46345 212 46401
rect 268 46345 289 46401
rect 191 46324 289 46345
rect 191 46085 289 46106
rect 191 46029 212 46085
rect 268 46029 289 46085
rect 191 46008 289 46029
rect 191 45848 289 45869
rect 191 45792 212 45848
rect 268 45792 289 45848
rect 191 45771 289 45792
rect 191 45611 289 45632
rect 191 45555 212 45611
rect 268 45555 289 45611
rect 191 45534 289 45555
rect 191 45295 289 45316
rect 191 45239 212 45295
rect 268 45239 289 45295
rect 191 45218 289 45239
rect 191 45058 289 45079
rect 191 45002 212 45058
rect 268 45002 289 45058
rect 191 44981 289 45002
rect 191 44821 289 44842
rect 191 44765 212 44821
rect 268 44765 289 44821
rect 191 44744 289 44765
rect 191 44505 289 44526
rect 191 44449 212 44505
rect 268 44449 289 44505
rect 191 44428 289 44449
rect 191 44268 289 44289
rect 191 44212 212 44268
rect 268 44212 289 44268
rect 191 44191 289 44212
rect 191 44031 289 44052
rect 191 43975 212 44031
rect 268 43975 289 44031
rect 191 43954 289 43975
rect 191 43715 289 43736
rect 191 43659 212 43715
rect 268 43659 289 43715
rect 191 43638 289 43659
rect 191 43478 289 43499
rect 191 43422 212 43478
rect 268 43422 289 43478
rect 191 43401 289 43422
rect 191 43241 289 43262
rect 191 43185 212 43241
rect 268 43185 289 43241
rect 191 43164 289 43185
rect 191 42925 289 42946
rect 191 42869 212 42925
rect 268 42869 289 42925
rect 191 42848 289 42869
rect 191 42688 289 42709
rect 191 42632 212 42688
rect 268 42632 289 42688
rect 191 42611 289 42632
rect 191 42451 289 42472
rect 191 42395 212 42451
rect 268 42395 289 42451
rect 191 42374 289 42395
rect 191 42135 289 42156
rect 191 42079 212 42135
rect 268 42079 289 42135
rect 191 42058 289 42079
rect 191 41898 289 41919
rect 191 41842 212 41898
rect 268 41842 289 41898
rect 191 41821 289 41842
rect 191 41661 289 41682
rect 191 41605 212 41661
rect 268 41605 289 41661
rect 191 41584 289 41605
rect 191 41345 289 41366
rect 191 41289 212 41345
rect 268 41289 289 41345
rect 191 41268 289 41289
rect 191 41108 289 41129
rect 191 41052 212 41108
rect 268 41052 289 41108
rect 191 41031 289 41052
rect 191 40871 289 40892
rect 191 40815 212 40871
rect 268 40815 289 40871
rect 191 40794 289 40815
rect 191 40555 289 40576
rect 191 40499 212 40555
rect 268 40499 289 40555
rect 191 40478 289 40499
rect 191 40318 289 40339
rect 191 40262 212 40318
rect 268 40262 289 40318
rect 191 40241 289 40262
rect 191 40081 289 40102
rect 191 40025 212 40081
rect 268 40025 289 40081
rect 191 40004 289 40025
rect 191 39765 289 39786
rect 191 39709 212 39765
rect 268 39709 289 39765
rect 191 39688 289 39709
rect 191 39528 289 39549
rect 191 39472 212 39528
rect 268 39472 289 39528
rect 191 39451 289 39472
rect 191 39291 289 39312
rect 191 39235 212 39291
rect 268 39235 289 39291
rect 191 39214 289 39235
rect 191 38975 289 38996
rect 191 38919 212 38975
rect 268 38919 289 38975
rect 191 38898 289 38919
rect 191 38738 289 38759
rect 191 38682 212 38738
rect 268 38682 289 38738
rect 191 38661 289 38682
rect 191 38501 289 38522
rect 191 38445 212 38501
rect 268 38445 289 38501
rect 191 38424 289 38445
rect 191 38185 289 38206
rect 191 38129 212 38185
rect 268 38129 289 38185
rect 191 38108 289 38129
rect 191 37948 289 37969
rect 191 37892 212 37948
rect 268 37892 289 37948
rect 191 37871 289 37892
rect 191 37711 289 37732
rect 191 37655 212 37711
rect 268 37655 289 37711
rect 191 37634 289 37655
rect 191 37395 289 37416
rect 191 37339 212 37395
rect 268 37339 289 37395
rect 191 37318 289 37339
rect 191 37158 289 37179
rect 191 37102 212 37158
rect 268 37102 289 37158
rect 191 37081 289 37102
rect 191 36921 289 36942
rect 191 36865 212 36921
rect 268 36865 289 36921
rect 191 36844 289 36865
rect 191 36605 289 36626
rect 191 36549 212 36605
rect 268 36549 289 36605
rect 191 36528 289 36549
rect 191 36368 289 36389
rect 191 36312 212 36368
rect 268 36312 289 36368
rect 191 36291 289 36312
rect 191 36131 289 36152
rect 191 36075 212 36131
rect 268 36075 289 36131
rect 191 36054 289 36075
rect 191 35815 289 35836
rect 191 35759 212 35815
rect 268 35759 289 35815
rect 191 35738 289 35759
rect 191 35578 289 35599
rect 191 35522 212 35578
rect 268 35522 289 35578
rect 191 35501 289 35522
rect 191 35341 289 35362
rect 191 35285 212 35341
rect 268 35285 289 35341
rect 191 35264 289 35285
rect 191 35025 289 35046
rect 191 34969 212 35025
rect 268 34969 289 35025
rect 191 34948 289 34969
rect 191 34788 289 34809
rect 191 34732 212 34788
rect 268 34732 289 34788
rect 191 34711 289 34732
rect 191 34551 289 34572
rect 191 34495 212 34551
rect 268 34495 289 34551
rect 191 34474 289 34495
rect 191 34235 289 34256
rect 191 34179 212 34235
rect 268 34179 289 34235
rect 191 34158 289 34179
rect 191 33998 289 34019
rect 191 33942 212 33998
rect 268 33942 289 33998
rect 191 33921 289 33942
rect 191 33761 289 33782
rect 191 33705 212 33761
rect 268 33705 289 33761
rect 191 33684 289 33705
rect 191 33445 289 33466
rect 191 33389 212 33445
rect 268 33389 289 33445
rect 191 33368 289 33389
rect 191 33208 289 33229
rect 191 33152 212 33208
rect 268 33152 289 33208
rect 191 33131 289 33152
rect 191 32971 289 32992
rect 191 32915 212 32971
rect 268 32915 289 32971
rect 191 32894 289 32915
rect 191 32655 289 32676
rect 191 32599 212 32655
rect 268 32599 289 32655
rect 191 32578 289 32599
rect 191 32418 289 32439
rect 191 32362 212 32418
rect 268 32362 289 32418
rect 191 32341 289 32362
rect 191 32181 289 32202
rect 191 32125 212 32181
rect 268 32125 289 32181
rect 191 32104 289 32125
rect 191 31865 289 31886
rect 191 31809 212 31865
rect 268 31809 289 31865
rect 191 31788 289 31809
rect 191 31628 289 31649
rect 191 31572 212 31628
rect 268 31572 289 31628
rect 191 31551 289 31572
rect 191 31391 289 31412
rect 191 31335 212 31391
rect 268 31335 289 31391
rect 191 31314 289 31335
rect 191 31075 289 31096
rect 191 31019 212 31075
rect 268 31019 289 31075
rect 191 30998 289 31019
rect 191 30838 289 30859
rect 191 30782 212 30838
rect 268 30782 289 30838
rect 191 30761 289 30782
rect 191 30601 289 30622
rect 191 30545 212 30601
rect 268 30545 289 30601
rect 191 30524 289 30545
rect 191 30285 289 30306
rect 191 30229 212 30285
rect 268 30229 289 30285
rect 191 30208 289 30229
rect 191 30048 289 30069
rect 191 29992 212 30048
rect 268 29992 289 30048
rect 191 29971 289 29992
rect 191 29811 289 29832
rect 191 29755 212 29811
rect 268 29755 289 29811
rect 191 29734 289 29755
rect 191 29495 289 29516
rect 191 29439 212 29495
rect 268 29439 289 29495
rect 191 29418 289 29439
rect 191 29258 289 29279
rect 191 29202 212 29258
rect 268 29202 289 29258
rect 191 29181 289 29202
rect 191 29021 289 29042
rect 191 28965 212 29021
rect 268 28965 289 29021
rect 191 28944 289 28965
rect 191 28705 289 28726
rect 191 28649 212 28705
rect 268 28649 289 28705
rect 191 28628 289 28649
rect 191 28468 289 28489
rect 191 28412 212 28468
rect 268 28412 289 28468
rect 191 28391 289 28412
rect 191 28231 289 28252
rect 191 28175 212 28231
rect 268 28175 289 28231
rect 191 28154 289 28175
rect 191 27915 289 27936
rect 191 27859 212 27915
rect 268 27859 289 27915
rect 191 27838 289 27859
rect 191 27678 289 27699
rect 191 27622 212 27678
rect 268 27622 289 27678
rect 191 27601 289 27622
rect 191 27441 289 27462
rect 191 27385 212 27441
rect 268 27385 289 27441
rect 191 27364 289 27385
rect 191 27125 289 27146
rect 191 27069 212 27125
rect 268 27069 289 27125
rect 191 27048 289 27069
rect 191 26888 289 26909
rect 191 26832 212 26888
rect 268 26832 289 26888
rect 191 26811 289 26832
rect 191 26651 289 26672
rect 191 26595 212 26651
rect 268 26595 289 26651
rect 191 26574 289 26595
rect 191 26335 289 26356
rect 191 26279 212 26335
rect 268 26279 289 26335
rect 191 26258 289 26279
rect 191 26098 289 26119
rect 191 26042 212 26098
rect 268 26042 289 26098
rect 191 26021 289 26042
rect 191 25861 289 25882
rect 191 25805 212 25861
rect 268 25805 289 25861
rect 191 25784 289 25805
rect 191 25545 289 25566
rect 191 25489 212 25545
rect 268 25489 289 25545
rect 191 25468 289 25489
rect 191 25308 289 25329
rect 191 25252 212 25308
rect 268 25252 289 25308
rect 191 25231 289 25252
rect 191 25071 289 25092
rect 191 25015 212 25071
rect 268 25015 289 25071
rect 191 24994 289 25015
rect 191 24755 289 24776
rect 191 24699 212 24755
rect 268 24699 289 24755
rect 191 24678 289 24699
rect 191 24518 289 24539
rect 191 24462 212 24518
rect 268 24462 289 24518
rect 191 24441 289 24462
rect 191 24281 289 24302
rect 191 24225 212 24281
rect 268 24225 289 24281
rect 191 24204 289 24225
rect 191 23965 289 23986
rect 191 23909 212 23965
rect 268 23909 289 23965
rect 191 23888 289 23909
rect 191 23728 289 23749
rect 191 23672 212 23728
rect 268 23672 289 23728
rect 191 23651 289 23672
rect 191 23491 289 23512
rect 191 23435 212 23491
rect 268 23435 289 23491
rect 191 23414 289 23435
rect 191 23175 289 23196
rect 191 23119 212 23175
rect 268 23119 289 23175
rect 191 23098 289 23119
rect 191 22938 289 22959
rect 191 22882 212 22938
rect 268 22882 289 22938
rect 191 22861 289 22882
rect 191 22701 289 22722
rect 191 22645 212 22701
rect 268 22645 289 22701
rect 191 22624 289 22645
rect 191 22385 289 22406
rect 191 22329 212 22385
rect 268 22329 289 22385
rect 191 22308 289 22329
rect 191 22148 289 22169
rect 191 22092 212 22148
rect 268 22092 289 22148
rect 191 22071 289 22092
rect 191 21911 289 21932
rect 191 21855 212 21911
rect 268 21855 289 21911
rect 191 21834 289 21855
rect 191 21595 289 21616
rect 191 21539 212 21595
rect 268 21539 289 21595
rect 191 21518 289 21539
rect 191 21358 289 21379
rect 191 21302 212 21358
rect 268 21302 289 21358
rect 191 21281 289 21302
rect 191 21121 289 21142
rect 191 21065 212 21121
rect 268 21065 289 21121
rect 191 21044 289 21065
rect 191 20805 289 20826
rect 191 20749 212 20805
rect 268 20749 289 20805
rect 191 20728 289 20749
rect 191 20568 289 20589
rect 191 20512 212 20568
rect 268 20512 289 20568
rect 191 20491 289 20512
rect 191 20331 289 20352
rect 191 20275 212 20331
rect 268 20275 289 20331
rect 191 20254 289 20275
rect 191 20015 289 20036
rect 191 19959 212 20015
rect 268 19959 289 20015
rect 191 19938 289 19959
rect 191 19778 289 19799
rect 191 19722 212 19778
rect 268 19722 289 19778
rect 191 19701 289 19722
rect 191 19541 289 19562
rect 191 19485 212 19541
rect 268 19485 289 19541
rect 191 19464 289 19485
rect 191 19225 289 19246
rect 191 19169 212 19225
rect 268 19169 289 19225
rect 191 19148 289 19169
rect 191 18988 289 19009
rect 191 18932 212 18988
rect 268 18932 289 18988
rect 191 18911 289 18932
rect 191 18751 289 18772
rect 191 18695 212 18751
rect 268 18695 289 18751
rect 191 18674 289 18695
rect 191 18435 289 18456
rect 191 18379 212 18435
rect 268 18379 289 18435
rect 191 18358 289 18379
rect 191 18198 289 18219
rect 191 18142 212 18198
rect 268 18142 289 18198
rect 191 18121 289 18142
rect 191 17961 289 17982
rect 191 17905 212 17961
rect 268 17905 289 17961
rect 191 17884 289 17905
rect 191 17645 289 17666
rect 191 17589 212 17645
rect 268 17589 289 17645
rect 191 17568 289 17589
rect 191 17408 289 17429
rect 191 17352 212 17408
rect 268 17352 289 17408
rect 191 17331 289 17352
rect 191 17171 289 17192
rect 191 17115 212 17171
rect 268 17115 289 17171
rect 191 17094 289 17115
rect 191 16855 289 16876
rect 191 16799 212 16855
rect 268 16799 289 16855
rect 191 16778 289 16799
rect 191 16618 289 16639
rect 191 16562 212 16618
rect 268 16562 289 16618
rect 191 16541 289 16562
rect 191 16381 289 16402
rect 191 16325 212 16381
rect 268 16325 289 16381
rect 191 16304 289 16325
rect 191 16065 289 16086
rect 191 16009 212 16065
rect 268 16009 289 16065
rect 191 15988 289 16009
rect 191 15828 289 15849
rect 191 15772 212 15828
rect 268 15772 289 15828
rect 191 15751 289 15772
rect 191 15591 289 15612
rect 191 15535 212 15591
rect 268 15535 289 15591
rect 191 15514 289 15535
rect 191 15275 289 15296
rect 191 15219 212 15275
rect 268 15219 289 15275
rect 191 15198 289 15219
rect 191 15038 289 15059
rect 191 14982 212 15038
rect 268 14982 289 15038
rect 191 14961 289 14982
rect 191 14801 289 14822
rect 191 14745 212 14801
rect 268 14745 289 14801
rect 191 14724 289 14745
rect 191 14485 289 14506
rect 191 14429 212 14485
rect 268 14429 289 14485
rect 191 14408 289 14429
rect 191 14248 289 14269
rect 191 14192 212 14248
rect 268 14192 289 14248
rect 191 14171 289 14192
rect 191 14011 289 14032
rect 191 13955 212 14011
rect 268 13955 289 14011
rect 191 13934 289 13955
rect 191 13695 289 13716
rect 191 13639 212 13695
rect 268 13639 289 13695
rect 191 13618 289 13639
rect 191 13458 289 13479
rect 191 13402 212 13458
rect 268 13402 289 13458
rect 191 13381 289 13402
rect 191 13221 289 13242
rect 191 13165 212 13221
rect 268 13165 289 13221
rect 191 13144 289 13165
rect 191 12905 289 12926
rect 191 12849 212 12905
rect 268 12849 289 12905
rect 191 12828 289 12849
rect 191 12668 289 12689
rect 191 12612 212 12668
rect 268 12612 289 12668
rect 191 12591 289 12612
rect 191 12431 289 12452
rect 191 12375 212 12431
rect 268 12375 289 12431
rect 191 12354 289 12375
rect 191 12115 289 12136
rect 191 12059 212 12115
rect 268 12059 289 12115
rect 191 12038 289 12059
rect 191 11878 289 11899
rect 191 11822 212 11878
rect 268 11822 289 11878
rect 191 11801 289 11822
rect 191 11641 289 11662
rect 191 11585 212 11641
rect 268 11585 289 11641
rect 191 11564 289 11585
rect 191 11325 289 11346
rect 191 11269 212 11325
rect 268 11269 289 11325
rect 191 11248 289 11269
rect 191 11088 289 11109
rect 191 11032 212 11088
rect 268 11032 289 11088
rect 191 11011 289 11032
rect 191 10851 289 10872
rect 191 10795 212 10851
rect 268 10795 289 10851
rect 191 10774 289 10795
rect 191 10535 289 10556
rect 191 10479 212 10535
rect 268 10479 289 10535
rect 191 10458 289 10479
rect 191 10298 289 10319
rect 191 10242 212 10298
rect 268 10242 289 10298
rect 191 10221 289 10242
rect 191 10061 289 10082
rect 191 10005 212 10061
rect 268 10005 289 10061
rect 191 9984 289 10005
rect 191 9745 289 9766
rect 191 9689 212 9745
rect 268 9689 289 9745
rect 191 9668 289 9689
rect 191 9508 289 9529
rect 191 9452 212 9508
rect 268 9452 289 9508
rect 191 9431 289 9452
rect 191 9271 289 9292
rect 191 9215 212 9271
rect 268 9215 289 9271
rect 191 9194 289 9215
rect 191 8955 289 8976
rect 191 8899 212 8955
rect 268 8899 289 8955
rect 191 8878 289 8899
rect 191 8718 289 8739
rect 191 8662 212 8718
rect 268 8662 289 8718
rect 191 8641 289 8662
rect 191 8481 289 8502
rect 191 8425 212 8481
rect 268 8425 289 8481
rect 191 8404 289 8425
rect 191 8165 289 8186
rect 191 8109 212 8165
rect 268 8109 289 8165
rect 191 8088 289 8109
rect 191 7928 289 7949
rect 191 7872 212 7928
rect 268 7872 289 7928
rect 191 7851 289 7872
rect 191 7691 289 7712
rect 191 7635 212 7691
rect 268 7635 289 7691
rect 191 7614 289 7635
rect 191 7375 289 7396
rect 191 7319 212 7375
rect 268 7319 289 7375
rect 191 7298 289 7319
rect 191 7138 289 7159
rect 191 7082 212 7138
rect 268 7082 289 7138
rect 191 7061 289 7082
rect 191 6901 289 6922
rect 191 6845 212 6901
rect 268 6845 289 6901
rect 191 6824 289 6845
rect 191 6585 289 6606
rect 191 6529 212 6585
rect 268 6529 289 6585
rect 191 6508 289 6529
rect 191 6348 289 6369
rect 191 6292 212 6348
rect 268 6292 289 6348
rect 191 6271 289 6292
rect 191 6111 289 6132
rect 191 6055 212 6111
rect 268 6055 289 6111
rect 191 6034 289 6055
rect 191 5795 289 5816
rect 191 5739 212 5795
rect 268 5739 289 5795
rect 191 5718 289 5739
rect 191 5558 289 5579
rect 191 5502 212 5558
rect 268 5502 289 5558
rect 191 5481 289 5502
rect 191 5321 289 5342
rect 191 5265 212 5321
rect 268 5265 289 5321
rect 191 5244 289 5265
rect 191 5005 289 5026
rect 191 4949 212 5005
rect 268 4949 289 5005
rect 191 4928 289 4949
rect 191 4768 289 4789
rect 191 4712 212 4768
rect 268 4712 289 4768
rect 191 4691 289 4712
rect 191 4531 289 4552
rect 191 4475 212 4531
rect 268 4475 289 4531
rect 191 4454 289 4475
rect 191 4215 289 4236
rect 191 4159 212 4215
rect 268 4159 289 4215
rect 191 4138 289 4159
rect 191 3978 289 3999
rect 191 3922 212 3978
rect 268 3922 289 3978
rect 191 3901 289 3922
rect 191 3741 289 3762
rect 191 3685 212 3741
rect 268 3685 289 3741
rect 191 3664 289 3685
rect 191 3425 289 3446
rect 191 3369 212 3425
rect 268 3369 289 3425
rect 191 3348 289 3369
rect 191 3188 289 3209
rect 191 3132 212 3188
rect 268 3132 289 3188
rect 191 3111 289 3132
rect 191 2951 289 2972
rect 191 2895 212 2951
rect 268 2895 289 2951
rect 191 2874 289 2895
rect 191 2635 289 2656
rect 191 2579 212 2635
rect 268 2579 289 2635
rect 191 2558 289 2579
rect 191 2398 289 2419
rect 191 2342 212 2398
rect 268 2342 289 2398
rect 191 2321 289 2342
rect 191 2161 289 2182
rect 191 2105 212 2161
rect 268 2105 289 2161
rect 191 2084 289 2105
rect 191 1845 289 1866
rect 191 1789 212 1845
rect 268 1789 289 1845
rect 191 1768 289 1789
rect 191 1608 289 1629
rect 191 1552 212 1608
rect 268 1552 289 1608
rect 191 1531 289 1552
rect 191 1371 289 1392
rect 191 1315 212 1371
rect 268 1315 289 1371
rect 191 1294 289 1315
rect 191 1055 289 1076
rect 191 999 212 1055
rect 268 999 289 1055
rect 191 978 289 999
rect 191 818 289 839
rect 191 762 212 818
rect 268 762 289 818
rect 191 741 289 762
rect 191 581 289 602
rect 191 525 212 581
rect 268 525 289 581
rect 191 504 289 525
use contact_9  contact_9_0
timestamp 1707688321
transform 1 0 207 0 1 516
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1707688321
transform 1 0 207 0 1 1306
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1707688321
transform 1 0 207 0 1 753
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1707688321
transform 1 0 207 0 1 990
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1707688321
transform 1 0 207 0 1 12840
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1707688321
transform 1 0 207 0 1 12603
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1707688321
transform 1 0 207 0 1 12366
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1707688321
transform 1 0 207 0 1 12050
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1707688321
transform 1 0 207 0 1 11813
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1707688321
transform 1 0 207 0 1 11576
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1707688321
transform 1 0 207 0 1 11260
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1707688321
transform 1 0 207 0 1 11023
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1707688321
transform 1 0 207 0 1 10786
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1707688321
transform 1 0 207 0 1 10470
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1707688321
transform 1 0 207 0 1 10233
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1707688321
transform 1 0 207 0 1 9996
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1707688321
transform 1 0 207 0 1 9680
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1707688321
transform 1 0 207 0 1 9443
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1707688321
transform 1 0 207 0 1 9206
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1707688321
transform 1 0 207 0 1 8890
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1707688321
transform 1 0 207 0 1 8653
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1707688321
transform 1 0 207 0 1 8416
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1707688321
transform 1 0 207 0 1 8100
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1707688321
transform 1 0 207 0 1 7863
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1707688321
transform 1 0 207 0 1 7626
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1707688321
transform 1 0 207 0 1 7310
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1707688321
transform 1 0 207 0 1 7073
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1707688321
transform 1 0 207 0 1 6836
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1707688321
transform 1 0 207 0 1 6520
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1707688321
transform 1 0 207 0 1 6283
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1707688321
transform 1 0 207 0 1 6046
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1707688321
transform 1 0 207 0 1 5730
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1707688321
transform 1 0 207 0 1 5493
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1707688321
transform 1 0 207 0 1 5256
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1707688321
transform 1 0 207 0 1 4940
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1707688321
transform 1 0 207 0 1 4703
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1707688321
transform 1 0 207 0 1 4466
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1707688321
transform 1 0 207 0 1 4150
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1707688321
transform 1 0 207 0 1 3913
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1707688321
transform 1 0 207 0 1 3676
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1707688321
transform 1 0 207 0 1 3360
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1707688321
transform 1 0 207 0 1 3123
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1707688321
transform 1 0 207 0 1 2886
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1707688321
transform 1 0 207 0 1 2570
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1707688321
transform 1 0 207 0 1 2333
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1707688321
transform 1 0 207 0 1 2096
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1707688321
transform 1 0 207 0 1 1780
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1707688321
transform 1 0 207 0 1 1543
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1707688321
transform 1 0 207 0 1 25796
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1707688321
transform 1 0 207 0 1 25480
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1707688321
transform 1 0 207 0 1 25243
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1707688321
transform 1 0 207 0 1 25006
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1707688321
transform 1 0 207 0 1 24690
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1707688321
transform 1 0 207 0 1 24453
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1707688321
transform 1 0 207 0 1 24216
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1707688321
transform 1 0 207 0 1 23900
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1707688321
transform 1 0 207 0 1 23663
box 0 0 1 1
use contact_9  contact_9_57
timestamp 1707688321
transform 1 0 207 0 1 23426
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1707688321
transform 1 0 207 0 1 23110
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1707688321
transform 1 0 207 0 1 22873
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1707688321
transform 1 0 207 0 1 22636
box 0 0 1 1
use contact_9  contact_9_61
timestamp 1707688321
transform 1 0 207 0 1 22320
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1707688321
transform 1 0 207 0 1 22083
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1707688321
transform 1 0 207 0 1 21846
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1707688321
transform 1 0 207 0 1 21530
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1707688321
transform 1 0 207 0 1 21293
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1707688321
transform 1 0 207 0 1 21056
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1707688321
transform 1 0 207 0 1 20740
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1707688321
transform 1 0 207 0 1 20503
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1707688321
transform 1 0 207 0 1 20266
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1707688321
transform 1 0 207 0 1 19950
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1707688321
transform 1 0 207 0 1 19713
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1707688321
transform 1 0 207 0 1 19476
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1707688321
transform 1 0 207 0 1 19160
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1707688321
transform 1 0 207 0 1 18923
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1707688321
transform 1 0 207 0 1 18686
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1707688321
transform 1 0 207 0 1 18370
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1707688321
transform 1 0 207 0 1 18133
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1707688321
transform 1 0 207 0 1 17896
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1707688321
transform 1 0 207 0 1 17580
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1707688321
transform 1 0 207 0 1 17343
box 0 0 1 1
use contact_9  contact_9_81
timestamp 1707688321
transform 1 0 207 0 1 17106
box 0 0 1 1
use contact_9  contact_9_82
timestamp 1707688321
transform 1 0 207 0 1 16790
box 0 0 1 1
use contact_9  contact_9_83
timestamp 1707688321
transform 1 0 207 0 1 16553
box 0 0 1 1
use contact_9  contact_9_84
timestamp 1707688321
transform 1 0 207 0 1 16316
box 0 0 1 1
use contact_9  contact_9_85
timestamp 1707688321
transform 1 0 207 0 1 16000
box 0 0 1 1
use contact_9  contact_9_86
timestamp 1707688321
transform 1 0 207 0 1 15763
box 0 0 1 1
use contact_9  contact_9_87
timestamp 1707688321
transform 1 0 207 0 1 15526
box 0 0 1 1
use contact_9  contact_9_88
timestamp 1707688321
transform 1 0 207 0 1 15210
box 0 0 1 1
use contact_9  contact_9_89
timestamp 1707688321
transform 1 0 207 0 1 14973
box 0 0 1 1
use contact_9  contact_9_90
timestamp 1707688321
transform 1 0 207 0 1 14736
box 0 0 1 1
use contact_9  contact_9_91
timestamp 1707688321
transform 1 0 207 0 1 14420
box 0 0 1 1
use contact_9  contact_9_92
timestamp 1707688321
transform 1 0 207 0 1 14183
box 0 0 1 1
use contact_9  contact_9_93
timestamp 1707688321
transform 1 0 207 0 1 13946
box 0 0 1 1
use contact_9  contact_9_94
timestamp 1707688321
transform 1 0 207 0 1 13630
box 0 0 1 1
use contact_9  contact_9_95
timestamp 1707688321
transform 1 0 207 0 1 13393
box 0 0 1 1
use contact_9  contact_9_96
timestamp 1707688321
transform 1 0 207 0 1 13156
box 0 0 1 1
use contact_9  contact_9_97
timestamp 1707688321
transform 1 0 207 0 1 26270
box 0 0 1 1
use contact_9  contact_9_98
timestamp 1707688321
transform 1 0 207 0 1 38673
box 0 0 1 1
use contact_9  contact_9_99
timestamp 1707688321
transform 1 0 207 0 1 38436
box 0 0 1 1
use contact_9  contact_9_100
timestamp 1707688321
transform 1 0 207 0 1 38120
box 0 0 1 1
use contact_9  contact_9_101
timestamp 1707688321
transform 1 0 207 0 1 37883
box 0 0 1 1
use contact_9  contact_9_102
timestamp 1707688321
transform 1 0 207 0 1 37646
box 0 0 1 1
use contact_9  contact_9_103
timestamp 1707688321
transform 1 0 207 0 1 37330
box 0 0 1 1
use contact_9  contact_9_104
timestamp 1707688321
transform 1 0 207 0 1 37093
box 0 0 1 1
use contact_9  contact_9_105
timestamp 1707688321
transform 1 0 207 0 1 36856
box 0 0 1 1
use contact_9  contact_9_106
timestamp 1707688321
transform 1 0 207 0 1 36540
box 0 0 1 1
use contact_9  contact_9_107
timestamp 1707688321
transform 1 0 207 0 1 36303
box 0 0 1 1
use contact_9  contact_9_108
timestamp 1707688321
transform 1 0 207 0 1 36066
box 0 0 1 1
use contact_9  contact_9_109
timestamp 1707688321
transform 1 0 207 0 1 35750
box 0 0 1 1
use contact_9  contact_9_110
timestamp 1707688321
transform 1 0 207 0 1 35513
box 0 0 1 1
use contact_9  contact_9_111
timestamp 1707688321
transform 1 0 207 0 1 35276
box 0 0 1 1
use contact_9  contact_9_112
timestamp 1707688321
transform 1 0 207 0 1 34960
box 0 0 1 1
use contact_9  contact_9_113
timestamp 1707688321
transform 1 0 207 0 1 34723
box 0 0 1 1
use contact_9  contact_9_114
timestamp 1707688321
transform 1 0 207 0 1 34486
box 0 0 1 1
use contact_9  contact_9_115
timestamp 1707688321
transform 1 0 207 0 1 34170
box 0 0 1 1
use contact_9  contact_9_116
timestamp 1707688321
transform 1 0 207 0 1 33933
box 0 0 1 1
use contact_9  contact_9_117
timestamp 1707688321
transform 1 0 207 0 1 33696
box 0 0 1 1
use contact_9  contact_9_118
timestamp 1707688321
transform 1 0 207 0 1 33380
box 0 0 1 1
use contact_9  contact_9_119
timestamp 1707688321
transform 1 0 207 0 1 33143
box 0 0 1 1
use contact_9  contact_9_120
timestamp 1707688321
transform 1 0 207 0 1 32906
box 0 0 1 1
use contact_9  contact_9_121
timestamp 1707688321
transform 1 0 207 0 1 32590
box 0 0 1 1
use contact_9  contact_9_122
timestamp 1707688321
transform 1 0 207 0 1 32353
box 0 0 1 1
use contact_9  contact_9_123
timestamp 1707688321
transform 1 0 207 0 1 32116
box 0 0 1 1
use contact_9  contact_9_124
timestamp 1707688321
transform 1 0 207 0 1 31800
box 0 0 1 1
use contact_9  contact_9_125
timestamp 1707688321
transform 1 0 207 0 1 31563
box 0 0 1 1
use contact_9  contact_9_126
timestamp 1707688321
transform 1 0 207 0 1 31326
box 0 0 1 1
use contact_9  contact_9_127
timestamp 1707688321
transform 1 0 207 0 1 31010
box 0 0 1 1
use contact_9  contact_9_128
timestamp 1707688321
transform 1 0 207 0 1 30773
box 0 0 1 1
use contact_9  contact_9_129
timestamp 1707688321
transform 1 0 207 0 1 30536
box 0 0 1 1
use contact_9  contact_9_130
timestamp 1707688321
transform 1 0 207 0 1 30220
box 0 0 1 1
use contact_9  contact_9_131
timestamp 1707688321
transform 1 0 207 0 1 29983
box 0 0 1 1
use contact_9  contact_9_132
timestamp 1707688321
transform 1 0 207 0 1 29746
box 0 0 1 1
use contact_9  contact_9_133
timestamp 1707688321
transform 1 0 207 0 1 29430
box 0 0 1 1
use contact_9  contact_9_134
timestamp 1707688321
transform 1 0 207 0 1 29193
box 0 0 1 1
use contact_9  contact_9_135
timestamp 1707688321
transform 1 0 207 0 1 28956
box 0 0 1 1
use contact_9  contact_9_136
timestamp 1707688321
transform 1 0 207 0 1 28640
box 0 0 1 1
use contact_9  contact_9_137
timestamp 1707688321
transform 1 0 207 0 1 28403
box 0 0 1 1
use contact_9  contact_9_138
timestamp 1707688321
transform 1 0 207 0 1 28166
box 0 0 1 1
use contact_9  contact_9_139
timestamp 1707688321
transform 1 0 207 0 1 27850
box 0 0 1 1
use contact_9  contact_9_140
timestamp 1707688321
transform 1 0 207 0 1 27613
box 0 0 1 1
use contact_9  contact_9_141
timestamp 1707688321
transform 1 0 207 0 1 27376
box 0 0 1 1
use contact_9  contact_9_142
timestamp 1707688321
transform 1 0 207 0 1 27060
box 0 0 1 1
use contact_9  contact_9_143
timestamp 1707688321
transform 1 0 207 0 1 26823
box 0 0 1 1
use contact_9  contact_9_144
timestamp 1707688321
transform 1 0 207 0 1 26586
box 0 0 1 1
use contact_9  contact_9_145
timestamp 1707688321
transform 1 0 207 0 1 51550
box 0 0 1 1
use contact_9  contact_9_146
timestamp 1707688321
transform 1 0 207 0 1 51313
box 0 0 1 1
use contact_9  contact_9_147
timestamp 1707688321
transform 1 0 207 0 1 51076
box 0 0 1 1
use contact_9  contact_9_148
timestamp 1707688321
transform 1 0 207 0 1 50760
box 0 0 1 1
use contact_9  contact_9_149
timestamp 1707688321
transform 1 0 207 0 1 50523
box 0 0 1 1
use contact_9  contact_9_150
timestamp 1707688321
transform 1 0 207 0 1 50286
box 0 0 1 1
use contact_9  contact_9_151
timestamp 1707688321
transform 1 0 207 0 1 49970
box 0 0 1 1
use contact_9  contact_9_152
timestamp 1707688321
transform 1 0 207 0 1 49733
box 0 0 1 1
use contact_9  contact_9_153
timestamp 1707688321
transform 1 0 207 0 1 49496
box 0 0 1 1
use contact_9  contact_9_154
timestamp 1707688321
transform 1 0 207 0 1 49180
box 0 0 1 1
use contact_9  contact_9_155
timestamp 1707688321
transform 1 0 207 0 1 48943
box 0 0 1 1
use contact_9  contact_9_156
timestamp 1707688321
transform 1 0 207 0 1 48706
box 0 0 1 1
use contact_9  contact_9_157
timestamp 1707688321
transform 1 0 207 0 1 48390
box 0 0 1 1
use contact_9  contact_9_158
timestamp 1707688321
transform 1 0 207 0 1 48153
box 0 0 1 1
use contact_9  contact_9_159
timestamp 1707688321
transform 1 0 207 0 1 47916
box 0 0 1 1
use contact_9  contact_9_160
timestamp 1707688321
transform 1 0 207 0 1 47600
box 0 0 1 1
use contact_9  contact_9_161
timestamp 1707688321
transform 1 0 207 0 1 47363
box 0 0 1 1
use contact_9  contact_9_162
timestamp 1707688321
transform 1 0 207 0 1 47126
box 0 0 1 1
use contact_9  contact_9_163
timestamp 1707688321
transform 1 0 207 0 1 46810
box 0 0 1 1
use contact_9  contact_9_164
timestamp 1707688321
transform 1 0 207 0 1 46573
box 0 0 1 1
use contact_9  contact_9_165
timestamp 1707688321
transform 1 0 207 0 1 46336
box 0 0 1 1
use contact_9  contact_9_166
timestamp 1707688321
transform 1 0 207 0 1 46020
box 0 0 1 1
use contact_9  contact_9_167
timestamp 1707688321
transform 1 0 207 0 1 45783
box 0 0 1 1
use contact_9  contact_9_168
timestamp 1707688321
transform 1 0 207 0 1 45546
box 0 0 1 1
use contact_9  contact_9_169
timestamp 1707688321
transform 1 0 207 0 1 45230
box 0 0 1 1
use contact_9  contact_9_170
timestamp 1707688321
transform 1 0 207 0 1 44993
box 0 0 1 1
use contact_9  contact_9_171
timestamp 1707688321
transform 1 0 207 0 1 44756
box 0 0 1 1
use contact_9  contact_9_172
timestamp 1707688321
transform 1 0 207 0 1 44440
box 0 0 1 1
use contact_9  contact_9_173
timestamp 1707688321
transform 1 0 207 0 1 44203
box 0 0 1 1
use contact_9  contact_9_174
timestamp 1707688321
transform 1 0 207 0 1 43966
box 0 0 1 1
use contact_9  contact_9_175
timestamp 1707688321
transform 1 0 207 0 1 43650
box 0 0 1 1
use contact_9  contact_9_176
timestamp 1707688321
transform 1 0 207 0 1 43413
box 0 0 1 1
use contact_9  contact_9_177
timestamp 1707688321
transform 1 0 207 0 1 43176
box 0 0 1 1
use contact_9  contact_9_178
timestamp 1707688321
transform 1 0 207 0 1 42860
box 0 0 1 1
use contact_9  contact_9_179
timestamp 1707688321
transform 1 0 207 0 1 42623
box 0 0 1 1
use contact_9  contact_9_180
timestamp 1707688321
transform 1 0 207 0 1 42386
box 0 0 1 1
use contact_9  contact_9_181
timestamp 1707688321
transform 1 0 207 0 1 42070
box 0 0 1 1
use contact_9  contact_9_182
timestamp 1707688321
transform 1 0 207 0 1 41833
box 0 0 1 1
use contact_9  contact_9_183
timestamp 1707688321
transform 1 0 207 0 1 41596
box 0 0 1 1
use contact_9  contact_9_184
timestamp 1707688321
transform 1 0 207 0 1 41280
box 0 0 1 1
use contact_9  contact_9_185
timestamp 1707688321
transform 1 0 207 0 1 41043
box 0 0 1 1
use contact_9  contact_9_186
timestamp 1707688321
transform 1 0 207 0 1 40806
box 0 0 1 1
use contact_9  contact_9_187
timestamp 1707688321
transform 1 0 207 0 1 40490
box 0 0 1 1
use contact_9  contact_9_188
timestamp 1707688321
transform 1 0 207 0 1 40253
box 0 0 1 1
use contact_9  contact_9_189
timestamp 1707688321
transform 1 0 207 0 1 40016
box 0 0 1 1
use contact_9  contact_9_190
timestamp 1707688321
transform 1 0 207 0 1 39700
box 0 0 1 1
use contact_9  contact_9_191
timestamp 1707688321
transform 1 0 207 0 1 39463
box 0 0 1 1
use contact_9  contact_9_192
timestamp 1707688321
transform 1 0 207 0 1 39226
box 0 0 1 1
use contact_9  contact_9_193
timestamp 1707688321
transform 1 0 207 0 1 38910
box 0 0 1 1
use contact_9  contact_9_194
timestamp 1707688321
transform 1 0 207 0 1 26033
box 0 0 1 1
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_0
timestamp 1707688321
transform 1 0 0 0 -1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_1
timestamp 1707688321
transform 1 0 0 0 -1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_2
timestamp 1707688321
transform 1 0 0 0 1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_3
timestamp 1707688321
transform 1 0 0 0 -1 1580
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_4
timestamp 1707688321
transform 1 0 0 0 1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_5
timestamp 1707688321
transform 1 0 0 0 -1 790
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_6
timestamp 1707688321
transform 1 0 0 0 1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_7
timestamp 1707688321
transform 1 0 0 0 -1 3950
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_8
timestamp 1707688321
transform 1 0 0 0 1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_9
timestamp 1707688321
transform 1 0 0 0 -1 3160
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_10
timestamp 1707688321
transform 1 0 0 0 1 2370
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_11
timestamp 1707688321
transform 1 0 0 0 1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_12
timestamp 1707688321
transform 1 0 0 0 -1 12640
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_13
timestamp 1707688321
transform 1 0 0 0 1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_14
timestamp 1707688321
transform 1 0 0 0 -1 11850
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_15
timestamp 1707688321
transform 1 0 0 0 1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_16
timestamp 1707688321
transform 1 0 0 0 -1 11060
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_17
timestamp 1707688321
transform 1 0 0 0 1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_18
timestamp 1707688321
transform 1 0 0 0 -1 10270
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_19
timestamp 1707688321
transform 1 0 0 0 1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_20
timestamp 1707688321
transform 1 0 0 0 -1 9480
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_21
timestamp 1707688321
transform 1 0 0 0 1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_22
timestamp 1707688321
transform 1 0 0 0 -1 8690
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_23
timestamp 1707688321
transform 1 0 0 0 1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_24
timestamp 1707688321
transform 1 0 0 0 -1 7900
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_25
timestamp 1707688321
transform 1 0 0 0 1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_26
timestamp 1707688321
transform 1 0 0 0 -1 7110
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_27
timestamp 1707688321
transform 1 0 0 0 1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_28
timestamp 1707688321
transform 1 0 0 0 -1 6320
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_29
timestamp 1707688321
transform 1 0 0 0 1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_30
timestamp 1707688321
transform 1 0 0 0 -1 5530
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_31
timestamp 1707688321
transform 1 0 0 0 1 4740
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_32
timestamp 1707688321
transform 1 0 0 0 1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_33
timestamp 1707688321
transform 1 0 0 0 1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_34
timestamp 1707688321
transform 1 0 0 0 -1 25280
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_35
timestamp 1707688321
transform 1 0 0 0 1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_36
timestamp 1707688321
transform 1 0 0 0 -1 24490
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_37
timestamp 1707688321
transform 1 0 0 0 1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_38
timestamp 1707688321
transform 1 0 0 0 -1 23700
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_39
timestamp 1707688321
transform 1 0 0 0 1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_40
timestamp 1707688321
transform 1 0 0 0 -1 22910
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_41
timestamp 1707688321
transform 1 0 0 0 1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_42
timestamp 1707688321
transform 1 0 0 0 -1 22120
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_43
timestamp 1707688321
transform 1 0 0 0 1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_44
timestamp 1707688321
transform 1 0 0 0 -1 21330
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_45
timestamp 1707688321
transform 1 0 0 0 1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_46
timestamp 1707688321
transform 1 0 0 0 -1 20540
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_47
timestamp 1707688321
transform 1 0 0 0 1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_48
timestamp 1707688321
transform 1 0 0 0 -1 19750
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_49
timestamp 1707688321
transform 1 0 0 0 1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_50
timestamp 1707688321
transform 1 0 0 0 -1 18960
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_51
timestamp 1707688321
transform 1 0 0 0 1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_52
timestamp 1707688321
transform 1 0 0 0 -1 18170
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_53
timestamp 1707688321
transform 1 0 0 0 1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_54
timestamp 1707688321
transform 1 0 0 0 -1 17380
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_55
timestamp 1707688321
transform 1 0 0 0 1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_56
timestamp 1707688321
transform 1 0 0 0 -1 16590
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_57
timestamp 1707688321
transform 1 0 0 0 1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_58
timestamp 1707688321
transform 1 0 0 0 -1 15800
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_59
timestamp 1707688321
transform 1 0 0 0 1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_60
timestamp 1707688321
transform 1 0 0 0 -1 15010
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_61
timestamp 1707688321
transform 1 0 0 0 1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_62
timestamp 1707688321
transform 1 0 0 0 -1 14220
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_63
timestamp 1707688321
transform 1 0 0 0 -1 13430
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_64
timestamp 1707688321
transform 1 0 0 0 -1 30020
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_65
timestamp 1707688321
transform 1 0 0 0 1 29230
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_66
timestamp 1707688321
transform 1 0 0 0 -1 29230
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_67
timestamp 1707688321
transform 1 0 0 0 1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_68
timestamp 1707688321
transform 1 0 0 0 -1 26860
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_69
timestamp 1707688321
transform 1 0 0 0 1 28440
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_70
timestamp 1707688321
transform 1 0 0 0 -1 28440
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_71
timestamp 1707688321
transform 1 0 0 0 1 27650
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_72
timestamp 1707688321
transform 1 0 0 0 -1 27650
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_73
timestamp 1707688321
transform 1 0 0 0 -1 38710
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_74
timestamp 1707688321
transform 1 0 0 0 1 37920
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_75
timestamp 1707688321
transform 1 0 0 0 -1 37920
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_76
timestamp 1707688321
transform 1 0 0 0 1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_77
timestamp 1707688321
transform 1 0 0 0 -1 37130
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_78
timestamp 1707688321
transform 1 0 0 0 1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_79
timestamp 1707688321
transform 1 0 0 0 -1 36340
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_80
timestamp 1707688321
transform 1 0 0 0 1 35550
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_81
timestamp 1707688321
transform 1 0 0 0 -1 35550
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_82
timestamp 1707688321
transform 1 0 0 0 1 34760
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_83
timestamp 1707688321
transform 1 0 0 0 -1 34760
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_84
timestamp 1707688321
transform 1 0 0 0 1 33970
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_85
timestamp 1707688321
transform 1 0 0 0 -1 33970
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_86
timestamp 1707688321
transform 1 0 0 0 1 33180
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_87
timestamp 1707688321
transform 1 0 0 0 -1 33180
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_88
timestamp 1707688321
transform 1 0 0 0 1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_89
timestamp 1707688321
transform 1 0 0 0 -1 32390
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_90
timestamp 1707688321
transform 1 0 0 0 1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_91
timestamp 1707688321
transform 1 0 0 0 -1 31600
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_92
timestamp 1707688321
transform 1 0 0 0 1 30810
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_93
timestamp 1707688321
transform 1 0 0 0 -1 30810
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_94
timestamp 1707688321
transform 1 0 0 0 1 30020
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_95
timestamp 1707688321
transform 1 0 0 0 -1 39500
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_96
timestamp 1707688321
transform 1 0 0 0 1 51350
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_97
timestamp 1707688321
transform 1 0 0 0 -1 51350
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_98
timestamp 1707688321
transform 1 0 0 0 1 50560
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_99
timestamp 1707688321
transform 1 0 0 0 -1 50560
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_100
timestamp 1707688321
transform 1 0 0 0 1 49770
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_101
timestamp 1707688321
transform 1 0 0 0 -1 49770
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_102
timestamp 1707688321
transform 1 0 0 0 1 48980
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_103
timestamp 1707688321
transform 1 0 0 0 -1 48980
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_104
timestamp 1707688321
transform 1 0 0 0 1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_105
timestamp 1707688321
transform 1 0 0 0 -1 48190
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_106
timestamp 1707688321
transform 1 0 0 0 1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_107
timestamp 1707688321
transform 1 0 0 0 -1 47400
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_108
timestamp 1707688321
transform 1 0 0 0 1 46610
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_109
timestamp 1707688321
transform 1 0 0 0 -1 46610
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_110
timestamp 1707688321
transform 1 0 0 0 1 45820
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_111
timestamp 1707688321
transform 1 0 0 0 -1 45820
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_112
timestamp 1707688321
transform 1 0 0 0 1 45030
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_113
timestamp 1707688321
transform 1 0 0 0 -1 45030
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_114
timestamp 1707688321
transform 1 0 0 0 1 44240
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_115
timestamp 1707688321
transform 1 0 0 0 -1 44240
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_116
timestamp 1707688321
transform 1 0 0 0 1 43450
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_117
timestamp 1707688321
transform 1 0 0 0 -1 43450
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_118
timestamp 1707688321
transform 1 0 0 0 1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_119
timestamp 1707688321
transform 1 0 0 0 -1 42660
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_120
timestamp 1707688321
transform 1 0 0 0 1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_121
timestamp 1707688321
transform 1 0 0 0 -1 41870
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_122
timestamp 1707688321
transform 1 0 0 0 1 41080
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_123
timestamp 1707688321
transform 1 0 0 0 -1 41080
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_124
timestamp 1707688321
transform 1 0 0 0 1 40290
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_125
timestamp 1707688321
transform 1 0 0 0 -1 40290
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_126
timestamp 1707688321
transform 1 0 0 0 1 39500
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_127
timestamp 1707688321
transform 1 0 0 0 1 38710
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_128
timestamp 1707688321
transform 1 0 0 0 1 26070
box -42 -55 624 371
use sky130_fd_bd_sram__openram_dp_cell_cap_row_3  sky130_fd_bd_sram__openram_dp_cell_cap_row_129
timestamp 1707688321
transform 1 0 0 0 -1 26070
box -42 -55 624 371
<< labels >>
rlabel metal2 s 312 40953 312 40953 4 wl1_103
port 1 nsew
rlabel metal2 s 312 46263 312 46263 4 wl0_117
port 2 nsew
rlabel metal2 s 312 48537 312 48537 4 wl0_122
port 3 nsew
rlabel metal2 s 312 39057 312 39057 4 wl0_98
port 4 nsew
rlabel metal2 s 312 47747 312 47747 4 wl0_120
port 5 nsew
rlabel metal2 s 312 39847 312 39847 4 wl0_100
port 6 nsew
rlabel metal2 s 312 44683 312 44683 4 wl0_113
port 7 nsew
rlabel metal2 s 312 42787 312 42787 4 wl1_108
port 8 nsew
rlabel metal2 s 312 50687 312 50687 4 wl1_128
port 9 nsew
rlabel metal2 s 312 47273 312 47273 4 wl1_119
port 10 nsew
rlabel metal2 s 312 39627 312 39627 4 wl1_100
port 11 nsew
rlabel metal2 s 312 43893 312 43893 4 wl0_111
port 12 nsew
rlabel metal2 s 312 45947 312 45947 4 wl1_116
port 13 nsew
rlabel metal2 s 312 39153 312 39153 4 wl0_99
port 14 nsew
rlabel metal2 s 312 51223 312 51223 4 wl1_129
port 15 nsew
rlabel metal2 s 312 51477 312 51477 4 wl1_130
port 16 nsew
rlabel metal2 s 312 48063 312 48063 4 wl1_121
port 17 nsew
rlabel metal2 s 312 43577 312 43577 4 wl1_110
port 18 nsew
rlabel metal2 s 312 49643 312 49643 4 wl1_125
port 19 nsew
rlabel metal2 s 312 44113 312 44113 4 wl1_111
port 20 nsew
rlabel metal2 s 312 41743 312 41743 4 wl1_105
port 21 nsew
rlabel metal2 s 312 44903 312 44903 4 wl1_113
port 22 nsew
rlabel metal2 s 312 49107 312 49107 4 wl1_124
port 23 nsew
rlabel metal2 s 312 50433 312 50433 4 wl1_127
port 24 nsew
rlabel metal2 s 312 49327 312 49327 4 wl0_124
port 25 nsew
rlabel metal2 s 312 43007 312 43007 4 wl0_108
port 26 nsew
rlabel metal2 s 312 50117 312 50117 4 wl0_126
port 27 nsew
rlabel metal2 s 312 40637 312 40637 4 wl0_102
port 28 nsew
rlabel metal2 s 312 45377 312 45377 4 wl0_114
port 29 nsew
rlabel metal2 s 312 42533 312 42533 4 wl1_107
port 30 nsew
rlabel metal2 s 312 48853 312 48853 4 wl1_123
port 31 nsew
rlabel metal2 s 312 40417 312 40417 4 wl1_102
port 32 nsew
rlabel metal2 s 312 47843 312 47843 4 wl0_121
port 33 nsew
rlabel metal2 s 312 46957 312 46957 4 wl0_118
port 34 nsew
rlabel metal2 s 312 41523 312 41523 4 wl0_105
port 35 nsew
rlabel metal2 s 312 43797 312 43797 4 wl0_110
port 36 nsew
rlabel metal2 s 312 45157 312 45157 4 wl1_114
port 37 nsew
rlabel metal2 s 312 44367 312 44367 4 wl1_112
port 38 nsew
rlabel metal2 s 312 51697 312 51697 4 wl0_130
port 39 nsew
rlabel metal2 s 312 45473 312 45473 4 wl0_115
port 40 nsew
rlabel metal2 s 312 41997 312 41997 4 wl1_106
port 41 nsew
rlabel metal2 s 312 48317 312 48317 4 wl1_122
port 42 nsew
rlabel metal2 s 312 51003 312 51003 4 wl0_129
port 43 nsew
rlabel metal2 s 312 40163 312 40163 4 wl1_101
port 44 nsew
rlabel metal2 s 312 50213 312 50213 4 wl0_127
port 45 nsew
rlabel metal2 s 312 50907 312 50907 4 wl0_128
port 46 nsew
rlabel metal2 s 312 43103 312 43103 4 wl0_109
port 47 nsew
rlabel metal2 s 312 45693 312 45693 4 wl1_115
port 48 nsew
rlabel metal2 s 312 46167 312 46167 4 wl0_116
port 49 nsew
rlabel metal2 s 312 46483 312 46483 4 wl1_117
port 50 nsew
rlabel metal2 s 312 46737 312 46737 4 wl1_118
port 51 nsew
rlabel metal2 s 312 39943 312 39943 4 wl0_101
port 52 nsew
rlabel metal2 s 312 47527 312 47527 4 wl1_120
port 53 nsew
rlabel metal2 s 312 40733 312 40733 4 wl0_103
port 54 nsew
rlabel metal2 s 312 41427 312 41427 4 wl0_104
port 55 nsew
rlabel metal2 s 312 39373 312 39373 4 wl1_99
port 56 nsew
rlabel metal2 s 312 47053 312 47053 4 wl0_119
port 57 nsew
rlabel metal2 s 312 49897 312 49897 4 wl1_126
port 58 nsew
rlabel metal2 s 312 44587 312 44587 4 wl0_112
port 59 nsew
rlabel metal2 s 312 42217 312 42217 4 wl0_106
port 60 nsew
rlabel metal2 s 312 49423 312 49423 4 wl0_125
port 61 nsew
rlabel metal2 s 312 42313 312 42313 4 wl0_107
port 62 nsew
rlabel metal2 s 312 48633 312 48633 4 wl0_123
port 63 nsew
rlabel metal2 s 312 43323 312 43323 4 wl1_109
port 64 nsew
rlabel metal2 s 312 41207 312 41207 4 wl1_104
port 65 nsew
rlabel metal2 s 312 27207 312 27207 4 wl0_68
port 66 nsew
rlabel metal2 s 312 30683 312 30683 4 wl1_77
port 67 nsew
rlabel metal2 s 312 28787 312 28787 4 wl0_72
port 68 nsew
rlabel metal2 s 312 31473 312 31473 4 wl1_79
port 69 nsew
rlabel metal2 s 312 37257 312 37257 4 wl1_94
port 70 nsew
rlabel metal2 s 312 36687 312 36687 4 wl0_92
port 71 nsew
rlabel metal2 s 312 26197 312 26197 4 wl1_66
port 72 nsew
rlabel metal2 s 312 26733 312 26733 4 wl1_67
port 73 nsew
rlabel metal2 s 312 36783 312 36783 4 wl0_93
port 74 nsew
rlabel metal2 s 312 31727 312 31727 4 wl1_80
port 75 nsew
rlabel metal2 s 312 30463 312 30463 4 wl0_77
port 76 nsew
rlabel metal2 s 312 28093 312 28093 4 wl0_71
port 77 nsew
rlabel metal2 s 312 35423 312 35423 4 wl1_89
port 78 nsew
rlabel metal2 s 312 38267 312 38267 4 wl0_96
port 79 nsew
rlabel metal2 s 312 32043 312 32043 4 wl0_81
port 80 nsew
rlabel metal2 s 312 35993 312 35993 4 wl0_91
port 81 nsew
rlabel metal2 s 312 38583 312 38583 4 wl1_97
port 82 nsew
rlabel metal2 s 312 33307 312 33307 4 wl1_84
port 83 nsew
rlabel metal2 s 312 29673 312 29673 4 wl0_75
port 84 nsew
rlabel metal2 s 312 36213 312 36213 4 wl1_91
port 85 nsew
rlabel metal2 s 312 29103 312 29103 4 wl1_73
port 86 nsew
rlabel metal2 s 312 29357 312 29357 4 wl1_74
port 87 nsew
rlabel metal2 s 312 33623 312 33623 4 wl0_85
port 88 nsew
rlabel metal2 s 312 34887 312 34887 4 wl1_88
port 89 nsew
rlabel metal2 s 312 38837 312 38837 4 wl1_98
port 90 nsew
rlabel metal2 s 312 35107 312 35107 4 wl0_88
port 91 nsew
rlabel metal2 s 312 35677 312 35677 4 wl1_90
port 92 nsew
rlabel metal2 s 312 27777 312 27777 4 wl1_70
port 93 nsew
rlabel metal2 s 312 37477 312 37477 4 wl0_94
port 94 nsew
rlabel metal2 s 312 26513 312 26513 4 wl0_67
port 95 nsew
rlabel metal2 s 312 30147 312 30147 4 wl1_76
port 96 nsew
rlabel metal2 s 312 32833 312 32833 4 wl0_83
port 97 nsew
rlabel metal2 s 312 28313 312 28313 4 wl1_71
port 98 nsew
rlabel metal2 s 312 38363 312 38363 4 wl0_97
port 99 nsew
rlabel metal2 s 312 35897 312 35897 4 wl0_90
port 100 nsew
rlabel metal2 s 312 33843 312 33843 4 wl1_85
port 101 nsew
rlabel metal2 s 312 26987 312 26987 4 wl1_68
port 102 nsew
rlabel metal2 s 312 33053 312 33053 4 wl1_83
port 103 nsew
rlabel metal2 s 312 32517 312 32517 4 wl1_82
port 104 nsew
rlabel metal2 s 312 31253 312 31253 4 wl0_79
port 105 nsew
rlabel metal2 s 312 32737 312 32737 4 wl0_82
port 106 nsew
rlabel metal2 s 312 34413 312 34413 4 wl0_87
port 107 nsew
rlabel metal2 s 312 31947 312 31947 4 wl0_80
port 108 nsew
rlabel metal2 s 312 34317 312 34317 4 wl0_86
port 109 nsew
rlabel metal2 s 312 28567 312 28567 4 wl1_72
port 110 nsew
rlabel metal2 s 312 28883 312 28883 4 wl0_73
port 111 nsew
rlabel metal2 s 312 37793 312 37793 4 wl1_95
port 112 nsew
rlabel metal2 s 312 38047 312 38047 4 wl1_96
port 113 nsew
rlabel metal2 s 312 27303 312 27303 4 wl0_69
port 114 nsew
rlabel metal2 s 312 37573 312 37573 4 wl0_95
port 115 nsew
rlabel metal2 s 312 29577 312 29577 4 wl0_74
port 116 nsew
rlabel metal2 s 312 35203 312 35203 4 wl0_89
port 117 nsew
rlabel metal2 s 312 34097 312 34097 4 wl1_86
port 118 nsew
rlabel metal2 s 312 27997 312 27997 4 wl0_70
port 119 nsew
rlabel metal2 s 312 32263 312 32263 4 wl1_81
port 120 nsew
rlabel metal2 s 312 30937 312 30937 4 wl1_78
port 121 nsew
rlabel metal2 s 312 29893 312 29893 4 wl1_75
port 122 nsew
rlabel metal2 s 312 37003 312 37003 4 wl1_93
port 123 nsew
rlabel metal2 s 312 27523 312 27523 4 wl1_69
port 124 nsew
rlabel metal2 s 312 36467 312 36467 4 wl1_92
port 125 nsew
rlabel metal2 s 312 26417 312 26417 4 wl0_66
port 126 nsew
rlabel metal2 s 312 33527 312 33527 4 wl0_84
port 127 nsew
rlabel metal2 s 312 34633 312 34633 4 wl1_87
port 128 nsew
rlabel metal2 s 312 30367 312 30367 4 wl0_76
port 129 nsew
rlabel metal2 s 312 31157 312 31157 4 wl0_78
port 130 nsew
rlabel metal2 s 312 15673 312 15673 4 wl1_39
port 131 nsew
rlabel metal2 s 312 24617 312 24617 4 wl1_62
port 132 nsew
rlabel metal2 s 312 14883 312 14883 4 wl1_37
port 133 nsew
rlabel metal2 s 312 19877 312 19877 4 wl1_50
port 134 nsew
rlabel metal2 s 312 20413 312 20413 4 wl1_51
port 135 nsew
rlabel metal2 s 312 16717 312 16717 4 wl1_42
port 136 nsew
rlabel metal2 s 312 23257 312 23257 4 wl0_58
port 137 nsew
rlabel metal2 s 312 18517 312 18517 4 wl0_46
port 138 nsew
rlabel metal2 s 312 22247 312 22247 4 wl1_56
port 139 nsew
rlabel metal2 s 312 25943 312 25943 4 wl1_65
port 140 nsew
rlabel metal2 s 312 13873 312 13873 4 wl0_35
port 141 nsew
rlabel metal2 s 312 24143 312 24143 4 wl0_61
port 142 nsew
rlabel metal2 s 312 18833 312 18833 4 wl1_47
port 143 nsew
rlabel metal2 s 312 15137 312 15137 4 wl1_38
port 144 nsew
rlabel metal2 s 312 14663 312 14663 4 wl0_37
port 145 nsew
rlabel metal2 s 312 21993 312 21993 4 wl1_55
port 146 nsew
rlabel metal2 s 312 23573 312 23573 4 wl1_59
port 147 nsew
rlabel metal2 s 312 21773 312 21773 4 wl0_55
port 148 nsew
rlabel metal2 s 312 23827 312 23827 4 wl1_60
port 149 nsew
rlabel metal2 s 312 17033 312 17033 4 wl0_43
port 150 nsew
rlabel metal2 s 312 15357 312 15357 4 wl0_38
port 151 nsew
rlabel metal2 s 312 16147 312 16147 4 wl0_40
port 152 nsew
rlabel metal2 s 312 25407 312 25407 4 wl1_64
port 153 nsew
rlabel metal2 s 312 17253 312 17253 4 wl1_43
port 154 nsew
rlabel metal2 s 312 20887 312 20887 4 wl0_52
port 155 nsew
rlabel metal2 s 312 18613 312 18613 4 wl0_47
port 156 nsew
rlabel metal2 s 312 16243 312 16243 4 wl0_41
port 157 nsew
rlabel metal2 s 312 17507 312 17507 4 wl1_44
port 158 nsew
rlabel metal2 s 312 23353 312 23353 4 wl0_59
port 159 nsew
rlabel metal2 s 312 23037 312 23037 4 wl1_58
port 160 nsew
rlabel metal2 s 312 20097 312 20097 4 wl0_50
port 161 nsew
rlabel metal2 s 312 19307 312 19307 4 wl0_48
port 162 nsew
rlabel metal2 s 312 22563 312 22563 4 wl0_57
port 163 nsew
rlabel metal2 s 312 13303 312 13303 4 wl1_33
port 164 nsew
rlabel metal2 s 312 15453 312 15453 4 wl0_39
port 165 nsew
rlabel metal2 s 312 18043 312 18043 4 wl1_45
port 166 nsew
rlabel metal2 s 312 19087 312 19087 4 wl1_48
port 167 nsew
rlabel metal2 s 312 19623 312 19623 4 wl1_49
port 168 nsew
rlabel metal2 s 312 20193 312 20193 4 wl0_51
port 169 nsew
rlabel metal2 s 312 24047 312 24047 4 wl0_60
port 170 nsew
rlabel metal2 s 312 20667 312 20667 4 wl1_52
port 171 nsew
rlabel metal2 s 312 14347 312 14347 4 wl1_36
port 172 nsew
rlabel metal2 s 312 19403 312 19403 4 wl0_49
port 173 nsew
rlabel metal2 s 312 21203 312 21203 4 wl1_53
port 174 nsew
rlabel metal2 s 312 15927 312 15927 4 wl1_40
port 175 nsew
rlabel metal2 s 312 17823 312 17823 4 wl0_45
port 176 nsew
rlabel metal2 s 312 13557 312 13557 4 wl1_34
port 177 nsew
rlabel metal2 s 312 25627 312 25627 4 wl0_64
port 178 nsew
rlabel metal2 s 312 21457 312 21457 4 wl1_54
port 179 nsew
rlabel metal2 s 312 17727 312 17727 4 wl0_44
port 180 nsew
rlabel metal2 s 312 25723 312 25723 4 wl0_65
port 181 nsew
rlabel metal2 s 312 16463 312 16463 4 wl1_41
port 182 nsew
rlabel metal2 s 312 18297 312 18297 4 wl1_46
port 183 nsew
rlabel metal2 s 312 24363 312 24363 4 wl1_61
port 184 nsew
rlabel metal2 s 312 22783 312 22783 4 wl1_57
port 185 nsew
rlabel metal2 s 312 25153 312 25153 4 wl1_63
port 186 nsew
rlabel metal2 s 312 16937 312 16937 4 wl0_42
port 187 nsew
rlabel metal2 s 312 14093 312 14093 4 wl1_35
port 188 nsew
rlabel metal2 s 312 14567 312 14567 4 wl0_36
port 189 nsew
rlabel metal2 s 312 24837 312 24837 4 wl0_62
port 190 nsew
rlabel metal2 s 312 20983 312 20983 4 wl0_53
port 191 nsew
rlabel metal2 s 312 22467 312 22467 4 wl0_56
port 192 nsew
rlabel metal2 s 312 24933 312 24933 4 wl0_63
port 193 nsew
rlabel metal2 s 312 13777 312 13777 4 wl0_34
port 194 nsew
rlabel metal2 s 312 21677 312 21677 4 wl0_54
port 195 nsew
rlabel metal2 s 312 9607 312 9607 4 wl1_24
port 196 nsew
rlabel metal2 s 312 9133 312 9133 4 wl0_23
port 197 nsew
rlabel metal2 s 312 1707 312 1707 4 wl1_4
port 198 nsew
rlabel metal2 s 312 1137 312 1137 4 wl0_2
port 199 nsew
rlabel metal2 s 312 8343 312 8343 4 wl0_21
port 200 nsew
rlabel metal2 s 312 9923 312 9923 4 wl0_25
port 201 nsew
rlabel metal2 s 312 6193 312 6193 4 wl1_15
port 202 nsew
rlabel metal2 s 312 10713 312 10713 4 wl0_27
port 203 nsew
rlabel metal2 s 312 1233 312 1233 4 wl0_3
port 204 nsew
rlabel metal2 s 312 10143 312 10143 4 wl1_25
port 205 nsew
rlabel metal2 s 312 3823 312 3823 4 wl1_9
port 206 nsew
rlabel metal2 s 312 11977 312 11977 4 wl1_30
port 207 nsew
rlabel metal2 s 312 7773 312 7773 4 wl1_19
port 208 nsew
rlabel metal2 s 312 13083 312 13083 4 wl0_33
port 209 nsew
rlabel metal2 s 312 6763 312 6763 4 wl0_17
port 210 nsew
rlabel metal2 s 312 2813 312 2813 4 wl0_7
port 211 nsew
rlabel metal2 s 312 443 312 443 4 wl0_1
port 212 nsew
rlabel metal2 s 312 5403 312 5403 4 wl1_13
port 213 nsew
rlabel metal2 s 312 7553 312 7553 4 wl0_19
port 214 nsew
rlabel metal2 s 312 5183 312 5183 4 wl0_13
port 215 nsew
rlabel metal2 s 312 1927 312 1927 4 wl0_4
port 216 nsew
rlabel metal2 s 312 12293 312 12293 4 wl0_31
port 217 nsew
rlabel metal2 s 312 9353 312 9353 4 wl1_23
port 218 nsew
rlabel metal2 s 312 3603 312 3603 4 wl0_9
port 219 nsew
rlabel metal2 s 312 8247 312 8247 4 wl0_20
port 220 nsew
rlabel metal2 s 312 12767 312 12767 4 wl1_32
port 221 nsew
rlabel metal2 s 312 12987 312 12987 4 wl0_32
port 222 nsew
rlabel metal2 s 312 6447 312 6447 4 wl1_16
port 223 nsew
rlabel metal2 s 312 1453 312 1453 4 wl1_3
port 224 nsew
rlabel metal2 s 312 3033 312 3033 4 wl1_7
port 225 nsew
rlabel metal2 s 312 4077 312 4077 4 wl1_10
port 226 nsew
rlabel metal2 s 312 8563 312 8563 4 wl1_21
port 227 nsew
rlabel metal2 s 312 10617 312 10617 4 wl0_26
port 228 nsew
rlabel metal2 s 312 5087 312 5087 4 wl0_12
port 229 nsew
rlabel metal2 s 312 4613 312 4613 4 wl1_11
port 230 nsew
rlabel metal2 s 312 11503 312 11503 4 wl0_29
port 231 nsew
rlabel metal2 s 312 8027 312 8027 4 wl1_20
port 232 nsew
rlabel metal2 s 312 5877 312 5877 4 wl0_14
port 233 nsew
rlabel metal2 s 312 2243 312 2243 4 wl1_5
port 234 nsew
rlabel metal2 s 312 7457 312 7457 4 wl0_18
port 235 nsew
rlabel metal2 s 312 10397 312 10397 4 wl1_26
port 236 nsew
rlabel metal2 s 312 12197 312 12197 4 wl0_30
port 237 nsew
rlabel metal2 s 312 5657 312 5657 4 wl1_14
port 238 nsew
rlabel metal2 s 312 7237 312 7237 4 wl1_18
port 239 nsew
rlabel metal2 s 312 12513 312 12513 4 wl1_31
port 240 nsew
rlabel metal2 s 312 2717 312 2717 4 wl0_6
port 241 nsew
rlabel metal2 s 312 9037 312 9037 4 wl0_22
port 242 nsew
rlabel metal2 s 312 2497 312 2497 4 wl1_6
port 243 nsew
rlabel metal2 s 312 3287 312 3287 4 wl1_8
port 244 nsew
rlabel metal2 s 312 11187 312 11187 4 wl1_28
port 245 nsew
rlabel metal2 s 312 3507 312 3507 4 wl0_8
port 246 nsew
rlabel metal2 s 312 917 312 917 4 wl1_2
port 247 nsew
rlabel metal2 s 312 6667 312 6667 4 wl0_16
port 248 nsew
rlabel metal2 s 312 4297 312 4297 4 wl0_10
port 249 nsew
rlabel metal2 s 312 2023 312 2023 4 wl0_5
port 250 nsew
rlabel metal2 s 312 4867 312 4867 4 wl1_12
port 251 nsew
rlabel metal2 s 312 11723 312 11723 4 wl1_29
port 252 nsew
rlabel metal2 s 312 663 312 663 4 wl1_1
port 253 nsew
rlabel metal2 s 312 11407 312 11407 4 wl0_28
port 254 nsew
rlabel metal2 s 312 6983 312 6983 4 wl1_17
port 255 nsew
rlabel metal2 s 312 5973 312 5973 4 wl0_15
port 256 nsew
rlabel metal2 s 312 9827 312 9827 4 wl0_24
port 257 nsew
rlabel metal2 s 312 8817 312 8817 4 wl1_22
port 258 nsew
rlabel metal2 s 312 4393 312 4393 4 wl0_11
port 259 nsew
rlabel metal2 s 312 10933 312 10933 4 wl1_27
port 260 nsew
rlabel metal3 s 240 33970 240 33970 4 gnd
port 261 nsew
rlabel metal3 s 240 48190 240 48190 4 gnd
port 261 nsew
rlabel metal3 s 240 43687 240 43687 4 gnd
port 261 nsew
rlabel metal3 s 240 34523 240 34523 4 gnd
port 261 nsew
rlabel metal3 s 240 48427 240 48427 4 gnd
port 261 nsew
rlabel metal3 s 240 29783 240 29783 4 gnd
port 261 nsew
rlabel metal3 s 240 31047 240 31047 4 gnd
port 261 nsew
rlabel metal3 s 240 40053 240 40053 4 gnd
port 261 nsew
rlabel metal3 s 240 44240 240 44240 4 gnd
port 261 nsew
rlabel metal3 s 240 32627 240 32627 4 gnd
port 261 nsew
rlabel metal3 s 240 49533 240 49533 4 gnd
port 261 nsew
rlabel metal3 s 240 48980 240 48980 4 gnd
port 261 nsew
rlabel metal3 s 240 36103 240 36103 4 gnd
port 261 nsew
rlabel metal3 s 240 35313 240 35313 4 gnd
port 261 nsew
rlabel metal3 s 240 34760 240 34760 4 gnd
port 261 nsew
rlabel metal3 s 240 37920 240 37920 4 gnd
port 261 nsew
rlabel metal3 s 240 35550 240 35550 4 gnd
port 261 nsew
rlabel metal3 s 240 51350 240 51350 4 gnd
port 261 nsew
rlabel metal3 s 240 35787 240 35787 4 gnd
port 261 nsew
rlabel metal3 s 240 43450 240 43450 4 gnd
port 261 nsew
rlabel metal3 s 240 37683 240 37683 4 gnd
port 261 nsew
rlabel metal3 s 240 43213 240 43213 4 gnd
port 261 nsew
rlabel metal3 s 240 27887 240 27887 4 gnd
port 261 nsew
rlabel metal3 s 240 32943 240 32943 4 gnd
port 261 nsew
rlabel metal3 s 240 41870 240 41870 4 gnd
port 261 nsew
rlabel metal3 s 240 45267 240 45267 4 gnd
port 261 nsew
rlabel metal3 s 240 29467 240 29467 4 gnd
port 261 nsew
rlabel metal3 s 240 40290 240 40290 4 gnd
port 261 nsew
rlabel metal3 s 240 46610 240 46610 4 gnd
port 261 nsew
rlabel metal3 s 240 42423 240 42423 4 gnd
port 261 nsew
rlabel metal3 s 240 47400 240 47400 4 gnd
port 261 nsew
rlabel metal3 s 240 28677 240 28677 4 gnd
port 261 nsew
rlabel metal3 s 240 50007 240 50007 4 gnd
port 261 nsew
rlabel metal3 s 240 32153 240 32153 4 gnd
port 261 nsew
rlabel metal3 s 240 27413 240 27413 4 gnd
port 261 nsew
rlabel metal3 s 240 40843 240 40843 4 gnd
port 261 nsew
rlabel metal3 s 240 38947 240 38947 4 gnd
port 261 nsew
rlabel metal3 s 240 29230 240 29230 4 gnd
port 261 nsew
rlabel metal3 s 240 33180 240 33180 4 gnd
port 261 nsew
rlabel metal3 s 240 47163 240 47163 4 gnd
port 261 nsew
rlabel metal3 s 240 34997 240 34997 4 gnd
port 261 nsew
rlabel metal3 s 240 37367 240 37367 4 gnd
port 261 nsew
rlabel metal3 s 240 27650 240 27650 4 gnd
port 261 nsew
rlabel metal3 s 240 42897 240 42897 4 gnd
port 261 nsew
rlabel metal3 s 240 32390 240 32390 4 gnd
port 261 nsew
rlabel metal3 s 240 26307 240 26307 4 gnd
port 261 nsew
rlabel metal3 s 240 46373 240 46373 4 gnd
port 261 nsew
rlabel metal3 s 240 44793 240 44793 4 gnd
port 261 nsew
rlabel metal3 s 240 31600 240 31600 4 gnd
port 261 nsew
rlabel metal3 s 240 44003 240 44003 4 gnd
port 261 nsew
rlabel metal3 s 240 37130 240 37130 4 gnd
port 261 nsew
rlabel metal3 s 240 47637 240 47637 4 gnd
port 261 nsew
rlabel metal3 s 240 28993 240 28993 4 gnd
port 261 nsew
rlabel metal3 s 240 33417 240 33417 4 gnd
port 261 nsew
rlabel metal3 s 240 38157 240 38157 4 gnd
port 261 nsew
rlabel metal3 s 240 39500 240 39500 4 gnd
port 261 nsew
rlabel metal3 s 240 30573 240 30573 4 gnd
port 261 nsew
rlabel metal3 s 240 41080 240 41080 4 gnd
port 261 nsew
rlabel metal3 s 240 38710 240 38710 4 gnd
port 261 nsew
rlabel metal3 s 240 39263 240 39263 4 gnd
port 261 nsew
rlabel metal3 s 240 44477 240 44477 4 gnd
port 261 nsew
rlabel metal3 s 240 34207 240 34207 4 gnd
port 261 nsew
rlabel metal3 s 240 28203 240 28203 4 gnd
port 261 nsew
rlabel metal3 s 240 30257 240 30257 4 gnd
port 261 nsew
rlabel metal3 s 240 45030 240 45030 4 gnd
port 261 nsew
rlabel metal3 s 240 47953 240 47953 4 gnd
port 261 nsew
rlabel metal3 s 240 27097 240 27097 4 gnd
port 261 nsew
rlabel metal3 s 240 51113 240 51113 4 gnd
port 261 nsew
rlabel metal3 s 240 26623 240 26623 4 gnd
port 261 nsew
rlabel metal3 s 240 45583 240 45583 4 gnd
port 261 nsew
rlabel metal3 s 240 36577 240 36577 4 gnd
port 261 nsew
rlabel metal3 s 240 42107 240 42107 4 gnd
port 261 nsew
rlabel metal3 s 240 30020 240 30020 4 gnd
port 261 nsew
rlabel metal3 s 240 40527 240 40527 4 gnd
port 261 nsew
rlabel metal3 s 240 46847 240 46847 4 gnd
port 261 nsew
rlabel metal3 s 240 48743 240 48743 4 gnd
port 261 nsew
rlabel metal3 s 240 38473 240 38473 4 gnd
port 261 nsew
rlabel metal3 s 240 49217 240 49217 4 gnd
port 261 nsew
rlabel metal3 s 240 31837 240 31837 4 gnd
port 261 nsew
rlabel metal3 s 240 42660 240 42660 4 gnd
port 261 nsew
rlabel metal3 s 240 30810 240 30810 4 gnd
port 261 nsew
rlabel metal3 s 240 41317 240 41317 4 gnd
port 261 nsew
rlabel metal3 s 240 36340 240 36340 4 gnd
port 261 nsew
rlabel metal3 s 240 46057 240 46057 4 gnd
port 261 nsew
rlabel metal3 s 240 49770 240 49770 4 gnd
port 261 nsew
rlabel metal3 s 240 41633 240 41633 4 gnd
port 261 nsew
rlabel metal3 s 240 50323 240 50323 4 gnd
port 261 nsew
rlabel metal3 s 240 45820 240 45820 4 gnd
port 261 nsew
rlabel metal3 s 240 33733 240 33733 4 gnd
port 261 nsew
rlabel metal3 s 240 50560 240 50560 4 gnd
port 261 nsew
rlabel metal3 s 240 51587 240 51587 4 gnd
port 261 nsew
rlabel metal3 s 240 50797 240 50797 4 gnd
port 261 nsew
rlabel metal3 s 240 39737 240 39737 4 gnd
port 261 nsew
rlabel metal3 s 240 28440 240 28440 4 gnd
port 261 nsew
rlabel metal3 s 240 26860 240 26860 4 gnd
port 261 nsew
rlabel metal3 s 240 36893 240 36893 4 gnd
port 261 nsew
rlabel metal3 s 240 31363 240 31363 4 gnd
port 261 nsew
rlabel metal3 s 240 19987 240 19987 4 gnd
port 261 nsew
rlabel metal3 s 240 20540 240 20540 4 gnd
port 261 nsew
rlabel metal3 s 240 21883 240 21883 4 gnd
port 261 nsew
rlabel metal3 s 240 7663 240 7663 4 gnd
port 261 nsew
rlabel metal3 s 240 18407 240 18407 4 gnd
port 261 nsew
rlabel metal3 s 240 16037 240 16037 4 gnd
port 261 nsew
rlabel metal3 s 240 4740 240 4740 4 gnd
port 261 nsew
rlabel metal3 s 240 5530 240 5530 4 gnd
port 261 nsew
rlabel metal3 s 240 24727 240 24727 4 gnd
port 261 nsew
rlabel metal3 s 240 9717 240 9717 4 gnd
port 261 nsew
rlabel metal3 s 240 3397 240 3397 4 gnd
port 261 nsew
rlabel metal3 s 240 12640 240 12640 4 gnd
port 261 nsew
rlabel metal3 s 240 25043 240 25043 4 gnd
port 261 nsew
rlabel metal3 s 240 3713 240 3713 4 gnd
port 261 nsew
rlabel metal3 s 240 5767 240 5767 4 gnd
port 261 nsew
rlabel metal3 s 240 11297 240 11297 4 gnd
port 261 nsew
rlabel metal3 s 240 18170 240 18170 4 gnd
port 261 nsew
rlabel metal3 s 240 1817 240 1817 4 gnd
port 261 nsew
rlabel metal3 s 240 17143 240 17143 4 gnd
port 261 nsew
rlabel metal3 s 240 10823 240 10823 4 gnd
port 261 nsew
rlabel metal3 s 240 4187 240 4187 4 gnd
port 261 nsew
rlabel metal3 s 240 23937 240 23937 4 gnd
port 261 nsew
rlabel metal3 s 240 25833 240 25833 4 gnd
port 261 nsew
rlabel metal3 s 240 21330 240 21330 4 gnd
port 261 nsew
rlabel metal3 s 240 23147 240 23147 4 gnd
port 261 nsew
rlabel metal3 s 240 8927 240 8927 4 gnd
port 261 nsew
rlabel metal3 s 240 20777 240 20777 4 gnd
port 261 nsew
rlabel metal3 s 240 6873 240 6873 4 gnd
port 261 nsew
rlabel metal3 s 240 11613 240 11613 4 gnd
port 261 nsew
rlabel metal3 s 240 17380 240 17380 4 gnd
port 261 nsew
rlabel metal3 s 240 12877 240 12877 4 gnd
port 261 nsew
rlabel metal3 s 240 17617 240 17617 4 gnd
port 261 nsew
rlabel metal3 s 240 15800 240 15800 4 gnd
port 261 nsew
rlabel metal3 s 240 10270 240 10270 4 gnd
port 261 nsew
rlabel metal3 s 240 2607 240 2607 4 gnd
port 261 nsew
rlabel metal3 s 240 19750 240 19750 4 gnd
port 261 nsew
rlabel metal3 s 240 14773 240 14773 4 gnd
port 261 nsew
rlabel metal3 s 240 2133 240 2133 4 gnd
port 261 nsew
rlabel metal3 s 240 6320 240 6320 4 gnd
port 261 nsew
rlabel metal3 s 240 25280 240 25280 4 gnd
port 261 nsew
rlabel metal3 s 240 15563 240 15563 4 gnd
port 261 nsew
rlabel metal3 s 240 19513 240 19513 4 gnd
port 261 nsew
rlabel metal3 s 240 20303 240 20303 4 gnd
port 261 nsew
rlabel metal3 s 240 4503 240 4503 4 gnd
port 261 nsew
rlabel metal3 s 240 4977 240 4977 4 gnd
port 261 nsew
rlabel metal3 s 240 18723 240 18723 4 gnd
port 261 nsew
rlabel metal3 s 240 13667 240 13667 4 gnd
port 261 nsew
rlabel metal3 s 240 7900 240 7900 4 gnd
port 261 nsew
rlabel metal3 s 240 9480 240 9480 4 gnd
port 261 nsew
rlabel metal3 s 240 19197 240 19197 4 gnd
port 261 nsew
rlabel metal3 s 240 16353 240 16353 4 gnd
port 261 nsew
rlabel metal3 s 240 13193 240 13193 4 gnd
port 261 nsew
rlabel metal3 s 240 22910 240 22910 4 gnd
port 261 nsew
rlabel metal3 s 240 7110 240 7110 4 gnd
port 261 nsew
rlabel metal3 s 240 1580 240 1580 4 gnd
port 261 nsew
rlabel metal3 s 240 3950 240 3950 4 gnd
port 261 nsew
rlabel metal3 s 240 15010 240 15010 4 gnd
port 261 nsew
rlabel metal3 s 240 13983 240 13983 4 gnd
port 261 nsew
rlabel metal3 s 240 22673 240 22673 4 gnd
port 261 nsew
rlabel metal3 s 240 16827 240 16827 4 gnd
port 261 nsew
rlabel metal3 s 240 22120 240 22120 4 gnd
port 261 nsew
rlabel metal3 s 240 10507 240 10507 4 gnd
port 261 nsew
rlabel metal3 s 240 25517 240 25517 4 gnd
port 261 nsew
rlabel metal3 s 240 26070 240 26070 4 gnd
port 261 nsew
rlabel metal3 s 240 15247 240 15247 4 gnd
port 261 nsew
rlabel metal3 s 240 24490 240 24490 4 gnd
port 261 nsew
rlabel metal3 s 240 553 240 553 4 gnd
port 261 nsew
rlabel metal3 s 240 3160 240 3160 4 gnd
port 261 nsew
rlabel metal3 s 240 1343 240 1343 4 gnd
port 261 nsew
rlabel metal3 s 240 8453 240 8453 4 gnd
port 261 nsew
rlabel metal3 s 240 1027 240 1027 4 gnd
port 261 nsew
rlabel metal3 s 240 11060 240 11060 4 gnd
port 261 nsew
rlabel metal3 s 240 21567 240 21567 4 gnd
port 261 nsew
rlabel metal3 s 240 21093 240 21093 4 gnd
port 261 nsew
rlabel metal3 s 240 22357 240 22357 4 gnd
port 261 nsew
rlabel metal3 s 240 2370 240 2370 4 gnd
port 261 nsew
rlabel metal3 s 240 2923 240 2923 4 gnd
port 261 nsew
rlabel metal3 s 240 23700 240 23700 4 gnd
port 261 nsew
rlabel metal3 s 240 7347 240 7347 4 gnd
port 261 nsew
rlabel metal3 s 240 23463 240 23463 4 gnd
port 261 nsew
rlabel metal3 s 240 16590 240 16590 4 gnd
port 261 nsew
rlabel metal3 s 240 13430 240 13430 4 gnd
port 261 nsew
rlabel metal3 s 240 8137 240 8137 4 gnd
port 261 nsew
rlabel metal3 s 240 9243 240 9243 4 gnd
port 261 nsew
rlabel metal3 s 240 11850 240 11850 4 gnd
port 261 nsew
rlabel metal3 s 240 12087 240 12087 4 gnd
port 261 nsew
rlabel metal3 s 240 6083 240 6083 4 gnd
port 261 nsew
rlabel metal3 s 240 24253 240 24253 4 gnd
port 261 nsew
rlabel metal3 s 240 790 240 790 4 gnd
port 261 nsew
rlabel metal3 s 240 18960 240 18960 4 gnd
port 261 nsew
rlabel metal3 s 240 14220 240 14220 4 gnd
port 261 nsew
rlabel metal3 s 240 5293 240 5293 4 gnd
port 261 nsew
rlabel metal3 s 240 8690 240 8690 4 gnd
port 261 nsew
rlabel metal3 s 240 6557 240 6557 4 gnd
port 261 nsew
rlabel metal3 s 240 12403 240 12403 4 gnd
port 261 nsew
rlabel metal3 s 240 14457 240 14457 4 gnd
port 261 nsew
rlabel metal3 s 240 17933 240 17933 4 gnd
port 261 nsew
rlabel metal3 s 240 10033 240 10033 4 gnd
port 261 nsew
<< properties >>
string FIXED_BBOX 0 0 624 52140
string GDS_END 4577438
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4503342
<< end >>
