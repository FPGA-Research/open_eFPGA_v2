magic
tech sky130A
magscale 1 2
timestamp 1707688321
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_1
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 20771116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 20770190
<< end >>
