##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 18:34:03 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S_term_single2
  CLASS BLOCK ;
  SIZE 240.1200 BY 30.2600 ;
  FOREIGN S_term_single2 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.282 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.9450 29.9300 14.1150 30.2600 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.9672 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 69.7585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.956 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 12.5650 29.9300 12.7350 30.2600 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 29.9300 11.3550 30.2600 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.3508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.008 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 29.9300 10.4350 30.2600 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.7868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 83.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 29.9300 25.1550 30.2600 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.606 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 23.6050 29.9300 23.7750 30.2600 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.472 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.2250 29.9300 22.3950 30.2600 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.072 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 29.9300 21.0150 30.2600 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7433 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.9778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.4958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.448 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 29.9300 19.6350 30.2600 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.097 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3888 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.8295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.67 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.0850 29.9300 18.2550 30.2600 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.0902 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 29.9300 16.8750 30.2600 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.631 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 29.9300 15.4950 30.2600 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.002 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 29.9300 35.7350 30.2600 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 29.9300 34.3550 30.2600 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.322 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 29.9300 33.4350 30.2600 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.308 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 31.8850 29.9300 32.0550 30.2600 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8377 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.0175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.336 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 30.5050 29.9300 30.6750 30.2600 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4017 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8375 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.0868 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.6 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 29.9300 29.2950 30.2600 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.3964 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.205 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.944 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 27.7450 29.9300 27.9150 30.2600 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9389 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 28.51 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 152.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 26.3650 29.9300 26.5350 30.2600 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.99025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.165 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.7904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 73.8745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.714 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.1850 29.9300 57.3550 30.2600 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.5132 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.33 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 29.9300 56.4350 30.2600 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.828 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 59.0625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3694 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.048 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.8850 29.9300 55.0550 30.2600 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.572 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.408 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.5050 29.9300 53.6750 30.2600 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7621 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.888 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.424 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 29.9300 52.2950 30.2600 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.584 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.8425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.7450 29.9300 50.9150 30.2600 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27925 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.505 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.1845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8856 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.31 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 49.3650 29.9300 49.5350 30.2600 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.39485 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.641 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.2548 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 81.1965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.868 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 29.9300 48.1550 30.2600 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 46.6050 29.9300 46.7750 30.2600 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.428 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.416 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.2250 29.9300 45.3950 30.2600 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.808 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 29.9300 44.0150 30.2600 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0256 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.01 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.4650 29.9300 42.6350 30.2600 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 41.0850 29.9300 41.2550 30.2600 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 29.9300 39.8750 30.2600 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 40.3025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 38.3250 29.9300 38.4950 30.2600 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.144 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.6425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4311 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 36.9450 29.9300 37.1150 30.2600 ;
    END
  END N4BEG[0]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 29.9300 79.4350 30.2600 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.8850 29.9300 78.0550 30.2600 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.0992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.4185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 29.9300 76.6750 30.2600 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 29.9300 75.2950 30.2600 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.594 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.7450 29.9300 73.9150 30.2600 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.897 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 29.9300 72.5350 30.2600 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.676 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 29.9300 71.1550 30.2600 ;
    END
  END NN4BEG[9]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9396 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.614 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.6050 29.9300 69.7750 30.2600 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.282 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 68.2250 29.9300 68.3950 30.2600 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 29.9300 67.0150 30.2600 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0099 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.0828 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.912 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 65.4650 29.9300 65.6350 30.2600 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.2788 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 61.3165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 64.0850 29.9300 64.2550 30.2600 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 29.9300 62.8750 30.2600 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7088 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.426 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.3250 29.9300 61.4950 30.2600 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.4388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 104.144 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 59.9450 29.9300 60.1150 30.2600 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.29665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.349 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.3338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.315 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 29.9300 58.7350 30.2600 ;
    END
  END NN4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.52785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.621 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.314 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.5418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.2013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 84.3250 29.9300 84.4950 30.2600 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.274 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 29.1355 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 136.324 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 82.9450 29.9300 83.1150 30.2600 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6173 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9155 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.09 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.7046 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 77.2481 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 413.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 81.5650 29.9300 81.7350 30.2600 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2316 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.0805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.798 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.3066 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.5094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 80.1850 29.9300 80.3550 30.2600 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.5997 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.9748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 105.9450 29.9300 106.1150 30.2600 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.064 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2055 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.39 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 104.5650 29.9300 104.7350 30.2600 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.368 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9733 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.4182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 103.1850 29.9300 103.3550 30.2600 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.524 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.9277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 102.2650 29.9300 102.4350 30.2600 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.4865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.5692 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 100.8850 29.9300 101.0550 30.2600 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7945 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.825 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.1552 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.376 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 50.2934 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 268.808 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 99.5050 29.9300 99.6750 30.2600 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.98645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.337 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.62 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.5519 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.7642 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 98.1250 29.9300 98.2950 30.2600 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8126 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.956 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.9705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.8211 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.8522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 96.7450 29.9300 96.9150 30.2600 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2968 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5833 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.20245 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.0396 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.152 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 50.6167 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 269.509 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 95.3650 29.9300 95.5350 30.2600 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.2575 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 120.94 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 93.9850 29.9300 94.1550 30.2600 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.9048 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5599 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.1648 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 69.0632 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 366.918 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 92.6050 29.9300 92.7750 30.2600 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0424 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.094 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.3805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 91.2250 29.9300 91.3950 30.2600 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3128 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.4865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.108 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2123 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.0377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 89.8450 29.9300 90.0150 30.2600 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.0096 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.812 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.2638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.129 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 88.4650 29.9300 88.6350 30.2600 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.2262 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.541 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 40.5079 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 195.547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 87.0850 29.9300 87.2550 30.2600 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.536 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0827 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.1604 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 85.7050 29.9300 85.8750 30.2600 ;
    END
  END S2END[0]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.846 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8348 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.056 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.1104 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.104 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 149.1850 29.9300 149.3550 30.2600 ;
    END
  END SS4END[15]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.891 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.0412 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.698 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 148.2650 29.9300 148.4350 30.2600 ;
    END
  END SS4END[14]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.0442 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 36.4651 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 203.594 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 146.8850 29.9300 147.0550 30.2600 ;
    END
  END SS4END[13]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.0739 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 55.9214 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 145.5050 29.9300 145.6750 30.2600 ;
    END
  END SS4END[12]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.18405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.25629 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.8333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 144.1250 29.9300 144.2950 30.2600 ;
    END
  END SS4END[11]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.58 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.3318 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.1855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 142.7450 29.9300 142.9150 30.2600 ;
    END
  END SS4END[10]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4842 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6167 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.623 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 141.3650 29.9300 141.5350 30.2600 ;
    END
  END SS4END[9]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.44 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.082 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1984 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.544 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 139.9850 29.9300 140.1550 30.2600 ;
    END
  END SS4END[8]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4188 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.858 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6777 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.783 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 138.6050 29.9300 138.7750 30.2600 ;
    END
  END SS4END[7]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.95 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.9418 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.2704 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 137.2250 29.9300 137.3950 30.2600 ;
    END
  END SS4END[6]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.99 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.6475 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.374 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 135.8450 29.9300 136.0150 30.2600 ;
    END
  END SS4END[5]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3252 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.85 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.014 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.8299 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.9591 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 134.4650 29.9300 134.6350 30.2600 ;
    END
  END SS4END[4]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.301 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.584 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 59.8179 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 314.019 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 133.0850 29.9300 133.2550 30.2600 ;
    END
  END SS4END[3]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.572 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 82.5346 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 131.7050 29.9300 131.8750 30.2600 ;
    END
  END SS4END[2]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.168 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.6626 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.5472 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 130.3250 29.9300 130.4950 30.2600 ;
    END
  END SS4END[1]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.492625 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.088 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2376 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 91.6091 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 489.799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 128.9450 29.9300 129.1150 30.2600 ;
    END
  END SS4END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.814 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.834 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 27.006 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.84 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 127.5650 29.9300 127.7350 30.2600 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.78 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.9909 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.5314 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 126.1850 29.9300 126.3550 30.2600 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.01625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.725 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2398 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.081 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.4362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.1572 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 125.2650 29.9300 125.4350 30.2600 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.7404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.6245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.8585 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 123.8850 29.9300 124.0550 30.2600 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.17685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.561 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.68 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.928 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 44.728 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 216.965 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 122.5050 29.9300 122.6750 30.2600 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.51725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.785 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.238 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.4651 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 111.33 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 121.1250 29.9300 121.2950 30.2600 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.1632 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 81.3679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 119.7450 29.9300 119.9150 30.2600 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.16705 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.373 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.69 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.5682 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.3931 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 118.3650 29.9300 118.5350 30.2600 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.972 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7016 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 26.9588 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 146.453 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 116.9850 29.9300 117.1550 30.2600 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.038 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.977 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.9528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 115.6050 29.9300 115.7750 30.2600 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.568 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6515 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.1858 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 76.4811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 114.2250 29.9300 114.3950 30.2600 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.558 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.1898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.713 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 28.6613 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 138.116 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 112.8450 29.9300 113.0150 30.2600 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.3134 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.331 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.7959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 112.494 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 111.4650 29.9300 111.6350 30.2600 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.208 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 78.7814 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 110.0850 29.9300 110.2550 30.2600 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0564 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.0935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8115 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 55.184 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 291.126 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 108.7050 29.9300 108.8750 30.2600 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.76245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.897 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.584 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9204 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 74.4119 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 107.3250 29.9300 107.4950 30.2600 ;
    END
  END S4END[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9068 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.4565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.68 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.5179 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 102.082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0672 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.432 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.3436 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.6405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.5386 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.48 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 95.1475 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 512.67 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3576 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 60.0274 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 292.431 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6014 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.884 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.0356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 55.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.858 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.818 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3242 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.3711 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.808 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.9625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.842 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 31.7846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 153.415 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8822 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 12.958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.0656 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.624 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 21.4909 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 116.664 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.7076 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 63.4235 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.499 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.6022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 23.5629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6675 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.737 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 82.6456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 440.547 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.697 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.82 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5028 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.4365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.932 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.07642 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 15.6164 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5823 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.7405 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.673 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 116.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8196 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 40.6204 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 213.314 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2753 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.934 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 101.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.6212 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 64.511 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 350.233 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4688 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.728 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.4444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.1445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.94 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0009 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 65.9811 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.7476 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.869 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 71.9777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 383.726 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.72 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.5225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.228 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.904 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6513 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.491 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.42245 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.497 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.2588 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 66.2165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0362 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.9906 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.5464 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.6545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.202 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.2601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.8522 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.938 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 53.5796 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 256.965 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.1495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6638 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.1918 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6641 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.92 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.04 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.9696 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 54.0569 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 290.818 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.411 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.58836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.0806 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 38.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 51.7695 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 273.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 77.038 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 380.805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9008 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.5956 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 115.032 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 609.132 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.662 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.45881 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.1667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6097 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.8875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 38.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 203.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 31.1642 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 165.928 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.6188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 110.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 69.4582 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 354.415 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1897 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.946 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.5582 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.192 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 80.4531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 437.541 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1175 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2506 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.8082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.776 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.3645 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.4686 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.758 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 20.8113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5985 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.9236 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.0755 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 20.2528 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 64.5022 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 327.657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7626 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.587 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 28.6600 240.1200 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3219 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 26.6200 240.1200 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.821 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 30.2448 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 161.776 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 24.9200 240.1200 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4866 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.089 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 22.8800 240.1200 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.716 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 21.1800 240.1200 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4064 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.806 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 19.1400 240.1200 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6844 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.078 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 17.4400 240.1200 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.3699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.5055 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 15.7400 240.1200 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8575 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 34.7826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.448 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 13.7000 240.1200 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6579 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.0635 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 12.0000 240.1200 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.1462 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.623 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 10.3000 240.1200 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 29.0508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 155.408 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 8.2600 240.1200 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.3728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 135.792 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 6.5600 240.1200 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.44 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 4.5200 240.1200 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2585 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 2.8200 240.1200 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7914 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.731 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 239.6350 1.1200 240.1200 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.4988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 77.4165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.592 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5858 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.928 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 27.6250 240.1200 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.0439 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.142 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.072 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 25.9250 240.1200 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.2264 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 56.0175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2972 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.368 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 24.2250 240.1200 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.9836 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.8405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.278 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 22.5250 240.1200 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.5196 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.5205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.38 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 20.8250 240.1200 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 160.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.3986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 120.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 19.1250 240.1200 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0094 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.364 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 10.2344 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.135 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 17.4250 240.1200 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1049 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.0748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.536 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 15.7250 240.1200 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.0688 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 60.2665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 14.0250 240.1200 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.5096 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 47.4705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.1245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.957 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.904 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.0338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.984 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 12.3250 240.1200 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.275 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 14.9192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 74.5185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 10.6250 240.1200 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.4152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.9985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0434 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.863 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 8.9250 240.1200 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3672 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.432 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 15.8208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 79.0265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 7.2250 240.1200 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 18.6016 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 92.8935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 5.5250 240.1200 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 16.1827 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 80.836 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 3.8250 240.1200 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.36465 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.429 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 13.0992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 65.4185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 239.7900 2.1250 240.1200 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6615 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.2154 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.9497 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 149.6600 0.0000 149.8000 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.1701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.6604 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 144.1400 0.0000 144.2800 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4531 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8035 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 26.8028 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 122.987 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 139.0800 0.0000 139.2200 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6349 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9485 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.1022 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 105.384 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 133.5600 0.0000 133.7000 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8215 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.3931 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 128.5000 0.0000 128.6400 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.233 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.229 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 57.7789 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 306.95 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 123.4400 0.0000 123.5800 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9535 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7852 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.7736 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 117.4600 0.0000 117.6000 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4995 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.6142 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.3679 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 112.8600 0.0000 113.0000 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.4934 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.7642 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 107.3400 0.0000 107.4800 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3425 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.5849 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 102.2800 0.0000 102.4200 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.7462 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 69.1887 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6808 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 98.8616 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 0.0000 91.8400 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.30849 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.4151 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 0.0000 86.7800 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8277 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9125 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.6381 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 107.258 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 81.5800 0.0000 81.7200 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4739 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7895 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.1978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.06 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 76.0600 0.0000 76.2000 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4805 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.2544 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 100.827 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 71.0000 0.0000 71.1400 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9383 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4655 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2569 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.9465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 65.9400 0.0000 66.0800 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.239 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 60.4200 0.0000 60.5600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4155 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.0947 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.3459 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 55.3600 0.0000 55.5000 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2955 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.6557 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 83.1509 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 50.3000 0.0000 50.4400 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1484 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.581 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 128.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.8754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 209.9200 29.7750 210.0600 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3015 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3995 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 206.7000 29.7750 206.8400 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 203.9400 29.7750 204.0800 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3326 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.384 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7898 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.016 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 201.1800 29.7750 201.3200 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9947 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7475 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 198.4200 29.7750 198.5600 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.38 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 33.1458 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.248 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 195.2000 29.7750 195.3400 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7299 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5415 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 192.4400 29.7750 192.5800 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 189.6800 29.7750 189.8200 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.829 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.6866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 186.9200 29.7750 187.0600 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3963 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.7555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 184.1600 29.7750 184.3000 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8375 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9615 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 180.9400 29.7750 181.0800 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 178.1800 29.7750 178.3200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.6131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 175.4200 29.7750 175.5600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5095 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 172.6600 29.7750 172.8000 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.177 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.724 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.311 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 169.9000 29.7750 170.0400 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6035 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 166.6800 29.7750 166.8200 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 163.9200 29.7750 164.0600 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 161.1600 29.7750 161.3000 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.098 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.2005 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 158.4000 29.7750 158.5400 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.8527 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 155.6400 29.7750 155.7800 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 234.5600 6.0700 ;
        RECT 5.5600 23.0000 234.5600 25.0000 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 232.5600 15.0600 234.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 232.5600 9.6200 234.5600 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 232.5600 20.5000 234.5600 20.9800 ;
      LAYER met4 ;
        RECT 232.5600 4.0700 234.5600 25.0000 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 237.5600 3.0700 ;
        RECT 2.5600 26.0000 237.5600 28.0000 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 235.5600 6.9000 237.5600 7.3800 ;
        RECT 235.5600 12.3400 237.5600 12.8200 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 235.5600 17.7800 237.5600 18.2600 ;
      LAYER met4 ;
        RECT 235.5600 1.0700 237.5600 28.0000 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 149.5250 29.7600 240.1200 30.2600 ;
      RECT 148.6050 29.7600 149.0150 30.2600 ;
      RECT 147.2250 29.7600 148.0950 30.2600 ;
      RECT 145.8450 29.7600 146.7150 30.2600 ;
      RECT 144.4650 29.7600 145.3350 30.2600 ;
      RECT 143.0850 29.7600 143.9550 30.2600 ;
      RECT 141.7050 29.7600 142.5750 30.2600 ;
      RECT 140.3250 29.7600 141.1950 30.2600 ;
      RECT 138.9450 29.7600 139.8150 30.2600 ;
      RECT 137.5650 29.7600 138.4350 30.2600 ;
      RECT 136.1850 29.7600 137.0550 30.2600 ;
      RECT 134.8050 29.7600 135.6750 30.2600 ;
      RECT 133.4250 29.7600 134.2950 30.2600 ;
      RECT 132.0450 29.7600 132.9150 30.2600 ;
      RECT 130.6650 29.7600 131.5350 30.2600 ;
      RECT 129.2850 29.7600 130.1550 30.2600 ;
      RECT 127.9050 29.7600 128.7750 30.2600 ;
      RECT 126.5250 29.7600 127.3950 30.2600 ;
      RECT 125.6050 29.7600 126.0150 30.2600 ;
      RECT 124.2250 29.7600 125.0950 30.2600 ;
      RECT 122.8450 29.7600 123.7150 30.2600 ;
      RECT 121.4650 29.7600 122.3350 30.2600 ;
      RECT 120.0850 29.7600 120.9550 30.2600 ;
      RECT 118.7050 29.7600 119.5750 30.2600 ;
      RECT 117.3250 29.7600 118.1950 30.2600 ;
      RECT 115.9450 29.7600 116.8150 30.2600 ;
      RECT 114.5650 29.7600 115.4350 30.2600 ;
      RECT 113.1850 29.7600 114.0550 30.2600 ;
      RECT 111.8050 29.7600 112.6750 30.2600 ;
      RECT 110.4250 29.7600 111.2950 30.2600 ;
      RECT 109.0450 29.7600 109.9150 30.2600 ;
      RECT 107.6650 29.7600 108.5350 30.2600 ;
      RECT 106.2850 29.7600 107.1550 30.2600 ;
      RECT 104.9050 29.7600 105.7750 30.2600 ;
      RECT 103.5250 29.7600 104.3950 30.2600 ;
      RECT 102.6050 29.7600 103.0150 30.2600 ;
      RECT 101.2250 29.7600 102.0950 30.2600 ;
      RECT 99.8450 29.7600 100.7150 30.2600 ;
      RECT 98.4650 29.7600 99.3350 30.2600 ;
      RECT 97.0850 29.7600 97.9550 30.2600 ;
      RECT 95.7050 29.7600 96.5750 30.2600 ;
      RECT 94.3250 29.7600 95.1950 30.2600 ;
      RECT 92.9450 29.7600 93.8150 30.2600 ;
      RECT 91.5650 29.7600 92.4350 30.2600 ;
      RECT 90.1850 29.7600 91.0550 30.2600 ;
      RECT 88.8050 29.7600 89.6750 30.2600 ;
      RECT 87.4250 29.7600 88.2950 30.2600 ;
      RECT 86.0450 29.7600 86.9150 30.2600 ;
      RECT 84.6650 29.7600 85.5350 30.2600 ;
      RECT 83.2850 29.7600 84.1550 30.2600 ;
      RECT 81.9050 29.7600 82.7750 30.2600 ;
      RECT 80.5250 29.7600 81.3950 30.2600 ;
      RECT 79.6050 29.7600 80.0150 30.2600 ;
      RECT 78.2250 29.7600 79.0950 30.2600 ;
      RECT 76.8450 29.7600 77.7150 30.2600 ;
      RECT 75.4650 29.7600 76.3350 30.2600 ;
      RECT 74.0850 29.7600 74.9550 30.2600 ;
      RECT 72.7050 29.7600 73.5750 30.2600 ;
      RECT 71.3250 29.7600 72.1950 30.2600 ;
      RECT 69.9450 29.7600 70.8150 30.2600 ;
      RECT 68.5650 29.7600 69.4350 30.2600 ;
      RECT 67.1850 29.7600 68.0550 30.2600 ;
      RECT 65.8050 29.7600 66.6750 30.2600 ;
      RECT 64.4250 29.7600 65.2950 30.2600 ;
      RECT 63.0450 29.7600 63.9150 30.2600 ;
      RECT 61.6650 29.7600 62.5350 30.2600 ;
      RECT 60.2850 29.7600 61.1550 30.2600 ;
      RECT 58.9050 29.7600 59.7750 30.2600 ;
      RECT 57.5250 29.7600 58.3950 30.2600 ;
      RECT 56.6050 29.7600 57.0150 30.2600 ;
      RECT 55.2250 29.7600 56.0950 30.2600 ;
      RECT 53.8450 29.7600 54.7150 30.2600 ;
      RECT 52.4650 29.7600 53.3350 30.2600 ;
      RECT 51.0850 29.7600 51.9550 30.2600 ;
      RECT 49.7050 29.7600 50.5750 30.2600 ;
      RECT 48.3250 29.7600 49.1950 30.2600 ;
      RECT 46.9450 29.7600 47.8150 30.2600 ;
      RECT 45.5650 29.7600 46.4350 30.2600 ;
      RECT 44.1850 29.7600 45.0550 30.2600 ;
      RECT 42.8050 29.7600 43.6750 30.2600 ;
      RECT 41.4250 29.7600 42.2950 30.2600 ;
      RECT 40.0450 29.7600 40.9150 30.2600 ;
      RECT 38.6650 29.7600 39.5350 30.2600 ;
      RECT 37.2850 29.7600 38.1550 30.2600 ;
      RECT 35.9050 29.7600 36.7750 30.2600 ;
      RECT 34.5250 29.7600 35.3950 30.2600 ;
      RECT 33.6050 29.7600 34.0150 30.2600 ;
      RECT 32.2250 29.7600 33.0950 30.2600 ;
      RECT 30.8450 29.7600 31.7150 30.2600 ;
      RECT 29.4650 29.7600 30.3350 30.2600 ;
      RECT 28.0850 29.7600 28.9550 30.2600 ;
      RECT 26.7050 29.7600 27.5750 30.2600 ;
      RECT 25.3250 29.7600 26.1950 30.2600 ;
      RECT 23.9450 29.7600 24.8150 30.2600 ;
      RECT 22.5650 29.7600 23.4350 30.2600 ;
      RECT 21.1850 29.7600 22.0550 30.2600 ;
      RECT 19.8050 29.7600 20.6750 30.2600 ;
      RECT 18.4250 29.7600 19.2950 30.2600 ;
      RECT 17.0450 29.7600 17.9150 30.2600 ;
      RECT 15.6650 29.7600 16.5350 30.2600 ;
      RECT 14.2850 29.7600 15.1550 30.2600 ;
      RECT 12.9050 29.7600 13.7750 30.2600 ;
      RECT 11.5250 29.7600 12.3950 30.2600 ;
      RECT 10.6050 29.7600 11.0150 30.2600 ;
      RECT 0.0000 29.7600 10.0950 30.2600 ;
      RECT 0.0000 28.9850 240.1200 29.7600 ;
      RECT 0.5000 28.4750 240.1200 28.9850 ;
      RECT 0.0000 27.9650 240.1200 28.4750 ;
      RECT 0.0000 27.4550 239.6200 27.9650 ;
      RECT 0.0000 26.9450 240.1200 27.4550 ;
      RECT 0.5000 26.4350 240.1200 26.9450 ;
      RECT 0.0000 26.2650 240.1200 26.4350 ;
      RECT 0.0000 25.7550 239.6200 26.2650 ;
      RECT 0.0000 25.2450 240.1200 25.7550 ;
      RECT 0.5000 24.7350 240.1200 25.2450 ;
      RECT 0.0000 24.5650 240.1200 24.7350 ;
      RECT 0.0000 24.0550 239.6200 24.5650 ;
      RECT 0.0000 23.2050 240.1200 24.0550 ;
      RECT 0.5000 22.8650 240.1200 23.2050 ;
      RECT 0.5000 22.6950 239.6200 22.8650 ;
      RECT 0.0000 22.3550 239.6200 22.6950 ;
      RECT 0.0000 21.5050 240.1200 22.3550 ;
      RECT 0.5000 21.1650 240.1200 21.5050 ;
      RECT 0.5000 20.9950 239.6200 21.1650 ;
      RECT 0.0000 20.6550 239.6200 20.9950 ;
      RECT 0.0000 19.4650 240.1200 20.6550 ;
      RECT 0.5000 18.9550 239.6200 19.4650 ;
      RECT 0.0000 17.7650 240.1200 18.9550 ;
      RECT 0.5000 17.2550 239.6200 17.7650 ;
      RECT 0.0000 16.0650 240.1200 17.2550 ;
      RECT 0.5000 15.5550 239.6200 16.0650 ;
      RECT 0.0000 14.3650 240.1200 15.5550 ;
      RECT 0.0000 14.0250 239.6200 14.3650 ;
      RECT 0.5000 13.8550 239.6200 14.0250 ;
      RECT 0.5000 13.5150 240.1200 13.8550 ;
      RECT 0.0000 12.6650 240.1200 13.5150 ;
      RECT 0.0000 12.3250 239.6200 12.6650 ;
      RECT 0.5000 12.1550 239.6200 12.3250 ;
      RECT 0.5000 11.8150 240.1200 12.1550 ;
      RECT 0.0000 10.9650 240.1200 11.8150 ;
      RECT 0.0000 10.6250 239.6200 10.9650 ;
      RECT 0.5000 10.4550 239.6200 10.6250 ;
      RECT 0.5000 10.1150 240.1200 10.4550 ;
      RECT 0.0000 9.2650 240.1200 10.1150 ;
      RECT 0.0000 8.7550 239.6200 9.2650 ;
      RECT 0.0000 8.5850 240.1200 8.7550 ;
      RECT 0.5000 8.0750 240.1200 8.5850 ;
      RECT 0.0000 7.5650 240.1200 8.0750 ;
      RECT 0.0000 7.0550 239.6200 7.5650 ;
      RECT 0.0000 6.8850 240.1200 7.0550 ;
      RECT 0.5000 6.3750 240.1200 6.8850 ;
      RECT 0.0000 5.8650 240.1200 6.3750 ;
      RECT 0.0000 5.3550 239.6200 5.8650 ;
      RECT 0.0000 4.8450 240.1200 5.3550 ;
      RECT 0.5000 4.3350 240.1200 4.8450 ;
      RECT 0.0000 4.1650 240.1200 4.3350 ;
      RECT 0.0000 3.6550 239.6200 4.1650 ;
      RECT 0.0000 3.1450 240.1200 3.6550 ;
      RECT 0.5000 2.6350 240.1200 3.1450 ;
      RECT 0.0000 2.4650 240.1200 2.6350 ;
      RECT 0.0000 1.9550 239.6200 2.4650 ;
      RECT 0.0000 1.4450 240.1200 1.9550 ;
      RECT 0.5000 0.9350 240.1200 1.4450 ;
      RECT 0.0000 0.0000 240.1200 0.9350 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 240.1200 30.2600 ;
    LAYER met2 ;
      RECT 210.2000 29.6350 240.1200 30.2600 ;
      RECT 206.9800 29.6350 209.7800 30.2600 ;
      RECT 204.2200 29.6350 206.5600 30.2600 ;
      RECT 201.4600 29.6350 203.8000 30.2600 ;
      RECT 198.7000 29.6350 201.0400 30.2600 ;
      RECT 195.4800 29.6350 198.2800 30.2600 ;
      RECT 192.7200 29.6350 195.0600 30.2600 ;
      RECT 189.9600 29.6350 192.3000 30.2600 ;
      RECT 187.2000 29.6350 189.5400 30.2600 ;
      RECT 184.4400 29.6350 186.7800 30.2600 ;
      RECT 181.2200 29.6350 184.0200 30.2600 ;
      RECT 178.4600 29.6350 180.8000 30.2600 ;
      RECT 175.7000 29.6350 178.0400 30.2600 ;
      RECT 172.9400 29.6350 175.2800 30.2600 ;
      RECT 170.1800 29.6350 172.5200 30.2600 ;
      RECT 166.9600 29.6350 169.7600 30.2600 ;
      RECT 164.2000 29.6350 166.5400 30.2600 ;
      RECT 161.4400 29.6350 163.7800 30.2600 ;
      RECT 158.6800 29.6350 161.0200 30.2600 ;
      RECT 155.9200 29.6350 158.2600 30.2600 ;
      RECT 0.0000 29.6350 155.5000 30.2600 ;
      RECT 0.0000 28.9400 240.1200 29.6350 ;
      RECT 0.0000 28.5200 239.4950 28.9400 ;
      RECT 0.0000 27.9200 240.1200 28.5200 ;
      RECT 0.6250 27.5000 240.1200 27.9200 ;
      RECT 0.0000 26.9000 240.1200 27.5000 ;
      RECT 0.0000 26.4800 239.4950 26.9000 ;
      RECT 0.0000 26.2200 240.1200 26.4800 ;
      RECT 0.6250 25.8000 240.1200 26.2200 ;
      RECT 0.0000 25.2000 240.1200 25.8000 ;
      RECT 0.0000 24.7800 239.4950 25.2000 ;
      RECT 0.0000 24.5200 240.1200 24.7800 ;
      RECT 0.6250 24.1000 240.1200 24.5200 ;
      RECT 0.0000 23.1600 240.1200 24.1000 ;
      RECT 0.0000 22.8200 239.4950 23.1600 ;
      RECT 0.6250 22.7400 239.4950 22.8200 ;
      RECT 0.6250 22.4000 240.1200 22.7400 ;
      RECT 0.0000 21.4600 240.1200 22.4000 ;
      RECT 0.0000 21.1200 239.4950 21.4600 ;
      RECT 0.6250 21.0400 239.4950 21.1200 ;
      RECT 0.6250 20.7000 240.1200 21.0400 ;
      RECT 0.0000 19.4200 240.1200 20.7000 ;
      RECT 0.6250 19.0000 239.4950 19.4200 ;
      RECT 0.0000 17.7200 240.1200 19.0000 ;
      RECT 0.6250 17.3000 239.4950 17.7200 ;
      RECT 0.0000 16.0200 240.1200 17.3000 ;
      RECT 0.6250 15.6000 239.4950 16.0200 ;
      RECT 0.0000 14.3200 240.1200 15.6000 ;
      RECT 0.6250 13.9800 240.1200 14.3200 ;
      RECT 0.6250 13.9000 239.4950 13.9800 ;
      RECT 0.0000 13.5600 239.4950 13.9000 ;
      RECT 0.0000 12.6200 240.1200 13.5600 ;
      RECT 0.6250 12.2800 240.1200 12.6200 ;
      RECT 0.6250 12.2000 239.4950 12.2800 ;
      RECT 0.0000 11.8600 239.4950 12.2000 ;
      RECT 0.0000 10.9200 240.1200 11.8600 ;
      RECT 0.6250 10.5800 240.1200 10.9200 ;
      RECT 0.6250 10.5000 239.4950 10.5800 ;
      RECT 0.0000 10.1600 239.4950 10.5000 ;
      RECT 0.0000 9.2200 240.1200 10.1600 ;
      RECT 0.6250 8.8000 240.1200 9.2200 ;
      RECT 0.0000 8.5400 240.1200 8.8000 ;
      RECT 0.0000 8.1200 239.4950 8.5400 ;
      RECT 0.0000 7.5200 240.1200 8.1200 ;
      RECT 0.6250 7.1000 240.1200 7.5200 ;
      RECT 0.0000 6.8400 240.1200 7.1000 ;
      RECT 0.0000 6.4200 239.4950 6.8400 ;
      RECT 0.0000 5.8200 240.1200 6.4200 ;
      RECT 0.6250 5.4000 240.1200 5.8200 ;
      RECT 0.0000 4.8000 240.1200 5.4000 ;
      RECT 0.0000 4.3800 239.4950 4.8000 ;
      RECT 0.0000 4.1200 240.1200 4.3800 ;
      RECT 0.6250 3.7000 240.1200 4.1200 ;
      RECT 0.0000 3.1000 240.1200 3.7000 ;
      RECT 0.0000 2.6800 239.4950 3.1000 ;
      RECT 0.0000 2.4200 240.1200 2.6800 ;
      RECT 0.6250 2.0000 240.1200 2.4200 ;
      RECT 0.0000 1.4000 240.1200 2.0000 ;
      RECT 0.0000 0.9800 239.4950 1.4000 ;
      RECT 0.0000 0.6250 240.1200 0.9800 ;
      RECT 149.9400 0.0000 240.1200 0.6250 ;
      RECT 144.4200 0.0000 149.5200 0.6250 ;
      RECT 139.3600 0.0000 144.0000 0.6250 ;
      RECT 133.8400 0.0000 138.9400 0.6250 ;
      RECT 128.7800 0.0000 133.4200 0.6250 ;
      RECT 123.7200 0.0000 128.3600 0.6250 ;
      RECT 117.7400 0.0000 123.3000 0.6250 ;
      RECT 113.1400 0.0000 117.3200 0.6250 ;
      RECT 107.6200 0.0000 112.7200 0.6250 ;
      RECT 102.5600 0.0000 107.2000 0.6250 ;
      RECT 97.0400 0.0000 102.1400 0.6250 ;
      RECT 91.9800 0.0000 96.6200 0.6250 ;
      RECT 86.9200 0.0000 91.5600 0.6250 ;
      RECT 81.8600 0.0000 86.5000 0.6250 ;
      RECT 76.3400 0.0000 81.4400 0.6250 ;
      RECT 71.2800 0.0000 75.9200 0.6250 ;
      RECT 66.2200 0.0000 70.8600 0.6250 ;
      RECT 60.7000 0.0000 65.8000 0.6250 ;
      RECT 55.6400 0.0000 60.2800 0.6250 ;
      RECT 50.5800 0.0000 55.2200 0.6250 ;
      RECT 0.0000 0.0000 50.1600 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 237.8600 25.7000 240.1200 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 240.1200 25.7000 ;
      RECT 234.8600 22.7000 240.1200 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 240.1200 22.7000 ;
      RECT 234.8600 20.2000 240.1200 21.2800 ;
      RECT 7.8600 20.2000 232.2600 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 240.1200 20.2000 ;
      RECT 237.8600 17.4800 240.1200 18.5600 ;
      RECT 4.8600 17.4800 235.2600 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 240.1200 17.4800 ;
      RECT 234.8600 14.7600 240.1200 15.8400 ;
      RECT 7.8600 14.7600 232.2600 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 240.1200 14.7600 ;
      RECT 237.8600 12.0400 240.1200 13.1200 ;
      RECT 4.8600 12.0400 235.2600 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 240.1200 12.0400 ;
      RECT 234.8600 9.3200 240.1200 10.4000 ;
      RECT 7.8600 9.3200 232.2600 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 240.1200 9.3200 ;
      RECT 237.8600 6.6000 240.1200 7.6800 ;
      RECT 4.8600 6.6000 235.2600 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 240.1200 6.6000 ;
      RECT 234.8600 3.7700 240.1200 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 240.1200 3.7700 ;
      RECT 237.8600 0.7700 240.1200 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 240.1200 30.2600 ;
      RECT 4.8600 25.3000 235.2600 28.3000 ;
      RECT 234.8600 3.7700 235.2600 25.3000 ;
      RECT 7.8600 3.7700 232.2600 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 237.8600 0.7700 240.1200 28.3000 ;
      RECT 4.8600 0.7700 235.2600 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 240.1200 0.7700 ;
  END
END S_term_single2

END LIBRARY
