magic
tech sky130B
timestamp 1707688321
<< obsli1 >>
rect 0 396 394 413
rect 0 343 27 396
rect 411 378 438 413
rect 44 361 438 378
rect 0 326 394 343
rect 0 273 27 326
rect 411 308 438 361
rect 44 291 438 308
rect 0 256 394 273
rect 0 203 27 256
rect 411 238 438 291
rect 44 221 438 238
rect 0 186 394 203
rect 0 133 27 186
rect 411 168 438 221
rect 44 151 438 168
rect 0 116 394 133
rect 0 63 27 116
rect 411 98 438 151
rect 44 81 438 98
rect 0 46 394 63
rect 411 46 438 81
rect 0 32 27 46
<< obsm1 >>
rect 0 427 438 459
rect 0 32 27 413
rect 44 32 58 413
rect 72 46 86 427
rect 100 32 114 413
rect 128 46 142 427
rect 156 32 170 413
rect 184 46 198 427
rect 212 32 226 413
rect 240 46 254 427
rect 268 32 282 413
rect 296 46 310 427
rect 324 32 338 413
rect 352 46 366 427
rect 380 32 394 413
rect 411 46 438 427
rect 0 0 438 32
<< obsm2 >>
rect 0 427 438 459
rect 0 32 27 413
rect 44 46 58 427
rect 72 32 86 413
rect 100 46 114 427
rect 128 32 142 413
rect 156 46 170 427
rect 184 32 198 413
rect 212 46 226 427
rect 240 32 254 413
rect 268 46 282 427
rect 296 32 310 413
rect 324 46 338 427
rect 352 32 366 413
rect 380 46 394 427
rect 411 46 438 427
rect 0 0 438 32
<< properties >>
string FIXED_BBOX 0 0 438 459
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 70294
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 60000
<< end >>
