magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 35896 -598 35946 -582
rect 35930 -632 35946 -598
rect 35896 -648 35946 -632
<< polycont >>
rect -34 16 0 50
rect 35896 -632 35930 -598
<< npolyres >>
rect 0 0 35946 66
rect 35880 -96 35946 0
rect -50 -162 35946 -96
rect -50 -258 16 -162
rect -50 -324 35946 -258
rect 35880 -420 35946 -324
rect -50 -486 35946 -420
rect -50 -582 16 -486
rect -50 -648 35896 -582
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 35896 -598 35930 -582
rect 35896 -648 35930 -632
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_0
timestamp 1707688321
transform 1 0 -50 0 1 0
box 0 0 1 1
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_1
timestamp 1707688321
transform 1 0 35880 0 1 -648
box 0 0 1 1
<< properties >>
string GDS_END 42930456
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42928884
<< end >>
