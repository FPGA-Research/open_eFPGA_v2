magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1451 203
rect 29 -17 63 21
<< locali >>
rect 787 323 837 425
rect 955 323 1005 425
rect 1123 323 1173 425
rect 1291 323 1341 425
rect 787 289 1455 323
rect 72 215 706 255
rect 760 215 1308 255
rect 1342 181 1455 289
rect 107 145 1455 181
rect 107 51 173 145
rect 275 51 341 145
rect 443 51 509 145
rect 611 51 677 145
rect 779 51 845 145
rect 947 51 1013 145
rect 1115 51 1181 145
rect 1283 51 1349 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 18 333 81 493
rect 115 367 165 527
rect 199 333 249 493
rect 283 367 333 527
rect 367 333 417 493
rect 451 367 501 527
rect 535 333 585 493
rect 619 367 669 527
rect 703 459 1425 493
rect 703 333 753 459
rect 18 291 753 333
rect 871 357 921 459
rect 1039 357 1089 459
rect 1207 357 1257 459
rect 1375 357 1425 459
rect 18 17 73 181
rect 207 17 241 111
rect 375 17 409 111
rect 543 17 577 111
rect 711 17 745 111
rect 879 17 913 111
rect 1047 17 1081 111
rect 1215 17 1249 111
rect 1383 17 1441 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 72 215 706 255 6 A
port 1 nsew signal input
rlabel locali s 760 215 1308 255 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1451 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1283 51 1349 145 6 Y
port 7 nsew signal output
rlabel locali s 1115 51 1181 145 6 Y
port 7 nsew signal output
rlabel locali s 947 51 1013 145 6 Y
port 7 nsew signal output
rlabel locali s 779 51 845 145 6 Y
port 7 nsew signal output
rlabel locali s 611 51 677 145 6 Y
port 7 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 7 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 7 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 7 nsew signal output
rlabel locali s 107 145 1455 181 6 Y
port 7 nsew signal output
rlabel locali s 1342 181 1455 289 6 Y
port 7 nsew signal output
rlabel locali s 787 289 1455 323 6 Y
port 7 nsew signal output
rlabel locali s 1291 323 1341 425 6 Y
port 7 nsew signal output
rlabel locali s 1123 323 1173 425 6 Y
port 7 nsew signal output
rlabel locali s 955 323 1005 425 6 Y
port 7 nsew signal output
rlabel locali s 787 323 837 425 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1976198
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1964800
<< end >>
