magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 538
rect 61 0 64 538
<< via1 >>
rect 3 0 61 538
<< metal2 >>
rect 0 0 3 538
rect 61 0 64 538
<< properties >>
string GDS_END 88151118
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88148810
<< end >>
