magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 10046 9692 10777 13218
rect 10193 8170 10245 8202
<< pwell >>
rect 11269 13766 11491 14904
rect 11092 13544 11491 13766
rect 10186 9832 10272 12934
<< mvpsubdiff >>
rect 11295 14854 11465 14878
rect 11329 14820 11363 14854
rect 11397 14820 11431 14854
rect 11295 14785 11465 14820
rect 11329 14751 11363 14785
rect 11397 14783 11465 14785
rect 11397 14751 11431 14783
rect 11295 14749 11431 14751
rect 11295 14716 11465 14749
rect 11329 14682 11363 14716
rect 11397 14712 11465 14716
rect 11397 14682 11431 14712
rect 11295 14678 11431 14682
rect 11295 14647 11465 14678
rect 11329 14613 11363 14647
rect 11397 14641 11465 14647
rect 11397 14613 11431 14641
rect 11295 14607 11431 14613
rect 11295 14578 11465 14607
rect 11329 14544 11363 14578
rect 11397 14570 11465 14578
rect 11397 14544 11431 14570
rect 11295 14536 11431 14544
rect 11295 14509 11465 14536
rect 11329 14475 11363 14509
rect 11397 14499 11465 14509
rect 11397 14475 11431 14499
rect 11295 14465 11431 14475
rect 11295 14440 11465 14465
rect 11329 14406 11363 14440
rect 11397 14428 11465 14440
rect 11397 14406 11431 14428
rect 11295 14394 11431 14406
rect 11295 14371 11465 14394
rect 11295 14370 11363 14371
rect 11329 14337 11363 14370
rect 11397 14357 11465 14371
rect 11397 14337 11431 14357
rect 11329 14336 11431 14337
rect 11295 14323 11431 14336
rect 11295 14302 11465 14323
rect 11295 14300 11363 14302
rect 11329 14268 11363 14300
rect 11397 14286 11465 14302
rect 11397 14268 11431 14286
rect 11329 14266 11431 14268
rect 11295 14252 11431 14266
rect 11295 14232 11465 14252
rect 11295 14230 11363 14232
rect 11329 14198 11363 14230
rect 11397 14214 11465 14232
rect 11397 14198 11431 14214
rect 11329 14196 11431 14198
rect 11295 14180 11431 14196
rect 11295 14162 11465 14180
rect 11295 14160 11363 14162
rect 11329 14128 11363 14160
rect 11397 14142 11465 14162
rect 11397 14128 11431 14142
rect 11329 14126 11431 14128
rect 11295 14108 11431 14126
rect 11295 14092 11465 14108
rect 11295 14090 11363 14092
rect 11329 14058 11363 14090
rect 11397 14070 11465 14092
rect 11397 14058 11431 14070
rect 11329 14056 11431 14058
rect 11295 14036 11431 14056
rect 11295 14022 11465 14036
rect 11295 14020 11363 14022
rect 11329 13988 11363 14020
rect 11397 13998 11465 14022
rect 11397 13988 11431 13998
rect 11329 13986 11431 13988
rect 11295 13964 11431 13986
rect 11295 13952 11465 13964
rect 11295 13950 11363 13952
rect 11329 13918 11363 13950
rect 11397 13926 11465 13952
rect 11397 13918 11431 13926
rect 11329 13916 11431 13918
rect 11295 13892 11431 13916
rect 11295 13882 11465 13892
rect 11295 13880 11363 13882
rect 11329 13848 11363 13880
rect 11397 13854 11465 13882
rect 11397 13848 11431 13854
rect 11329 13846 11431 13848
rect 11295 13820 11431 13846
rect 11295 13812 11465 13820
rect 11295 13810 11363 13812
rect 11329 13778 11363 13810
rect 11397 13782 11465 13812
rect 11397 13778 11431 13782
rect 11329 13776 11431 13778
rect 11295 13748 11431 13776
rect 11295 13742 11465 13748
rect 11295 13740 11363 13742
rect 11118 13706 11142 13740
rect 11176 13706 11219 13740
rect 11253 13706 11295 13740
rect 11329 13708 11363 13740
rect 11397 13710 11465 13742
rect 11397 13708 11431 13710
rect 11329 13706 11431 13708
rect 11118 13676 11431 13706
rect 11118 13672 11465 13676
rect 11118 13638 11142 13672
rect 11176 13638 11216 13672
rect 11250 13638 11290 13672
rect 11324 13638 11363 13672
rect 11397 13638 11465 13672
rect 11118 13604 11431 13638
rect 11118 13570 11142 13604
rect 11176 13570 11223 13604
rect 11257 13570 11304 13604
rect 11338 13570 11465 13604
rect 10212 12884 10246 12908
rect 10212 9916 10246 12850
rect 10212 9858 10246 9882
<< mvpsubdiffcont >>
rect 11295 14820 11329 14854
rect 11363 14820 11397 14854
rect 11431 14820 11465 14854
rect 11295 14751 11329 14785
rect 11363 14751 11397 14785
rect 11431 14749 11465 14783
rect 11295 14682 11329 14716
rect 11363 14682 11397 14716
rect 11431 14678 11465 14712
rect 11295 14613 11329 14647
rect 11363 14613 11397 14647
rect 11431 14607 11465 14641
rect 11295 14544 11329 14578
rect 11363 14544 11397 14578
rect 11431 14536 11465 14570
rect 11295 14475 11329 14509
rect 11363 14475 11397 14509
rect 11431 14465 11465 14499
rect 11295 14406 11329 14440
rect 11363 14406 11397 14440
rect 11431 14394 11465 14428
rect 11295 14336 11329 14370
rect 11363 14337 11397 14371
rect 11431 14323 11465 14357
rect 11295 14266 11329 14300
rect 11363 14268 11397 14302
rect 11431 14252 11465 14286
rect 11295 14196 11329 14230
rect 11363 14198 11397 14232
rect 11431 14180 11465 14214
rect 11295 14126 11329 14160
rect 11363 14128 11397 14162
rect 11431 14108 11465 14142
rect 11295 14056 11329 14090
rect 11363 14058 11397 14092
rect 11431 14036 11465 14070
rect 11295 13986 11329 14020
rect 11363 13988 11397 14022
rect 11431 13964 11465 13998
rect 11295 13916 11329 13950
rect 11363 13918 11397 13952
rect 11431 13892 11465 13926
rect 11295 13846 11329 13880
rect 11363 13848 11397 13882
rect 11431 13820 11465 13854
rect 11295 13776 11329 13810
rect 11363 13778 11397 13812
rect 11431 13748 11465 13782
rect 11142 13706 11176 13740
rect 11219 13706 11253 13740
rect 11295 13706 11329 13740
rect 11363 13708 11397 13742
rect 11431 13676 11465 13710
rect 11142 13638 11176 13672
rect 11216 13638 11250 13672
rect 11290 13638 11324 13672
rect 11363 13638 11397 13672
rect 11431 13604 11465 13638
rect 11142 13570 11176 13604
rect 11223 13570 11257 13604
rect 11304 13570 11338 13604
rect 10212 12850 10246 12884
rect 10212 9882 10246 9916
<< poly >>
rect 10983 15574 11055 15590
rect 10983 15540 11005 15574
rect 11039 15540 11055 15574
rect 10983 15503 11055 15540
rect 10983 15470 11005 15503
rect 10989 15469 11005 15470
rect 11039 15469 11055 15503
rect 10989 15432 11055 15469
rect 10989 15414 11005 15432
rect 10983 15398 11005 15414
rect 11039 15398 11055 15432
rect 10983 15361 11055 15398
rect 10983 15327 11005 15361
rect 11039 15327 11055 15361
rect 10983 15294 11055 15327
rect 10989 15290 11055 15294
rect 10989 15256 11005 15290
rect 11039 15256 11055 15290
rect 10989 15238 11055 15256
rect 10983 15219 11055 15238
rect 10983 15185 11005 15219
rect 11039 15185 11055 15219
rect 10983 15148 11055 15185
rect 10983 15118 11005 15148
rect 10989 15114 11005 15118
rect 11039 15114 11055 15148
rect 10989 15077 11055 15114
rect 10989 15062 11005 15077
rect 10983 15043 11005 15062
rect 11039 15043 11055 15077
rect 10983 15006 11055 15043
rect 10983 14972 11005 15006
rect 11039 14972 11055 15006
rect 10983 14942 11055 14972
rect 10989 14935 11055 14942
rect 10989 14901 11005 14935
rect 11039 14901 11055 14935
rect 10989 14886 11055 14901
rect 10983 14864 11055 14886
rect 10983 14830 11005 14864
rect 11039 14830 11055 14864
rect 10983 14792 11055 14830
rect 10983 14766 11005 14792
rect 10989 14758 11005 14766
rect 11039 14758 11055 14792
rect 10989 14720 11055 14758
rect 10989 14710 11005 14720
rect 10983 14686 11005 14710
rect 11039 14686 11055 14720
rect 10983 14648 11055 14686
rect 10983 14614 11005 14648
rect 11039 14614 11055 14648
rect 10983 14590 11055 14614
rect 10989 14576 11055 14590
rect 10989 14542 11005 14576
rect 11039 14542 11055 14576
rect 10989 14534 11055 14542
rect 10983 14504 11055 14534
rect 10983 14470 11005 14504
rect 11039 14470 11055 14504
rect 10983 14432 11055 14470
rect 10983 14414 11005 14432
rect 10989 14398 11005 14414
rect 11039 14398 11055 14432
rect 10989 14360 11055 14398
rect 10989 14358 11005 14360
rect 10983 14326 11005 14358
rect 11039 14326 11055 14360
rect 10983 14288 11055 14326
rect 10983 14254 11005 14288
rect 11039 14254 11055 14288
rect 10983 14238 11055 14254
rect 10989 14182 11055 14196
rect 10983 14180 11055 14182
rect 10983 14146 11005 14180
rect 11039 14146 11055 14180
rect 10983 14112 11055 14146
rect 10983 14078 11005 14112
rect 11039 14078 11055 14112
rect 10983 14062 11055 14078
rect 10370 12823 10504 12839
rect 10370 12789 10386 12823
rect 10420 12789 10454 12823
rect 10488 12789 10504 12823
rect 10370 12773 10504 12789
rect 10373 12766 10493 12773
<< polycont >>
rect 11005 15540 11039 15574
rect 11005 15469 11039 15503
rect 11005 15398 11039 15432
rect 11005 15327 11039 15361
rect 11005 15256 11039 15290
rect 11005 15185 11039 15219
rect 11005 15114 11039 15148
rect 11005 15043 11039 15077
rect 11005 14972 11039 15006
rect 11005 14901 11039 14935
rect 11005 14830 11039 14864
rect 11005 14758 11039 14792
rect 11005 14686 11039 14720
rect 11005 14614 11039 14648
rect 11005 14542 11039 14576
rect 11005 14470 11039 14504
rect 11005 14398 11039 14432
rect 11005 14326 11039 14360
rect 11005 14254 11039 14288
rect 11005 14146 11039 14180
rect 11005 14078 11039 14112
rect 10386 12789 10420 12823
rect 10454 12789 10488 12823
<< locali >>
rect 10314 15601 10354 15635
rect 10388 15601 10428 15635
rect 10462 15601 10502 15635
rect 10536 15601 10576 15635
rect 10610 15601 10650 15635
rect 10684 15601 10723 15635
rect 10757 15601 10796 15635
rect 10830 15601 10869 15635
rect 11037 15574 11039 15590
rect 11003 15540 11005 15556
rect 11003 15517 11039 15540
rect 11037 15503 11039 15517
rect 11003 15469 11005 15483
rect 9983 15425 10024 15459
rect 10058 15425 10099 15459
rect 10133 15425 10174 15459
rect 10208 15425 10249 15459
rect 10283 15425 10323 15459
rect 10357 15425 10397 15459
rect 10431 15425 10471 15459
rect 11003 15444 11039 15469
rect 11037 15432 11039 15444
rect 11003 15398 11005 15410
rect 11003 15371 11039 15398
rect 11037 15361 11039 15371
rect 11003 15327 11005 15337
rect 11003 15298 11039 15327
rect 11037 15290 11039 15298
rect 10314 15249 10354 15283
rect 10388 15249 10428 15283
rect 10462 15249 10502 15283
rect 10536 15249 10576 15283
rect 10610 15249 10650 15283
rect 10684 15249 10723 15283
rect 10757 15249 10796 15283
rect 10830 15249 10869 15283
rect 11003 15256 11005 15264
rect 11003 15225 11039 15256
rect 11037 15219 11039 15225
rect 11003 15185 11005 15191
rect 11003 15152 11039 15185
rect 11037 15148 11039 15152
rect 11003 15114 11005 15118
rect 9983 15073 10024 15107
rect 10058 15073 10099 15107
rect 10133 15073 10174 15107
rect 10208 15073 10249 15107
rect 10283 15073 10323 15107
rect 10357 15073 10397 15107
rect 10431 15073 10471 15107
rect 11003 15079 11039 15114
rect 11037 15077 11039 15079
rect 11003 15043 11005 15045
rect 11003 15006 11039 15043
rect 11003 14935 11039 14972
rect 11003 14933 11005 14935
rect 10314 14897 10354 14931
rect 10388 14897 10428 14931
rect 10462 14897 10502 14931
rect 10536 14897 10576 14931
rect 10610 14897 10650 14931
rect 10684 14897 10723 14931
rect 10757 14897 10796 14931
rect 10830 14897 10869 14931
rect 11037 14899 11039 14901
rect 11003 14864 11039 14899
rect 11003 14860 11005 14864
rect 11037 14826 11039 14830
rect 11003 14792 11039 14826
rect 11003 14788 11005 14792
rect 9983 14721 10024 14755
rect 10058 14721 10099 14755
rect 10133 14721 10174 14755
rect 10208 14721 10249 14755
rect 10283 14721 10323 14755
rect 10357 14721 10397 14755
rect 10431 14721 10471 14755
rect 11037 14754 11039 14758
rect 11003 14720 11039 14754
rect 11003 14716 11005 14720
rect 11037 14682 11039 14686
rect 11003 14648 11039 14682
rect 11003 14644 11005 14648
rect 11037 14610 11039 14614
rect 10314 14545 10354 14579
rect 10388 14545 10428 14579
rect 10462 14545 10502 14579
rect 10536 14545 10576 14579
rect 10610 14545 10650 14579
rect 10684 14545 10723 14579
rect 10757 14545 10796 14579
rect 10830 14545 10869 14579
rect 11003 14576 11039 14610
rect 11003 14572 11005 14576
rect 11037 14538 11039 14542
rect 11003 14504 11039 14538
rect 11003 14500 11005 14504
rect 11037 14466 11039 14470
rect 11003 14432 11039 14466
rect 11003 14428 11005 14432
rect 9983 14369 10024 14403
rect 10058 14369 10099 14403
rect 10133 14369 10174 14403
rect 10208 14369 10249 14403
rect 10283 14369 10323 14403
rect 10357 14369 10397 14403
rect 10431 14369 10471 14403
rect 11037 14394 11039 14398
rect 11003 14360 11039 14394
rect 11003 14356 11005 14360
rect 11037 14322 11039 14326
rect 11003 14288 11039 14322
rect 11003 14284 11005 14288
rect 11037 14250 11039 14254
rect 11005 14238 11039 14250
rect 11295 14854 11465 14878
rect 11329 14820 11363 14854
rect 11397 14820 11431 14854
rect 11295 14785 11465 14820
rect 11329 14751 11363 14785
rect 11397 14783 11465 14785
rect 11397 14751 11431 14783
rect 11295 14749 11431 14751
rect 11295 14716 11465 14749
rect 11329 14682 11363 14716
rect 11397 14712 11465 14716
rect 11397 14682 11431 14712
rect 11295 14678 11431 14682
rect 11295 14647 11465 14678
rect 11329 14613 11363 14647
rect 11397 14641 11465 14647
rect 11397 14613 11431 14641
rect 11295 14607 11431 14613
rect 11295 14578 11465 14607
rect 11329 14544 11363 14578
rect 11397 14570 11465 14578
rect 11397 14544 11431 14570
rect 11295 14536 11431 14544
rect 11295 14509 11465 14536
rect 11329 14475 11363 14509
rect 11397 14499 11465 14509
rect 11397 14475 11431 14499
rect 11295 14465 11431 14475
rect 11295 14440 11465 14465
rect 11329 14406 11363 14440
rect 11397 14428 11465 14440
rect 11397 14406 11431 14428
rect 11295 14394 11431 14406
rect 11295 14371 11465 14394
rect 11295 14370 11363 14371
rect 11329 14337 11363 14370
rect 11397 14357 11465 14371
rect 11397 14337 11431 14357
rect 11329 14336 11431 14337
rect 11295 14323 11431 14336
rect 11295 14302 11465 14323
rect 11295 14300 11363 14302
rect 11329 14268 11363 14300
rect 11397 14286 11465 14302
rect 11397 14268 11431 14286
rect 11329 14266 11431 14268
rect 11295 14252 11431 14266
rect 11295 14232 11465 14252
rect 11295 14230 11363 14232
rect 10314 14193 10360 14227
rect 10394 14193 10440 14227
rect 10474 14193 10520 14227
rect 10554 14193 10600 14227
rect 10634 14193 10680 14227
rect 10714 14193 10759 14227
rect 10793 14193 10838 14227
rect 11329 14198 11363 14230
rect 11397 14214 11465 14232
rect 11397 14198 11431 14214
rect 11329 14196 11431 14198
rect 11005 14184 11039 14196
rect 11037 14180 11039 14184
rect 11003 14146 11005 14150
rect 11003 14112 11039 14146
rect 11003 14104 11005 14112
rect 11037 14070 11039 14078
rect 11005 14062 11039 14070
rect 11295 14180 11431 14196
rect 11295 14162 11465 14180
rect 11295 14160 11363 14162
rect 11329 14128 11363 14160
rect 11397 14142 11465 14162
rect 11397 14128 11431 14142
rect 11329 14126 11431 14128
rect 11295 14108 11431 14126
rect 11295 14092 11465 14108
rect 11295 14090 11363 14092
rect 11329 14058 11363 14090
rect 11397 14070 11465 14092
rect 11397 14058 11431 14070
rect 11329 14056 11431 14058
rect 10003 14017 10044 14051
rect 10078 14017 10119 14051
rect 10153 14017 10194 14051
rect 10228 14017 10269 14051
rect 10303 14017 10344 14051
rect 10378 14017 10419 14051
rect 10453 14017 10494 14051
rect 10528 14017 10569 14051
rect 10603 14017 10644 14051
rect 10678 14017 10719 14051
rect 10753 14017 10794 14051
rect 10828 14017 10869 14051
rect 11295 14036 11431 14056
rect 11295 14022 11465 14036
rect 11295 14020 11363 14022
rect 11329 13988 11363 14020
rect 11397 13998 11465 14022
rect 11397 13988 11431 13998
rect 11329 13986 11431 13988
rect 11295 13964 11431 13986
rect 11295 13952 11465 13964
rect 11295 13950 11363 13952
rect 11329 13918 11363 13950
rect 11397 13926 11465 13952
rect 11397 13918 11431 13926
rect 11329 13916 11431 13918
rect 11295 13892 11431 13916
rect 11295 13882 11465 13892
rect 11295 13880 11363 13882
rect 11329 13848 11363 13880
rect 11397 13854 11465 13882
rect 11397 13848 11431 13854
rect 11329 13846 11431 13848
rect 11295 13820 11431 13846
rect 11295 13812 11465 13820
rect 11295 13810 11363 13812
rect 11329 13778 11363 13810
rect 11397 13782 11465 13812
rect 11397 13778 11431 13782
rect 11329 13776 11431 13778
rect 11295 13748 11431 13776
rect 11295 13742 11465 13748
rect 11295 13740 11363 13742
rect 11118 13706 11142 13740
rect 11176 13706 11219 13740
rect 11253 13706 11295 13740
rect 11329 13708 11363 13740
rect 11397 13710 11465 13742
rect 11397 13708 11431 13710
rect 11329 13706 11431 13708
rect 11118 13676 11431 13706
rect 11118 13672 11465 13676
rect 11118 13638 11142 13672
rect 11176 13638 11216 13672
rect 11250 13638 11290 13672
rect 11324 13638 11363 13672
rect 11397 13638 11465 13672
rect 11118 13604 11431 13638
rect 11118 13570 11142 13604
rect 11176 13570 11223 13604
rect 11257 13570 11304 13604
rect 11338 13570 11465 13604
rect 10212 12884 10246 12908
rect 10212 12836 10246 12850
rect 10212 12762 10246 12802
rect 10370 12789 10386 12823
rect 10420 12811 10454 12823
rect 10436 12789 10454 12811
rect 10488 12789 10504 12823
rect 10212 9916 10246 12728
rect 10402 12731 10436 12777
rect 10328 12616 10362 12655
rect 10328 12543 10362 12582
rect 10328 12470 10362 12509
rect 10328 12397 10362 12436
rect 10328 12324 10362 12363
rect 10328 12252 10362 12290
rect 10328 12180 10362 12218
rect 10504 12616 10538 12655
rect 10504 12543 10538 12582
rect 10504 12470 10538 12509
rect 10504 12397 10538 12436
rect 10504 12324 10538 12363
rect 10504 12252 10538 12290
rect 10504 12180 10538 12218
rect 10212 9858 10246 9882
<< viali >>
rect 10280 15601 10314 15635
rect 10354 15601 10388 15635
rect 10428 15601 10462 15635
rect 10502 15601 10536 15635
rect 10576 15601 10610 15635
rect 10650 15601 10684 15635
rect 10723 15601 10757 15635
rect 10796 15601 10830 15635
rect 10869 15601 10903 15635
rect 11003 15574 11037 15590
rect 11003 15556 11005 15574
rect 11005 15556 11037 15574
rect 11003 15503 11037 15517
rect 11003 15483 11005 15503
rect 11005 15483 11037 15503
rect 9949 15425 9983 15459
rect 10024 15425 10058 15459
rect 10099 15425 10133 15459
rect 10174 15425 10208 15459
rect 10249 15425 10283 15459
rect 10323 15425 10357 15459
rect 10397 15425 10431 15459
rect 10471 15425 10505 15459
rect 11003 15432 11037 15444
rect 11003 15410 11005 15432
rect 11005 15410 11037 15432
rect 11003 15361 11037 15371
rect 11003 15337 11005 15361
rect 11005 15337 11037 15361
rect 11003 15290 11037 15298
rect 10280 15249 10314 15283
rect 10354 15249 10388 15283
rect 10428 15249 10462 15283
rect 10502 15249 10536 15283
rect 10576 15249 10610 15283
rect 10650 15249 10684 15283
rect 10723 15249 10757 15283
rect 10796 15249 10830 15283
rect 10869 15249 10903 15283
rect 11003 15264 11005 15290
rect 11005 15264 11037 15290
rect 11003 15219 11037 15225
rect 11003 15191 11005 15219
rect 11005 15191 11037 15219
rect 11003 15148 11037 15152
rect 11003 15118 11005 15148
rect 11005 15118 11037 15148
rect 9949 15073 9983 15107
rect 10024 15073 10058 15107
rect 10099 15073 10133 15107
rect 10174 15073 10208 15107
rect 10249 15073 10283 15107
rect 10323 15073 10357 15107
rect 10397 15073 10431 15107
rect 10471 15073 10505 15107
rect 11003 15077 11037 15079
rect 11003 15045 11005 15077
rect 11005 15045 11037 15077
rect 11003 14972 11005 15006
rect 11005 14972 11037 15006
rect 10280 14897 10314 14931
rect 10354 14897 10388 14931
rect 10428 14897 10462 14931
rect 10502 14897 10536 14931
rect 10576 14897 10610 14931
rect 10650 14897 10684 14931
rect 10723 14897 10757 14931
rect 10796 14897 10830 14931
rect 10869 14897 10903 14931
rect 11003 14901 11005 14933
rect 11005 14901 11037 14933
rect 11003 14899 11037 14901
rect 11003 14830 11005 14860
rect 11005 14830 11037 14860
rect 11003 14826 11037 14830
rect 11003 14758 11005 14788
rect 11005 14758 11037 14788
rect 9949 14721 9983 14755
rect 10024 14721 10058 14755
rect 10099 14721 10133 14755
rect 10174 14721 10208 14755
rect 10249 14721 10283 14755
rect 10323 14721 10357 14755
rect 10397 14721 10431 14755
rect 10471 14721 10505 14755
rect 11003 14754 11037 14758
rect 11003 14686 11005 14716
rect 11005 14686 11037 14716
rect 11003 14682 11037 14686
rect 11003 14614 11005 14644
rect 11005 14614 11037 14644
rect 11003 14610 11037 14614
rect 10280 14545 10314 14579
rect 10354 14545 10388 14579
rect 10428 14545 10462 14579
rect 10502 14545 10536 14579
rect 10576 14545 10610 14579
rect 10650 14545 10684 14579
rect 10723 14545 10757 14579
rect 10796 14545 10830 14579
rect 10869 14545 10903 14579
rect 11003 14542 11005 14572
rect 11005 14542 11037 14572
rect 11003 14538 11037 14542
rect 11003 14470 11005 14500
rect 11005 14470 11037 14500
rect 11003 14466 11037 14470
rect 9949 14369 9983 14403
rect 10024 14369 10058 14403
rect 10099 14369 10133 14403
rect 10174 14369 10208 14403
rect 10249 14369 10283 14403
rect 10323 14369 10357 14403
rect 10397 14369 10431 14403
rect 10471 14369 10505 14403
rect 11003 14398 11005 14428
rect 11005 14398 11037 14428
rect 11003 14394 11037 14398
rect 11003 14326 11005 14356
rect 11005 14326 11037 14356
rect 11003 14322 11037 14326
rect 11003 14254 11005 14284
rect 11005 14254 11037 14284
rect 11003 14250 11037 14254
rect 10280 14193 10314 14227
rect 10360 14193 10394 14227
rect 10440 14193 10474 14227
rect 10520 14193 10554 14227
rect 10600 14193 10634 14227
rect 10680 14193 10714 14227
rect 10759 14193 10793 14227
rect 10838 14193 10872 14227
rect 11003 14180 11037 14184
rect 11003 14150 11005 14180
rect 11005 14150 11037 14180
rect 11003 14078 11005 14104
rect 11005 14078 11037 14104
rect 11003 14070 11037 14078
rect 9969 14017 10003 14051
rect 10044 14017 10078 14051
rect 10119 14017 10153 14051
rect 10194 14017 10228 14051
rect 10269 14017 10303 14051
rect 10344 14017 10378 14051
rect 10419 14017 10453 14051
rect 10494 14017 10528 14051
rect 10569 14017 10603 14051
rect 10644 14017 10678 14051
rect 10719 14017 10753 14051
rect 10794 14017 10828 14051
rect 10869 14017 10903 14051
rect 10212 12802 10246 12836
rect 10402 12789 10420 12811
rect 10420 12789 10436 12811
rect 10212 12728 10246 12762
rect 10402 12777 10436 12789
rect 10402 12697 10436 12731
rect 10328 12655 10362 12689
rect 10328 12582 10362 12616
rect 10328 12509 10362 12543
rect 10328 12436 10362 12470
rect 10328 12363 10362 12397
rect 10328 12290 10362 12324
rect 10328 12218 10362 12252
rect 10328 12146 10362 12180
rect 10504 12655 10538 12689
rect 10504 12582 10538 12616
rect 10504 12509 10538 12543
rect 10504 12436 10538 12470
rect 10504 12363 10538 12397
rect 10504 12290 10538 12324
rect 10504 12218 10538 12252
rect 10504 12146 10538 12180
<< metal1 >>
tri 10538 15738 10563 15763 ne
tri 10538 15641 10563 15666 se
rect 10563 15641 10915 15763
tri 10915 15738 10940 15763 nw
rect 10268 15635 10915 15641
rect 10268 15601 10280 15635
rect 10314 15601 10354 15635
rect 10388 15601 10428 15635
rect 10462 15601 10502 15635
rect 10536 15601 10576 15635
rect 10610 15601 10650 15635
rect 10684 15601 10723 15635
rect 10757 15601 10796 15635
rect 10830 15601 10869 15635
rect 10903 15601 10915 15635
rect 10268 15595 10915 15601
tri 10538 15590 10543 15595 ne
rect 10543 15590 10915 15595
tri 10543 15570 10563 15590 ne
rect 9937 15459 10517 15465
rect 9937 15425 9949 15459
rect 9983 15425 10024 15459
rect 10058 15425 10099 15459
rect 10133 15425 10174 15459
rect 10208 15425 10249 15459
rect 10283 15425 10323 15459
rect 10357 15425 10397 15459
rect 10431 15425 10471 15459
rect 10505 15425 10517 15459
rect 9937 15419 10517 15425
rect 9937 15410 10238 15419
tri 10238 15410 10247 15419 nw
rect 9937 15402 10230 15410
tri 10230 15402 10238 15410 nw
rect 9937 15396 10222 15402
rect 9937 15344 9947 15396
rect 9999 15344 10011 15396
rect 10063 15344 10075 15396
rect 10127 15344 10222 15396
tri 10222 15394 10230 15402 nw
rect 10563 15396 10915 15590
rect 9937 15329 10222 15344
rect 9937 15277 9947 15329
rect 9999 15277 10011 15329
rect 10063 15277 10075 15329
rect 10127 15277 10222 15329
rect 10563 15344 10616 15396
rect 10668 15344 10680 15396
rect 10732 15344 10744 15396
rect 10796 15344 10808 15396
rect 10860 15344 10915 15396
rect 10563 15329 10915 15344
tri 10547 15298 10563 15314 se
rect 10563 15298 10616 15329
tri 10538 15289 10547 15298 se
rect 10547 15289 10616 15298
rect 9937 15262 10222 15277
rect 9937 15210 9947 15262
rect 9999 15210 10011 15262
rect 10063 15210 10075 15262
rect 10127 15210 10222 15262
rect 10268 15283 10616 15289
rect 10668 15283 10680 15329
rect 10732 15283 10744 15329
rect 10796 15283 10808 15329
rect 10860 15283 10915 15329
rect 10268 15249 10280 15283
rect 10314 15249 10354 15283
rect 10388 15249 10428 15283
rect 10462 15249 10502 15283
rect 10536 15249 10576 15283
rect 10610 15277 10616 15283
rect 10860 15277 10869 15283
rect 10610 15262 10650 15277
rect 10684 15262 10723 15277
rect 10757 15262 10796 15277
rect 10830 15262 10869 15277
rect 10610 15249 10616 15262
rect 10860 15249 10869 15262
rect 10903 15249 10915 15283
rect 10268 15243 10616 15249
tri 10538 15225 10556 15243 ne
rect 10556 15225 10616 15243
tri 10556 15218 10563 15225 ne
rect 9937 15195 10222 15210
rect 9937 15143 9947 15195
rect 9999 15143 10011 15195
rect 10063 15143 10075 15195
rect 10127 15143 10222 15195
rect 9937 15128 10222 15143
rect 10563 15210 10616 15225
rect 10668 15210 10680 15249
rect 10732 15210 10744 15249
rect 10796 15210 10808 15249
rect 10860 15210 10915 15249
rect 10563 15195 10915 15210
rect 10563 15143 10616 15195
rect 10668 15143 10680 15195
rect 10732 15143 10744 15195
rect 10796 15143 10808 15195
rect 10860 15143 10915 15195
rect 9937 15076 9947 15128
rect 9999 15076 10011 15128
rect 10063 15076 10075 15128
rect 10127 15118 10222 15128
tri 10222 15118 10242 15138 sw
rect 10563 15128 10915 15143
rect 10127 15113 10242 15118
tri 10242 15113 10247 15118 sw
rect 10127 15107 10517 15113
rect 9937 15073 9949 15076
rect 9983 15073 10024 15076
rect 10058 15073 10099 15076
rect 10133 15073 10174 15107
rect 10208 15073 10249 15107
rect 10283 15073 10323 15107
rect 10357 15073 10397 15107
rect 10431 15073 10471 15107
rect 10505 15073 10517 15107
rect 9937 15067 10517 15073
rect 10563 15076 10616 15128
rect 10668 15076 10680 15128
rect 10732 15076 10744 15128
rect 10796 15076 10808 15128
rect 10860 15076 10915 15128
rect 9937 15060 10225 15067
rect 9937 15008 9947 15060
rect 9999 15008 10011 15060
rect 10063 15008 10075 15060
rect 10127 15045 10225 15060
tri 10225 15045 10247 15067 nw
rect 10563 15061 10915 15076
rect 10127 15008 10222 15045
tri 10222 15042 10225 15045 nw
rect 9937 14992 10222 15008
rect 9937 14940 9947 14992
rect 9999 14940 10011 14992
rect 10063 14940 10075 14992
rect 10127 14940 10222 14992
rect 10563 15009 10616 15061
rect 10668 15009 10680 15061
rect 10732 15009 10744 15061
rect 10796 15009 10808 15061
rect 10860 15009 10915 15061
rect 10563 14994 10915 15009
rect 9937 14924 10222 14940
tri 10538 14937 10563 14962 se
rect 10563 14942 10616 14994
rect 10668 14942 10680 14994
rect 10732 14942 10744 14994
rect 10796 14942 10808 14994
rect 10860 14942 10915 14994
rect 10563 14937 10915 14942
rect 9937 14872 9947 14924
rect 9999 14872 10011 14924
rect 10063 14872 10075 14924
rect 10127 14872 10222 14924
rect 10268 14931 10915 14937
rect 10268 14897 10280 14931
rect 10314 14897 10354 14931
rect 10388 14897 10428 14931
rect 10462 14897 10502 14931
rect 10536 14897 10576 14931
rect 10610 14927 10650 14931
rect 10684 14927 10723 14931
rect 10757 14927 10796 14931
rect 10830 14927 10869 14931
rect 10610 14897 10616 14927
rect 10860 14897 10869 14927
rect 10903 14897 10915 14931
rect 10268 14891 10616 14897
rect 9937 14856 10222 14872
tri 10538 14866 10563 14891 ne
rect 10563 14875 10616 14891
rect 10668 14875 10680 14897
rect 10732 14875 10744 14897
rect 10796 14875 10808 14897
rect 10860 14875 10915 14897
rect 9937 14804 9947 14856
rect 9999 14804 10011 14856
rect 10063 14804 10075 14856
rect 10127 14804 10222 14856
rect 9937 14788 10222 14804
rect 9937 14736 9947 14788
rect 9999 14736 10011 14788
rect 10063 14736 10075 14788
rect 10127 14761 10222 14788
rect 10563 14860 10915 14875
rect 10563 14808 10616 14860
rect 10668 14808 10680 14860
rect 10732 14808 10744 14860
rect 10796 14808 10808 14860
rect 10860 14808 10915 14860
rect 10563 14792 10915 14808
tri 10222 14761 10247 14786 sw
rect 10127 14755 10517 14761
rect 9937 14721 9949 14736
rect 9983 14721 10024 14736
rect 10058 14721 10099 14736
rect 10133 14721 10174 14755
rect 10208 14721 10249 14755
rect 10283 14721 10323 14755
rect 10357 14721 10397 14755
rect 10431 14721 10471 14755
rect 10505 14721 10517 14755
rect 9937 14720 10517 14721
rect 9937 14668 9947 14720
rect 9999 14668 10011 14720
rect 10063 14668 10075 14720
rect 10127 14715 10517 14720
rect 10563 14740 10616 14792
rect 10668 14740 10680 14792
rect 10732 14740 10744 14792
rect 10796 14740 10808 14792
rect 10860 14740 10915 14792
rect 10563 14724 10915 14740
rect 10127 14668 10222 14715
tri 10222 14690 10247 14715 nw
rect 9937 14652 10222 14668
rect 9937 14600 9947 14652
rect 9999 14600 10011 14652
rect 10063 14600 10075 14652
rect 10127 14600 10222 14652
rect 10563 14672 10616 14724
rect 10668 14672 10680 14724
rect 10732 14672 10744 14724
rect 10796 14672 10808 14724
rect 10860 14672 10915 14724
rect 10563 14656 10915 14672
rect 9937 14584 10222 14600
tri 10538 14585 10563 14610 se
rect 10563 14604 10616 14656
rect 10668 14604 10680 14656
rect 10732 14604 10744 14656
rect 10796 14604 10808 14656
rect 10860 14604 10915 14656
rect 10563 14588 10915 14604
rect 10563 14585 10616 14588
rect 9937 14532 9947 14584
rect 9999 14532 10011 14584
rect 10063 14532 10075 14584
rect 10127 14532 10222 14584
rect 10268 14579 10616 14585
rect 10668 14579 10680 14588
rect 10732 14579 10744 14588
rect 10796 14579 10808 14588
rect 10860 14579 10915 14588
rect 10268 14545 10280 14579
rect 10314 14545 10354 14579
rect 10388 14545 10428 14579
rect 10462 14545 10502 14579
rect 10536 14545 10576 14579
rect 10610 14545 10616 14579
rect 10860 14545 10869 14579
rect 10903 14545 10915 14579
rect 10268 14539 10616 14545
tri 10538 14538 10539 14539 ne
rect 10539 14538 10616 14539
rect 9937 14428 10222 14532
tri 10539 14530 10547 14538 ne
rect 10547 14536 10616 14538
rect 10668 14536 10680 14545
rect 10732 14536 10744 14545
rect 10796 14536 10808 14545
rect 10860 14536 10915 14545
rect 10547 14530 10915 14536
tri 10547 14514 10563 14530 ne
tri 10222 14428 10228 14434 sw
rect 9937 14409 10228 14428
tri 10228 14409 10247 14428 sw
rect 9937 14403 10517 14409
rect 9937 14369 9949 14403
rect 9983 14369 10024 14403
rect 10058 14369 10099 14403
rect 10133 14369 10174 14403
rect 10208 14369 10249 14403
rect 10283 14369 10323 14403
rect 10357 14369 10397 14403
rect 10431 14369 10471 14403
rect 10505 14369 10517 14403
rect 9937 14363 10517 14369
rect 9937 14356 10240 14363
tri 10240 14356 10247 14363 nw
rect 9937 14201 10222 14356
tri 10222 14338 10240 14356 nw
rect 10563 14330 10915 14530
rect 10563 14325 10910 14330
tri 10910 14325 10915 14330 nw
rect 10997 15590 11043 15602
rect 10997 15556 11003 15590
rect 11037 15556 11043 15590
rect 10997 15517 11043 15556
rect 10997 15483 11003 15517
rect 11037 15483 11043 15517
rect 10997 15444 11043 15483
rect 10997 15410 11003 15444
rect 11037 15410 11043 15444
rect 10997 15371 11043 15410
rect 10997 15337 11003 15371
rect 11037 15337 11043 15371
rect 10997 15298 11043 15337
rect 10997 15264 11003 15298
rect 11037 15264 11043 15298
rect 10997 15225 11043 15264
rect 10997 15191 11003 15225
rect 11037 15191 11043 15225
rect 10997 15152 11043 15191
rect 10997 15118 11003 15152
rect 11037 15118 11043 15152
rect 10997 15079 11043 15118
rect 10997 15045 11003 15079
rect 11037 15045 11043 15079
rect 10997 15006 11043 15045
rect 10997 14972 11003 15006
rect 11037 14972 11043 15006
rect 10997 14933 11043 14972
rect 10997 14899 11003 14933
rect 11037 14899 11043 14933
rect 10997 14860 11043 14899
rect 10997 14826 11003 14860
rect 11037 14826 11043 14860
rect 10997 14788 11043 14826
rect 10997 14754 11003 14788
rect 11037 14754 11043 14788
rect 10997 14716 11043 14754
rect 10997 14682 11003 14716
rect 11037 14682 11043 14716
rect 10997 14644 11043 14682
rect 10997 14610 11003 14644
rect 11037 14610 11043 14644
rect 10997 14572 11043 14610
rect 10997 14538 11003 14572
rect 11037 14538 11043 14572
rect 10997 14500 11043 14538
rect 10997 14466 11003 14500
rect 11037 14466 11043 14500
rect 10997 14428 11043 14466
rect 10997 14394 11003 14428
rect 11037 14394 11043 14428
rect 10997 14356 11043 14394
rect 10563 14322 10907 14325
tri 10907 14322 10910 14325 nw
tri 10996 14322 10997 14323 se
rect 10997 14322 11003 14356
rect 11037 14322 11043 14356
tri 10555 14250 10563 14258 se
rect 10563 14250 10884 14322
tri 10884 14299 10907 14322 nw
tri 10973 14299 10996 14322 se
rect 10996 14299 11043 14322
tri 10958 14284 10973 14299 se
rect 10973 14284 11043 14299
tri 10924 14250 10958 14284 se
rect 10958 14250 11003 14284
rect 11037 14250 11043 14284
tri 10538 14233 10555 14250 se
rect 10555 14233 10884 14250
rect 10268 14227 10884 14233
rect 10268 14193 10280 14227
rect 10314 14193 10360 14227
rect 10394 14193 10440 14227
rect 10474 14193 10520 14227
rect 10554 14193 10600 14227
rect 10634 14193 10680 14227
rect 10714 14193 10759 14227
rect 10793 14193 10838 14227
rect 10872 14193 10884 14227
rect 10268 14187 10884 14193
tri 10912 14238 10924 14250 se
rect 10924 14238 11043 14250
rect 11239 15396 11505 15402
rect 11239 15344 11250 15396
rect 11302 15344 11314 15396
rect 11366 15344 11378 15396
rect 11430 15344 11442 15396
rect 11494 15344 11505 15396
rect 11239 15329 11505 15344
rect 11239 15277 11250 15329
rect 11302 15277 11314 15329
rect 11366 15277 11378 15329
rect 11430 15277 11442 15329
rect 11494 15277 11505 15329
rect 11239 15262 11505 15277
rect 11239 15210 11250 15262
rect 11302 15210 11314 15262
rect 11366 15210 11378 15262
rect 11430 15210 11442 15262
rect 11494 15210 11505 15262
rect 11239 15195 11505 15210
rect 11239 15143 11250 15195
rect 11302 15143 11314 15195
rect 11366 15143 11378 15195
rect 11430 15143 11442 15195
rect 11494 15143 11505 15195
rect 11239 15128 11505 15143
rect 11239 15076 11250 15128
rect 11302 15076 11314 15128
rect 11366 15076 11378 15128
rect 11430 15076 11442 15128
rect 11494 15076 11505 15128
rect 11239 15061 11505 15076
rect 11239 15009 11250 15061
rect 11302 15009 11314 15061
rect 11366 15009 11378 15061
rect 11430 15009 11442 15061
rect 11494 15009 11505 15061
rect 11239 14994 11505 15009
rect 11239 14942 11250 14994
rect 11302 14942 11314 14994
rect 11366 14942 11378 14994
rect 11430 14942 11442 14994
rect 11494 14942 11505 14994
rect 11239 14927 11505 14942
rect 11239 14875 11250 14927
rect 11302 14875 11314 14927
rect 11366 14875 11378 14927
rect 11430 14875 11442 14927
rect 11494 14875 11505 14927
rect 11239 14860 11505 14875
rect 11239 14808 11250 14860
rect 11302 14808 11314 14860
rect 11366 14808 11378 14860
rect 11430 14808 11442 14860
rect 11494 14808 11505 14860
rect 11239 14792 11505 14808
rect 11239 14740 11250 14792
rect 11302 14740 11314 14792
rect 11366 14740 11378 14792
rect 11430 14740 11442 14792
rect 11494 14740 11505 14792
rect 11239 14724 11505 14740
rect 11239 14672 11250 14724
rect 11302 14672 11314 14724
rect 11366 14672 11378 14724
rect 11430 14672 11442 14724
rect 11494 14672 11505 14724
rect 11239 14656 11505 14672
rect 11239 14604 11250 14656
rect 11302 14604 11314 14656
rect 11366 14604 11378 14656
rect 11430 14604 11442 14656
rect 11494 14604 11505 14656
rect 11239 14588 11505 14604
rect 11239 14536 11250 14588
rect 11302 14536 11314 14588
rect 11366 14536 11378 14588
rect 11430 14536 11442 14588
rect 11494 14536 11505 14588
tri 10900 14070 10912 14082 se
rect 10912 14070 10958 14238
tri 10958 14213 10983 14238 nw
tri 10888 14058 10900 14070 se
rect 10900 14058 10958 14070
tri 10887 14057 10888 14058 se
rect 10888 14057 10958 14058
rect 9957 14051 10236 14057
rect 10288 14051 10310 14057
rect 10362 14051 10958 14057
rect 9957 14017 9969 14051
rect 10003 14017 10044 14051
rect 10078 14017 10119 14051
rect 10153 14017 10194 14051
rect 10228 14017 10236 14051
rect 10303 14017 10310 14051
rect 10378 14017 10419 14051
rect 10453 14017 10494 14051
rect 10528 14017 10569 14051
rect 10603 14017 10644 14051
rect 10678 14017 10719 14051
rect 10753 14017 10794 14051
rect 10828 14017 10869 14051
rect 10903 14046 10958 14051
rect 10903 14017 10923 14046
rect 9957 14005 10236 14017
rect 10288 14005 10310 14017
rect 10362 14011 10923 14017
tri 10923 14011 10958 14046 nw
rect 10991 14190 11043 14196
rect 10991 14116 11043 14138
rect 10362 14005 10368 14011
tri 10368 14005 10374 14011 nw
tri 10967 13881 10991 13905 se
rect 10991 13886 11043 14064
rect 10991 13881 11034 13886
rect 9243 13829 9249 13881
rect 9301 13829 9313 13881
rect 9365 13829 9371 13881
rect 10230 13829 10236 13881
rect 10288 13829 10310 13881
rect 10362 13829 10368 13881
tri 10963 13877 10967 13881 se
rect 10967 13877 11034 13881
tri 11034 13877 11043 13886 nw
tri 7463 12972 7469 12978 nw
rect 7686 6286 7810 6673
tri 9236 2435 9243 2442 se
rect 9243 2435 9295 13829
tri 9295 13804 9320 13829 nw
tri 10297 13804 10322 13829 ne
rect 10090 12836 10252 12914
rect 10090 12802 10212 12836
rect 10246 12802 10252 12836
rect 10090 12762 10252 12802
rect 10090 12728 10212 12762
rect 10246 12728 10252 12762
rect 10090 10115 10252 12728
rect 10322 12689 10368 13829
rect 10322 12655 10328 12689
rect 10362 12655 10368 12689
rect 10396 13831 10988 13877
tri 10988 13831 11034 13877 nw
rect 10396 13829 10469 13831
tri 10469 13829 10471 13831 nw
rect 10396 13804 10444 13829
tri 10444 13804 10469 13829 nw
rect 10396 12811 10442 13804
tri 10442 13802 10444 13804 nw
rect 11239 13489 11505 14536
rect 11239 13437 11250 13489
rect 11302 13437 11314 13489
rect 11366 13437 11378 13489
rect 11430 13437 11442 13489
rect 11494 13437 11505 13489
rect 11239 13416 11505 13437
rect 11239 13364 11250 13416
rect 11302 13364 11314 13416
rect 11366 13364 11378 13416
rect 11430 13364 11442 13416
rect 11494 13364 11505 13416
rect 11239 13342 11505 13364
rect 11239 13290 11250 13342
rect 11302 13290 11314 13342
rect 11366 13290 11378 13342
rect 11430 13290 11442 13342
rect 11494 13290 11505 13342
rect 11239 13268 11505 13290
rect 11239 13216 11250 13268
rect 11302 13216 11314 13268
rect 11366 13216 11378 13268
rect 11430 13216 11442 13268
rect 11494 13216 11505 13268
rect 11239 13194 11505 13216
rect 11239 13142 11250 13194
rect 11302 13142 11314 13194
rect 11366 13142 11378 13194
rect 11430 13142 11442 13194
rect 11494 13142 11505 13194
rect 11239 13120 11505 13142
rect 11239 13068 11250 13120
rect 11302 13068 11314 13120
rect 11366 13068 11378 13120
rect 11430 13068 11442 13120
rect 11494 13068 11505 13120
rect 11239 13062 11505 13068
rect 10396 12777 10402 12811
rect 10436 12777 10442 12811
rect 10396 12731 10442 12777
rect 10396 12697 10402 12731
rect 10436 12697 10442 12731
rect 10396 12685 10442 12697
rect 10498 12689 10660 12914
rect 10322 12616 10368 12655
rect 10322 12582 10328 12616
rect 10362 12582 10368 12616
rect 10322 12543 10368 12582
rect 10322 12509 10328 12543
rect 10362 12509 10368 12543
rect 10322 12470 10368 12509
rect 10322 12436 10328 12470
rect 10362 12436 10368 12470
rect 10322 12397 10368 12436
rect 10322 12363 10328 12397
rect 10362 12363 10368 12397
rect 10322 12324 10368 12363
rect 10322 12290 10328 12324
rect 10362 12290 10368 12324
rect 10322 12252 10368 12290
rect 10322 12218 10328 12252
rect 10362 12218 10368 12252
rect 10322 12180 10368 12218
rect 10322 12146 10328 12180
rect 10362 12146 10368 12180
rect 10322 12134 10368 12146
rect 10498 12655 10504 12689
rect 10538 12655 10660 12689
rect 10498 12616 10660 12655
rect 10498 12582 10504 12616
rect 10538 12582 10660 12616
rect 10498 12543 10660 12582
rect 10498 12509 10504 12543
rect 10538 12509 10660 12543
rect 10498 12470 10660 12509
rect 10498 12436 10504 12470
rect 10538 12436 10660 12470
rect 10498 12397 10660 12436
rect 10498 12363 10504 12397
rect 10538 12363 10660 12397
rect 10498 12324 10660 12363
rect 10498 12290 10504 12324
rect 10538 12290 10660 12324
rect 10498 12252 10660 12290
rect 10498 12218 10504 12252
rect 10538 12218 10660 12252
rect 10498 12180 10660 12218
rect 10498 12146 10504 12180
rect 10538 12146 10660 12180
tri 10252 10115 10277 10140 sw
tri 10473 10115 10498 10140 se
rect 10498 10115 10660 12146
rect 10090 10063 10215 10115
rect 10267 10063 10280 10115
rect 10332 10063 10345 10115
rect 10397 10063 10410 10115
rect 10090 10051 10410 10063
rect 10090 9999 10215 10051
rect 10267 9999 10280 10051
rect 10332 9999 10345 10051
rect 10397 9999 10410 10051
rect 10090 9987 10410 9999
rect 10090 9935 10215 9987
rect 10267 9935 10280 9987
rect 10332 9935 10345 9987
rect 10397 9935 10410 9987
rect 10654 9935 10660 10115
rect 10090 9875 10660 9935
rect 10090 9850 10303 9875
tri 10303 9850 10328 9875 nw
tri 10448 9850 10473 9875 ne
rect 10473 9850 10660 9875
rect 10090 8911 10277 9850
tri 10277 9824 10303 9850 nw
tri 10277 9280 10302 9305 sw
tri 10277 9209 10302 9234 nw
rect 10090 8859 10097 8911
rect 10149 8859 10277 8911
rect 10090 8847 10277 8859
rect 10090 8795 10097 8847
rect 10149 8795 10277 8847
rect 10090 8783 10277 8795
rect 10090 8731 10097 8783
rect 10149 8731 10277 8783
rect 10090 8388 10277 8731
rect 10090 8336 10097 8388
rect 10149 8336 10277 8388
rect 10090 8324 10277 8336
rect 10090 8272 10097 8324
rect 10149 8272 10277 8324
rect 10090 8260 10277 8272
rect 10090 8208 10097 8260
rect 10149 8208 10277 8260
rect 10090 8202 10277 8208
tri 10161 8170 10193 8202 ne
tri 10245 8170 10277 8202 nw
tri 7557 2417 7575 2435 se
tri 9218 2417 9236 2435 se
rect 9236 2417 9295 2435
rect 7505 2365 7511 2417
rect 7563 2365 7575 2417
rect 7627 2365 7633 2417
rect 9167 2365 9173 2417
rect 9225 2365 9237 2417
rect 9289 2365 9295 2417
tri 7550 2340 7575 2365 ne
<< via1 >>
rect 9947 15344 9999 15396
rect 10011 15344 10063 15396
rect 10075 15344 10127 15396
rect 9947 15277 9999 15329
rect 10011 15277 10063 15329
rect 10075 15277 10127 15329
rect 10616 15344 10668 15396
rect 10680 15344 10732 15396
rect 10744 15344 10796 15396
rect 10808 15344 10860 15396
rect 9947 15210 9999 15262
rect 10011 15210 10063 15262
rect 10075 15210 10127 15262
rect 10616 15283 10668 15329
rect 10680 15283 10732 15329
rect 10744 15283 10796 15329
rect 10808 15283 10860 15329
rect 10616 15277 10650 15283
rect 10650 15277 10668 15283
rect 10680 15277 10684 15283
rect 10684 15277 10723 15283
rect 10723 15277 10732 15283
rect 10744 15277 10757 15283
rect 10757 15277 10796 15283
rect 10808 15277 10830 15283
rect 10830 15277 10860 15283
rect 10616 15249 10650 15262
rect 10650 15249 10668 15262
rect 10680 15249 10684 15262
rect 10684 15249 10723 15262
rect 10723 15249 10732 15262
rect 10744 15249 10757 15262
rect 10757 15249 10796 15262
rect 10808 15249 10830 15262
rect 10830 15249 10860 15262
rect 9947 15143 9999 15195
rect 10011 15143 10063 15195
rect 10075 15143 10127 15195
rect 10616 15210 10668 15249
rect 10680 15210 10732 15249
rect 10744 15210 10796 15249
rect 10808 15210 10860 15249
rect 10616 15143 10668 15195
rect 10680 15143 10732 15195
rect 10744 15143 10796 15195
rect 10808 15143 10860 15195
rect 9947 15107 9999 15128
rect 9947 15076 9949 15107
rect 9949 15076 9983 15107
rect 9983 15076 9999 15107
rect 10011 15107 10063 15128
rect 10011 15076 10024 15107
rect 10024 15076 10058 15107
rect 10058 15076 10063 15107
rect 10075 15107 10127 15128
rect 10075 15076 10099 15107
rect 10099 15076 10127 15107
rect 10616 15076 10668 15128
rect 10680 15076 10732 15128
rect 10744 15076 10796 15128
rect 10808 15076 10860 15128
rect 9947 15008 9999 15060
rect 10011 15008 10063 15060
rect 10075 15008 10127 15060
rect 9947 14940 9999 14992
rect 10011 14940 10063 14992
rect 10075 14940 10127 14992
rect 10616 15009 10668 15061
rect 10680 15009 10732 15061
rect 10744 15009 10796 15061
rect 10808 15009 10860 15061
rect 10616 14942 10668 14994
rect 10680 14942 10732 14994
rect 10744 14942 10796 14994
rect 10808 14942 10860 14994
rect 9947 14872 9999 14924
rect 10011 14872 10063 14924
rect 10075 14872 10127 14924
rect 10616 14897 10650 14927
rect 10650 14897 10668 14927
rect 10680 14897 10684 14927
rect 10684 14897 10723 14927
rect 10723 14897 10732 14927
rect 10744 14897 10757 14927
rect 10757 14897 10796 14927
rect 10808 14897 10830 14927
rect 10830 14897 10860 14927
rect 10616 14875 10668 14897
rect 10680 14875 10732 14897
rect 10744 14875 10796 14897
rect 10808 14875 10860 14897
rect 9947 14804 9999 14856
rect 10011 14804 10063 14856
rect 10075 14804 10127 14856
rect 9947 14755 9999 14788
rect 9947 14736 9949 14755
rect 9949 14736 9983 14755
rect 9983 14736 9999 14755
rect 10011 14755 10063 14788
rect 10011 14736 10024 14755
rect 10024 14736 10058 14755
rect 10058 14736 10063 14755
rect 10075 14755 10127 14788
rect 10616 14808 10668 14860
rect 10680 14808 10732 14860
rect 10744 14808 10796 14860
rect 10808 14808 10860 14860
rect 10075 14736 10099 14755
rect 10099 14736 10127 14755
rect 9947 14668 9999 14720
rect 10011 14668 10063 14720
rect 10075 14668 10127 14720
rect 10616 14740 10668 14792
rect 10680 14740 10732 14792
rect 10744 14740 10796 14792
rect 10808 14740 10860 14792
rect 9947 14600 9999 14652
rect 10011 14600 10063 14652
rect 10075 14600 10127 14652
rect 10616 14672 10668 14724
rect 10680 14672 10732 14724
rect 10744 14672 10796 14724
rect 10808 14672 10860 14724
rect 10616 14604 10668 14656
rect 10680 14604 10732 14656
rect 10744 14604 10796 14656
rect 10808 14604 10860 14656
rect 9947 14532 9999 14584
rect 10011 14532 10063 14584
rect 10075 14532 10127 14584
rect 10616 14579 10668 14588
rect 10680 14579 10732 14588
rect 10744 14579 10796 14588
rect 10808 14579 10860 14588
rect 10616 14545 10650 14579
rect 10650 14545 10668 14579
rect 10680 14545 10684 14579
rect 10684 14545 10723 14579
rect 10723 14545 10732 14579
rect 10744 14545 10757 14579
rect 10757 14545 10796 14579
rect 10808 14545 10830 14579
rect 10830 14545 10860 14579
rect 10616 14536 10668 14545
rect 10680 14536 10732 14545
rect 10744 14536 10796 14545
rect 10808 14536 10860 14545
rect 11250 15344 11302 15396
rect 11314 15344 11366 15396
rect 11378 15344 11430 15396
rect 11442 15344 11494 15396
rect 11250 15277 11302 15329
rect 11314 15277 11366 15329
rect 11378 15277 11430 15329
rect 11442 15277 11494 15329
rect 11250 15210 11302 15262
rect 11314 15210 11366 15262
rect 11378 15210 11430 15262
rect 11442 15210 11494 15262
rect 11250 15143 11302 15195
rect 11314 15143 11366 15195
rect 11378 15143 11430 15195
rect 11442 15143 11494 15195
rect 11250 15076 11302 15128
rect 11314 15076 11366 15128
rect 11378 15076 11430 15128
rect 11442 15076 11494 15128
rect 11250 15009 11302 15061
rect 11314 15009 11366 15061
rect 11378 15009 11430 15061
rect 11442 15009 11494 15061
rect 11250 14942 11302 14994
rect 11314 14942 11366 14994
rect 11378 14942 11430 14994
rect 11442 14942 11494 14994
rect 11250 14875 11302 14927
rect 11314 14875 11366 14927
rect 11378 14875 11430 14927
rect 11442 14875 11494 14927
rect 11250 14808 11302 14860
rect 11314 14808 11366 14860
rect 11378 14808 11430 14860
rect 11442 14808 11494 14860
rect 11250 14740 11302 14792
rect 11314 14740 11366 14792
rect 11378 14740 11430 14792
rect 11442 14740 11494 14792
rect 11250 14672 11302 14724
rect 11314 14672 11366 14724
rect 11378 14672 11430 14724
rect 11442 14672 11494 14724
rect 11250 14604 11302 14656
rect 11314 14604 11366 14656
rect 11378 14604 11430 14656
rect 11442 14604 11494 14656
rect 11250 14536 11302 14588
rect 11314 14536 11366 14588
rect 11378 14536 11430 14588
rect 11442 14536 11494 14588
rect 10236 14051 10288 14057
rect 10310 14051 10362 14057
rect 10236 14017 10269 14051
rect 10269 14017 10288 14051
rect 10310 14017 10344 14051
rect 10344 14017 10362 14051
rect 10236 14005 10288 14017
rect 10310 14005 10362 14017
rect 10991 14184 11043 14190
rect 10991 14150 11003 14184
rect 11003 14150 11037 14184
rect 11037 14150 11043 14184
rect 10991 14138 11043 14150
rect 10991 14104 11043 14116
rect 10991 14070 11003 14104
rect 11003 14070 11037 14104
rect 11037 14070 11043 14104
rect 10991 14064 11043 14070
rect 9249 13829 9301 13881
rect 9313 13829 9365 13881
rect 10236 13829 10288 13881
rect 10310 13829 10362 13881
rect 11250 13437 11302 13489
rect 11314 13437 11366 13489
rect 11378 13437 11430 13489
rect 11442 13437 11494 13489
rect 11250 13364 11302 13416
rect 11314 13364 11366 13416
rect 11378 13364 11430 13416
rect 11442 13364 11494 13416
rect 11250 13290 11302 13342
rect 11314 13290 11366 13342
rect 11378 13290 11430 13342
rect 11442 13290 11494 13342
rect 11250 13216 11302 13268
rect 11314 13216 11366 13268
rect 11378 13216 11430 13268
rect 11442 13216 11494 13268
rect 11250 13142 11302 13194
rect 11314 13142 11366 13194
rect 11378 13142 11430 13194
rect 11442 13142 11494 13194
rect 11250 13068 11302 13120
rect 11314 13068 11366 13120
rect 11378 13068 11430 13120
rect 11442 13068 11494 13120
rect 10215 10063 10267 10115
rect 10280 10063 10332 10115
rect 10345 10063 10397 10115
rect 10215 9999 10267 10051
rect 10280 9999 10332 10051
rect 10345 9999 10397 10051
rect 10215 9935 10267 9987
rect 10280 9935 10332 9987
rect 10345 9935 10397 9987
rect 10410 9935 10654 10115
rect 10097 8859 10149 8911
rect 10097 8795 10149 8847
rect 10097 8731 10149 8783
rect 10097 8336 10149 8388
rect 10097 8272 10149 8324
rect 10097 8208 10149 8260
rect 7511 2365 7563 2417
rect 7575 2365 7627 2417
rect 9173 2365 9225 2417
rect 9237 2365 9289 2417
<< metal2 >>
rect 9947 15396 10127 15402
rect 9999 15344 10011 15396
rect 10063 15344 10075 15396
rect 9947 15329 10127 15344
rect 9999 15277 10011 15329
rect 10063 15277 10075 15329
rect 9947 15262 10127 15277
rect 9999 15210 10011 15262
rect 10063 15210 10075 15262
rect 9947 15195 10127 15210
rect 9999 15143 10011 15195
rect 10063 15143 10075 15195
rect 9947 15128 10127 15143
rect 9999 15076 10011 15128
rect 10063 15076 10075 15128
rect 9947 15074 10127 15076
tri 9922 15061 9935 15074 ne
rect 9935 15061 10127 15074
tri 9935 15060 9936 15061 ne
rect 9936 15060 10127 15061
tri 9936 15049 9947 15060 ne
rect 9999 15008 10011 15060
rect 10063 15008 10075 15060
rect 9947 14992 10127 15008
rect 9999 14940 10011 14992
rect 10063 14940 10075 14992
rect 9947 14924 10127 14940
rect 9999 14872 10011 14924
rect 10063 14872 10075 14924
rect 9947 14856 10127 14872
rect 9999 14804 10011 14856
rect 10063 14804 10075 14856
rect 9947 14788 10127 14804
rect 9999 14736 10011 14788
rect 10063 14736 10075 14788
rect 9947 14720 10127 14736
rect 9999 14668 10011 14720
rect 10063 14668 10075 14720
rect 9947 14652 10127 14668
rect 9999 14600 10011 14652
rect 10063 14600 10075 14652
rect 9947 14584 10127 14600
rect 9999 14532 10011 14584
rect 10063 14532 10075 14584
rect 9947 14526 10127 14532
rect 10605 15396 11505 15402
rect 10605 15344 10616 15396
rect 10668 15344 10680 15396
rect 10732 15344 10744 15396
rect 10796 15344 10808 15396
rect 10860 15344 11250 15396
rect 11302 15344 11314 15396
rect 11366 15344 11378 15396
rect 11430 15344 11442 15396
rect 11494 15344 11505 15396
rect 10605 15329 11505 15344
rect 10605 15277 10616 15329
rect 10668 15277 10680 15329
rect 10732 15277 10744 15329
rect 10796 15277 10808 15329
rect 10860 15277 11250 15329
rect 11302 15277 11314 15329
rect 11366 15277 11378 15329
rect 11430 15277 11442 15329
rect 11494 15277 11505 15329
rect 10605 15262 11505 15277
rect 10605 15210 10616 15262
rect 10668 15210 10680 15262
rect 10732 15210 10744 15262
rect 10796 15210 10808 15262
rect 10860 15210 11250 15262
rect 11302 15210 11314 15262
rect 11366 15210 11378 15262
rect 11430 15210 11442 15262
rect 11494 15210 11505 15262
rect 10605 15195 11505 15210
rect 10605 15143 10616 15195
rect 10668 15143 10680 15195
rect 10732 15143 10744 15195
rect 10796 15143 10808 15195
rect 10860 15143 11250 15195
rect 11302 15143 11314 15195
rect 11366 15143 11378 15195
rect 11430 15143 11442 15195
rect 11494 15143 11505 15195
rect 10605 15128 11505 15143
rect 10605 15076 10616 15128
rect 10668 15076 10680 15128
rect 10732 15076 10744 15128
rect 10796 15076 10808 15128
rect 10860 15076 11250 15128
rect 11302 15076 11314 15128
rect 11366 15076 11378 15128
rect 11430 15076 11442 15128
rect 11494 15076 11505 15128
rect 10605 15061 11505 15076
rect 10605 15009 10616 15061
rect 10668 15009 10680 15061
rect 10732 15009 10744 15061
rect 10796 15009 10808 15061
rect 10860 15009 11250 15061
rect 11302 15009 11314 15061
rect 11366 15009 11378 15061
rect 11430 15009 11442 15061
rect 11494 15009 11505 15061
rect 10605 14994 11505 15009
rect 10605 14942 10616 14994
rect 10668 14942 10680 14994
rect 10732 14942 10744 14994
rect 10796 14942 10808 14994
rect 10860 14942 11250 14994
rect 11302 14942 11314 14994
rect 11366 14942 11378 14994
rect 11430 14942 11442 14994
rect 11494 14942 11505 14994
rect 10605 14927 11505 14942
rect 10605 14875 10616 14927
rect 10668 14875 10680 14927
rect 10732 14875 10744 14927
rect 10796 14875 10808 14927
rect 10860 14875 11250 14927
rect 11302 14875 11314 14927
rect 11366 14875 11378 14927
rect 11430 14875 11442 14927
rect 11494 14875 11505 14927
rect 10605 14860 11505 14875
rect 10605 14808 10616 14860
rect 10668 14808 10680 14860
rect 10732 14808 10744 14860
rect 10796 14808 10808 14860
rect 10860 14808 11250 14860
rect 11302 14808 11314 14860
rect 11366 14808 11378 14860
rect 11430 14808 11442 14860
rect 11494 14808 11505 14860
rect 10605 14792 11505 14808
rect 10605 14740 10616 14792
rect 10668 14740 10680 14792
rect 10732 14740 10744 14792
rect 10796 14740 10808 14792
rect 10860 14740 11250 14792
rect 11302 14740 11314 14792
rect 11366 14740 11378 14792
rect 11430 14740 11442 14792
rect 11494 14740 11505 14792
rect 10605 14724 11505 14740
rect 10605 14672 10616 14724
rect 10668 14672 10680 14724
rect 10732 14672 10744 14724
rect 10796 14672 10808 14724
rect 10860 14672 11250 14724
rect 11302 14672 11314 14724
rect 11366 14672 11378 14724
rect 11430 14672 11442 14724
rect 11494 14672 11505 14724
rect 10605 14656 11505 14672
rect 10605 14604 10616 14656
rect 10668 14604 10680 14656
rect 10732 14604 10744 14656
rect 10796 14604 10808 14656
rect 10860 14604 11250 14656
rect 11302 14604 11314 14656
rect 11366 14604 11378 14656
rect 11430 14604 11442 14656
rect 11494 14604 11505 14656
rect 10605 14588 11505 14604
rect 10605 14536 10616 14588
rect 10668 14536 10680 14588
rect 10732 14536 10744 14588
rect 10796 14536 10808 14588
rect 10860 14536 11250 14588
rect 11302 14536 11314 14588
rect 11366 14536 11378 14588
rect 11430 14536 11442 14588
rect 11494 14536 11505 14588
rect 10605 14530 11505 14536
rect 1202 14274 9783 14326
tri 9761 14270 9765 14274 ne
rect 9765 14270 9783 14274
tri 9783 14270 9839 14326 sw
tri 9765 14252 9783 14270 ne
rect 9783 14252 9839 14270
tri 9783 14196 9839 14252 ne
tri 9839 14196 9913 14270 sw
tri 9839 14190 9845 14196 ne
rect 9845 14190 11043 14196
tri 9845 14144 9891 14190 ne
rect 9891 14144 10991 14190
tri 10905 14138 10911 14144 ne
rect 10911 14138 10991 14144
tri 10911 14116 10933 14138 ne
rect 10933 14116 11043 14138
tri 10933 14064 10985 14116 ne
rect 10985 14064 10991 14116
tri 10985 14058 10991 14064 ne
rect 10991 14058 11043 14064
rect 10230 14005 10236 14057
rect 10288 14005 10310 14057
rect 10362 14005 10368 14057
rect 1202 13888 9165 13940
tri 9143 13881 9150 13888 ne
rect 9150 13881 9165 13888
tri 9165 13881 9224 13940 sw
tri 10205 13881 10230 13906 se
rect 10230 13881 10368 14005
rect 13182 13925 13266 14055
tri 9150 13866 9165 13881 ne
rect 9165 13866 9249 13881
tri 9165 13829 9202 13866 ne
rect 9202 13829 9249 13866
rect 9301 13829 9313 13881
rect 9365 13829 10236 13881
rect 10288 13829 10310 13881
rect 10362 13829 10368 13881
rect 13182 13739 13266 13869
rect 11239 13489 11505 13495
rect 11239 13437 11250 13489
rect 11302 13437 11314 13489
rect 11366 13437 11378 13489
rect 11430 13437 11442 13489
rect 11494 13437 11505 13489
rect 11239 13416 11505 13437
rect 11239 13364 11250 13416
rect 11302 13364 11314 13416
rect 11366 13364 11378 13416
rect 11430 13364 11442 13416
rect 11494 13364 11505 13416
rect 11239 13342 11505 13364
rect 11239 13290 11250 13342
rect 11302 13290 11314 13342
rect 11366 13290 11378 13342
rect 11430 13290 11442 13342
rect 11494 13290 11505 13342
rect 11239 13268 11505 13290
rect 11239 13216 11250 13268
rect 11302 13216 11314 13268
rect 11366 13216 11378 13268
rect 11430 13216 11442 13268
rect 11494 13216 11505 13268
rect 11239 13194 11505 13216
rect 11239 13142 11250 13194
rect 11302 13142 11314 13194
rect 11366 13142 11378 13194
rect 11430 13142 11442 13194
rect 11494 13142 11505 13194
rect 11239 13120 11505 13142
rect 11239 13068 11250 13120
rect 11302 13068 11314 13120
rect 11366 13068 11378 13120
rect 11430 13068 11442 13120
rect 11494 13068 11505 13120
rect 11239 13062 11505 13068
tri 1176 12978 1179 12981 ne
rect 1117 11625 1149 11818
rect 1117 10799 1152 11083
rect 1117 9849 1151 10115
rect 10206 10063 10215 10115
rect 10267 10063 10280 10115
rect 10332 10063 10345 10115
rect 10397 10063 10410 10115
rect 10206 10051 10410 10063
rect 10206 9999 10215 10051
rect 10267 9999 10280 10051
rect 10332 9999 10345 10051
rect 10397 9999 10410 10051
rect 10206 9987 10410 9999
rect 10206 9935 10215 9987
rect 10267 9935 10280 9987
rect 10332 9935 10345 9987
rect 10397 9935 10410 9987
rect 10654 9935 10660 10115
rect 10206 9849 10660 9935
rect 1117 9528 1145 9721
rect 12797 9209 12868 9339
rect 1117 8724 1148 8916
rect 10091 8859 10097 8911
rect 10149 8859 10155 8911
rect 10091 8847 10155 8859
rect 10091 8795 10097 8847
rect 10149 8795 10155 8847
rect 10091 8783 10155 8795
rect 10091 8731 10097 8783
rect 10149 8731 10155 8783
rect 1117 8202 1150 8394
rect 10091 8336 10097 8388
rect 10149 8336 10155 8388
rect 10091 8324 10155 8336
rect 10091 8272 10097 8324
rect 10149 8272 10155 8324
rect 10091 8260 10155 8272
rect 10091 8208 10097 8260
rect 10149 8208 10155 8260
rect 1117 7021 1150 7213
rect 4290 6727 4348 6857
rect 1117 6325 1144 6455
rect 1117 5586 1150 5778
rect 1117 3315 9308 3641
rect 1117 2816 8809 3315
tri 8809 2816 9308 3315 nw
rect 7505 2365 7511 2417
rect 7563 2365 7575 2417
rect 7627 2365 9173 2417
rect 9225 2365 9237 2417
rect 9289 2365 9295 2417
rect 1119 2114 1164 2166
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 9371 0 1 13829
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 9295 0 1 2365
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 7633 0 1 2365
box 0 0 1 1
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1707688321
transform -1 0 10493 0 1 12151
box -79 -26 199 626
use pfet_CDNS_52468879185313  pfet_CDNS_52468879185313_0
timestamp 1707688321
transform 0 1 9957 -1 0 14182
box -119 -66 239 1066
use pfet_CDNS_524688791851645  pfet_CDNS_524688791851645_0
timestamp 1707688321
transform 0 1 9957 1 0 14238
box -119 -66 1471 1066
use sky130_fd_io__sio_opamp_stage_c_c  sky130_fd_io__sio_opamp_stage_c_c_0
timestamp 1707688321
transform 1 0 0 0 1 1569
box 1022 -289 13266 14527
<< labels >>
flabel comment s 9723 2618 9723 2618 0 FreeSans 100 270 0 0 li_jumper_ok
flabel comment s 1410 2603 1410 2603 0 FreeSans 100 270 0 0 li_jumper_ok
flabel metal1 s 7686 6286 7810 6673 0 FreeSans 1000 90 0 0 fb_out
port 2 nsew
flabel metal2 s 1202 14274 1237 14326 0 FreeSans 200 0 0 0 vreg_en_h
port 3 nsew
flabel metal2 s 13182 13925 13266 14055 0 FreeSans 200 0 0 0 refleak_bias
port 4 nsew
flabel metal2 s 1202 13888 1237 13940 0 FreeSans 200 0 0 0 vreg_en_h_n
port 5 nsew
flabel metal2 s 1117 11625 1149 11818 0 FreeSans 200 0 0 0 vcc_io
port 6 nsew
flabel metal2 s 1119 2114 1164 2166 0 FreeSans 200 0 0 0 en_hicc
port 7 nsew
flabel metal2 s 1117 9528 1145 9721 0 FreeSans 200 0 0 0 vcc_io
port 6 nsew
flabel metal2 s 1117 6325 1144 6455 0 FreeSans 200 0 0 0 vcc_io
port 6 nsew
flabel metal2 s 1117 5586 1150 5778 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 7021 1150 7213 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 8202 1150 8394 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 8724 1148 8916 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 9849 1151 10115 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 10799 1152 11083 0 FreeSans 200 0 0 0 vgnd
port 8 nsew
flabel metal2 s 1117 2816 1399 3641 0 FreeSans 1000 90 0 0 vgnd
port 8 nsew
flabel metal2 s 4290 6727 4348 6857 0 FreeSans 1000 90 0 0 fb_in
port 9 nsew
flabel metal2 s 13182 13739 13266 13869 0 FreeSans 200 0 0 0 voutref
port 10 nsew
flabel metal2 s 12797 9209 12868 9339 0 FreeSans 200 0 0 0 fb_out
port 2 nsew
<< properties >>
string GDS_END 97340834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97303580
string path 259.200 346.375 255.750 346.375 
<< end >>
