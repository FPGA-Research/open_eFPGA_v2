magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 0 0 472 3549
<< ndiff >>
rect 26 3515 86 3523
rect 26 3481 39 3515
rect 73 3481 86 3515
rect 26 3447 86 3481
rect 26 3413 39 3447
rect 73 3413 86 3447
rect 386 3515 446 3523
rect 386 3481 399 3515
rect 433 3481 446 3515
rect 386 3447 446 3481
rect 386 3413 399 3447
rect 433 3413 446 3447
<< ndiffc >>
rect 39 3481 73 3515
rect 39 3413 73 3447
rect 399 3481 433 3515
rect 399 3413 433 3447
<< ndiffres >>
rect 26 86 86 3413
rect 146 3463 326 3523
rect 146 86 206 3463
rect 26 26 206 86
rect 266 86 326 3463
rect 386 86 446 3413
rect 266 26 446 86
<< locali >>
rect 23 3481 39 3515
rect 73 3481 89 3515
rect 23 3447 89 3481
rect 23 3413 39 3447
rect 73 3413 89 3447
rect 383 3481 399 3515
rect 433 3481 449 3515
rect 383 3447 449 3481
rect 383 3413 399 3447
rect 433 3413 449 3447
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform 0 1 387 -1 0 3455
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 0 1 27 -1 0 3523
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1707688321
transform 0 1 387 -1 0 3523
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1707688321
transform 0 1 27 -1 0 3455
box 0 0 1 1
<< properties >>
string GDS_END 6670932
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6669320
<< end >>
