magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< locali >>
rect 0 2861 300 3000
rect 0 2827 133 2861
rect 167 2827 300 2861
rect 0 2765 300 2827
rect 0 2731 133 2765
rect 167 2731 300 2765
rect 0 2669 300 2731
rect 0 2635 133 2669
rect 167 2635 300 2669
rect 0 2573 300 2635
rect 0 2539 133 2573
rect 167 2539 300 2573
rect 0 2477 300 2539
rect 0 2443 133 2477
rect 167 2443 300 2477
rect 0 2381 300 2443
rect 0 2347 133 2381
rect 167 2347 300 2381
rect 0 2285 300 2347
rect 0 2251 133 2285
rect 167 2251 300 2285
rect 0 2189 300 2251
rect 0 2155 133 2189
rect 167 2155 300 2189
rect 0 2093 300 2155
rect 0 2059 133 2093
rect 167 2059 300 2093
rect 0 1997 300 2059
rect 0 1963 133 1997
rect 167 1963 300 1997
rect 0 1901 300 1963
rect 0 1867 133 1901
rect 167 1867 300 1901
rect 0 1805 300 1867
rect 0 1771 133 1805
rect 167 1771 300 1805
rect 0 1709 300 1771
rect 0 1675 133 1709
rect 167 1675 300 1709
rect 0 1613 300 1675
rect 0 1579 133 1613
rect 167 1579 300 1613
rect 0 1517 300 1579
rect 0 1483 133 1517
rect 167 1483 300 1517
rect 0 1421 300 1483
rect 0 1387 133 1421
rect 167 1387 300 1421
rect 0 1325 300 1387
rect 0 1291 133 1325
rect 167 1291 300 1325
rect 0 1229 300 1291
rect 0 1195 133 1229
rect 167 1195 300 1229
rect 0 1133 300 1195
rect 0 1099 133 1133
rect 167 1099 300 1133
rect 0 1037 300 1099
rect 0 1003 133 1037
rect 167 1003 300 1037
rect 0 941 300 1003
rect 0 907 133 941
rect 167 907 300 941
rect 0 845 300 907
rect 0 811 133 845
rect 167 811 300 845
rect 0 749 300 811
rect 0 715 133 749
rect 167 715 300 749
rect 0 653 300 715
rect 0 619 133 653
rect 167 619 300 653
rect 0 557 300 619
rect 0 523 133 557
rect 167 523 300 557
rect 0 461 300 523
rect 0 427 133 461
rect 167 427 300 461
rect 0 365 300 427
rect 0 331 133 365
rect 167 331 300 365
rect 0 269 300 331
rect 0 235 133 269
rect 167 235 300 269
rect 0 173 300 235
rect 0 139 133 173
rect 167 139 300 173
rect 0 0 300 139
<< viali >>
rect 133 2827 167 2861
rect 133 2731 167 2765
rect 133 2635 167 2669
rect 133 2539 167 2573
rect 133 2443 167 2477
rect 133 2347 167 2381
rect 133 2251 167 2285
rect 133 2155 167 2189
rect 133 2059 167 2093
rect 133 1963 167 1997
rect 133 1867 167 1901
rect 133 1771 167 1805
rect 133 1675 167 1709
rect 133 1579 167 1613
rect 133 1483 167 1517
rect 133 1387 167 1421
rect 133 1291 167 1325
rect 133 1195 167 1229
rect 133 1099 167 1133
rect 133 1003 167 1037
rect 133 907 167 941
rect 133 811 167 845
rect 133 715 167 749
rect 133 619 167 653
rect 133 523 167 557
rect 133 427 167 461
rect 133 331 167 365
rect 133 235 167 269
rect 133 139 167 173
<< metal1 >>
tri 0 2940 60 3000 se
rect 60 2940 240 3000
tri 240 2940 300 3000 sw
rect 0 2861 300 2940
rect 0 2827 133 2861
rect 167 2827 300 2861
rect 0 2765 300 2827
rect 0 2731 133 2765
rect 167 2731 300 2765
rect 0 2669 300 2731
rect 0 2635 133 2669
rect 167 2635 300 2669
rect 0 2573 300 2635
rect 0 2539 133 2573
rect 167 2539 300 2573
rect 0 2477 300 2539
rect 0 2443 133 2477
rect 167 2443 300 2477
rect 0 2381 300 2443
rect 0 2347 133 2381
rect 167 2347 300 2381
rect 0 2285 300 2347
rect 0 2251 133 2285
rect 167 2251 300 2285
rect 0 2189 300 2251
rect 0 2155 133 2189
rect 167 2155 300 2189
rect 0 2093 300 2155
rect 0 2059 133 2093
rect 167 2059 300 2093
rect 0 1997 300 2059
rect 0 1963 133 1997
rect 167 1963 300 1997
rect 0 1901 300 1963
rect 0 1867 133 1901
rect 167 1867 300 1901
rect 0 1805 300 1867
rect 0 1771 133 1805
rect 167 1771 300 1805
rect 0 1709 300 1771
rect 0 1675 133 1709
rect 167 1675 300 1709
rect 0 1613 300 1675
rect 0 1579 133 1613
rect 167 1579 300 1613
rect 0 1517 300 1579
rect 0 1483 133 1517
rect 167 1483 300 1517
rect 0 1421 300 1483
rect 0 1387 133 1421
rect 167 1387 300 1421
rect 0 1325 300 1387
rect 0 1291 133 1325
rect 167 1291 300 1325
rect 0 1229 300 1291
rect 0 1195 133 1229
rect 167 1195 300 1229
rect 0 1133 300 1195
rect 0 1099 133 1133
rect 167 1099 300 1133
rect 0 1037 300 1099
rect 0 1003 133 1037
rect 167 1003 300 1037
rect 0 941 300 1003
rect 0 907 133 941
rect 167 907 300 941
rect 0 845 300 907
rect 0 811 133 845
rect 167 811 300 845
rect 0 749 300 811
rect 0 715 133 749
rect 167 715 300 749
rect 0 653 300 715
rect 0 619 133 653
rect 167 619 300 653
rect 0 557 300 619
rect 0 523 133 557
rect 167 523 300 557
rect 0 461 300 523
rect 0 427 133 461
rect 167 427 300 461
rect 0 365 300 427
rect 0 331 133 365
rect 167 331 300 365
rect 0 269 300 331
rect 0 235 133 269
rect 167 235 300 269
rect 0 173 300 235
rect 0 139 133 173
rect 167 139 300 173
rect 0 60 300 139
tri 0 0 60 60 ne
rect 60 0 240 60
tri 240 0 300 60 nw
use L1M1_CDNS_55959141808683  L1M1_CDNS_55959141808683_0
timestamp 1707688321
transform 1 0 61 0 1 139
box -12 -6 190 2728
<< properties >>
string GDS_END 42971096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42958020
<< end >>
