magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -133 -66 236 666
<< mvpmos >>
rect 0 0 120 600
<< mvpdiff >>
rect -50 0 0 600
rect 120 0 170 600
<< poly >>
rect 0 600 120 626
rect 0 -26 120 0
<< locali >>
rect -59 -4 -25 538
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_0
timestamp 1707688321
transform -1 0 -14 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -42 267 -42 267 0 FreeSans 300 0 0 0 S
flabel comment s 145 300 145 300 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 67709588
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 67708622
<< end >>
