
module eFPGA_top (I_top, T_top, O_top, A_config_C, B_config_C, CLK, SelfWriteStrobe, SelfWriteData, Rx, ComActive, ReceiveLED, s_clk, s_data);
	// External USER ports 
	//inout [16-1:0] PAD; // these are for Dirk and go to the pad ring
	output [24-1:0] I_top; 
	output [24-1:0] T_top;
	input  [24-1:0] O_top;
	output [48-1:0] A_config_C;
	output [48-1:0] B_config_C;

	input CLK; // This clock can go to the CPU (connects to the fabric LUT output flops

	// CPU configuration port
	input SelfWriteStrobe; // must decode address and write enable
	input [32-1:0] SelfWriteData; // configuration data write port

	// UART configuration port
	input Rx;
	output ComActive;
	output ReceiveLED;

	// BitBang configuration port
	input s_clk;
	input s_data;

	parameter include_eFPGA = 1;
	parameter NumberOfRows = 12;
	parameter NumberOfCols = 14;
	parameter FrameBitsPerRow = 32;
	parameter MaxFramesPerCol = 20;
	parameter desync_flag = 20;
	parameter FrameSelectWidth = 5;
	parameter RowSelectWidth = 5;

	//BlockRAM ports
	wire [180-1:0] RAM2FAB_D;
	wire [192-1:0] FAB2RAM_D;
	wire [96-1:0] FAB2RAM_A;
	wire [48-1:0] FAB2RAM_C;
	wire [48-1:0] Config_accessC;

	// Signal declarations
	wire [(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;

	wire [(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;

	wire [(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;

	wire [FrameBitsPerRow-1:0] FrameAddressRegister;
	wire LongFrameStrobe;
	wire [31:0] LocalWriteData;
	wire LocalWriteStrobe;
	wire [RowSelectWidth-1:0] RowSelect;


Config Config_inst (
	.CLK(CLK),
	.Rx(Rx),
	.ComActive(ComActive),
	.ReceiveLED(ReceiveLED),
	.s_clk(s_clk),
	.s_data(s_data),
	.SelfWriteData(SelfWriteData),
	.SelfWriteStrobe(SelfWriteStrobe),
	
	.ConfigWriteData(LocalWriteData),
	.ConfigWriteStrobe(LocalWriteStrobe),
	
	.FrameAddressRegister(FrameAddressRegister),
	.LongFrameStrobe(LongFrameStrobe),
	.RowSelect(RowSelect)
);


	// L: if include_eFPGA = 1 generate

	Frame_Data_Reg_0 Inst_Frame_Data_Reg_0 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[0*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_1 Inst_Frame_Data_Reg_1 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[1*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_2 Inst_Frame_Data_Reg_2 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[2*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_3 Inst_Frame_Data_Reg_3 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[3*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_4 Inst_Frame_Data_Reg_4 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[4*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_5 Inst_Frame_Data_Reg_5 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[5*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_6 Inst_Frame_Data_Reg_6 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[6*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_7 Inst_Frame_Data_Reg_7 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[7*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_8 Inst_Frame_Data_Reg_8 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[8*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_9 Inst_Frame_Data_Reg_9 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[9*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_10 Inst_Frame_Data_Reg_10 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[10*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Data_Reg_11 Inst_Frame_Data_Reg_11 (
	.FrameData_I(LocalWriteData),
	.FrameData_O(FrameRegister[11*FrameBitsPerRow+:FrameBitsPerRow]),
	.RowSelect(RowSelect),
	.CLK(CLK)
	);

	Frame_Select_0 Inst_Frame_Select_0 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[0*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_1 Inst_Frame_Select_1 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[1*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_2 Inst_Frame_Select_2 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[2*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_3 Inst_Frame_Select_3 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[3*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_4 Inst_Frame_Select_4 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[4*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_5 Inst_Frame_Select_5 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[5*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_6 Inst_Frame_Select_6 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[6*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_7 Inst_Frame_Select_7 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[7*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_8 Inst_Frame_Select_8 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[8*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_9 Inst_Frame_Select_9 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[9*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_10 Inst_Frame_Select_10 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[10*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_11 Inst_Frame_Select_11 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[11*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_12 Inst_Frame_Select_12 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[12*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	Frame_Select_13 Inst_Frame_Select_13 (
	.FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
	.FrameStrobe_O(FrameSelect[13*MaxFramesPerCol +: MaxFramesPerCol]),
	.FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-(FrameSelectWidth)]),
	.FrameStrobe(LongFrameStrobe)
	);

	wire [11:0] dump;

	eFPGA Inst_eFPGA(
	.Tile_X0Y1_A_I_top(I_top[23]),
	.Tile_X0Y1_B_I_top(I_top[22]),
	.Tile_X0Y2_A_I_top(I_top[21]),
	.Tile_X0Y2_B_I_top(I_top[20]),
	.Tile_X0Y3_A_I_top(I_top[19]),
	.Tile_X0Y3_B_I_top(I_top[18]),
	.Tile_X0Y4_A_I_top(I_top[17]),
	.Tile_X0Y4_B_I_top(I_top[16]),
	.Tile_X0Y5_A_I_top(I_top[15]),
	.Tile_X0Y5_B_I_top(I_top[14]),
	.Tile_X0Y6_A_I_top(I_top[13]),
	.Tile_X0Y6_B_I_top(I_top[12]),
	.Tile_X0Y7_A_I_top(I_top[11]),
	.Tile_X0Y7_B_I_top(I_top[10]),
	.Tile_X0Y8_A_I_top(I_top[9]),
	.Tile_X0Y8_B_I_top(I_top[8]),
	.Tile_X0Y9_A_I_top(I_top[7]),
	.Tile_X0Y9_B_I_top(I_top[6]),
	.Tile_X0Y10_A_I_top(I_top[5]),
	.Tile_X0Y10_B_I_top(I_top[4]),
	.Tile_X0Y11_A_I_top(I_top[3]),
	.Tile_X0Y11_B_I_top(I_top[2]),
	.Tile_X0Y12_A_I_top(I_top[1]),
	.Tile_X0Y12_B_I_top(I_top[0]),

	.Tile_X0Y1_A_T_top(T_top[23]),
	.Tile_X0Y1_B_T_top(T_top[22]),
	.Tile_X0Y2_A_T_top(T_top[21]),
	.Tile_X0Y2_B_T_top(T_top[20]),
	.Tile_X0Y3_A_T_top(T_top[19]),
	.Tile_X0Y3_B_T_top(T_top[18]),
	.Tile_X0Y4_A_T_top(T_top[17]),
	.Tile_X0Y4_B_T_top(T_top[16]),
	.Tile_X0Y5_A_T_top(T_top[15]),
	.Tile_X0Y5_B_T_top(T_top[14]),
	.Tile_X0Y6_A_T_top(T_top[13]),
	.Tile_X0Y6_B_T_top(T_top[12]),
	.Tile_X0Y7_A_T_top(T_top[11]),
	.Tile_X0Y7_B_T_top(T_top[10]),
	.Tile_X0Y8_A_T_top(T_top[9]),
	.Tile_X0Y8_B_T_top(T_top[8]),
	.Tile_X0Y9_A_T_top(T_top[7]),
	.Tile_X0Y9_B_T_top(T_top[6]),
	.Tile_X0Y10_A_T_top(T_top[5]),
	.Tile_X0Y10_B_T_top(T_top[4]),
	.Tile_X0Y11_A_T_top(T_top[3]),
	.Tile_X0Y11_B_T_top(T_top[2]),
	.Tile_X0Y12_A_T_top(T_top[1]),
	.Tile_X0Y12_B_T_top(T_top[0]),

	.Tile_X0Y1_A_O_top(O_top[23]),
	.Tile_X0Y1_B_O_top(O_top[22]),
	.Tile_X0Y2_A_O_top(O_top[21]),
	.Tile_X0Y2_B_O_top(O_top[20]),
	.Tile_X0Y3_A_O_top(O_top[19]),
	.Tile_X0Y3_B_O_top(O_top[18]),
	.Tile_X0Y4_A_O_top(O_top[17]),
	.Tile_X0Y4_B_O_top(O_top[16]),
	.Tile_X0Y5_A_O_top(O_top[15]),
	.Tile_X0Y5_B_O_top(O_top[14]),
	.Tile_X0Y6_A_O_top(O_top[13]),
	.Tile_X0Y6_B_O_top(O_top[12]),
	.Tile_X0Y7_A_O_top(O_top[11]),
	.Tile_X0Y7_B_O_top(O_top[10]),
	.Tile_X0Y8_A_O_top(O_top[9]),
	.Tile_X0Y8_B_O_top(O_top[8]),
	.Tile_X0Y9_A_O_top(O_top[7]),
	.Tile_X0Y9_B_O_top(O_top[6]),
	.Tile_X0Y10_A_O_top(O_top[5]),
	.Tile_X0Y10_B_O_top(O_top[4]),
	.Tile_X0Y11_A_O_top(O_top[3]),
	.Tile_X0Y11_B_O_top(O_top[2]),
	.Tile_X0Y12_A_O_top(O_top[1]),
	.Tile_X0Y12_B_O_top(O_top[0]),

	.Tile_X0Y1_A_config_C_bit0(A_config_C[47]),
	.Tile_X0Y1_A_config_C_bit1(A_config_C[46]),
	.Tile_X0Y1_A_config_C_bit2(A_config_C[45]),
	.Tile_X0Y1_A_config_C_bit3(A_config_C[44]),
	.Tile_X0Y2_A_config_C_bit0(A_config_C[43]),
	.Tile_X0Y2_A_config_C_bit1(A_config_C[42]),
	.Tile_X0Y2_A_config_C_bit2(A_config_C[41]),
	.Tile_X0Y2_A_config_C_bit3(A_config_C[40]),
	.Tile_X0Y3_A_config_C_bit0(A_config_C[39]),
	.Tile_X0Y3_A_config_C_bit1(A_config_C[38]),
	.Tile_X0Y3_A_config_C_bit2(A_config_C[37]),
	.Tile_X0Y3_A_config_C_bit3(A_config_C[36]),
	.Tile_X0Y4_A_config_C_bit0(A_config_C[35]),
	.Tile_X0Y4_A_config_C_bit1(A_config_C[34]),
	.Tile_X0Y4_A_config_C_bit2(A_config_C[33]),
	.Tile_X0Y4_A_config_C_bit3(A_config_C[32]),
	.Tile_X0Y5_A_config_C_bit0(A_config_C[31]),
	.Tile_X0Y5_A_config_C_bit1(A_config_C[30]),
	.Tile_X0Y5_A_config_C_bit2(A_config_C[29]),
	.Tile_X0Y5_A_config_C_bit3(A_config_C[28]),
	.Tile_X0Y6_A_config_C_bit0(A_config_C[27]),
	.Tile_X0Y6_A_config_C_bit1(A_config_C[26]),
	.Tile_X0Y6_A_config_C_bit2(A_config_C[25]),
	.Tile_X0Y6_A_config_C_bit3(A_config_C[24]),
	.Tile_X0Y7_A_config_C_bit0(A_config_C[23]),
	.Tile_X0Y7_A_config_C_bit1(A_config_C[22]),
	.Tile_X0Y7_A_config_C_bit2(A_config_C[21]),
	.Tile_X0Y7_A_config_C_bit3(A_config_C[20]),
	.Tile_X0Y8_A_config_C_bit0(A_config_C[19]),
	.Tile_X0Y8_A_config_C_bit1(A_config_C[18]),
	.Tile_X0Y8_A_config_C_bit2(A_config_C[17]),
	.Tile_X0Y8_A_config_C_bit3(A_config_C[16]),
	.Tile_X0Y9_A_config_C_bit0(A_config_C[15]),
	.Tile_X0Y9_A_config_C_bit1(A_config_C[14]),
	.Tile_X0Y9_A_config_C_bit2(A_config_C[13]),
	.Tile_X0Y9_A_config_C_bit3(A_config_C[12]),
	.Tile_X0Y10_A_config_C_bit0(A_config_C[11]),
	.Tile_X0Y10_A_config_C_bit1(A_config_C[10]),
	.Tile_X0Y10_A_config_C_bit2(A_config_C[9]),
	.Tile_X0Y10_A_config_C_bit3(A_config_C[8]),
	.Tile_X0Y11_A_config_C_bit0(A_config_C[7]),
	.Tile_X0Y11_A_config_C_bit1(A_config_C[6]),
	.Tile_X0Y11_A_config_C_bit2(A_config_C[5]),
	.Tile_X0Y11_A_config_C_bit3(A_config_C[4]),
	.Tile_X0Y12_A_config_C_bit0(A_config_C[3]),
	.Tile_X0Y12_A_config_C_bit1(A_config_C[2]),
	.Tile_X0Y12_A_config_C_bit2(A_config_C[1]),
	.Tile_X0Y12_A_config_C_bit3(A_config_C[0]),

	.Tile_X0Y1_B_config_C_bit0(B_config_C[47]),
	.Tile_X0Y1_B_config_C_bit1(B_config_C[46]),
	.Tile_X0Y1_B_config_C_bit2(B_config_C[45]),
	.Tile_X0Y1_B_config_C_bit3(B_config_C[44]),
	.Tile_X0Y2_B_config_C_bit0(B_config_C[43]),
	.Tile_X0Y2_B_config_C_bit1(B_config_C[42]),
	.Tile_X0Y2_B_config_C_bit2(B_config_C[41]),
	.Tile_X0Y2_B_config_C_bit3(B_config_C[40]),
	.Tile_X0Y3_B_config_C_bit0(B_config_C[39]),
	.Tile_X0Y3_B_config_C_bit1(B_config_C[38]),
	.Tile_X0Y3_B_config_C_bit2(B_config_C[37]),
	.Tile_X0Y3_B_config_C_bit3(B_config_C[36]),
	.Tile_X0Y4_B_config_C_bit0(B_config_C[35]),
	.Tile_X0Y4_B_config_C_bit1(B_config_C[34]),
	.Tile_X0Y4_B_config_C_bit2(B_config_C[33]),
	.Tile_X0Y4_B_config_C_bit3(B_config_C[32]),
	.Tile_X0Y5_B_config_C_bit0(B_config_C[31]),
	.Tile_X0Y5_B_config_C_bit1(B_config_C[30]),
	.Tile_X0Y5_B_config_C_bit2(B_config_C[29]),
	.Tile_X0Y5_B_config_C_bit3(B_config_C[28]),
	.Tile_X0Y6_B_config_C_bit0(B_config_C[27]),
	.Tile_X0Y6_B_config_C_bit1(B_config_C[26]),
	.Tile_X0Y6_B_config_C_bit2(B_config_C[25]),
	.Tile_X0Y6_B_config_C_bit3(B_config_C[24]),
	.Tile_X0Y7_B_config_C_bit0(B_config_C[23]),
	.Tile_X0Y7_B_config_C_bit1(B_config_C[22]),
	.Tile_X0Y7_B_config_C_bit2(B_config_C[21]),
	.Tile_X0Y7_B_config_C_bit3(B_config_C[20]),
	.Tile_X0Y8_B_config_C_bit0(B_config_C[19]),
	.Tile_X0Y8_B_config_C_bit1(B_config_C[18]),
	.Tile_X0Y8_B_config_C_bit2(B_config_C[17]),
	.Tile_X0Y8_B_config_C_bit3(B_config_C[16]),
	.Tile_X0Y9_B_config_C_bit0(B_config_C[15]),
	.Tile_X0Y9_B_config_C_bit1(B_config_C[14]),
	.Tile_X0Y9_B_config_C_bit2(B_config_C[13]),
	.Tile_X0Y9_B_config_C_bit3(B_config_C[12]),
	.Tile_X0Y10_B_config_C_bit0(B_config_C[11]),
	.Tile_X0Y10_B_config_C_bit1(B_config_C[10]),
	.Tile_X0Y10_B_config_C_bit2(B_config_C[9]),
	.Tile_X0Y10_B_config_C_bit3(B_config_C[8]),
	.Tile_X0Y11_B_config_C_bit0(B_config_C[7]),
	.Tile_X0Y11_B_config_C_bit1(B_config_C[6]),
	.Tile_X0Y11_B_config_C_bit2(B_config_C[5]),
	.Tile_X0Y11_B_config_C_bit3(B_config_C[4]),
	.Tile_X0Y12_B_config_C_bit0(B_config_C[3]),
	.Tile_X0Y12_B_config_C_bit1(B_config_C[2]),
	.Tile_X0Y12_B_config_C_bit2(B_config_C[1]),
	.Tile_X0Y12_B_config_C_bit3(B_config_C[0]),

	.Tile_X13Y1_RAM2FAB_D0_I0(RAM2FAB_D[179]),
	.Tile_X13Y1_RAM2FAB_D0_I1(RAM2FAB_D[178]),
	.Tile_X13Y1_RAM2FAB_D0_I2(RAM2FAB_D[177]),
	.Tile_X13Y1_RAM2FAB_D0_I3(RAM2FAB_D[176]),
	.Tile_X13Y1_RAM2FAB_D1_I0(RAM2FAB_D[175]),
	.Tile_X13Y1_RAM2FAB_D1_I1(RAM2FAB_D[174]),
	.Tile_X13Y1_RAM2FAB_D1_I2(dump[11]),
	.Tile_X13Y1_RAM2FAB_D1_I3(RAM2FAB_D[173]),
	.Tile_X13Y1_RAM2FAB_D2_I0(RAM2FAB_D[172]),
	.Tile_X13Y1_RAM2FAB_D2_I1(RAM2FAB_D[171]),
	.Tile_X13Y1_RAM2FAB_D2_I2(RAM2FAB_D[170]),
	.Tile_X13Y1_RAM2FAB_D2_I3(RAM2FAB_D[169]),
	.Tile_X13Y1_RAM2FAB_D3_I0(RAM2FAB_D[168]),
	.Tile_X13Y1_RAM2FAB_D3_I1(RAM2FAB_D[167]),
	.Tile_X13Y1_RAM2FAB_D3_I2(RAM2FAB_D[166]),
	.Tile_X13Y1_RAM2FAB_D3_I3(RAM2FAB_D[165]),
	.Tile_X13Y2_RAM2FAB_D0_I0(RAM2FAB_D[164]),
	.Tile_X13Y2_RAM2FAB_D0_I1(RAM2FAB_D[163]),
	.Tile_X13Y2_RAM2FAB_D0_I2(RAM2FAB_D[162]),
	.Tile_X13Y2_RAM2FAB_D0_I3(RAM2FAB_D[161]),
	.Tile_X13Y2_RAM2FAB_D1_I0(RAM2FAB_D[160]),
	.Tile_X13Y2_RAM2FAB_D1_I1(RAM2FAB_D[159]),
	.Tile_X13Y2_RAM2FAB_D1_I2(dump[10]),
	.Tile_X13Y2_RAM2FAB_D1_I3(RAM2FAB_D[158]),
	.Tile_X13Y2_RAM2FAB_D2_I0(RAM2FAB_D[157]),
	.Tile_X13Y2_RAM2FAB_D2_I1(RAM2FAB_D[156]),
	.Tile_X13Y2_RAM2FAB_D2_I2(RAM2FAB_D[155]),
	.Tile_X13Y2_RAM2FAB_D2_I3(RAM2FAB_D[154]),
	.Tile_X13Y2_RAM2FAB_D3_I0(RAM2FAB_D[153]),
	.Tile_X13Y2_RAM2FAB_D3_I1(RAM2FAB_D[152]),
	.Tile_X13Y2_RAM2FAB_D3_I2(RAM2FAB_D[151]),
	.Tile_X13Y2_RAM2FAB_D3_I3(RAM2FAB_D[150]),
	.Tile_X13Y3_RAM2FAB_D0_I0(RAM2FAB_D[149]),
	.Tile_X13Y3_RAM2FAB_D0_I1(RAM2FAB_D[148]),
	.Tile_X13Y3_RAM2FAB_D0_I2(RAM2FAB_D[147]),
	.Tile_X13Y3_RAM2FAB_D0_I3(RAM2FAB_D[146]),
	.Tile_X13Y3_RAM2FAB_D1_I0(RAM2FAB_D[145]),
	.Tile_X13Y3_RAM2FAB_D1_I1(RAM2FAB_D[144]),
	.Tile_X13Y3_RAM2FAB_D1_I2(dump[9]),
	.Tile_X13Y3_RAM2FAB_D1_I3(RAM2FAB_D[143]),
	.Tile_X13Y3_RAM2FAB_D2_I0(RAM2FAB_D[142]),
	.Tile_X13Y3_RAM2FAB_D2_I1(RAM2FAB_D[141]),
	.Tile_X13Y3_RAM2FAB_D2_I2(RAM2FAB_D[140]),
	.Tile_X13Y3_RAM2FAB_D2_I3(RAM2FAB_D[139]),
	.Tile_X13Y3_RAM2FAB_D3_I0(RAM2FAB_D[138]),
	.Tile_X13Y3_RAM2FAB_D3_I1(RAM2FAB_D[137]),
	.Tile_X13Y3_RAM2FAB_D3_I2(RAM2FAB_D[136]),
	.Tile_X13Y3_RAM2FAB_D3_I3(RAM2FAB_D[135]),
	.Tile_X13Y4_RAM2FAB_D0_I0(RAM2FAB_D[134]),
	.Tile_X13Y4_RAM2FAB_D0_I1(RAM2FAB_D[133]),
	.Tile_X13Y4_RAM2FAB_D0_I2(RAM2FAB_D[132]),
	.Tile_X13Y4_RAM2FAB_D0_I3(RAM2FAB_D[131]),
	.Tile_X13Y4_RAM2FAB_D1_I0(RAM2FAB_D[130]),
	.Tile_X13Y4_RAM2FAB_D1_I1(RAM2FAB_D[129]),
	.Tile_X13Y4_RAM2FAB_D1_I2(dump[8]),
	.Tile_X13Y4_RAM2FAB_D1_I3(RAM2FAB_D[128]),
	.Tile_X13Y4_RAM2FAB_D2_I0(RAM2FAB_D[127]),
	.Tile_X13Y4_RAM2FAB_D2_I1(RAM2FAB_D[126]),
	.Tile_X13Y4_RAM2FAB_D2_I2(RAM2FAB_D[125]),
	.Tile_X13Y4_RAM2FAB_D2_I3(RAM2FAB_D[124]),
	.Tile_X13Y4_RAM2FAB_D3_I0(RAM2FAB_D[123]),
	.Tile_X13Y4_RAM2FAB_D3_I1(RAM2FAB_D[122]),
	.Tile_X13Y4_RAM2FAB_D3_I2(RAM2FAB_D[121]),
	.Tile_X13Y4_RAM2FAB_D3_I3(RAM2FAB_D[120]),
	.Tile_X13Y5_RAM2FAB_D0_I0(RAM2FAB_D[119]),
	.Tile_X13Y5_RAM2FAB_D0_I1(RAM2FAB_D[118]),
	.Tile_X13Y5_RAM2FAB_D0_I2(RAM2FAB_D[117]),
	.Tile_X13Y5_RAM2FAB_D0_I3(RAM2FAB_D[116]),
	.Tile_X13Y5_RAM2FAB_D1_I0(RAM2FAB_D[115]),
	.Tile_X13Y5_RAM2FAB_D1_I1(RAM2FAB_D[114]),
	.Tile_X13Y5_RAM2FAB_D1_I2(dump[7]),
	.Tile_X13Y5_RAM2FAB_D1_I3(RAM2FAB_D[113]),
	.Tile_X13Y5_RAM2FAB_D2_I0(RAM2FAB_D[112]),
	.Tile_X13Y5_RAM2FAB_D2_I1(RAM2FAB_D[111]),
	.Tile_X13Y5_RAM2FAB_D2_I2(RAM2FAB_D[110]),
	.Tile_X13Y5_RAM2FAB_D2_I3(RAM2FAB_D[109]),
	.Tile_X13Y5_RAM2FAB_D3_I0(RAM2FAB_D[108]),
	.Tile_X13Y5_RAM2FAB_D3_I1(RAM2FAB_D[107]),
	.Tile_X13Y5_RAM2FAB_D3_I2(RAM2FAB_D[106]),
	.Tile_X13Y5_RAM2FAB_D3_I3(RAM2FAB_D[105]),
	.Tile_X13Y6_RAM2FAB_D0_I0(RAM2FAB_D[104]),
	.Tile_X13Y6_RAM2FAB_D0_I1(RAM2FAB_D[103]),
	.Tile_X13Y6_RAM2FAB_D0_I2(RAM2FAB_D[102]),
	.Tile_X13Y6_RAM2FAB_D0_I3(RAM2FAB_D[101]),
	.Tile_X13Y6_RAM2FAB_D1_I0(RAM2FAB_D[100]),
	.Tile_X13Y6_RAM2FAB_D1_I1(RAM2FAB_D[99]),
	.Tile_X13Y6_RAM2FAB_D1_I2(dump[6]),
	.Tile_X13Y6_RAM2FAB_D1_I3(RAM2FAB_D[98]),
	.Tile_X13Y6_RAM2FAB_D2_I0(RAM2FAB_D[97]),
	.Tile_X13Y6_RAM2FAB_D2_I1(RAM2FAB_D[96]),
	.Tile_X13Y6_RAM2FAB_D2_I2(RAM2FAB_D[95]),
	.Tile_X13Y6_RAM2FAB_D2_I3(RAM2FAB_D[94]),
	.Tile_X13Y6_RAM2FAB_D3_I0(RAM2FAB_D[93]),
	.Tile_X13Y6_RAM2FAB_D3_I1(RAM2FAB_D[92]),
	.Tile_X13Y6_RAM2FAB_D3_I2(RAM2FAB_D[91]),
	.Tile_X13Y6_RAM2FAB_D3_I3(RAM2FAB_D[90]),
	.Tile_X13Y7_RAM2FAB_D0_I0(RAM2FAB_D[89]),
	.Tile_X13Y7_RAM2FAB_D0_I1(RAM2FAB_D[88]),
	.Tile_X13Y7_RAM2FAB_D0_I2(RAM2FAB_D[87]),
	.Tile_X13Y7_RAM2FAB_D0_I3(RAM2FAB_D[86]),
	.Tile_X13Y7_RAM2FAB_D1_I0(RAM2FAB_D[85]),
	.Tile_X13Y7_RAM2FAB_D1_I1(RAM2FAB_D[84]),
	.Tile_X13Y7_RAM2FAB_D1_I2(dump[5]),
	.Tile_X13Y7_RAM2FAB_D1_I3(RAM2FAB_D[83]),
	.Tile_X13Y7_RAM2FAB_D2_I0(RAM2FAB_D[82]),
	.Tile_X13Y7_RAM2FAB_D2_I1(RAM2FAB_D[81]),
	.Tile_X13Y7_RAM2FAB_D2_I2(RAM2FAB_D[80]),
	.Tile_X13Y7_RAM2FAB_D2_I3(RAM2FAB_D[79]),
	.Tile_X13Y7_RAM2FAB_D3_I0(RAM2FAB_D[78]),
	.Tile_X13Y7_RAM2FAB_D3_I1(RAM2FAB_D[77]),
	.Tile_X13Y7_RAM2FAB_D3_I2(RAM2FAB_D[76]),
	.Tile_X13Y7_RAM2FAB_D3_I3(RAM2FAB_D[75]),
	.Tile_X13Y8_RAM2FAB_D0_I0(RAM2FAB_D[74]),
	.Tile_X13Y8_RAM2FAB_D0_I1(RAM2FAB_D[73]),
	.Tile_X13Y8_RAM2FAB_D0_I2(RAM2FAB_D[72]),
	.Tile_X13Y8_RAM2FAB_D0_I3(RAM2FAB_D[71]),
	.Tile_X13Y8_RAM2FAB_D1_I0(RAM2FAB_D[70]),
	.Tile_X13Y8_RAM2FAB_D1_I1(RAM2FAB_D[69]),
	.Tile_X13Y8_RAM2FAB_D1_I2(dump[4]),
	.Tile_X13Y8_RAM2FAB_D1_I3(RAM2FAB_D[68]),
	.Tile_X13Y8_RAM2FAB_D2_I0(RAM2FAB_D[67]),
	.Tile_X13Y8_RAM2FAB_D2_I1(RAM2FAB_D[66]),
	.Tile_X13Y8_RAM2FAB_D2_I2(RAM2FAB_D[65]),
	.Tile_X13Y8_RAM2FAB_D2_I3(RAM2FAB_D[64]),
	.Tile_X13Y8_RAM2FAB_D3_I0(RAM2FAB_D[63]),
	.Tile_X13Y8_RAM2FAB_D3_I1(RAM2FAB_D[62]),
	.Tile_X13Y8_RAM2FAB_D3_I2(RAM2FAB_D[61]),
	.Tile_X13Y8_RAM2FAB_D3_I3(RAM2FAB_D[60]),
	.Tile_X13Y9_RAM2FAB_D0_I0(RAM2FAB_D[59]),
	.Tile_X13Y9_RAM2FAB_D0_I1(RAM2FAB_D[58]),
	.Tile_X13Y9_RAM2FAB_D0_I2(RAM2FAB_D[57]),
	.Tile_X13Y9_RAM2FAB_D0_I3(RAM2FAB_D[56]),
	.Tile_X13Y9_RAM2FAB_D1_I0(RAM2FAB_D[55]),
	.Tile_X13Y9_RAM2FAB_D1_I1(RAM2FAB_D[54]),
	.Tile_X13Y9_RAM2FAB_D1_I2(dump[3]),
	.Tile_X13Y9_RAM2FAB_D1_I3(RAM2FAB_D[53]),
	.Tile_X13Y9_RAM2FAB_D2_I0(RAM2FAB_D[52]),
	.Tile_X13Y9_RAM2FAB_D2_I1(RAM2FAB_D[51]),
	.Tile_X13Y9_RAM2FAB_D2_I2(RAM2FAB_D[50]),
	.Tile_X13Y9_RAM2FAB_D2_I3(RAM2FAB_D[49]),
	.Tile_X13Y9_RAM2FAB_D3_I0(RAM2FAB_D[48]),
	.Tile_X13Y9_RAM2FAB_D3_I1(RAM2FAB_D[47]),
	.Tile_X13Y9_RAM2FAB_D3_I2(RAM2FAB_D[46]),
	.Tile_X13Y9_RAM2FAB_D3_I3(RAM2FAB_D[45]),
	.Tile_X13Y10_RAM2FAB_D0_I0(RAM2FAB_D[44]),
	.Tile_X13Y10_RAM2FAB_D0_I1(RAM2FAB_D[43]),
	.Tile_X13Y10_RAM2FAB_D0_I2(RAM2FAB_D[42]),
	.Tile_X13Y10_RAM2FAB_D0_I3(RAM2FAB_D[41]),
	.Tile_X13Y10_RAM2FAB_D1_I0(RAM2FAB_D[40]),
	.Tile_X13Y10_RAM2FAB_D1_I1(RAM2FAB_D[39]),
	.Tile_X13Y10_RAM2FAB_D1_I2(dump[2]),
	.Tile_X13Y10_RAM2FAB_D1_I3(RAM2FAB_D[38]),
	.Tile_X13Y10_RAM2FAB_D2_I0(RAM2FAB_D[37]),
	.Tile_X13Y10_RAM2FAB_D2_I1(RAM2FAB_D[36]),
	.Tile_X13Y10_RAM2FAB_D2_I2(RAM2FAB_D[35]),
	.Tile_X13Y10_RAM2FAB_D2_I3(RAM2FAB_D[34]),
	.Tile_X13Y10_RAM2FAB_D3_I0(RAM2FAB_D[33]),
	.Tile_X13Y10_RAM2FAB_D3_I1(RAM2FAB_D[32]),
	.Tile_X13Y10_RAM2FAB_D3_I2(RAM2FAB_D[31]),
	.Tile_X13Y10_RAM2FAB_D3_I3(RAM2FAB_D[30]),
	.Tile_X13Y11_RAM2FAB_D0_I0(RAM2FAB_D[29]),
	.Tile_X13Y11_RAM2FAB_D0_I1(RAM2FAB_D[28]),
	.Tile_X13Y11_RAM2FAB_D0_I2(RAM2FAB_D[27]),
	.Tile_X13Y11_RAM2FAB_D0_I3(RAM2FAB_D[26]),
	.Tile_X13Y11_RAM2FAB_D1_I0(RAM2FAB_D[25]),
	.Tile_X13Y11_RAM2FAB_D1_I1(RAM2FAB_D[24]),
	.Tile_X13Y11_RAM2FAB_D1_I2(dump[1]),
	.Tile_X13Y11_RAM2FAB_D1_I3(RAM2FAB_D[23]),
	.Tile_X13Y11_RAM2FAB_D2_I0(RAM2FAB_D[22]),
	.Tile_X13Y11_RAM2FAB_D2_I1(RAM2FAB_D[21]),
	.Tile_X13Y11_RAM2FAB_D2_I2(RAM2FAB_D[20]),
	.Tile_X13Y11_RAM2FAB_D2_I3(RAM2FAB_D[19]),
	.Tile_X13Y11_RAM2FAB_D3_I0(RAM2FAB_D[18]),
	.Tile_X13Y11_RAM2FAB_D3_I1(RAM2FAB_D[17]),
	.Tile_X13Y11_RAM2FAB_D3_I2(RAM2FAB_D[16]),
	.Tile_X13Y11_RAM2FAB_D3_I3(RAM2FAB_D[15]),
	.Tile_X13Y12_RAM2FAB_D0_I0(RAM2FAB_D[14]),
	.Tile_X13Y12_RAM2FAB_D0_I1(RAM2FAB_D[13]),
	.Tile_X13Y12_RAM2FAB_D0_I2(RAM2FAB_D[12]),
	.Tile_X13Y12_RAM2FAB_D0_I3(RAM2FAB_D[11]),
	.Tile_X13Y12_RAM2FAB_D1_I0(RAM2FAB_D[10]),
	.Tile_X13Y12_RAM2FAB_D1_I1(RAM2FAB_D[9]),
	.Tile_X13Y12_RAM2FAB_D1_I2(dump[0]),
	.Tile_X13Y12_RAM2FAB_D1_I3(RAM2FAB_D[8]),
	.Tile_X13Y12_RAM2FAB_D2_I0(RAM2FAB_D[7]),
	.Tile_X13Y12_RAM2FAB_D2_I1(RAM2FAB_D[6]),
	.Tile_X13Y12_RAM2FAB_D2_I2(RAM2FAB_D[5]),
	.Tile_X13Y12_RAM2FAB_D2_I3(RAM2FAB_D[4]),
	.Tile_X13Y12_RAM2FAB_D3_I0(RAM2FAB_D[3]),
	.Tile_X13Y12_RAM2FAB_D3_I1(RAM2FAB_D[2]),
	.Tile_X13Y12_RAM2FAB_D3_I2(RAM2FAB_D[1]),
	.Tile_X13Y12_RAM2FAB_D3_I3(RAM2FAB_D[0]),

	.Tile_X13Y1_FAB2RAM_D0_O0(FAB2RAM_D[191]),
	.Tile_X13Y1_FAB2RAM_D0_O1(FAB2RAM_D[190]),
	.Tile_X13Y1_FAB2RAM_D0_O2(FAB2RAM_D[189]),
	.Tile_X13Y1_FAB2RAM_D0_O3(FAB2RAM_D[188]),
	.Tile_X13Y1_FAB2RAM_D1_O0(FAB2RAM_D[187]),
	.Tile_X13Y1_FAB2RAM_D1_O1(FAB2RAM_D[186]),
	.Tile_X13Y1_FAB2RAM_D1_O2(FAB2RAM_D[185]),
	.Tile_X13Y1_FAB2RAM_D1_O3(FAB2RAM_D[184]),
	.Tile_X13Y1_FAB2RAM_D2_O0(FAB2RAM_D[183]),
	.Tile_X13Y1_FAB2RAM_D2_O1(FAB2RAM_D[182]),
	.Tile_X13Y1_FAB2RAM_D2_O2(FAB2RAM_D[181]),
	.Tile_X13Y1_FAB2RAM_D2_O3(FAB2RAM_D[180]),
	.Tile_X13Y1_FAB2RAM_D3_O0(FAB2RAM_D[179]),
	.Tile_X13Y1_FAB2RAM_D3_O1(FAB2RAM_D[178]),
	.Tile_X13Y1_FAB2RAM_D3_O2(FAB2RAM_D[177]),
	.Tile_X13Y1_FAB2RAM_D3_O3(FAB2RAM_D[176]),
	.Tile_X13Y2_FAB2RAM_D0_O0(FAB2RAM_D[175]),
	.Tile_X13Y2_FAB2RAM_D0_O1(FAB2RAM_D[174]),
	.Tile_X13Y2_FAB2RAM_D0_O2(FAB2RAM_D[173]),
	.Tile_X13Y2_FAB2RAM_D0_O3(FAB2RAM_D[172]),
	.Tile_X13Y2_FAB2RAM_D1_O0(FAB2RAM_D[171]),
	.Tile_X13Y2_FAB2RAM_D1_O1(FAB2RAM_D[170]),
	.Tile_X13Y2_FAB2RAM_D1_O2(FAB2RAM_D[169]),
	.Tile_X13Y2_FAB2RAM_D1_O3(FAB2RAM_D[168]),
	.Tile_X13Y2_FAB2RAM_D2_O0(FAB2RAM_D[167]),
	.Tile_X13Y2_FAB2RAM_D2_O1(FAB2RAM_D[166]),
	.Tile_X13Y2_FAB2RAM_D2_O2(FAB2RAM_D[165]),
	.Tile_X13Y2_FAB2RAM_D2_O3(FAB2RAM_D[164]),
	.Tile_X13Y2_FAB2RAM_D3_O0(FAB2RAM_D[163]),
	.Tile_X13Y2_FAB2RAM_D3_O1(FAB2RAM_D[162]),
	.Tile_X13Y2_FAB2RAM_D3_O2(FAB2RAM_D[161]),
	.Tile_X13Y2_FAB2RAM_D3_O3(FAB2RAM_D[160]),
	.Tile_X13Y3_FAB2RAM_D0_O0(FAB2RAM_D[159]),
	.Tile_X13Y3_FAB2RAM_D0_O1(FAB2RAM_D[158]),
	.Tile_X13Y3_FAB2RAM_D0_O2(FAB2RAM_D[157]),
	.Tile_X13Y3_FAB2RAM_D0_O3(FAB2RAM_D[156]),
	.Tile_X13Y3_FAB2RAM_D1_O0(FAB2RAM_D[155]),
	.Tile_X13Y3_FAB2RAM_D1_O1(FAB2RAM_D[154]),
	.Tile_X13Y3_FAB2RAM_D1_O2(FAB2RAM_D[153]),
	.Tile_X13Y3_FAB2RAM_D1_O3(FAB2RAM_D[152]),
	.Tile_X13Y3_FAB2RAM_D2_O0(FAB2RAM_D[151]),
	.Tile_X13Y3_FAB2RAM_D2_O1(FAB2RAM_D[150]),
	.Tile_X13Y3_FAB2RAM_D2_O2(FAB2RAM_D[149]),
	.Tile_X13Y3_FAB2RAM_D2_O3(FAB2RAM_D[148]),
	.Tile_X13Y3_FAB2RAM_D3_O0(FAB2RAM_D[147]),
	.Tile_X13Y3_FAB2RAM_D3_O1(FAB2RAM_D[146]),
	.Tile_X13Y3_FAB2RAM_D3_O2(FAB2RAM_D[145]),
	.Tile_X13Y3_FAB2RAM_D3_O3(FAB2RAM_D[144]),
	.Tile_X13Y4_FAB2RAM_D0_O0(FAB2RAM_D[143]),
	.Tile_X13Y4_FAB2RAM_D0_O1(FAB2RAM_D[142]),
	.Tile_X13Y4_FAB2RAM_D0_O2(FAB2RAM_D[141]),
	.Tile_X13Y4_FAB2RAM_D0_O3(FAB2RAM_D[140]),
	.Tile_X13Y4_FAB2RAM_D1_O0(FAB2RAM_D[139]),
	.Tile_X13Y4_FAB2RAM_D1_O1(FAB2RAM_D[138]),
	.Tile_X13Y4_FAB2RAM_D1_O2(FAB2RAM_D[137]),
	.Tile_X13Y4_FAB2RAM_D1_O3(FAB2RAM_D[136]),
	.Tile_X13Y4_FAB2RAM_D2_O0(FAB2RAM_D[135]),
	.Tile_X13Y4_FAB2RAM_D2_O1(FAB2RAM_D[134]),
	.Tile_X13Y4_FAB2RAM_D2_O2(FAB2RAM_D[133]),
	.Tile_X13Y4_FAB2RAM_D2_O3(FAB2RAM_D[132]),
	.Tile_X13Y4_FAB2RAM_D3_O0(FAB2RAM_D[131]),
	.Tile_X13Y4_FAB2RAM_D3_O1(FAB2RAM_D[130]),
	.Tile_X13Y4_FAB2RAM_D3_O2(FAB2RAM_D[129]),
	.Tile_X13Y4_FAB2RAM_D3_O3(FAB2RAM_D[128]),
	.Tile_X13Y5_FAB2RAM_D0_O0(FAB2RAM_D[127]),
	.Tile_X13Y5_FAB2RAM_D0_O1(FAB2RAM_D[126]),
	.Tile_X13Y5_FAB2RAM_D0_O2(FAB2RAM_D[125]),
	.Tile_X13Y5_FAB2RAM_D0_O3(FAB2RAM_D[124]),
	.Tile_X13Y5_FAB2RAM_D1_O0(FAB2RAM_D[123]),
	.Tile_X13Y5_FAB2RAM_D1_O1(FAB2RAM_D[122]),
	.Tile_X13Y5_FAB2RAM_D1_O2(FAB2RAM_D[121]),
	.Tile_X13Y5_FAB2RAM_D1_O3(FAB2RAM_D[120]),
	.Tile_X13Y5_FAB2RAM_D2_O0(FAB2RAM_D[119]),
	.Tile_X13Y5_FAB2RAM_D2_O1(FAB2RAM_D[118]),
	.Tile_X13Y5_FAB2RAM_D2_O2(FAB2RAM_D[117]),
	.Tile_X13Y5_FAB2RAM_D2_O3(FAB2RAM_D[116]),
	.Tile_X13Y5_FAB2RAM_D3_O0(FAB2RAM_D[115]),
	.Tile_X13Y5_FAB2RAM_D3_O1(FAB2RAM_D[114]),
	.Tile_X13Y5_FAB2RAM_D3_O2(FAB2RAM_D[113]),
	.Tile_X13Y5_FAB2RAM_D3_O3(FAB2RAM_D[112]),
	.Tile_X13Y6_FAB2RAM_D0_O0(FAB2RAM_D[111]),
	.Tile_X13Y6_FAB2RAM_D0_O1(FAB2RAM_D[110]),
	.Tile_X13Y6_FAB2RAM_D0_O2(FAB2RAM_D[109]),
	.Tile_X13Y6_FAB2RAM_D0_O3(FAB2RAM_D[108]),
	.Tile_X13Y6_FAB2RAM_D1_O0(FAB2RAM_D[107]),
	.Tile_X13Y6_FAB2RAM_D1_O1(FAB2RAM_D[106]),
	.Tile_X13Y6_FAB2RAM_D1_O2(FAB2RAM_D[105]),
	.Tile_X13Y6_FAB2RAM_D1_O3(FAB2RAM_D[104]),
	.Tile_X13Y6_FAB2RAM_D2_O0(FAB2RAM_D[103]),
	.Tile_X13Y6_FAB2RAM_D2_O1(FAB2RAM_D[102]),
	.Tile_X13Y6_FAB2RAM_D2_O2(FAB2RAM_D[101]),
	.Tile_X13Y6_FAB2RAM_D2_O3(FAB2RAM_D[100]),
	.Tile_X13Y6_FAB2RAM_D3_O0(FAB2RAM_D[99]),
	.Tile_X13Y6_FAB2RAM_D3_O1(FAB2RAM_D[98]),
	.Tile_X13Y6_FAB2RAM_D3_O2(FAB2RAM_D[97]),
	.Tile_X13Y6_FAB2RAM_D3_O3(FAB2RAM_D[96]),
	.Tile_X13Y7_FAB2RAM_D0_O0(FAB2RAM_D[95]),
	.Tile_X13Y7_FAB2RAM_D0_O1(FAB2RAM_D[94]),
	.Tile_X13Y7_FAB2RAM_D0_O2(FAB2RAM_D[93]),
	.Tile_X13Y7_FAB2RAM_D0_O3(FAB2RAM_D[92]),
	.Tile_X13Y7_FAB2RAM_D1_O0(FAB2RAM_D[91]),
	.Tile_X13Y7_FAB2RAM_D1_O1(FAB2RAM_D[90]),
	.Tile_X13Y7_FAB2RAM_D1_O2(FAB2RAM_D[89]),
	.Tile_X13Y7_FAB2RAM_D1_O3(FAB2RAM_D[88]),
	.Tile_X13Y7_FAB2RAM_D2_O0(FAB2RAM_D[87]),
	.Tile_X13Y7_FAB2RAM_D2_O1(FAB2RAM_D[86]),
	.Tile_X13Y7_FAB2RAM_D2_O2(FAB2RAM_D[85]),
	.Tile_X13Y7_FAB2RAM_D2_O3(FAB2RAM_D[84]),
	.Tile_X13Y7_FAB2RAM_D3_O0(FAB2RAM_D[83]),
	.Tile_X13Y7_FAB2RAM_D3_O1(FAB2RAM_D[82]),
	.Tile_X13Y7_FAB2RAM_D3_O2(FAB2RAM_D[81]),
	.Tile_X13Y7_FAB2RAM_D3_O3(FAB2RAM_D[80]),
	.Tile_X13Y8_FAB2RAM_D0_O0(FAB2RAM_D[79]),
	.Tile_X13Y8_FAB2RAM_D0_O1(FAB2RAM_D[78]),
	.Tile_X13Y8_FAB2RAM_D0_O2(FAB2RAM_D[77]),
	.Tile_X13Y8_FAB2RAM_D0_O3(FAB2RAM_D[76]),
	.Tile_X13Y8_FAB2RAM_D1_O0(FAB2RAM_D[75]),
	.Tile_X13Y8_FAB2RAM_D1_O1(FAB2RAM_D[74]),
	.Tile_X13Y8_FAB2RAM_D1_O2(FAB2RAM_D[73]),
	.Tile_X13Y8_FAB2RAM_D1_O3(FAB2RAM_D[72]),
	.Tile_X13Y8_FAB2RAM_D2_O0(FAB2RAM_D[71]),
	.Tile_X13Y8_FAB2RAM_D2_O1(FAB2RAM_D[70]),
	.Tile_X13Y8_FAB2RAM_D2_O2(FAB2RAM_D[69]),
	.Tile_X13Y8_FAB2RAM_D2_O3(FAB2RAM_D[68]),
	.Tile_X13Y8_FAB2RAM_D3_O0(FAB2RAM_D[67]),
	.Tile_X13Y8_FAB2RAM_D3_O1(FAB2RAM_D[66]),
	.Tile_X13Y8_FAB2RAM_D3_O2(FAB2RAM_D[65]),
	.Tile_X13Y8_FAB2RAM_D3_O3(FAB2RAM_D[64]),
	.Tile_X13Y9_FAB2RAM_D0_O0(FAB2RAM_D[63]),
	.Tile_X13Y9_FAB2RAM_D0_O1(FAB2RAM_D[62]),
	.Tile_X13Y9_FAB2RAM_D0_O2(FAB2RAM_D[61]),
	.Tile_X13Y9_FAB2RAM_D0_O3(FAB2RAM_D[60]),
	.Tile_X13Y9_FAB2RAM_D1_O0(FAB2RAM_D[59]),
	.Tile_X13Y9_FAB2RAM_D1_O1(FAB2RAM_D[58]),
	.Tile_X13Y9_FAB2RAM_D1_O2(FAB2RAM_D[57]),
	.Tile_X13Y9_FAB2RAM_D1_O3(FAB2RAM_D[56]),
	.Tile_X13Y9_FAB2RAM_D2_O0(FAB2RAM_D[55]),
	.Tile_X13Y9_FAB2RAM_D2_O1(FAB2RAM_D[54]),
	.Tile_X13Y9_FAB2RAM_D2_O2(FAB2RAM_D[53]),
	.Tile_X13Y9_FAB2RAM_D2_O3(FAB2RAM_D[52]),
	.Tile_X13Y9_FAB2RAM_D3_O0(FAB2RAM_D[51]),
	.Tile_X13Y9_FAB2RAM_D3_O1(FAB2RAM_D[50]),
	.Tile_X13Y9_FAB2RAM_D3_O2(FAB2RAM_D[49]),
	.Tile_X13Y9_FAB2RAM_D3_O3(FAB2RAM_D[48]),
	.Tile_X13Y10_FAB2RAM_D0_O0(FAB2RAM_D[47]),
	.Tile_X13Y10_FAB2RAM_D0_O1(FAB2RAM_D[46]),
	.Tile_X13Y10_FAB2RAM_D0_O2(FAB2RAM_D[45]),
	.Tile_X13Y10_FAB2RAM_D0_O3(FAB2RAM_D[44]),
	.Tile_X13Y10_FAB2RAM_D1_O0(FAB2RAM_D[43]),
	.Tile_X13Y10_FAB2RAM_D1_O1(FAB2RAM_D[42]),
	.Tile_X13Y10_FAB2RAM_D1_O2(FAB2RAM_D[41]),
	.Tile_X13Y10_FAB2RAM_D1_O3(FAB2RAM_D[40]),
	.Tile_X13Y10_FAB2RAM_D2_O0(FAB2RAM_D[39]),
	.Tile_X13Y10_FAB2RAM_D2_O1(FAB2RAM_D[38]),
	.Tile_X13Y10_FAB2RAM_D2_O2(FAB2RAM_D[37]),
	.Tile_X13Y10_FAB2RAM_D2_O3(FAB2RAM_D[36]),
	.Tile_X13Y10_FAB2RAM_D3_O0(FAB2RAM_D[35]),
	.Tile_X13Y10_FAB2RAM_D3_O1(FAB2RAM_D[34]),
	.Tile_X13Y10_FAB2RAM_D3_O2(FAB2RAM_D[33]),
	.Tile_X13Y10_FAB2RAM_D3_O3(FAB2RAM_D[32]),
	.Tile_X13Y11_FAB2RAM_D0_O0(FAB2RAM_D[31]),
	.Tile_X13Y11_FAB2RAM_D0_O1(FAB2RAM_D[30]),
	.Tile_X13Y11_FAB2RAM_D0_O2(FAB2RAM_D[29]),
	.Tile_X13Y11_FAB2RAM_D0_O3(FAB2RAM_D[28]),
	.Tile_X13Y11_FAB2RAM_D1_O0(FAB2RAM_D[27]),
	.Tile_X13Y11_FAB2RAM_D1_O1(FAB2RAM_D[26]),
	.Tile_X13Y11_FAB2RAM_D1_O2(FAB2RAM_D[25]),
	.Tile_X13Y11_FAB2RAM_D1_O3(FAB2RAM_D[24]),
	.Tile_X13Y11_FAB2RAM_D2_O0(FAB2RAM_D[23]),
	.Tile_X13Y11_FAB2RAM_D2_O1(FAB2RAM_D[22]),
	.Tile_X13Y11_FAB2RAM_D2_O2(FAB2RAM_D[21]),
	.Tile_X13Y11_FAB2RAM_D2_O3(FAB2RAM_D[20]),
	.Tile_X13Y11_FAB2RAM_D3_O0(FAB2RAM_D[19]),
	.Tile_X13Y11_FAB2RAM_D3_O1(FAB2RAM_D[18]),
	.Tile_X13Y11_FAB2RAM_D3_O2(FAB2RAM_D[17]),
	.Tile_X13Y11_FAB2RAM_D3_O3(FAB2RAM_D[16]),
	.Tile_X13Y12_FAB2RAM_D0_O0(FAB2RAM_D[15]),
	.Tile_X13Y12_FAB2RAM_D0_O1(FAB2RAM_D[14]),
	.Tile_X13Y12_FAB2RAM_D0_O2(FAB2RAM_D[13]),
	.Tile_X13Y12_FAB2RAM_D0_O3(FAB2RAM_D[12]),
	.Tile_X13Y12_FAB2RAM_D1_O0(FAB2RAM_D[11]),
	.Tile_X13Y12_FAB2RAM_D1_O1(FAB2RAM_D[10]),
	.Tile_X13Y12_FAB2RAM_D1_O2(FAB2RAM_D[9]),
	.Tile_X13Y12_FAB2RAM_D1_O3(FAB2RAM_D[8]),
	.Tile_X13Y12_FAB2RAM_D2_O0(FAB2RAM_D[7]),
	.Tile_X13Y12_FAB2RAM_D2_O1(FAB2RAM_D[6]),
	.Tile_X13Y12_FAB2RAM_D2_O2(FAB2RAM_D[5]),
	.Tile_X13Y12_FAB2RAM_D2_O3(FAB2RAM_D[4]),
	.Tile_X13Y12_FAB2RAM_D3_O0(FAB2RAM_D[3]),
	.Tile_X13Y12_FAB2RAM_D3_O1(FAB2RAM_D[2]),
	.Tile_X13Y12_FAB2RAM_D3_O2(FAB2RAM_D[1]),
	.Tile_X13Y12_FAB2RAM_D3_O3(FAB2RAM_D[0]),

	.Tile_X13Y1_FAB2RAM_A0_O0(FAB2RAM_A[95]),
	.Tile_X13Y1_FAB2RAM_A0_O1(FAB2RAM_A[94]),
	.Tile_X13Y1_FAB2RAM_A0_O2(FAB2RAM_A[93]),
	.Tile_X13Y1_FAB2RAM_A0_O3(FAB2RAM_A[92]),
	.Tile_X13Y1_FAB2RAM_A1_O0(FAB2RAM_A[91]),
	.Tile_X13Y1_FAB2RAM_A1_O1(FAB2RAM_A[90]),
	.Tile_X13Y1_FAB2RAM_A1_O2(FAB2RAM_A[89]),
	.Tile_X13Y1_FAB2RAM_A1_O3(FAB2RAM_A[88]),
	.Tile_X13Y2_FAB2RAM_A0_O0(FAB2RAM_A[87]),
	.Tile_X13Y2_FAB2RAM_A0_O1(FAB2RAM_A[86]),
	.Tile_X13Y2_FAB2RAM_A0_O2(FAB2RAM_A[85]),
	.Tile_X13Y2_FAB2RAM_A0_O3(FAB2RAM_A[84]),
	.Tile_X13Y2_FAB2RAM_A1_O0(FAB2RAM_A[83]),
	.Tile_X13Y2_FAB2RAM_A1_O1(FAB2RAM_A[82]),
	.Tile_X13Y2_FAB2RAM_A1_O2(FAB2RAM_A[81]),
	.Tile_X13Y2_FAB2RAM_A1_O3(FAB2RAM_A[80]),
	.Tile_X13Y3_FAB2RAM_A0_O0(FAB2RAM_A[79]),
	.Tile_X13Y3_FAB2RAM_A0_O1(FAB2RAM_A[78]),
	.Tile_X13Y3_FAB2RAM_A0_O2(FAB2RAM_A[77]),
	.Tile_X13Y3_FAB2RAM_A0_O3(FAB2RAM_A[76]),
	.Tile_X13Y3_FAB2RAM_A1_O0(FAB2RAM_A[75]),
	.Tile_X13Y3_FAB2RAM_A1_O1(FAB2RAM_A[74]),
	.Tile_X13Y3_FAB2RAM_A1_O2(FAB2RAM_A[73]),
	.Tile_X13Y3_FAB2RAM_A1_O3(FAB2RAM_A[72]),
	.Tile_X13Y4_FAB2RAM_A0_O0(FAB2RAM_A[71]),
	.Tile_X13Y4_FAB2RAM_A0_O1(FAB2RAM_A[70]),
	.Tile_X13Y4_FAB2RAM_A0_O2(FAB2RAM_A[69]),
	.Tile_X13Y4_FAB2RAM_A0_O3(FAB2RAM_A[68]),
	.Tile_X13Y4_FAB2RAM_A1_O0(FAB2RAM_A[67]),
	.Tile_X13Y4_FAB2RAM_A1_O1(FAB2RAM_A[66]),
	.Tile_X13Y4_FAB2RAM_A1_O2(FAB2RAM_A[65]),
	.Tile_X13Y4_FAB2RAM_A1_O3(FAB2RAM_A[64]),
	.Tile_X13Y5_FAB2RAM_A0_O0(FAB2RAM_A[63]),
	.Tile_X13Y5_FAB2RAM_A0_O1(FAB2RAM_A[62]),
	.Tile_X13Y5_FAB2RAM_A0_O2(FAB2RAM_A[61]),
	.Tile_X13Y5_FAB2RAM_A0_O3(FAB2RAM_A[60]),
	.Tile_X13Y5_FAB2RAM_A1_O0(FAB2RAM_A[59]),
	.Tile_X13Y5_FAB2RAM_A1_O1(FAB2RAM_A[58]),
	.Tile_X13Y5_FAB2RAM_A1_O2(FAB2RAM_A[57]),
	.Tile_X13Y5_FAB2RAM_A1_O3(FAB2RAM_A[56]),
	.Tile_X13Y6_FAB2RAM_A0_O0(FAB2RAM_A[55]),
	.Tile_X13Y6_FAB2RAM_A0_O1(FAB2RAM_A[54]),
	.Tile_X13Y6_FAB2RAM_A0_O2(FAB2RAM_A[53]),
	.Tile_X13Y6_FAB2RAM_A0_O3(FAB2RAM_A[52]),
	.Tile_X13Y6_FAB2RAM_A1_O0(FAB2RAM_A[51]),
	.Tile_X13Y6_FAB2RAM_A1_O1(FAB2RAM_A[50]),
	.Tile_X13Y6_FAB2RAM_A1_O2(FAB2RAM_A[49]),
	.Tile_X13Y6_FAB2RAM_A1_O3(FAB2RAM_A[48]),
	.Tile_X13Y7_FAB2RAM_A0_O0(FAB2RAM_A[47]),
	.Tile_X13Y7_FAB2RAM_A0_O1(FAB2RAM_A[46]),
	.Tile_X13Y7_FAB2RAM_A0_O2(FAB2RAM_A[45]),
	.Tile_X13Y7_FAB2RAM_A0_O3(FAB2RAM_A[44]),
	.Tile_X13Y7_FAB2RAM_A1_O0(FAB2RAM_A[43]),
	.Tile_X13Y7_FAB2RAM_A1_O1(FAB2RAM_A[42]),
	.Tile_X13Y7_FAB2RAM_A1_O2(FAB2RAM_A[41]),
	.Tile_X13Y7_FAB2RAM_A1_O3(FAB2RAM_A[40]),
	.Tile_X13Y8_FAB2RAM_A0_O0(FAB2RAM_A[39]),
	.Tile_X13Y8_FAB2RAM_A0_O1(FAB2RAM_A[38]),
	.Tile_X13Y8_FAB2RAM_A0_O2(FAB2RAM_A[37]),
	.Tile_X13Y8_FAB2RAM_A0_O3(FAB2RAM_A[36]),
	.Tile_X13Y8_FAB2RAM_A1_O0(FAB2RAM_A[35]),
	.Tile_X13Y8_FAB2RAM_A1_O1(FAB2RAM_A[34]),
	.Tile_X13Y8_FAB2RAM_A1_O2(FAB2RAM_A[33]),
	.Tile_X13Y8_FAB2RAM_A1_O3(FAB2RAM_A[32]),
	.Tile_X13Y9_FAB2RAM_A0_O0(FAB2RAM_A[31]),
	.Tile_X13Y9_FAB2RAM_A0_O1(FAB2RAM_A[30]),
	.Tile_X13Y9_FAB2RAM_A0_O2(FAB2RAM_A[29]),
	.Tile_X13Y9_FAB2RAM_A0_O3(FAB2RAM_A[28]),
	.Tile_X13Y9_FAB2RAM_A1_O0(FAB2RAM_A[27]),
	.Tile_X13Y9_FAB2RAM_A1_O1(FAB2RAM_A[26]),
	.Tile_X13Y9_FAB2RAM_A1_O2(FAB2RAM_A[25]),
	.Tile_X13Y9_FAB2RAM_A1_O3(FAB2RAM_A[24]),
	.Tile_X13Y10_FAB2RAM_A0_O0(FAB2RAM_A[23]),
	.Tile_X13Y10_FAB2RAM_A0_O1(FAB2RAM_A[22]),
	.Tile_X13Y10_FAB2RAM_A0_O2(FAB2RAM_A[21]),
	.Tile_X13Y10_FAB2RAM_A0_O3(FAB2RAM_A[20]),
	.Tile_X13Y10_FAB2RAM_A1_O0(FAB2RAM_A[19]),
	.Tile_X13Y10_FAB2RAM_A1_O1(FAB2RAM_A[18]),
	.Tile_X13Y10_FAB2RAM_A1_O2(FAB2RAM_A[17]),
	.Tile_X13Y10_FAB2RAM_A1_O3(FAB2RAM_A[16]),
	.Tile_X13Y11_FAB2RAM_A0_O0(FAB2RAM_A[15]),
	.Tile_X13Y11_FAB2RAM_A0_O1(FAB2RAM_A[14]),
	.Tile_X13Y11_FAB2RAM_A0_O2(FAB2RAM_A[13]),
	.Tile_X13Y11_FAB2RAM_A0_O3(FAB2RAM_A[12]),
	.Tile_X13Y11_FAB2RAM_A1_O0(FAB2RAM_A[11]),
	.Tile_X13Y11_FAB2RAM_A1_O1(FAB2RAM_A[10]),
	.Tile_X13Y11_FAB2RAM_A1_O2(FAB2RAM_A[9]),
	.Tile_X13Y11_FAB2RAM_A1_O3(FAB2RAM_A[8]),
	.Tile_X13Y12_FAB2RAM_A0_O0(FAB2RAM_A[7]),
	.Tile_X13Y12_FAB2RAM_A0_O1(FAB2RAM_A[6]),
	.Tile_X13Y12_FAB2RAM_A0_O2(FAB2RAM_A[5]),
	.Tile_X13Y12_FAB2RAM_A0_O3(FAB2RAM_A[4]),
	.Tile_X13Y12_FAB2RAM_A1_O0(FAB2RAM_A[3]),
	.Tile_X13Y12_FAB2RAM_A1_O1(FAB2RAM_A[2]),
	.Tile_X13Y12_FAB2RAM_A1_O2(FAB2RAM_A[1]),
	.Tile_X13Y12_FAB2RAM_A1_O3(FAB2RAM_A[0]),

	.Tile_X13Y1_FAB2RAM_C_O0(FAB2RAM_C[47]),
	.Tile_X13Y1_FAB2RAM_C_O1(FAB2RAM_C[46]),
	.Tile_X13Y1_FAB2RAM_C_O2(FAB2RAM_C[45]),
	.Tile_X13Y1_FAB2RAM_C_O3(FAB2RAM_C[44]),
	.Tile_X13Y2_FAB2RAM_C_O0(FAB2RAM_C[43]),
	.Tile_X13Y2_FAB2RAM_C_O1(FAB2RAM_C[42]),
	.Tile_X13Y2_FAB2RAM_C_O2(FAB2RAM_C[41]),
	.Tile_X13Y2_FAB2RAM_C_O3(FAB2RAM_C[40]),
	.Tile_X13Y3_FAB2RAM_C_O0(FAB2RAM_C[39]),
	.Tile_X13Y3_FAB2RAM_C_O1(FAB2RAM_C[38]),
	.Tile_X13Y3_FAB2RAM_C_O2(FAB2RAM_C[37]),
	.Tile_X13Y3_FAB2RAM_C_O3(FAB2RAM_C[36]),
	.Tile_X13Y4_FAB2RAM_C_O0(FAB2RAM_C[35]),
	.Tile_X13Y4_FAB2RAM_C_O1(FAB2RAM_C[34]),
	.Tile_X13Y4_FAB2RAM_C_O2(FAB2RAM_C[33]),
	.Tile_X13Y4_FAB2RAM_C_O3(FAB2RAM_C[32]),
	.Tile_X13Y5_FAB2RAM_C_O0(FAB2RAM_C[31]),
	.Tile_X13Y5_FAB2RAM_C_O1(FAB2RAM_C[30]),
	.Tile_X13Y5_FAB2RAM_C_O2(FAB2RAM_C[29]),
	.Tile_X13Y5_FAB2RAM_C_O3(FAB2RAM_C[28]),
	.Tile_X13Y6_FAB2RAM_C_O0(FAB2RAM_C[27]),
	.Tile_X13Y6_FAB2RAM_C_O1(FAB2RAM_C[26]),
	.Tile_X13Y6_FAB2RAM_C_O2(FAB2RAM_C[25]),
	.Tile_X13Y6_FAB2RAM_C_O3(FAB2RAM_C[24]),
	.Tile_X13Y7_FAB2RAM_C_O0(FAB2RAM_C[23]),
	.Tile_X13Y7_FAB2RAM_C_O1(FAB2RAM_C[22]),
	.Tile_X13Y7_FAB2RAM_C_O2(FAB2RAM_C[21]),
	.Tile_X13Y7_FAB2RAM_C_O3(FAB2RAM_C[20]),
	.Tile_X13Y8_FAB2RAM_C_O0(FAB2RAM_C[19]),
	.Tile_X13Y8_FAB2RAM_C_O1(FAB2RAM_C[18]),
	.Tile_X13Y8_FAB2RAM_C_O2(FAB2RAM_C[17]),
	.Tile_X13Y8_FAB2RAM_C_O3(FAB2RAM_C[16]),
	.Tile_X13Y9_FAB2RAM_C_O0(FAB2RAM_C[15]),
	.Tile_X13Y9_FAB2RAM_C_O1(FAB2RAM_C[14]),
	.Tile_X13Y9_FAB2RAM_C_O2(FAB2RAM_C[13]),
	.Tile_X13Y9_FAB2RAM_C_O3(FAB2RAM_C[12]),
	.Tile_X13Y10_FAB2RAM_C_O0(FAB2RAM_C[11]),
	.Tile_X13Y10_FAB2RAM_C_O1(FAB2RAM_C[10]),
	.Tile_X13Y10_FAB2RAM_C_O2(FAB2RAM_C[9]),
	.Tile_X13Y10_FAB2RAM_C_O3(FAB2RAM_C[8]),
	.Tile_X13Y11_FAB2RAM_C_O0(FAB2RAM_C[7]),
	.Tile_X13Y11_FAB2RAM_C_O1(FAB2RAM_C[6]),
	.Tile_X13Y11_FAB2RAM_C_O2(FAB2RAM_C[5]),
	.Tile_X13Y11_FAB2RAM_C_O3(FAB2RAM_C[4]),
	.Tile_X13Y12_FAB2RAM_C_O0(FAB2RAM_C[3]),
	.Tile_X13Y12_FAB2RAM_C_O1(FAB2RAM_C[2]),
	.Tile_X13Y12_FAB2RAM_C_O2(FAB2RAM_C[1]),
	.Tile_X13Y12_FAB2RAM_C_O3(FAB2RAM_C[0]),

	.Tile_X13Y1_Config_accessC_bit0(Config_accessC[47]),
	.Tile_X13Y1_Config_accessC_bit1(Config_accessC[46]),
	.Tile_X13Y1_Config_accessC_bit2(Config_accessC[45]),
	.Tile_X13Y1_Config_accessC_bit3(Config_accessC[44]),
	.Tile_X13Y2_Config_accessC_bit0(Config_accessC[43]),
	.Tile_X13Y2_Config_accessC_bit1(Config_accessC[42]),
	.Tile_X13Y2_Config_accessC_bit2(Config_accessC[41]),
	.Tile_X13Y2_Config_accessC_bit3(Config_accessC[40]),
	.Tile_X13Y3_Config_accessC_bit0(Config_accessC[39]),
	.Tile_X13Y3_Config_accessC_bit1(Config_accessC[38]),
	.Tile_X13Y3_Config_accessC_bit2(Config_accessC[37]),
	.Tile_X13Y3_Config_accessC_bit3(Config_accessC[36]),
	.Tile_X13Y4_Config_accessC_bit0(Config_accessC[35]),
	.Tile_X13Y4_Config_accessC_bit1(Config_accessC[34]),
	.Tile_X13Y4_Config_accessC_bit2(Config_accessC[33]),
	.Tile_X13Y4_Config_accessC_bit3(Config_accessC[32]),
	.Tile_X13Y5_Config_accessC_bit0(Config_accessC[31]),
	.Tile_X13Y5_Config_accessC_bit1(Config_accessC[30]),
	.Tile_X13Y5_Config_accessC_bit2(Config_accessC[29]),
	.Tile_X13Y5_Config_accessC_bit3(Config_accessC[28]),
	.Tile_X13Y6_Config_accessC_bit0(Config_accessC[27]),
	.Tile_X13Y6_Config_accessC_bit1(Config_accessC[26]),
	.Tile_X13Y6_Config_accessC_bit2(Config_accessC[25]),
	.Tile_X13Y6_Config_accessC_bit3(Config_accessC[24]),
	.Tile_X13Y7_Config_accessC_bit0(Config_accessC[23]),
	.Tile_X13Y7_Config_accessC_bit1(Config_accessC[22]),
	.Tile_X13Y7_Config_accessC_bit2(Config_accessC[21]),
	.Tile_X13Y7_Config_accessC_bit3(Config_accessC[20]),
	.Tile_X13Y8_Config_accessC_bit0(Config_accessC[19]),
	.Tile_X13Y8_Config_accessC_bit1(Config_accessC[18]),
	.Tile_X13Y8_Config_accessC_bit2(Config_accessC[17]),
	.Tile_X13Y8_Config_accessC_bit3(Config_accessC[16]),
	.Tile_X13Y9_Config_accessC_bit0(Config_accessC[15]),
	.Tile_X13Y9_Config_accessC_bit1(Config_accessC[14]),
	.Tile_X13Y9_Config_accessC_bit2(Config_accessC[13]),
	.Tile_X13Y9_Config_accessC_bit3(Config_accessC[12]),
	.Tile_X13Y10_Config_accessC_bit0(Config_accessC[11]),
	.Tile_X13Y10_Config_accessC_bit1(Config_accessC[10]),
	.Tile_X13Y10_Config_accessC_bit2(Config_accessC[9]),
	.Tile_X13Y10_Config_accessC_bit3(Config_accessC[8]),
	.Tile_X13Y11_Config_accessC_bit0(Config_accessC[7]),
	.Tile_X13Y11_Config_accessC_bit1(Config_accessC[6]),
	.Tile_X13Y11_Config_accessC_bit2(Config_accessC[5]),
	.Tile_X13Y11_Config_accessC_bit3(Config_accessC[4]),
	.Tile_X13Y12_Config_accessC_bit0(Config_accessC[3]),
	.Tile_X13Y12_Config_accessC_bit1(Config_accessC[2]),
	.Tile_X13Y12_Config_accessC_bit2(Config_accessC[1]),
	.Tile_X13Y12_Config_accessC_bit3(Config_accessC[0]),

	//declarations
	.UserCLK(CLK),
	.FrameData(FrameData),
	.FrameStrobe(FrameSelect)
	);

	BlockRAM_2KB Inst_BlockRAM_0 (
	.rd_clk(CLK),
	.rd_addr(FAB2RAM_A[10:0]),
	.rd_data(RAM2FAB_D[31:0]),
	.wr_clk(CLK),
	.wr_en(FAB2RAM_C[0]),
	.wr_addr(FAB2RAM_A[21:11]),
	.wr_data(FAB2RAM_D[31:0]),
	.C0(Config_accessC[0]),
	.C1(Config_accessC[1]),
	.C2(Config_accessC[2]),
	.C3(Config_accessC[3]),
	.C4(Config_accessC[4])
	);

	BlockRAM_2KB Inst_BlockRAM_1 (
	.rd_clk(CLK),
	.rd_addr(FAB2RAM_A[34:24]),
	.rd_data(RAM2FAB_D[79:48]),
	.wr_clk(CLK),
	.wr_en(FAB2RAM_C[12]),
	.wr_addr(FAB2RAM_A[45:35]),
	.wr_data(FAB2RAM_D[79:48]),
	.C0(Config_accessC[12]),
	.C1(Config_accessC[13]),
	.C2(Config_accessC[14]),
	.C3(Config_accessC[15]),
	.C4(Config_accessC[16])
	);

	BlockRAM_2KB Inst_BlockRAM_2 (
	.rd_clk(CLK),
	.rd_addr(FAB2RAM_A[58:48]),
	.rd_data(RAM2FAB_D[127:96]),
	.wr_clk(CLK),
	.wr_en(FAB2RAM_C[24]),
	.wr_addr(FAB2RAM_A[69:59]),
	.wr_data(FAB2RAM_D[127:96]),
	.C0(Config_accessC[24]),
	.C1(Config_accessC[25]),
	.C2(Config_accessC[26]),
	.C3(Config_accessC[27]),
	.C4(Config_accessC[28])
	);

	BlockRAM_2KB Inst_BlockRAM_3 (
	.rd_clk(CLK),
	.rd_addr(FAB2RAM_A[82:72]),
	.rd_data(RAM2FAB_D[175:144]),
	.wr_clk(CLK),
	.wr_en(FAB2RAM_C[36]),
	.wr_addr(FAB2RAM_A[93:83]),
	.wr_data(FAB2RAM_D[175:144]),
	.C0(Config_accessC[36]),
	.C1(Config_accessC[37]),
	.C2(Config_accessC[38]),
	.C3(Config_accessC[39]),
	.C4(Config_accessC[40])
	);

	assign FrameData = {32'h12345678,FrameRegister,32'h12345678};

endmodule

