magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 122
rect 285 0 288 122
<< via1 >>
rect 3 0 285 122
<< metal2 >>
rect 0 0 3 122
rect 285 0 288 122
<< properties >>
string GDS_END 88153612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88151176
<< end >>
